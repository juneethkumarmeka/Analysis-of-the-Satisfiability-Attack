module basic_2500_25000_3000_8_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_1533,In_195);
and U1 (N_1,In_219,In_1936);
nor U2 (N_2,In_718,In_589);
nor U3 (N_3,In_999,In_1415);
nand U4 (N_4,In_507,In_1485);
and U5 (N_5,In_248,In_391);
or U6 (N_6,In_1978,In_2391);
nand U7 (N_7,In_828,In_1159);
and U8 (N_8,In_1905,In_124);
nor U9 (N_9,In_1557,In_852);
nand U10 (N_10,In_111,In_809);
or U11 (N_11,In_1002,In_2366);
or U12 (N_12,In_1968,In_657);
nor U13 (N_13,In_1755,In_2053);
or U14 (N_14,In_1898,In_2140);
nor U15 (N_15,In_2193,In_155);
nand U16 (N_16,In_1388,In_1665);
xor U17 (N_17,In_1961,In_636);
nand U18 (N_18,In_1039,In_5);
or U19 (N_19,In_1028,In_868);
xnor U20 (N_20,In_821,In_632);
and U21 (N_21,In_2388,In_453);
or U22 (N_22,In_487,In_2418);
xor U23 (N_23,In_1561,In_922);
or U24 (N_24,In_1814,In_2258);
and U25 (N_25,In_479,In_932);
nand U26 (N_26,In_1107,In_1053);
nand U27 (N_27,In_186,In_2412);
and U28 (N_28,In_2332,In_1193);
nor U29 (N_29,In_1863,In_1141);
or U30 (N_30,In_28,In_1307);
nand U31 (N_31,In_713,In_936);
nor U32 (N_32,In_2044,In_1651);
or U33 (N_33,In_2325,In_1095);
and U34 (N_34,In_247,In_796);
and U35 (N_35,In_2381,In_2077);
nor U36 (N_36,In_1985,In_2274);
and U37 (N_37,In_2459,In_388);
nor U38 (N_38,In_2447,In_1687);
and U39 (N_39,In_593,In_798);
nand U40 (N_40,In_496,In_559);
or U41 (N_41,In_2179,In_1883);
and U42 (N_42,In_409,In_1316);
and U43 (N_43,In_849,In_2370);
nor U44 (N_44,In_1330,In_1829);
nor U45 (N_45,In_482,In_2331);
nor U46 (N_46,In_728,In_333);
nand U47 (N_47,In_164,In_1369);
nor U48 (N_48,In_1737,In_1641);
and U49 (N_49,In_2365,In_1270);
or U50 (N_50,In_2008,In_1045);
xnor U51 (N_51,In_710,In_1527);
xnor U52 (N_52,In_2334,In_1373);
xor U53 (N_53,In_1643,In_2143);
nand U54 (N_54,In_624,In_822);
and U55 (N_55,In_2424,In_1387);
nand U56 (N_56,In_1713,In_696);
nor U57 (N_57,In_781,In_446);
nand U58 (N_58,In_677,In_1627);
or U59 (N_59,In_855,In_907);
nor U60 (N_60,In_178,In_1171);
or U61 (N_61,In_64,In_2011);
xor U62 (N_62,In_1066,In_2453);
nand U63 (N_63,In_1470,In_1337);
and U64 (N_64,In_586,In_1495);
xor U65 (N_65,In_344,In_990);
nand U66 (N_66,In_580,In_38);
nand U67 (N_67,In_658,In_1513);
or U68 (N_68,In_1418,In_2121);
or U69 (N_69,In_764,In_403);
nand U70 (N_70,In_293,In_1626);
or U71 (N_71,In_628,In_91);
nor U72 (N_72,In_1758,In_635);
nand U73 (N_73,In_1433,In_2451);
nand U74 (N_74,In_1482,In_1069);
and U75 (N_75,In_913,In_70);
and U76 (N_76,In_996,In_1283);
nor U77 (N_77,In_1220,In_993);
and U78 (N_78,In_2180,In_1182);
or U79 (N_79,In_935,In_714);
nor U80 (N_80,In_704,In_158);
or U81 (N_81,In_90,In_1531);
and U82 (N_82,In_1299,In_1413);
nor U83 (N_83,In_2488,In_399);
nor U84 (N_84,In_241,In_1902);
nor U85 (N_85,In_323,In_39);
and U86 (N_86,In_199,In_2495);
nor U87 (N_87,In_524,In_2378);
or U88 (N_88,In_2050,In_221);
nor U89 (N_89,In_641,In_638);
xnor U90 (N_90,In_1650,In_401);
nor U91 (N_91,In_1734,In_674);
nand U92 (N_92,In_1680,In_23);
nor U93 (N_93,In_663,In_2435);
or U94 (N_94,In_1587,In_160);
xor U95 (N_95,In_450,In_502);
and U96 (N_96,In_168,In_891);
and U97 (N_97,In_1313,In_2368);
nor U98 (N_98,In_901,In_1279);
or U99 (N_99,In_1483,In_1952);
nand U100 (N_100,In_918,In_800);
nor U101 (N_101,In_1449,In_542);
and U102 (N_102,In_722,In_2494);
and U103 (N_103,In_1191,In_1026);
nor U104 (N_104,In_610,In_434);
and U105 (N_105,In_2014,In_1260);
nand U106 (N_106,In_1020,In_1402);
and U107 (N_107,In_2001,In_2146);
and U108 (N_108,In_625,In_816);
nor U109 (N_109,In_335,In_2300);
nand U110 (N_110,In_501,In_1659);
nor U111 (N_111,In_357,In_390);
nor U112 (N_112,In_1216,In_972);
and U113 (N_113,In_1731,In_2197);
nand U114 (N_114,In_861,In_940);
nor U115 (N_115,In_2278,In_379);
and U116 (N_116,In_1132,In_2081);
nor U117 (N_117,In_2428,In_1882);
nand U118 (N_118,In_1931,In_2027);
or U119 (N_119,In_1785,In_956);
or U120 (N_120,In_371,In_698);
or U121 (N_121,In_2246,In_430);
nor U122 (N_122,In_1027,In_1808);
and U123 (N_123,In_1516,In_252);
nand U124 (N_124,In_1981,In_1743);
nor U125 (N_125,In_418,In_157);
and U126 (N_126,In_2042,In_95);
or U127 (N_127,In_2188,In_777);
nand U128 (N_128,In_1078,In_1001);
nor U129 (N_129,In_2189,In_1560);
or U130 (N_130,In_108,In_1632);
xor U131 (N_131,In_1621,In_2088);
or U132 (N_132,In_601,In_544);
nand U133 (N_133,In_2000,In_2323);
nand U134 (N_134,In_2203,In_1572);
and U135 (N_135,In_135,In_460);
xor U136 (N_136,In_2032,In_533);
nand U137 (N_137,In_1768,In_2313);
nor U138 (N_138,In_1872,In_412);
xnor U139 (N_139,In_1007,In_1293);
nor U140 (N_140,In_1221,In_1897);
or U141 (N_141,In_385,In_961);
or U142 (N_142,In_2136,In_1528);
and U143 (N_143,In_170,In_311);
nor U144 (N_144,In_2449,In_2497);
or U145 (N_145,In_1727,In_517);
and U146 (N_146,In_753,In_2327);
xnor U147 (N_147,In_1416,In_948);
nor U148 (N_148,In_1467,In_448);
and U149 (N_149,In_1615,In_2359);
and U150 (N_150,In_1630,In_963);
nor U151 (N_151,In_1033,In_975);
xor U152 (N_152,In_1946,In_2306);
and U153 (N_153,In_1878,In_1228);
or U154 (N_154,In_1181,In_1784);
nor U155 (N_155,In_969,In_60);
or U156 (N_156,In_4,In_202);
and U157 (N_157,In_668,In_2322);
or U158 (N_158,In_478,In_667);
nand U159 (N_159,In_1261,In_237);
and U160 (N_160,In_2466,In_1035);
and U161 (N_161,In_953,In_1044);
or U162 (N_162,In_2375,In_1376);
and U163 (N_163,In_691,In_1301);
nand U164 (N_164,In_86,In_1851);
nand U165 (N_165,In_1813,In_1894);
nor U166 (N_166,In_122,In_1018);
and U167 (N_167,In_1631,In_58);
or U168 (N_168,In_84,In_2054);
xor U169 (N_169,In_1083,In_461);
or U170 (N_170,In_943,In_1236);
nor U171 (N_171,In_1274,In_1438);
or U172 (N_172,In_1804,In_1569);
nand U173 (N_173,In_2031,In_772);
and U174 (N_174,In_1363,In_1917);
nor U175 (N_175,In_459,In_2217);
nor U176 (N_176,In_686,In_1606);
or U177 (N_177,In_1267,In_620);
nand U178 (N_178,In_730,In_2083);
or U179 (N_179,In_1389,In_350);
or U180 (N_180,In_511,In_766);
and U181 (N_181,In_181,In_1396);
nand U182 (N_182,In_795,In_2160);
nor U183 (N_183,In_2299,In_264);
nand U184 (N_184,In_504,In_1541);
or U185 (N_185,In_1195,In_48);
and U186 (N_186,In_910,In_1318);
and U187 (N_187,In_1282,In_2478);
nand U188 (N_188,In_228,In_373);
and U189 (N_189,In_1778,In_1545);
nor U190 (N_190,In_213,In_1789);
or U191 (N_191,In_49,In_2177);
nor U192 (N_192,In_1967,In_272);
nand U193 (N_193,In_1,In_176);
or U194 (N_194,In_1328,In_314);
nor U195 (N_195,In_1099,In_805);
and U196 (N_196,In_532,In_204);
nand U197 (N_197,In_729,In_1435);
and U198 (N_198,In_1984,In_1234);
xnor U199 (N_199,In_2085,In_1303);
nor U200 (N_200,In_267,In_1353);
and U201 (N_201,In_640,In_185);
nor U202 (N_202,In_1745,In_1792);
and U203 (N_203,In_2404,In_2319);
nand U204 (N_204,In_1423,In_1884);
nor U205 (N_205,In_683,In_2123);
nand U206 (N_206,In_1716,In_527);
and U207 (N_207,In_365,In_1311);
or U208 (N_208,In_2390,In_1788);
or U209 (N_209,In_1060,In_484);
xor U210 (N_210,In_1497,In_1252);
or U211 (N_211,In_872,In_397);
nand U212 (N_212,In_361,In_1079);
nor U213 (N_213,In_2150,In_94);
or U214 (N_214,In_1317,In_1243);
or U215 (N_215,In_1006,In_147);
nand U216 (N_216,In_454,In_682);
and U217 (N_217,In_1447,In_2457);
or U218 (N_218,In_1886,In_472);
or U219 (N_219,In_747,In_2096);
nor U220 (N_220,In_950,In_1793);
and U221 (N_221,In_232,In_1380);
xor U222 (N_222,In_804,In_2316);
or U223 (N_223,In_2154,In_467);
and U224 (N_224,In_456,In_436);
nor U225 (N_225,In_678,In_2012);
nor U226 (N_226,In_782,In_1178);
nor U227 (N_227,In_1479,In_1455);
xnor U228 (N_228,In_1584,In_914);
or U229 (N_229,In_286,In_2392);
nand U230 (N_230,In_2344,In_1964);
or U231 (N_231,In_2089,In_848);
or U232 (N_232,In_196,In_191);
and U233 (N_233,In_885,In_2496);
nor U234 (N_234,In_2164,In_672);
and U235 (N_235,In_1896,In_964);
or U236 (N_236,In_905,In_1583);
nor U237 (N_237,In_949,In_194);
nor U238 (N_238,In_2196,In_536);
or U239 (N_239,In_2341,In_223);
and U240 (N_240,In_540,In_1932);
nand U241 (N_241,In_761,In_47);
nor U242 (N_242,In_954,In_1692);
and U243 (N_243,In_1055,In_316);
and U244 (N_244,In_226,In_1971);
xnor U245 (N_245,In_8,In_2234);
xor U246 (N_246,In_1566,In_1408);
nand U247 (N_247,In_421,In_701);
nand U248 (N_248,In_1766,In_419);
nor U249 (N_249,In_992,In_2290);
nor U250 (N_250,In_606,In_818);
or U251 (N_251,In_616,In_653);
xnor U252 (N_252,In_2132,In_1104);
nor U253 (N_253,In_1573,In_2200);
and U254 (N_254,In_2367,In_1577);
and U255 (N_255,In_132,In_2460);
and U256 (N_256,In_1254,In_1070);
and U257 (N_257,In_1288,In_346);
nand U258 (N_258,In_239,In_244);
and U259 (N_259,In_1726,In_1771);
nand U260 (N_260,In_1865,In_2315);
and U261 (N_261,In_1364,In_1982);
nand U262 (N_262,In_2294,In_2099);
xor U263 (N_263,In_1595,In_1400);
nand U264 (N_264,In_836,In_1063);
and U265 (N_265,In_133,In_1124);
and U266 (N_266,In_880,In_1036);
or U267 (N_267,In_1204,In_2280);
or U268 (N_268,In_493,In_1544);
and U269 (N_269,In_1300,In_50);
and U270 (N_270,In_945,In_285);
nand U271 (N_271,In_2402,In_508);
and U272 (N_272,In_1724,In_97);
nor U273 (N_273,In_908,In_930);
or U274 (N_274,In_1853,In_2417);
xor U275 (N_275,In_1277,In_1492);
or U276 (N_276,In_767,In_1258);
or U277 (N_277,In_291,In_19);
or U278 (N_278,In_1197,In_2006);
nand U279 (N_279,In_2307,In_2257);
nand U280 (N_280,In_2144,In_2041);
nand U281 (N_281,In_916,In_2361);
or U282 (N_282,In_1014,In_612);
and U283 (N_283,In_680,In_1266);
and U284 (N_284,In_1707,In_1453);
nand U285 (N_285,In_2128,In_1564);
nand U286 (N_286,In_599,In_1576);
nor U287 (N_287,In_750,In_2218);
nor U288 (N_288,In_1515,In_2397);
and U289 (N_289,In_971,In_1892);
or U290 (N_290,In_358,In_1333);
xor U291 (N_291,In_684,In_1670);
nand U292 (N_292,In_2467,In_519);
and U293 (N_293,In_378,In_510);
and U294 (N_294,In_1845,In_1164);
nor U295 (N_295,In_627,In_442);
or U296 (N_296,In_1466,In_1226);
nor U297 (N_297,In_2318,In_895);
and U298 (N_298,In_1410,In_1673);
or U299 (N_299,In_2051,In_1163);
nand U300 (N_300,In_166,In_1401);
nor U301 (N_301,In_1996,In_1691);
nand U302 (N_302,In_400,In_2239);
and U303 (N_303,In_25,In_831);
or U304 (N_304,In_887,In_12);
xor U305 (N_305,In_2236,In_843);
or U306 (N_306,In_2036,In_1654);
nand U307 (N_307,In_1137,In_1944);
nor U308 (N_308,In_2183,In_919);
nand U309 (N_309,In_2285,In_1382);
and U310 (N_310,In_2022,In_2104);
nand U311 (N_311,In_2276,In_1695);
or U312 (N_312,In_671,In_554);
nor U313 (N_313,In_1888,In_925);
nor U314 (N_314,In_3,In_538);
nor U315 (N_315,In_1499,In_334);
nand U316 (N_316,In_2118,In_1098);
nand U317 (N_317,In_1432,In_1786);
nand U318 (N_318,In_1347,In_1925);
and U319 (N_319,In_1272,In_670);
and U320 (N_320,In_514,In_2463);
or U321 (N_321,In_2034,In_2176);
nor U322 (N_322,In_1686,In_2350);
xor U323 (N_323,In_471,In_380);
or U324 (N_324,In_1381,In_1222);
or U325 (N_325,In_1976,In_180);
or U326 (N_326,In_1550,In_2329);
nor U327 (N_327,In_1911,In_2263);
nand U328 (N_328,In_1218,In_1802);
and U329 (N_329,In_1180,In_1175);
xor U330 (N_330,In_1153,In_1965);
or U331 (N_331,In_2298,In_1822);
nand U332 (N_332,In_1304,In_1714);
and U333 (N_333,In_1502,In_1783);
nand U334 (N_334,In_1797,In_2374);
or U335 (N_335,In_1209,In_1145);
or U336 (N_336,In_1004,In_1478);
or U337 (N_337,In_1958,In_773);
nand U338 (N_338,In_277,In_1312);
or U339 (N_339,In_1648,In_317);
nor U340 (N_340,In_1231,In_2019);
or U341 (N_341,In_1238,In_740);
and U342 (N_342,In_1477,In_130);
or U343 (N_343,In_149,In_1796);
nor U344 (N_344,In_1585,In_2030);
xor U345 (N_345,In_309,In_741);
and U346 (N_346,In_322,In_690);
nor U347 (N_347,In_468,In_2066);
nor U348 (N_348,In_1975,In_477);
nor U349 (N_349,In_847,In_2283);
or U350 (N_350,In_475,In_812);
and U351 (N_351,In_2261,In_1223);
nor U352 (N_352,In_2312,In_569);
xnor U353 (N_353,In_1953,In_1712);
nor U354 (N_354,In_2288,In_1355);
nor U355 (N_355,In_1049,In_1919);
and U356 (N_356,In_1281,In_1828);
or U357 (N_357,In_1994,In_1235);
nand U358 (N_358,In_211,In_2486);
nor U359 (N_359,In_1161,In_1242);
and U360 (N_360,In_437,In_598);
nor U361 (N_361,In_1278,In_279);
nand U362 (N_362,In_1950,In_2065);
nand U363 (N_363,In_495,In_148);
and U364 (N_364,In_384,In_525);
or U365 (N_365,In_283,In_2208);
nor U366 (N_366,In_1407,In_318);
nand U367 (N_367,In_153,In_1653);
nand U368 (N_368,In_783,In_1885);
and U369 (N_369,In_937,In_1676);
nor U370 (N_370,In_832,In_1914);
nand U371 (N_371,In_96,In_159);
nor U372 (N_372,In_844,In_1273);
nor U373 (N_373,In_473,In_2221);
nor U374 (N_374,In_985,In_571);
or U375 (N_375,In_1546,In_152);
nand U376 (N_376,In_1203,In_441);
xnor U377 (N_377,In_1463,In_222);
and U378 (N_378,In_2335,In_1620);
and U379 (N_379,In_520,In_217);
and U380 (N_380,In_2147,In_1593);
nor U381 (N_381,In_1773,In_1361);
nor U382 (N_382,In_808,In_2450);
or U383 (N_383,In_2337,In_699);
and U384 (N_384,In_794,In_934);
xor U385 (N_385,In_575,In_63);
and U386 (N_386,In_1397,In_2352);
or U387 (N_387,In_1761,In_1979);
nand U388 (N_388,In_360,In_476);
or U389 (N_389,In_1215,In_1841);
and U390 (N_390,In_1563,In_1484);
nand U391 (N_391,In_2343,In_1118);
or U392 (N_392,In_2267,In_888);
or U393 (N_393,In_853,In_2068);
nor U394 (N_394,In_235,In_1875);
and U395 (N_395,In_803,In_1781);
or U396 (N_396,In_899,In_2170);
nor U397 (N_397,In_1915,In_1062);
and U398 (N_398,In_1704,In_970);
nor U399 (N_399,In_1559,In_1824);
nor U400 (N_400,In_2046,In_2191);
or U401 (N_401,In_765,In_406);
or U402 (N_402,In_2481,In_80);
nor U403 (N_403,In_1777,In_1420);
nand U404 (N_404,In_208,In_2371);
and U405 (N_405,In_271,In_1729);
nor U406 (N_406,In_1846,In_1443);
nor U407 (N_407,In_2410,In_1454);
and U408 (N_408,In_1139,In_1959);
or U409 (N_409,In_428,In_744);
nand U410 (N_410,In_1790,In_838);
nand U411 (N_411,In_1100,In_2268);
or U412 (N_412,In_2358,In_1217);
or U413 (N_413,In_2023,In_743);
nor U414 (N_414,In_2145,In_1618);
nand U415 (N_415,In_187,In_1876);
nor U416 (N_416,In_1068,In_425);
xor U417 (N_417,In_2364,In_581);
nand U418 (N_418,In_1444,In_107);
and U419 (N_419,In_1094,In_1090);
or U420 (N_420,In_561,In_1310);
nand U421 (N_421,In_611,In_2212);
nor U422 (N_422,In_303,In_1377);
or U423 (N_423,In_329,In_2106);
nor U424 (N_424,In_2259,In_862);
nor U425 (N_425,In_112,In_1605);
nor U426 (N_426,In_123,In_2029);
nand U427 (N_427,In_1057,In_1506);
nor U428 (N_428,In_1963,In_912);
and U429 (N_429,In_1920,In_1294);
nor U430 (N_430,In_555,In_1728);
xnor U431 (N_431,In_1929,In_359);
nor U432 (N_432,In_509,In_320);
and U433 (N_433,In_1772,In_2185);
nor U434 (N_434,In_917,In_529);
nor U435 (N_435,In_464,In_75);
nand U436 (N_436,In_2204,In_2305);
or U437 (N_437,In_617,In_1344);
and U438 (N_438,In_1900,In_2195);
or U439 (N_439,In_1947,In_2311);
nor U440 (N_440,In_1669,In_583);
xor U441 (N_441,In_1746,In_52);
and U442 (N_442,In_2125,In_1085);
xnor U443 (N_443,In_579,In_404);
nand U444 (N_444,In_431,In_1750);
or U445 (N_445,In_339,In_1591);
nand U446 (N_446,In_1112,In_1023);
nor U447 (N_447,In_1038,In_382);
nand U448 (N_448,In_1534,In_1948);
and U449 (N_449,In_1103,In_2250);
nand U450 (N_450,In_763,In_42);
nor U451 (N_451,In_1855,In_1108);
and U452 (N_452,In_1526,In_29);
nor U453 (N_453,In_1297,In_2333);
or U454 (N_454,In_982,In_370);
nor U455 (N_455,In_522,In_2465);
and U456 (N_456,In_494,In_354);
nand U457 (N_457,In_1000,In_1548);
nor U458 (N_458,In_652,In_1690);
nor U459 (N_459,In_1080,In_2079);
nand U460 (N_460,In_325,In_1880);
nand U461 (N_461,In_881,In_659);
nor U462 (N_462,In_1903,In_2482);
nand U463 (N_463,In_2211,In_470);
or U464 (N_464,In_543,In_681);
nand U465 (N_465,In_405,In_2010);
or U466 (N_466,In_197,In_2168);
or U467 (N_467,In_1839,In_110);
nor U468 (N_468,In_845,In_1798);
or U469 (N_469,In_1398,In_364);
and U470 (N_470,In_1343,In_1858);
xor U471 (N_471,In_381,In_2171);
and U472 (N_472,In_1458,In_1956);
nand U473 (N_473,In_432,In_1165);
xnor U474 (N_474,In_989,In_1464);
nand U475 (N_475,In_88,In_1657);
or U476 (N_476,In_817,In_1156);
nand U477 (N_477,In_2296,In_238);
xnor U478 (N_478,In_2252,In_1417);
or U479 (N_479,In_2349,In_893);
nand U480 (N_480,In_1819,In_1030);
and U481 (N_481,In_732,In_2013);
nand U482 (N_482,In_1763,In_131);
or U483 (N_483,In_1491,In_1185);
or U484 (N_484,In_372,In_2394);
and U485 (N_485,In_1954,In_1120);
xor U486 (N_486,In_469,In_994);
or U487 (N_487,In_965,In_1024);
or U488 (N_488,In_1168,In_256);
nand U489 (N_489,In_491,In_1993);
and U490 (N_490,In_2105,In_860);
and U491 (N_491,In_1076,In_1543);
nand U492 (N_492,In_2187,In_1445);
and U493 (N_493,In_1940,In_41);
xor U494 (N_494,In_1757,In_20);
or U495 (N_495,In_54,In_79);
nand U496 (N_496,In_2039,In_2425);
or U497 (N_497,In_2468,In_1565);
nand U498 (N_498,In_1610,In_1612);
nor U499 (N_499,In_1157,In_2214);
and U500 (N_500,In_1206,In_1113);
and U501 (N_501,In_214,In_1805);
nand U502 (N_502,In_837,In_497);
or U503 (N_503,In_2162,In_2120);
nor U504 (N_504,In_1529,In_2438);
nor U505 (N_505,In_1422,In_646);
and U506 (N_506,In_161,In_2131);
and U507 (N_507,In_553,In_234);
and U508 (N_508,In_2336,In_2009);
nand U509 (N_509,In_900,In_1655);
nand U510 (N_510,In_305,In_1460);
or U511 (N_511,In_140,In_1741);
nand U512 (N_512,In_1607,In_1826);
nor U513 (N_513,In_423,In_1324);
or U514 (N_514,In_1162,In_859);
nor U515 (N_515,In_1342,In_902);
xor U516 (N_516,In_1166,In_121);
nor U517 (N_517,In_331,In_2255);
nand U518 (N_518,In_911,In_2427);
xnor U519 (N_519,In_2209,In_921);
or U520 (N_520,In_216,In_1096);
nand U521 (N_521,In_2277,In_2169);
nor U522 (N_522,In_1187,In_142);
or U523 (N_523,In_2225,In_18);
nand U524 (N_524,In_146,In_2219);
or U525 (N_525,In_2379,In_547);
nand U526 (N_526,In_814,In_1537);
nor U527 (N_527,In_2115,In_645);
nor U528 (N_528,In_560,In_1977);
and U529 (N_529,In_1472,In_1451);
xnor U530 (N_530,In_1015,In_731);
nand U531 (N_531,In_1174,In_190);
nor U532 (N_532,In_1640,In_2469);
or U533 (N_533,In_1322,In_2492);
nand U534 (N_534,In_2064,In_1290);
xnor U535 (N_535,In_257,In_1250);
xnor U536 (N_536,In_595,In_2385);
or U537 (N_537,In_462,In_503);
or U538 (N_538,In_506,In_537);
nor U539 (N_539,In_393,In_1708);
and U540 (N_540,In_693,In_505);
and U541 (N_541,In_2202,In_1280);
nand U542 (N_542,In_2498,In_661);
or U543 (N_543,In_929,In_1715);
and U544 (N_544,In_2279,In_2247);
or U545 (N_545,In_1151,In_723);
or U546 (N_546,In_1379,In_1683);
or U547 (N_547,In_1645,In_68);
or U548 (N_548,In_603,In_1291);
or U549 (N_549,In_719,In_1775);
nor U550 (N_550,In_414,In_1867);
nand U551 (N_551,In_138,In_2251);
and U552 (N_552,In_1469,In_251);
nor U553 (N_553,In_262,In_1521);
nand U554 (N_554,In_2439,In_778);
nor U555 (N_555,In_1625,In_2100);
nand U556 (N_556,In_1685,In_2080);
nor U557 (N_557,In_1922,In_631);
nor U558 (N_558,In_534,In_243);
and U559 (N_559,In_1081,In_2487);
and U560 (N_560,In_78,In_869);
nor U561 (N_561,In_76,In_1072);
nand U562 (N_562,In_550,In_2458);
and U563 (N_563,In_1341,In_2002);
xnor U564 (N_564,In_1633,In_163);
nor U565 (N_565,In_995,In_144);
xor U566 (N_566,In_1973,In_1092);
nor U567 (N_567,In_21,In_716);
nor U568 (N_568,In_266,In_1891);
or U569 (N_569,In_1701,In_830);
nand U570 (N_570,In_1667,In_101);
nand U571 (N_571,In_363,In_1893);
and U572 (N_572,In_1399,In_2192);
or U573 (N_573,In_134,In_2303);
and U574 (N_574,In_878,In_104);
and U575 (N_575,In_2297,In_1200);
or U576 (N_576,In_733,In_34);
nor U577 (N_577,In_1732,In_955);
nor U578 (N_578,In_1169,In_1320);
nor U579 (N_579,In_897,In_326);
or U580 (N_580,In_530,In_1762);
or U581 (N_581,In_633,In_345);
nor U582 (N_582,In_1285,In_7);
nor U583 (N_583,In_870,In_1934);
xor U584 (N_584,In_184,In_2491);
nor U585 (N_585,In_762,In_751);
nor U586 (N_586,In_725,In_2456);
and U587 (N_587,In_894,In_1866);
xnor U588 (N_588,In_1425,In_1663);
or U589 (N_589,In_957,In_236);
or U590 (N_590,In_819,In_2472);
and U591 (N_591,In_1998,In_1327);
nor U592 (N_592,In_207,In_11);
and U593 (N_593,In_877,In_1065);
nor U594 (N_594,In_2021,In_2007);
nor U595 (N_595,In_1111,In_2090);
and U596 (N_596,In_387,In_1144);
and U597 (N_597,In_1459,In_2224);
nor U598 (N_598,In_600,In_2153);
nand U599 (N_599,In_2320,In_1287);
nor U600 (N_600,In_2287,In_2493);
or U601 (N_601,In_136,In_556);
nand U602 (N_602,In_2440,In_874);
nand U603 (N_603,In_1214,In_1186);
nor U604 (N_604,In_892,In_656);
nor U605 (N_605,In_1452,In_2098);
nor U606 (N_606,In_366,In_1496);
nor U607 (N_607,In_1611,In_1589);
or U608 (N_608,In_879,In_647);
and U609 (N_609,In_398,In_1760);
nand U610 (N_610,In_1357,In_928);
nand U611 (N_611,In_1248,In_2207);
nor U612 (N_612,In_1597,In_596);
xnor U613 (N_613,In_974,In_790);
nor U614 (N_614,In_639,In_1602);
nand U615 (N_615,In_1158,In_1674);
and U616 (N_616,In_1152,In_2354);
nor U617 (N_617,In_1930,In_206);
nor U618 (N_618,In_1668,In_1329);
nor U619 (N_619,In_1879,In_1913);
and U620 (N_620,In_1562,In_623);
xor U621 (N_621,In_2351,In_2380);
or U622 (N_622,In_1769,In_1647);
and U623 (N_623,In_1599,In_1087);
nor U624 (N_624,In_71,In_987);
xnor U625 (N_625,In_1908,In_2243);
nor U626 (N_626,In_774,In_210);
or U627 (N_627,In_962,In_1512);
and U628 (N_628,In_1756,In_1918);
nand U629 (N_629,In_1747,In_1424);
or U630 (N_630,In_1061,In_2330);
nand U631 (N_631,In_977,In_951);
or U632 (N_632,In_174,In_127);
nand U633 (N_633,In_93,In_1753);
and U634 (N_634,In_2190,In_2420);
nor U635 (N_635,In_1490,In_2446);
and U636 (N_636,In_592,In_585);
nor U637 (N_637,In_1321,In_61);
nand U638 (N_638,In_53,In_1689);
nand U639 (N_639,In_1613,In_1859);
or U640 (N_640,In_1335,In_1409);
or U641 (N_641,In_634,In_906);
nor U642 (N_642,In_1532,In_1530);
nor U643 (N_643,In_643,In_1077);
nor U644 (N_644,In_2205,In_145);
or U645 (N_645,In_2223,In_2265);
or U646 (N_646,In_1489,In_1916);
nor U647 (N_647,In_780,In_702);
xnor U648 (N_648,In_1508,In_1703);
and U649 (N_649,In_1688,In_1056);
or U650 (N_650,In_1245,In_1847);
nor U651 (N_651,In_858,In_481);
or U652 (N_652,In_2338,In_1514);
nor U653 (N_653,In_1969,In_840);
nor U654 (N_654,In_2445,In_1336);
nor U655 (N_655,In_1907,In_1698);
nand U656 (N_656,In_1179,In_1538);
nand U657 (N_657,In_1849,In_260);
and U658 (N_658,In_169,In_1149);
xor U659 (N_659,In_2016,In_100);
nor U660 (N_660,In_205,In_2360);
and U661 (N_661,In_2119,In_1050);
or U662 (N_662,In_362,In_1127);
or U663 (N_663,In_2133,In_1807);
xnor U664 (N_664,In_712,In_1170);
nand U665 (N_665,In_1871,In_662);
xor U666 (N_666,In_2215,In_250);
xnor U667 (N_667,In_2238,In_1390);
nor U668 (N_668,In_535,In_1213);
and U669 (N_669,In_2199,In_2422);
and U670 (N_670,In_443,In_2406);
or U671 (N_671,In_2230,In_1962);
nor U672 (N_672,In_2093,In_545);
nor U673 (N_673,In_1553,In_1494);
nor U674 (N_674,In_630,In_2082);
xor U675 (N_675,In_2455,In_490);
nor U676 (N_676,In_2222,In_2063);
nor U677 (N_677,In_1933,In_394);
and U678 (N_678,In_754,In_2389);
nor U679 (N_679,In_2377,In_201);
or U680 (N_680,In_1468,In_1748);
nand U681 (N_681,In_1323,In_1522);
nand U682 (N_682,In_188,In_1440);
nand U683 (N_683,In_1910,In_1210);
nor U684 (N_684,In_1202,In_1131);
or U685 (N_685,In_810,In_1198);
or U686 (N_686,In_825,In_770);
xor U687 (N_687,In_410,In_1710);
nor U688 (N_688,In_1405,In_255);
or U689 (N_689,In_947,In_2231);
and U690 (N_690,In_1268,In_2087);
xor U691 (N_691,In_2292,In_2441);
nand U692 (N_692,In_474,In_629);
nor U693 (N_693,In_1012,In_2442);
and U694 (N_694,In_274,In_183);
or U695 (N_695,In_1115,In_597);
nor U696 (N_696,In_1086,In_444);
and U697 (N_697,In_1349,In_1385);
xor U698 (N_698,In_2092,In_621);
and U699 (N_699,In_1212,In_1598);
xor U700 (N_700,In_1619,In_1071);
or U701 (N_701,In_771,In_2175);
nor U702 (N_702,In_2461,In_1367);
xor U703 (N_703,In_1244,In_73);
nand U704 (N_704,In_2384,In_1121);
nand U705 (N_705,In_1816,In_1684);
or U706 (N_706,In_31,In_215);
nor U707 (N_707,In_489,In_227);
nand U708 (N_708,In_2241,In_2045);
xnor U709 (N_709,In_1264,In_62);
xor U710 (N_710,In_2067,In_1540);
or U711 (N_711,In_1624,In_198);
nor U712 (N_712,In_1992,In_1105);
or U713 (N_713,In_1302,In_15);
or U714 (N_714,In_1227,In_694);
nor U715 (N_715,In_1173,In_515);
nor U716 (N_716,In_141,In_952);
and U717 (N_717,In_1421,In_1374);
or U718 (N_718,In_2073,In_27);
nor U719 (N_719,In_1208,In_1836);
nand U720 (N_720,In_1147,In_2382);
nand U721 (N_721,In_1271,In_294);
nand U722 (N_722,In_465,In_1767);
nor U723 (N_723,In_2353,In_304);
and U724 (N_724,In_755,In_2226);
xor U725 (N_725,In_203,In_1500);
and U726 (N_726,In_2436,In_1835);
xnor U727 (N_727,In_313,In_1326);
or U728 (N_728,In_1251,In_116);
or U729 (N_729,In_499,In_1656);
nand U730 (N_730,In_841,In_336);
and U731 (N_731,In_2248,In_1989);
nand U732 (N_732,In_1465,In_775);
nand U733 (N_733,In_2097,In_1140);
or U734 (N_734,In_1661,In_1991);
xor U735 (N_735,In_319,In_1356);
xnor U736 (N_736,In_230,In_1097);
nand U737 (N_737,In_1308,In_1742);
or U738 (N_738,In_1412,In_851);
or U739 (N_739,In_67,In_1029);
or U740 (N_740,In_1869,In_785);
nor U741 (N_741,In_1549,In_1392);
xnor U742 (N_742,In_1838,In_1255);
or U743 (N_743,In_787,In_246);
and U744 (N_744,In_452,In_619);
xnor U745 (N_745,In_1276,In_1809);
nand U746 (N_746,In_968,In_2108);
nor U747 (N_747,In_449,In_991);
and U748 (N_748,In_376,In_1372);
nor U749 (N_749,In_1365,In_263);
nand U750 (N_750,In_2057,In_669);
and U751 (N_751,In_2172,In_2138);
and U752 (N_752,In_1779,In_1581);
or U753 (N_753,In_797,In_1675);
nor U754 (N_754,In_106,In_523);
nand U755 (N_755,In_2142,In_1176);
and U756 (N_756,In_875,In_1359);
nor U757 (N_757,In_613,In_59);
or U758 (N_758,In_776,In_1857);
or U759 (N_759,In_609,In_1046);
or U760 (N_760,In_480,In_967);
or U761 (N_761,In_389,In_1194);
nand U762 (N_762,In_429,In_1448);
or U763 (N_763,In_129,In_14);
or U764 (N_764,In_531,In_602);
and U765 (N_765,In_2048,In_439);
or U766 (N_766,In_167,In_2254);
and U767 (N_767,In_1555,In_752);
and U768 (N_768,In_2056,In_1517);
or U769 (N_769,In_269,In_1844);
xor U770 (N_770,In_1941,In_2273);
and U771 (N_771,In_119,In_162);
or U772 (N_772,In_1609,In_2431);
nand U773 (N_773,In_1629,In_1504);
nand U774 (N_774,In_463,In_2071);
or U775 (N_775,In_2373,In_1723);
nand U776 (N_776,In_551,In_2076);
nor U777 (N_777,In_1820,In_587);
nor U778 (N_778,In_1441,In_44);
nor U779 (N_779,In_518,In_253);
or U780 (N_780,In_1803,In_2163);
nor U781 (N_781,In_736,In_1325);
and U782 (N_782,In_1064,In_1601);
or U783 (N_783,In_1988,In_570);
nand U784 (N_784,In_150,In_1721);
and U785 (N_785,In_1172,In_426);
nand U786 (N_786,In_2095,In_815);
xor U787 (N_787,In_1129,In_607);
and U788 (N_788,In_1436,In_1309);
xnor U789 (N_789,In_1022,In_192);
and U790 (N_790,In_552,In_330);
nand U791 (N_791,In_2411,In_1350);
or U792 (N_792,In_618,In_1718);
nor U793 (N_793,In_2433,In_1945);
nand U794 (N_794,In_1133,In_2122);
nor U795 (N_795,In_2363,In_2237);
nor U796 (N_796,In_2286,In_1275);
nand U797 (N_797,In_128,In_2152);
nand U798 (N_798,In_541,In_676);
or U799 (N_799,In_1427,In_2139);
or U800 (N_800,In_2452,In_2489);
xnor U801 (N_801,In_0,In_1787);
nor U802 (N_802,In_769,In_1233);
nand U803 (N_803,In_2194,In_614);
nand U804 (N_804,In_1476,In_498);
and U805 (N_805,In_573,In_865);
or U806 (N_806,In_292,In_2471);
and U807 (N_807,In_2260,In_1776);
nor U808 (N_808,In_786,In_791);
and U809 (N_809,In_485,In_377);
and U810 (N_810,In_1265,In_175);
xnor U811 (N_811,In_2018,In_2072);
xnor U812 (N_812,In_1678,In_1256);
nor U813 (N_813,In_568,In_748);
nor U814 (N_814,In_402,In_2025);
or U815 (N_815,In_1935,In_546);
and U816 (N_816,In_424,In_1378);
xnor U817 (N_817,In_513,In_1642);
and U818 (N_818,In_165,In_2228);
nor U819 (N_819,In_1507,In_1800);
nand U820 (N_820,In_734,In_2432);
and U821 (N_821,In_2116,In_2091);
nor U822 (N_822,In_973,In_2281);
nor U823 (N_823,In_1224,In_2270);
or U824 (N_824,In_927,In_2284);
nand U825 (N_825,In_1138,In_2233);
or U826 (N_826,In_1031,In_1346);
xor U827 (N_827,In_720,In_2245);
nor U828 (N_828,In_289,In_1780);
and U829 (N_829,In_466,In_679);
xor U830 (N_830,In_310,In_2340);
nand U831 (N_831,In_2086,In_1697);
nor U832 (N_832,In_2107,In_259);
xor U833 (N_833,In_648,In_306);
nand U834 (N_834,In_811,In_1547);
nor U835 (N_835,In_2216,In_2117);
and U836 (N_836,In_1571,In_369);
nor U837 (N_837,In_1519,In_622);
nor U838 (N_838,In_1520,In_675);
nor U839 (N_839,In_1983,In_278);
and U840 (N_840,In_1295,In_1366);
nor U841 (N_841,In_2405,In_2301);
or U842 (N_842,In_1644,In_1493);
nand U843 (N_843,In_57,In_695);
nor U844 (N_844,In_321,In_1551);
and U845 (N_845,In_1128,In_209);
and U846 (N_846,In_451,In_938);
or U847 (N_847,In_1972,In_1906);
nand U848 (N_848,In_1338,In_2124);
or U849 (N_849,In_1815,In_1360);
or U850 (N_850,In_1759,In_26);
nand U851 (N_851,In_856,In_2109);
nor U852 (N_852,In_2186,In_959);
or U853 (N_853,In_1649,In_66);
and U854 (N_854,In_820,In_2362);
and U855 (N_855,In_1881,In_823);
nand U856 (N_856,In_1119,In_2302);
nand U857 (N_857,In_966,In_717);
and U858 (N_858,In_1262,In_1525);
nor U859 (N_859,In_1636,In_2272);
nand U860 (N_860,In_1475,In_341);
or U861 (N_861,In_1339,In_1025);
or U862 (N_862,In_1628,In_565);
and U863 (N_863,In_1662,In_1912);
nand U864 (N_864,In_1136,In_114);
nor U865 (N_865,In_2182,In_2414);
nand U866 (N_866,In_2304,In_280);
nor U867 (N_867,In_2314,In_528);
and U868 (N_868,In_367,In_1021);
nor U869 (N_869,In_2490,In_1205);
nor U870 (N_870,In_2137,In_2347);
nand U871 (N_871,In_2035,In_1837);
or U872 (N_872,In_37,In_1818);
and U873 (N_873,In_16,In_156);
nand U874 (N_874,In_1765,In_941);
or U875 (N_875,In_2477,In_1928);
or U876 (N_876,In_1117,In_1314);
nand U877 (N_877,In_1671,In_757);
nor U878 (N_878,In_408,In_1660);
and U879 (N_879,In_1146,In_2220);
nor U880 (N_880,In_229,In_1431);
or U881 (N_881,In_1511,In_154);
and U882 (N_882,In_1634,In_557);
nand U883 (N_883,In_1503,In_483);
nor U884 (N_884,In_526,In_2242);
nor U885 (N_885,In_1125,In_1830);
or U886 (N_886,In_1411,In_864);
or U887 (N_887,In_245,In_1319);
nand U888 (N_888,In_1130,In_768);
nor U889 (N_889,In_1637,In_997);
xor U890 (N_890,In_2156,In_558);
or U891 (N_891,In_113,In_1744);
nor U892 (N_892,In_1505,In_871);
xnor U893 (N_893,In_2229,In_2396);
nand U894 (N_894,In_758,In_1840);
nand U895 (N_895,In_2158,In_1143);
and U896 (N_896,In_958,In_1854);
nor U897 (N_897,In_1943,In_1150);
nand U898 (N_898,In_788,In_1658);
nor U899 (N_899,In_637,In_978);
nor U900 (N_900,In_883,In_700);
nor U901 (N_901,In_650,In_854);
nor U902 (N_902,In_2227,In_83);
and U903 (N_903,In_749,In_759);
or U904 (N_904,In_392,In_1823);
nand U905 (N_905,In_1340,In_890);
or U906 (N_906,In_539,In_413);
or U907 (N_907,In_1608,In_1375);
nand U908 (N_908,In_802,In_721);
or U909 (N_909,In_1498,In_193);
nand U910 (N_910,In_1801,In_857);
or U911 (N_911,In_1009,In_1730);
nand U912 (N_912,In_258,In_1600);
nand U913 (N_913,In_81,In_1048);
nor U914 (N_914,In_433,In_2094);
nor U915 (N_915,In_981,In_660);
and U916 (N_916,In_1101,In_98);
nand U917 (N_917,In_2293,In_298);
and U918 (N_918,In_886,In_2101);
xnor U919 (N_919,In_548,In_2159);
nor U920 (N_920,In_2112,In_846);
and U921 (N_921,In_1456,In_2102);
nand U922 (N_922,In_942,In_2157);
or U923 (N_923,In_976,In_931);
or U924 (N_924,In_1782,In_572);
or U925 (N_925,In_1588,In_2317);
or U926 (N_926,In_1554,In_2434);
and U927 (N_927,In_1462,In_2309);
and U928 (N_928,In_1568,In_301);
xor U929 (N_929,In_1201,In_1088);
and U930 (N_930,In_1966,In_2473);
or U931 (N_931,In_1093,In_1617);
or U932 (N_932,In_2024,In_850);
or U933 (N_933,In_177,In_1949);
nand U934 (N_934,In_417,In_1059);
nor U935 (N_935,In_1873,In_1395);
or U936 (N_936,In_1594,In_300);
xnor U937 (N_937,In_435,In_281);
nand U938 (N_938,In_2235,In_120);
nand U939 (N_939,In_566,In_2400);
nand U940 (N_940,In_1842,In_1923);
or U941 (N_941,In_1582,In_2005);
nor U942 (N_942,In_242,In_353);
nor U943 (N_943,In_447,In_608);
nor U944 (N_944,In_1990,In_139);
or U945 (N_945,In_1764,In_882);
nand U946 (N_946,In_2356,In_1123);
nor U947 (N_947,In_276,In_1177);
and U948 (N_948,In_1899,In_488);
and U949 (N_949,In_863,In_2348);
nor U950 (N_950,In_1740,In_1539);
nor U951 (N_951,In_2126,In_876);
nand U952 (N_952,In_1016,In_2416);
and U953 (N_953,In_1122,In_1799);
nor U954 (N_954,In_348,In_1895);
or U955 (N_955,In_2269,In_697);
nor U956 (N_956,In_1189,In_337);
nand U957 (N_957,In_1699,In_2475);
and U958 (N_958,In_903,In_2266);
nand U959 (N_959,In_1393,In_349);
or U960 (N_960,In_1754,In_807);
or U961 (N_961,In_2339,In_1230);
nor U962 (N_962,In_1269,In_254);
nand U963 (N_963,In_89,In_1909);
xnor U964 (N_964,In_2075,In_2372);
nand U965 (N_965,In_567,In_2443);
nand U966 (N_966,In_324,In_143);
nor U967 (N_967,In_1666,In_898);
or U968 (N_968,In_793,In_1586);
nor U969 (N_969,In_1446,In_563);
xnor U970 (N_970,In_486,In_1501);
or U971 (N_971,In_2069,In_2419);
nor U972 (N_972,In_82,In_826);
xor U973 (N_973,In_2244,In_1722);
or U974 (N_974,In_1480,In_915);
or U975 (N_975,In_1084,In_2357);
nand U976 (N_976,In_2184,In_1253);
and U977 (N_977,In_1827,In_760);
nor U978 (N_978,In_562,In_604);
or U979 (N_979,In_1904,In_909);
nor U980 (N_980,In_2017,In_1306);
or U981 (N_981,In_45,In_118);
nand U982 (N_982,In_2476,In_249);
and U983 (N_983,In_2326,In_1679);
and U984 (N_984,In_69,In_1239);
nor U985 (N_985,In_1524,In_2409);
xor U986 (N_986,In_1106,In_2401);
nand U987 (N_987,In_109,In_1148);
nand U988 (N_988,In_1974,In_2155);
nor U989 (N_989,In_705,In_584);
or U990 (N_990,In_1289,In_779);
or U991 (N_991,In_2423,In_200);
nor U992 (N_992,In_1623,In_979);
nor U993 (N_993,In_1510,In_1856);
and U994 (N_994,In_1705,In_1739);
or U995 (N_995,In_2355,In_1832);
or U996 (N_996,In_2129,In_1810);
nor U997 (N_997,In_654,In_1091);
and U998 (N_998,In_1134,In_1368);
xor U999 (N_999,In_1430,In_386);
nor U1000 (N_1000,In_1383,In_1032);
nand U1001 (N_1001,In_1575,In_2004);
nand U1002 (N_1002,In_2062,In_6);
nand U1003 (N_1003,In_218,In_1938);
nor U1004 (N_1004,In_2232,In_1019);
nor U1005 (N_1005,In_1700,In_2253);
nor U1006 (N_1006,In_792,In_687);
and U1007 (N_1007,In_2127,In_103);
nand U1008 (N_1008,In_2342,In_2070);
nand U1009 (N_1009,In_2149,In_2262);
nor U1010 (N_1010,In_2198,In_1074);
nand U1011 (N_1011,In_99,In_1237);
or U1012 (N_1012,In_1862,In_1394);
nand U1013 (N_1013,In_1719,In_72);
and U1014 (N_1014,In_784,In_923);
nand U1015 (N_1015,In_1384,In_1603);
xor U1016 (N_1016,In_2049,In_1155);
nor U1017 (N_1017,In_1457,In_87);
nor U1018 (N_1018,In_512,In_383);
nor U1019 (N_1019,In_1864,In_1008);
nor U1020 (N_1020,In_2020,In_1518);
and U1021 (N_1021,In_1725,In_2474);
nand U1022 (N_1022,In_1404,In_1037);
xor U1023 (N_1023,In_2321,In_302);
nand U1024 (N_1024,In_1752,In_835);
nand U1025 (N_1025,In_275,In_2399);
and U1026 (N_1026,In_1812,In_2178);
nor U1027 (N_1027,In_1184,In_1054);
nor U1028 (N_1028,In_17,In_742);
nor U1029 (N_1029,In_328,In_492);
or U1030 (N_1030,In_261,In_1939);
nand U1031 (N_1031,In_739,In_1580);
nor U1032 (N_1032,In_1980,In_43);
and U1033 (N_1033,In_1488,In_220);
or U1034 (N_1034,In_746,In_284);
nor U1035 (N_1035,In_240,In_2462);
nor U1036 (N_1036,In_1736,In_1870);
and U1037 (N_1037,In_2415,In_1075);
xor U1038 (N_1038,In_564,In_173);
or U1039 (N_1039,In_1694,In_1791);
or U1040 (N_1040,In_2408,In_1556);
nor U1041 (N_1041,In_1696,In_1806);
or U1042 (N_1042,In_1622,In_1471);
and U1043 (N_1043,In_2395,In_1414);
or U1044 (N_1044,In_2484,In_332);
or U1045 (N_1045,In_171,In_1817);
or U1046 (N_1046,In_2141,In_839);
nor U1047 (N_1047,In_273,In_1542);
and U1048 (N_1048,In_1334,In_1733);
nand U1049 (N_1049,In_2181,In_2103);
and U1050 (N_1050,In_1286,In_1860);
nand U1051 (N_1051,In_833,In_440);
xnor U1052 (N_1052,In_1219,In_2047);
nand U1053 (N_1053,In_1439,In_2289);
and U1054 (N_1054,In_873,In_2033);
or U1055 (N_1055,In_889,In_896);
or U1056 (N_1056,In_268,In_706);
xnor U1057 (N_1057,In_1955,In_2015);
and U1058 (N_1058,In_673,In_1051);
nor U1059 (N_1059,In_1473,In_2282);
or U1060 (N_1060,In_1795,In_2376);
nor U1061 (N_1061,In_342,In_1461);
or U1062 (N_1062,In_455,In_1042);
nor U1063 (N_1063,In_1257,In_1167);
xnor U1064 (N_1064,In_2055,In_1889);
or U1065 (N_1065,In_1646,In_2114);
and U1066 (N_1066,In_1190,In_352);
and U1067 (N_1067,In_1154,In_1639);
xnor U1068 (N_1068,In_1135,In_1614);
and U1069 (N_1069,In_1058,In_1196);
nand U1070 (N_1070,In_1142,In_1921);
nand U1071 (N_1071,In_2264,In_1850);
or U1072 (N_1072,In_834,In_1034);
nor U1073 (N_1073,In_225,In_827);
nand U1074 (N_1074,In_1284,In_986);
and U1075 (N_1075,In_2206,In_1579);
and U1076 (N_1076,In_40,In_2383);
or U1077 (N_1077,In_813,In_842);
nand U1078 (N_1078,In_35,In_1843);
and U1079 (N_1079,In_231,In_2037);
nand U1080 (N_1080,In_1887,In_1821);
xor U1081 (N_1081,In_172,In_1616);
nand U1082 (N_1082,In_1811,In_1354);
nand U1083 (N_1083,In_582,In_1749);
or U1084 (N_1084,In_1709,In_688);
or U1085 (N_1085,In_1315,In_1536);
nand U1086 (N_1086,In_117,In_65);
nand U1087 (N_1087,In_10,In_1774);
nand U1088 (N_1088,In_1578,In_709);
nor U1089 (N_1089,In_1693,In_287);
or U1090 (N_1090,In_2078,In_56);
nand U1091 (N_1091,In_2499,In_1706);
nand U1092 (N_1092,In_1677,In_1043);
nand U1093 (N_1093,In_1951,In_1635);
nand U1094 (N_1094,In_1751,In_295);
nand U1095 (N_1095,In_2061,In_1861);
nor U1096 (N_1096,In_924,In_137);
nor U1097 (N_1097,In_983,In_2201);
nand U1098 (N_1098,In_2346,In_806);
nand U1099 (N_1099,In_2295,In_591);
or U1100 (N_1100,In_422,In_368);
nor U1101 (N_1101,In_576,In_1852);
or U1102 (N_1102,In_396,In_1358);
nor U1103 (N_1103,In_1296,In_1010);
and U1104 (N_1104,In_2464,In_737);
and U1105 (N_1105,In_46,In_343);
xnor U1106 (N_1106,In_375,In_2166);
and U1107 (N_1107,In_420,In_1672);
and U1108 (N_1108,In_2369,In_1429);
nor U1109 (N_1109,In_1877,In_884);
nor U1110 (N_1110,In_1720,In_1292);
nand U1111 (N_1111,In_2398,In_233);
xor U1112 (N_1112,In_998,In_1552);
nor U1113 (N_1113,In_946,In_1428);
and U1114 (N_1114,In_74,In_307);
or U1115 (N_1115,In_212,In_1192);
xnor U1116 (N_1116,In_282,In_1109);
and U1117 (N_1117,In_1970,In_1702);
nor U1118 (N_1118,In_2060,In_1874);
nor U1119 (N_1119,In_2052,In_666);
nor U1120 (N_1120,In_1419,In_594);
nor U1121 (N_1121,In_988,In_2151);
nor U1122 (N_1122,In_726,In_1188);
and U1123 (N_1123,In_2483,In_445);
or U1124 (N_1124,In_2074,In_1834);
nand U1125 (N_1125,In_1211,In_1681);
nand U1126 (N_1126,In_2470,In_1073);
nand U1127 (N_1127,In_1362,In_1590);
and U1128 (N_1128,In_745,In_1082);
xor U1129 (N_1129,In_1570,In_2134);
nor U1130 (N_1130,In_799,In_1403);
or U1131 (N_1131,In_904,In_1199);
or U1132 (N_1132,In_655,In_1574);
nor U1133 (N_1133,In_1126,In_1298);
and U1134 (N_1134,In_1942,In_605);
and U1135 (N_1135,In_312,In_32);
nor U1136 (N_1136,In_642,In_2240);
and U1137 (N_1137,In_265,In_395);
nor U1138 (N_1138,In_427,In_411);
nand U1139 (N_1139,In_2386,In_1604);
nor U1140 (N_1140,In_126,In_1370);
nor U1141 (N_1141,In_1890,In_1426);
or U1142 (N_1142,In_1263,In_2393);
xnor U1143 (N_1143,In_33,In_13);
and U1144 (N_1144,In_1406,In_2043);
xnor U1145 (N_1145,In_980,In_1901);
and U1146 (N_1146,In_85,In_356);
or U1147 (N_1147,In_2110,In_1305);
nand U1148 (N_1148,In_867,In_2480);
and U1149 (N_1149,In_1246,In_1638);
or U1150 (N_1150,In_9,In_270);
and U1151 (N_1151,In_296,In_151);
or U1152 (N_1152,In_500,In_944);
nor U1153 (N_1153,In_703,In_2271);
or U1154 (N_1154,In_1831,In_1450);
nor U1155 (N_1155,In_1332,In_2421);
nor U1156 (N_1156,In_1437,In_1391);
nor U1157 (N_1157,In_125,In_738);
xor U1158 (N_1158,In_1926,In_1596);
or U1159 (N_1159,In_297,In_2413);
or U1160 (N_1160,In_1249,In_24);
and U1161 (N_1161,In_182,In_2059);
and U1162 (N_1162,In_574,In_2174);
xor U1163 (N_1163,In_926,In_2485);
or U1164 (N_1164,In_735,In_685);
nor U1165 (N_1165,In_2148,In_588);
nand U1166 (N_1166,In_2173,In_2275);
or U1167 (N_1167,In_2324,In_549);
nand U1168 (N_1168,In_939,In_1183);
nor U1169 (N_1169,In_457,In_829);
and U1170 (N_1170,In_1352,In_1937);
and U1171 (N_1171,In_1005,In_1535);
or U1172 (N_1172,In_340,In_2058);
nand U1173 (N_1173,In_36,In_689);
and U1174 (N_1174,In_1442,In_179);
nor U1175 (N_1175,In_105,In_1229);
nand U1176 (N_1176,In_2256,In_1997);
or U1177 (N_1177,In_2444,In_615);
nand U1178 (N_1178,In_2310,In_1110);
nand U1179 (N_1179,In_1848,In_438);
or U1180 (N_1180,In_1509,In_1351);
nand U1181 (N_1181,In_299,In_1474);
or U1182 (N_1182,In_1247,In_2430);
nor U1183 (N_1183,In_1664,In_1089);
and U1184 (N_1184,In_1434,In_1371);
nor U1185 (N_1185,In_2249,In_1999);
or U1186 (N_1186,In_590,In_1041);
xor U1187 (N_1187,In_2038,In_1011);
or U1188 (N_1188,In_1232,In_102);
and U1189 (N_1189,In_347,In_1348);
nand U1190 (N_1190,In_2426,In_1682);
nor U1191 (N_1191,In_1868,In_1995);
nor U1192 (N_1192,In_665,In_1957);
xnor U1193 (N_1193,In_189,In_727);
or U1194 (N_1194,In_1986,In_1770);
nand U1195 (N_1195,In_1738,In_2454);
xor U1196 (N_1196,In_2328,In_2387);
nand U1197 (N_1197,In_1592,In_1116);
nand U1198 (N_1198,In_1052,In_2448);
or U1199 (N_1199,In_2028,In_2167);
nor U1200 (N_1200,In_960,In_1486);
nand U1201 (N_1201,In_2161,In_789);
nor U1202 (N_1202,In_577,In_374);
and U1203 (N_1203,In_2437,In_1345);
and U1204 (N_1204,In_626,In_724);
and U1205 (N_1205,In_290,In_664);
and U1206 (N_1206,In_1114,In_416);
nand U1207 (N_1207,In_30,In_458);
or U1208 (N_1208,In_715,In_692);
nor U1209 (N_1209,In_2213,In_2130);
nor U1210 (N_1210,In_1102,In_2040);
nand U1211 (N_1211,In_1003,In_415);
nor U1212 (N_1212,In_1735,In_1481);
and U1213 (N_1213,In_327,In_866);
xor U1214 (N_1214,In_2111,In_1067);
and U1215 (N_1215,In_920,In_2429);
nand U1216 (N_1216,In_2165,In_711);
and U1217 (N_1217,In_1567,In_338);
and U1218 (N_1218,In_1259,In_115);
nand U1219 (N_1219,In_1240,In_2407);
nand U1220 (N_1220,In_1487,In_1960);
or U1221 (N_1221,In_2308,In_1225);
and U1222 (N_1222,In_1717,In_1794);
or U1223 (N_1223,In_1987,In_2);
nand U1224 (N_1224,In_2113,In_224);
or U1225 (N_1225,In_1927,In_1017);
and U1226 (N_1226,In_1386,In_824);
and U1227 (N_1227,In_1711,In_22);
nand U1228 (N_1228,In_51,In_644);
or U1229 (N_1229,In_2345,In_1652);
nand U1230 (N_1230,In_578,In_1825);
xor U1231 (N_1231,In_651,In_77);
nand U1232 (N_1232,In_1331,In_2084);
nand U1233 (N_1233,In_521,In_355);
nand U1234 (N_1234,In_1040,In_1523);
nor U1235 (N_1235,In_2135,In_2026);
or U1236 (N_1236,In_801,In_707);
or U1237 (N_1237,In_516,In_1207);
nand U1238 (N_1238,In_351,In_2210);
xor U1239 (N_1239,In_1833,In_288);
nor U1240 (N_1240,In_649,In_2403);
nand U1241 (N_1241,In_308,In_2291);
nor U1242 (N_1242,In_1013,In_2003);
nor U1243 (N_1243,In_92,In_984);
nor U1244 (N_1244,In_407,In_933);
nand U1245 (N_1245,In_1924,In_1047);
nor U1246 (N_1246,In_315,In_55);
or U1247 (N_1247,In_1241,In_2479);
nand U1248 (N_1248,In_1160,In_756);
and U1249 (N_1249,In_708,In_1558);
or U1250 (N_1250,In_318,In_1657);
nand U1251 (N_1251,In_2259,In_2475);
or U1252 (N_1252,In_825,In_2005);
nor U1253 (N_1253,In_1741,In_2259);
and U1254 (N_1254,In_15,In_2365);
and U1255 (N_1255,In_1519,In_594);
and U1256 (N_1256,In_223,In_440);
nor U1257 (N_1257,In_790,In_1803);
and U1258 (N_1258,In_861,In_1257);
nor U1259 (N_1259,In_1747,In_1507);
and U1260 (N_1260,In_1316,In_788);
xor U1261 (N_1261,In_711,In_1661);
nor U1262 (N_1262,In_67,In_1639);
or U1263 (N_1263,In_1693,In_924);
or U1264 (N_1264,In_101,In_257);
xnor U1265 (N_1265,In_563,In_194);
and U1266 (N_1266,In_1307,In_1482);
xor U1267 (N_1267,In_1168,In_2264);
nor U1268 (N_1268,In_2189,In_15);
and U1269 (N_1269,In_1912,In_104);
nor U1270 (N_1270,In_2470,In_16);
nor U1271 (N_1271,In_485,In_2464);
and U1272 (N_1272,In_266,In_2159);
and U1273 (N_1273,In_1566,In_1330);
nor U1274 (N_1274,In_1530,In_2476);
nand U1275 (N_1275,In_63,In_1954);
nand U1276 (N_1276,In_762,In_2396);
and U1277 (N_1277,In_1723,In_288);
and U1278 (N_1278,In_621,In_1859);
nand U1279 (N_1279,In_1603,In_1431);
or U1280 (N_1280,In_1621,In_522);
and U1281 (N_1281,In_2062,In_1625);
and U1282 (N_1282,In_1534,In_817);
nor U1283 (N_1283,In_574,In_1030);
or U1284 (N_1284,In_817,In_1440);
or U1285 (N_1285,In_899,In_372);
nor U1286 (N_1286,In_488,In_2270);
nand U1287 (N_1287,In_276,In_906);
nor U1288 (N_1288,In_1268,In_1377);
nand U1289 (N_1289,In_1243,In_2051);
nand U1290 (N_1290,In_991,In_763);
or U1291 (N_1291,In_2348,In_461);
and U1292 (N_1292,In_203,In_260);
nand U1293 (N_1293,In_1484,In_1412);
and U1294 (N_1294,In_1965,In_1688);
nor U1295 (N_1295,In_395,In_451);
nor U1296 (N_1296,In_1893,In_803);
nor U1297 (N_1297,In_2206,In_2240);
or U1298 (N_1298,In_756,In_1494);
and U1299 (N_1299,In_1826,In_797);
nor U1300 (N_1300,In_2139,In_2062);
nor U1301 (N_1301,In_1412,In_1083);
nor U1302 (N_1302,In_2411,In_2032);
or U1303 (N_1303,In_1553,In_1757);
and U1304 (N_1304,In_64,In_383);
nand U1305 (N_1305,In_1595,In_1880);
nor U1306 (N_1306,In_1712,In_1620);
nand U1307 (N_1307,In_246,In_895);
and U1308 (N_1308,In_1222,In_526);
nand U1309 (N_1309,In_1367,In_1285);
nor U1310 (N_1310,In_2190,In_662);
nand U1311 (N_1311,In_960,In_1740);
nand U1312 (N_1312,In_1096,In_2251);
nand U1313 (N_1313,In_1857,In_656);
xor U1314 (N_1314,In_883,In_664);
nand U1315 (N_1315,In_2249,In_1151);
or U1316 (N_1316,In_182,In_1325);
and U1317 (N_1317,In_634,In_1895);
nand U1318 (N_1318,In_1641,In_600);
nor U1319 (N_1319,In_2192,In_904);
and U1320 (N_1320,In_1473,In_1166);
nand U1321 (N_1321,In_357,In_1072);
xnor U1322 (N_1322,In_123,In_2440);
and U1323 (N_1323,In_1215,In_1890);
nand U1324 (N_1324,In_312,In_652);
or U1325 (N_1325,In_303,In_45);
nand U1326 (N_1326,In_2272,In_2033);
and U1327 (N_1327,In_1650,In_477);
nand U1328 (N_1328,In_2135,In_1620);
nand U1329 (N_1329,In_1290,In_934);
nand U1330 (N_1330,In_1418,In_2467);
and U1331 (N_1331,In_2302,In_1426);
and U1332 (N_1332,In_232,In_1240);
xnor U1333 (N_1333,In_1897,In_2480);
xnor U1334 (N_1334,In_2332,In_2316);
xnor U1335 (N_1335,In_105,In_1879);
nor U1336 (N_1336,In_915,In_2455);
nor U1337 (N_1337,In_1029,In_387);
nand U1338 (N_1338,In_2439,In_290);
nand U1339 (N_1339,In_2172,In_863);
or U1340 (N_1340,In_955,In_2011);
and U1341 (N_1341,In_118,In_531);
xnor U1342 (N_1342,In_1259,In_1092);
nor U1343 (N_1343,In_265,In_1232);
or U1344 (N_1344,In_1411,In_277);
xnor U1345 (N_1345,In_1530,In_27);
nand U1346 (N_1346,In_1959,In_409);
nand U1347 (N_1347,In_1835,In_392);
nor U1348 (N_1348,In_1346,In_544);
or U1349 (N_1349,In_1608,In_2054);
nor U1350 (N_1350,In_2148,In_1624);
nor U1351 (N_1351,In_1673,In_94);
nor U1352 (N_1352,In_1968,In_2210);
nand U1353 (N_1353,In_51,In_1916);
or U1354 (N_1354,In_306,In_1744);
nand U1355 (N_1355,In_1230,In_1956);
nand U1356 (N_1356,In_213,In_1243);
xor U1357 (N_1357,In_1468,In_937);
nand U1358 (N_1358,In_687,In_1512);
and U1359 (N_1359,In_714,In_1881);
nand U1360 (N_1360,In_401,In_301);
or U1361 (N_1361,In_2495,In_272);
and U1362 (N_1362,In_1419,In_1873);
and U1363 (N_1363,In_1493,In_909);
or U1364 (N_1364,In_2321,In_1828);
or U1365 (N_1365,In_1585,In_1338);
or U1366 (N_1366,In_2112,In_16);
and U1367 (N_1367,In_394,In_486);
nand U1368 (N_1368,In_206,In_2379);
or U1369 (N_1369,In_2344,In_536);
nand U1370 (N_1370,In_1942,In_103);
and U1371 (N_1371,In_1139,In_1902);
or U1372 (N_1372,In_1498,In_2105);
nand U1373 (N_1373,In_1831,In_1053);
nand U1374 (N_1374,In_263,In_1236);
nor U1375 (N_1375,In_1380,In_2334);
xor U1376 (N_1376,In_728,In_311);
nand U1377 (N_1377,In_1839,In_192);
or U1378 (N_1378,In_2130,In_175);
and U1379 (N_1379,In_516,In_248);
and U1380 (N_1380,In_1305,In_386);
or U1381 (N_1381,In_1043,In_1372);
or U1382 (N_1382,In_1004,In_816);
or U1383 (N_1383,In_1379,In_2150);
nand U1384 (N_1384,In_508,In_1203);
nand U1385 (N_1385,In_1036,In_652);
or U1386 (N_1386,In_2482,In_92);
nor U1387 (N_1387,In_1935,In_1866);
and U1388 (N_1388,In_1512,In_62);
or U1389 (N_1389,In_875,In_1168);
nand U1390 (N_1390,In_2255,In_2034);
nor U1391 (N_1391,In_99,In_2058);
nor U1392 (N_1392,In_2294,In_1823);
nor U1393 (N_1393,In_2026,In_2425);
nand U1394 (N_1394,In_2254,In_1060);
nor U1395 (N_1395,In_744,In_354);
xnor U1396 (N_1396,In_1704,In_1521);
xnor U1397 (N_1397,In_633,In_1773);
and U1398 (N_1398,In_2269,In_2417);
xnor U1399 (N_1399,In_435,In_649);
and U1400 (N_1400,In_646,In_1989);
nor U1401 (N_1401,In_1821,In_2029);
or U1402 (N_1402,In_2399,In_1299);
or U1403 (N_1403,In_1417,In_52);
nor U1404 (N_1404,In_1184,In_823);
or U1405 (N_1405,In_2499,In_1819);
nor U1406 (N_1406,In_732,In_1314);
and U1407 (N_1407,In_757,In_1264);
and U1408 (N_1408,In_1690,In_213);
or U1409 (N_1409,In_2435,In_1595);
nor U1410 (N_1410,In_530,In_240);
or U1411 (N_1411,In_1621,In_293);
xnor U1412 (N_1412,In_1841,In_886);
or U1413 (N_1413,In_1337,In_1762);
and U1414 (N_1414,In_2212,In_1509);
nand U1415 (N_1415,In_234,In_409);
nor U1416 (N_1416,In_890,In_180);
and U1417 (N_1417,In_47,In_1717);
or U1418 (N_1418,In_1651,In_424);
and U1419 (N_1419,In_1405,In_779);
or U1420 (N_1420,In_2422,In_1313);
nor U1421 (N_1421,In_2106,In_1636);
and U1422 (N_1422,In_67,In_493);
xor U1423 (N_1423,In_1605,In_2373);
nand U1424 (N_1424,In_727,In_142);
and U1425 (N_1425,In_1760,In_1862);
nor U1426 (N_1426,In_1081,In_1201);
or U1427 (N_1427,In_54,In_1948);
nor U1428 (N_1428,In_453,In_2333);
nor U1429 (N_1429,In_775,In_1676);
nor U1430 (N_1430,In_2467,In_34);
or U1431 (N_1431,In_1891,In_1449);
and U1432 (N_1432,In_762,In_1786);
and U1433 (N_1433,In_760,In_883);
or U1434 (N_1434,In_854,In_1233);
nand U1435 (N_1435,In_1686,In_2042);
nor U1436 (N_1436,In_1623,In_1557);
xor U1437 (N_1437,In_1452,In_378);
nand U1438 (N_1438,In_919,In_208);
or U1439 (N_1439,In_2270,In_557);
and U1440 (N_1440,In_885,In_1085);
and U1441 (N_1441,In_770,In_2133);
nand U1442 (N_1442,In_806,In_1426);
nor U1443 (N_1443,In_448,In_256);
nor U1444 (N_1444,In_1511,In_2129);
nor U1445 (N_1445,In_1434,In_1141);
nor U1446 (N_1446,In_2298,In_1367);
nor U1447 (N_1447,In_476,In_613);
xor U1448 (N_1448,In_242,In_1753);
nand U1449 (N_1449,In_497,In_2391);
or U1450 (N_1450,In_515,In_631);
nand U1451 (N_1451,In_498,In_1203);
nand U1452 (N_1452,In_1840,In_684);
nor U1453 (N_1453,In_916,In_1604);
nor U1454 (N_1454,In_588,In_1199);
nor U1455 (N_1455,In_1587,In_61);
or U1456 (N_1456,In_737,In_2308);
nor U1457 (N_1457,In_66,In_1917);
xor U1458 (N_1458,In_1040,In_2179);
or U1459 (N_1459,In_375,In_1966);
xnor U1460 (N_1460,In_933,In_2228);
or U1461 (N_1461,In_2071,In_1551);
nor U1462 (N_1462,In_1612,In_2229);
or U1463 (N_1463,In_835,In_1749);
nor U1464 (N_1464,In_1190,In_696);
nand U1465 (N_1465,In_366,In_1000);
xnor U1466 (N_1466,In_1640,In_36);
or U1467 (N_1467,In_1362,In_1213);
or U1468 (N_1468,In_1992,In_2133);
nor U1469 (N_1469,In_1094,In_2128);
nor U1470 (N_1470,In_1240,In_2210);
nor U1471 (N_1471,In_2269,In_1381);
xnor U1472 (N_1472,In_616,In_142);
nor U1473 (N_1473,In_1057,In_1123);
or U1474 (N_1474,In_1019,In_1785);
and U1475 (N_1475,In_1184,In_840);
and U1476 (N_1476,In_553,In_317);
nor U1477 (N_1477,In_1809,In_2348);
nand U1478 (N_1478,In_1049,In_1953);
and U1479 (N_1479,In_1613,In_1070);
nor U1480 (N_1480,In_702,In_2);
and U1481 (N_1481,In_1080,In_96);
or U1482 (N_1482,In_628,In_1376);
and U1483 (N_1483,In_2145,In_1545);
nand U1484 (N_1484,In_1714,In_543);
and U1485 (N_1485,In_1156,In_116);
or U1486 (N_1486,In_2067,In_347);
or U1487 (N_1487,In_249,In_1586);
nor U1488 (N_1488,In_659,In_955);
and U1489 (N_1489,In_791,In_55);
and U1490 (N_1490,In_1572,In_959);
nor U1491 (N_1491,In_279,In_1429);
and U1492 (N_1492,In_757,In_1847);
and U1493 (N_1493,In_868,In_62);
nand U1494 (N_1494,In_385,In_578);
xnor U1495 (N_1495,In_468,In_20);
nand U1496 (N_1496,In_475,In_1295);
and U1497 (N_1497,In_1228,In_859);
and U1498 (N_1498,In_2188,In_865);
nor U1499 (N_1499,In_1496,In_1885);
nand U1500 (N_1500,In_1649,In_365);
or U1501 (N_1501,In_236,In_1295);
or U1502 (N_1502,In_1450,In_1692);
nor U1503 (N_1503,In_48,In_1536);
xor U1504 (N_1504,In_15,In_1439);
nand U1505 (N_1505,In_1668,In_1944);
nor U1506 (N_1506,In_603,In_2344);
nand U1507 (N_1507,In_1117,In_1600);
nor U1508 (N_1508,In_1565,In_335);
nand U1509 (N_1509,In_1741,In_2481);
nand U1510 (N_1510,In_839,In_16);
nand U1511 (N_1511,In_1928,In_2489);
xor U1512 (N_1512,In_1484,In_2096);
and U1513 (N_1513,In_2156,In_1798);
nand U1514 (N_1514,In_2490,In_649);
xor U1515 (N_1515,In_1751,In_1985);
nand U1516 (N_1516,In_999,In_93);
and U1517 (N_1517,In_850,In_1511);
nor U1518 (N_1518,In_51,In_2286);
or U1519 (N_1519,In_1348,In_870);
or U1520 (N_1520,In_1468,In_84);
nor U1521 (N_1521,In_1777,In_862);
nand U1522 (N_1522,In_1085,In_2042);
nand U1523 (N_1523,In_1829,In_529);
or U1524 (N_1524,In_2258,In_1297);
or U1525 (N_1525,In_1738,In_210);
or U1526 (N_1526,In_1766,In_2470);
nand U1527 (N_1527,In_229,In_2427);
and U1528 (N_1528,In_2334,In_2418);
xnor U1529 (N_1529,In_897,In_1896);
nor U1530 (N_1530,In_2326,In_318);
or U1531 (N_1531,In_1943,In_364);
or U1532 (N_1532,In_266,In_2487);
and U1533 (N_1533,In_2321,In_1426);
and U1534 (N_1534,In_697,In_250);
xnor U1535 (N_1535,In_583,In_1262);
nand U1536 (N_1536,In_180,In_1075);
or U1537 (N_1537,In_1755,In_2305);
nor U1538 (N_1538,In_2109,In_782);
nand U1539 (N_1539,In_2169,In_483);
and U1540 (N_1540,In_1592,In_2451);
and U1541 (N_1541,In_1316,In_1017);
nand U1542 (N_1542,In_1600,In_2014);
nand U1543 (N_1543,In_692,In_544);
or U1544 (N_1544,In_538,In_640);
or U1545 (N_1545,In_1774,In_2466);
nand U1546 (N_1546,In_472,In_1322);
nand U1547 (N_1547,In_1614,In_888);
or U1548 (N_1548,In_1707,In_1008);
or U1549 (N_1549,In_180,In_1570);
xor U1550 (N_1550,In_1947,In_628);
and U1551 (N_1551,In_1213,In_2021);
xor U1552 (N_1552,In_747,In_39);
xor U1553 (N_1553,In_1192,In_518);
nor U1554 (N_1554,In_267,In_1669);
nor U1555 (N_1555,In_983,In_1365);
nor U1556 (N_1556,In_1050,In_1104);
nor U1557 (N_1557,In_394,In_700);
and U1558 (N_1558,In_1957,In_2350);
and U1559 (N_1559,In_1048,In_1086);
or U1560 (N_1560,In_644,In_1648);
or U1561 (N_1561,In_2317,In_1602);
nand U1562 (N_1562,In_1589,In_511);
or U1563 (N_1563,In_1707,In_306);
and U1564 (N_1564,In_1410,In_1650);
nand U1565 (N_1565,In_197,In_873);
nand U1566 (N_1566,In_435,In_1881);
or U1567 (N_1567,In_2481,In_1814);
nand U1568 (N_1568,In_1433,In_798);
and U1569 (N_1569,In_2378,In_1377);
and U1570 (N_1570,In_1486,In_90);
or U1571 (N_1571,In_1479,In_931);
nor U1572 (N_1572,In_1729,In_2145);
or U1573 (N_1573,In_2023,In_1839);
nand U1574 (N_1574,In_274,In_2105);
or U1575 (N_1575,In_675,In_2423);
and U1576 (N_1576,In_1133,In_1603);
nand U1577 (N_1577,In_956,In_241);
xnor U1578 (N_1578,In_1118,In_1122);
nor U1579 (N_1579,In_164,In_1807);
xnor U1580 (N_1580,In_220,In_318);
xnor U1581 (N_1581,In_1033,In_1175);
or U1582 (N_1582,In_1503,In_1365);
or U1583 (N_1583,In_1461,In_1602);
or U1584 (N_1584,In_2420,In_1928);
or U1585 (N_1585,In_930,In_1585);
nand U1586 (N_1586,In_1742,In_1424);
xnor U1587 (N_1587,In_735,In_2079);
and U1588 (N_1588,In_2254,In_1275);
and U1589 (N_1589,In_779,In_1939);
nand U1590 (N_1590,In_943,In_2392);
xnor U1591 (N_1591,In_633,In_706);
and U1592 (N_1592,In_1655,In_458);
nor U1593 (N_1593,In_1675,In_2491);
or U1594 (N_1594,In_2296,In_2248);
and U1595 (N_1595,In_2475,In_1100);
and U1596 (N_1596,In_1789,In_1942);
or U1597 (N_1597,In_2182,In_2151);
and U1598 (N_1598,In_389,In_1564);
xor U1599 (N_1599,In_1573,In_1773);
and U1600 (N_1600,In_2042,In_283);
and U1601 (N_1601,In_379,In_2191);
nor U1602 (N_1602,In_1316,In_2224);
xor U1603 (N_1603,In_991,In_834);
or U1604 (N_1604,In_326,In_97);
xnor U1605 (N_1605,In_1852,In_1769);
and U1606 (N_1606,In_2253,In_2112);
nor U1607 (N_1607,In_1775,In_200);
and U1608 (N_1608,In_2065,In_1857);
nand U1609 (N_1609,In_422,In_1828);
and U1610 (N_1610,In_29,In_1726);
or U1611 (N_1611,In_375,In_651);
nand U1612 (N_1612,In_720,In_1439);
nor U1613 (N_1613,In_2184,In_876);
or U1614 (N_1614,In_1902,In_555);
and U1615 (N_1615,In_29,In_1097);
nor U1616 (N_1616,In_2189,In_2243);
or U1617 (N_1617,In_1749,In_1644);
nor U1618 (N_1618,In_1079,In_2450);
nor U1619 (N_1619,In_1089,In_1763);
and U1620 (N_1620,In_883,In_2334);
nand U1621 (N_1621,In_32,In_696);
nand U1622 (N_1622,In_1124,In_667);
nand U1623 (N_1623,In_2005,In_767);
and U1624 (N_1624,In_418,In_2358);
or U1625 (N_1625,In_2341,In_2453);
nand U1626 (N_1626,In_2379,In_2437);
and U1627 (N_1627,In_2020,In_1594);
and U1628 (N_1628,In_1986,In_2466);
xor U1629 (N_1629,In_2281,In_266);
or U1630 (N_1630,In_910,In_542);
nor U1631 (N_1631,In_1526,In_1788);
or U1632 (N_1632,In_2054,In_1842);
nor U1633 (N_1633,In_1830,In_1820);
or U1634 (N_1634,In_2250,In_1832);
or U1635 (N_1635,In_2210,In_266);
nand U1636 (N_1636,In_664,In_524);
and U1637 (N_1637,In_202,In_2052);
and U1638 (N_1638,In_421,In_1614);
and U1639 (N_1639,In_2210,In_1593);
nor U1640 (N_1640,In_890,In_512);
nand U1641 (N_1641,In_2140,In_1496);
nand U1642 (N_1642,In_2002,In_358);
nor U1643 (N_1643,In_592,In_2335);
or U1644 (N_1644,In_164,In_211);
and U1645 (N_1645,In_471,In_1643);
nand U1646 (N_1646,In_1840,In_1938);
nor U1647 (N_1647,In_892,In_1271);
or U1648 (N_1648,In_1751,In_1827);
nand U1649 (N_1649,In_915,In_2048);
nor U1650 (N_1650,In_975,In_2312);
or U1651 (N_1651,In_1725,In_2123);
and U1652 (N_1652,In_890,In_452);
nand U1653 (N_1653,In_1377,In_1292);
or U1654 (N_1654,In_1274,In_299);
nand U1655 (N_1655,In_2031,In_1049);
or U1656 (N_1656,In_1550,In_1858);
and U1657 (N_1657,In_1868,In_1045);
or U1658 (N_1658,In_503,In_988);
nand U1659 (N_1659,In_2467,In_413);
and U1660 (N_1660,In_1953,In_2438);
nor U1661 (N_1661,In_69,In_2236);
nand U1662 (N_1662,In_446,In_1306);
and U1663 (N_1663,In_2273,In_2240);
nand U1664 (N_1664,In_2319,In_1454);
xor U1665 (N_1665,In_608,In_1355);
nand U1666 (N_1666,In_1174,In_1098);
and U1667 (N_1667,In_534,In_1333);
nand U1668 (N_1668,In_2421,In_393);
or U1669 (N_1669,In_1407,In_2464);
xnor U1670 (N_1670,In_766,In_1464);
xor U1671 (N_1671,In_1516,In_1339);
nand U1672 (N_1672,In_1456,In_2160);
xor U1673 (N_1673,In_2182,In_2025);
and U1674 (N_1674,In_566,In_1741);
nand U1675 (N_1675,In_37,In_2235);
and U1676 (N_1676,In_1477,In_866);
and U1677 (N_1677,In_639,In_429);
or U1678 (N_1678,In_2341,In_1982);
nor U1679 (N_1679,In_210,In_1161);
nor U1680 (N_1680,In_292,In_2381);
and U1681 (N_1681,In_1059,In_424);
and U1682 (N_1682,In_1645,In_416);
nand U1683 (N_1683,In_1156,In_341);
nand U1684 (N_1684,In_384,In_709);
nand U1685 (N_1685,In_1315,In_1852);
and U1686 (N_1686,In_1945,In_1463);
nor U1687 (N_1687,In_1902,In_1603);
or U1688 (N_1688,In_1856,In_544);
nor U1689 (N_1689,In_574,In_558);
and U1690 (N_1690,In_1010,In_56);
nor U1691 (N_1691,In_555,In_1113);
nor U1692 (N_1692,In_1607,In_1918);
or U1693 (N_1693,In_1526,In_778);
xnor U1694 (N_1694,In_2183,In_235);
nor U1695 (N_1695,In_2485,In_662);
nor U1696 (N_1696,In_193,In_305);
nand U1697 (N_1697,In_1930,In_2402);
and U1698 (N_1698,In_2380,In_179);
nand U1699 (N_1699,In_2220,In_1516);
or U1700 (N_1700,In_2383,In_2489);
xor U1701 (N_1701,In_2158,In_448);
nor U1702 (N_1702,In_503,In_1642);
or U1703 (N_1703,In_803,In_557);
and U1704 (N_1704,In_1062,In_296);
and U1705 (N_1705,In_1697,In_2053);
and U1706 (N_1706,In_1470,In_921);
nand U1707 (N_1707,In_1867,In_808);
nor U1708 (N_1708,In_2346,In_1498);
xor U1709 (N_1709,In_141,In_646);
and U1710 (N_1710,In_1388,In_1519);
nor U1711 (N_1711,In_40,In_173);
or U1712 (N_1712,In_1174,In_715);
and U1713 (N_1713,In_1761,In_706);
or U1714 (N_1714,In_366,In_721);
and U1715 (N_1715,In_1808,In_1576);
nor U1716 (N_1716,In_1776,In_196);
or U1717 (N_1717,In_688,In_1153);
and U1718 (N_1718,In_1923,In_2038);
nor U1719 (N_1719,In_256,In_1688);
or U1720 (N_1720,In_2272,In_1499);
or U1721 (N_1721,In_2045,In_2383);
or U1722 (N_1722,In_2070,In_1433);
and U1723 (N_1723,In_1151,In_666);
nand U1724 (N_1724,In_1758,In_1890);
or U1725 (N_1725,In_1386,In_1399);
xor U1726 (N_1726,In_2145,In_308);
or U1727 (N_1727,In_960,In_921);
nand U1728 (N_1728,In_1554,In_433);
nor U1729 (N_1729,In_1969,In_1165);
nor U1730 (N_1730,In_2030,In_1942);
or U1731 (N_1731,In_894,In_543);
and U1732 (N_1732,In_527,In_1688);
nand U1733 (N_1733,In_1468,In_2188);
nor U1734 (N_1734,In_2058,In_652);
and U1735 (N_1735,In_436,In_2377);
nand U1736 (N_1736,In_1674,In_571);
or U1737 (N_1737,In_1249,In_1991);
or U1738 (N_1738,In_537,In_1267);
and U1739 (N_1739,In_2137,In_745);
and U1740 (N_1740,In_1713,In_273);
nand U1741 (N_1741,In_177,In_2443);
xnor U1742 (N_1742,In_701,In_1286);
nor U1743 (N_1743,In_1523,In_1910);
or U1744 (N_1744,In_223,In_158);
nand U1745 (N_1745,In_1228,In_601);
nand U1746 (N_1746,In_1389,In_139);
or U1747 (N_1747,In_1062,In_645);
and U1748 (N_1748,In_628,In_1490);
xor U1749 (N_1749,In_900,In_1645);
and U1750 (N_1750,In_2063,In_833);
and U1751 (N_1751,In_138,In_221);
nand U1752 (N_1752,In_97,In_340);
or U1753 (N_1753,In_1992,In_1158);
xnor U1754 (N_1754,In_1421,In_2194);
nand U1755 (N_1755,In_659,In_2375);
nand U1756 (N_1756,In_2048,In_86);
and U1757 (N_1757,In_1008,In_236);
nand U1758 (N_1758,In_706,In_642);
nand U1759 (N_1759,In_642,In_717);
xor U1760 (N_1760,In_147,In_1209);
or U1761 (N_1761,In_1676,In_1952);
xnor U1762 (N_1762,In_993,In_990);
xnor U1763 (N_1763,In_111,In_1178);
nand U1764 (N_1764,In_87,In_2054);
or U1765 (N_1765,In_2125,In_1694);
xor U1766 (N_1766,In_637,In_1758);
xor U1767 (N_1767,In_1864,In_106);
nor U1768 (N_1768,In_2300,In_1185);
or U1769 (N_1769,In_549,In_1577);
or U1770 (N_1770,In_2035,In_1404);
nor U1771 (N_1771,In_252,In_2389);
and U1772 (N_1772,In_1744,In_1622);
or U1773 (N_1773,In_2002,In_1612);
nand U1774 (N_1774,In_1260,In_572);
and U1775 (N_1775,In_562,In_2003);
and U1776 (N_1776,In_2155,In_917);
nor U1777 (N_1777,In_538,In_1730);
nand U1778 (N_1778,In_420,In_1072);
and U1779 (N_1779,In_1858,In_1270);
nand U1780 (N_1780,In_473,In_573);
or U1781 (N_1781,In_277,In_1269);
or U1782 (N_1782,In_835,In_2272);
xor U1783 (N_1783,In_2172,In_964);
nand U1784 (N_1784,In_2382,In_409);
and U1785 (N_1785,In_1940,In_254);
or U1786 (N_1786,In_1007,In_1888);
or U1787 (N_1787,In_2172,In_48);
or U1788 (N_1788,In_1106,In_1606);
and U1789 (N_1789,In_383,In_156);
and U1790 (N_1790,In_1041,In_139);
or U1791 (N_1791,In_2059,In_691);
nor U1792 (N_1792,In_1713,In_453);
or U1793 (N_1793,In_1571,In_1671);
nand U1794 (N_1794,In_1909,In_2259);
xnor U1795 (N_1795,In_740,In_650);
nand U1796 (N_1796,In_1993,In_563);
or U1797 (N_1797,In_772,In_2394);
nand U1798 (N_1798,In_2133,In_743);
or U1799 (N_1799,In_1582,In_1395);
xor U1800 (N_1800,In_265,In_831);
and U1801 (N_1801,In_1904,In_1629);
nand U1802 (N_1802,In_329,In_1611);
nor U1803 (N_1803,In_468,In_1437);
nand U1804 (N_1804,In_1759,In_62);
nand U1805 (N_1805,In_2411,In_416);
or U1806 (N_1806,In_556,In_2268);
nand U1807 (N_1807,In_254,In_246);
nor U1808 (N_1808,In_665,In_1080);
nand U1809 (N_1809,In_2491,In_936);
nor U1810 (N_1810,In_208,In_104);
and U1811 (N_1811,In_1748,In_651);
nor U1812 (N_1812,In_424,In_1140);
nand U1813 (N_1813,In_867,In_2287);
and U1814 (N_1814,In_1059,In_1758);
or U1815 (N_1815,In_665,In_686);
nor U1816 (N_1816,In_458,In_1309);
nor U1817 (N_1817,In_583,In_935);
and U1818 (N_1818,In_43,In_1056);
nand U1819 (N_1819,In_2402,In_1565);
and U1820 (N_1820,In_2066,In_959);
xnor U1821 (N_1821,In_372,In_141);
nand U1822 (N_1822,In_860,In_1446);
nor U1823 (N_1823,In_16,In_2421);
and U1824 (N_1824,In_1200,In_1537);
nand U1825 (N_1825,In_594,In_9);
nand U1826 (N_1826,In_974,In_537);
or U1827 (N_1827,In_1891,In_1791);
nor U1828 (N_1828,In_2318,In_927);
or U1829 (N_1829,In_923,In_355);
xnor U1830 (N_1830,In_1264,In_303);
nand U1831 (N_1831,In_822,In_2471);
or U1832 (N_1832,In_76,In_940);
or U1833 (N_1833,In_128,In_392);
nand U1834 (N_1834,In_13,In_1326);
or U1835 (N_1835,In_179,In_101);
nor U1836 (N_1836,In_654,In_2267);
nor U1837 (N_1837,In_888,In_474);
and U1838 (N_1838,In_73,In_2173);
xor U1839 (N_1839,In_1068,In_2256);
and U1840 (N_1840,In_2266,In_500);
or U1841 (N_1841,In_636,In_2280);
xor U1842 (N_1842,In_1537,In_398);
and U1843 (N_1843,In_1556,In_1766);
and U1844 (N_1844,In_82,In_881);
xor U1845 (N_1845,In_1933,In_1443);
and U1846 (N_1846,In_1578,In_125);
and U1847 (N_1847,In_1076,In_2215);
and U1848 (N_1848,In_373,In_143);
and U1849 (N_1849,In_759,In_1692);
nor U1850 (N_1850,In_1624,In_2424);
xnor U1851 (N_1851,In_2212,In_1333);
nor U1852 (N_1852,In_1371,In_720);
nand U1853 (N_1853,In_1389,In_2354);
nand U1854 (N_1854,In_2196,In_2185);
and U1855 (N_1855,In_814,In_131);
or U1856 (N_1856,In_1209,In_1881);
xor U1857 (N_1857,In_2035,In_2128);
nand U1858 (N_1858,In_708,In_1162);
xor U1859 (N_1859,In_1607,In_850);
nor U1860 (N_1860,In_1134,In_1250);
and U1861 (N_1861,In_2048,In_1094);
or U1862 (N_1862,In_949,In_76);
nand U1863 (N_1863,In_2396,In_719);
or U1864 (N_1864,In_1163,In_339);
nand U1865 (N_1865,In_1529,In_1944);
nor U1866 (N_1866,In_1497,In_280);
or U1867 (N_1867,In_1782,In_120);
or U1868 (N_1868,In_476,In_2362);
nor U1869 (N_1869,In_546,In_604);
nor U1870 (N_1870,In_872,In_2002);
xor U1871 (N_1871,In_1090,In_629);
nor U1872 (N_1872,In_163,In_507);
or U1873 (N_1873,In_2315,In_1552);
nor U1874 (N_1874,In_1712,In_718);
or U1875 (N_1875,In_1639,In_378);
nor U1876 (N_1876,In_633,In_1336);
and U1877 (N_1877,In_1757,In_866);
nor U1878 (N_1878,In_369,In_1659);
nor U1879 (N_1879,In_984,In_923);
nor U1880 (N_1880,In_1151,In_2491);
and U1881 (N_1881,In_1696,In_1694);
nor U1882 (N_1882,In_1341,In_2073);
and U1883 (N_1883,In_787,In_1397);
and U1884 (N_1884,In_438,In_1373);
and U1885 (N_1885,In_2037,In_2284);
nor U1886 (N_1886,In_987,In_832);
nor U1887 (N_1887,In_1200,In_1960);
nor U1888 (N_1888,In_1324,In_813);
and U1889 (N_1889,In_2107,In_89);
nor U1890 (N_1890,In_2359,In_444);
xnor U1891 (N_1891,In_707,In_2424);
xor U1892 (N_1892,In_2010,In_434);
nand U1893 (N_1893,In_557,In_614);
nand U1894 (N_1894,In_2412,In_363);
nand U1895 (N_1895,In_2025,In_608);
nor U1896 (N_1896,In_722,In_169);
and U1897 (N_1897,In_1672,In_550);
xnor U1898 (N_1898,In_2330,In_2483);
nor U1899 (N_1899,In_369,In_185);
nor U1900 (N_1900,In_1364,In_358);
and U1901 (N_1901,In_499,In_1434);
nor U1902 (N_1902,In_672,In_1103);
and U1903 (N_1903,In_1701,In_2007);
nand U1904 (N_1904,In_1218,In_2384);
or U1905 (N_1905,In_1159,In_2319);
and U1906 (N_1906,In_1425,In_2129);
nand U1907 (N_1907,In_737,In_1889);
and U1908 (N_1908,In_244,In_2387);
and U1909 (N_1909,In_1181,In_1058);
and U1910 (N_1910,In_1182,In_717);
or U1911 (N_1911,In_249,In_2344);
nor U1912 (N_1912,In_2263,In_52);
xor U1913 (N_1913,In_1126,In_1634);
and U1914 (N_1914,In_713,In_517);
nand U1915 (N_1915,In_568,In_2370);
xnor U1916 (N_1916,In_2166,In_1121);
or U1917 (N_1917,In_680,In_1341);
xnor U1918 (N_1918,In_42,In_2423);
xnor U1919 (N_1919,In_928,In_2249);
nor U1920 (N_1920,In_1906,In_815);
nand U1921 (N_1921,In_1568,In_2453);
and U1922 (N_1922,In_2358,In_1635);
nor U1923 (N_1923,In_2180,In_2380);
nor U1924 (N_1924,In_891,In_1404);
or U1925 (N_1925,In_2032,In_2392);
and U1926 (N_1926,In_1391,In_225);
nor U1927 (N_1927,In_929,In_175);
xor U1928 (N_1928,In_1723,In_1258);
nand U1929 (N_1929,In_2474,In_1362);
and U1930 (N_1930,In_524,In_881);
nor U1931 (N_1931,In_191,In_2179);
and U1932 (N_1932,In_2150,In_312);
and U1933 (N_1933,In_1454,In_687);
and U1934 (N_1934,In_1204,In_1553);
and U1935 (N_1935,In_390,In_1202);
nand U1936 (N_1936,In_2355,In_65);
or U1937 (N_1937,In_1783,In_1287);
and U1938 (N_1938,In_2043,In_2458);
nor U1939 (N_1939,In_950,In_2403);
nand U1940 (N_1940,In_758,In_1575);
xnor U1941 (N_1941,In_1602,In_2000);
and U1942 (N_1942,In_1414,In_990);
or U1943 (N_1943,In_699,In_2138);
nand U1944 (N_1944,In_1128,In_1195);
nand U1945 (N_1945,In_2322,In_2219);
xor U1946 (N_1946,In_718,In_2093);
xor U1947 (N_1947,In_170,In_532);
or U1948 (N_1948,In_754,In_1809);
nor U1949 (N_1949,In_1079,In_1142);
nor U1950 (N_1950,In_2195,In_1302);
xnor U1951 (N_1951,In_2441,In_1402);
and U1952 (N_1952,In_1284,In_1425);
nand U1953 (N_1953,In_643,In_1133);
nand U1954 (N_1954,In_892,In_1963);
or U1955 (N_1955,In_1759,In_210);
nor U1956 (N_1956,In_1889,In_576);
nor U1957 (N_1957,In_820,In_9);
nor U1958 (N_1958,In_1220,In_957);
nor U1959 (N_1959,In_1065,In_205);
nand U1960 (N_1960,In_1570,In_1281);
xnor U1961 (N_1961,In_178,In_2235);
and U1962 (N_1962,In_795,In_30);
or U1963 (N_1963,In_842,In_1916);
or U1964 (N_1964,In_604,In_502);
and U1965 (N_1965,In_1819,In_2309);
or U1966 (N_1966,In_1747,In_964);
nor U1967 (N_1967,In_781,In_1327);
nand U1968 (N_1968,In_2343,In_1454);
or U1969 (N_1969,In_659,In_231);
nand U1970 (N_1970,In_1403,In_2399);
and U1971 (N_1971,In_717,In_162);
nor U1972 (N_1972,In_1713,In_2259);
nand U1973 (N_1973,In_1929,In_1829);
nor U1974 (N_1974,In_1428,In_1004);
nand U1975 (N_1975,In_2114,In_1444);
or U1976 (N_1976,In_2123,In_703);
nand U1977 (N_1977,In_323,In_1638);
nor U1978 (N_1978,In_1774,In_1388);
xnor U1979 (N_1979,In_2178,In_215);
nand U1980 (N_1980,In_2301,In_568);
nor U1981 (N_1981,In_37,In_599);
nor U1982 (N_1982,In_755,In_1247);
or U1983 (N_1983,In_2216,In_1095);
or U1984 (N_1984,In_238,In_396);
and U1985 (N_1985,In_1083,In_1322);
and U1986 (N_1986,In_2462,In_1688);
nand U1987 (N_1987,In_130,In_2029);
and U1988 (N_1988,In_1318,In_390);
nand U1989 (N_1989,In_1802,In_1391);
nor U1990 (N_1990,In_1068,In_650);
or U1991 (N_1991,In_1663,In_689);
and U1992 (N_1992,In_2061,In_533);
nor U1993 (N_1993,In_140,In_2422);
and U1994 (N_1994,In_651,In_702);
or U1995 (N_1995,In_51,In_2491);
nor U1996 (N_1996,In_1864,In_616);
and U1997 (N_1997,In_1836,In_1065);
nand U1998 (N_1998,In_1291,In_1599);
xor U1999 (N_1999,In_1114,In_1904);
nand U2000 (N_2000,In_697,In_739);
xnor U2001 (N_2001,In_2485,In_1109);
or U2002 (N_2002,In_456,In_2129);
and U2003 (N_2003,In_1086,In_1877);
nor U2004 (N_2004,In_1641,In_2402);
nand U2005 (N_2005,In_290,In_1972);
or U2006 (N_2006,In_2471,In_1738);
or U2007 (N_2007,In_105,In_429);
or U2008 (N_2008,In_1572,In_993);
nand U2009 (N_2009,In_1192,In_1214);
xnor U2010 (N_2010,In_2361,In_1522);
nand U2011 (N_2011,In_404,In_1732);
nand U2012 (N_2012,In_2001,In_759);
nand U2013 (N_2013,In_1769,In_1306);
and U2014 (N_2014,In_2313,In_1047);
nor U2015 (N_2015,In_2251,In_482);
nand U2016 (N_2016,In_347,In_1951);
xor U2017 (N_2017,In_2157,In_1539);
nand U2018 (N_2018,In_2117,In_1800);
xnor U2019 (N_2019,In_1644,In_2065);
and U2020 (N_2020,In_1534,In_780);
or U2021 (N_2021,In_1543,In_1422);
or U2022 (N_2022,In_2491,In_196);
nor U2023 (N_2023,In_2451,In_1607);
nand U2024 (N_2024,In_706,In_676);
nand U2025 (N_2025,In_2218,In_2069);
nor U2026 (N_2026,In_1819,In_1273);
nand U2027 (N_2027,In_1152,In_2083);
or U2028 (N_2028,In_991,In_1404);
nand U2029 (N_2029,In_21,In_2021);
and U2030 (N_2030,In_1838,In_2184);
nor U2031 (N_2031,In_846,In_1489);
and U2032 (N_2032,In_703,In_1163);
nor U2033 (N_2033,In_1089,In_2371);
or U2034 (N_2034,In_404,In_2282);
nor U2035 (N_2035,In_1427,In_902);
and U2036 (N_2036,In_1868,In_361);
and U2037 (N_2037,In_2176,In_742);
nor U2038 (N_2038,In_2331,In_192);
or U2039 (N_2039,In_2492,In_640);
or U2040 (N_2040,In_2493,In_2421);
or U2041 (N_2041,In_2022,In_2430);
or U2042 (N_2042,In_953,In_639);
xnor U2043 (N_2043,In_1686,In_1582);
or U2044 (N_2044,In_2022,In_2210);
or U2045 (N_2045,In_1808,In_1148);
nand U2046 (N_2046,In_198,In_297);
and U2047 (N_2047,In_1277,In_2266);
or U2048 (N_2048,In_1424,In_2085);
and U2049 (N_2049,In_1431,In_292);
nand U2050 (N_2050,In_2328,In_1577);
and U2051 (N_2051,In_304,In_1045);
nand U2052 (N_2052,In_314,In_240);
xnor U2053 (N_2053,In_1172,In_1029);
nand U2054 (N_2054,In_2325,In_538);
nand U2055 (N_2055,In_795,In_790);
nand U2056 (N_2056,In_984,In_399);
or U2057 (N_2057,In_1044,In_631);
and U2058 (N_2058,In_1779,In_1815);
and U2059 (N_2059,In_1506,In_570);
and U2060 (N_2060,In_1883,In_835);
and U2061 (N_2061,In_1919,In_1033);
nor U2062 (N_2062,In_1633,In_2363);
nor U2063 (N_2063,In_2388,In_1772);
or U2064 (N_2064,In_1634,In_1992);
and U2065 (N_2065,In_439,In_1806);
nor U2066 (N_2066,In_2440,In_825);
nor U2067 (N_2067,In_573,In_2486);
nor U2068 (N_2068,In_1241,In_623);
and U2069 (N_2069,In_751,In_956);
nor U2070 (N_2070,In_1475,In_909);
xnor U2071 (N_2071,In_901,In_1232);
nand U2072 (N_2072,In_148,In_1097);
nor U2073 (N_2073,In_1343,In_1823);
and U2074 (N_2074,In_1414,In_1597);
nor U2075 (N_2075,In_1606,In_2007);
or U2076 (N_2076,In_2058,In_1683);
and U2077 (N_2077,In_2419,In_1282);
nand U2078 (N_2078,In_2065,In_1349);
nor U2079 (N_2079,In_160,In_2481);
xor U2080 (N_2080,In_1287,In_1753);
nand U2081 (N_2081,In_75,In_996);
xnor U2082 (N_2082,In_2298,In_1095);
and U2083 (N_2083,In_2028,In_1069);
nor U2084 (N_2084,In_1410,In_1235);
and U2085 (N_2085,In_1455,In_2233);
nor U2086 (N_2086,In_2124,In_2356);
nor U2087 (N_2087,In_1870,In_1951);
xnor U2088 (N_2088,In_0,In_371);
nand U2089 (N_2089,In_1227,In_1192);
nand U2090 (N_2090,In_911,In_1936);
nor U2091 (N_2091,In_118,In_2120);
and U2092 (N_2092,In_1233,In_1741);
and U2093 (N_2093,In_1980,In_1408);
xnor U2094 (N_2094,In_1500,In_844);
and U2095 (N_2095,In_500,In_1471);
nand U2096 (N_2096,In_127,In_1970);
and U2097 (N_2097,In_2013,In_2366);
or U2098 (N_2098,In_177,In_1912);
or U2099 (N_2099,In_1782,In_469);
and U2100 (N_2100,In_1780,In_1706);
or U2101 (N_2101,In_2316,In_2053);
and U2102 (N_2102,In_123,In_670);
xnor U2103 (N_2103,In_1184,In_1938);
nor U2104 (N_2104,In_2074,In_480);
nor U2105 (N_2105,In_330,In_1064);
xor U2106 (N_2106,In_264,In_978);
nand U2107 (N_2107,In_1109,In_1779);
or U2108 (N_2108,In_1930,In_980);
or U2109 (N_2109,In_1317,In_271);
or U2110 (N_2110,In_1468,In_1348);
and U2111 (N_2111,In_247,In_719);
nor U2112 (N_2112,In_250,In_1992);
nand U2113 (N_2113,In_1323,In_1113);
nand U2114 (N_2114,In_83,In_1228);
nand U2115 (N_2115,In_1375,In_2495);
nand U2116 (N_2116,In_662,In_1050);
and U2117 (N_2117,In_1372,In_677);
or U2118 (N_2118,In_1754,In_656);
and U2119 (N_2119,In_1857,In_2391);
nor U2120 (N_2120,In_452,In_2233);
nor U2121 (N_2121,In_2389,In_1645);
nand U2122 (N_2122,In_2175,In_813);
or U2123 (N_2123,In_58,In_1183);
or U2124 (N_2124,In_1440,In_1230);
or U2125 (N_2125,In_91,In_1336);
nand U2126 (N_2126,In_1954,In_1618);
nor U2127 (N_2127,In_157,In_1348);
and U2128 (N_2128,In_822,In_1817);
nor U2129 (N_2129,In_2269,In_2383);
or U2130 (N_2130,In_1284,In_2009);
and U2131 (N_2131,In_2383,In_1600);
or U2132 (N_2132,In_1747,In_361);
nor U2133 (N_2133,In_698,In_2198);
nor U2134 (N_2134,In_510,In_1009);
or U2135 (N_2135,In_1611,In_690);
or U2136 (N_2136,In_1859,In_762);
nand U2137 (N_2137,In_124,In_1454);
or U2138 (N_2138,In_2282,In_391);
nor U2139 (N_2139,In_2277,In_179);
and U2140 (N_2140,In_2280,In_1603);
xor U2141 (N_2141,In_1339,In_343);
nand U2142 (N_2142,In_174,In_1293);
xnor U2143 (N_2143,In_588,In_1562);
and U2144 (N_2144,In_2156,In_1392);
nand U2145 (N_2145,In_1807,In_1065);
and U2146 (N_2146,In_2444,In_1997);
nor U2147 (N_2147,In_1379,In_1932);
or U2148 (N_2148,In_1931,In_83);
nand U2149 (N_2149,In_1535,In_2185);
nor U2150 (N_2150,In_2283,In_2246);
and U2151 (N_2151,In_2008,In_1260);
xor U2152 (N_2152,In_2376,In_1135);
and U2153 (N_2153,In_734,In_304);
nand U2154 (N_2154,In_308,In_773);
and U2155 (N_2155,In_206,In_841);
nor U2156 (N_2156,In_260,In_1574);
nor U2157 (N_2157,In_2445,In_494);
nand U2158 (N_2158,In_1864,In_185);
nor U2159 (N_2159,In_1422,In_1934);
or U2160 (N_2160,In_1632,In_2328);
nand U2161 (N_2161,In_1295,In_1873);
nand U2162 (N_2162,In_1329,In_909);
or U2163 (N_2163,In_990,In_1336);
and U2164 (N_2164,In_887,In_856);
or U2165 (N_2165,In_1545,In_715);
or U2166 (N_2166,In_1163,In_64);
nor U2167 (N_2167,In_1660,In_1646);
or U2168 (N_2168,In_1996,In_1539);
and U2169 (N_2169,In_1607,In_1430);
and U2170 (N_2170,In_2167,In_235);
or U2171 (N_2171,In_412,In_548);
nand U2172 (N_2172,In_1259,In_2399);
and U2173 (N_2173,In_1788,In_1311);
nand U2174 (N_2174,In_2393,In_705);
nand U2175 (N_2175,In_2299,In_943);
nand U2176 (N_2176,In_547,In_1816);
or U2177 (N_2177,In_1423,In_858);
nor U2178 (N_2178,In_288,In_1063);
nand U2179 (N_2179,In_787,In_533);
or U2180 (N_2180,In_2145,In_2476);
and U2181 (N_2181,In_2331,In_1120);
or U2182 (N_2182,In_383,In_2483);
or U2183 (N_2183,In_1772,In_1114);
or U2184 (N_2184,In_834,In_642);
nor U2185 (N_2185,In_1696,In_548);
nor U2186 (N_2186,In_1819,In_1209);
or U2187 (N_2187,In_961,In_1246);
xor U2188 (N_2188,In_345,In_1289);
xor U2189 (N_2189,In_1843,In_2078);
nor U2190 (N_2190,In_392,In_1751);
and U2191 (N_2191,In_2018,In_2402);
and U2192 (N_2192,In_1295,In_1448);
nor U2193 (N_2193,In_1897,In_1389);
or U2194 (N_2194,In_1039,In_1122);
nand U2195 (N_2195,In_1594,In_513);
nor U2196 (N_2196,In_2352,In_2061);
and U2197 (N_2197,In_1850,In_1235);
xnor U2198 (N_2198,In_2,In_436);
and U2199 (N_2199,In_964,In_1144);
nor U2200 (N_2200,In_1823,In_2385);
or U2201 (N_2201,In_949,In_1511);
nor U2202 (N_2202,In_1913,In_1764);
nor U2203 (N_2203,In_599,In_1533);
xor U2204 (N_2204,In_1314,In_884);
and U2205 (N_2205,In_193,In_1430);
and U2206 (N_2206,In_1067,In_1138);
nand U2207 (N_2207,In_613,In_1442);
nor U2208 (N_2208,In_2138,In_1848);
or U2209 (N_2209,In_418,In_340);
and U2210 (N_2210,In_1279,In_2306);
xor U2211 (N_2211,In_1895,In_762);
or U2212 (N_2212,In_1491,In_193);
or U2213 (N_2213,In_2261,In_2170);
and U2214 (N_2214,In_700,In_867);
nor U2215 (N_2215,In_2151,In_247);
xor U2216 (N_2216,In_2003,In_1006);
nand U2217 (N_2217,In_601,In_550);
nand U2218 (N_2218,In_2130,In_1004);
xor U2219 (N_2219,In_2155,In_1555);
xor U2220 (N_2220,In_2167,In_2277);
nor U2221 (N_2221,In_604,In_930);
nor U2222 (N_2222,In_1013,In_1617);
or U2223 (N_2223,In_2417,In_1343);
nand U2224 (N_2224,In_1924,In_2149);
and U2225 (N_2225,In_1535,In_2498);
nand U2226 (N_2226,In_873,In_228);
nand U2227 (N_2227,In_389,In_618);
or U2228 (N_2228,In_1441,In_1757);
nand U2229 (N_2229,In_2381,In_187);
nand U2230 (N_2230,In_347,In_874);
or U2231 (N_2231,In_1894,In_1082);
nand U2232 (N_2232,In_2177,In_452);
xor U2233 (N_2233,In_1092,In_1893);
or U2234 (N_2234,In_32,In_138);
and U2235 (N_2235,In_1272,In_1025);
or U2236 (N_2236,In_1954,In_2148);
or U2237 (N_2237,In_1123,In_1744);
and U2238 (N_2238,In_1511,In_2314);
and U2239 (N_2239,In_2403,In_1511);
or U2240 (N_2240,In_2301,In_923);
nand U2241 (N_2241,In_2285,In_91);
and U2242 (N_2242,In_368,In_1270);
nor U2243 (N_2243,In_621,In_362);
or U2244 (N_2244,In_463,In_1916);
or U2245 (N_2245,In_493,In_955);
and U2246 (N_2246,In_1520,In_1042);
nand U2247 (N_2247,In_280,In_2306);
and U2248 (N_2248,In_1101,In_590);
nor U2249 (N_2249,In_1607,In_1994);
or U2250 (N_2250,In_1762,In_145);
or U2251 (N_2251,In_2456,In_2060);
nand U2252 (N_2252,In_2122,In_2302);
nand U2253 (N_2253,In_546,In_2335);
nor U2254 (N_2254,In_1940,In_50);
or U2255 (N_2255,In_358,In_1400);
nand U2256 (N_2256,In_1221,In_355);
and U2257 (N_2257,In_1922,In_1183);
or U2258 (N_2258,In_1410,In_2355);
nor U2259 (N_2259,In_1555,In_73);
nor U2260 (N_2260,In_1863,In_1922);
nor U2261 (N_2261,In_735,In_1934);
and U2262 (N_2262,In_2126,In_906);
xor U2263 (N_2263,In_246,In_1264);
nand U2264 (N_2264,In_516,In_2111);
nand U2265 (N_2265,In_1752,In_604);
nand U2266 (N_2266,In_2105,In_371);
nand U2267 (N_2267,In_156,In_879);
nor U2268 (N_2268,In_1376,In_386);
or U2269 (N_2269,In_906,In_1186);
or U2270 (N_2270,In_1426,In_2460);
and U2271 (N_2271,In_516,In_244);
or U2272 (N_2272,In_505,In_1225);
nor U2273 (N_2273,In_835,In_358);
or U2274 (N_2274,In_874,In_1378);
nor U2275 (N_2275,In_985,In_1100);
nand U2276 (N_2276,In_183,In_1233);
and U2277 (N_2277,In_699,In_1551);
nor U2278 (N_2278,In_746,In_253);
nor U2279 (N_2279,In_1635,In_736);
nor U2280 (N_2280,In_180,In_1672);
nand U2281 (N_2281,In_1508,In_882);
and U2282 (N_2282,In_2207,In_2061);
nand U2283 (N_2283,In_754,In_278);
or U2284 (N_2284,In_510,In_2491);
xor U2285 (N_2285,In_1892,In_1257);
and U2286 (N_2286,In_944,In_299);
nor U2287 (N_2287,In_1588,In_1141);
xor U2288 (N_2288,In_1251,In_2225);
nand U2289 (N_2289,In_284,In_1227);
nor U2290 (N_2290,In_764,In_492);
or U2291 (N_2291,In_847,In_2470);
nor U2292 (N_2292,In_710,In_44);
nor U2293 (N_2293,In_2107,In_271);
and U2294 (N_2294,In_1930,In_402);
or U2295 (N_2295,In_257,In_1027);
nand U2296 (N_2296,In_337,In_958);
xnor U2297 (N_2297,In_1715,In_916);
and U2298 (N_2298,In_2126,In_1369);
and U2299 (N_2299,In_1312,In_423);
or U2300 (N_2300,In_2307,In_1623);
or U2301 (N_2301,In_1628,In_1790);
or U2302 (N_2302,In_1980,In_1608);
nand U2303 (N_2303,In_2193,In_776);
nand U2304 (N_2304,In_1273,In_2378);
or U2305 (N_2305,In_1668,In_1798);
or U2306 (N_2306,In_1325,In_147);
nor U2307 (N_2307,In_2338,In_1355);
and U2308 (N_2308,In_594,In_1936);
or U2309 (N_2309,In_20,In_2478);
or U2310 (N_2310,In_1728,In_2496);
or U2311 (N_2311,In_571,In_1694);
and U2312 (N_2312,In_1133,In_1336);
nor U2313 (N_2313,In_1684,In_1515);
and U2314 (N_2314,In_1157,In_262);
or U2315 (N_2315,In_991,In_2432);
or U2316 (N_2316,In_1601,In_1119);
nor U2317 (N_2317,In_1423,In_1639);
and U2318 (N_2318,In_2188,In_1071);
and U2319 (N_2319,In_1308,In_557);
or U2320 (N_2320,In_1067,In_432);
or U2321 (N_2321,In_1567,In_2459);
or U2322 (N_2322,In_1922,In_1889);
or U2323 (N_2323,In_2302,In_550);
nor U2324 (N_2324,In_1643,In_742);
or U2325 (N_2325,In_1112,In_1491);
nor U2326 (N_2326,In_1561,In_1250);
or U2327 (N_2327,In_1211,In_1945);
nand U2328 (N_2328,In_2189,In_1267);
nand U2329 (N_2329,In_1028,In_1875);
nor U2330 (N_2330,In_1210,In_1222);
nand U2331 (N_2331,In_358,In_336);
nor U2332 (N_2332,In_164,In_2380);
nor U2333 (N_2333,In_1842,In_1202);
xor U2334 (N_2334,In_971,In_158);
nor U2335 (N_2335,In_1436,In_578);
and U2336 (N_2336,In_139,In_1187);
nor U2337 (N_2337,In_1832,In_1667);
nand U2338 (N_2338,In_2167,In_510);
nor U2339 (N_2339,In_1645,In_1830);
nor U2340 (N_2340,In_1188,In_1414);
xnor U2341 (N_2341,In_624,In_1762);
xor U2342 (N_2342,In_1821,In_1174);
xor U2343 (N_2343,In_814,In_1659);
and U2344 (N_2344,In_0,In_1513);
nor U2345 (N_2345,In_1538,In_479);
xnor U2346 (N_2346,In_2034,In_1511);
nor U2347 (N_2347,In_439,In_709);
nand U2348 (N_2348,In_1874,In_770);
xnor U2349 (N_2349,In_1351,In_1323);
xnor U2350 (N_2350,In_503,In_1369);
nor U2351 (N_2351,In_1857,In_2123);
xor U2352 (N_2352,In_115,In_470);
nand U2353 (N_2353,In_2374,In_1199);
xnor U2354 (N_2354,In_1050,In_1237);
xor U2355 (N_2355,In_51,In_1387);
nor U2356 (N_2356,In_856,In_63);
xor U2357 (N_2357,In_2098,In_286);
and U2358 (N_2358,In_2210,In_1542);
nor U2359 (N_2359,In_1073,In_1363);
or U2360 (N_2360,In_863,In_864);
or U2361 (N_2361,In_1981,In_2341);
nor U2362 (N_2362,In_2069,In_923);
xnor U2363 (N_2363,In_1793,In_1359);
nor U2364 (N_2364,In_475,In_324);
or U2365 (N_2365,In_1857,In_2366);
and U2366 (N_2366,In_756,In_798);
or U2367 (N_2367,In_1349,In_2215);
and U2368 (N_2368,In_327,In_808);
or U2369 (N_2369,In_1092,In_1890);
nor U2370 (N_2370,In_2397,In_1639);
nand U2371 (N_2371,In_1128,In_1339);
nand U2372 (N_2372,In_1934,In_298);
and U2373 (N_2373,In_1076,In_677);
nand U2374 (N_2374,In_688,In_916);
nor U2375 (N_2375,In_86,In_1645);
and U2376 (N_2376,In_583,In_2017);
nand U2377 (N_2377,In_360,In_2036);
nand U2378 (N_2378,In_2452,In_2058);
nor U2379 (N_2379,In_2249,In_354);
or U2380 (N_2380,In_607,In_207);
nor U2381 (N_2381,In_1222,In_2483);
nor U2382 (N_2382,In_1668,In_272);
nand U2383 (N_2383,In_2049,In_1898);
nor U2384 (N_2384,In_2349,In_1909);
or U2385 (N_2385,In_14,In_0);
xor U2386 (N_2386,In_1048,In_1438);
nor U2387 (N_2387,In_1857,In_2081);
xor U2388 (N_2388,In_91,In_1213);
or U2389 (N_2389,In_1044,In_1798);
nand U2390 (N_2390,In_2176,In_318);
or U2391 (N_2391,In_1340,In_2308);
xor U2392 (N_2392,In_582,In_2463);
and U2393 (N_2393,In_2407,In_1469);
and U2394 (N_2394,In_771,In_2054);
nand U2395 (N_2395,In_2208,In_1534);
nand U2396 (N_2396,In_2344,In_993);
nor U2397 (N_2397,In_1757,In_1351);
or U2398 (N_2398,In_710,In_1079);
nor U2399 (N_2399,In_300,In_2095);
xnor U2400 (N_2400,In_1998,In_1496);
and U2401 (N_2401,In_761,In_2229);
nand U2402 (N_2402,In_1620,In_933);
or U2403 (N_2403,In_1390,In_2254);
nor U2404 (N_2404,In_1126,In_429);
nand U2405 (N_2405,In_542,In_736);
nor U2406 (N_2406,In_997,In_1752);
xnor U2407 (N_2407,In_1900,In_822);
xnor U2408 (N_2408,In_2345,In_770);
and U2409 (N_2409,In_2227,In_2051);
and U2410 (N_2410,In_926,In_838);
and U2411 (N_2411,In_2232,In_962);
nand U2412 (N_2412,In_2034,In_1893);
nor U2413 (N_2413,In_1912,In_1112);
or U2414 (N_2414,In_116,In_73);
and U2415 (N_2415,In_150,In_47);
nor U2416 (N_2416,In_1619,In_2106);
xnor U2417 (N_2417,In_809,In_1948);
nand U2418 (N_2418,In_2405,In_246);
nand U2419 (N_2419,In_551,In_2231);
or U2420 (N_2420,In_1334,In_2035);
xnor U2421 (N_2421,In_63,In_1830);
xor U2422 (N_2422,In_8,In_1392);
or U2423 (N_2423,In_2464,In_508);
or U2424 (N_2424,In_1894,In_417);
nand U2425 (N_2425,In_2356,In_373);
nor U2426 (N_2426,In_2472,In_1683);
and U2427 (N_2427,In_602,In_2400);
nand U2428 (N_2428,In_1880,In_909);
or U2429 (N_2429,In_246,In_1017);
or U2430 (N_2430,In_2207,In_2349);
xor U2431 (N_2431,In_315,In_666);
or U2432 (N_2432,In_766,In_214);
nor U2433 (N_2433,In_884,In_642);
or U2434 (N_2434,In_2261,In_1836);
or U2435 (N_2435,In_1926,In_1271);
nor U2436 (N_2436,In_2021,In_1614);
nand U2437 (N_2437,In_44,In_1680);
and U2438 (N_2438,In_1958,In_1157);
and U2439 (N_2439,In_504,In_1334);
or U2440 (N_2440,In_2141,In_1984);
and U2441 (N_2441,In_58,In_73);
nor U2442 (N_2442,In_2421,In_361);
or U2443 (N_2443,In_1017,In_183);
or U2444 (N_2444,In_1470,In_1477);
nand U2445 (N_2445,In_1111,In_91);
nor U2446 (N_2446,In_1881,In_449);
nor U2447 (N_2447,In_1202,In_92);
and U2448 (N_2448,In_1393,In_685);
or U2449 (N_2449,In_1662,In_576);
nor U2450 (N_2450,In_213,In_1687);
nor U2451 (N_2451,In_1047,In_868);
nor U2452 (N_2452,In_1800,In_2464);
nor U2453 (N_2453,In_466,In_1457);
nand U2454 (N_2454,In_1357,In_1139);
nand U2455 (N_2455,In_609,In_2077);
nor U2456 (N_2456,In_226,In_868);
nor U2457 (N_2457,In_2062,In_1618);
nand U2458 (N_2458,In_2482,In_1368);
and U2459 (N_2459,In_2030,In_2010);
or U2460 (N_2460,In_562,In_2383);
nor U2461 (N_2461,In_1998,In_1278);
or U2462 (N_2462,In_17,In_665);
nor U2463 (N_2463,In_1362,In_1913);
nand U2464 (N_2464,In_1565,In_558);
xor U2465 (N_2465,In_1698,In_955);
and U2466 (N_2466,In_2202,In_310);
or U2467 (N_2467,In_1036,In_1975);
nand U2468 (N_2468,In_351,In_135);
and U2469 (N_2469,In_1332,In_1137);
xnor U2470 (N_2470,In_2048,In_1811);
and U2471 (N_2471,In_2282,In_1302);
xnor U2472 (N_2472,In_620,In_1596);
or U2473 (N_2473,In_1513,In_687);
or U2474 (N_2474,In_1155,In_1834);
or U2475 (N_2475,In_2314,In_934);
xnor U2476 (N_2476,In_2141,In_1988);
and U2477 (N_2477,In_1846,In_1339);
nor U2478 (N_2478,In_2329,In_514);
nand U2479 (N_2479,In_410,In_1567);
xor U2480 (N_2480,In_2299,In_918);
xor U2481 (N_2481,In_659,In_566);
and U2482 (N_2482,In_964,In_1826);
nand U2483 (N_2483,In_270,In_1335);
or U2484 (N_2484,In_1256,In_432);
nor U2485 (N_2485,In_1108,In_746);
nor U2486 (N_2486,In_2319,In_409);
xor U2487 (N_2487,In_1899,In_1248);
or U2488 (N_2488,In_1972,In_5);
or U2489 (N_2489,In_2497,In_1198);
xnor U2490 (N_2490,In_2285,In_1427);
nand U2491 (N_2491,In_2338,In_20);
or U2492 (N_2492,In_2484,In_416);
nand U2493 (N_2493,In_2232,In_1799);
nand U2494 (N_2494,In_1768,In_610);
or U2495 (N_2495,In_1024,In_1271);
xnor U2496 (N_2496,In_2354,In_1392);
or U2497 (N_2497,In_2499,In_2351);
xnor U2498 (N_2498,In_1039,In_2037);
or U2499 (N_2499,In_53,In_1593);
nand U2500 (N_2500,In_1198,In_73);
xnor U2501 (N_2501,In_37,In_802);
or U2502 (N_2502,In_2255,In_1291);
and U2503 (N_2503,In_1207,In_855);
nor U2504 (N_2504,In_2046,In_1500);
nor U2505 (N_2505,In_2371,In_1570);
or U2506 (N_2506,In_48,In_2430);
or U2507 (N_2507,In_2438,In_1945);
or U2508 (N_2508,In_2097,In_389);
xnor U2509 (N_2509,In_2482,In_791);
nor U2510 (N_2510,In_1866,In_416);
or U2511 (N_2511,In_453,In_968);
and U2512 (N_2512,In_776,In_2189);
nor U2513 (N_2513,In_121,In_1078);
nand U2514 (N_2514,In_1737,In_2250);
or U2515 (N_2515,In_2264,In_885);
nor U2516 (N_2516,In_2117,In_1540);
xnor U2517 (N_2517,In_150,In_2288);
and U2518 (N_2518,In_1543,In_1744);
xor U2519 (N_2519,In_945,In_521);
nand U2520 (N_2520,In_1395,In_624);
or U2521 (N_2521,In_2428,In_753);
nor U2522 (N_2522,In_1075,In_2007);
and U2523 (N_2523,In_1721,In_2260);
nand U2524 (N_2524,In_1299,In_254);
nand U2525 (N_2525,In_67,In_1891);
or U2526 (N_2526,In_1092,In_2226);
or U2527 (N_2527,In_282,In_1254);
or U2528 (N_2528,In_374,In_167);
nor U2529 (N_2529,In_124,In_893);
and U2530 (N_2530,In_1211,In_476);
nor U2531 (N_2531,In_2457,In_935);
and U2532 (N_2532,In_1209,In_2461);
or U2533 (N_2533,In_2448,In_1662);
or U2534 (N_2534,In_2196,In_1296);
or U2535 (N_2535,In_303,In_753);
or U2536 (N_2536,In_2368,In_2286);
and U2537 (N_2537,In_1445,In_382);
or U2538 (N_2538,In_563,In_1543);
and U2539 (N_2539,In_2302,In_2305);
and U2540 (N_2540,In_227,In_2305);
nand U2541 (N_2541,In_2157,In_144);
and U2542 (N_2542,In_1997,In_2198);
nor U2543 (N_2543,In_2340,In_1917);
nor U2544 (N_2544,In_266,In_278);
nand U2545 (N_2545,In_2421,In_1291);
nor U2546 (N_2546,In_2494,In_2281);
and U2547 (N_2547,In_1412,In_1727);
xor U2548 (N_2548,In_682,In_712);
or U2549 (N_2549,In_1923,In_2474);
nor U2550 (N_2550,In_1121,In_116);
or U2551 (N_2551,In_625,In_1357);
xor U2552 (N_2552,In_2223,In_2167);
nand U2553 (N_2553,In_2344,In_1022);
nor U2554 (N_2554,In_2379,In_2312);
nor U2555 (N_2555,In_62,In_33);
or U2556 (N_2556,In_2071,In_688);
and U2557 (N_2557,In_2130,In_2160);
or U2558 (N_2558,In_2144,In_2072);
nand U2559 (N_2559,In_956,In_252);
nand U2560 (N_2560,In_103,In_991);
nand U2561 (N_2561,In_2455,In_1605);
or U2562 (N_2562,In_1008,In_611);
and U2563 (N_2563,In_853,In_2147);
or U2564 (N_2564,In_176,In_1574);
and U2565 (N_2565,In_1095,In_1513);
nor U2566 (N_2566,In_1004,In_2360);
and U2567 (N_2567,In_1243,In_2397);
and U2568 (N_2568,In_1555,In_296);
and U2569 (N_2569,In_1457,In_192);
nor U2570 (N_2570,In_795,In_590);
or U2571 (N_2571,In_64,In_890);
nor U2572 (N_2572,In_2354,In_1171);
or U2573 (N_2573,In_32,In_721);
and U2574 (N_2574,In_769,In_1315);
nor U2575 (N_2575,In_1272,In_2404);
nor U2576 (N_2576,In_1509,In_1707);
xor U2577 (N_2577,In_2056,In_368);
or U2578 (N_2578,In_1021,In_1149);
and U2579 (N_2579,In_2005,In_1685);
nor U2580 (N_2580,In_1122,In_1179);
or U2581 (N_2581,In_908,In_1462);
or U2582 (N_2582,In_1017,In_986);
nand U2583 (N_2583,In_1842,In_2053);
or U2584 (N_2584,In_1403,In_1491);
xnor U2585 (N_2585,In_1047,In_139);
nand U2586 (N_2586,In_886,In_1462);
nor U2587 (N_2587,In_2446,In_450);
nand U2588 (N_2588,In_1231,In_130);
and U2589 (N_2589,In_1637,In_335);
and U2590 (N_2590,In_936,In_2166);
xor U2591 (N_2591,In_831,In_1757);
and U2592 (N_2592,In_1959,In_345);
or U2593 (N_2593,In_955,In_678);
nor U2594 (N_2594,In_1380,In_596);
and U2595 (N_2595,In_2230,In_1901);
or U2596 (N_2596,In_1572,In_2151);
and U2597 (N_2597,In_554,In_1208);
nand U2598 (N_2598,In_232,In_1463);
nor U2599 (N_2599,In_1047,In_2433);
nor U2600 (N_2600,In_186,In_333);
and U2601 (N_2601,In_493,In_669);
or U2602 (N_2602,In_2171,In_2446);
and U2603 (N_2603,In_1252,In_319);
nor U2604 (N_2604,In_402,In_229);
or U2605 (N_2605,In_654,In_1053);
and U2606 (N_2606,In_2307,In_1269);
xnor U2607 (N_2607,In_889,In_1181);
and U2608 (N_2608,In_1553,In_1309);
nor U2609 (N_2609,In_1952,In_200);
nor U2610 (N_2610,In_1293,In_687);
or U2611 (N_2611,In_1839,In_350);
or U2612 (N_2612,In_929,In_2229);
nand U2613 (N_2613,In_733,In_844);
and U2614 (N_2614,In_793,In_121);
or U2615 (N_2615,In_841,In_1948);
nand U2616 (N_2616,In_766,In_1865);
nor U2617 (N_2617,In_1392,In_1768);
and U2618 (N_2618,In_186,In_1136);
nand U2619 (N_2619,In_334,In_218);
or U2620 (N_2620,In_1444,In_1450);
nor U2621 (N_2621,In_327,In_1763);
or U2622 (N_2622,In_1091,In_1438);
nand U2623 (N_2623,In_745,In_960);
nand U2624 (N_2624,In_845,In_2208);
and U2625 (N_2625,In_1135,In_274);
and U2626 (N_2626,In_563,In_1976);
or U2627 (N_2627,In_536,In_1496);
nand U2628 (N_2628,In_889,In_2236);
xor U2629 (N_2629,In_2164,In_859);
or U2630 (N_2630,In_876,In_1746);
nand U2631 (N_2631,In_1254,In_1185);
nor U2632 (N_2632,In_1476,In_430);
nand U2633 (N_2633,In_125,In_28);
or U2634 (N_2634,In_1635,In_1226);
nand U2635 (N_2635,In_388,In_2300);
or U2636 (N_2636,In_181,In_2425);
nor U2637 (N_2637,In_1473,In_1764);
and U2638 (N_2638,In_627,In_805);
and U2639 (N_2639,In_284,In_420);
nor U2640 (N_2640,In_2280,In_627);
or U2641 (N_2641,In_1057,In_2326);
nand U2642 (N_2642,In_1884,In_1917);
nand U2643 (N_2643,In_922,In_1164);
nor U2644 (N_2644,In_2455,In_2471);
or U2645 (N_2645,In_677,In_1989);
nor U2646 (N_2646,In_2302,In_1783);
nand U2647 (N_2647,In_1769,In_2038);
or U2648 (N_2648,In_97,In_1213);
nand U2649 (N_2649,In_731,In_258);
nor U2650 (N_2650,In_1865,In_253);
nor U2651 (N_2651,In_1537,In_2343);
nor U2652 (N_2652,In_626,In_1019);
nor U2653 (N_2653,In_1384,In_1411);
and U2654 (N_2654,In_454,In_934);
nor U2655 (N_2655,In_32,In_1357);
nand U2656 (N_2656,In_1815,In_2123);
and U2657 (N_2657,In_1666,In_1493);
nand U2658 (N_2658,In_451,In_692);
or U2659 (N_2659,In_1242,In_57);
nor U2660 (N_2660,In_402,In_1660);
nor U2661 (N_2661,In_2109,In_135);
nor U2662 (N_2662,In_490,In_205);
and U2663 (N_2663,In_1242,In_2479);
nand U2664 (N_2664,In_2282,In_2021);
nand U2665 (N_2665,In_589,In_2057);
xor U2666 (N_2666,In_646,In_1709);
or U2667 (N_2667,In_296,In_1741);
or U2668 (N_2668,In_726,In_895);
or U2669 (N_2669,In_150,In_2247);
nor U2670 (N_2670,In_1417,In_2014);
or U2671 (N_2671,In_2443,In_2225);
and U2672 (N_2672,In_980,In_2053);
nor U2673 (N_2673,In_503,In_1215);
or U2674 (N_2674,In_529,In_1668);
nand U2675 (N_2675,In_1199,In_88);
nor U2676 (N_2676,In_248,In_934);
xor U2677 (N_2677,In_1101,In_1146);
nand U2678 (N_2678,In_289,In_695);
nor U2679 (N_2679,In_1147,In_1014);
and U2680 (N_2680,In_210,In_1881);
nor U2681 (N_2681,In_189,In_461);
or U2682 (N_2682,In_2004,In_768);
or U2683 (N_2683,In_708,In_1959);
or U2684 (N_2684,In_2377,In_1151);
and U2685 (N_2685,In_1464,In_424);
nand U2686 (N_2686,In_475,In_1434);
nor U2687 (N_2687,In_882,In_1489);
nor U2688 (N_2688,In_163,In_1244);
or U2689 (N_2689,In_2280,In_966);
or U2690 (N_2690,In_262,In_612);
or U2691 (N_2691,In_1926,In_405);
nand U2692 (N_2692,In_2190,In_2416);
nor U2693 (N_2693,In_1816,In_1024);
nor U2694 (N_2694,In_936,In_74);
nand U2695 (N_2695,In_2294,In_515);
or U2696 (N_2696,In_1021,In_1684);
nand U2697 (N_2697,In_436,In_1417);
and U2698 (N_2698,In_1725,In_1074);
and U2699 (N_2699,In_1600,In_1987);
or U2700 (N_2700,In_336,In_1771);
nor U2701 (N_2701,In_1384,In_859);
nor U2702 (N_2702,In_942,In_1292);
or U2703 (N_2703,In_161,In_1665);
nand U2704 (N_2704,In_834,In_372);
or U2705 (N_2705,In_580,In_558);
and U2706 (N_2706,In_1002,In_2152);
nor U2707 (N_2707,In_770,In_564);
and U2708 (N_2708,In_1589,In_628);
or U2709 (N_2709,In_837,In_693);
nor U2710 (N_2710,In_541,In_272);
and U2711 (N_2711,In_1552,In_151);
and U2712 (N_2712,In_620,In_2479);
and U2713 (N_2713,In_354,In_165);
or U2714 (N_2714,In_504,In_633);
or U2715 (N_2715,In_607,In_796);
nand U2716 (N_2716,In_2315,In_738);
xor U2717 (N_2717,In_1399,In_149);
nand U2718 (N_2718,In_425,In_2299);
or U2719 (N_2719,In_2313,In_1401);
and U2720 (N_2720,In_1565,In_1860);
xor U2721 (N_2721,In_2054,In_973);
nand U2722 (N_2722,In_880,In_1422);
nor U2723 (N_2723,In_15,In_1584);
and U2724 (N_2724,In_1544,In_384);
nand U2725 (N_2725,In_2200,In_1318);
and U2726 (N_2726,In_320,In_759);
nand U2727 (N_2727,In_1710,In_1781);
and U2728 (N_2728,In_2304,In_406);
nor U2729 (N_2729,In_339,In_597);
nand U2730 (N_2730,In_2407,In_1084);
or U2731 (N_2731,In_2087,In_488);
xnor U2732 (N_2732,In_64,In_638);
nor U2733 (N_2733,In_548,In_872);
and U2734 (N_2734,In_739,In_1402);
nor U2735 (N_2735,In_1132,In_2181);
or U2736 (N_2736,In_393,In_1234);
and U2737 (N_2737,In_2196,In_800);
and U2738 (N_2738,In_845,In_1047);
xor U2739 (N_2739,In_1244,In_2245);
xnor U2740 (N_2740,In_101,In_626);
xnor U2741 (N_2741,In_871,In_1896);
and U2742 (N_2742,In_1667,In_735);
nor U2743 (N_2743,In_793,In_875);
or U2744 (N_2744,In_1865,In_141);
or U2745 (N_2745,In_396,In_1047);
xor U2746 (N_2746,In_1879,In_296);
or U2747 (N_2747,In_751,In_740);
xor U2748 (N_2748,In_1786,In_1522);
or U2749 (N_2749,In_816,In_1093);
and U2750 (N_2750,In_960,In_2162);
nor U2751 (N_2751,In_303,In_838);
nand U2752 (N_2752,In_469,In_1609);
nand U2753 (N_2753,In_520,In_1344);
nand U2754 (N_2754,In_1359,In_612);
nor U2755 (N_2755,In_250,In_2037);
nor U2756 (N_2756,In_1844,In_780);
nand U2757 (N_2757,In_583,In_2246);
nor U2758 (N_2758,In_93,In_1373);
nand U2759 (N_2759,In_747,In_1241);
nor U2760 (N_2760,In_773,In_1259);
nor U2761 (N_2761,In_154,In_1475);
nand U2762 (N_2762,In_1309,In_221);
nand U2763 (N_2763,In_1156,In_986);
or U2764 (N_2764,In_1856,In_58);
nand U2765 (N_2765,In_1776,In_1164);
nand U2766 (N_2766,In_795,In_899);
or U2767 (N_2767,In_1496,In_2392);
nor U2768 (N_2768,In_83,In_2175);
nor U2769 (N_2769,In_146,In_375);
nand U2770 (N_2770,In_1595,In_2195);
nor U2771 (N_2771,In_2083,In_477);
or U2772 (N_2772,In_832,In_1360);
nand U2773 (N_2773,In_1380,In_517);
nor U2774 (N_2774,In_2295,In_266);
and U2775 (N_2775,In_2035,In_1106);
and U2776 (N_2776,In_214,In_514);
and U2777 (N_2777,In_1292,In_1973);
nor U2778 (N_2778,In_1187,In_113);
xnor U2779 (N_2779,In_1330,In_217);
xnor U2780 (N_2780,In_1345,In_552);
nand U2781 (N_2781,In_383,In_1775);
or U2782 (N_2782,In_1871,In_150);
and U2783 (N_2783,In_35,In_1233);
and U2784 (N_2784,In_2420,In_895);
and U2785 (N_2785,In_119,In_2064);
or U2786 (N_2786,In_1363,In_1039);
nor U2787 (N_2787,In_1369,In_2196);
nor U2788 (N_2788,In_2051,In_264);
nor U2789 (N_2789,In_293,In_2319);
nor U2790 (N_2790,In_2095,In_1234);
nand U2791 (N_2791,In_2010,In_1235);
or U2792 (N_2792,In_1913,In_289);
nand U2793 (N_2793,In_1519,In_405);
nor U2794 (N_2794,In_1434,In_181);
nand U2795 (N_2795,In_2347,In_760);
or U2796 (N_2796,In_1619,In_271);
nor U2797 (N_2797,In_630,In_546);
and U2798 (N_2798,In_1944,In_2378);
xnor U2799 (N_2799,In_1691,In_2353);
nor U2800 (N_2800,In_1430,In_840);
and U2801 (N_2801,In_963,In_1142);
xor U2802 (N_2802,In_428,In_1358);
and U2803 (N_2803,In_2415,In_1677);
xor U2804 (N_2804,In_1985,In_1649);
xnor U2805 (N_2805,In_2405,In_200);
xor U2806 (N_2806,In_509,In_1674);
nand U2807 (N_2807,In_1798,In_1347);
and U2808 (N_2808,In_1357,In_540);
nor U2809 (N_2809,In_1936,In_386);
and U2810 (N_2810,In_1153,In_1019);
or U2811 (N_2811,In_1303,In_719);
or U2812 (N_2812,In_1122,In_234);
and U2813 (N_2813,In_642,In_2124);
nand U2814 (N_2814,In_269,In_507);
nor U2815 (N_2815,In_384,In_932);
and U2816 (N_2816,In_843,In_1869);
or U2817 (N_2817,In_2404,In_1977);
nand U2818 (N_2818,In_1238,In_2218);
or U2819 (N_2819,In_1803,In_616);
nand U2820 (N_2820,In_145,In_1799);
or U2821 (N_2821,In_1676,In_212);
and U2822 (N_2822,In_2038,In_1843);
nand U2823 (N_2823,In_481,In_406);
nand U2824 (N_2824,In_1090,In_1647);
nor U2825 (N_2825,In_1042,In_1215);
and U2826 (N_2826,In_498,In_441);
and U2827 (N_2827,In_2242,In_1578);
or U2828 (N_2828,In_28,In_2378);
and U2829 (N_2829,In_2359,In_526);
nand U2830 (N_2830,In_1515,In_2216);
nand U2831 (N_2831,In_250,In_2412);
nor U2832 (N_2832,In_83,In_1708);
or U2833 (N_2833,In_650,In_2300);
nand U2834 (N_2834,In_1730,In_1754);
nand U2835 (N_2835,In_103,In_1335);
or U2836 (N_2836,In_420,In_496);
nor U2837 (N_2837,In_916,In_609);
nand U2838 (N_2838,In_2284,In_1223);
or U2839 (N_2839,In_533,In_255);
and U2840 (N_2840,In_2251,In_2457);
and U2841 (N_2841,In_884,In_1716);
or U2842 (N_2842,In_1952,In_505);
or U2843 (N_2843,In_553,In_448);
nor U2844 (N_2844,In_2294,In_1277);
nor U2845 (N_2845,In_1671,In_2122);
nand U2846 (N_2846,In_1888,In_1008);
nand U2847 (N_2847,In_480,In_888);
nor U2848 (N_2848,In_1540,In_169);
or U2849 (N_2849,In_194,In_1986);
and U2850 (N_2850,In_383,In_1914);
or U2851 (N_2851,In_1676,In_1243);
or U2852 (N_2852,In_761,In_1522);
and U2853 (N_2853,In_443,In_2050);
xor U2854 (N_2854,In_2089,In_89);
xnor U2855 (N_2855,In_708,In_1410);
nor U2856 (N_2856,In_33,In_1176);
nand U2857 (N_2857,In_1610,In_959);
and U2858 (N_2858,In_519,In_1039);
nor U2859 (N_2859,In_466,In_1049);
and U2860 (N_2860,In_1358,In_1737);
nor U2861 (N_2861,In_2134,In_2347);
and U2862 (N_2862,In_1828,In_994);
or U2863 (N_2863,In_209,In_1698);
and U2864 (N_2864,In_1583,In_1651);
or U2865 (N_2865,In_1629,In_474);
nor U2866 (N_2866,In_394,In_1457);
or U2867 (N_2867,In_2467,In_2276);
nand U2868 (N_2868,In_1684,In_441);
and U2869 (N_2869,In_115,In_1352);
or U2870 (N_2870,In_265,In_2219);
nand U2871 (N_2871,In_1298,In_325);
and U2872 (N_2872,In_1407,In_73);
or U2873 (N_2873,In_1034,In_388);
nor U2874 (N_2874,In_2096,In_156);
nor U2875 (N_2875,In_1563,In_1261);
or U2876 (N_2876,In_649,In_763);
and U2877 (N_2877,In_1680,In_1232);
nor U2878 (N_2878,In_1371,In_2385);
or U2879 (N_2879,In_18,In_1796);
nand U2880 (N_2880,In_1815,In_1214);
and U2881 (N_2881,In_2027,In_2165);
xor U2882 (N_2882,In_2074,In_2488);
nor U2883 (N_2883,In_2348,In_869);
nor U2884 (N_2884,In_2360,In_1218);
or U2885 (N_2885,In_1804,In_1559);
nand U2886 (N_2886,In_1191,In_621);
and U2887 (N_2887,In_2342,In_1637);
or U2888 (N_2888,In_76,In_1524);
or U2889 (N_2889,In_1012,In_885);
or U2890 (N_2890,In_924,In_1256);
or U2891 (N_2891,In_1511,In_2242);
or U2892 (N_2892,In_1916,In_1913);
or U2893 (N_2893,In_757,In_2060);
nor U2894 (N_2894,In_1745,In_2034);
or U2895 (N_2895,In_1923,In_2104);
xnor U2896 (N_2896,In_1430,In_1174);
nand U2897 (N_2897,In_654,In_1317);
nor U2898 (N_2898,In_1323,In_2017);
or U2899 (N_2899,In_1671,In_122);
nand U2900 (N_2900,In_364,In_1901);
or U2901 (N_2901,In_1821,In_2102);
and U2902 (N_2902,In_2499,In_84);
or U2903 (N_2903,In_1765,In_1510);
nand U2904 (N_2904,In_992,In_1867);
and U2905 (N_2905,In_442,In_2109);
nand U2906 (N_2906,In_2153,In_1895);
xnor U2907 (N_2907,In_1228,In_314);
xnor U2908 (N_2908,In_1686,In_20);
or U2909 (N_2909,In_2495,In_2044);
nand U2910 (N_2910,In_2005,In_1284);
and U2911 (N_2911,In_1067,In_51);
and U2912 (N_2912,In_213,In_2461);
xnor U2913 (N_2913,In_971,In_82);
and U2914 (N_2914,In_2047,In_1583);
xor U2915 (N_2915,In_966,In_1514);
nand U2916 (N_2916,In_1668,In_238);
xor U2917 (N_2917,In_2000,In_1396);
nand U2918 (N_2918,In_1842,In_277);
nand U2919 (N_2919,In_1733,In_189);
nand U2920 (N_2920,In_1221,In_89);
and U2921 (N_2921,In_2380,In_1737);
nand U2922 (N_2922,In_477,In_1040);
or U2923 (N_2923,In_371,In_651);
nand U2924 (N_2924,In_1620,In_1894);
nor U2925 (N_2925,In_310,In_1727);
nand U2926 (N_2926,In_1018,In_541);
xor U2927 (N_2927,In_1913,In_868);
or U2928 (N_2928,In_131,In_1081);
nand U2929 (N_2929,In_306,In_435);
xor U2930 (N_2930,In_1955,In_1239);
and U2931 (N_2931,In_635,In_405);
or U2932 (N_2932,In_93,In_1453);
xor U2933 (N_2933,In_1687,In_914);
or U2934 (N_2934,In_1581,In_1021);
and U2935 (N_2935,In_1344,In_914);
or U2936 (N_2936,In_160,In_532);
nor U2937 (N_2937,In_1266,In_951);
and U2938 (N_2938,In_586,In_1218);
and U2939 (N_2939,In_1088,In_1146);
or U2940 (N_2940,In_146,In_1889);
or U2941 (N_2941,In_904,In_205);
nand U2942 (N_2942,In_1615,In_2419);
or U2943 (N_2943,In_1003,In_148);
or U2944 (N_2944,In_2432,In_816);
and U2945 (N_2945,In_1993,In_209);
nor U2946 (N_2946,In_293,In_2342);
nand U2947 (N_2947,In_562,In_336);
xnor U2948 (N_2948,In_2229,In_649);
and U2949 (N_2949,In_2430,In_1131);
nor U2950 (N_2950,In_1140,In_2379);
xor U2951 (N_2951,In_1148,In_2211);
and U2952 (N_2952,In_1655,In_1874);
or U2953 (N_2953,In_534,In_2247);
and U2954 (N_2954,In_1266,In_573);
or U2955 (N_2955,In_960,In_8);
nand U2956 (N_2956,In_2392,In_1642);
nand U2957 (N_2957,In_938,In_1671);
or U2958 (N_2958,In_942,In_1920);
nor U2959 (N_2959,In_343,In_1311);
or U2960 (N_2960,In_2415,In_1375);
nand U2961 (N_2961,In_2434,In_2384);
and U2962 (N_2962,In_966,In_651);
nand U2963 (N_2963,In_332,In_1842);
nand U2964 (N_2964,In_1024,In_566);
and U2965 (N_2965,In_2401,In_1149);
xnor U2966 (N_2966,In_1645,In_1079);
xnor U2967 (N_2967,In_2064,In_757);
or U2968 (N_2968,In_284,In_1137);
nor U2969 (N_2969,In_494,In_1259);
xnor U2970 (N_2970,In_1402,In_714);
and U2971 (N_2971,In_120,In_2467);
nor U2972 (N_2972,In_2325,In_113);
xor U2973 (N_2973,In_113,In_1712);
nor U2974 (N_2974,In_1439,In_1486);
and U2975 (N_2975,In_2377,In_1514);
nor U2976 (N_2976,In_942,In_1788);
and U2977 (N_2977,In_1154,In_1847);
nand U2978 (N_2978,In_955,In_1601);
or U2979 (N_2979,In_2400,In_711);
nand U2980 (N_2980,In_1970,In_137);
or U2981 (N_2981,In_659,In_2247);
and U2982 (N_2982,In_2248,In_2122);
nand U2983 (N_2983,In_1198,In_1479);
or U2984 (N_2984,In_1325,In_1525);
xor U2985 (N_2985,In_2078,In_286);
nor U2986 (N_2986,In_2021,In_1825);
xnor U2987 (N_2987,In_643,In_831);
and U2988 (N_2988,In_24,In_2224);
xor U2989 (N_2989,In_827,In_1391);
nand U2990 (N_2990,In_1185,In_1114);
or U2991 (N_2991,In_2094,In_420);
or U2992 (N_2992,In_1125,In_806);
or U2993 (N_2993,In_874,In_1041);
xnor U2994 (N_2994,In_2213,In_1051);
nor U2995 (N_2995,In_1214,In_1568);
nand U2996 (N_2996,In_517,In_2174);
and U2997 (N_2997,In_469,In_1908);
or U2998 (N_2998,In_1360,In_267);
xor U2999 (N_2999,In_96,In_521);
nand U3000 (N_3000,In_1261,In_1133);
and U3001 (N_3001,In_920,In_2304);
nand U3002 (N_3002,In_998,In_2265);
nor U3003 (N_3003,In_2016,In_756);
nor U3004 (N_3004,In_1007,In_2469);
xnor U3005 (N_3005,In_455,In_2174);
and U3006 (N_3006,In_2298,In_2195);
nor U3007 (N_3007,In_297,In_339);
and U3008 (N_3008,In_1608,In_857);
and U3009 (N_3009,In_40,In_1759);
and U3010 (N_3010,In_1934,In_621);
and U3011 (N_3011,In_2096,In_1005);
or U3012 (N_3012,In_1432,In_1992);
nor U3013 (N_3013,In_398,In_1486);
xor U3014 (N_3014,In_945,In_2029);
nand U3015 (N_3015,In_553,In_886);
nand U3016 (N_3016,In_88,In_1372);
nor U3017 (N_3017,In_2424,In_1982);
xor U3018 (N_3018,In_241,In_2475);
or U3019 (N_3019,In_386,In_1544);
nand U3020 (N_3020,In_965,In_212);
nand U3021 (N_3021,In_612,In_92);
or U3022 (N_3022,In_1718,In_2130);
nor U3023 (N_3023,In_2046,In_1401);
and U3024 (N_3024,In_187,In_1549);
nor U3025 (N_3025,In_1509,In_1571);
nor U3026 (N_3026,In_1007,In_1193);
nand U3027 (N_3027,In_1197,In_802);
or U3028 (N_3028,In_1653,In_33);
nor U3029 (N_3029,In_1565,In_334);
nor U3030 (N_3030,In_2456,In_683);
nor U3031 (N_3031,In_807,In_733);
or U3032 (N_3032,In_1434,In_1566);
nand U3033 (N_3033,In_1591,In_2394);
nand U3034 (N_3034,In_148,In_618);
and U3035 (N_3035,In_363,In_2281);
or U3036 (N_3036,In_643,In_2318);
or U3037 (N_3037,In_522,In_596);
xor U3038 (N_3038,In_2359,In_2313);
nand U3039 (N_3039,In_1230,In_247);
and U3040 (N_3040,In_415,In_524);
or U3041 (N_3041,In_542,In_1595);
or U3042 (N_3042,In_1269,In_1451);
or U3043 (N_3043,In_120,In_2317);
and U3044 (N_3044,In_1171,In_1890);
nand U3045 (N_3045,In_1460,In_991);
nand U3046 (N_3046,In_775,In_695);
and U3047 (N_3047,In_2211,In_1857);
or U3048 (N_3048,In_88,In_1624);
and U3049 (N_3049,In_784,In_1016);
nand U3050 (N_3050,In_2412,In_1961);
nor U3051 (N_3051,In_2372,In_1220);
or U3052 (N_3052,In_1309,In_1537);
or U3053 (N_3053,In_1238,In_2277);
and U3054 (N_3054,In_2071,In_71);
nor U3055 (N_3055,In_1795,In_1769);
nor U3056 (N_3056,In_1996,In_651);
or U3057 (N_3057,In_951,In_623);
nor U3058 (N_3058,In_415,In_2240);
or U3059 (N_3059,In_2095,In_1550);
nor U3060 (N_3060,In_1329,In_2008);
or U3061 (N_3061,In_1409,In_996);
and U3062 (N_3062,In_775,In_556);
nor U3063 (N_3063,In_206,In_923);
or U3064 (N_3064,In_715,In_1534);
nor U3065 (N_3065,In_835,In_668);
nor U3066 (N_3066,In_882,In_1976);
nor U3067 (N_3067,In_1924,In_1316);
and U3068 (N_3068,In_1967,In_1045);
nand U3069 (N_3069,In_223,In_1348);
or U3070 (N_3070,In_1366,In_1380);
or U3071 (N_3071,In_1331,In_2371);
and U3072 (N_3072,In_251,In_1722);
xor U3073 (N_3073,In_2075,In_334);
and U3074 (N_3074,In_852,In_300);
xnor U3075 (N_3075,In_2235,In_1940);
and U3076 (N_3076,In_2381,In_1127);
or U3077 (N_3077,In_1481,In_1979);
nand U3078 (N_3078,In_2423,In_1271);
or U3079 (N_3079,In_1640,In_244);
nand U3080 (N_3080,In_1268,In_348);
nor U3081 (N_3081,In_2431,In_2047);
nor U3082 (N_3082,In_1689,In_1621);
or U3083 (N_3083,In_872,In_971);
nand U3084 (N_3084,In_803,In_742);
nand U3085 (N_3085,In_2313,In_1638);
and U3086 (N_3086,In_1490,In_1169);
xor U3087 (N_3087,In_17,In_401);
nor U3088 (N_3088,In_1700,In_1424);
or U3089 (N_3089,In_228,In_140);
nand U3090 (N_3090,In_1788,In_2159);
and U3091 (N_3091,In_114,In_2407);
or U3092 (N_3092,In_2249,In_2299);
and U3093 (N_3093,In_1965,In_1909);
nor U3094 (N_3094,In_286,In_478);
or U3095 (N_3095,In_266,In_1610);
nand U3096 (N_3096,In_373,In_1571);
nand U3097 (N_3097,In_624,In_1846);
or U3098 (N_3098,In_1315,In_2338);
or U3099 (N_3099,In_453,In_1220);
and U3100 (N_3100,In_31,In_629);
nand U3101 (N_3101,In_19,In_1563);
nor U3102 (N_3102,In_2046,In_1051);
and U3103 (N_3103,In_1098,In_1793);
and U3104 (N_3104,In_809,In_332);
or U3105 (N_3105,In_2077,In_1333);
xnor U3106 (N_3106,In_1046,In_1297);
nor U3107 (N_3107,In_564,In_2275);
or U3108 (N_3108,In_1296,In_87);
and U3109 (N_3109,In_1904,In_947);
xnor U3110 (N_3110,In_465,In_1448);
and U3111 (N_3111,In_107,In_17);
nor U3112 (N_3112,In_275,In_1456);
or U3113 (N_3113,In_1424,In_992);
and U3114 (N_3114,In_96,In_2255);
xnor U3115 (N_3115,In_2417,In_902);
and U3116 (N_3116,In_1406,In_483);
nand U3117 (N_3117,In_1900,In_1659);
or U3118 (N_3118,In_1541,In_903);
nand U3119 (N_3119,In_1837,In_1971);
nand U3120 (N_3120,In_920,In_552);
or U3121 (N_3121,In_137,In_1706);
nand U3122 (N_3122,In_1679,In_1199);
xnor U3123 (N_3123,In_2256,In_744);
nand U3124 (N_3124,In_1275,In_228);
and U3125 (N_3125,N_788,N_1746);
and U3126 (N_3126,N_31,N_2280);
nand U3127 (N_3127,N_2148,N_2165);
xor U3128 (N_3128,N_2955,N_1594);
xnor U3129 (N_3129,N_1936,N_2839);
or U3130 (N_3130,N_1090,N_0);
nand U3131 (N_3131,N_2994,N_125);
nor U3132 (N_3132,N_275,N_1792);
or U3133 (N_3133,N_1557,N_1303);
or U3134 (N_3134,N_2670,N_2264);
nand U3135 (N_3135,N_1293,N_2471);
nand U3136 (N_3136,N_1730,N_422);
and U3137 (N_3137,N_833,N_2926);
or U3138 (N_3138,N_2145,N_1353);
xor U3139 (N_3139,N_898,N_826);
nand U3140 (N_3140,N_507,N_289);
xnor U3141 (N_3141,N_1677,N_554);
and U3142 (N_3142,N_984,N_27);
nor U3143 (N_3143,N_115,N_2474);
or U3144 (N_3144,N_1050,N_2430);
and U3145 (N_3145,N_2940,N_2971);
nand U3146 (N_3146,N_659,N_2056);
and U3147 (N_3147,N_1211,N_685);
or U3148 (N_3148,N_2563,N_1933);
nand U3149 (N_3149,N_1672,N_2228);
or U3150 (N_3150,N_609,N_356);
or U3151 (N_3151,N_2000,N_1925);
nand U3152 (N_3152,N_1100,N_2151);
nand U3153 (N_3153,N_2390,N_2395);
or U3154 (N_3154,N_1463,N_2028);
and U3155 (N_3155,N_2797,N_1983);
nor U3156 (N_3156,N_2951,N_1567);
nand U3157 (N_3157,N_305,N_658);
nand U3158 (N_3158,N_1629,N_2365);
nand U3159 (N_3159,N_1054,N_2686);
nor U3160 (N_3160,N_46,N_2210);
and U3161 (N_3161,N_1878,N_1262);
nand U3162 (N_3162,N_1882,N_2531);
and U3163 (N_3163,N_2335,N_583);
and U3164 (N_3164,N_1074,N_974);
xnor U3165 (N_3165,N_2302,N_1501);
nand U3166 (N_3166,N_936,N_1214);
and U3167 (N_3167,N_357,N_2241);
nor U3168 (N_3168,N_727,N_2178);
xnor U3169 (N_3169,N_1381,N_1717);
nor U3170 (N_3170,N_1448,N_116);
nand U3171 (N_3171,N_436,N_1450);
or U3172 (N_3172,N_1078,N_2041);
nand U3173 (N_3173,N_1409,N_2019);
nand U3174 (N_3174,N_418,N_1583);
and U3175 (N_3175,N_1135,N_267);
xnor U3176 (N_3176,N_2642,N_816);
nand U3177 (N_3177,N_1774,N_2158);
nand U3178 (N_3178,N_339,N_1888);
nand U3179 (N_3179,N_1053,N_2063);
nand U3180 (N_3180,N_2776,N_2924);
nor U3181 (N_3181,N_1979,N_142);
or U3182 (N_3182,N_3101,N_183);
and U3183 (N_3183,N_99,N_1119);
xor U3184 (N_3184,N_1616,N_2164);
nand U3185 (N_3185,N_128,N_725);
nor U3186 (N_3186,N_465,N_2293);
nand U3187 (N_3187,N_251,N_1109);
or U3188 (N_3188,N_603,N_2976);
and U3189 (N_3189,N_838,N_1222);
nand U3190 (N_3190,N_2123,N_1977);
nand U3191 (N_3191,N_1121,N_1230);
nor U3192 (N_3192,N_2345,N_3002);
nand U3193 (N_3193,N_2634,N_208);
nor U3194 (N_3194,N_943,N_1292);
nand U3195 (N_3195,N_225,N_3042);
nand U3196 (N_3196,N_2486,N_3009);
or U3197 (N_3197,N_491,N_1867);
nand U3198 (N_3198,N_1043,N_2785);
or U3199 (N_3199,N_1428,N_2403);
nor U3200 (N_3200,N_317,N_1896);
nand U3201 (N_3201,N_3046,N_229);
nor U3202 (N_3202,N_2074,N_1005);
and U3203 (N_3203,N_1974,N_2009);
nand U3204 (N_3204,N_2016,N_878);
and U3205 (N_3205,N_162,N_469);
nand U3206 (N_3206,N_2918,N_1963);
nand U3207 (N_3207,N_735,N_1953);
nand U3208 (N_3208,N_1511,N_672);
nor U3209 (N_3209,N_1732,N_1505);
nor U3210 (N_3210,N_1604,N_1270);
nand U3211 (N_3211,N_2549,N_828);
and U3212 (N_3212,N_230,N_2472);
nor U3213 (N_3213,N_3112,N_2844);
and U3214 (N_3214,N_2411,N_560);
xor U3215 (N_3215,N_1092,N_2595);
nand U3216 (N_3216,N_261,N_1171);
nor U3217 (N_3217,N_1662,N_856);
nand U3218 (N_3218,N_997,N_2792);
nor U3219 (N_3219,N_1601,N_693);
and U3220 (N_3220,N_1724,N_2653);
xnor U3221 (N_3221,N_873,N_463);
nand U3222 (N_3222,N_568,N_2666);
nand U3223 (N_3223,N_596,N_1151);
or U3224 (N_3224,N_3033,N_2214);
or U3225 (N_3225,N_2993,N_790);
and U3226 (N_3226,N_2155,N_3060);
nor U3227 (N_3227,N_2311,N_384);
nor U3228 (N_3228,N_2484,N_1081);
and U3229 (N_3229,N_493,N_2870);
xnor U3230 (N_3230,N_487,N_1734);
nand U3231 (N_3231,N_2194,N_3084);
nor U3232 (N_3232,N_1679,N_412);
nand U3233 (N_3233,N_1834,N_1909);
or U3234 (N_3234,N_1014,N_2259);
nand U3235 (N_3235,N_3068,N_1346);
and U3236 (N_3236,N_1651,N_846);
or U3237 (N_3237,N_2017,N_626);
xor U3238 (N_3238,N_450,N_1153);
or U3239 (N_3239,N_1449,N_1653);
and U3240 (N_3240,N_2719,N_777);
xnor U3241 (N_3241,N_695,N_1465);
and U3242 (N_3242,N_1299,N_1503);
nor U3243 (N_3243,N_2314,N_2227);
nor U3244 (N_3244,N_2256,N_2287);
xor U3245 (N_3245,N_2824,N_530);
nand U3246 (N_3246,N_879,N_241);
nor U3247 (N_3247,N_1605,N_2677);
nand U3248 (N_3248,N_3080,N_2469);
xnor U3249 (N_3249,N_243,N_1026);
and U3250 (N_3250,N_660,N_591);
and U3251 (N_3251,N_2764,N_158);
or U3252 (N_3252,N_831,N_616);
nand U3253 (N_3253,N_783,N_2551);
nand U3254 (N_3254,N_716,N_209);
or U3255 (N_3255,N_2803,N_3119);
and U3256 (N_3256,N_175,N_1545);
and U3257 (N_3257,N_57,N_1281);
nand U3258 (N_3258,N_2275,N_2527);
nand U3259 (N_3259,N_499,N_1420);
nand U3260 (N_3260,N_96,N_1782);
or U3261 (N_3261,N_2750,N_1149);
or U3262 (N_3262,N_2147,N_1415);
xor U3263 (N_3263,N_1033,N_2351);
nor U3264 (N_3264,N_1472,N_2692);
and U3265 (N_3265,N_2959,N_618);
and U3266 (N_3266,N_2729,N_2929);
nand U3267 (N_3267,N_1015,N_2811);
and U3268 (N_3268,N_2691,N_1948);
nor U3269 (N_3269,N_2808,N_1273);
nand U3270 (N_3270,N_68,N_2582);
xor U3271 (N_3271,N_2783,N_1370);
nor U3272 (N_3272,N_859,N_1426);
and U3273 (N_3273,N_1533,N_2629);
xor U3274 (N_3274,N_3007,N_822);
nand U3275 (N_3275,N_2861,N_2829);
nor U3276 (N_3276,N_2204,N_1890);
and U3277 (N_3277,N_1970,N_324);
xnor U3278 (N_3278,N_227,N_1831);
and U3279 (N_3279,N_649,N_2613);
and U3280 (N_3280,N_2752,N_2172);
xnor U3281 (N_3281,N_667,N_1253);
nor U3282 (N_3282,N_2543,N_2628);
nor U3283 (N_3283,N_1279,N_945);
and U3284 (N_3284,N_19,N_653);
nand U3285 (N_3285,N_501,N_2047);
or U3286 (N_3286,N_1167,N_2186);
nor U3287 (N_3287,N_2967,N_191);
or U3288 (N_3288,N_1659,N_1676);
and U3289 (N_3289,N_2508,N_2916);
and U3290 (N_3290,N_2413,N_2745);
nor U3291 (N_3291,N_1927,N_1161);
nand U3292 (N_3292,N_1124,N_127);
or U3293 (N_3293,N_726,N_2076);
or U3294 (N_3294,N_222,N_2420);
and U3295 (N_3295,N_1328,N_1061);
or U3296 (N_3296,N_2415,N_3093);
xor U3297 (N_3297,N_2012,N_160);
nand U3298 (N_3298,N_2272,N_1249);
nand U3299 (N_3299,N_836,N_448);
or U3300 (N_3300,N_1769,N_470);
or U3301 (N_3301,N_2910,N_2466);
and U3302 (N_3302,N_1203,N_2325);
and U3303 (N_3303,N_781,N_1291);
and U3304 (N_3304,N_2029,N_2944);
nor U3305 (N_3305,N_181,N_1787);
or U3306 (N_3306,N_1194,N_1064);
xnor U3307 (N_3307,N_1147,N_425);
nor U3308 (N_3308,N_2922,N_2648);
or U3309 (N_3309,N_1714,N_2310);
nand U3310 (N_3310,N_925,N_546);
nor U3311 (N_3311,N_2289,N_1775);
xnor U3312 (N_3312,N_3074,N_1471);
or U3313 (N_3313,N_3024,N_2689);
xor U3314 (N_3314,N_1245,N_2079);
or U3315 (N_3315,N_544,N_1178);
nor U3316 (N_3316,N_865,N_1911);
nor U3317 (N_3317,N_2840,N_2826);
and U3318 (N_3318,N_3057,N_671);
nor U3319 (N_3319,N_2675,N_2759);
nor U3320 (N_3320,N_304,N_3012);
or U3321 (N_3321,N_2298,N_1688);
xnor U3322 (N_3322,N_2377,N_1785);
or U3323 (N_3323,N_2442,N_114);
nand U3324 (N_3324,N_565,N_611);
and U3325 (N_3325,N_1767,N_402);
and U3326 (N_3326,N_576,N_488);
nor U3327 (N_3327,N_1550,N_1524);
and U3328 (N_3328,N_1352,N_2733);
nor U3329 (N_3329,N_1058,N_2331);
nor U3330 (N_3330,N_1267,N_2159);
nor U3331 (N_3331,N_1210,N_1294);
and U3332 (N_3332,N_1703,N_919);
nand U3333 (N_3333,N_526,N_33);
nand U3334 (N_3334,N_2682,N_745);
or U3335 (N_3335,N_1591,N_636);
nand U3336 (N_3336,N_1197,N_1514);
nand U3337 (N_3337,N_2893,N_1117);
nor U3338 (N_3338,N_1917,N_399);
nand U3339 (N_3339,N_1941,N_219);
nand U3340 (N_3340,N_2412,N_1059);
nand U3341 (N_3341,N_2681,N_170);
or U3342 (N_3342,N_109,N_1846);
and U3343 (N_3343,N_1452,N_458);
and U3344 (N_3344,N_2268,N_542);
nor U3345 (N_3345,N_2226,N_1455);
or U3346 (N_3346,N_255,N_1172);
or U3347 (N_3347,N_1981,N_2905);
and U3348 (N_3348,N_3066,N_1742);
and U3349 (N_3349,N_521,N_2815);
and U3350 (N_3350,N_3117,N_1099);
and U3351 (N_3351,N_1154,N_1393);
nand U3352 (N_3352,N_2878,N_2044);
or U3353 (N_3353,N_1741,N_3000);
nand U3354 (N_3354,N_2175,N_703);
nor U3355 (N_3355,N_1069,N_361);
or U3356 (N_3356,N_1424,N_2282);
and U3357 (N_3357,N_1362,N_2344);
or U3358 (N_3358,N_2478,N_553);
and U3359 (N_3359,N_510,N_1971);
nand U3360 (N_3360,N_1924,N_1108);
or U3361 (N_3361,N_2769,N_90);
or U3362 (N_3362,N_1592,N_2424);
or U3363 (N_3363,N_627,N_299);
nand U3364 (N_3364,N_1079,N_2939);
and U3365 (N_3365,N_45,N_2771);
nor U3366 (N_3366,N_931,N_2376);
and U3367 (N_3367,N_2132,N_2872);
and U3368 (N_3368,N_1887,N_1634);
or U3369 (N_3369,N_1858,N_2470);
and U3370 (N_3370,N_2234,N_2972);
nand U3371 (N_3371,N_166,N_1182);
or U3372 (N_3372,N_2532,N_1699);
and U3373 (N_3373,N_126,N_1803);
nand U3374 (N_3374,N_247,N_767);
and U3375 (N_3375,N_203,N_400);
nor U3376 (N_3376,N_145,N_497);
and U3377 (N_3377,N_338,N_2945);
nor U3378 (N_3378,N_2251,N_2312);
nand U3379 (N_3379,N_582,N_65);
or U3380 (N_3380,N_2617,N_902);
and U3381 (N_3381,N_364,N_1901);
nor U3382 (N_3382,N_891,N_1287);
and U3383 (N_3383,N_2419,N_4);
xor U3384 (N_3384,N_2193,N_3086);
and U3385 (N_3385,N_1793,N_1563);
nor U3386 (N_3386,N_1619,N_2254);
or U3387 (N_3387,N_2748,N_2949);
nand U3388 (N_3388,N_1635,N_1935);
nand U3389 (N_3389,N_2743,N_993);
and U3390 (N_3390,N_721,N_625);
or U3391 (N_3391,N_140,N_1146);
or U3392 (N_3392,N_2477,N_2989);
and U3393 (N_3393,N_2676,N_1670);
or U3394 (N_3394,N_2581,N_2011);
nor U3395 (N_3395,N_2913,N_2589);
nor U3396 (N_3396,N_11,N_1928);
nand U3397 (N_3397,N_2524,N_1906);
xnor U3398 (N_3398,N_1736,N_1814);
and U3399 (N_3399,N_2946,N_2979);
and U3400 (N_3400,N_646,N_88);
and U3401 (N_3401,N_2075,N_337);
or U3402 (N_3402,N_2775,N_3105);
and U3403 (N_3403,N_2115,N_3035);
xnor U3404 (N_3404,N_2552,N_870);
nand U3405 (N_3405,N_713,N_82);
and U3406 (N_3406,N_682,N_2257);
or U3407 (N_3407,N_743,N_1068);
or U3408 (N_3408,N_1019,N_608);
and U3409 (N_3409,N_832,N_1470);
nor U3410 (N_3410,N_478,N_848);
nand U3411 (N_3411,N_1722,N_2665);
nand U3412 (N_3412,N_100,N_498);
nand U3413 (N_3413,N_2970,N_2805);
or U3414 (N_3414,N_1645,N_1978);
and U3415 (N_3415,N_2146,N_1160);
nor U3416 (N_3416,N_540,N_2458);
nand U3417 (N_3417,N_843,N_1950);
or U3418 (N_3418,N_1145,N_2343);
nand U3419 (N_3419,N_1038,N_1300);
nand U3420 (N_3420,N_306,N_1157);
and U3421 (N_3421,N_1159,N_2822);
nor U3422 (N_3422,N_2947,N_683);
or U3423 (N_3423,N_2643,N_1200);
nor U3424 (N_3424,N_1016,N_2170);
xnor U3425 (N_3425,N_1175,N_1812);
or U3426 (N_3426,N_426,N_2909);
or U3427 (N_3427,N_1044,N_246);
or U3428 (N_3428,N_1401,N_957);
and U3429 (N_3429,N_3071,N_60);
nand U3430 (N_3430,N_679,N_1341);
nand U3431 (N_3431,N_877,N_1045);
and U3432 (N_3432,N_1949,N_2207);
xor U3433 (N_3433,N_1333,N_2723);
and U3434 (N_3434,N_2435,N_1283);
nand U3435 (N_3435,N_2454,N_277);
nor U3436 (N_3436,N_912,N_1542);
xor U3437 (N_3437,N_1539,N_808);
nor U3438 (N_3438,N_852,N_2473);
nor U3439 (N_3439,N_1566,N_1892);
nor U3440 (N_3440,N_2751,N_168);
and U3441 (N_3441,N_737,N_2206);
or U3442 (N_3442,N_1274,N_2190);
nand U3443 (N_3443,N_533,N_2284);
nand U3444 (N_3444,N_427,N_2927);
nor U3445 (N_3445,N_2183,N_2977);
nand U3446 (N_3446,N_1847,N_1894);
or U3447 (N_3447,N_941,N_1838);
and U3448 (N_3448,N_1719,N_2656);
nand U3449 (N_3449,N_2818,N_575);
nor U3450 (N_3450,N_350,N_2867);
nand U3451 (N_3451,N_634,N_1359);
and U3452 (N_3452,N_1460,N_2574);
or U3453 (N_3453,N_824,N_1883);
nor U3454 (N_3454,N_2295,N_702);
and U3455 (N_3455,N_397,N_1349);
nand U3456 (N_3456,N_1740,N_1013);
nor U3457 (N_3457,N_85,N_428);
nor U3458 (N_3458,N_599,N_2778);
xnor U3459 (N_3459,N_2220,N_2460);
and U3460 (N_3460,N_2702,N_1739);
and U3461 (N_3461,N_217,N_1073);
nor U3462 (N_3462,N_1868,N_2630);
nor U3463 (N_3463,N_1399,N_2966);
and U3464 (N_3464,N_269,N_319);
and U3465 (N_3465,N_2627,N_2375);
or U3466 (N_3466,N_1041,N_897);
xnor U3467 (N_3467,N_2746,N_2489);
or U3468 (N_3468,N_1084,N_1482);
nor U3469 (N_3469,N_1585,N_2570);
nand U3470 (N_3470,N_1276,N_651);
nand U3471 (N_3471,N_437,N_975);
nand U3472 (N_3472,N_1029,N_2704);
nand U3473 (N_3473,N_3124,N_91);
nand U3474 (N_3474,N_2038,N_2902);
or U3475 (N_3475,N_2931,N_815);
nand U3476 (N_3476,N_1599,N_2058);
nor U3477 (N_3477,N_2493,N_1086);
nor U3478 (N_3478,N_2736,N_678);
nor U3479 (N_3479,N_503,N_1205);
or U3480 (N_3480,N_869,N_691);
nand U3481 (N_3481,N_791,N_1902);
nand U3482 (N_3482,N_1648,N_2523);
or U3483 (N_3483,N_360,N_2936);
or U3484 (N_3484,N_334,N_189);
and U3485 (N_3485,N_1817,N_2128);
nor U3486 (N_3486,N_1560,N_2305);
or U3487 (N_3487,N_1819,N_2757);
or U3488 (N_3488,N_373,N_2984);
nand U3489 (N_3489,N_871,N_2481);
nor U3490 (N_3490,N_143,N_2758);
and U3491 (N_3491,N_2669,N_1515);
or U3492 (N_3492,N_333,N_2232);
xnor U3493 (N_3493,N_2001,N_742);
nor U3494 (N_3494,N_2651,N_1444);
nand U3495 (N_3495,N_1179,N_1326);
nor U3496 (N_3496,N_761,N_2113);
nor U3497 (N_3497,N_2592,N_2594);
nor U3498 (N_3498,N_2361,N_766);
xnor U3499 (N_3499,N_2754,N_250);
nand U3500 (N_3500,N_1640,N_951);
nand U3501 (N_3501,N_1395,N_2942);
nand U3502 (N_3502,N_2566,N_1708);
nand U3503 (N_3503,N_2536,N_2933);
and U3504 (N_3504,N_163,N_3038);
nor U3505 (N_3505,N_592,N_950);
nand U3506 (N_3506,N_2299,N_963);
and U3507 (N_3507,N_366,N_2036);
nand U3508 (N_3508,N_252,N_2786);
and U3509 (N_3509,N_259,N_3067);
nand U3510 (N_3510,N_1541,N_988);
nor U3511 (N_3511,N_1419,N_2427);
nand U3512 (N_3512,N_2447,N_1036);
nor U3513 (N_3513,N_628,N_3118);
nand U3514 (N_3514,N_1307,N_271);
xnor U3515 (N_3515,N_2187,N_2568);
or U3516 (N_3516,N_1710,N_2231);
nor U3517 (N_3517,N_1011,N_1852);
nor U3518 (N_3518,N_1572,N_2340);
or U3519 (N_3519,N_1034,N_3055);
nor U3520 (N_3520,N_2717,N_2548);
or U3521 (N_3521,N_340,N_1956);
and U3522 (N_3522,N_2690,N_729);
nor U3523 (N_3523,N_1697,N_570);
or U3524 (N_3524,N_823,N_442);
or U3525 (N_3525,N_1323,N_3085);
and U3526 (N_3526,N_1675,N_249);
xnor U3527 (N_3527,N_1586,N_2810);
or U3528 (N_3528,N_39,N_1298);
nand U3529 (N_3529,N_1748,N_2384);
xnor U3530 (N_3530,N_1116,N_2124);
and U3531 (N_3531,N_2911,N_1822);
nor U3532 (N_3532,N_1989,N_2858);
and U3533 (N_3533,N_2890,N_1666);
and U3534 (N_3534,N_1798,N_1305);
nor U3535 (N_3535,N_3082,N_1313);
and U3536 (N_3536,N_1646,N_971);
nor U3537 (N_3537,N_1423,N_1707);
or U3538 (N_3538,N_1582,N_961);
or U3539 (N_3539,N_665,N_2740);
xor U3540 (N_3540,N_1735,N_2097);
xnor U3541 (N_3541,N_287,N_17);
or U3542 (N_3542,N_2386,N_2042);
and U3543 (N_3543,N_803,N_110);
or U3544 (N_3544,N_2812,N_489);
nor U3545 (N_3545,N_2958,N_1327);
nor U3546 (N_3546,N_2995,N_3083);
xnor U3547 (N_3547,N_2294,N_612);
xor U3548 (N_3548,N_1952,N_2080);
and U3549 (N_3549,N_1148,N_1723);
or U3550 (N_3550,N_1136,N_1255);
and U3551 (N_3551,N_2276,N_1510);
and U3552 (N_3552,N_1277,N_1637);
nand U3553 (N_3553,N_3072,N_2306);
or U3554 (N_3554,N_2117,N_3039);
xor U3555 (N_3555,N_192,N_899);
nand U3556 (N_3556,N_419,N_2426);
xnor U3557 (N_3557,N_1198,N_1229);
nand U3558 (N_3558,N_347,N_780);
nor U3559 (N_3559,N_1414,N_2002);
nor U3560 (N_3560,N_1031,N_2610);
and U3561 (N_3561,N_380,N_2333);
nor U3562 (N_3562,N_365,N_2197);
or U3563 (N_3563,N_1919,N_2108);
nand U3564 (N_3564,N_1508,N_2842);
or U3565 (N_3565,N_2860,N_802);
or U3566 (N_3566,N_779,N_632);
nand U3567 (N_3567,N_1168,N_441);
nor U3568 (N_3568,N_129,N_1296);
or U3569 (N_3569,N_2322,N_1573);
and U3570 (N_3570,N_631,N_1521);
or U3571 (N_3571,N_1966,N_2171);
nor U3572 (N_3572,N_439,N_1371);
and U3573 (N_3573,N_918,N_2485);
nand U3574 (N_3574,N_2587,N_104);
and U3575 (N_3575,N_1664,N_711);
nand U3576 (N_3576,N_475,N_1481);
or U3577 (N_3577,N_650,N_2596);
nand U3578 (N_3578,N_937,N_1318);
and U3579 (N_3579,N_2347,N_904);
nand U3580 (N_3580,N_2919,N_174);
or U3581 (N_3581,N_1209,N_1627);
nor U3582 (N_3582,N_457,N_2832);
nor U3583 (N_3583,N_494,N_296);
nor U3584 (N_3584,N_597,N_744);
nor U3585 (N_3585,N_1569,N_2537);
nand U3586 (N_3586,N_1489,N_699);
nor U3587 (N_3587,N_106,N_923);
xnor U3588 (N_3588,N_2843,N_1944);
or U3589 (N_3589,N_2092,N_2957);
xor U3590 (N_3590,N_1795,N_1526);
or U3591 (N_3591,N_118,N_452);
or U3592 (N_3592,N_960,N_1347);
or U3593 (N_3593,N_2006,N_362);
or U3594 (N_3594,N_1926,N_2585);
nor U3595 (N_3595,N_483,N_895);
nor U3596 (N_3596,N_2650,N_484);
nand U3597 (N_3597,N_2897,N_1791);
and U3598 (N_3598,N_1777,N_1558);
nor U3599 (N_3599,N_1330,N_6);
and U3600 (N_3600,N_358,N_2327);
or U3601 (N_3601,N_2281,N_811);
xor U3602 (N_3602,N_50,N_2678);
and U3603 (N_3603,N_325,N_1856);
nor U3604 (N_3604,N_1727,N_537);
nand U3605 (N_3605,N_1478,N_2088);
or U3606 (N_3606,N_1725,N_161);
or U3607 (N_3607,N_2359,N_2865);
or U3608 (N_3608,N_654,N_2433);
nand U3609 (N_3609,N_2766,N_1325);
nor U3610 (N_3610,N_1243,N_1130);
or U3611 (N_3611,N_607,N_1163);
nand U3612 (N_3612,N_2189,N_1506);
or U3613 (N_3613,N_41,N_928);
xor U3614 (N_3614,N_1995,N_2889);
and U3615 (N_3615,N_2948,N_1874);
and U3616 (N_3616,N_1403,N_1378);
nand U3617 (N_3617,N_2176,N_297);
and U3618 (N_3618,N_817,N_176);
and U3619 (N_3619,N_758,N_1991);
nand U3620 (N_3620,N_837,N_1096);
and U3621 (N_3621,N_69,N_177);
or U3622 (N_3622,N_1260,N_1170);
nor U3623 (N_3623,N_313,N_1354);
or U3624 (N_3624,N_1006,N_980);
or U3625 (N_3625,N_541,N_1516);
nand U3626 (N_3626,N_1564,N_2631);
nand U3627 (N_3627,N_1618,N_1898);
nand U3628 (N_3628,N_2987,N_288);
nor U3629 (N_3629,N_1755,N_1879);
nand U3630 (N_3630,N_2937,N_1982);
and U3631 (N_3631,N_866,N_2875);
nor U3632 (N_3632,N_966,N_283);
and U3633 (N_3633,N_2160,N_2087);
or U3634 (N_3634,N_1959,N_2608);
nand U3635 (N_3635,N_2065,N_2816);
nor U3636 (N_3636,N_119,N_1242);
or U3637 (N_3637,N_3054,N_2782);
nand U3638 (N_3638,N_2448,N_572);
and U3639 (N_3639,N_2985,N_1110);
xor U3640 (N_3640,N_992,N_958);
nand U3641 (N_3641,N_1338,N_468);
and U3642 (N_3642,N_420,N_2601);
nand U3643 (N_3643,N_1224,N_2795);
nand U3644 (N_3644,N_689,N_1351);
nand U3645 (N_3645,N_1113,N_1310);
or U3646 (N_3646,N_3047,N_2161);
nand U3647 (N_3647,N_14,N_1150);
nor U3648 (N_3648,N_1630,N_2698);
xor U3649 (N_3649,N_1467,N_1308);
and U3650 (N_3650,N_1189,N_1588);
nor U3651 (N_3651,N_71,N_2247);
nand U3652 (N_3652,N_2607,N_1837);
or U3653 (N_3653,N_2658,N_1195);
nand U3654 (N_3654,N_1208,N_316);
nand U3655 (N_3655,N_509,N_1228);
nand U3656 (N_3656,N_552,N_1875);
nand U3657 (N_3657,N_390,N_147);
or U3658 (N_3658,N_1825,N_896);
xnor U3659 (N_3659,N_872,N_1366);
nand U3660 (N_3660,N_30,N_605);
nor U3661 (N_3661,N_2456,N_2188);
xor U3662 (N_3662,N_3077,N_240);
nand U3663 (N_3663,N_2506,N_1844);
nor U3664 (N_3664,N_2564,N_2032);
nor U3665 (N_3665,N_3058,N_2881);
nor U3666 (N_3666,N_946,N_1993);
nor U3667 (N_3667,N_675,N_137);
nor U3668 (N_3668,N_2457,N_444);
or U3669 (N_3669,N_2242,N_2779);
and U3670 (N_3670,N_2827,N_1386);
or U3671 (N_3671,N_2049,N_1413);
and U3672 (N_3672,N_1022,N_1114);
nand U3673 (N_3673,N_2154,N_2106);
xor U3674 (N_3674,N_640,N_471);
or U3675 (N_3675,N_124,N_2418);
xnor U3676 (N_3676,N_467,N_1387);
nor U3677 (N_3677,N_738,N_2250);
and U3678 (N_3678,N_1832,N_320);
or U3679 (N_3679,N_1553,N_388);
nor U3680 (N_3680,N_581,N_1028);
nand U3681 (N_3681,N_2646,N_409);
nor U3682 (N_3682,N_778,N_2514);
nand U3683 (N_3683,N_2923,N_1373);
and U3684 (N_3684,N_1805,N_2975);
and U3685 (N_3685,N_1221,N_345);
and U3686 (N_3686,N_310,N_807);
and U3687 (N_3687,N_2475,N_97);
nand U3688 (N_3688,N_890,N_1020);
xor U3689 (N_3689,N_1060,N_970);
or U3690 (N_3690,N_37,N_2372);
or U3691 (N_3691,N_917,N_3051);
nor U3692 (N_3692,N_211,N_1931);
and U3693 (N_3693,N_3026,N_224);
nor U3694 (N_3694,N_1237,N_242);
nand U3695 (N_3695,N_1869,N_1713);
nor U3696 (N_3696,N_461,N_2078);
and U3697 (N_3697,N_2848,N_1065);
or U3698 (N_3698,N_1633,N_2104);
nand U3699 (N_3699,N_1561,N_2405);
or U3700 (N_3700,N_3019,N_1383);
nand U3701 (N_3701,N_2142,N_500);
xor U3702 (N_3702,N_3106,N_1416);
or U3703 (N_3703,N_2730,N_2960);
or U3704 (N_3704,N_2899,N_314);
and U3705 (N_3705,N_1483,N_538);
xor U3706 (N_3706,N_585,N_804);
nor U3707 (N_3707,N_1565,N_1271);
nor U3708 (N_3708,N_2496,N_1280);
and U3709 (N_3709,N_1269,N_1976);
or U3710 (N_3710,N_800,N_854);
and U3711 (N_3711,N_905,N_2892);
or U3712 (N_3712,N_580,N_232);
or U3713 (N_3713,N_1631,N_22);
nand U3714 (N_3714,N_886,N_1304);
or U3715 (N_3715,N_2233,N_1910);
and U3716 (N_3716,N_740,N_929);
and U3717 (N_3717,N_2144,N_121);
nand U3718 (N_3718,N_1744,N_1192);
and U3719 (N_3719,N_1891,N_201);
or U3720 (N_3720,N_1886,N_1042);
xor U3721 (N_3721,N_237,N_2640);
nand U3722 (N_3722,N_1263,N_474);
xor U3723 (N_3723,N_281,N_3064);
nand U3724 (N_3724,N_1355,N_2432);
nand U3725 (N_3725,N_2917,N_141);
and U3726 (N_3726,N_2674,N_2394);
xor U3727 (N_3727,N_1796,N_1201);
or U3728 (N_3728,N_534,N_1864);
or U3729 (N_3729,N_138,N_1456);
nand U3730 (N_3730,N_1219,N_1760);
nand U3731 (N_3731,N_1914,N_2201);
nand U3732 (N_3732,N_3069,N_2554);
or U3733 (N_3733,N_231,N_1518);
or U3734 (N_3734,N_2152,N_1322);
nand U3735 (N_3735,N_254,N_995);
nand U3736 (N_3736,N_2023,N_2744);
nor U3737 (N_3737,N_1829,N_2290);
xnor U3738 (N_3738,N_892,N_861);
and U3739 (N_3739,N_2540,N_2838);
and U3740 (N_3740,N_1118,N_2930);
nand U3741 (N_3741,N_2143,N_2724);
nand U3742 (N_3742,N_2334,N_1309);
nand U3743 (N_3743,N_749,N_372);
nand U3744 (N_3744,N_2304,N_396);
nor U3745 (N_3745,N_792,N_590);
nor U3746 (N_3746,N_2181,N_2163);
or U3747 (N_3747,N_2436,N_2991);
nor U3748 (N_3748,N_1504,N_2659);
or U3749 (N_3749,N_1836,N_1799);
nor U3750 (N_3750,N_619,N_690);
xor U3751 (N_3751,N_2586,N_1334);
nand U3752 (N_3752,N_2755,N_89);
nor U3753 (N_3753,N_708,N_1070);
nand U3754 (N_3754,N_733,N_2051);
nor U3755 (N_3755,N_2813,N_370);
or U3756 (N_3756,N_1965,N_855);
and U3757 (N_3757,N_2423,N_719);
nor U3758 (N_3758,N_2279,N_3062);
nand U3759 (N_3759,N_291,N_2525);
nor U3760 (N_3760,N_433,N_1407);
nor U3761 (N_3761,N_1385,N_548);
or U3762 (N_3762,N_2066,N_875);
nor U3763 (N_3763,N_2439,N_1750);
and U3764 (N_3764,N_1809,N_173);
and U3765 (N_3765,N_2992,N_629);
or U3766 (N_3766,N_1636,N_2301);
and U3767 (N_3767,N_2391,N_1442);
nand U3768 (N_3768,N_1112,N_20);
nand U3769 (N_3769,N_2480,N_736);
nor U3770 (N_3770,N_391,N_2777);
nand U3771 (N_3771,N_2535,N_985);
nor U3772 (N_3772,N_1839,N_307);
xnor U3773 (N_3773,N_1134,N_1529);
and U3774 (N_3774,N_1626,N_2003);
nor U3775 (N_3775,N_3029,N_2252);
xor U3776 (N_3776,N_21,N_344);
nand U3777 (N_3777,N_3023,N_1821);
nand U3778 (N_3778,N_2297,N_911);
nor U3779 (N_3779,N_2800,N_1227);
or U3780 (N_3780,N_186,N_234);
and U3781 (N_3781,N_857,N_2672);
xor U3782 (N_3782,N_184,N_1088);
nand U3783 (N_3783,N_1693,N_387);
and U3784 (N_3784,N_1964,N_446);
and U3785 (N_3785,N_600,N_2440);
nand U3786 (N_3786,N_1379,N_2084);
and U3787 (N_3787,N_1238,N_785);
nand U3788 (N_3788,N_561,N_2073);
and U3789 (N_3789,N_87,N_2762);
nor U3790 (N_3790,N_1613,N_180);
or U3791 (N_3791,N_323,N_2738);
and U3792 (N_3792,N_1315,N_2071);
and U3793 (N_3793,N_154,N_2632);
and U3794 (N_3794,N_2468,N_773);
nor U3795 (N_3795,N_1344,N_80);
nor U3796 (N_3796,N_2638,N_680);
nand U3797 (N_3797,N_587,N_797);
and U3798 (N_3798,N_1772,N_579);
nand U3799 (N_3799,N_260,N_1376);
and U3800 (N_3800,N_1556,N_2626);
and U3801 (N_3801,N_1311,N_1876);
or U3802 (N_3802,N_98,N_1716);
nand U3803 (N_3803,N_3008,N_2083);
nand U3804 (N_3804,N_2027,N_706);
nor U3805 (N_3805,N_2168,N_624);
or U3806 (N_3806,N_3004,N_2445);
nand U3807 (N_3807,N_2520,N_511);
or U3808 (N_3808,N_2647,N_1432);
nand U3809 (N_3809,N_2950,N_1780);
nand U3810 (N_3810,N_760,N_2982);
nand U3811 (N_3811,N_2753,N_2379);
nor U3812 (N_3812,N_1845,N_438);
or U3813 (N_3813,N_1412,N_1388);
or U3814 (N_3814,N_2664,N_2560);
xnor U3815 (N_3815,N_701,N_1174);
nor U3816 (N_3816,N_1535,N_1190);
and U3817 (N_3817,N_944,N_2662);
or U3818 (N_3818,N_2920,N_1921);
or U3819 (N_3819,N_1830,N_1234);
nand U3820 (N_3820,N_1431,N_1536);
and U3821 (N_3821,N_2696,N_1903);
and U3822 (N_3822,N_1579,N_190);
xnor U3823 (N_3823,N_1468,N_1581);
or U3824 (N_3824,N_2732,N_2487);
nand U3825 (N_3825,N_1144,N_1486);
nand U3826 (N_3826,N_1236,N_933);
nor U3827 (N_3827,N_1361,N_1040);
xnor U3828 (N_3828,N_1212,N_1623);
and U3829 (N_3829,N_329,N_105);
nand U3830 (N_3830,N_903,N_371);
nor U3831 (N_3831,N_54,N_3102);
nand U3832 (N_3832,N_2368,N_967);
nand U3833 (N_3833,N_171,N_516);
xnor U3834 (N_3834,N_1823,N_477);
nand U3835 (N_3835,N_1870,N_2884);
or U3836 (N_3836,N_1430,N_2238);
nand U3837 (N_3837,N_2374,N_1781);
nand U3838 (N_3838,N_1968,N_383);
and U3839 (N_3839,N_1226,N_1638);
and U3840 (N_3840,N_92,N_1973);
nand U3841 (N_3841,N_1106,N_1196);
and U3842 (N_3842,N_1316,N_741);
or U3843 (N_3843,N_593,N_3114);
nor U3844 (N_3844,N_482,N_2680);
nand U3845 (N_3845,N_676,N_2342);
and U3846 (N_3846,N_1816,N_3099);
or U3847 (N_3847,N_2693,N_1806);
and U3848 (N_3848,N_2321,N_1686);
nand U3849 (N_3849,N_1986,N_207);
nor U3850 (N_3850,N_601,N_464);
and U3851 (N_3851,N_753,N_858);
or U3852 (N_3852,N_152,N_3049);
nor U3853 (N_3853,N_1225,N_1000);
or U3854 (N_3854,N_2761,N_1669);
and U3855 (N_3855,N_2410,N_1815);
nor U3856 (N_3856,N_976,N_1595);
nand U3857 (N_3857,N_1895,N_1389);
and U3858 (N_3858,N_2094,N_1446);
and U3859 (N_3859,N_2015,N_549);
nand U3860 (N_3860,N_723,N_1286);
xor U3861 (N_3861,N_2500,N_2635);
and U3862 (N_3862,N_2547,N_2541);
nor U3863 (N_3863,N_2034,N_38);
nand U3864 (N_3864,N_2369,N_1375);
nand U3865 (N_3865,N_2406,N_429);
nor U3866 (N_3866,N_2973,N_2273);
nand U3867 (N_3867,N_40,N_1589);
and U3868 (N_3868,N_3018,N_2774);
and U3869 (N_3869,N_1247,N_821);
nor U3870 (N_3870,N_673,N_2018);
nor U3871 (N_3871,N_2048,N_414);
and U3872 (N_3872,N_2599,N_2184);
and U3873 (N_3873,N_914,N_775);
nand U3874 (N_3874,N_2820,N_2851);
xor U3875 (N_3875,N_1337,N_215);
nand U3876 (N_3876,N_2072,N_2713);
or U3877 (N_3877,N_952,N_2718);
nand U3878 (N_3878,N_633,N_1487);
nor U3879 (N_3879,N_66,N_2326);
nor U3880 (N_3880,N_2059,N_70);
and U3881 (N_3881,N_1984,N_1548);
or U3882 (N_3882,N_617,N_1988);
xnor U3883 (N_3883,N_1493,N_1216);
nand U3884 (N_3884,N_556,N_2804);
or U3885 (N_3885,N_2542,N_1275);
nand U3886 (N_3886,N_2590,N_55);
xor U3887 (N_3887,N_401,N_2313);
or U3888 (N_3888,N_3020,N_2482);
nand U3889 (N_3889,N_2192,N_1922);
or U3890 (N_3890,N_1920,N_172);
nor U3891 (N_3891,N_3090,N_2615);
and U3892 (N_3892,N_2641,N_704);
xor U3893 (N_3893,N_1055,N_1720);
nand U3894 (N_3894,N_2502,N_2396);
nand U3895 (N_3895,N_2383,N_1075);
and U3896 (N_3896,N_1840,N_1377);
xnor U3897 (N_3897,N_2687,N_924);
nand U3898 (N_3898,N_1418,N_2577);
nor U3899 (N_3899,N_2303,N_2025);
nand U3900 (N_3900,N_2417,N_1833);
nor U3901 (N_3901,N_3027,N_2216);
xnor U3902 (N_3902,N_1102,N_1574);
and U3903 (N_3903,N_2307,N_1811);
nand U3904 (N_3904,N_2528,N_3103);
and U3905 (N_3905,N_717,N_301);
nor U3906 (N_3906,N_3036,N_2999);
nor U3907 (N_3907,N_2954,N_2434);
and U3908 (N_3908,N_117,N_1773);
or U3909 (N_3909,N_1621,N_2246);
or U3910 (N_3910,N_732,N_3097);
or U3911 (N_3911,N_2512,N_1751);
or U3912 (N_3912,N_934,N_2900);
and U3913 (N_3913,N_1990,N_424);
and U3914 (N_3914,N_2236,N_3073);
and U3915 (N_3915,N_1682,N_1165);
and U3916 (N_3916,N_1786,N_1458);
or U3917 (N_3917,N_3031,N_1319);
and U3918 (N_3918,N_2567,N_1600);
nand U3919 (N_3919,N_795,N_2364);
nor U3920 (N_3920,N_2358,N_1578);
and U3921 (N_3921,N_3048,N_2126);
and U3922 (N_3922,N_1547,N_280);
or U3923 (N_3923,N_2618,N_204);
or U3924 (N_3924,N_2798,N_2401);
nor U3925 (N_3925,N_2180,N_1698);
nand U3926 (N_3926,N_876,N_51);
nor U3927 (N_3927,N_979,N_226);
or U3928 (N_3928,N_432,N_647);
nand U3929 (N_3929,N_2784,N_1164);
nand U3930 (N_3930,N_466,N_328);
xnor U3931 (N_3931,N_1860,N_2963);
nand U3932 (N_3932,N_563,N_1872);
nand U3933 (N_3933,N_520,N_1241);
nand U3934 (N_3934,N_375,N_2429);
nor U3935 (N_3935,N_1398,N_1810);
and U3936 (N_3936,N_1571,N_2780);
or U3937 (N_3937,N_2291,N_2725);
and U3938 (N_3938,N_2362,N_2852);
and U3939 (N_3939,N_2491,N_282);
or U3940 (N_3940,N_1461,N_354);
or U3941 (N_3941,N_1961,N_83);
nand U3942 (N_3942,N_1731,N_2773);
and U3943 (N_3943,N_386,N_1527);
nand U3944 (N_3944,N_1357,N_2407);
and U3945 (N_3945,N_1665,N_1800);
nor U3946 (N_3946,N_793,N_1332);
nor U3947 (N_3947,N_2845,N_2219);
nor U3948 (N_3948,N_829,N_2455);
and U3949 (N_3949,N_2320,N_1400);
nand U3950 (N_3950,N_1718,N_1904);
or U3951 (N_3951,N_505,N_2134);
and U3952 (N_3952,N_28,N_2091);
and U3953 (N_3953,N_1266,N_3052);
nand U3954 (N_3954,N_81,N_2370);
xnor U3955 (N_3955,N_1656,N_529);
nor U3956 (N_3956,N_1813,N_2530);
nand U3957 (N_3957,N_2428,N_2224);
nand U3958 (N_3958,N_981,N_2953);
nand U3959 (N_3959,N_61,N_2082);
and U3960 (N_3960,N_2459,N_746);
nor U3961 (N_3961,N_1188,N_2479);
nor U3962 (N_3962,N_1609,N_998);
or U3963 (N_3963,N_3006,N_1559);
nand U3964 (N_3964,N_2120,N_2855);
or U3965 (N_3965,N_1702,N_1779);
and U3966 (N_3966,N_2726,N_244);
and U3967 (N_3967,N_2399,N_2278);
nor U3968 (N_3968,N_1733,N_3096);
nor U3969 (N_3969,N_3022,N_786);
and U3970 (N_3970,N_1543,N_652);
xor U3971 (N_3971,N_755,N_1753);
and U3972 (N_3972,N_2422,N_502);
and U3973 (N_3973,N_2561,N_2781);
nand U3974 (N_3974,N_2612,N_2414);
nand U3975 (N_3975,N_1,N_769);
xor U3976 (N_3976,N_661,N_1177);
nor U3977 (N_3977,N_1853,N_1808);
or U3978 (N_3978,N_1459,N_1663);
and U3979 (N_3979,N_136,N_968);
nand U3980 (N_3980,N_378,N_962);
xnor U3981 (N_3981,N_2712,N_1137);
or U3982 (N_3982,N_1111,N_2346);
and U3983 (N_3983,N_798,N_195);
xnor U3984 (N_3984,N_238,N_1562);
or U3985 (N_3985,N_2,N_2045);
nor U3986 (N_3986,N_1912,N_3059);
or U3987 (N_3987,N_2476,N_410);
xnor U3988 (N_3988,N_972,N_485);
nor U3989 (N_3989,N_2043,N_1080);
or U3990 (N_3990,N_2389,N_1485);
and U3991 (N_3991,N_2230,N_2196);
nor U3992 (N_3992,N_2064,N_1035);
or U3993 (N_3993,N_165,N_2862);
xor U3994 (N_3994,N_1801,N_1003);
and U3995 (N_3995,N_2107,N_1321);
nand U3996 (N_3996,N_2300,N_2602);
or U3997 (N_3997,N_193,N_293);
nor U3998 (N_3998,N_302,N_930);
and U3999 (N_3999,N_2138,N_3065);
and U4000 (N_4000,N_348,N_2830);
nor U4001 (N_4001,N_336,N_72);
and U4002 (N_4002,N_2727,N_2619);
xor U4003 (N_4003,N_1162,N_1537);
and U4004 (N_4004,N_2622,N_543);
nand U4005 (N_4005,N_1655,N_257);
xor U4006 (N_4006,N_1339,N_2185);
nor U4007 (N_4007,N_1457,N_2465);
nor U4008 (N_4008,N_403,N_2382);
nand U4009 (N_4009,N_1598,N_2240);
nand U4010 (N_4010,N_1268,N_889);
and U4011 (N_4011,N_200,N_12);
nand U4012 (N_4012,N_430,N_2162);
nor U4013 (N_4013,N_2518,N_2173);
nand U4014 (N_4014,N_58,N_1480);
nor U4015 (N_4015,N_2720,N_1835);
and U4016 (N_4016,N_78,N_2199);
nor U4017 (N_4017,N_598,N_2055);
or U4018 (N_4018,N_199,N_964);
or U4019 (N_4019,N_276,N_36);
and U4020 (N_4020,N_1185,N_1012);
or U4021 (N_4021,N_714,N_513);
and U4022 (N_4022,N_1009,N_1939);
xnor U4023 (N_4023,N_2952,N_2381);
xor U4024 (N_4024,N_1360,N_722);
xnor U4025 (N_4025,N_1048,N_1700);
and U4026 (N_4026,N_1523,N_2061);
or U4027 (N_4027,N_947,N_1364);
nand U4028 (N_4028,N_982,N_1643);
and U4029 (N_4029,N_512,N_2292);
or U4030 (N_4030,N_1580,N_292);
and U4031 (N_4031,N_1406,N_1960);
and U4032 (N_4032,N_614,N_2262);
or U4033 (N_4033,N_2895,N_1384);
nand U4034 (N_4034,N_2504,N_2062);
or U4035 (N_4035,N_1125,N_2317);
and U4036 (N_4036,N_253,N_536);
nor U4037 (N_4037,N_2492,N_2366);
xnor U4038 (N_4038,N_440,N_635);
nor U4039 (N_4039,N_2367,N_862);
nor U4040 (N_4040,N_1089,N_95);
nand U4041 (N_4041,N_1923,N_2888);
and U4042 (N_4042,N_2912,N_1538);
or U4043 (N_4043,N_389,N_10);
nand U4044 (N_4044,N_1802,N_52);
or U4045 (N_4045,N_2052,N_2050);
nand U4046 (N_4046,N_710,N_2039);
nor U4047 (N_4047,N_1477,N_188);
or U4048 (N_4048,N_2116,N_1850);
or U4049 (N_4049,N_2533,N_2022);
nand U4050 (N_4050,N_1394,N_621);
or U4051 (N_4051,N_1690,N_734);
nor U4052 (N_4052,N_2081,N_2980);
or U4053 (N_4053,N_2501,N_1076);
nor U4054 (N_4054,N_1715,N_1103);
xor U4055 (N_4055,N_1940,N_794);
nand U4056 (N_4056,N_2336,N_2887);
or U4057 (N_4057,N_153,N_1052);
or U4058 (N_4058,N_1660,N_2683);
nor U4059 (N_4059,N_2885,N_376);
nand U4060 (N_4060,N_2085,N_2253);
nor U4061 (N_4061,N_3122,N_1010);
nand U4062 (N_4062,N_1295,N_133);
and U4063 (N_4063,N_868,N_1235);
nand U4064 (N_4064,N_1577,N_1687);
and U4065 (N_4065,N_1658,N_2639);
nor U4066 (N_4066,N_2265,N_1597);
or U4067 (N_4067,N_806,N_3070);
or U4068 (N_4068,N_615,N_2637);
nand U4069 (N_4069,N_1306,N_1402);
or U4070 (N_4070,N_270,N_278);
or U4071 (N_4071,N_1889,N_2673);
or U4072 (N_4072,N_2452,N_2633);
and U4073 (N_4073,N_2571,N_9);
nand U4074 (N_4074,N_2285,N_1842);
or U4075 (N_4075,N_2007,N_1987);
nor U4076 (N_4076,N_1290,N_2266);
nor U4077 (N_4077,N_2519,N_1763);
and U4078 (N_4078,N_1143,N_169);
and U4079 (N_4079,N_776,N_1752);
or U4080 (N_4080,N_2385,N_2943);
xor U4081 (N_4081,N_2338,N_472);
and U4082 (N_4082,N_1804,N_1985);
nor U4083 (N_4083,N_1855,N_1611);
nor U4084 (N_4084,N_495,N_435);
and U4085 (N_4085,N_131,N_2245);
or U4086 (N_4086,N_2212,N_451);
and U4087 (N_4087,N_2229,N_2685);
xnor U4088 (N_4088,N_907,N_2102);
xnor U4089 (N_4089,N_381,N_545);
nand U4090 (N_4090,N_29,N_3005);
nor U4091 (N_4091,N_885,N_2679);
xnor U4092 (N_4092,N_3016,N_1951);
and U4093 (N_4093,N_894,N_148);
or U4094 (N_4094,N_1039,N_367);
and U4095 (N_4095,N_569,N_2894);
xnor U4096 (N_4096,N_3021,N_965);
and U4097 (N_4097,N_1141,N_2609);
nand U4098 (N_4098,N_2330,N_1972);
xor U4099 (N_4099,N_43,N_1437);
xor U4100 (N_4100,N_1391,N_2915);
or U4101 (N_4101,N_379,N_198);
nor U4102 (N_4102,N_2139,N_1706);
nand U4103 (N_4103,N_595,N_1417);
nor U4104 (N_4104,N_657,N_2965);
and U4105 (N_4105,N_1343,N_1859);
nor U4106 (N_4106,N_2825,N_2077);
and U4107 (N_4107,N_490,N_2127);
nor U4108 (N_4108,N_2271,N_263);
xor U4109 (N_4109,N_434,N_2555);
nand U4110 (N_4110,N_2070,N_1272);
nand U4111 (N_4111,N_2249,N_648);
nor U4112 (N_4112,N_3028,N_1632);
nor U4113 (N_4113,N_1180,N_1849);
and U4114 (N_4114,N_2416,N_2288);
and U4115 (N_4115,N_2921,N_916);
nor U4116 (N_4116,N_84,N_523);
and U4117 (N_4117,N_983,N_368);
nor U4118 (N_4118,N_2089,N_2516);
or U4119 (N_4119,N_1422,N_2809);
or U4120 (N_4120,N_1411,N_1498);
nor U4121 (N_4121,N_881,N_2763);
nor U4122 (N_4122,N_2741,N_2057);
and U4123 (N_4123,N_801,N_311);
nor U4124 (N_4124,N_2998,N_2174);
and U4125 (N_4125,N_2109,N_2604);
nor U4126 (N_4126,N_1369,N_239);
or U4127 (N_4127,N_2636,N_1317);
and U4128 (N_4128,N_1607,N_2398);
and U4129 (N_4129,N_564,N_768);
nor U4130 (N_4130,N_550,N_1827);
and U4131 (N_4131,N_417,N_1021);
nor U4132 (N_4132,N_2558,N_2462);
or U4133 (N_4133,N_2467,N_1674);
or U4134 (N_4134,N_1445,N_1083);
nand U4135 (N_4135,N_2371,N_1397);
or U4136 (N_4136,N_547,N_3075);
or U4137 (N_4137,N_2296,N_2934);
nand U4138 (N_4138,N_642,N_987);
nor U4139 (N_4139,N_1425,N_3025);
nand U4140 (N_4140,N_431,N_1916);
nand U4141 (N_4141,N_2096,N_216);
and U4142 (N_4142,N_1085,N_1246);
or U4143 (N_4143,N_1957,N_309);
and U4144 (N_4144,N_2828,N_2166);
or U4145 (N_4145,N_7,N_2575);
nor U4146 (N_4146,N_103,N_2715);
or U4147 (N_4147,N_1434,N_1288);
or U4148 (N_4148,N_774,N_3014);
and U4149 (N_4149,N_2538,N_1479);
xor U4150 (N_4150,N_662,N_1929);
nand U4151 (N_4151,N_202,N_285);
and U4152 (N_4152,N_986,N_245);
nor U4153 (N_4153,N_638,N_2749);
nand U4154 (N_4154,N_64,N_284);
or U4155 (N_4155,N_1217,N_462);
or U4156 (N_4156,N_2794,N_3011);
nand U4157 (N_4157,N_517,N_214);
and U4158 (N_4158,N_2544,N_935);
xor U4159 (N_4159,N_2623,N_3061);
nor U4160 (N_4160,N_2928,N_2941);
and U4161 (N_4161,N_830,N_525);
nor U4162 (N_4162,N_1593,N_2150);
nand U4163 (N_4163,N_825,N_318);
xor U4164 (N_4164,N_2668,N_2806);
nor U4165 (N_4165,N_2801,N_1231);
or U4166 (N_4166,N_901,N_863);
and U4167 (N_4167,N_2453,N_527);
and U4168 (N_4168,N_2722,N_1057);
nand U4169 (N_4169,N_2329,N_2620);
and U4170 (N_4170,N_449,N_2461);
xnor U4171 (N_4171,N_1642,N_1335);
and U4172 (N_4172,N_939,N_492);
xor U4173 (N_4173,N_2136,N_2195);
nand U4174 (N_4174,N_1513,N_2969);
nand U4175 (N_4175,N_2425,N_1608);
and U4176 (N_4176,N_1584,N_577);
and U4177 (N_4177,N_332,N_1429);
and U4178 (N_4178,N_1213,N_1071);
xnor U4179 (N_4179,N_342,N_1756);
nor U4180 (N_4180,N_1497,N_1297);
nor U4181 (N_4181,N_3109,N_712);
nor U4182 (N_4182,N_2315,N_139);
and U4183 (N_4183,N_2739,N_294);
nand U4184 (N_4184,N_2261,N_909);
nor U4185 (N_4185,N_1880,N_2463);
nand U4186 (N_4186,N_1790,N_1094);
nor U4187 (N_4187,N_913,N_844);
or U4188 (N_4188,N_3030,N_1215);
and U4189 (N_4189,N_840,N_1522);
and U4190 (N_4190,N_1199,N_771);
and U4191 (N_4191,N_423,N_2898);
xor U4192 (N_4192,N_639,N_2645);
or U4193 (N_4193,N_108,N_2728);
nor U4194 (N_4194,N_2876,N_990);
nor U4195 (N_4195,N_2559,N_1937);
xor U4196 (N_4196,N_1768,N_888);
nor U4197 (N_4197,N_1789,N_2248);
or U4198 (N_4198,N_2841,N_2380);
nor U4199 (N_4199,N_2823,N_955);
and U4200 (N_4200,N_443,N_2534);
and U4201 (N_4201,N_820,N_2026);
and U4202 (N_4202,N_1181,N_1372);
nor U4203 (N_4203,N_883,N_1881);
and U4204 (N_4204,N_1025,N_2157);
and U4205 (N_4205,N_2767,N_1367);
nor U4206 (N_4206,N_2483,N_1251);
nor U4207 (N_4207,N_2846,N_455);
nand U4208 (N_4208,N_146,N_2731);
nand U4209 (N_4209,N_2874,N_1438);
or U4210 (N_4210,N_2539,N_1683);
and U4211 (N_4211,N_2037,N_1072);
nand U4212 (N_4212,N_1930,N_1770);
or U4213 (N_4213,N_185,N_3095);
xnor U4214 (N_4214,N_496,N_518);
or U4215 (N_4215,N_1534,N_2409);
nand U4216 (N_4216,N_2182,N_1712);
nand U4217 (N_4217,N_2709,N_1495);
nor U4218 (N_4218,N_1152,N_1861);
nand U4219 (N_4219,N_694,N_2119);
nor U4220 (N_4220,N_1158,N_15);
nor U4221 (N_4221,N_2332,N_1488);
nor U4222 (N_4222,N_2974,N_2387);
xor U4223 (N_4223,N_1784,N_2901);
xnor U4224 (N_4224,N_1899,N_2983);
or U4225 (N_4225,N_1166,N_2010);
or U4226 (N_4226,N_2938,N_1138);
nor U4227 (N_4227,N_3089,N_2796);
xnor U4228 (N_4228,N_2509,N_1549);
nand U4229 (N_4229,N_818,N_47);
nand U4230 (N_4230,N_2588,N_2444);
nand U4231 (N_4231,N_1077,N_1826);
nand U4232 (N_4232,N_2177,N_757);
and U4233 (N_4233,N_2024,N_2255);
or U4234 (N_4234,N_842,N_2112);
and U4235 (N_4235,N_1254,N_2449);
and U4236 (N_4236,N_79,N_731);
or U4237 (N_4237,N_3113,N_1509);
or U4238 (N_4238,N_2060,N_1129);
nand U4239 (N_4239,N_206,N_2202);
and U4240 (N_4240,N_2244,N_3037);
nand U4241 (N_4241,N_3123,N_2821);
nor U4242 (N_4242,N_1173,N_827);
and U4243 (N_4243,N_2149,N_2603);
xor U4244 (N_4244,N_2956,N_2760);
and U4245 (N_4245,N_841,N_1002);
nor U4246 (N_4246,N_954,N_404);
nand U4247 (N_4247,N_233,N_586);
or U4248 (N_4248,N_2118,N_999);
xor U4249 (N_4249,N_24,N_799);
or U4250 (N_4250,N_2807,N_2437);
or U4251 (N_4251,N_2886,N_1218);
nand U4252 (N_4252,N_835,N_2130);
and U4253 (N_4253,N_197,N_1622);
nor U4254 (N_4254,N_3013,N_2125);
and U4255 (N_4255,N_351,N_1701);
nor U4256 (N_4256,N_2864,N_1183);
nor U4257 (N_4257,N_1066,N_2277);
and U4258 (N_4258,N_2833,N_2925);
nor U4259 (N_4259,N_1749,N_1696);
nand U4260 (N_4260,N_558,N_2323);
xnor U4261 (N_4261,N_1095,N_312);
and U4262 (N_4262,N_1427,N_1340);
nor U4263 (N_4263,N_2529,N_2621);
or U4264 (N_4264,N_2616,N_2606);
or U4265 (N_4265,N_2316,N_346);
or U4266 (N_4266,N_566,N_2961);
or U4267 (N_4267,N_623,N_956);
nor U4268 (N_4268,N_1729,N_2856);
or U4269 (N_4269,N_655,N_1024);
or U4270 (N_4270,N_812,N_295);
nand U4271 (N_4271,N_2393,N_1206);
nor U4272 (N_4272,N_2579,N_212);
nor U4273 (N_4273,N_1678,N_2614);
or U4274 (N_4274,N_645,N_2111);
nand U4275 (N_4275,N_1433,N_2446);
and U4276 (N_4276,N_1758,N_2770);
nor U4277 (N_4277,N_2573,N_392);
xor U4278 (N_4278,N_2004,N_2799);
and U4279 (N_4279,N_1759,N_940);
nand U4280 (N_4280,N_759,N_1128);
and U4281 (N_4281,N_2701,N_594);
xnor U4282 (N_4282,N_1176,N_363);
or U4283 (N_4283,N_213,N_707);
or U4284 (N_4284,N_1278,N_167);
and U4285 (N_4285,N_3078,N_1107);
and U4286 (N_4286,N_1499,N_1302);
or U4287 (N_4287,N_1602,N_1841);
nor U4288 (N_4288,N_1258,N_385);
nor U4289 (N_4289,N_2790,N_2788);
or U4290 (N_4290,N_2873,N_1494);
nand U4291 (N_4291,N_1440,N_164);
nand U4292 (N_4292,N_1186,N_1848);
nor U4293 (N_4293,N_335,N_1587);
nand U4294 (N_4294,N_2583,N_221);
or U4295 (N_4295,N_864,N_2499);
xor U4296 (N_4296,N_359,N_2392);
or U4297 (N_4297,N_112,N_1843);
nor U4298 (N_4298,N_1336,N_2443);
and U4299 (N_4299,N_130,N_1410);
nand U4300 (N_4300,N_1528,N_2221);
nand U4301 (N_4301,N_2879,N_94);
nand U4302 (N_4302,N_3032,N_2068);
nand U4303 (N_4303,N_2644,N_867);
xor U4304 (N_4304,N_1202,N_2488);
and U4305 (N_4305,N_1695,N_1828);
and U4306 (N_4306,N_16,N_1250);
or U4307 (N_4307,N_927,N_2660);
xnor U4308 (N_4308,N_157,N_1023);
xnor U4309 (N_4309,N_1570,N_298);
nor U4310 (N_4310,N_330,N_1647);
xor U4311 (N_4311,N_2708,N_3087);
nor U4312 (N_4312,N_1807,N_1131);
nand U4313 (N_4313,N_991,N_959);
or U4314 (N_4314,N_1893,N_135);
nor U4315 (N_4315,N_1962,N_1918);
and U4316 (N_4316,N_2866,N_2624);
nor U4317 (N_4317,N_796,N_2318);
and U4318 (N_4318,N_2836,N_750);
nand U4319 (N_4319,N_2868,N_395);
and U4320 (N_4320,N_1603,N_2450);
and U4321 (N_4321,N_1575,N_2215);
nand U4322 (N_4322,N_355,N_1232);
xor U4323 (N_4323,N_1067,N_1532);
and U4324 (N_4324,N_1492,N_2348);
nand U4325 (N_4325,N_2522,N_880);
nor U4326 (N_4326,N_1624,N_1443);
nor U4327 (N_4327,N_1474,N_3);
xor U4328 (N_4328,N_574,N_641);
nand U4329 (N_4329,N_1257,N_144);
and U4330 (N_4330,N_3121,N_49);
nor U4331 (N_4331,N_559,N_3115);
and U4332 (N_4332,N_1204,N_996);
and U4333 (N_4333,N_681,N_343);
xnor U4334 (N_4334,N_2611,N_1975);
and U4335 (N_4335,N_666,N_1169);
xor U4336 (N_4336,N_3041,N_2515);
xor U4337 (N_4337,N_480,N_1436);
nor U4338 (N_4338,N_2835,N_1969);
or U4339 (N_4339,N_479,N_1046);
nand U4340 (N_4340,N_2225,N_73);
and U4341 (N_4341,N_2768,N_1123);
or U4342 (N_4342,N_2505,N_2421);
nor U4343 (N_4343,N_2200,N_2657);
xor U4344 (N_4344,N_2906,N_2101);
nand U4345 (N_4345,N_3110,N_1142);
and U4346 (N_4346,N_1738,N_2243);
xor U4347 (N_4347,N_2258,N_1252);
xnor U4348 (N_4348,N_1244,N_445);
nand U4349 (N_4349,N_349,N_460);
nor U4350 (N_4350,N_1617,N_1942);
or U4351 (N_4351,N_1256,N_1320);
xor U4352 (N_4352,N_2098,N_74);
and U4353 (N_4353,N_1728,N_2133);
xor U4354 (N_4354,N_264,N_2896);
nand U4355 (N_4355,N_1788,N_3050);
nand U4356 (N_4356,N_1871,N_2546);
or U4357 (N_4357,N_134,N_2008);
and U4358 (N_4358,N_926,N_2020);
or U4359 (N_4359,N_2853,N_1650);
or U4360 (N_4360,N_2402,N_1754);
and U4361 (N_4361,N_1018,N_1943);
nand U4362 (N_4362,N_809,N_1685);
and U4363 (N_4363,N_1115,N_2847);
nand U4364 (N_4364,N_1101,N_1711);
nor U4365 (N_4365,N_2854,N_2267);
or U4366 (N_4366,N_2756,N_1284);
and U4367 (N_4367,N_279,N_2337);
or U4368 (N_4368,N_53,N_814);
or U4369 (N_4369,N_2235,N_698);
nor U4370 (N_4370,N_2711,N_1091);
or U4371 (N_4371,N_2869,N_1454);
nand U4372 (N_4372,N_326,N_26);
or U4373 (N_4373,N_2697,N_2511);
nor U4374 (N_4374,N_2521,N_3120);
or U4375 (N_4375,N_578,N_910);
or U4376 (N_4376,N_1764,N_262);
and U4377 (N_4377,N_2849,N_834);
or U4378 (N_4378,N_1517,N_2495);
nor U4379 (N_4379,N_1441,N_2131);
nor U4380 (N_4380,N_2714,N_1126);
and U4381 (N_4381,N_2814,N_1525);
and U4382 (N_4382,N_453,N_674);
and U4383 (N_4383,N_353,N_2105);
nand U4384 (N_4384,N_1997,N_2578);
nand U4385 (N_4385,N_1999,N_1778);
and U4386 (N_4386,N_2308,N_196);
nor U4387 (N_4387,N_1857,N_2986);
nor U4388 (N_4388,N_1063,N_2198);
and U4389 (N_4389,N_2211,N_1265);
and U4390 (N_4390,N_266,N_476);
nor U4391 (N_4391,N_382,N_1610);
xnor U4392 (N_4392,N_1862,N_2494);
or U4393 (N_4393,N_2907,N_1540);
nand U4394 (N_4394,N_1184,N_887);
nand U4395 (N_4395,N_248,N_3100);
nand U4396 (N_4396,N_2716,N_1820);
nor U4397 (N_4397,N_504,N_643);
nand U4398 (N_4398,N_405,N_2503);
xnor U4399 (N_4399,N_849,N_1766);
nor U4400 (N_4400,N_2834,N_2153);
nor U4401 (N_4401,N_1743,N_1967);
nor U4402 (N_4402,N_35,N_2373);
nand U4403 (N_4403,N_2706,N_2684);
nor U4404 (N_4404,N_1897,N_2122);
nor U4405 (N_4405,N_2205,N_588);
nand U4406 (N_4406,N_2513,N_1453);
or U4407 (N_4407,N_1680,N_1264);
nor U4408 (N_4408,N_2932,N_1884);
nor U4409 (N_4409,N_1590,N_2397);
nor U4410 (N_4410,N_2747,N_413);
nand U4411 (N_4411,N_1530,N_406);
nor U4412 (N_4412,N_1691,N_8);
xor U4413 (N_4413,N_751,N_2721);
and U4414 (N_4414,N_715,N_1104);
and U4415 (N_4415,N_1421,N_2914);
nor U4416 (N_4416,N_535,N_265);
or U4417 (N_4417,N_1187,N_1958);
xor U4418 (N_4418,N_2121,N_2129);
or U4419 (N_4419,N_2700,N_770);
nand U4420 (N_4420,N_273,N_2260);
nor U4421 (N_4421,N_111,N_3010);
nor U4422 (N_4422,N_1644,N_1824);
and U4423 (N_4423,N_473,N_2054);
and U4424 (N_4424,N_1946,N_730);
and U4425 (N_4425,N_1007,N_953);
xnor U4426 (N_4426,N_1661,N_2352);
and U4427 (N_4427,N_459,N_1191);
and U4428 (N_4428,N_1469,N_2877);
nor U4429 (N_4429,N_369,N_1908);
nor U4430 (N_4430,N_1475,N_860);
nor U4431 (N_4431,N_2625,N_1405);
nand U4432 (N_4432,N_3015,N_2787);
nor U4433 (N_4433,N_1133,N_1671);
and U4434 (N_4434,N_1451,N_1994);
or U4435 (N_4435,N_1905,N_506);
xnor U4436 (N_4436,N_2328,N_2438);
xor U4437 (N_4437,N_696,N_393);
nor U4438 (N_4438,N_948,N_3017);
nor U4439 (N_4439,N_700,N_2968);
or U4440 (N_4440,N_63,N_156);
nand U4441 (N_4441,N_1721,N_567);
or U4442 (N_4442,N_688,N_1056);
and U4443 (N_4443,N_2014,N_1484);
and U4444 (N_4444,N_2360,N_2600);
nand U4445 (N_4445,N_942,N_2021);
nor U4446 (N_4446,N_421,N_2964);
or U4447 (N_4447,N_765,N_754);
or U4448 (N_4448,N_3092,N_2400);
and U4449 (N_4449,N_932,N_720);
nor U4450 (N_4450,N_327,N_539);
nand U4451 (N_4451,N_2103,N_853);
and U4452 (N_4452,N_610,N_2591);
nand U4453 (N_4453,N_1289,N_2451);
nor U4454 (N_4454,N_272,N_709);
xor U4455 (N_4455,N_906,N_2349);
or U4456 (N_4456,N_223,N_3081);
and U4457 (N_4457,N_1998,N_42);
nand U4458 (N_4458,N_2694,N_1345);
and U4459 (N_4459,N_2213,N_1863);
nor U4460 (N_4460,N_752,N_1771);
or U4461 (N_4461,N_1954,N_2565);
nand U4462 (N_4462,N_2341,N_352);
nor U4463 (N_4463,N_3003,N_220);
and U4464 (N_4464,N_2069,N_1464);
nor U4465 (N_4465,N_2735,N_1667);
nor U4466 (N_4466,N_1098,N_1239);
or U4467 (N_4467,N_2649,N_1794);
nor U4468 (N_4468,N_149,N_1496);
and U4469 (N_4469,N_845,N_2033);
nand U4470 (N_4470,N_839,N_3044);
nor U4471 (N_4471,N_2339,N_620);
and U4472 (N_4472,N_571,N_2688);
and U4473 (N_4473,N_2095,N_528);
or U4474 (N_4474,N_1356,N_101);
and U4475 (N_4475,N_1105,N_1520);
nand U4476 (N_4476,N_1004,N_1854);
nor U4477 (N_4477,N_2013,N_159);
or U4478 (N_4478,N_555,N_1314);
xnor U4479 (N_4479,N_1207,N_2903);
or U4480 (N_4480,N_1030,N_908);
xor U4481 (N_4481,N_2772,N_1127);
nand U4482 (N_4482,N_2562,N_25);
and U4483 (N_4483,N_122,N_2908);
nor U4484 (N_4484,N_637,N_3040);
nor U4485 (N_4485,N_1140,N_67);
nor U4486 (N_4486,N_2793,N_5);
or U4487 (N_4487,N_3076,N_1396);
nand U4488 (N_4488,N_179,N_3056);
or U4489 (N_4489,N_2663,N_1500);
or U4490 (N_4490,N_268,N_1681);
and U4491 (N_4491,N_1502,N_1363);
nand U4492 (N_4492,N_1747,N_2904);
and U4493 (N_4493,N_2208,N_602);
nand U4494 (N_4494,N_2431,N_2661);
xor U4495 (N_4495,N_1704,N_2030);
or U4496 (N_4496,N_1439,N_2110);
nand U4497 (N_4497,N_1552,N_884);
and U4498 (N_4498,N_978,N_584);
or U4499 (N_4499,N_132,N_1761);
nor U4500 (N_4500,N_920,N_589);
nor U4501 (N_4501,N_2357,N_1082);
xor U4502 (N_4502,N_1606,N_2880);
nand U4503 (N_4503,N_1365,N_669);
and U4504 (N_4504,N_1390,N_613);
or U4505 (N_4505,N_2671,N_1947);
nor U4506 (N_4506,N_2167,N_1757);
and U4507 (N_4507,N_772,N_2237);
and U4508 (N_4508,N_1654,N_1087);
and U4509 (N_4509,N_56,N_2545);
nand U4510 (N_4510,N_573,N_847);
and U4511 (N_4511,N_1466,N_663);
nor U4512 (N_4512,N_644,N_2765);
or U4513 (N_4513,N_2093,N_1866);
or U4514 (N_4514,N_1008,N_1462);
nand U4515 (N_4515,N_2557,N_236);
nand U4516 (N_4516,N_2441,N_1652);
or U4517 (N_4517,N_1612,N_18);
nand U4518 (N_4518,N_2222,N_2605);
and U4519 (N_4519,N_1628,N_2137);
or U4520 (N_4520,N_2837,N_1139);
or U4521 (N_4521,N_123,N_2883);
and U4522 (N_4522,N_2707,N_2156);
nand U4523 (N_4523,N_2576,N_2550);
and U4524 (N_4524,N_1001,N_1342);
and U4525 (N_4525,N_2263,N_1865);
nor U4526 (N_4526,N_3045,N_3107);
xor U4527 (N_4527,N_1554,N_2269);
xnor U4528 (N_4528,N_341,N_218);
nand U4529 (N_4529,N_1301,N_686);
nor U4530 (N_4530,N_1900,N_2710);
and U4531 (N_4531,N_1037,N_1240);
and U4532 (N_4532,N_2223,N_1615);
and U4533 (N_4533,N_256,N_1380);
and U4534 (N_4534,N_2699,N_2517);
nor U4535 (N_4535,N_1546,N_1762);
and U4536 (N_4536,N_1374,N_1705);
nor U4537 (N_4537,N_1507,N_1915);
and U4538 (N_4538,N_1223,N_1531);
and U4539 (N_4539,N_3108,N_2114);
nor U4540 (N_4540,N_606,N_1368);
or U4541 (N_4541,N_2507,N_1551);
xnor U4542 (N_4542,N_994,N_1193);
nand U4543 (N_4543,N_274,N_1555);
and U4544 (N_4544,N_2695,N_2490);
and U4545 (N_4545,N_1932,N_178);
nand U4546 (N_4546,N_3001,N_407);
nor U4547 (N_4547,N_531,N_2498);
or U4548 (N_4548,N_2283,N_2553);
nor U4549 (N_4549,N_2703,N_205);
xor U4550 (N_4550,N_394,N_59);
and U4551 (N_4551,N_2742,N_2819);
nor U4552 (N_4552,N_604,N_1473);
nor U4553 (N_4553,N_1907,N_3043);
nand U4554 (N_4554,N_1596,N_519);
nor U4555 (N_4555,N_2526,N_76);
nand U4556 (N_4556,N_303,N_893);
xnor U4557 (N_4557,N_2572,N_2962);
or U4558 (N_4558,N_2598,N_1938);
or U4559 (N_4559,N_1955,N_2654);
nand U4560 (N_4560,N_2388,N_764);
and U4561 (N_4561,N_508,N_524);
nor U4562 (N_4562,N_2791,N_813);
nor U4563 (N_4563,N_2169,N_3091);
nor U4564 (N_4564,N_3111,N_1491);
nand U4565 (N_4565,N_454,N_1435);
nand U4566 (N_4566,N_2996,N_416);
nor U4567 (N_4567,N_810,N_2005);
nand U4568 (N_4568,N_1032,N_113);
nand U4569 (N_4569,N_718,N_1490);
nor U4570 (N_4570,N_989,N_2086);
nor U4571 (N_4571,N_1568,N_1614);
or U4572 (N_4572,N_2378,N_2356);
or U4573 (N_4573,N_1348,N_1062);
nor U4574 (N_4574,N_2209,N_86);
nand U4575 (N_4575,N_1673,N_2191);
nor U4576 (N_4576,N_1980,N_1913);
and U4577 (N_4577,N_2802,N_1797);
nand U4578 (N_4578,N_656,N_2734);
xor U4579 (N_4579,N_2737,N_1382);
and U4580 (N_4580,N_874,N_922);
nand U4581 (N_4581,N_321,N_1726);
xnor U4582 (N_4582,N_1649,N_1392);
nor U4583 (N_4583,N_1851,N_850);
nor U4584 (N_4584,N_684,N_739);
and U4585 (N_4585,N_1097,N_1657);
nor U4586 (N_4586,N_2988,N_1641);
or U4587 (N_4587,N_2031,N_1408);
nor U4588 (N_4588,N_2655,N_900);
nor U4589 (N_4589,N_1934,N_1358);
nand U4590 (N_4590,N_1285,N_107);
and U4591 (N_4591,N_3104,N_551);
and U4592 (N_4592,N_514,N_2891);
nand U4593 (N_4593,N_1689,N_557);
nor U4594 (N_4594,N_805,N_2354);
nand U4595 (N_4595,N_2408,N_2099);
nand U4596 (N_4596,N_62,N_1684);
xnor U4597 (N_4597,N_23,N_2935);
nand U4598 (N_4598,N_1776,N_1122);
nor U4599 (N_4599,N_2789,N_2324);
or U4600 (N_4600,N_2067,N_3079);
xor U4601 (N_4601,N_1156,N_2140);
and U4602 (N_4602,N_1992,N_2859);
nand U4603 (N_4603,N_1324,N_1350);
nand U4604 (N_4604,N_1877,N_1120);
nand U4605 (N_4605,N_1668,N_2652);
or U4606 (N_4606,N_2309,N_2363);
and U4607 (N_4607,N_1519,N_2053);
nand U4608 (N_4608,N_705,N_915);
nor U4609 (N_4609,N_2090,N_2510);
nor U4610 (N_4610,N_1017,N_1709);
and U4611 (N_4611,N_408,N_1476);
and U4612 (N_4612,N_3116,N_2882);
and U4613 (N_4613,N_2135,N_3094);
or U4614 (N_4614,N_1783,N_2850);
nand U4615 (N_4615,N_532,N_1873);
or U4616 (N_4616,N_228,N_150);
nor U4617 (N_4617,N_374,N_377);
and U4618 (N_4618,N_977,N_1047);
or U4619 (N_4619,N_286,N_1447);
or U4620 (N_4620,N_151,N_692);
or U4621 (N_4621,N_1220,N_481);
nand U4622 (N_4622,N_756,N_728);
and U4623 (N_4623,N_486,N_331);
and U4624 (N_4624,N_32,N_1261);
nand U4625 (N_4625,N_1093,N_1945);
xnor U4626 (N_4626,N_2203,N_2404);
nand U4627 (N_4627,N_697,N_938);
nor U4628 (N_4628,N_2239,N_2355);
nand U4629 (N_4629,N_921,N_1233);
nand U4630 (N_4630,N_2990,N_3098);
and U4631 (N_4631,N_668,N_630);
nor U4632 (N_4632,N_210,N_664);
nand U4633 (N_4633,N_1051,N_93);
or U4634 (N_4634,N_2217,N_182);
nand U4635 (N_4635,N_3034,N_763);
nand U4636 (N_4636,N_290,N_2350);
or U4637 (N_4637,N_670,N_2981);
nand U4638 (N_4638,N_789,N_1049);
or U4639 (N_4639,N_2179,N_13);
nand U4640 (N_4640,N_34,N_2997);
and U4641 (N_4641,N_398,N_2497);
and U4642 (N_4642,N_1765,N_2046);
xor U4643 (N_4643,N_784,N_2597);
nor U4644 (N_4644,N_2270,N_748);
nand U4645 (N_4645,N_1885,N_819);
xor U4646 (N_4646,N_120,N_1620);
and U4647 (N_4647,N_2100,N_562);
nor U4648 (N_4648,N_1331,N_187);
or U4649 (N_4649,N_2464,N_787);
nor U4650 (N_4650,N_155,N_3063);
and U4651 (N_4651,N_300,N_1745);
nor U4652 (N_4652,N_2569,N_2580);
and U4653 (N_4653,N_969,N_1692);
and U4654 (N_4654,N_1132,N_1576);
nor U4655 (N_4655,N_48,N_1155);
or U4656 (N_4656,N_456,N_1312);
nand U4657 (N_4657,N_1404,N_522);
and U4658 (N_4658,N_2667,N_1544);
nor U4659 (N_4659,N_415,N_2817);
and U4660 (N_4660,N_3088,N_882);
and U4661 (N_4661,N_1512,N_102);
or U4662 (N_4662,N_782,N_2141);
or U4663 (N_4663,N_1694,N_2593);
nor U4664 (N_4664,N_622,N_2831);
and U4665 (N_4665,N_258,N_687);
and U4666 (N_4666,N_2863,N_1282);
nor U4667 (N_4667,N_851,N_1996);
nand U4668 (N_4668,N_447,N_2871);
and U4669 (N_4669,N_1737,N_2857);
nor U4670 (N_4670,N_308,N_1329);
and U4671 (N_4671,N_2978,N_973);
xor U4672 (N_4672,N_44,N_77);
or U4673 (N_4673,N_1818,N_724);
or U4674 (N_4674,N_1639,N_2584);
or U4675 (N_4675,N_677,N_235);
or U4676 (N_4676,N_2035,N_949);
or U4677 (N_4677,N_75,N_2218);
or U4678 (N_4678,N_515,N_747);
nor U4679 (N_4679,N_3053,N_2286);
or U4680 (N_4680,N_194,N_1259);
and U4681 (N_4681,N_1027,N_762);
nor U4682 (N_4682,N_2319,N_1248);
and U4683 (N_4683,N_2040,N_315);
nor U4684 (N_4684,N_2705,N_2556);
nor U4685 (N_4685,N_2274,N_2353);
nand U4686 (N_4686,N_1625,N_411);
and U4687 (N_4687,N_322,N_2192);
nor U4688 (N_4688,N_1486,N_26);
and U4689 (N_4689,N_2023,N_961);
or U4690 (N_4690,N_1831,N_514);
xor U4691 (N_4691,N_2137,N_1419);
nor U4692 (N_4692,N_659,N_2311);
nand U4693 (N_4693,N_3008,N_346);
nor U4694 (N_4694,N_2144,N_1565);
or U4695 (N_4695,N_2560,N_513);
and U4696 (N_4696,N_1843,N_1286);
nor U4697 (N_4697,N_1477,N_1388);
or U4698 (N_4698,N_2908,N_1586);
nand U4699 (N_4699,N_1315,N_1477);
and U4700 (N_4700,N_1552,N_1134);
or U4701 (N_4701,N_141,N_1667);
xnor U4702 (N_4702,N_370,N_217);
and U4703 (N_4703,N_331,N_1767);
nand U4704 (N_4704,N_1355,N_943);
nor U4705 (N_4705,N_1049,N_2166);
or U4706 (N_4706,N_811,N_316);
and U4707 (N_4707,N_604,N_317);
nor U4708 (N_4708,N_2757,N_2297);
nand U4709 (N_4709,N_2365,N_1186);
nand U4710 (N_4710,N_2319,N_2682);
or U4711 (N_4711,N_958,N_672);
nand U4712 (N_4712,N_629,N_990);
and U4713 (N_4713,N_2983,N_3041);
and U4714 (N_4714,N_2706,N_1741);
xnor U4715 (N_4715,N_1813,N_2261);
nor U4716 (N_4716,N_599,N_1596);
nor U4717 (N_4717,N_1772,N_2129);
or U4718 (N_4718,N_2632,N_1717);
nand U4719 (N_4719,N_303,N_839);
or U4720 (N_4720,N_2722,N_1223);
xnor U4721 (N_4721,N_1581,N_350);
nor U4722 (N_4722,N_1205,N_283);
xnor U4723 (N_4723,N_1840,N_644);
nor U4724 (N_4724,N_805,N_2405);
and U4725 (N_4725,N_1983,N_1716);
or U4726 (N_4726,N_2792,N_1879);
nand U4727 (N_4727,N_2399,N_2180);
or U4728 (N_4728,N_1059,N_583);
nand U4729 (N_4729,N_1469,N_1729);
nand U4730 (N_4730,N_1660,N_1668);
nor U4731 (N_4731,N_3030,N_2725);
xnor U4732 (N_4732,N_6,N_1441);
xnor U4733 (N_4733,N_16,N_137);
nand U4734 (N_4734,N_883,N_2079);
nor U4735 (N_4735,N_2685,N_1255);
nor U4736 (N_4736,N_2080,N_532);
nor U4737 (N_4737,N_2009,N_2795);
and U4738 (N_4738,N_2348,N_2005);
and U4739 (N_4739,N_88,N_2611);
or U4740 (N_4740,N_994,N_668);
or U4741 (N_4741,N_2800,N_2840);
xor U4742 (N_4742,N_108,N_1209);
and U4743 (N_4743,N_1065,N_2294);
or U4744 (N_4744,N_1381,N_1915);
and U4745 (N_4745,N_2674,N_2615);
xnor U4746 (N_4746,N_2589,N_2968);
and U4747 (N_4747,N_755,N_2249);
nand U4748 (N_4748,N_18,N_3052);
nor U4749 (N_4749,N_456,N_855);
nand U4750 (N_4750,N_1683,N_2994);
or U4751 (N_4751,N_375,N_2419);
and U4752 (N_4752,N_2724,N_827);
nand U4753 (N_4753,N_1798,N_614);
and U4754 (N_4754,N_1697,N_1461);
xor U4755 (N_4755,N_1053,N_2443);
nor U4756 (N_4756,N_1090,N_409);
or U4757 (N_4757,N_2277,N_1518);
nor U4758 (N_4758,N_123,N_187);
nor U4759 (N_4759,N_1768,N_1955);
and U4760 (N_4760,N_2559,N_716);
or U4761 (N_4761,N_1944,N_1789);
nand U4762 (N_4762,N_1359,N_2307);
or U4763 (N_4763,N_2936,N_1777);
and U4764 (N_4764,N_977,N_420);
nor U4765 (N_4765,N_489,N_944);
nor U4766 (N_4766,N_2887,N_1951);
nand U4767 (N_4767,N_1348,N_1009);
nor U4768 (N_4768,N_2839,N_817);
or U4769 (N_4769,N_2046,N_1194);
nor U4770 (N_4770,N_502,N_2641);
and U4771 (N_4771,N_1175,N_725);
and U4772 (N_4772,N_2197,N_86);
xnor U4773 (N_4773,N_1103,N_629);
and U4774 (N_4774,N_361,N_1050);
and U4775 (N_4775,N_356,N_1422);
nor U4776 (N_4776,N_2173,N_445);
or U4777 (N_4777,N_1869,N_2782);
nand U4778 (N_4778,N_3075,N_1948);
nor U4779 (N_4779,N_2041,N_2067);
nor U4780 (N_4780,N_2926,N_2643);
or U4781 (N_4781,N_1735,N_150);
nand U4782 (N_4782,N_864,N_323);
nand U4783 (N_4783,N_2833,N_1689);
nand U4784 (N_4784,N_1645,N_1525);
and U4785 (N_4785,N_2820,N_178);
nor U4786 (N_4786,N_2967,N_2135);
or U4787 (N_4787,N_1549,N_2813);
nand U4788 (N_4788,N_1884,N_167);
nand U4789 (N_4789,N_73,N_225);
nand U4790 (N_4790,N_1549,N_631);
nor U4791 (N_4791,N_1236,N_1368);
nand U4792 (N_4792,N_2706,N_1931);
or U4793 (N_4793,N_191,N_2257);
or U4794 (N_4794,N_2413,N_137);
nand U4795 (N_4795,N_55,N_1198);
nor U4796 (N_4796,N_748,N_3104);
or U4797 (N_4797,N_3065,N_1567);
and U4798 (N_4798,N_2530,N_2181);
and U4799 (N_4799,N_819,N_2836);
nor U4800 (N_4800,N_1681,N_960);
nand U4801 (N_4801,N_1441,N_1432);
and U4802 (N_4802,N_2796,N_2706);
or U4803 (N_4803,N_242,N_2779);
or U4804 (N_4804,N_3061,N_1418);
xor U4805 (N_4805,N_1256,N_958);
and U4806 (N_4806,N_1340,N_602);
or U4807 (N_4807,N_336,N_2646);
nand U4808 (N_4808,N_1490,N_1100);
nor U4809 (N_4809,N_1930,N_2727);
or U4810 (N_4810,N_3090,N_2339);
nand U4811 (N_4811,N_283,N_1326);
or U4812 (N_4812,N_613,N_1586);
nor U4813 (N_4813,N_1065,N_395);
or U4814 (N_4814,N_394,N_835);
nand U4815 (N_4815,N_474,N_2167);
nor U4816 (N_4816,N_1727,N_719);
nand U4817 (N_4817,N_3035,N_1033);
xnor U4818 (N_4818,N_2836,N_456);
xor U4819 (N_4819,N_1245,N_2753);
nor U4820 (N_4820,N_777,N_2857);
and U4821 (N_4821,N_1201,N_2072);
nand U4822 (N_4822,N_541,N_596);
and U4823 (N_4823,N_353,N_129);
nand U4824 (N_4824,N_2631,N_3046);
and U4825 (N_4825,N_3002,N_2974);
and U4826 (N_4826,N_1947,N_244);
nand U4827 (N_4827,N_2793,N_2417);
and U4828 (N_4828,N_1873,N_183);
or U4829 (N_4829,N_1653,N_1957);
nor U4830 (N_4830,N_348,N_1141);
and U4831 (N_4831,N_2139,N_59);
nor U4832 (N_4832,N_1621,N_2883);
or U4833 (N_4833,N_395,N_2373);
nor U4834 (N_4834,N_2352,N_2925);
xor U4835 (N_4835,N_1989,N_1836);
nand U4836 (N_4836,N_1204,N_2410);
or U4837 (N_4837,N_2319,N_2848);
or U4838 (N_4838,N_1440,N_1717);
nor U4839 (N_4839,N_1015,N_1764);
and U4840 (N_4840,N_1765,N_532);
xor U4841 (N_4841,N_1816,N_2174);
or U4842 (N_4842,N_2509,N_28);
and U4843 (N_4843,N_1777,N_1891);
nand U4844 (N_4844,N_1750,N_2380);
nand U4845 (N_4845,N_2113,N_970);
nand U4846 (N_4846,N_1727,N_594);
nor U4847 (N_4847,N_870,N_1380);
nand U4848 (N_4848,N_1056,N_1349);
and U4849 (N_4849,N_1055,N_1321);
or U4850 (N_4850,N_403,N_1199);
and U4851 (N_4851,N_2093,N_951);
nor U4852 (N_4852,N_290,N_443);
or U4853 (N_4853,N_2201,N_2127);
nor U4854 (N_4854,N_2058,N_1756);
nor U4855 (N_4855,N_829,N_2876);
nand U4856 (N_4856,N_1468,N_345);
or U4857 (N_4857,N_1116,N_1299);
nor U4858 (N_4858,N_2513,N_751);
or U4859 (N_4859,N_2466,N_2823);
nand U4860 (N_4860,N_789,N_794);
or U4861 (N_4861,N_2546,N_84);
and U4862 (N_4862,N_2537,N_87);
nor U4863 (N_4863,N_457,N_684);
xor U4864 (N_4864,N_961,N_1962);
or U4865 (N_4865,N_558,N_839);
or U4866 (N_4866,N_2131,N_2792);
or U4867 (N_4867,N_1996,N_459);
and U4868 (N_4868,N_2925,N_79);
xor U4869 (N_4869,N_2616,N_1150);
nand U4870 (N_4870,N_851,N_625);
or U4871 (N_4871,N_1214,N_1724);
nor U4872 (N_4872,N_2668,N_310);
and U4873 (N_4873,N_1638,N_82);
nor U4874 (N_4874,N_413,N_2015);
nor U4875 (N_4875,N_1926,N_904);
nor U4876 (N_4876,N_418,N_1181);
nand U4877 (N_4877,N_1929,N_1506);
and U4878 (N_4878,N_1553,N_866);
or U4879 (N_4879,N_1056,N_1958);
and U4880 (N_4880,N_1745,N_1775);
and U4881 (N_4881,N_38,N_2264);
nor U4882 (N_4882,N_479,N_2900);
nor U4883 (N_4883,N_740,N_1358);
nor U4884 (N_4884,N_2812,N_620);
nand U4885 (N_4885,N_2096,N_822);
nand U4886 (N_4886,N_1025,N_2997);
xor U4887 (N_4887,N_877,N_2523);
and U4888 (N_4888,N_938,N_37);
nand U4889 (N_4889,N_2294,N_1945);
and U4890 (N_4890,N_1025,N_1844);
and U4891 (N_4891,N_899,N_925);
xnor U4892 (N_4892,N_445,N_2379);
and U4893 (N_4893,N_364,N_936);
nor U4894 (N_4894,N_194,N_1669);
and U4895 (N_4895,N_3093,N_731);
or U4896 (N_4896,N_451,N_2701);
or U4897 (N_4897,N_2123,N_1398);
and U4898 (N_4898,N_337,N_2979);
nand U4899 (N_4899,N_1855,N_2196);
or U4900 (N_4900,N_446,N_2058);
nand U4901 (N_4901,N_1683,N_189);
xnor U4902 (N_4902,N_2889,N_2365);
or U4903 (N_4903,N_745,N_288);
xor U4904 (N_4904,N_1480,N_1384);
nand U4905 (N_4905,N_544,N_617);
nand U4906 (N_4906,N_1037,N_939);
or U4907 (N_4907,N_2529,N_3084);
nand U4908 (N_4908,N_2946,N_2859);
nor U4909 (N_4909,N_634,N_2635);
and U4910 (N_4910,N_3045,N_3039);
and U4911 (N_4911,N_1502,N_1971);
and U4912 (N_4912,N_2044,N_1942);
and U4913 (N_4913,N_964,N_2317);
nor U4914 (N_4914,N_2090,N_501);
and U4915 (N_4915,N_2154,N_1560);
and U4916 (N_4916,N_2763,N_617);
or U4917 (N_4917,N_1810,N_715);
nand U4918 (N_4918,N_3,N_1807);
or U4919 (N_4919,N_700,N_2980);
and U4920 (N_4920,N_509,N_907);
or U4921 (N_4921,N_579,N_2090);
nor U4922 (N_4922,N_374,N_1777);
nand U4923 (N_4923,N_1123,N_1823);
and U4924 (N_4924,N_1073,N_3067);
nand U4925 (N_4925,N_1622,N_2004);
nor U4926 (N_4926,N_1179,N_2445);
or U4927 (N_4927,N_1236,N_1199);
and U4928 (N_4928,N_505,N_28);
nand U4929 (N_4929,N_1955,N_281);
nand U4930 (N_4930,N_447,N_1739);
or U4931 (N_4931,N_2154,N_548);
and U4932 (N_4932,N_292,N_2939);
xnor U4933 (N_4933,N_1013,N_2782);
xnor U4934 (N_4934,N_373,N_438);
and U4935 (N_4935,N_1471,N_2233);
or U4936 (N_4936,N_778,N_2270);
nand U4937 (N_4937,N_2249,N_185);
nor U4938 (N_4938,N_551,N_2930);
or U4939 (N_4939,N_1947,N_435);
or U4940 (N_4940,N_950,N_2567);
nand U4941 (N_4941,N_138,N_10);
nor U4942 (N_4942,N_368,N_21);
nor U4943 (N_4943,N_1283,N_1032);
nand U4944 (N_4944,N_960,N_2493);
and U4945 (N_4945,N_1499,N_821);
nand U4946 (N_4946,N_1455,N_582);
nor U4947 (N_4947,N_1940,N_3108);
nor U4948 (N_4948,N_1442,N_2732);
nand U4949 (N_4949,N_666,N_2076);
nor U4950 (N_4950,N_413,N_1831);
and U4951 (N_4951,N_565,N_1807);
and U4952 (N_4952,N_2513,N_463);
and U4953 (N_4953,N_1747,N_1821);
nand U4954 (N_4954,N_585,N_2421);
nor U4955 (N_4955,N_446,N_1755);
nand U4956 (N_4956,N_153,N_1681);
or U4957 (N_4957,N_791,N_2760);
or U4958 (N_4958,N_691,N_2269);
nand U4959 (N_4959,N_2160,N_2678);
xor U4960 (N_4960,N_1569,N_542);
or U4961 (N_4961,N_184,N_2117);
or U4962 (N_4962,N_3107,N_444);
nor U4963 (N_4963,N_1181,N_764);
nand U4964 (N_4964,N_2144,N_2364);
nand U4965 (N_4965,N_625,N_2367);
nand U4966 (N_4966,N_663,N_1153);
or U4967 (N_4967,N_1742,N_2677);
nor U4968 (N_4968,N_2472,N_2230);
nand U4969 (N_4969,N_2351,N_2511);
nor U4970 (N_4970,N_1854,N_2826);
and U4971 (N_4971,N_2271,N_2808);
nand U4972 (N_4972,N_3093,N_193);
nand U4973 (N_4973,N_1649,N_588);
and U4974 (N_4974,N_262,N_1232);
and U4975 (N_4975,N_272,N_2566);
or U4976 (N_4976,N_2636,N_2390);
or U4977 (N_4977,N_676,N_1650);
and U4978 (N_4978,N_2462,N_2146);
or U4979 (N_4979,N_956,N_2805);
nand U4980 (N_4980,N_776,N_203);
nand U4981 (N_4981,N_1119,N_2822);
nand U4982 (N_4982,N_2969,N_930);
xor U4983 (N_4983,N_2968,N_1110);
nor U4984 (N_4984,N_1910,N_2531);
nand U4985 (N_4985,N_2343,N_296);
xnor U4986 (N_4986,N_418,N_774);
or U4987 (N_4987,N_2642,N_1844);
and U4988 (N_4988,N_2381,N_424);
and U4989 (N_4989,N_1228,N_2223);
xnor U4990 (N_4990,N_2003,N_1727);
nor U4991 (N_4991,N_2634,N_734);
or U4992 (N_4992,N_2261,N_2561);
and U4993 (N_4993,N_1674,N_3040);
and U4994 (N_4994,N_1021,N_768);
and U4995 (N_4995,N_1382,N_2580);
nor U4996 (N_4996,N_2491,N_1272);
xor U4997 (N_4997,N_3021,N_2233);
nor U4998 (N_4998,N_3102,N_2588);
or U4999 (N_4999,N_691,N_1487);
xnor U5000 (N_5000,N_1550,N_2951);
xnor U5001 (N_5001,N_3042,N_2833);
and U5002 (N_5002,N_356,N_57);
or U5003 (N_5003,N_2663,N_2384);
nand U5004 (N_5004,N_2382,N_2715);
nor U5005 (N_5005,N_2901,N_1130);
nand U5006 (N_5006,N_1017,N_1137);
or U5007 (N_5007,N_838,N_2194);
xor U5008 (N_5008,N_1326,N_2206);
or U5009 (N_5009,N_1418,N_933);
nor U5010 (N_5010,N_643,N_700);
and U5011 (N_5011,N_415,N_2825);
nand U5012 (N_5012,N_2019,N_797);
or U5013 (N_5013,N_1900,N_769);
or U5014 (N_5014,N_2055,N_2935);
nor U5015 (N_5015,N_2919,N_681);
or U5016 (N_5016,N_2983,N_189);
xor U5017 (N_5017,N_318,N_2101);
or U5018 (N_5018,N_2950,N_490);
or U5019 (N_5019,N_1674,N_512);
and U5020 (N_5020,N_1297,N_1452);
nand U5021 (N_5021,N_540,N_1903);
nand U5022 (N_5022,N_609,N_2053);
or U5023 (N_5023,N_958,N_3069);
nand U5024 (N_5024,N_1155,N_1121);
nor U5025 (N_5025,N_1686,N_277);
nand U5026 (N_5026,N_1630,N_1221);
nor U5027 (N_5027,N_2443,N_2606);
and U5028 (N_5028,N_848,N_1070);
and U5029 (N_5029,N_1217,N_2363);
and U5030 (N_5030,N_2569,N_139);
and U5031 (N_5031,N_2151,N_301);
nor U5032 (N_5032,N_22,N_1750);
and U5033 (N_5033,N_61,N_1569);
nand U5034 (N_5034,N_2151,N_3008);
nand U5035 (N_5035,N_1025,N_342);
nand U5036 (N_5036,N_947,N_1776);
and U5037 (N_5037,N_2251,N_2843);
nor U5038 (N_5038,N_1353,N_2241);
xor U5039 (N_5039,N_412,N_721);
nor U5040 (N_5040,N_2163,N_1172);
and U5041 (N_5041,N_3122,N_567);
or U5042 (N_5042,N_184,N_1924);
and U5043 (N_5043,N_1546,N_559);
nor U5044 (N_5044,N_1301,N_3040);
or U5045 (N_5045,N_1514,N_874);
nand U5046 (N_5046,N_2922,N_1447);
and U5047 (N_5047,N_808,N_170);
nor U5048 (N_5048,N_1525,N_987);
nor U5049 (N_5049,N_1519,N_1129);
nand U5050 (N_5050,N_495,N_1792);
nor U5051 (N_5051,N_2250,N_618);
and U5052 (N_5052,N_2492,N_1939);
nand U5053 (N_5053,N_1777,N_2411);
nand U5054 (N_5054,N_1657,N_1678);
and U5055 (N_5055,N_1073,N_213);
nor U5056 (N_5056,N_1261,N_2790);
nor U5057 (N_5057,N_503,N_1725);
or U5058 (N_5058,N_899,N_1640);
nand U5059 (N_5059,N_1375,N_2943);
or U5060 (N_5060,N_2822,N_114);
and U5061 (N_5061,N_782,N_318);
xor U5062 (N_5062,N_2125,N_2863);
and U5063 (N_5063,N_1777,N_2011);
nor U5064 (N_5064,N_520,N_1411);
and U5065 (N_5065,N_1139,N_2259);
nor U5066 (N_5066,N_3004,N_1269);
nand U5067 (N_5067,N_508,N_847);
nand U5068 (N_5068,N_748,N_2848);
and U5069 (N_5069,N_1654,N_1642);
and U5070 (N_5070,N_1147,N_2785);
nor U5071 (N_5071,N_850,N_1210);
and U5072 (N_5072,N_1352,N_2247);
nor U5073 (N_5073,N_1876,N_1364);
nor U5074 (N_5074,N_1881,N_1113);
and U5075 (N_5075,N_2228,N_862);
or U5076 (N_5076,N_589,N_821);
xor U5077 (N_5077,N_1998,N_1344);
and U5078 (N_5078,N_2460,N_1484);
or U5079 (N_5079,N_2875,N_1217);
or U5080 (N_5080,N_2911,N_263);
and U5081 (N_5081,N_2666,N_497);
and U5082 (N_5082,N_1279,N_1530);
nand U5083 (N_5083,N_60,N_304);
and U5084 (N_5084,N_1811,N_757);
and U5085 (N_5085,N_790,N_113);
or U5086 (N_5086,N_2618,N_1640);
nor U5087 (N_5087,N_151,N_1639);
nand U5088 (N_5088,N_467,N_1878);
and U5089 (N_5089,N_354,N_2274);
nand U5090 (N_5090,N_1011,N_2506);
and U5091 (N_5091,N_949,N_2052);
and U5092 (N_5092,N_421,N_2200);
and U5093 (N_5093,N_694,N_798);
nor U5094 (N_5094,N_816,N_1471);
and U5095 (N_5095,N_777,N_1035);
nand U5096 (N_5096,N_821,N_968);
nor U5097 (N_5097,N_102,N_2492);
or U5098 (N_5098,N_1903,N_1471);
nand U5099 (N_5099,N_167,N_587);
xor U5100 (N_5100,N_1443,N_637);
xnor U5101 (N_5101,N_2536,N_741);
and U5102 (N_5102,N_472,N_1852);
nor U5103 (N_5103,N_1035,N_2172);
nand U5104 (N_5104,N_2496,N_3103);
nand U5105 (N_5105,N_869,N_1418);
and U5106 (N_5106,N_2726,N_2921);
nor U5107 (N_5107,N_2169,N_2625);
or U5108 (N_5108,N_422,N_2606);
nand U5109 (N_5109,N_777,N_2762);
nor U5110 (N_5110,N_1676,N_968);
or U5111 (N_5111,N_2869,N_2406);
or U5112 (N_5112,N_1112,N_1704);
and U5113 (N_5113,N_7,N_220);
nor U5114 (N_5114,N_2372,N_960);
and U5115 (N_5115,N_2726,N_269);
xor U5116 (N_5116,N_2573,N_3105);
and U5117 (N_5117,N_1782,N_2808);
nand U5118 (N_5118,N_1874,N_103);
or U5119 (N_5119,N_1631,N_2966);
nor U5120 (N_5120,N_1367,N_299);
nor U5121 (N_5121,N_1251,N_2114);
and U5122 (N_5122,N_1909,N_1272);
nor U5123 (N_5123,N_1704,N_1665);
or U5124 (N_5124,N_1666,N_2358);
or U5125 (N_5125,N_87,N_1216);
or U5126 (N_5126,N_2549,N_676);
nor U5127 (N_5127,N_1343,N_1291);
or U5128 (N_5128,N_1671,N_1457);
and U5129 (N_5129,N_2670,N_1901);
nor U5130 (N_5130,N_538,N_1620);
nor U5131 (N_5131,N_2326,N_1766);
xor U5132 (N_5132,N_379,N_1311);
xnor U5133 (N_5133,N_2628,N_550);
nor U5134 (N_5134,N_1126,N_1495);
xnor U5135 (N_5135,N_1422,N_1162);
or U5136 (N_5136,N_2194,N_862);
nand U5137 (N_5137,N_490,N_3053);
nand U5138 (N_5138,N_2384,N_99);
and U5139 (N_5139,N_2318,N_1179);
or U5140 (N_5140,N_473,N_2875);
nand U5141 (N_5141,N_2118,N_477);
nor U5142 (N_5142,N_2022,N_99);
nand U5143 (N_5143,N_1474,N_2697);
and U5144 (N_5144,N_197,N_2007);
or U5145 (N_5145,N_3098,N_2528);
nor U5146 (N_5146,N_2028,N_1972);
nand U5147 (N_5147,N_988,N_2591);
xnor U5148 (N_5148,N_162,N_977);
nand U5149 (N_5149,N_560,N_2002);
nand U5150 (N_5150,N_1102,N_1700);
nand U5151 (N_5151,N_793,N_3035);
or U5152 (N_5152,N_2224,N_1113);
or U5153 (N_5153,N_2086,N_1987);
nand U5154 (N_5154,N_1382,N_1446);
and U5155 (N_5155,N_1575,N_631);
or U5156 (N_5156,N_2798,N_1215);
xnor U5157 (N_5157,N_2200,N_797);
and U5158 (N_5158,N_2249,N_267);
or U5159 (N_5159,N_2682,N_2594);
and U5160 (N_5160,N_2547,N_2685);
and U5161 (N_5161,N_513,N_589);
and U5162 (N_5162,N_1835,N_712);
nand U5163 (N_5163,N_2888,N_1503);
and U5164 (N_5164,N_1099,N_2907);
nand U5165 (N_5165,N_1715,N_1925);
nand U5166 (N_5166,N_53,N_2833);
and U5167 (N_5167,N_248,N_1275);
and U5168 (N_5168,N_2935,N_2193);
xnor U5169 (N_5169,N_1068,N_2902);
and U5170 (N_5170,N_1436,N_797);
nor U5171 (N_5171,N_3037,N_315);
or U5172 (N_5172,N_2797,N_1920);
or U5173 (N_5173,N_1225,N_2961);
or U5174 (N_5174,N_97,N_632);
and U5175 (N_5175,N_2001,N_3000);
nand U5176 (N_5176,N_2375,N_942);
nor U5177 (N_5177,N_1940,N_2739);
nor U5178 (N_5178,N_2534,N_1291);
nor U5179 (N_5179,N_1629,N_236);
nand U5180 (N_5180,N_2558,N_386);
and U5181 (N_5181,N_690,N_222);
nor U5182 (N_5182,N_79,N_1482);
nand U5183 (N_5183,N_958,N_1008);
or U5184 (N_5184,N_952,N_2079);
and U5185 (N_5185,N_2699,N_1389);
nand U5186 (N_5186,N_1947,N_2918);
or U5187 (N_5187,N_2253,N_2602);
nor U5188 (N_5188,N_311,N_1593);
and U5189 (N_5189,N_1754,N_2802);
or U5190 (N_5190,N_428,N_1166);
nand U5191 (N_5191,N_3028,N_2874);
nand U5192 (N_5192,N_1772,N_2821);
nor U5193 (N_5193,N_2635,N_803);
nor U5194 (N_5194,N_550,N_1592);
nand U5195 (N_5195,N_2569,N_209);
or U5196 (N_5196,N_167,N_2317);
and U5197 (N_5197,N_1736,N_409);
and U5198 (N_5198,N_2290,N_1536);
nor U5199 (N_5199,N_1279,N_985);
nor U5200 (N_5200,N_553,N_1620);
and U5201 (N_5201,N_2682,N_477);
nor U5202 (N_5202,N_2095,N_2730);
nand U5203 (N_5203,N_386,N_2971);
nor U5204 (N_5204,N_1606,N_1829);
nor U5205 (N_5205,N_1314,N_1241);
and U5206 (N_5206,N_1385,N_2153);
or U5207 (N_5207,N_1164,N_2676);
nor U5208 (N_5208,N_234,N_1801);
or U5209 (N_5209,N_2819,N_970);
nor U5210 (N_5210,N_2954,N_657);
or U5211 (N_5211,N_2899,N_1192);
xor U5212 (N_5212,N_1360,N_3118);
and U5213 (N_5213,N_134,N_2731);
and U5214 (N_5214,N_2966,N_718);
nand U5215 (N_5215,N_291,N_868);
and U5216 (N_5216,N_2915,N_676);
nor U5217 (N_5217,N_1788,N_913);
nor U5218 (N_5218,N_2481,N_2542);
and U5219 (N_5219,N_3015,N_2384);
and U5220 (N_5220,N_1224,N_60);
nand U5221 (N_5221,N_2216,N_1964);
and U5222 (N_5222,N_741,N_2641);
and U5223 (N_5223,N_408,N_277);
nor U5224 (N_5224,N_236,N_1640);
nor U5225 (N_5225,N_1544,N_1077);
nor U5226 (N_5226,N_89,N_2265);
and U5227 (N_5227,N_2133,N_1504);
nand U5228 (N_5228,N_3002,N_1560);
or U5229 (N_5229,N_2833,N_1089);
and U5230 (N_5230,N_1467,N_2872);
and U5231 (N_5231,N_788,N_680);
xnor U5232 (N_5232,N_1943,N_2667);
nor U5233 (N_5233,N_60,N_839);
and U5234 (N_5234,N_1927,N_1531);
nor U5235 (N_5235,N_2252,N_2496);
or U5236 (N_5236,N_1611,N_1773);
and U5237 (N_5237,N_2272,N_1198);
and U5238 (N_5238,N_1474,N_2583);
nand U5239 (N_5239,N_2227,N_2185);
and U5240 (N_5240,N_2901,N_416);
or U5241 (N_5241,N_1811,N_732);
nor U5242 (N_5242,N_464,N_1680);
nand U5243 (N_5243,N_3086,N_1759);
xnor U5244 (N_5244,N_2515,N_2262);
and U5245 (N_5245,N_2948,N_595);
nor U5246 (N_5246,N_334,N_1335);
xor U5247 (N_5247,N_2701,N_1393);
and U5248 (N_5248,N_1858,N_937);
or U5249 (N_5249,N_1546,N_3057);
xor U5250 (N_5250,N_3068,N_2068);
nor U5251 (N_5251,N_1761,N_1168);
or U5252 (N_5252,N_1646,N_1921);
nor U5253 (N_5253,N_354,N_857);
or U5254 (N_5254,N_1427,N_2997);
or U5255 (N_5255,N_1375,N_2479);
or U5256 (N_5256,N_1707,N_1652);
nor U5257 (N_5257,N_348,N_1683);
and U5258 (N_5258,N_2151,N_1515);
nand U5259 (N_5259,N_546,N_753);
or U5260 (N_5260,N_2239,N_633);
xnor U5261 (N_5261,N_1920,N_819);
nand U5262 (N_5262,N_2227,N_2297);
and U5263 (N_5263,N_2329,N_1779);
or U5264 (N_5264,N_1394,N_1);
or U5265 (N_5265,N_1672,N_404);
or U5266 (N_5266,N_2816,N_1829);
or U5267 (N_5267,N_1150,N_372);
or U5268 (N_5268,N_1880,N_966);
or U5269 (N_5269,N_2801,N_2354);
nand U5270 (N_5270,N_2691,N_1504);
and U5271 (N_5271,N_2392,N_505);
and U5272 (N_5272,N_2513,N_320);
nor U5273 (N_5273,N_2598,N_828);
nor U5274 (N_5274,N_482,N_696);
nand U5275 (N_5275,N_1204,N_1777);
and U5276 (N_5276,N_1969,N_2892);
and U5277 (N_5277,N_1367,N_2469);
or U5278 (N_5278,N_2905,N_1728);
xnor U5279 (N_5279,N_1459,N_1777);
nor U5280 (N_5280,N_1647,N_2860);
nand U5281 (N_5281,N_488,N_675);
nand U5282 (N_5282,N_2344,N_1593);
nand U5283 (N_5283,N_1288,N_1864);
xnor U5284 (N_5284,N_1456,N_746);
or U5285 (N_5285,N_1653,N_1981);
nor U5286 (N_5286,N_155,N_1216);
nand U5287 (N_5287,N_974,N_1548);
and U5288 (N_5288,N_3068,N_2278);
and U5289 (N_5289,N_878,N_1149);
nand U5290 (N_5290,N_623,N_296);
xor U5291 (N_5291,N_1494,N_1145);
or U5292 (N_5292,N_2118,N_327);
and U5293 (N_5293,N_117,N_1978);
or U5294 (N_5294,N_3061,N_1297);
and U5295 (N_5295,N_2633,N_2661);
or U5296 (N_5296,N_961,N_1560);
nor U5297 (N_5297,N_1580,N_1193);
xor U5298 (N_5298,N_1538,N_1457);
nor U5299 (N_5299,N_1365,N_563);
nand U5300 (N_5300,N_2877,N_2963);
nand U5301 (N_5301,N_1780,N_32);
nand U5302 (N_5302,N_2929,N_2609);
nand U5303 (N_5303,N_1342,N_3051);
and U5304 (N_5304,N_1414,N_715);
and U5305 (N_5305,N_828,N_2515);
and U5306 (N_5306,N_2814,N_2811);
and U5307 (N_5307,N_2776,N_23);
and U5308 (N_5308,N_2377,N_1510);
or U5309 (N_5309,N_688,N_1303);
nand U5310 (N_5310,N_438,N_2717);
nor U5311 (N_5311,N_2463,N_1685);
or U5312 (N_5312,N_126,N_693);
nand U5313 (N_5313,N_2749,N_2524);
and U5314 (N_5314,N_269,N_2196);
and U5315 (N_5315,N_2375,N_3049);
and U5316 (N_5316,N_724,N_1609);
nor U5317 (N_5317,N_1045,N_2076);
xnor U5318 (N_5318,N_2936,N_1663);
nand U5319 (N_5319,N_838,N_2805);
or U5320 (N_5320,N_2398,N_1862);
nand U5321 (N_5321,N_2558,N_2003);
or U5322 (N_5322,N_420,N_2511);
xnor U5323 (N_5323,N_2664,N_2060);
and U5324 (N_5324,N_1276,N_1648);
nand U5325 (N_5325,N_1655,N_1526);
nand U5326 (N_5326,N_2231,N_1120);
nand U5327 (N_5327,N_382,N_2869);
or U5328 (N_5328,N_1353,N_270);
nand U5329 (N_5329,N_883,N_1858);
xor U5330 (N_5330,N_2372,N_784);
nand U5331 (N_5331,N_197,N_668);
nand U5332 (N_5332,N_917,N_2141);
nand U5333 (N_5333,N_1202,N_1264);
nor U5334 (N_5334,N_1718,N_146);
nand U5335 (N_5335,N_699,N_3036);
xnor U5336 (N_5336,N_426,N_13);
nor U5337 (N_5337,N_1382,N_1154);
and U5338 (N_5338,N_2899,N_2671);
nand U5339 (N_5339,N_659,N_235);
nand U5340 (N_5340,N_2759,N_2013);
or U5341 (N_5341,N_1584,N_3110);
and U5342 (N_5342,N_2285,N_2707);
nand U5343 (N_5343,N_161,N_2661);
and U5344 (N_5344,N_2566,N_196);
or U5345 (N_5345,N_2100,N_1083);
or U5346 (N_5346,N_1902,N_581);
or U5347 (N_5347,N_439,N_3027);
or U5348 (N_5348,N_2168,N_2102);
xor U5349 (N_5349,N_713,N_102);
xnor U5350 (N_5350,N_2293,N_2542);
or U5351 (N_5351,N_717,N_2614);
or U5352 (N_5352,N_2613,N_2312);
nor U5353 (N_5353,N_2996,N_2931);
nor U5354 (N_5354,N_2964,N_1117);
and U5355 (N_5355,N_57,N_1933);
or U5356 (N_5356,N_2236,N_917);
or U5357 (N_5357,N_2125,N_2261);
and U5358 (N_5358,N_1455,N_1977);
and U5359 (N_5359,N_187,N_2817);
nand U5360 (N_5360,N_3078,N_367);
nand U5361 (N_5361,N_49,N_1296);
or U5362 (N_5362,N_2937,N_2378);
or U5363 (N_5363,N_745,N_1103);
xnor U5364 (N_5364,N_2727,N_2437);
nand U5365 (N_5365,N_556,N_851);
and U5366 (N_5366,N_478,N_1693);
xnor U5367 (N_5367,N_181,N_2278);
nand U5368 (N_5368,N_2331,N_2317);
nand U5369 (N_5369,N_2235,N_2303);
xnor U5370 (N_5370,N_644,N_1211);
nand U5371 (N_5371,N_1147,N_3028);
nand U5372 (N_5372,N_2843,N_240);
or U5373 (N_5373,N_2764,N_692);
nor U5374 (N_5374,N_857,N_1543);
and U5375 (N_5375,N_2161,N_1034);
nand U5376 (N_5376,N_2102,N_1007);
nor U5377 (N_5377,N_1144,N_760);
or U5378 (N_5378,N_2382,N_625);
nor U5379 (N_5379,N_490,N_2318);
and U5380 (N_5380,N_1804,N_2494);
or U5381 (N_5381,N_391,N_2892);
or U5382 (N_5382,N_2257,N_1630);
nor U5383 (N_5383,N_2962,N_1253);
or U5384 (N_5384,N_1001,N_2254);
or U5385 (N_5385,N_106,N_294);
and U5386 (N_5386,N_734,N_988);
nor U5387 (N_5387,N_2914,N_240);
nor U5388 (N_5388,N_2193,N_465);
nor U5389 (N_5389,N_2968,N_1269);
nand U5390 (N_5390,N_3052,N_1998);
or U5391 (N_5391,N_2854,N_2635);
nor U5392 (N_5392,N_2921,N_1031);
nor U5393 (N_5393,N_2967,N_817);
nor U5394 (N_5394,N_1762,N_2139);
and U5395 (N_5395,N_738,N_720);
nand U5396 (N_5396,N_1665,N_2258);
nor U5397 (N_5397,N_2701,N_763);
nor U5398 (N_5398,N_2449,N_1418);
and U5399 (N_5399,N_626,N_1062);
and U5400 (N_5400,N_1169,N_2528);
and U5401 (N_5401,N_687,N_2772);
nand U5402 (N_5402,N_2551,N_694);
or U5403 (N_5403,N_1393,N_1644);
nand U5404 (N_5404,N_1601,N_49);
nand U5405 (N_5405,N_1337,N_2041);
and U5406 (N_5406,N_1763,N_2280);
and U5407 (N_5407,N_508,N_2342);
xnor U5408 (N_5408,N_97,N_2977);
xnor U5409 (N_5409,N_1816,N_1961);
nand U5410 (N_5410,N_2320,N_1893);
xnor U5411 (N_5411,N_2747,N_228);
and U5412 (N_5412,N_2664,N_2399);
and U5413 (N_5413,N_521,N_2178);
nand U5414 (N_5414,N_1424,N_2301);
and U5415 (N_5415,N_478,N_1362);
or U5416 (N_5416,N_2847,N_1424);
and U5417 (N_5417,N_1000,N_2707);
nor U5418 (N_5418,N_1109,N_2908);
and U5419 (N_5419,N_703,N_123);
xnor U5420 (N_5420,N_152,N_2060);
nand U5421 (N_5421,N_42,N_2291);
nand U5422 (N_5422,N_3086,N_589);
nor U5423 (N_5423,N_2901,N_3024);
nand U5424 (N_5424,N_892,N_1975);
nor U5425 (N_5425,N_410,N_343);
nor U5426 (N_5426,N_2975,N_245);
xor U5427 (N_5427,N_2078,N_1891);
or U5428 (N_5428,N_3027,N_1210);
nand U5429 (N_5429,N_195,N_2124);
and U5430 (N_5430,N_794,N_326);
nor U5431 (N_5431,N_1923,N_2847);
nor U5432 (N_5432,N_1191,N_1070);
xor U5433 (N_5433,N_2682,N_958);
nor U5434 (N_5434,N_1112,N_2158);
xnor U5435 (N_5435,N_1024,N_1908);
nor U5436 (N_5436,N_2200,N_2497);
nor U5437 (N_5437,N_1,N_2845);
xnor U5438 (N_5438,N_3046,N_3038);
nor U5439 (N_5439,N_1880,N_2051);
nand U5440 (N_5440,N_999,N_2663);
nor U5441 (N_5441,N_691,N_2872);
nand U5442 (N_5442,N_653,N_1525);
and U5443 (N_5443,N_2411,N_250);
or U5444 (N_5444,N_2613,N_1025);
nor U5445 (N_5445,N_646,N_2741);
nand U5446 (N_5446,N_522,N_593);
xnor U5447 (N_5447,N_1605,N_2413);
nand U5448 (N_5448,N_2753,N_180);
nand U5449 (N_5449,N_601,N_323);
nand U5450 (N_5450,N_509,N_72);
and U5451 (N_5451,N_2993,N_720);
and U5452 (N_5452,N_2925,N_1609);
or U5453 (N_5453,N_1370,N_2406);
nand U5454 (N_5454,N_1051,N_18);
xnor U5455 (N_5455,N_823,N_1016);
or U5456 (N_5456,N_995,N_1877);
or U5457 (N_5457,N_48,N_2223);
or U5458 (N_5458,N_1230,N_1562);
nor U5459 (N_5459,N_2077,N_2997);
nand U5460 (N_5460,N_1300,N_2207);
and U5461 (N_5461,N_3034,N_2747);
nor U5462 (N_5462,N_1703,N_1546);
nor U5463 (N_5463,N_536,N_1696);
and U5464 (N_5464,N_782,N_356);
and U5465 (N_5465,N_569,N_1719);
xor U5466 (N_5466,N_2,N_1493);
nand U5467 (N_5467,N_525,N_1056);
nor U5468 (N_5468,N_615,N_475);
nor U5469 (N_5469,N_1236,N_1245);
xnor U5470 (N_5470,N_130,N_761);
and U5471 (N_5471,N_537,N_2485);
nor U5472 (N_5472,N_2928,N_1343);
nor U5473 (N_5473,N_441,N_495);
nand U5474 (N_5474,N_689,N_1626);
nor U5475 (N_5475,N_1566,N_3120);
and U5476 (N_5476,N_2268,N_958);
nor U5477 (N_5477,N_520,N_2007);
nor U5478 (N_5478,N_2680,N_2387);
nand U5479 (N_5479,N_3023,N_1917);
nand U5480 (N_5480,N_2580,N_3031);
nor U5481 (N_5481,N_1628,N_2611);
or U5482 (N_5482,N_2022,N_2493);
nand U5483 (N_5483,N_518,N_594);
and U5484 (N_5484,N_1317,N_1736);
nand U5485 (N_5485,N_2649,N_2181);
and U5486 (N_5486,N_474,N_1617);
or U5487 (N_5487,N_354,N_2808);
nand U5488 (N_5488,N_1887,N_3064);
xnor U5489 (N_5489,N_1942,N_3046);
nand U5490 (N_5490,N_1082,N_2230);
nand U5491 (N_5491,N_2019,N_554);
nor U5492 (N_5492,N_861,N_1151);
or U5493 (N_5493,N_717,N_2186);
nand U5494 (N_5494,N_30,N_850);
nand U5495 (N_5495,N_142,N_3026);
nor U5496 (N_5496,N_2866,N_2325);
nor U5497 (N_5497,N_941,N_2331);
nor U5498 (N_5498,N_187,N_2399);
and U5499 (N_5499,N_980,N_3071);
nor U5500 (N_5500,N_2458,N_2362);
nor U5501 (N_5501,N_654,N_1804);
nor U5502 (N_5502,N_3075,N_2754);
or U5503 (N_5503,N_756,N_2187);
nor U5504 (N_5504,N_2396,N_1196);
and U5505 (N_5505,N_196,N_2890);
and U5506 (N_5506,N_813,N_199);
nor U5507 (N_5507,N_1082,N_308);
nor U5508 (N_5508,N_1550,N_823);
nand U5509 (N_5509,N_1937,N_855);
nand U5510 (N_5510,N_118,N_751);
nor U5511 (N_5511,N_194,N_753);
nand U5512 (N_5512,N_529,N_3093);
or U5513 (N_5513,N_2284,N_2066);
or U5514 (N_5514,N_371,N_2454);
xor U5515 (N_5515,N_3063,N_2005);
xnor U5516 (N_5516,N_2485,N_1002);
nand U5517 (N_5517,N_1217,N_658);
xnor U5518 (N_5518,N_53,N_2445);
nor U5519 (N_5519,N_2262,N_1536);
and U5520 (N_5520,N_1577,N_368);
nor U5521 (N_5521,N_2878,N_1110);
nor U5522 (N_5522,N_375,N_2343);
nand U5523 (N_5523,N_209,N_2979);
and U5524 (N_5524,N_3040,N_46);
xnor U5525 (N_5525,N_501,N_1857);
or U5526 (N_5526,N_3028,N_2403);
nand U5527 (N_5527,N_1405,N_1394);
nand U5528 (N_5528,N_2785,N_232);
or U5529 (N_5529,N_259,N_2213);
or U5530 (N_5530,N_821,N_2539);
nor U5531 (N_5531,N_384,N_1267);
nor U5532 (N_5532,N_136,N_940);
or U5533 (N_5533,N_2606,N_1923);
or U5534 (N_5534,N_132,N_339);
nor U5535 (N_5535,N_237,N_470);
and U5536 (N_5536,N_1235,N_842);
and U5537 (N_5537,N_288,N_957);
and U5538 (N_5538,N_2353,N_1253);
nand U5539 (N_5539,N_377,N_2294);
and U5540 (N_5540,N_2665,N_2454);
or U5541 (N_5541,N_2348,N_1640);
nand U5542 (N_5542,N_1246,N_989);
nand U5543 (N_5543,N_2411,N_1206);
nand U5544 (N_5544,N_3026,N_2077);
nand U5545 (N_5545,N_2651,N_1082);
and U5546 (N_5546,N_3045,N_3089);
nor U5547 (N_5547,N_125,N_2811);
nand U5548 (N_5548,N_643,N_1002);
and U5549 (N_5549,N_1284,N_3108);
or U5550 (N_5550,N_532,N_1332);
or U5551 (N_5551,N_1073,N_425);
and U5552 (N_5552,N_3106,N_2556);
nand U5553 (N_5553,N_508,N_2278);
nor U5554 (N_5554,N_1948,N_1427);
xor U5555 (N_5555,N_2846,N_1067);
xnor U5556 (N_5556,N_3105,N_816);
or U5557 (N_5557,N_381,N_451);
nand U5558 (N_5558,N_2249,N_2267);
nor U5559 (N_5559,N_1986,N_2164);
or U5560 (N_5560,N_1388,N_1916);
nand U5561 (N_5561,N_1023,N_1693);
nand U5562 (N_5562,N_2627,N_285);
or U5563 (N_5563,N_196,N_1722);
and U5564 (N_5564,N_944,N_1055);
nor U5565 (N_5565,N_660,N_2015);
or U5566 (N_5566,N_2588,N_1166);
and U5567 (N_5567,N_1332,N_349);
nor U5568 (N_5568,N_1543,N_105);
nand U5569 (N_5569,N_648,N_975);
nand U5570 (N_5570,N_2960,N_1451);
nor U5571 (N_5571,N_258,N_2808);
nand U5572 (N_5572,N_2867,N_2);
nand U5573 (N_5573,N_327,N_2985);
nor U5574 (N_5574,N_362,N_1111);
and U5575 (N_5575,N_1270,N_2957);
nand U5576 (N_5576,N_1469,N_2668);
nor U5577 (N_5577,N_2033,N_1167);
or U5578 (N_5578,N_839,N_2501);
and U5579 (N_5579,N_3094,N_1744);
nand U5580 (N_5580,N_1012,N_145);
nand U5581 (N_5581,N_1066,N_3085);
nand U5582 (N_5582,N_2131,N_2767);
and U5583 (N_5583,N_2274,N_948);
or U5584 (N_5584,N_1338,N_662);
nand U5585 (N_5585,N_2530,N_2984);
nor U5586 (N_5586,N_1904,N_871);
nor U5587 (N_5587,N_1704,N_2319);
and U5588 (N_5588,N_1807,N_1301);
nand U5589 (N_5589,N_1274,N_835);
or U5590 (N_5590,N_112,N_2663);
nand U5591 (N_5591,N_1862,N_1888);
or U5592 (N_5592,N_2707,N_553);
and U5593 (N_5593,N_1889,N_1885);
nand U5594 (N_5594,N_1347,N_727);
or U5595 (N_5595,N_1449,N_1931);
and U5596 (N_5596,N_1661,N_2262);
nand U5597 (N_5597,N_1729,N_395);
xor U5598 (N_5598,N_424,N_948);
or U5599 (N_5599,N_28,N_1938);
nand U5600 (N_5600,N_2588,N_1327);
nor U5601 (N_5601,N_1176,N_205);
and U5602 (N_5602,N_701,N_2038);
and U5603 (N_5603,N_2607,N_72);
nor U5604 (N_5604,N_2739,N_2056);
or U5605 (N_5605,N_2731,N_750);
and U5606 (N_5606,N_409,N_780);
nor U5607 (N_5607,N_2935,N_2238);
nor U5608 (N_5608,N_2520,N_977);
and U5609 (N_5609,N_925,N_441);
nor U5610 (N_5610,N_321,N_793);
and U5611 (N_5611,N_2296,N_3083);
nor U5612 (N_5612,N_2489,N_287);
nand U5613 (N_5613,N_374,N_58);
or U5614 (N_5614,N_2356,N_2657);
or U5615 (N_5615,N_11,N_1373);
or U5616 (N_5616,N_2911,N_2357);
and U5617 (N_5617,N_2055,N_1226);
or U5618 (N_5618,N_2855,N_3059);
or U5619 (N_5619,N_1832,N_1924);
nor U5620 (N_5620,N_759,N_2259);
nand U5621 (N_5621,N_1200,N_63);
and U5622 (N_5622,N_1004,N_2961);
and U5623 (N_5623,N_20,N_360);
xnor U5624 (N_5624,N_1675,N_1868);
and U5625 (N_5625,N_2297,N_1792);
and U5626 (N_5626,N_902,N_2502);
nand U5627 (N_5627,N_1133,N_999);
nand U5628 (N_5628,N_1124,N_1763);
xnor U5629 (N_5629,N_303,N_843);
or U5630 (N_5630,N_955,N_478);
and U5631 (N_5631,N_1875,N_1608);
or U5632 (N_5632,N_365,N_1726);
or U5633 (N_5633,N_2021,N_2440);
and U5634 (N_5634,N_2767,N_878);
or U5635 (N_5635,N_2985,N_660);
nor U5636 (N_5636,N_204,N_574);
nand U5637 (N_5637,N_1003,N_286);
xor U5638 (N_5638,N_938,N_587);
xor U5639 (N_5639,N_2548,N_357);
nand U5640 (N_5640,N_1436,N_28);
or U5641 (N_5641,N_1067,N_2438);
or U5642 (N_5642,N_1432,N_1870);
nor U5643 (N_5643,N_2648,N_135);
nor U5644 (N_5644,N_663,N_1539);
and U5645 (N_5645,N_1511,N_44);
nor U5646 (N_5646,N_979,N_1974);
xor U5647 (N_5647,N_534,N_1800);
nor U5648 (N_5648,N_1159,N_2756);
or U5649 (N_5649,N_1365,N_1161);
nand U5650 (N_5650,N_295,N_748);
and U5651 (N_5651,N_1196,N_2821);
nand U5652 (N_5652,N_1225,N_525);
and U5653 (N_5653,N_2690,N_1560);
nor U5654 (N_5654,N_2331,N_1340);
and U5655 (N_5655,N_884,N_1097);
and U5656 (N_5656,N_1943,N_1241);
xnor U5657 (N_5657,N_1340,N_1770);
and U5658 (N_5658,N_1668,N_1706);
nand U5659 (N_5659,N_504,N_70);
nor U5660 (N_5660,N_1385,N_2075);
or U5661 (N_5661,N_705,N_768);
nor U5662 (N_5662,N_2013,N_908);
nand U5663 (N_5663,N_3045,N_1247);
xnor U5664 (N_5664,N_2405,N_3015);
or U5665 (N_5665,N_993,N_451);
nor U5666 (N_5666,N_1929,N_2081);
nand U5667 (N_5667,N_1827,N_3027);
and U5668 (N_5668,N_2945,N_2192);
nor U5669 (N_5669,N_2057,N_2785);
or U5670 (N_5670,N_1890,N_1682);
or U5671 (N_5671,N_910,N_2163);
or U5672 (N_5672,N_2009,N_2344);
nand U5673 (N_5673,N_1440,N_540);
and U5674 (N_5674,N_445,N_1168);
and U5675 (N_5675,N_602,N_3091);
nor U5676 (N_5676,N_2617,N_1478);
and U5677 (N_5677,N_362,N_2265);
nand U5678 (N_5678,N_2787,N_1147);
or U5679 (N_5679,N_919,N_1538);
or U5680 (N_5680,N_1859,N_838);
and U5681 (N_5681,N_2287,N_1243);
nor U5682 (N_5682,N_2983,N_309);
or U5683 (N_5683,N_2146,N_3094);
or U5684 (N_5684,N_1580,N_1353);
xnor U5685 (N_5685,N_1119,N_345);
or U5686 (N_5686,N_390,N_352);
or U5687 (N_5687,N_3030,N_1885);
nand U5688 (N_5688,N_2315,N_1240);
and U5689 (N_5689,N_544,N_1211);
nand U5690 (N_5690,N_2995,N_1222);
nand U5691 (N_5691,N_1519,N_2508);
xnor U5692 (N_5692,N_875,N_837);
nand U5693 (N_5693,N_2944,N_1631);
nor U5694 (N_5694,N_1162,N_383);
or U5695 (N_5695,N_2726,N_914);
nand U5696 (N_5696,N_2114,N_2731);
nor U5697 (N_5697,N_286,N_174);
or U5698 (N_5698,N_1660,N_1459);
nor U5699 (N_5699,N_467,N_2446);
and U5700 (N_5700,N_1138,N_862);
or U5701 (N_5701,N_2991,N_252);
or U5702 (N_5702,N_3055,N_1802);
and U5703 (N_5703,N_2346,N_2092);
nor U5704 (N_5704,N_2011,N_2064);
or U5705 (N_5705,N_1930,N_1423);
nand U5706 (N_5706,N_2930,N_2797);
or U5707 (N_5707,N_251,N_2188);
or U5708 (N_5708,N_1161,N_164);
nand U5709 (N_5709,N_2457,N_212);
xnor U5710 (N_5710,N_2346,N_1305);
xnor U5711 (N_5711,N_1199,N_1655);
nand U5712 (N_5712,N_1771,N_2493);
or U5713 (N_5713,N_988,N_551);
and U5714 (N_5714,N_156,N_2258);
nor U5715 (N_5715,N_2038,N_737);
nand U5716 (N_5716,N_2340,N_2944);
nand U5717 (N_5717,N_1837,N_457);
and U5718 (N_5718,N_2364,N_1483);
nand U5719 (N_5719,N_2552,N_2439);
and U5720 (N_5720,N_1668,N_2917);
nor U5721 (N_5721,N_1559,N_2813);
and U5722 (N_5722,N_464,N_837);
and U5723 (N_5723,N_108,N_927);
or U5724 (N_5724,N_681,N_2248);
nand U5725 (N_5725,N_541,N_2930);
and U5726 (N_5726,N_15,N_1854);
or U5727 (N_5727,N_3075,N_277);
and U5728 (N_5728,N_3073,N_1809);
nor U5729 (N_5729,N_569,N_2388);
xor U5730 (N_5730,N_2798,N_1629);
nand U5731 (N_5731,N_929,N_845);
nor U5732 (N_5732,N_2857,N_433);
or U5733 (N_5733,N_2320,N_541);
and U5734 (N_5734,N_1086,N_2201);
nand U5735 (N_5735,N_1324,N_383);
and U5736 (N_5736,N_2960,N_2517);
nor U5737 (N_5737,N_2950,N_2148);
nor U5738 (N_5738,N_2317,N_1558);
and U5739 (N_5739,N_2196,N_2331);
xor U5740 (N_5740,N_2009,N_1864);
nand U5741 (N_5741,N_1371,N_1731);
or U5742 (N_5742,N_800,N_980);
and U5743 (N_5743,N_2187,N_1310);
nand U5744 (N_5744,N_2156,N_76);
nand U5745 (N_5745,N_778,N_409);
and U5746 (N_5746,N_2588,N_2728);
nor U5747 (N_5747,N_2783,N_805);
or U5748 (N_5748,N_1736,N_2248);
and U5749 (N_5749,N_1984,N_2803);
xor U5750 (N_5750,N_1529,N_1241);
nand U5751 (N_5751,N_682,N_1793);
or U5752 (N_5752,N_1281,N_545);
nor U5753 (N_5753,N_2468,N_651);
or U5754 (N_5754,N_20,N_588);
and U5755 (N_5755,N_2616,N_3078);
nand U5756 (N_5756,N_1507,N_1514);
nand U5757 (N_5757,N_2837,N_847);
nor U5758 (N_5758,N_812,N_1839);
nor U5759 (N_5759,N_694,N_967);
nor U5760 (N_5760,N_1787,N_1619);
nor U5761 (N_5761,N_1574,N_568);
xnor U5762 (N_5762,N_2189,N_1828);
nor U5763 (N_5763,N_34,N_1070);
xor U5764 (N_5764,N_2080,N_2486);
or U5765 (N_5765,N_2913,N_2368);
nor U5766 (N_5766,N_2499,N_1918);
xor U5767 (N_5767,N_1303,N_1334);
and U5768 (N_5768,N_2284,N_2455);
and U5769 (N_5769,N_1050,N_2403);
nand U5770 (N_5770,N_933,N_1472);
or U5771 (N_5771,N_258,N_2795);
nor U5772 (N_5772,N_2677,N_2710);
nand U5773 (N_5773,N_2591,N_253);
and U5774 (N_5774,N_2964,N_2942);
or U5775 (N_5775,N_734,N_820);
or U5776 (N_5776,N_3014,N_2768);
nand U5777 (N_5777,N_2779,N_1181);
nand U5778 (N_5778,N_1873,N_68);
xnor U5779 (N_5779,N_911,N_2050);
or U5780 (N_5780,N_1158,N_2825);
nand U5781 (N_5781,N_3095,N_1758);
nor U5782 (N_5782,N_1273,N_1664);
or U5783 (N_5783,N_2091,N_1086);
nor U5784 (N_5784,N_2446,N_2190);
and U5785 (N_5785,N_1389,N_124);
and U5786 (N_5786,N_3005,N_190);
or U5787 (N_5787,N_2634,N_2084);
nand U5788 (N_5788,N_2559,N_3124);
or U5789 (N_5789,N_1499,N_1107);
nand U5790 (N_5790,N_420,N_573);
nor U5791 (N_5791,N_1953,N_99);
nor U5792 (N_5792,N_754,N_566);
nand U5793 (N_5793,N_805,N_675);
nand U5794 (N_5794,N_1310,N_629);
and U5795 (N_5795,N_568,N_738);
and U5796 (N_5796,N_2686,N_856);
or U5797 (N_5797,N_482,N_531);
or U5798 (N_5798,N_1596,N_945);
nor U5799 (N_5799,N_449,N_2179);
or U5800 (N_5800,N_1457,N_3019);
nor U5801 (N_5801,N_1008,N_1615);
nand U5802 (N_5802,N_2936,N_1472);
nand U5803 (N_5803,N_2147,N_1500);
nor U5804 (N_5804,N_1846,N_830);
xnor U5805 (N_5805,N_1238,N_834);
nand U5806 (N_5806,N_304,N_2542);
nor U5807 (N_5807,N_551,N_744);
and U5808 (N_5808,N_1352,N_2573);
or U5809 (N_5809,N_2537,N_2080);
nor U5810 (N_5810,N_3041,N_2761);
xnor U5811 (N_5811,N_2755,N_2832);
nand U5812 (N_5812,N_2849,N_2975);
or U5813 (N_5813,N_1255,N_1813);
xor U5814 (N_5814,N_1400,N_249);
or U5815 (N_5815,N_2487,N_586);
nor U5816 (N_5816,N_1204,N_1538);
or U5817 (N_5817,N_1492,N_393);
or U5818 (N_5818,N_679,N_405);
nor U5819 (N_5819,N_723,N_856);
and U5820 (N_5820,N_1333,N_2976);
xor U5821 (N_5821,N_2023,N_2978);
and U5822 (N_5822,N_1664,N_305);
and U5823 (N_5823,N_427,N_757);
nor U5824 (N_5824,N_2978,N_855);
or U5825 (N_5825,N_752,N_3061);
nand U5826 (N_5826,N_2639,N_1079);
and U5827 (N_5827,N_2247,N_3066);
or U5828 (N_5828,N_2329,N_2725);
and U5829 (N_5829,N_3041,N_1922);
or U5830 (N_5830,N_2958,N_2327);
nor U5831 (N_5831,N_3071,N_1502);
and U5832 (N_5832,N_2729,N_2661);
and U5833 (N_5833,N_512,N_1444);
nor U5834 (N_5834,N_2364,N_1252);
and U5835 (N_5835,N_357,N_2576);
or U5836 (N_5836,N_517,N_2980);
xnor U5837 (N_5837,N_1448,N_1168);
nor U5838 (N_5838,N_1059,N_1924);
and U5839 (N_5839,N_2959,N_699);
nor U5840 (N_5840,N_1837,N_295);
nor U5841 (N_5841,N_1562,N_2152);
nor U5842 (N_5842,N_2461,N_2782);
or U5843 (N_5843,N_51,N_958);
and U5844 (N_5844,N_3036,N_2763);
nand U5845 (N_5845,N_3120,N_344);
or U5846 (N_5846,N_2123,N_1317);
nand U5847 (N_5847,N_2538,N_1849);
and U5848 (N_5848,N_2559,N_2108);
or U5849 (N_5849,N_2363,N_1591);
nand U5850 (N_5850,N_1703,N_63);
nand U5851 (N_5851,N_2550,N_648);
nand U5852 (N_5852,N_2090,N_1332);
and U5853 (N_5853,N_516,N_2676);
or U5854 (N_5854,N_1373,N_843);
nor U5855 (N_5855,N_1782,N_934);
or U5856 (N_5856,N_820,N_2516);
nand U5857 (N_5857,N_2807,N_1636);
and U5858 (N_5858,N_2604,N_1778);
nand U5859 (N_5859,N_1521,N_142);
or U5860 (N_5860,N_1779,N_2793);
nor U5861 (N_5861,N_1083,N_1743);
xor U5862 (N_5862,N_2051,N_2588);
or U5863 (N_5863,N_2745,N_2991);
or U5864 (N_5864,N_2684,N_1652);
nor U5865 (N_5865,N_2794,N_2030);
nand U5866 (N_5866,N_2189,N_2925);
xnor U5867 (N_5867,N_2543,N_827);
or U5868 (N_5868,N_1195,N_995);
nand U5869 (N_5869,N_2193,N_645);
nand U5870 (N_5870,N_1105,N_1735);
or U5871 (N_5871,N_1957,N_1538);
and U5872 (N_5872,N_2441,N_386);
nor U5873 (N_5873,N_2017,N_2610);
nand U5874 (N_5874,N_341,N_2764);
nand U5875 (N_5875,N_1039,N_2198);
xor U5876 (N_5876,N_220,N_1793);
or U5877 (N_5877,N_985,N_1285);
nand U5878 (N_5878,N_2973,N_2041);
or U5879 (N_5879,N_2122,N_2168);
nand U5880 (N_5880,N_1749,N_2682);
or U5881 (N_5881,N_1944,N_704);
nand U5882 (N_5882,N_679,N_2297);
nand U5883 (N_5883,N_905,N_743);
nand U5884 (N_5884,N_2700,N_2026);
nor U5885 (N_5885,N_2912,N_1254);
and U5886 (N_5886,N_2192,N_1540);
or U5887 (N_5887,N_2531,N_2943);
nand U5888 (N_5888,N_2187,N_39);
nand U5889 (N_5889,N_464,N_2205);
nand U5890 (N_5890,N_3003,N_1234);
nand U5891 (N_5891,N_1811,N_2462);
nand U5892 (N_5892,N_3090,N_1749);
nor U5893 (N_5893,N_810,N_421);
or U5894 (N_5894,N_3061,N_2862);
or U5895 (N_5895,N_89,N_611);
nor U5896 (N_5896,N_283,N_2436);
nand U5897 (N_5897,N_139,N_1234);
or U5898 (N_5898,N_2972,N_334);
nand U5899 (N_5899,N_2116,N_703);
xor U5900 (N_5900,N_419,N_1524);
or U5901 (N_5901,N_526,N_792);
nand U5902 (N_5902,N_405,N_196);
or U5903 (N_5903,N_218,N_238);
nor U5904 (N_5904,N_2749,N_1315);
xnor U5905 (N_5905,N_2780,N_1204);
xnor U5906 (N_5906,N_2132,N_385);
nand U5907 (N_5907,N_2386,N_1097);
nand U5908 (N_5908,N_734,N_2410);
or U5909 (N_5909,N_1160,N_1995);
nand U5910 (N_5910,N_3032,N_2274);
nor U5911 (N_5911,N_329,N_1836);
nand U5912 (N_5912,N_420,N_945);
nand U5913 (N_5913,N_959,N_1683);
or U5914 (N_5914,N_2541,N_979);
nand U5915 (N_5915,N_1885,N_265);
xnor U5916 (N_5916,N_3074,N_523);
xnor U5917 (N_5917,N_2829,N_1364);
or U5918 (N_5918,N_2270,N_573);
or U5919 (N_5919,N_739,N_2758);
nand U5920 (N_5920,N_0,N_2976);
or U5921 (N_5921,N_556,N_1084);
nor U5922 (N_5922,N_167,N_82);
nand U5923 (N_5923,N_1220,N_2155);
or U5924 (N_5924,N_1798,N_98);
xnor U5925 (N_5925,N_1275,N_1915);
nor U5926 (N_5926,N_2484,N_1323);
nor U5927 (N_5927,N_2173,N_1827);
nor U5928 (N_5928,N_279,N_2136);
and U5929 (N_5929,N_2795,N_544);
and U5930 (N_5930,N_288,N_161);
and U5931 (N_5931,N_1912,N_2187);
and U5932 (N_5932,N_1710,N_2695);
nand U5933 (N_5933,N_2643,N_1565);
nand U5934 (N_5934,N_1063,N_1141);
or U5935 (N_5935,N_2683,N_1148);
xnor U5936 (N_5936,N_2392,N_1007);
nor U5937 (N_5937,N_1684,N_2886);
nand U5938 (N_5938,N_1859,N_1129);
and U5939 (N_5939,N_2238,N_2162);
and U5940 (N_5940,N_1790,N_587);
xor U5941 (N_5941,N_2140,N_2974);
or U5942 (N_5942,N_1707,N_2359);
nor U5943 (N_5943,N_276,N_2984);
or U5944 (N_5944,N_1874,N_698);
and U5945 (N_5945,N_344,N_2418);
xor U5946 (N_5946,N_759,N_293);
and U5947 (N_5947,N_557,N_1759);
nor U5948 (N_5948,N_274,N_1352);
nor U5949 (N_5949,N_7,N_837);
nor U5950 (N_5950,N_869,N_49);
nand U5951 (N_5951,N_2043,N_2455);
nor U5952 (N_5952,N_1295,N_911);
nor U5953 (N_5953,N_59,N_510);
and U5954 (N_5954,N_1401,N_553);
and U5955 (N_5955,N_827,N_542);
and U5956 (N_5956,N_1852,N_1565);
and U5957 (N_5957,N_2090,N_2092);
nor U5958 (N_5958,N_996,N_255);
and U5959 (N_5959,N_1833,N_1886);
or U5960 (N_5960,N_1059,N_1211);
nand U5961 (N_5961,N_1649,N_741);
nor U5962 (N_5962,N_275,N_109);
and U5963 (N_5963,N_1763,N_1402);
and U5964 (N_5964,N_891,N_1818);
nand U5965 (N_5965,N_1809,N_3016);
nand U5966 (N_5966,N_2751,N_10);
xor U5967 (N_5967,N_2910,N_2212);
nand U5968 (N_5968,N_2077,N_2554);
nor U5969 (N_5969,N_1434,N_1199);
nor U5970 (N_5970,N_317,N_1950);
and U5971 (N_5971,N_2936,N_855);
nor U5972 (N_5972,N_947,N_670);
xnor U5973 (N_5973,N_1599,N_351);
and U5974 (N_5974,N_1537,N_1746);
or U5975 (N_5975,N_1972,N_1825);
nor U5976 (N_5976,N_2476,N_664);
nor U5977 (N_5977,N_111,N_744);
and U5978 (N_5978,N_1696,N_582);
and U5979 (N_5979,N_216,N_60);
xnor U5980 (N_5980,N_2630,N_47);
nor U5981 (N_5981,N_1952,N_1549);
nand U5982 (N_5982,N_2160,N_616);
nor U5983 (N_5983,N_253,N_1796);
nor U5984 (N_5984,N_1254,N_1962);
nor U5985 (N_5985,N_16,N_1131);
and U5986 (N_5986,N_1874,N_389);
and U5987 (N_5987,N_141,N_307);
nor U5988 (N_5988,N_1342,N_2235);
nor U5989 (N_5989,N_1913,N_2021);
nor U5990 (N_5990,N_1263,N_2111);
nor U5991 (N_5991,N_1066,N_1154);
nand U5992 (N_5992,N_1640,N_1893);
nand U5993 (N_5993,N_2023,N_680);
or U5994 (N_5994,N_1101,N_1231);
and U5995 (N_5995,N_3004,N_1898);
and U5996 (N_5996,N_1815,N_1206);
or U5997 (N_5997,N_2447,N_2713);
nor U5998 (N_5998,N_225,N_499);
nand U5999 (N_5999,N_3028,N_920);
and U6000 (N_6000,N_1161,N_2013);
or U6001 (N_6001,N_1377,N_2858);
and U6002 (N_6002,N_915,N_1164);
and U6003 (N_6003,N_1169,N_2134);
xor U6004 (N_6004,N_974,N_1022);
or U6005 (N_6005,N_955,N_1760);
and U6006 (N_6006,N_2578,N_1376);
nor U6007 (N_6007,N_167,N_901);
or U6008 (N_6008,N_257,N_3093);
and U6009 (N_6009,N_2116,N_784);
or U6010 (N_6010,N_1704,N_1957);
nand U6011 (N_6011,N_196,N_1453);
nand U6012 (N_6012,N_1028,N_395);
or U6013 (N_6013,N_1227,N_260);
or U6014 (N_6014,N_1295,N_2039);
nor U6015 (N_6015,N_1201,N_528);
or U6016 (N_6016,N_2443,N_2656);
nor U6017 (N_6017,N_2701,N_1213);
xor U6018 (N_6018,N_147,N_504);
and U6019 (N_6019,N_1499,N_1058);
xnor U6020 (N_6020,N_2921,N_1377);
nand U6021 (N_6021,N_907,N_1212);
nor U6022 (N_6022,N_52,N_2839);
nor U6023 (N_6023,N_2828,N_3112);
and U6024 (N_6024,N_1921,N_2714);
nand U6025 (N_6025,N_345,N_1532);
xor U6026 (N_6026,N_1866,N_1351);
nand U6027 (N_6027,N_853,N_2445);
nor U6028 (N_6028,N_1363,N_911);
xnor U6029 (N_6029,N_1056,N_567);
or U6030 (N_6030,N_1716,N_2036);
and U6031 (N_6031,N_1086,N_241);
nand U6032 (N_6032,N_1752,N_706);
nor U6033 (N_6033,N_1103,N_1449);
nand U6034 (N_6034,N_3124,N_245);
nand U6035 (N_6035,N_153,N_2513);
and U6036 (N_6036,N_2228,N_1109);
nor U6037 (N_6037,N_3112,N_2169);
or U6038 (N_6038,N_273,N_3060);
or U6039 (N_6039,N_465,N_762);
nor U6040 (N_6040,N_3098,N_2477);
or U6041 (N_6041,N_2640,N_1700);
or U6042 (N_6042,N_168,N_1399);
xnor U6043 (N_6043,N_1907,N_2440);
nor U6044 (N_6044,N_2944,N_1645);
nor U6045 (N_6045,N_978,N_1325);
nand U6046 (N_6046,N_2157,N_437);
nor U6047 (N_6047,N_2554,N_2873);
nor U6048 (N_6048,N_2917,N_1985);
and U6049 (N_6049,N_3115,N_848);
and U6050 (N_6050,N_1491,N_713);
nand U6051 (N_6051,N_405,N_1565);
nor U6052 (N_6052,N_2067,N_92);
xnor U6053 (N_6053,N_465,N_2626);
xor U6054 (N_6054,N_2872,N_669);
nand U6055 (N_6055,N_946,N_1234);
or U6056 (N_6056,N_2755,N_796);
and U6057 (N_6057,N_540,N_1039);
or U6058 (N_6058,N_1000,N_1608);
nand U6059 (N_6059,N_1471,N_2287);
xnor U6060 (N_6060,N_2848,N_1304);
nor U6061 (N_6061,N_625,N_416);
nand U6062 (N_6062,N_1949,N_981);
nand U6063 (N_6063,N_763,N_810);
and U6064 (N_6064,N_438,N_282);
xnor U6065 (N_6065,N_3039,N_2779);
or U6066 (N_6066,N_1261,N_2460);
nor U6067 (N_6067,N_883,N_767);
or U6068 (N_6068,N_1347,N_876);
nor U6069 (N_6069,N_442,N_295);
nor U6070 (N_6070,N_520,N_144);
or U6071 (N_6071,N_1294,N_3109);
nand U6072 (N_6072,N_1956,N_229);
xnor U6073 (N_6073,N_670,N_1285);
nand U6074 (N_6074,N_2689,N_704);
and U6075 (N_6075,N_64,N_1977);
nand U6076 (N_6076,N_2650,N_2479);
or U6077 (N_6077,N_616,N_1873);
and U6078 (N_6078,N_2129,N_1470);
xnor U6079 (N_6079,N_1403,N_1580);
nand U6080 (N_6080,N_4,N_784);
and U6081 (N_6081,N_467,N_1985);
xnor U6082 (N_6082,N_209,N_3051);
xnor U6083 (N_6083,N_36,N_1468);
nand U6084 (N_6084,N_2586,N_339);
or U6085 (N_6085,N_2045,N_2737);
nand U6086 (N_6086,N_1459,N_2045);
nor U6087 (N_6087,N_1259,N_885);
nor U6088 (N_6088,N_416,N_2477);
nor U6089 (N_6089,N_800,N_1056);
or U6090 (N_6090,N_2799,N_2443);
nor U6091 (N_6091,N_3025,N_3042);
xnor U6092 (N_6092,N_60,N_2396);
nor U6093 (N_6093,N_576,N_2021);
and U6094 (N_6094,N_1601,N_1931);
nor U6095 (N_6095,N_766,N_2502);
and U6096 (N_6096,N_2077,N_2991);
nor U6097 (N_6097,N_1312,N_2935);
nor U6098 (N_6098,N_3028,N_292);
and U6099 (N_6099,N_257,N_1056);
nand U6100 (N_6100,N_245,N_2352);
or U6101 (N_6101,N_392,N_2112);
or U6102 (N_6102,N_639,N_2207);
and U6103 (N_6103,N_2147,N_1362);
xor U6104 (N_6104,N_616,N_1420);
xor U6105 (N_6105,N_3053,N_275);
or U6106 (N_6106,N_2026,N_2341);
nand U6107 (N_6107,N_1151,N_1738);
or U6108 (N_6108,N_2377,N_974);
nand U6109 (N_6109,N_2848,N_570);
nand U6110 (N_6110,N_289,N_2983);
or U6111 (N_6111,N_975,N_1828);
nand U6112 (N_6112,N_2837,N_1236);
nand U6113 (N_6113,N_1059,N_135);
xor U6114 (N_6114,N_117,N_1165);
or U6115 (N_6115,N_1729,N_1779);
and U6116 (N_6116,N_336,N_416);
nor U6117 (N_6117,N_44,N_196);
nor U6118 (N_6118,N_356,N_1925);
nor U6119 (N_6119,N_2436,N_1903);
nor U6120 (N_6120,N_401,N_803);
and U6121 (N_6121,N_1340,N_2156);
nand U6122 (N_6122,N_674,N_1977);
and U6123 (N_6123,N_1896,N_2609);
nor U6124 (N_6124,N_1623,N_859);
or U6125 (N_6125,N_2032,N_971);
and U6126 (N_6126,N_2143,N_2204);
nor U6127 (N_6127,N_937,N_272);
and U6128 (N_6128,N_951,N_1270);
and U6129 (N_6129,N_2320,N_2189);
nand U6130 (N_6130,N_1153,N_215);
nand U6131 (N_6131,N_2931,N_706);
xor U6132 (N_6132,N_1318,N_2365);
nand U6133 (N_6133,N_473,N_2128);
and U6134 (N_6134,N_272,N_1916);
or U6135 (N_6135,N_887,N_3055);
xnor U6136 (N_6136,N_2909,N_2353);
or U6137 (N_6137,N_2305,N_35);
or U6138 (N_6138,N_1477,N_2082);
nand U6139 (N_6139,N_2688,N_602);
and U6140 (N_6140,N_1435,N_2360);
nor U6141 (N_6141,N_2646,N_2565);
nand U6142 (N_6142,N_338,N_136);
nor U6143 (N_6143,N_2625,N_810);
and U6144 (N_6144,N_2934,N_1588);
or U6145 (N_6145,N_317,N_1971);
nand U6146 (N_6146,N_341,N_746);
or U6147 (N_6147,N_2662,N_2125);
and U6148 (N_6148,N_787,N_1323);
and U6149 (N_6149,N_331,N_1989);
and U6150 (N_6150,N_1834,N_17);
xor U6151 (N_6151,N_1014,N_1857);
or U6152 (N_6152,N_870,N_2699);
nor U6153 (N_6153,N_2592,N_2866);
xor U6154 (N_6154,N_452,N_597);
nand U6155 (N_6155,N_2427,N_774);
nand U6156 (N_6156,N_2594,N_2347);
xnor U6157 (N_6157,N_1415,N_386);
nand U6158 (N_6158,N_2687,N_2067);
and U6159 (N_6159,N_1166,N_1877);
nand U6160 (N_6160,N_1934,N_431);
nor U6161 (N_6161,N_2219,N_2405);
or U6162 (N_6162,N_1758,N_1576);
xor U6163 (N_6163,N_2235,N_1096);
nor U6164 (N_6164,N_236,N_1231);
xnor U6165 (N_6165,N_2771,N_2553);
and U6166 (N_6166,N_2791,N_372);
or U6167 (N_6167,N_2301,N_1494);
nor U6168 (N_6168,N_335,N_2759);
nand U6169 (N_6169,N_2806,N_1869);
nand U6170 (N_6170,N_2074,N_1033);
or U6171 (N_6171,N_2680,N_723);
or U6172 (N_6172,N_2723,N_647);
and U6173 (N_6173,N_442,N_372);
and U6174 (N_6174,N_3029,N_349);
xor U6175 (N_6175,N_2185,N_405);
and U6176 (N_6176,N_2532,N_2653);
nor U6177 (N_6177,N_1879,N_415);
nand U6178 (N_6178,N_2881,N_1537);
or U6179 (N_6179,N_2769,N_695);
nand U6180 (N_6180,N_813,N_494);
and U6181 (N_6181,N_120,N_861);
nor U6182 (N_6182,N_1457,N_192);
or U6183 (N_6183,N_1097,N_661);
nor U6184 (N_6184,N_194,N_1614);
or U6185 (N_6185,N_806,N_2106);
xnor U6186 (N_6186,N_1971,N_1265);
xnor U6187 (N_6187,N_2955,N_1454);
nand U6188 (N_6188,N_1697,N_1714);
or U6189 (N_6189,N_3088,N_2132);
xnor U6190 (N_6190,N_600,N_2834);
or U6191 (N_6191,N_2155,N_1509);
or U6192 (N_6192,N_549,N_1258);
or U6193 (N_6193,N_2477,N_2197);
nor U6194 (N_6194,N_189,N_1524);
nor U6195 (N_6195,N_1191,N_1503);
and U6196 (N_6196,N_1850,N_2612);
nor U6197 (N_6197,N_2681,N_2706);
nand U6198 (N_6198,N_2837,N_1153);
nand U6199 (N_6199,N_3067,N_613);
nor U6200 (N_6200,N_643,N_2369);
nand U6201 (N_6201,N_525,N_1473);
or U6202 (N_6202,N_869,N_2366);
xor U6203 (N_6203,N_468,N_2901);
or U6204 (N_6204,N_2029,N_921);
nor U6205 (N_6205,N_1580,N_2565);
and U6206 (N_6206,N_641,N_2425);
nand U6207 (N_6207,N_2473,N_1066);
nand U6208 (N_6208,N_1102,N_134);
and U6209 (N_6209,N_1825,N_3099);
and U6210 (N_6210,N_157,N_105);
xor U6211 (N_6211,N_1337,N_1010);
nor U6212 (N_6212,N_2625,N_553);
nand U6213 (N_6213,N_2827,N_1040);
or U6214 (N_6214,N_843,N_1732);
or U6215 (N_6215,N_102,N_441);
or U6216 (N_6216,N_2593,N_1423);
nor U6217 (N_6217,N_1000,N_1053);
nor U6218 (N_6218,N_1054,N_1347);
xnor U6219 (N_6219,N_2419,N_2735);
or U6220 (N_6220,N_434,N_1114);
nand U6221 (N_6221,N_1998,N_654);
or U6222 (N_6222,N_1662,N_2703);
xnor U6223 (N_6223,N_1780,N_634);
and U6224 (N_6224,N_225,N_163);
nor U6225 (N_6225,N_659,N_2018);
nor U6226 (N_6226,N_1175,N_840);
nor U6227 (N_6227,N_96,N_1245);
nor U6228 (N_6228,N_1488,N_1022);
xnor U6229 (N_6229,N_1231,N_1303);
or U6230 (N_6230,N_2209,N_2464);
nand U6231 (N_6231,N_3000,N_2495);
nor U6232 (N_6232,N_3049,N_1726);
xor U6233 (N_6233,N_2644,N_1591);
or U6234 (N_6234,N_2671,N_2715);
nor U6235 (N_6235,N_2505,N_322);
nand U6236 (N_6236,N_2047,N_257);
nor U6237 (N_6237,N_1904,N_2290);
xnor U6238 (N_6238,N_1456,N_1842);
and U6239 (N_6239,N_2193,N_614);
nor U6240 (N_6240,N_2735,N_2354);
xnor U6241 (N_6241,N_3117,N_2816);
xnor U6242 (N_6242,N_1749,N_3086);
xor U6243 (N_6243,N_1524,N_1383);
nand U6244 (N_6244,N_1018,N_2753);
nor U6245 (N_6245,N_3017,N_599);
nor U6246 (N_6246,N_2821,N_2771);
and U6247 (N_6247,N_124,N_822);
nand U6248 (N_6248,N_1511,N_1012);
and U6249 (N_6249,N_2797,N_2401);
nor U6250 (N_6250,N_5997,N_4941);
nor U6251 (N_6251,N_5255,N_4853);
nand U6252 (N_6252,N_3133,N_4308);
xor U6253 (N_6253,N_4358,N_4498);
and U6254 (N_6254,N_5204,N_4045);
nand U6255 (N_6255,N_5798,N_4126);
nor U6256 (N_6256,N_5631,N_4894);
xnor U6257 (N_6257,N_5550,N_5589);
or U6258 (N_6258,N_4887,N_6170);
and U6259 (N_6259,N_3642,N_5858);
and U6260 (N_6260,N_3312,N_4106);
nor U6261 (N_6261,N_3988,N_3405);
nand U6262 (N_6262,N_6247,N_3180);
nor U6263 (N_6263,N_4344,N_4008);
nor U6264 (N_6264,N_4871,N_5021);
or U6265 (N_6265,N_6192,N_4018);
and U6266 (N_6266,N_3281,N_4702);
or U6267 (N_6267,N_5657,N_5496);
and U6268 (N_6268,N_4841,N_5555);
xnor U6269 (N_6269,N_4290,N_4738);
nand U6270 (N_6270,N_6124,N_4671);
nor U6271 (N_6271,N_4957,N_3655);
or U6272 (N_6272,N_3840,N_3130);
nand U6273 (N_6273,N_3709,N_3350);
nand U6274 (N_6274,N_4513,N_5075);
xor U6275 (N_6275,N_5375,N_3975);
and U6276 (N_6276,N_5837,N_5775);
xnor U6277 (N_6277,N_5179,N_5231);
xor U6278 (N_6278,N_3858,N_5150);
nand U6279 (N_6279,N_3168,N_3558);
nand U6280 (N_6280,N_3538,N_4087);
and U6281 (N_6281,N_5392,N_3569);
nor U6282 (N_6282,N_4166,N_3607);
nor U6283 (N_6283,N_4028,N_4701);
and U6284 (N_6284,N_4915,N_3458);
and U6285 (N_6285,N_4333,N_5915);
or U6286 (N_6286,N_4378,N_3227);
or U6287 (N_6287,N_5245,N_5801);
xor U6288 (N_6288,N_3377,N_4985);
and U6289 (N_6289,N_5730,N_5558);
nand U6290 (N_6290,N_5346,N_3690);
nand U6291 (N_6291,N_4418,N_5403);
or U6292 (N_6292,N_3695,N_3157);
nand U6293 (N_6293,N_5493,N_4973);
nor U6294 (N_6294,N_3364,N_4713);
nand U6295 (N_6295,N_5632,N_4961);
xor U6296 (N_6296,N_3597,N_3480);
xor U6297 (N_6297,N_3796,N_4219);
or U6298 (N_6298,N_3708,N_5729);
or U6299 (N_6299,N_3266,N_4754);
nand U6300 (N_6300,N_3459,N_3342);
nand U6301 (N_6301,N_3927,N_5124);
or U6302 (N_6302,N_6132,N_5752);
nor U6303 (N_6303,N_4710,N_3600);
nand U6304 (N_6304,N_5739,N_3523);
nor U6305 (N_6305,N_5166,N_3482);
xor U6306 (N_6306,N_5673,N_4934);
nand U6307 (N_6307,N_3286,N_4616);
nand U6308 (N_6308,N_5622,N_3518);
and U6309 (N_6309,N_5593,N_3905);
or U6310 (N_6310,N_3341,N_4238);
or U6311 (N_6311,N_3940,N_4584);
or U6312 (N_6312,N_3551,N_3224);
nand U6313 (N_6313,N_3176,N_3825);
nor U6314 (N_6314,N_5289,N_6195);
and U6315 (N_6315,N_5241,N_4505);
nor U6316 (N_6316,N_3931,N_4542);
or U6317 (N_6317,N_3403,N_4861);
and U6318 (N_6318,N_5867,N_5158);
nand U6319 (N_6319,N_5036,N_4406);
and U6320 (N_6320,N_5859,N_4469);
or U6321 (N_6321,N_5749,N_3831);
xnor U6322 (N_6322,N_4003,N_5476);
nand U6323 (N_6323,N_5282,N_3680);
xnor U6324 (N_6324,N_5843,N_3914);
nor U6325 (N_6325,N_3230,N_5051);
or U6326 (N_6326,N_3501,N_4775);
or U6327 (N_6327,N_4092,N_4299);
nor U6328 (N_6328,N_3800,N_5616);
xnor U6329 (N_6329,N_5287,N_3702);
nand U6330 (N_6330,N_5154,N_3284);
nor U6331 (N_6331,N_5503,N_4494);
nand U6332 (N_6332,N_3252,N_3356);
nand U6333 (N_6333,N_5236,N_4407);
nand U6334 (N_6334,N_4569,N_6108);
nand U6335 (N_6335,N_5178,N_3485);
xor U6336 (N_6336,N_6034,N_6164);
xor U6337 (N_6337,N_3460,N_3641);
nand U6338 (N_6338,N_3219,N_5740);
nand U6339 (N_6339,N_3468,N_3141);
and U6340 (N_6340,N_5436,N_4236);
nor U6341 (N_6341,N_4493,N_5006);
nand U6342 (N_6342,N_3369,N_5328);
nor U6343 (N_6343,N_3378,N_6137);
nor U6344 (N_6344,N_4764,N_4518);
nand U6345 (N_6345,N_5463,N_4482);
nor U6346 (N_6346,N_4086,N_4517);
nor U6347 (N_6347,N_5746,N_3615);
nand U6348 (N_6348,N_4611,N_5385);
nor U6349 (N_6349,N_5055,N_4351);
or U6350 (N_6350,N_3241,N_5391);
and U6351 (N_6351,N_3235,N_6152);
xor U6352 (N_6352,N_5337,N_4676);
or U6353 (N_6353,N_3838,N_5104);
nand U6354 (N_6354,N_5620,N_3409);
xor U6355 (N_6355,N_6048,N_3763);
nand U6356 (N_6356,N_5102,N_5786);
nand U6357 (N_6357,N_3986,N_4085);
nand U6358 (N_6358,N_5790,N_4684);
nor U6359 (N_6359,N_5086,N_5454);
or U6360 (N_6360,N_3321,N_5895);
xor U6361 (N_6361,N_4162,N_5572);
nand U6362 (N_6362,N_5660,N_3787);
and U6363 (N_6363,N_5052,N_4121);
and U6364 (N_6364,N_3135,N_5306);
and U6365 (N_6365,N_5418,N_4474);
nor U6366 (N_6366,N_3171,N_3414);
nand U6367 (N_6367,N_3146,N_5647);
or U6368 (N_6368,N_4873,N_3140);
xor U6369 (N_6369,N_3408,N_5251);
or U6370 (N_6370,N_3764,N_5240);
and U6371 (N_6371,N_6127,N_4081);
nand U6372 (N_6372,N_4682,N_4888);
nor U6373 (N_6373,N_3593,N_3445);
nor U6374 (N_6374,N_5666,N_6135);
and U6375 (N_6375,N_4382,N_3779);
nand U6376 (N_6376,N_5935,N_6190);
nor U6377 (N_6377,N_3344,N_3532);
or U6378 (N_6378,N_6091,N_3239);
nand U6379 (N_6379,N_4901,N_5203);
or U6380 (N_6380,N_5165,N_4047);
and U6381 (N_6381,N_4264,N_4917);
nor U6382 (N_6382,N_5186,N_3706);
and U6383 (N_6383,N_4163,N_3714);
xnor U6384 (N_6384,N_3812,N_5344);
and U6385 (N_6385,N_6215,N_5380);
nor U6386 (N_6386,N_5275,N_4441);
or U6387 (N_6387,N_3349,N_4457);
xor U6388 (N_6388,N_3736,N_5597);
nand U6389 (N_6389,N_5121,N_6074);
xnor U6390 (N_6390,N_4788,N_5253);
nand U6391 (N_6391,N_4763,N_5683);
or U6392 (N_6392,N_6008,N_4878);
xor U6393 (N_6393,N_3254,N_4907);
or U6394 (N_6394,N_3343,N_5049);
xor U6395 (N_6395,N_4144,N_3841);
nand U6396 (N_6396,N_3487,N_4113);
xor U6397 (N_6397,N_5119,N_5926);
nand U6398 (N_6398,N_3871,N_4249);
nor U6399 (N_6399,N_4134,N_3739);
nand U6400 (N_6400,N_4452,N_4943);
nor U6401 (N_6401,N_5108,N_4490);
nand U6402 (N_6402,N_3605,N_5111);
or U6403 (N_6403,N_5308,N_4847);
or U6404 (N_6404,N_3731,N_3131);
or U6405 (N_6405,N_4252,N_5031);
and U6406 (N_6406,N_4362,N_3126);
or U6407 (N_6407,N_4443,N_3769);
and U6408 (N_6408,N_6204,N_4412);
xnor U6409 (N_6409,N_4263,N_5794);
xor U6410 (N_6410,N_6196,N_3911);
nor U6411 (N_6411,N_4533,N_5639);
and U6412 (N_6412,N_5387,N_4237);
and U6413 (N_6413,N_4751,N_6066);
and U6414 (N_6414,N_5143,N_4603);
and U6415 (N_6415,N_5812,N_4638);
nand U6416 (N_6416,N_5291,N_4535);
nor U6417 (N_6417,N_5132,N_5233);
nor U6418 (N_6418,N_4034,N_6177);
and U6419 (N_6419,N_5074,N_5654);
nor U6420 (N_6420,N_5553,N_6154);
nand U6421 (N_6421,N_4507,N_4834);
nand U6422 (N_6422,N_4810,N_3910);
and U6423 (N_6423,N_5462,N_5294);
nand U6424 (N_6424,N_5741,N_3339);
or U6425 (N_6425,N_4555,N_3775);
or U6426 (N_6426,N_6227,N_5062);
xor U6427 (N_6427,N_5636,N_5960);
or U6428 (N_6428,N_4963,N_3493);
nand U6429 (N_6429,N_4316,N_3951);
nor U6430 (N_6430,N_5142,N_5085);
and U6431 (N_6431,N_5089,N_5367);
and U6432 (N_6432,N_3232,N_4591);
and U6433 (N_6433,N_6014,N_3370);
nor U6434 (N_6434,N_3301,N_4348);
or U6435 (N_6435,N_4430,N_3550);
or U6436 (N_6436,N_5839,N_5713);
and U6437 (N_6437,N_4207,N_4192);
or U6438 (N_6438,N_6069,N_5548);
nand U6439 (N_6439,N_6222,N_3228);
nor U6440 (N_6440,N_4280,N_4779);
nand U6441 (N_6441,N_4064,N_3952);
nor U6442 (N_6442,N_4795,N_4026);
nor U6443 (N_6443,N_5637,N_6005);
and U6444 (N_6444,N_6083,N_3283);
nand U6445 (N_6445,N_6021,N_6093);
nor U6446 (N_6446,N_3566,N_3999);
nor U6447 (N_6447,N_5678,N_6232);
nor U6448 (N_6448,N_3696,N_5721);
and U6449 (N_6449,N_4697,N_6136);
nor U6450 (N_6450,N_3937,N_5906);
nor U6451 (N_6451,N_3194,N_5448);
nand U6452 (N_6452,N_5516,N_4213);
or U6453 (N_6453,N_4169,N_4090);
nand U6454 (N_6454,N_5875,N_4948);
nor U6455 (N_6455,N_3272,N_5680);
or U6456 (N_6456,N_5948,N_4870);
or U6457 (N_6457,N_4534,N_4341);
and U6458 (N_6458,N_3520,N_5214);
nor U6459 (N_6459,N_5568,N_4544);
nand U6460 (N_6460,N_5930,N_4700);
nor U6461 (N_6461,N_5412,N_3991);
or U6462 (N_6462,N_5822,N_5382);
xor U6463 (N_6463,N_3323,N_3306);
nor U6464 (N_6464,N_5726,N_4402);
and U6465 (N_6465,N_6111,N_3694);
nand U6466 (N_6466,N_5663,N_6140);
nor U6467 (N_6467,N_4874,N_3865);
nor U6468 (N_6468,N_4755,N_5866);
and U6469 (N_6469,N_3397,N_5748);
and U6470 (N_6470,N_5706,N_5148);
or U6471 (N_6471,N_5478,N_6033);
nor U6472 (N_6472,N_6020,N_4691);
xor U6473 (N_6473,N_4501,N_3505);
or U6474 (N_6474,N_5943,N_4271);
and U6475 (N_6475,N_4230,N_3427);
nor U6476 (N_6476,N_3782,N_3287);
or U6477 (N_6477,N_5013,N_4078);
nand U6478 (N_6478,N_4913,N_3436);
nor U6479 (N_6479,N_6178,N_5044);
nor U6480 (N_6480,N_5697,N_4208);
nor U6481 (N_6481,N_3928,N_5507);
nand U6482 (N_6482,N_3648,N_3365);
and U6483 (N_6483,N_6027,N_3293);
and U6484 (N_6484,N_3472,N_5932);
nand U6485 (N_6485,N_4578,N_4596);
and U6486 (N_6486,N_5582,N_4675);
and U6487 (N_6487,N_3795,N_4845);
xnor U6488 (N_6488,N_3936,N_4686);
nor U6489 (N_6489,N_3134,N_3852);
or U6490 (N_6490,N_4612,N_5625);
nor U6491 (N_6491,N_4746,N_4389);
nand U6492 (N_6492,N_3688,N_5796);
nor U6493 (N_6493,N_5987,N_4562);
and U6494 (N_6494,N_4373,N_5410);
or U6495 (N_6495,N_5197,N_4397);
nor U6496 (N_6496,N_3837,N_4286);
or U6497 (N_6497,N_5343,N_4849);
or U6498 (N_6498,N_3616,N_3554);
or U6499 (N_6499,N_6028,N_5621);
and U6500 (N_6500,N_4979,N_5038);
or U6501 (N_6501,N_3514,N_5146);
or U6502 (N_6502,N_4854,N_3467);
nor U6503 (N_6503,N_6026,N_5365);
nand U6504 (N_6504,N_4458,N_3751);
or U6505 (N_6505,N_3741,N_3274);
and U6506 (N_6506,N_4575,N_3900);
xor U6507 (N_6507,N_3816,N_5147);
nor U6508 (N_6508,N_6173,N_5850);
xor U6509 (N_6509,N_3955,N_3643);
or U6510 (N_6510,N_5844,N_4273);
nor U6511 (N_6511,N_3440,N_4855);
and U6512 (N_6512,N_3476,N_5904);
or U6513 (N_6513,N_4274,N_4978);
nand U6514 (N_6514,N_3964,N_4019);
nor U6515 (N_6515,N_3412,N_5945);
nor U6516 (N_6516,N_3529,N_3296);
nor U6517 (N_6517,N_4525,N_3510);
nor U6518 (N_6518,N_4939,N_5633);
or U6519 (N_6519,N_5341,N_4602);
or U6520 (N_6520,N_5902,N_4868);
or U6521 (N_6521,N_3161,N_6166);
nand U6522 (N_6522,N_3165,N_4265);
or U6523 (N_6523,N_6015,N_3475);
nor U6524 (N_6524,N_5851,N_5198);
nor U6525 (N_6525,N_3139,N_5816);
and U6526 (N_6526,N_4567,N_4075);
or U6527 (N_6527,N_4622,N_3229);
nor U6528 (N_6528,N_3868,N_3579);
or U6529 (N_6529,N_4381,N_3572);
or U6530 (N_6530,N_5059,N_5724);
and U6531 (N_6531,N_5345,N_5520);
or U6532 (N_6532,N_3374,N_3760);
and U6533 (N_6533,N_4224,N_3155);
or U6534 (N_6534,N_3954,N_5468);
nor U6535 (N_6535,N_3417,N_4410);
and U6536 (N_6536,N_4395,N_5262);
nand U6537 (N_6537,N_3638,N_5682);
or U6538 (N_6538,N_4905,N_5514);
and U6539 (N_6539,N_5457,N_3701);
nand U6540 (N_6540,N_5878,N_5508);
nor U6541 (N_6541,N_3953,N_4541);
xnor U6542 (N_6542,N_5787,N_5040);
xnor U6543 (N_6543,N_6003,N_5598);
and U6544 (N_6544,N_5070,N_4666);
or U6545 (N_6545,N_3899,N_3639);
nor U6546 (N_6546,N_3742,N_3687);
or U6547 (N_6547,N_4516,N_4711);
nor U6548 (N_6548,N_5669,N_4226);
nand U6549 (N_6549,N_3150,N_5979);
xnor U6550 (N_6550,N_5171,N_3767);
xor U6551 (N_6551,N_5750,N_4023);
nand U6552 (N_6552,N_3512,N_5848);
nor U6553 (N_6553,N_5982,N_4212);
or U6554 (N_6554,N_4970,N_5248);
and U6555 (N_6555,N_4718,N_3710);
nand U6556 (N_6556,N_5975,N_4315);
nand U6557 (N_6557,N_5309,N_3861);
nor U6558 (N_6558,N_3732,N_4731);
xnor U6559 (N_6559,N_5641,N_4789);
or U6560 (N_6560,N_3471,N_5889);
or U6561 (N_6561,N_5250,N_5224);
or U6562 (N_6562,N_5082,N_6145);
nor U6563 (N_6563,N_4532,N_4173);
nor U6564 (N_6564,N_5474,N_5076);
xnor U6565 (N_6565,N_4745,N_4929);
nand U6566 (N_6566,N_6209,N_4466);
and U6567 (N_6567,N_4222,N_3362);
nand U6568 (N_6568,N_4831,N_5400);
and U6569 (N_6569,N_4479,N_6009);
nand U6570 (N_6570,N_5128,N_4806);
nor U6571 (N_6571,N_4447,N_4962);
and U6572 (N_6572,N_5529,N_3231);
or U6573 (N_6573,N_3746,N_3586);
nor U6574 (N_6574,N_3172,N_4988);
and U6575 (N_6575,N_4220,N_3531);
nor U6576 (N_6576,N_4820,N_6131);
and U6577 (N_6577,N_3158,N_5937);
nor U6578 (N_6578,N_5939,N_3368);
and U6579 (N_6579,N_3355,N_6105);
xnor U6580 (N_6580,N_6202,N_4445);
and U6581 (N_6581,N_5718,N_4122);
nand U6582 (N_6582,N_3777,N_4423);
nor U6583 (N_6583,N_5556,N_6133);
and U6584 (N_6584,N_6063,N_4215);
or U6585 (N_6585,N_5916,N_4323);
nand U6586 (N_6586,N_3903,N_5467);
and U6587 (N_6587,N_4583,N_5317);
nor U6588 (N_6588,N_4598,N_5766);
and U6589 (N_6589,N_4640,N_4646);
and U6590 (N_6590,N_3498,N_4703);
or U6591 (N_6591,N_4270,N_4214);
or U6592 (N_6592,N_3195,N_4354);
and U6593 (N_6593,N_6045,N_3208);
nand U6594 (N_6594,N_5145,N_6042);
or U6595 (N_6595,N_4422,N_3889);
xnor U6596 (N_6596,N_5684,N_5999);
nor U6597 (N_6597,N_4794,N_4922);
nor U6598 (N_6598,N_3389,N_4179);
and U6599 (N_6599,N_5757,N_6119);
or U6600 (N_6600,N_5411,N_4604);
nor U6601 (N_6601,N_5498,N_5643);
nor U6602 (N_6602,N_3477,N_5484);
nor U6603 (N_6603,N_5709,N_6090);
and U6604 (N_6604,N_5745,N_4097);
xnor U6605 (N_6605,N_3411,N_4866);
nor U6606 (N_6606,N_3949,N_5303);
and U6607 (N_6607,N_4773,N_4859);
or U6608 (N_6608,N_4677,N_5492);
and U6609 (N_6609,N_4167,N_5295);
nand U6610 (N_6610,N_4770,N_4771);
nor U6611 (N_6611,N_4679,N_3466);
nor U6612 (N_6612,N_5826,N_3177);
nand U6613 (N_6613,N_4564,N_3138);
nor U6614 (N_6614,N_4170,N_3624);
xnor U6615 (N_6615,N_3430,N_5627);
or U6616 (N_6616,N_4437,N_5435);
or U6617 (N_6617,N_3401,N_3443);
nand U6618 (N_6618,N_4560,N_3300);
and U6619 (N_6619,N_5857,N_4049);
or U6620 (N_6620,N_4031,N_4054);
or U6621 (N_6621,N_4478,N_4428);
nand U6622 (N_6622,N_5327,N_6084);
and U6623 (N_6623,N_4637,N_3193);
or U6624 (N_6624,N_4625,N_4974);
or U6625 (N_6625,N_3773,N_3259);
and U6626 (N_6626,N_5969,N_3515);
nand U6627 (N_6627,N_5640,N_5398);
or U6628 (N_6628,N_3380,N_5704);
nand U6629 (N_6629,N_5347,N_3620);
xor U6630 (N_6630,N_3473,N_4938);
nand U6631 (N_6631,N_5200,N_4360);
and U6632 (N_6632,N_5330,N_5004);
nor U6633 (N_6633,N_5422,N_4601);
nand U6634 (N_6634,N_4895,N_4607);
and U6635 (N_6635,N_5383,N_4937);
and U6636 (N_6636,N_5202,N_3291);
and U6637 (N_6637,N_3938,N_3273);
and U6638 (N_6638,N_3977,N_5116);
nand U6639 (N_6639,N_3850,N_3214);
nand U6640 (N_6640,N_5360,N_5319);
or U6641 (N_6641,N_3926,N_3497);
nor U6642 (N_6642,N_5190,N_4649);
nand U6643 (N_6643,N_3400,N_4643);
xnor U6644 (N_6644,N_4661,N_5456);
and U6645 (N_6645,N_5105,N_3464);
nor U6646 (N_6646,N_4982,N_4843);
nor U6647 (N_6647,N_5974,N_3814);
or U6648 (N_6648,N_4955,N_5307);
nand U6649 (N_6649,N_4449,N_4319);
xnor U6650 (N_6650,N_4296,N_5695);
nand U6651 (N_6651,N_3757,N_4060);
nand U6652 (N_6652,N_5993,N_4862);
or U6653 (N_6653,N_6078,N_4815);
or U6654 (N_6654,N_4150,N_5494);
nand U6655 (N_6655,N_5043,N_3961);
nand U6656 (N_6656,N_3869,N_3329);
xor U6657 (N_6657,N_4235,N_5151);
or U6658 (N_6658,N_5928,N_4648);
and U6659 (N_6659,N_6022,N_4037);
nor U6660 (N_6660,N_3262,N_4599);
and U6661 (N_6661,N_5434,N_4073);
and U6662 (N_6662,N_4821,N_4337);
nor U6663 (N_6663,N_5769,N_3244);
nor U6664 (N_6664,N_5127,N_5106);
and U6665 (N_6665,N_3817,N_4694);
and U6666 (N_6666,N_4109,N_6087);
xor U6667 (N_6667,N_5862,N_5183);
nor U6668 (N_6668,N_4211,N_4906);
or U6669 (N_6669,N_6126,N_4898);
nor U6670 (N_6670,N_5814,N_5071);
nand U6671 (N_6671,N_5808,N_3338);
and U6672 (N_6672,N_6000,N_4807);
or U6673 (N_6673,N_5656,N_4281);
or U6674 (N_6674,N_3242,N_5451);
or U6675 (N_6675,N_3912,N_5648);
nand U6676 (N_6676,N_5838,N_5429);
and U6677 (N_6677,N_5167,N_5919);
and U6678 (N_6678,N_5182,N_4370);
or U6679 (N_6679,N_4093,N_4084);
nor U6680 (N_6680,N_3125,N_3363);
or U6681 (N_6681,N_4608,N_3653);
and U6682 (N_6682,N_4043,N_4151);
and U6683 (N_6683,N_4867,N_4940);
nor U6684 (N_6684,N_4016,N_4180);
nor U6685 (N_6685,N_5714,N_6184);
nor U6686 (N_6686,N_4971,N_4152);
xor U6687 (N_6687,N_6102,N_3504);
and U6688 (N_6688,N_3454,N_3491);
and U6689 (N_6689,N_4690,N_3879);
or U6690 (N_6690,N_3483,N_5762);
nand U6691 (N_6691,N_5791,N_5716);
nand U6692 (N_6692,N_5000,N_4266);
and U6693 (N_6693,N_3644,N_4155);
or U6694 (N_6694,N_3740,N_4153);
nand U6695 (N_6695,N_5334,N_6031);
nor U6696 (N_6696,N_5504,N_3722);
and U6697 (N_6697,N_6110,N_4617);
and U6698 (N_6698,N_4431,N_3860);
nor U6699 (N_6699,N_3353,N_3884);
nor U6700 (N_6700,N_3629,N_5849);
or U6701 (N_6701,N_5531,N_5285);
nor U6702 (N_6702,N_3189,N_5349);
xor U6703 (N_6703,N_5966,N_4720);
xnor U6704 (N_6704,N_4994,N_4835);
and U6705 (N_6705,N_5546,N_5313);
and U6706 (N_6706,N_4865,N_6198);
nand U6707 (N_6707,N_5103,N_4946);
nand U6708 (N_6708,N_4302,N_3151);
or U6709 (N_6709,N_3453,N_5359);
and U6710 (N_6710,N_5783,N_5747);
or U6711 (N_6711,N_3908,N_4546);
nand U6712 (N_6712,N_3856,N_3891);
xnor U6713 (N_6713,N_5544,N_3539);
and U6714 (N_6714,N_3809,N_5778);
nand U6715 (N_6715,N_3830,N_3589);
xnor U6716 (N_6716,N_3508,N_5026);
nor U6717 (N_6717,N_3528,N_3859);
nor U6718 (N_6718,N_6249,N_5078);
or U6719 (N_6719,N_4719,N_4554);
nor U6720 (N_6720,N_4413,N_4804);
and U6721 (N_6721,N_4645,N_6013);
or U6722 (N_6722,N_4379,N_6006);
nand U6723 (N_6723,N_4394,N_5338);
nor U6724 (N_6724,N_5634,N_4058);
nand U6725 (N_6725,N_3700,N_5962);
nand U6726 (N_6726,N_5624,N_3990);
and U6727 (N_6727,N_4247,N_3849);
and U6728 (N_6728,N_3661,N_3679);
and U6729 (N_6729,N_3906,N_4332);
nor U6730 (N_6730,N_5855,N_4053);
nand U6731 (N_6731,N_4128,N_4130);
or U6732 (N_6732,N_4965,N_3144);
and U6733 (N_6733,N_5094,N_3933);
or U6734 (N_6734,N_6176,N_5908);
nand U6735 (N_6735,N_3627,N_3917);
nor U6736 (N_6736,N_5180,N_5355);
xnor U6737 (N_6737,N_3810,N_3628);
xnor U6738 (N_6738,N_5736,N_4811);
or U6739 (N_6739,N_3402,N_3270);
and U6740 (N_6740,N_5354,N_3206);
nor U6741 (N_6741,N_3308,N_5259);
and U6742 (N_6742,N_4190,N_4784);
or U6743 (N_6743,N_5562,N_6081);
nor U6744 (N_6744,N_3654,N_5755);
and U6745 (N_6745,N_3540,N_4605);
xnor U6746 (N_6746,N_6123,N_5153);
or U6747 (N_6747,N_4914,N_4129);
xnor U6748 (N_6748,N_5773,N_6242);
and U6749 (N_6749,N_4899,N_5139);
and U6750 (N_6750,N_3724,N_4276);
or U6751 (N_6751,N_3452,N_5237);
and U6752 (N_6752,N_5316,N_3275);
and U6753 (N_6753,N_3129,N_5793);
or U6754 (N_6754,N_4580,N_5041);
and U6755 (N_6755,N_4925,N_3184);
nor U6756 (N_6756,N_5888,N_4864);
nor U6757 (N_6757,N_5988,N_4262);
nor U6758 (N_6758,N_5950,N_4805);
nand U6759 (N_6759,N_4248,N_3429);
or U6760 (N_6760,N_3240,N_4156);
and U6761 (N_6761,N_5010,N_5499);
and U6762 (N_6762,N_6076,N_3753);
nor U6763 (N_6763,N_5600,N_6100);
or U6764 (N_6764,N_5617,N_3147);
and U6765 (N_6765,N_4730,N_5221);
nand U6766 (N_6766,N_4477,N_5109);
nor U6767 (N_6767,N_4244,N_4692);
xnor U6768 (N_6768,N_5271,N_4068);
and U6769 (N_6769,N_5008,N_4522);
xor U6770 (N_6770,N_5163,N_5861);
or U6771 (N_6771,N_6079,N_6189);
nor U6772 (N_6772,N_3222,N_5077);
nand U6773 (N_6773,N_3559,N_3652);
or U6774 (N_6774,N_5865,N_5232);
and U6775 (N_6775,N_5545,N_4374);
nand U6776 (N_6776,N_4030,N_3581);
nand U6777 (N_6777,N_3633,N_4935);
nor U6778 (N_6778,N_4797,N_5575);
nor U6779 (N_6779,N_4732,N_6125);
nor U6780 (N_6780,N_5486,N_5276);
nor U6781 (N_6781,N_5399,N_4257);
nand U6782 (N_6782,N_6114,N_3994);
nand U6783 (N_6783,N_4421,N_3367);
nor U6784 (N_6784,N_5570,N_4665);
and U6785 (N_6785,N_4371,N_4356);
and U6786 (N_6786,N_5065,N_4198);
and U6787 (N_6787,N_4653,N_4400);
nand U6788 (N_6788,N_5097,N_5967);
nand U6789 (N_6789,N_3373,N_5426);
or U6790 (N_6790,N_4708,N_4585);
nand U6791 (N_6791,N_3220,N_3944);
and U6792 (N_6792,N_4353,N_4102);
or U6793 (N_6793,N_5811,N_4398);
xor U6794 (N_6794,N_4140,N_4590);
nand U6795 (N_6795,N_5439,N_3295);
or U6796 (N_6796,N_4006,N_4455);
nand U6797 (N_6797,N_3780,N_5452);
or U6798 (N_6798,N_4436,N_3234);
nand U6799 (N_6799,N_4947,N_5610);
nor U6800 (N_6800,N_5577,N_3238);
or U6801 (N_6801,N_5017,N_6118);
nor U6802 (N_6802,N_4147,N_6099);
and U6803 (N_6803,N_3170,N_4499);
or U6804 (N_6804,N_4089,N_4284);
nor U6805 (N_6805,N_4987,N_5110);
and U6806 (N_6806,N_4334,N_3956);
nand U6807 (N_6807,N_3358,N_6153);
or U6808 (N_6808,N_6047,N_3390);
nand U6809 (N_6809,N_5856,N_5366);
and U6810 (N_6810,N_5131,N_5405);
nand U6811 (N_6811,N_3828,N_3196);
or U6812 (N_6812,N_5419,N_3136);
or U6813 (N_6813,N_4620,N_4514);
or U6814 (N_6814,N_4768,N_3328);
or U6815 (N_6815,N_4320,N_5441);
xor U6816 (N_6816,N_3213,N_4002);
nand U6817 (N_6817,N_4258,N_3697);
nand U6818 (N_6818,N_5300,N_5469);
and U6819 (N_6819,N_3167,N_4869);
or U6820 (N_6820,N_4786,N_3386);
and U6821 (N_6821,N_3243,N_3744);
and U6822 (N_6822,N_5893,N_5650);
nor U6823 (N_6823,N_4495,N_4715);
and U6824 (N_6824,N_4067,N_5130);
or U6825 (N_6825,N_5990,N_3299);
nand U6826 (N_6826,N_4877,N_5364);
nand U6827 (N_6827,N_3216,N_4707);
and U6828 (N_6828,N_6055,N_3711);
nor U6829 (N_6829,N_3606,N_5918);
nor U6830 (N_6830,N_3507,N_5623);
and U6831 (N_6831,N_4952,N_4921);
nand U6832 (N_6832,N_5207,N_5540);
nand U6833 (N_6833,N_3997,N_3210);
and U6834 (N_6834,N_5281,N_6072);
or U6835 (N_6835,N_5079,N_4434);
xnor U6836 (N_6836,N_6051,N_4722);
nor U6837 (N_6837,N_3603,N_3320);
nor U6838 (N_6838,N_3251,N_4662);
nand U6839 (N_6839,N_3340,N_4448);
nor U6840 (N_6840,N_5952,N_3748);
or U6841 (N_6841,N_4798,N_3319);
nor U6842 (N_6842,N_3516,N_5042);
and U6843 (N_6843,N_4650,N_5560);
nor U6844 (N_6844,N_4042,N_4814);
nor U6845 (N_6845,N_4012,N_4343);
or U6846 (N_6846,N_5495,N_5871);
and U6847 (N_6847,N_3199,N_3896);
nor U6848 (N_6848,N_5819,N_3667);
and U6849 (N_6849,N_5473,N_3943);
nor U6850 (N_6850,N_4107,N_5835);
nand U6851 (N_6851,N_6057,N_5506);
and U6852 (N_6852,N_6181,N_4829);
nand U6853 (N_6853,N_6044,N_5402);
xor U6854 (N_6854,N_5587,N_3256);
nand U6855 (N_6855,N_3413,N_6213);
and U6856 (N_6856,N_3560,N_4920);
nand U6857 (N_6857,N_3704,N_6201);
and U6858 (N_6858,N_6120,N_6156);
nand U6859 (N_6859,N_4227,N_3137);
or U6860 (N_6860,N_3823,N_4325);
nor U6861 (N_6861,N_3392,N_4767);
and U6862 (N_6862,N_4483,N_3183);
nor U6863 (N_6863,N_6186,N_5482);
xor U6864 (N_6864,N_4099,N_5003);
nor U6865 (N_6865,N_5743,N_5388);
and U6866 (N_6866,N_4892,N_5115);
or U6867 (N_6867,N_3960,N_5831);
and U6868 (N_6868,N_4912,N_6217);
nand U6869 (N_6869,N_4295,N_5907);
nand U6870 (N_6870,N_4189,N_4769);
xor U6871 (N_6871,N_5421,N_6160);
and U6872 (N_6872,N_4743,N_5828);
nand U6873 (N_6873,N_3737,N_5376);
and U6874 (N_6874,N_3771,N_5242);
nand U6875 (N_6875,N_4217,N_5113);
nand U6876 (N_6876,N_5881,N_3492);
or U6877 (N_6877,N_3939,N_4573);
nand U6878 (N_6878,N_5804,N_5981);
nand U6879 (N_6879,N_5315,N_4204);
or U6880 (N_6880,N_5428,N_5258);
nor U6881 (N_6881,N_5257,N_4318);
and U6882 (N_6882,N_4285,N_4832);
or U6883 (N_6883,N_3182,N_6151);
and U6884 (N_6884,N_3438,N_4218);
xor U6885 (N_6885,N_5764,N_5566);
and U6886 (N_6886,N_4880,N_5226);
and U6887 (N_6887,N_4556,N_4059);
nand U6888 (N_6888,N_4655,N_5220);
nor U6889 (N_6889,N_5712,N_4813);
nor U6890 (N_6890,N_3451,N_5063);
or U6891 (N_6891,N_5222,N_3596);
and U6892 (N_6892,N_5088,N_6062);
and U6893 (N_6893,N_5170,N_4446);
and U6894 (N_6894,N_3185,N_4468);
or U6895 (N_6895,N_5715,N_5260);
and U6896 (N_6896,N_5708,N_4311);
nor U6897 (N_6897,N_3576,N_3250);
nand U6898 (N_6898,N_3713,N_3406);
and U6899 (N_6899,N_5585,N_5369);
nand U6900 (N_6900,N_4626,N_4052);
xor U6901 (N_6901,N_6001,N_4799);
nor U6902 (N_6902,N_4496,N_3307);
and U6903 (N_6903,N_5523,N_3826);
or U6904 (N_6904,N_3618,N_5135);
and U6905 (N_6905,N_4021,N_4651);
or U6906 (N_6906,N_4124,N_4330);
nand U6907 (N_6907,N_4793,N_5466);
nor U6908 (N_6908,N_5005,N_4762);
and U6909 (N_6909,N_3298,N_4540);
nor U6910 (N_6910,N_4464,N_4013);
and U6911 (N_6911,N_5490,N_4621);
nor U6912 (N_6912,N_3651,N_4138);
or U6913 (N_6913,N_4275,N_5920);
xor U6914 (N_6914,N_4372,N_5933);
nand U6915 (N_6915,N_3893,N_6097);
and U6916 (N_6916,N_5710,N_4277);
and U6917 (N_6917,N_6179,N_4716);
xor U6918 (N_6918,N_6224,N_5921);
nand U6919 (N_6919,N_6054,N_3449);
or U6920 (N_6920,N_5032,N_3422);
nor U6921 (N_6921,N_6168,N_5393);
or U6922 (N_6922,N_4444,N_3792);
xnor U6923 (N_6923,N_5619,N_4071);
nand U6924 (N_6924,N_3257,N_4897);
nor U6925 (N_6925,N_6207,N_4142);
nand U6926 (N_6926,N_5984,N_4737);
nand U6927 (N_6927,N_3945,N_3882);
nor U6928 (N_6928,N_4061,N_3621);
nor U6929 (N_6929,N_5465,N_5483);
xor U6930 (N_6930,N_3426,N_5235);
and U6931 (N_6931,N_4680,N_5693);
xor U6932 (N_6932,N_3573,N_3853);
nand U6933 (N_6933,N_4688,N_4891);
or U6934 (N_6934,N_5256,N_3957);
nand U6935 (N_6935,N_5318,N_5530);
and U6936 (N_6936,N_4949,N_4486);
nand U6937 (N_6937,N_3571,N_3315);
nand U6938 (N_6938,N_5863,N_5264);
or U6939 (N_6939,N_5581,N_5266);
xor U6940 (N_6940,N_5357,N_6024);
nor U6941 (N_6941,N_4307,N_5956);
and U6942 (N_6942,N_5827,N_6052);
nand U6943 (N_6943,N_4900,N_3236);
nand U6944 (N_6944,N_5156,N_5035);
nor U6945 (N_6945,N_6117,N_3890);
nand U6946 (N_6946,N_4736,N_4191);
and U6947 (N_6947,N_3676,N_5929);
nor U6948 (N_6948,N_5547,N_5213);
or U6949 (N_6949,N_5813,N_4440);
xnor U6950 (N_6950,N_4100,N_6130);
nand U6951 (N_6951,N_4069,N_4916);
nor U6952 (N_6952,N_5157,N_5776);
nand U6953 (N_6953,N_4568,N_5297);
nand U6954 (N_6954,N_6228,N_3590);
or U6955 (N_6955,N_5014,N_5563);
nor U6956 (N_6956,N_4234,N_3885);
or U6957 (N_6957,N_5539,N_5368);
or U6958 (N_6958,N_5754,N_3970);
or U6959 (N_6959,N_5509,N_5007);
and U6960 (N_6960,N_6129,N_6162);
nand U6961 (N_6961,N_3857,N_3872);
nand U6962 (N_6962,N_4678,N_5965);
and U6963 (N_6963,N_5057,N_3292);
nor U6964 (N_6964,N_3756,N_3870);
nor U6965 (N_6965,N_4659,N_3658);
and U6966 (N_6966,N_6010,N_4693);
or U6967 (N_6967,N_3502,N_5302);
or U6968 (N_6968,N_6038,N_3749);
or U6969 (N_6969,N_5832,N_3984);
xor U6970 (N_6970,N_3985,N_6075);
and U6971 (N_6971,N_3425,N_4055);
or U6972 (N_6972,N_5025,N_5949);
xor U6973 (N_6973,N_5215,N_4808);
or U6974 (N_6974,N_5126,N_5719);
or U6975 (N_6975,N_3381,N_5940);
or U6976 (N_6976,N_3264,N_6187);
nand U6977 (N_6977,N_3447,N_3934);
or U6978 (N_6978,N_5665,N_3759);
and U6979 (N_6979,N_4357,N_3707);
nor U6980 (N_6980,N_3657,N_5358);
or U6981 (N_6981,N_5442,N_4586);
nor U6982 (N_6982,N_5460,N_5187);
nand U6983 (N_6983,N_4827,N_6218);
nand U6984 (N_6984,N_5134,N_3824);
nor U6985 (N_6985,N_4077,N_4328);
and U6986 (N_6986,N_5842,N_4964);
nand U6987 (N_6987,N_4223,N_6161);
nor U6988 (N_6988,N_3778,N_5272);
and U6989 (N_6989,N_3574,N_5868);
or U6990 (N_6990,N_4705,N_5395);
and U6991 (N_6991,N_5066,N_5459);
nand U6992 (N_6992,N_3191,N_3922);
nor U6993 (N_6993,N_6144,N_5912);
and U6994 (N_6994,N_5525,N_4576);
nor U6995 (N_6995,N_3173,N_4687);
and U6996 (N_6996,N_3203,N_3790);
nand U6997 (N_6997,N_4391,N_5175);
nor U6998 (N_6998,N_4120,N_5537);
or U6999 (N_6999,N_4383,N_3594);
xor U7000 (N_7000,N_5011,N_4403);
nor U7001 (N_7001,N_3279,N_3563);
nor U7002 (N_7002,N_5825,N_4041);
nor U7003 (N_7003,N_3181,N_5759);
nand U7004 (N_7004,N_3781,N_4139);
nand U7005 (N_7005,N_5475,N_3490);
nand U7006 (N_7006,N_5958,N_4324);
or U7007 (N_7007,N_3280,N_3612);
or U7008 (N_7008,N_4565,N_5686);
nand U7009 (N_7009,N_4463,N_4322);
or U7010 (N_7010,N_6122,N_3552);
and U7011 (N_7011,N_4209,N_5155);
and U7012 (N_7012,N_3484,N_6167);
or U7013 (N_7013,N_3217,N_6210);
nand U7014 (N_7014,N_4765,N_5261);
nor U7015 (N_7015,N_5642,N_5588);
nand U7016 (N_7016,N_5996,N_4511);
xnor U7017 (N_7017,N_5314,N_4597);
xor U7018 (N_7018,N_3248,N_4384);
or U7019 (N_7019,N_3604,N_4176);
xor U7020 (N_7020,N_3820,N_5980);
nand U7021 (N_7021,N_5247,N_5394);
or U7022 (N_7022,N_6096,N_3916);
or U7023 (N_7023,N_5350,N_6165);
or U7024 (N_7024,N_4046,N_5961);
and U7025 (N_7025,N_3245,N_4088);
nand U7026 (N_7026,N_5019,N_3610);
nor U7027 (N_7027,N_5033,N_4112);
or U7028 (N_7028,N_4654,N_5322);
xor U7029 (N_7029,N_4740,N_5101);
nand U7030 (N_7030,N_3768,N_6214);
or U7031 (N_7031,N_4136,N_4902);
nor U7032 (N_7032,N_4986,N_3384);
and U7033 (N_7033,N_3276,N_3419);
nand U7034 (N_7034,N_3950,N_3774);
nor U7035 (N_7035,N_5733,N_6041);
and U7036 (N_7036,N_5977,N_6243);
nand U7037 (N_7037,N_4840,N_3979);
and U7038 (N_7038,N_5817,N_4566);
xnor U7039 (N_7039,N_5497,N_5853);
xor U7040 (N_7040,N_5707,N_4036);
xor U7041 (N_7041,N_5022,N_5717);
or U7042 (N_7042,N_3288,N_6231);
and U7043 (N_7043,N_3348,N_5941);
and U7044 (N_7044,N_5847,N_3684);
nand U7045 (N_7045,N_5596,N_6205);
nand U7046 (N_7046,N_3650,N_4893);
nor U7047 (N_7047,N_4581,N_4174);
and U7048 (N_7048,N_4930,N_5413);
nand U7049 (N_7049,N_3354,N_5181);
and U7050 (N_7050,N_6169,N_4577);
nand U7051 (N_7051,N_5205,N_6088);
xnor U7052 (N_7052,N_3941,N_4137);
nor U7053 (N_7053,N_3424,N_4639);
nand U7054 (N_7054,N_4812,N_4245);
nand U7055 (N_7055,N_3717,N_4287);
or U7056 (N_7056,N_5136,N_5536);
or U7057 (N_7057,N_6175,N_3862);
nand U7058 (N_7058,N_6061,N_4386);
or U7059 (N_7059,N_5732,N_4510);
and U7060 (N_7060,N_4735,N_5924);
or U7061 (N_7061,N_3148,N_4748);
nor U7062 (N_7062,N_5872,N_3303);
or U7063 (N_7063,N_5534,N_4414);
nor U7064 (N_7064,N_5885,N_5053);
or U7065 (N_7065,N_4051,N_4618);
or U7066 (N_7066,N_5860,N_3544);
or U7067 (N_7067,N_3673,N_5018);
or U7068 (N_7068,N_4255,N_3439);
or U7069 (N_7069,N_4559,N_4459);
nor U7070 (N_7070,N_3399,N_6200);
xnor U7071 (N_7071,N_4792,N_3670);
and U7072 (N_7072,N_3310,N_3524);
or U7073 (N_7073,N_4945,N_6188);
nor U7074 (N_7074,N_4127,N_5645);
or U7075 (N_7075,N_4216,N_4818);
or U7076 (N_7076,N_3223,N_5505);
or U7077 (N_7077,N_4819,N_4526);
xor U7078 (N_7078,N_3691,N_5100);
nor U7079 (N_7079,N_3500,N_5321);
nor U7080 (N_7080,N_4298,N_5277);
nor U7081 (N_7081,N_5605,N_5661);
nand U7082 (N_7082,N_3553,N_3179);
or U7083 (N_7083,N_5274,N_5430);
and U7084 (N_7084,N_3818,N_4904);
or U7085 (N_7085,N_4177,N_3963);
nand U7086 (N_7086,N_5675,N_4802);
nor U7087 (N_7087,N_6103,N_5614);
nand U7088 (N_7088,N_4200,N_5608);
nand U7089 (N_7089,N_4967,N_3675);
nand U7090 (N_7090,N_3410,N_4256);
and U7091 (N_7091,N_4539,N_4928);
or U7092 (N_7092,N_5607,N_4632);
nor U7093 (N_7093,N_4080,N_4909);
nor U7094 (N_7094,N_3267,N_5886);
or U7095 (N_7095,N_4193,N_4537);
and U7096 (N_7096,N_4953,N_6104);
nor U7097 (N_7097,N_4062,N_5630);
and U7098 (N_7098,N_3798,N_5149);
nand U7099 (N_7099,N_5687,N_3186);
and U7100 (N_7100,N_5658,N_4473);
xor U7101 (N_7101,N_4549,N_3677);
nor U7102 (N_7102,N_4453,N_4185);
or U7103 (N_7103,N_5332,N_4594);
and U7104 (N_7104,N_5362,N_5381);
nand U7105 (N_7105,N_5840,N_5903);
or U7106 (N_7106,N_5061,N_6116);
or U7107 (N_7107,N_4876,N_6146);
nand U7108 (N_7108,N_6229,N_4890);
or U7109 (N_7109,N_5613,N_3334);
or U7110 (N_7110,N_5068,N_4221);
and U7111 (N_7111,N_6233,N_5331);
nand U7112 (N_7112,N_3806,N_3346);
nand U7113 (N_7113,N_5887,N_3821);
or U7114 (N_7114,N_4165,N_4304);
and U7115 (N_7115,N_4149,N_4563);
or U7116 (N_7116,N_5738,N_3918);
nor U7117 (N_7117,N_6089,N_6053);
nand U7118 (N_7118,N_5927,N_4635);
and U7119 (N_7119,N_5761,N_4571);
and U7120 (N_7120,N_5976,N_3803);
or U7121 (N_7121,N_3801,N_6211);
or U7122 (N_7122,N_4774,N_3433);
nor U7123 (N_7123,N_6147,N_5883);
nor U7124 (N_7124,N_3783,N_4942);
and U7125 (N_7125,N_3664,N_3442);
or U7126 (N_7126,N_4131,N_3435);
nor U7127 (N_7127,N_5934,N_6106);
or U7128 (N_7128,N_4657,N_6199);
xnor U7129 (N_7129,N_5649,N_4997);
xor U7130 (N_7130,N_6112,N_5809);
xnor U7131 (N_7131,N_3925,N_4520);
and U7132 (N_7132,N_5532,N_4429);
and U7133 (N_7133,N_6068,N_5760);
nor U7134 (N_7134,N_4314,N_5758);
nand U7135 (N_7135,N_3894,N_3333);
or U7136 (N_7136,N_4558,N_3847);
xor U7137 (N_7137,N_6223,N_4766);
nand U7138 (N_7138,N_3253,N_4306);
xnor U7139 (N_7139,N_5323,N_3888);
nor U7140 (N_7140,N_3297,N_4785);
or U7141 (N_7141,N_6197,N_5290);
and U7142 (N_7142,N_3942,N_3143);
or U7143 (N_7143,N_4613,N_5192);
and U7144 (N_7144,N_6220,N_5821);
or U7145 (N_7145,N_5060,N_4926);
and U7146 (N_7146,N_4432,N_4500);
nor U7147 (N_7147,N_5438,N_5799);
and U7148 (N_7148,N_5407,N_5188);
and U7149 (N_7149,N_6040,N_4588);
or U7150 (N_7150,N_3947,N_3898);
nor U7151 (N_7151,N_4408,N_5162);
and U7152 (N_7152,N_4652,N_3794);
or U7153 (N_7153,N_4609,N_5280);
xor U7154 (N_7154,N_6239,N_5023);
or U7155 (N_7155,N_5283,N_3474);
and U7156 (N_7156,N_4022,N_5194);
or U7157 (N_7157,N_4630,N_3437);
nand U7158 (N_7158,N_4822,N_3218);
nor U7159 (N_7159,N_5882,N_4141);
and U7160 (N_7160,N_3815,N_5440);
and U7161 (N_7161,N_4817,N_4365);
xnor U7162 (N_7162,N_4033,N_4582);
or U7163 (N_7163,N_5189,N_4572);
and U7164 (N_7164,N_4543,N_3163);
nand U7165 (N_7165,N_5579,N_5084);
or U7166 (N_7166,N_5172,N_3237);
and U7167 (N_7167,N_4160,N_3204);
nor U7168 (N_7168,N_3915,N_4133);
and U7169 (N_7169,N_5731,N_5644);
nor U7170 (N_7170,N_5090,N_5638);
or U7171 (N_7171,N_6237,N_4996);
or U7172 (N_7172,N_4689,N_4579);
xnor U7173 (N_7173,N_6094,N_5526);
nor U7174 (N_7174,N_3725,N_4574);
nand U7175 (N_7175,N_3761,N_3376);
and U7176 (N_7176,N_4634,N_5168);
or U7177 (N_7177,N_4194,N_5737);
nor U7178 (N_7178,N_4503,N_3883);
or U7179 (N_7179,N_4592,N_4728);
nor U7180 (N_7180,N_5805,N_3324);
nand U7181 (N_7181,N_5443,N_3535);
nor U7182 (N_7182,N_5092,N_3260);
and U7183 (N_7183,N_4531,N_4641);
xor U7184 (N_7184,N_4345,N_5989);
nor U7185 (N_7185,N_3635,N_3561);
nor U7186 (N_7186,N_5571,N_5095);
nand U7187 (N_7187,N_3517,N_4725);
nand U7188 (N_7188,N_4910,N_4239);
nor U7189 (N_7189,N_3263,N_5679);
nand U7190 (N_7190,N_4240,N_3462);
and U7191 (N_7191,N_4101,N_3920);
and U7192 (N_7192,N_5176,N_3989);
nor U7193 (N_7193,N_3521,N_3387);
nand U7194 (N_7194,N_3623,N_4512);
nor U7195 (N_7195,N_5140,N_3611);
or U7196 (N_7196,N_4027,N_3522);
xor U7197 (N_7197,N_6134,N_3391);
nor U7198 (N_7198,N_3149,N_5371);
or U7199 (N_7199,N_3534,N_3415);
nor U7200 (N_7200,N_3747,N_4475);
and U7201 (N_7201,N_3683,N_4673);
nand U7202 (N_7202,N_3754,N_5963);
or U7203 (N_7203,N_4199,N_4672);
nor U7204 (N_7204,N_5864,N_6071);
nor U7205 (N_7205,N_4739,N_3261);
and U7206 (N_7206,N_4168,N_6216);
nand U7207 (N_7207,N_3978,N_4695);
nand U7208 (N_7208,N_5925,N_5951);
nor U7209 (N_7209,N_4415,N_3662);
and U7210 (N_7210,N_5072,N_4698);
or U7211 (N_7211,N_3745,N_3456);
or U7212 (N_7212,N_5339,N_5971);
nand U7213 (N_7213,N_5286,N_5986);
or U7214 (N_7214,N_3313,N_3221);
nor U7215 (N_7215,N_4492,N_3345);
nor U7216 (N_7216,N_4723,N_5164);
nand U7217 (N_7217,N_3998,N_5401);
nor U7218 (N_7218,N_4419,N_3446);
nand U7219 (N_7219,N_4561,N_4628);
nor U7220 (N_7220,N_4329,N_4860);
nand U7221 (N_7221,N_4206,N_3526);
nand U7222 (N_7222,N_3733,N_3656);
nand U7223 (N_7223,N_5565,N_5159);
or U7224 (N_7224,N_3921,N_5409);
nor U7225 (N_7225,N_3127,N_3200);
or U7226 (N_7226,N_4427,N_3546);
and U7227 (N_7227,N_3330,N_4135);
nor U7228 (N_7228,N_3577,N_6025);
nor U7229 (N_7229,N_3463,N_3705);
and U7230 (N_7230,N_4932,N_4015);
and U7231 (N_7231,N_3770,N_5073);
and U7232 (N_7232,N_3567,N_5777);
nor U7233 (N_7233,N_5774,N_4110);
nor U7234 (N_7234,N_6203,N_3617);
xnor U7235 (N_7235,N_4615,N_4366);
nor U7236 (N_7236,N_3530,N_3547);
or U7237 (N_7237,N_6070,N_5890);
xnor U7238 (N_7238,N_4310,N_5542);
and U7239 (N_7239,N_4405,N_5711);
nor U7240 (N_7240,N_3613,N_4188);
nand U7241 (N_7241,N_3337,N_3983);
nand U7242 (N_7242,N_3269,N_3637);
nand U7243 (N_7243,N_5045,N_3557);
or U7244 (N_7244,N_3630,N_4758);
nor U7245 (N_7245,N_4039,N_4606);
or U7246 (N_7246,N_4484,N_3735);
nor U7247 (N_7247,N_4035,N_5522);
or U7248 (N_7248,N_5219,N_3302);
or U7249 (N_7249,N_3591,N_4401);
or U7250 (N_7250,N_4201,N_5107);
xor U7251 (N_7251,N_3958,N_5690);
and U7252 (N_7252,N_5305,N_5767);
nand U7253 (N_7253,N_4714,N_4595);
nand U7254 (N_7254,N_3314,N_5144);
and U7255 (N_7255,N_5972,N_4456);
nor U7256 (N_7256,N_5611,N_5602);
nor U7257 (N_7257,N_3851,N_5845);
and U7258 (N_7258,N_6221,N_6064);
or U7259 (N_7259,N_3562,N_3686);
and U7260 (N_7260,N_3209,N_5521);
or U7261 (N_7261,N_4830,N_5599);
and U7262 (N_7262,N_4886,N_6182);
nand U7263 (N_7263,N_5458,N_4642);
xor U7264 (N_7264,N_4681,N_5954);
or U7265 (N_7265,N_3525,N_3470);
nor U7266 (N_7266,N_6163,N_5470);
nor U7267 (N_7267,N_4593,N_3864);
and U7268 (N_7268,N_5501,N_4000);
nor U7269 (N_7269,N_5433,N_6149);
or U7270 (N_7270,N_4487,N_4114);
nor U7271 (N_7271,N_5922,N_5576);
nor U7272 (N_7272,N_6049,N_5771);
or U7273 (N_7273,N_4726,N_5720);
or U7274 (N_7274,N_4289,N_4250);
or U7275 (N_7275,N_4232,N_5029);
nand U7276 (N_7276,N_5590,N_4704);
and U7277 (N_7277,N_5420,N_4119);
nand U7278 (N_7278,N_5324,N_5445);
nor U7279 (N_7279,N_4658,N_3738);
nor U7280 (N_7280,N_5612,N_3361);
and U7281 (N_7281,N_5396,N_6241);
nor U7282 (N_7282,N_5549,N_5161);
or U7283 (N_7283,N_3555,N_4610);
nor U7284 (N_7284,N_5342,N_4251);
nor U7285 (N_7285,N_5193,N_4709);
nand U7286 (N_7286,N_5326,N_4780);
nor U7287 (N_7287,N_3626,N_3372);
or U7288 (N_7288,N_5001,N_3226);
nand U7289 (N_7289,N_5824,N_5676);
and U7290 (N_7290,N_4376,N_4683);
or U7291 (N_7291,N_3634,N_6058);
nand U7292 (N_7292,N_5453,N_6086);
and U7293 (N_7293,N_3887,N_5034);
and U7294 (N_7294,N_4787,N_5039);
nand U7295 (N_7295,N_5028,N_6150);
and U7296 (N_7296,N_3904,N_4954);
and U7297 (N_7297,N_5361,N_3875);
and U7298 (N_7298,N_4300,N_5820);
nor U7299 (N_7299,N_5243,N_5009);
and U7300 (N_7300,N_5228,N_5936);
nor U7301 (N_7301,N_4433,N_4007);
nor U7302 (N_7302,N_4148,N_5722);
or U7303 (N_7303,N_3598,N_5087);
nand U7304 (N_7304,N_5512,N_4696);
or U7305 (N_7305,N_4364,N_5770);
or U7306 (N_7306,N_4809,N_4647);
and U7307 (N_7307,N_5320,N_3929);
or U7308 (N_7308,N_4919,N_5129);
or U7309 (N_7309,N_3211,N_5234);
and U7310 (N_7310,N_4753,N_5699);
xnor U7311 (N_7311,N_3835,N_3880);
xor U7312 (N_7312,N_4741,N_4506);
xor U7313 (N_7313,N_4936,N_5551);
and U7314 (N_7314,N_5554,N_4663);
and U7315 (N_7315,N_3479,N_6109);
and U7316 (N_7316,N_5329,N_5117);
and U7317 (N_7317,N_5668,N_5199);
and U7318 (N_7318,N_5333,N_4664);
nor U7319 (N_7319,N_5080,N_4883);
xor U7320 (N_7320,N_5378,N_4347);
or U7321 (N_7321,N_4116,N_4547);
nor U7322 (N_7322,N_6238,N_5894);
and U7323 (N_7323,N_4981,N_5174);
or U7324 (N_7324,N_3396,N_5946);
or U7325 (N_7325,N_5450,N_4272);
and U7326 (N_7326,N_3174,N_4409);
nand U7327 (N_7327,N_5696,N_4203);
nand U7328 (N_7328,N_5635,N_3128);
and U7329 (N_7329,N_3907,N_3382);
nor U7330 (N_7330,N_4184,N_4733);
or U7331 (N_7331,N_3335,N_5414);
and U7332 (N_7332,N_3663,N_4108);
or U7333 (N_7333,N_5177,N_4095);
and U7334 (N_7334,N_6095,N_6012);
nand U7335 (N_7335,N_5725,N_4029);
and U7336 (N_7336,N_4392,N_3819);
xnor U7337 (N_7337,N_3595,N_5870);
nand U7338 (N_7338,N_6234,N_3311);
and U7339 (N_7339,N_5959,N_3968);
and U7340 (N_7340,N_5681,N_4956);
and U7341 (N_7341,N_4388,N_3974);
or U7342 (N_7342,N_4772,N_3488);
and U7343 (N_7343,N_3212,N_4260);
nand U7344 (N_7344,N_5800,N_6155);
and U7345 (N_7345,N_3854,N_5056);
or U7346 (N_7346,N_4291,N_3791);
nand U7347 (N_7347,N_5461,N_6174);
nor U7348 (N_7348,N_4667,N_4816);
and U7349 (N_7349,N_6159,N_5114);
nand U7350 (N_7350,N_5659,N_5874);
nor U7351 (N_7351,N_5160,N_4259);
and U7352 (N_7352,N_6092,N_6158);
nor U7353 (N_7353,N_3752,N_5896);
xnor U7354 (N_7354,N_4712,N_4014);
and U7355 (N_7355,N_5216,N_4960);
or U7356 (N_7356,N_4065,N_5901);
nand U7357 (N_7357,N_5304,N_3448);
and U7358 (N_7358,N_3874,N_3421);
or U7359 (N_7359,N_4368,N_5455);
xor U7360 (N_7360,N_3693,N_6194);
and U7361 (N_7361,N_5561,N_5756);
nand U7362 (N_7362,N_5836,N_5578);
or U7363 (N_7363,N_6060,N_4633);
nor U7364 (N_7364,N_5348,N_4063);
nand U7365 (N_7365,N_5653,N_5584);
xnor U7366 (N_7366,N_5914,N_3285);
nor U7367 (N_7367,N_4614,N_5879);
and U7368 (N_7368,N_4297,N_5688);
or U7369 (N_7369,N_5416,N_5701);
and U7370 (N_7370,N_4267,N_4083);
and U7371 (N_7371,N_3202,N_4181);
or U7372 (N_7372,N_4756,N_3668);
and U7373 (N_7373,N_3587,N_5209);
nor U7374 (N_7374,N_5795,N_5500);
nor U7375 (N_7375,N_3316,N_5609);
nand U7376 (N_7376,N_5024,N_5252);
nand U7377 (N_7377,N_6056,N_6007);
nor U7378 (N_7378,N_4527,N_3317);
nand U7379 (N_7379,N_4066,N_4497);
nor U7380 (N_7380,N_5552,N_5884);
nor U7381 (N_7381,N_5446,N_3489);
xor U7382 (N_7382,N_4801,N_5591);
xnor U7383 (N_7383,N_5246,N_3602);
and U7384 (N_7384,N_4791,N_3309);
xor U7385 (N_7385,N_3666,N_5797);
xor U7386 (N_7386,N_3536,N_5373);
nor U7387 (N_7387,N_5677,N_4872);
or U7388 (N_7388,N_4335,N_4313);
and U7389 (N_7389,N_4485,N_3729);
nand U7390 (N_7390,N_3393,N_3967);
nor U7391 (N_7391,N_5535,N_4462);
or U7392 (N_7392,N_3715,N_4004);
or U7393 (N_7393,N_5763,N_3789);
and U7394 (N_7394,N_4519,N_5911);
xor U7395 (N_7395,N_5511,N_4523);
xor U7396 (N_7396,N_5742,N_5892);
nor U7397 (N_7397,N_4674,N_3327);
nor U7398 (N_7398,N_4828,N_4178);
or U7399 (N_7399,N_5431,N_4972);
or U7400 (N_7400,N_6235,N_5270);
nand U7401 (N_7401,N_5541,N_6246);
or U7402 (N_7402,N_3162,N_5807);
and U7403 (N_7403,N_4488,N_3169);
and U7404 (N_7404,N_5211,N_5652);
and U7405 (N_7405,N_5123,N_5269);
nand U7406 (N_7406,N_4724,N_5768);
or U7407 (N_7407,N_5876,N_3366);
nor U7408 (N_7408,N_3619,N_5626);
nand U7409 (N_7409,N_3154,N_3457);
nor U7410 (N_7410,N_5229,N_3537);
and U7411 (N_7411,N_5296,N_5691);
and U7412 (N_7412,N_4435,N_5298);
and U7413 (N_7413,N_5370,N_5118);
nor U7414 (N_7414,N_5481,N_5938);
or U7415 (N_7415,N_5067,N_4186);
nor U7416 (N_7416,N_5818,N_4305);
xnor U7417 (N_7417,N_4243,N_4995);
xnor U7418 (N_7418,N_4623,N_5254);
nor U7419 (N_7419,N_3799,N_3659);
or U7420 (N_7420,N_4346,N_3892);
and U7421 (N_7421,N_3580,N_3542);
and U7422 (N_7422,N_5628,N_4024);
and U7423 (N_7423,N_3583,N_5427);
and U7424 (N_7424,N_5909,N_3197);
nand U7425 (N_7425,N_6225,N_4349);
or U7426 (N_7426,N_5301,N_5942);
and U7427 (N_7427,N_3478,N_4857);
nor U7428 (N_7428,N_4082,N_5789);
nand U7429 (N_7429,N_4038,N_4552);
and U7430 (N_7430,N_4292,N_5651);
xnor U7431 (N_7431,N_6050,N_4105);
or U7432 (N_7432,N_3543,N_4451);
nor U7433 (N_7433,N_5196,N_3727);
nor U7434 (N_7434,N_5694,N_5137);
and U7435 (N_7435,N_4851,N_4538);
and U7436 (N_7436,N_5218,N_4959);
nor U7437 (N_7437,N_5744,N_3640);
and U7438 (N_7438,N_3142,N_3966);
xor U7439 (N_7439,N_5432,N_6191);
nand U7440 (N_7440,N_3420,N_3188);
xnor U7441 (N_7441,N_5833,N_4759);
or U7442 (N_7442,N_5698,N_5397);
and U7443 (N_7443,N_3494,N_4528);
and U7444 (N_7444,N_6208,N_5230);
nor U7445 (N_7445,N_5406,N_4685);
nor U7446 (N_7446,N_4025,N_3712);
xnor U7447 (N_7447,N_4202,N_5823);
xor U7448 (N_7448,N_5606,N_5880);
and U7449 (N_7449,N_4524,N_4931);
and U7450 (N_7450,N_4393,N_5788);
nor U7451 (N_7451,N_4465,N_5386);
or U7452 (N_7452,N_3418,N_3503);
nor U7453 (N_7453,N_4668,N_5477);
xnor U7454 (N_7454,N_4057,N_3132);
nor U7455 (N_7455,N_5604,N_6128);
nor U7456 (N_7456,N_4856,N_4783);
or U7457 (N_7457,N_3919,N_4187);
nor U7458 (N_7458,N_3632,N_3359);
and U7459 (N_7459,N_5417,N_4196);
nor U7460 (N_7460,N_4750,N_4924);
or U7461 (N_7461,N_4118,N_3878);
and U7462 (N_7462,N_4481,N_6002);
nand U7463 (N_7463,N_3867,N_4670);
xor U7464 (N_7464,N_4001,N_5533);
nand U7465 (N_7465,N_3305,N_5510);
or U7466 (N_7466,N_5734,N_5781);
xnor U7467 (N_7467,N_3511,N_4161);
and U7468 (N_7468,N_3692,N_3855);
and U7469 (N_7469,N_3318,N_4303);
nor U7470 (N_7470,N_3277,N_6011);
and U7471 (N_7471,N_3660,N_4369);
nor U7472 (N_7472,N_5784,N_3282);
or U7473 (N_7473,N_3946,N_5047);
or U7474 (N_7474,N_5310,N_4717);
and U7475 (N_7475,N_4557,N_4999);
nor U7476 (N_7476,N_5325,N_3646);
nand U7477 (N_7477,N_4992,N_4508);
and U7478 (N_7478,N_3336,N_3881);
and U7479 (N_7479,N_5480,N_6212);
xor U7480 (N_7480,N_5335,N_5408);
or U7481 (N_7481,N_3568,N_5779);
nor U7482 (N_7482,N_3836,N_5279);
nor U7483 (N_7483,N_5583,N_5293);
nand U7484 (N_7484,N_4387,N_3866);
and U7485 (N_7485,N_3404,N_5655);
nor U7486 (N_7486,N_4399,N_3614);
nor U7487 (N_7487,N_5299,N_4420);
nand U7488 (N_7488,N_5702,N_5356);
and U7489 (N_7489,N_4903,N_5141);
nand U7490 (N_7490,N_3996,N_4660);
and U7491 (N_7491,N_6244,N_4461);
and U7492 (N_7492,N_4115,N_5288);
nand U7493 (N_7493,N_4933,N_6036);
xor U7494 (N_7494,N_5815,N_4439);
nor U7495 (N_7495,N_3811,N_5225);
nor U7496 (N_7496,N_5058,N_5703);
nand U7497 (N_7497,N_6032,N_4480);
nor U7498 (N_7498,N_4491,N_3265);
or U7499 (N_7499,N_4278,N_4529);
nor U7500 (N_7500,N_3388,N_4923);
nand U7501 (N_7501,N_4205,N_5802);
nand U7502 (N_7502,N_5212,N_4426);
nand U7503 (N_7503,N_5670,N_4375);
nand U7504 (N_7504,N_4233,N_3233);
nand U7505 (N_7505,N_4340,N_5027);
nor U7506 (N_7506,N_3822,N_3431);
xor U7507 (N_7507,N_4111,N_3444);
or U7508 (N_7508,N_3465,N_3608);
nand U7509 (N_7509,N_3246,N_4803);
or U7510 (N_7510,N_5278,N_4079);
nand U7511 (N_7511,N_6035,N_3750);
nor U7512 (N_7512,N_3145,N_3428);
and U7513 (N_7513,N_4145,N_4103);
xnor U7514 (N_7514,N_5064,N_5873);
and U7515 (N_7515,N_3720,N_4396);
xnor U7516 (N_7516,N_6113,N_5877);
nor U7517 (N_7517,N_3873,N_4476);
and U7518 (N_7518,N_5268,N_4117);
nor U7519 (N_7519,N_4644,N_3788);
nor U7520 (N_7520,N_4254,N_3834);
nand U7521 (N_7521,N_3351,N_4172);
nor U7522 (N_7522,N_5978,N_4850);
nand U7523 (N_7523,N_4619,N_4927);
nor U7524 (N_7524,N_5098,N_3805);
and U7525 (N_7525,N_4879,N_4706);
nand U7526 (N_7526,N_4968,N_5618);
and U7527 (N_7527,N_3326,N_5352);
nand U7528 (N_7528,N_5994,N_6004);
nand U7529 (N_7529,N_5518,N_5728);
and U7530 (N_7530,N_4350,N_5249);
or U7531 (N_7531,N_3995,N_5905);
nor U7532 (N_7532,N_6230,N_5464);
or U7533 (N_7533,N_3863,N_6185);
nand U7534 (N_7534,N_5830,N_5753);
nor U7535 (N_7535,N_4044,N_4727);
or U7536 (N_7536,N_3845,N_5449);
or U7537 (N_7537,N_5910,N_5351);
or U7538 (N_7538,N_4450,N_5727);
nor U7539 (N_7539,N_4157,N_3625);
and U7540 (N_7540,N_5185,N_4125);
nand U7541 (N_7541,N_4800,N_5968);
nor U7542 (N_7542,N_3469,N_5692);
and U7543 (N_7543,N_5900,N_6082);
nand U7544 (N_7544,N_5615,N_6248);
nor U7545 (N_7545,N_3848,N_4454);
or U7546 (N_7546,N_4159,N_5841);
nand U7547 (N_7547,N_3383,N_4269);
nand U7548 (N_7548,N_6059,N_3423);
xor U7549 (N_7549,N_4460,N_3682);
or U7550 (N_7550,N_3192,N_6085);
nand U7551 (N_7551,N_4229,N_5569);
and U7552 (N_7552,N_4467,N_4361);
nor U7553 (N_7553,N_4355,N_5502);
and U7554 (N_7554,N_3582,N_4242);
and U7555 (N_7555,N_5336,N_3441);
nor U7556 (N_7556,N_5629,N_3827);
nand U7557 (N_7557,N_4975,N_5834);
nand U7558 (N_7558,N_4336,N_4631);
and U7559 (N_7559,N_3187,N_5543);
xor U7560 (N_7560,N_3570,N_3331);
nor U7561 (N_7561,N_4863,N_3304);
and U7562 (N_7562,N_3699,N_3674);
or U7563 (N_7563,N_3728,N_5415);
or U7564 (N_7564,N_5050,N_5685);
or U7565 (N_7565,N_5538,N_5125);
and U7566 (N_7566,N_3813,N_4833);
nand U7567 (N_7567,N_5970,N_5037);
or U7568 (N_7568,N_5173,N_6077);
nand U7569 (N_7569,N_4846,N_4825);
and U7570 (N_7570,N_5363,N_3772);
nor U7571 (N_7571,N_4331,N_4536);
or U7572 (N_7572,N_5953,N_6143);
nand U7573 (N_7573,N_5664,N_6107);
nand U7574 (N_7574,N_5227,N_4390);
nand U7575 (N_7575,N_3527,N_4380);
and U7576 (N_7576,N_4990,N_5311);
and U7577 (N_7577,N_4076,N_4950);
and U7578 (N_7578,N_3726,N_3371);
and U7579 (N_7579,N_4339,N_6023);
or U7580 (N_7580,N_3698,N_3672);
nand U7581 (N_7581,N_5425,N_3159);
nor U7582 (N_7582,N_5689,N_5700);
nor U7583 (N_7583,N_4848,N_3886);
or U7584 (N_7584,N_4545,N_4424);
nor U7585 (N_7585,N_4246,N_3375);
or U7586 (N_7586,N_3166,N_3533);
xor U7587 (N_7587,N_3545,N_3394);
or U7588 (N_7588,N_3509,N_4983);
and U7589 (N_7589,N_5782,N_6172);
or U7590 (N_7590,N_3290,N_4844);
or U7591 (N_7591,N_4548,N_4472);
and U7592 (N_7592,N_4094,N_5353);
or U7593 (N_7593,N_3549,N_5479);
nor U7594 (N_7594,N_5973,N_5944);
xor U7595 (N_7595,N_5244,N_4839);
nand U7596 (N_7596,N_4020,N_4570);
and U7597 (N_7597,N_4363,N_5217);
and U7598 (N_7598,N_4070,N_5002);
nor U7599 (N_7599,N_6067,N_5772);
nor U7600 (N_7600,N_4998,N_5206);
or U7601 (N_7601,N_4777,N_5389);
or U7602 (N_7602,N_5015,N_5191);
nor U7603 (N_7603,N_4966,N_3793);
nand U7604 (N_7604,N_3909,N_3993);
nor U7605 (N_7605,N_6206,N_6183);
nand U7606 (N_7606,N_3519,N_4553);
xnor U7607 (N_7607,N_4005,N_4404);
and U7608 (N_7608,N_3765,N_5559);
nand U7609 (N_7609,N_3495,N_5580);
nand U7610 (N_7610,N_5444,N_3723);
or U7611 (N_7611,N_4048,N_6101);
nor U7612 (N_7612,N_5955,N_4091);
nor U7613 (N_7613,N_6171,N_3190);
and U7614 (N_7614,N_3584,N_3962);
or U7615 (N_7615,N_4776,N_5957);
and U7616 (N_7616,N_5785,N_6019);
nor U7617 (N_7617,N_4991,N_3948);
or U7618 (N_7618,N_4530,N_3156);
nand U7619 (N_7619,N_6018,N_3599);
xor U7620 (N_7620,N_4911,N_3645);
nand U7621 (N_7621,N_3969,N_3205);
nand U7622 (N_7622,N_3981,N_4377);
nor U7623 (N_7623,N_3160,N_4104);
or U7624 (N_7624,N_4896,N_6240);
or U7625 (N_7625,N_6138,N_5267);
nor U7626 (N_7626,N_4338,N_6065);
nand U7627 (N_7627,N_4509,N_5792);
nand U7628 (N_7628,N_5573,N_4796);
nand U7629 (N_7629,N_6245,N_3647);
or U7630 (N_7630,N_3776,N_3450);
and U7631 (N_7631,N_4183,N_4757);
and U7632 (N_7632,N_4993,N_5527);
or U7633 (N_7633,N_5898,N_4636);
and U7634 (N_7634,N_4210,N_5223);
xnor U7635 (N_7635,N_3992,N_5210);
nor U7636 (N_7636,N_3721,N_4197);
nor U7637 (N_7637,N_6080,N_5515);
and U7638 (N_7638,N_4749,N_4600);
and U7639 (N_7639,N_3902,N_4317);
xnor U7640 (N_7640,N_5081,N_3649);
nand U7641 (N_7641,N_4442,N_4842);
and U7642 (N_7642,N_3578,N_4969);
nand U7643 (N_7643,N_4782,N_5374);
xor U7644 (N_7644,N_3785,N_4417);
or U7645 (N_7645,N_6141,N_5574);
nand U7646 (N_7646,N_4367,N_4438);
and U7647 (N_7647,N_4425,N_5138);
nand U7648 (N_7648,N_4778,N_4098);
xnor U7649 (N_7649,N_3506,N_5765);
xor U7650 (N_7650,N_5646,N_5133);
nand U7651 (N_7651,N_5899,N_4032);
nand U7652 (N_7652,N_5273,N_6226);
or U7653 (N_7653,N_3385,N_5829);
nor U7654 (N_7654,N_3972,N_3575);
and U7655 (N_7655,N_3271,N_5096);
nor U7656 (N_7656,N_5603,N_5284);
or U7657 (N_7657,N_4175,N_4551);
nand U7658 (N_7658,N_4882,N_4908);
nor U7659 (N_7659,N_3976,N_3395);
xnor U7660 (N_7660,N_4359,N_5913);
xor U7661 (N_7661,N_3901,N_3689);
or U7662 (N_7662,N_3496,N_4721);
xnor U7663 (N_7663,N_4228,N_4624);
nor U7664 (N_7664,N_4072,N_5377);
nand U7665 (N_7665,N_5998,N_4164);
nor U7666 (N_7666,N_4321,N_3755);
xor U7667 (N_7667,N_5751,N_4123);
xor U7668 (N_7668,N_6037,N_6098);
nor U7669 (N_7669,N_3548,N_3294);
and U7670 (N_7670,N_4884,N_4146);
nand U7671 (N_7671,N_3434,N_5595);
nand U7672 (N_7672,N_4301,N_5586);
and U7673 (N_7673,N_3766,N_5923);
nand U7674 (N_7674,N_4976,N_4261);
nand U7675 (N_7675,N_5917,N_4989);
nand U7676 (N_7676,N_4918,N_3665);
nand U7677 (N_7677,N_3347,N_5491);
nand U7678 (N_7678,N_3207,N_5723);
nor U7679 (N_7679,N_4288,N_6121);
xnor U7680 (N_7680,N_3877,N_3416);
nand U7681 (N_7681,N_5667,N_3289);
xor U7682 (N_7682,N_5093,N_5263);
nor U7683 (N_7683,N_3432,N_4837);
nand U7684 (N_7684,N_4074,N_4309);
nand U7685 (N_7685,N_5340,N_5120);
or U7686 (N_7686,N_3201,N_4096);
nand U7687 (N_7687,N_5404,N_3153);
nand U7688 (N_7688,N_4282,N_3786);
nor U7689 (N_7689,N_6157,N_3804);
and U7690 (N_7690,N_4342,N_3669);
and U7691 (N_7691,N_5083,N_5069);
nor U7692 (N_7692,N_5869,N_6030);
or U7693 (N_7693,N_3982,N_3685);
nor U7694 (N_7694,N_3332,N_3398);
nand U7695 (N_7695,N_3585,N_4881);
and U7696 (N_7696,N_4889,N_3833);
nor U7697 (N_7697,N_5016,N_5513);
nand U7698 (N_7698,N_3762,N_3730);
xor U7699 (N_7699,N_5594,N_4761);
nand U7700 (N_7700,N_5854,N_4225);
or U7701 (N_7701,N_5671,N_4656);
and U7702 (N_7702,N_3379,N_5995);
nand U7703 (N_7703,N_4010,N_4326);
and U7704 (N_7704,N_3843,N_5992);
nor U7705 (N_7705,N_4781,N_3832);
xor U7706 (N_7706,N_6115,N_6017);
or U7707 (N_7707,N_3322,N_5991);
and U7708 (N_7708,N_4629,N_6219);
xor U7709 (N_7709,N_3980,N_5931);
and U7710 (N_7710,N_5312,N_3897);
nor U7711 (N_7711,N_3178,N_5891);
xnor U7712 (N_7712,N_5048,N_4132);
and U7713 (N_7713,N_4742,N_4283);
nor U7714 (N_7714,N_4587,N_5169);
nor U7715 (N_7715,N_4195,N_3932);
or U7716 (N_7716,N_5488,N_3807);
and U7717 (N_7717,N_3247,N_5810);
nor U7718 (N_7718,N_4515,N_5705);
nor U7719 (N_7719,N_3198,N_3360);
nor U7720 (N_7720,N_5112,N_5672);
nand U7721 (N_7721,N_4171,N_4747);
nand U7722 (N_7722,N_3844,N_3923);
and U7723 (N_7723,N_3541,N_3842);
and U7724 (N_7724,N_3681,N_3930);
nor U7725 (N_7725,N_4744,N_4312);
or U7726 (N_7726,N_3486,N_4984);
xnor U7727 (N_7727,N_5292,N_3987);
or U7728 (N_7728,N_4268,N_5471);
and U7729 (N_7729,N_3631,N_4154);
or U7730 (N_7730,N_3278,N_5238);
or U7731 (N_7731,N_4504,N_5390);
or U7732 (N_7732,N_4470,N_5524);
xor U7733 (N_7733,N_3588,N_4521);
nor U7734 (N_7734,N_4231,N_4858);
nand U7735 (N_7735,N_3513,N_4143);
or U7736 (N_7736,N_4489,N_5437);
nor U7737 (N_7737,N_3935,N_5735);
nor U7738 (N_7738,N_4056,N_4182);
or U7739 (N_7739,N_5519,N_5674);
nor U7740 (N_7740,N_5846,N_4416);
and U7741 (N_7741,N_3784,N_6016);
nor U7742 (N_7742,N_5020,N_4352);
nor U7743 (N_7743,N_3758,N_5384);
nand U7744 (N_7744,N_6039,N_4852);
and U7745 (N_7745,N_4550,N_3461);
nand U7746 (N_7746,N_4411,N_6148);
or U7747 (N_7747,N_5152,N_3965);
nand U7748 (N_7748,N_4951,N_5239);
nand U7749 (N_7749,N_3499,N_5372);
and U7750 (N_7750,N_3352,N_3971);
xnor U7751 (N_7751,N_6046,N_6142);
nor U7752 (N_7752,N_3258,N_4826);
or U7753 (N_7753,N_5091,N_4293);
nor U7754 (N_7754,N_5201,N_5803);
nand U7755 (N_7755,N_5487,N_3152);
or U7756 (N_7756,N_5964,N_5567);
nor U7757 (N_7757,N_3455,N_3718);
nor U7758 (N_7758,N_4823,N_5557);
nand U7759 (N_7759,N_3564,N_4627);
nor U7760 (N_7760,N_5601,N_4158);
and U7761 (N_7761,N_3164,N_3743);
nor U7762 (N_7762,N_5379,N_3407);
nor U7763 (N_7763,N_5485,N_4253);
or U7764 (N_7764,N_6029,N_4734);
nand U7765 (N_7765,N_3876,N_4836);
or U7766 (N_7766,N_5983,N_3215);
nor U7767 (N_7767,N_5472,N_3601);
nor U7768 (N_7768,N_3671,N_3839);
nand U7769 (N_7769,N_4040,N_6236);
or U7770 (N_7770,N_3734,N_5054);
and U7771 (N_7771,N_4958,N_3249);
nand U7772 (N_7772,N_3225,N_4977);
or U7773 (N_7773,N_3895,N_4752);
nor U7774 (N_7774,N_6073,N_4838);
nor U7775 (N_7775,N_5099,N_3357);
nor U7776 (N_7776,N_3829,N_5184);
nand U7777 (N_7777,N_5012,N_5046);
nor U7778 (N_7778,N_4944,N_4790);
and U7779 (N_7779,N_4502,N_3846);
nor U7780 (N_7780,N_5517,N_4385);
nand U7781 (N_7781,N_6180,N_4011);
nand U7782 (N_7782,N_3802,N_3973);
and U7783 (N_7783,N_3636,N_4050);
nand U7784 (N_7784,N_4279,N_3622);
nor U7785 (N_7785,N_5489,N_5564);
or U7786 (N_7786,N_3808,N_3592);
nor U7787 (N_7787,N_3175,N_3556);
nor U7788 (N_7788,N_6193,N_3703);
nor U7789 (N_7789,N_3609,N_3481);
nand U7790 (N_7790,N_5447,N_4327);
nor U7791 (N_7791,N_4471,N_3719);
and U7792 (N_7792,N_3268,N_3325);
nor U7793 (N_7793,N_3678,N_4729);
nor U7794 (N_7794,N_4885,N_4760);
nor U7795 (N_7795,N_5897,N_4824);
nor U7796 (N_7796,N_5780,N_3797);
nand U7797 (N_7797,N_5985,N_4980);
xnor U7798 (N_7798,N_4875,N_6043);
nand U7799 (N_7799,N_5122,N_3913);
nand U7800 (N_7800,N_4589,N_3255);
nor U7801 (N_7801,N_5592,N_4669);
nand U7802 (N_7802,N_3959,N_5030);
xnor U7803 (N_7803,N_5424,N_5947);
and U7804 (N_7804,N_6139,N_3716);
xor U7805 (N_7805,N_3565,N_4699);
or U7806 (N_7806,N_5852,N_4017);
or U7807 (N_7807,N_5662,N_3924);
nand U7808 (N_7808,N_5265,N_4009);
nor U7809 (N_7809,N_5195,N_4294);
and U7810 (N_7810,N_5528,N_4241);
or U7811 (N_7811,N_5423,N_5806);
nand U7812 (N_7812,N_5208,N_5661);
or U7813 (N_7813,N_4349,N_3816);
or U7814 (N_7814,N_5526,N_5748);
and U7815 (N_7815,N_3263,N_3787);
or U7816 (N_7816,N_5047,N_5954);
and U7817 (N_7817,N_3184,N_5167);
xor U7818 (N_7818,N_4625,N_5274);
and U7819 (N_7819,N_4630,N_4370);
and U7820 (N_7820,N_3507,N_5487);
xnor U7821 (N_7821,N_3295,N_5293);
nand U7822 (N_7822,N_4428,N_5829);
or U7823 (N_7823,N_3265,N_4895);
or U7824 (N_7824,N_4377,N_3856);
or U7825 (N_7825,N_3718,N_4585);
nand U7826 (N_7826,N_4811,N_5028);
or U7827 (N_7827,N_5725,N_4989);
and U7828 (N_7828,N_3539,N_3485);
or U7829 (N_7829,N_5605,N_3712);
xor U7830 (N_7830,N_5916,N_5617);
and U7831 (N_7831,N_4391,N_4963);
nor U7832 (N_7832,N_4478,N_3927);
nand U7833 (N_7833,N_4416,N_5319);
nor U7834 (N_7834,N_4667,N_3143);
and U7835 (N_7835,N_5243,N_4224);
nor U7836 (N_7836,N_4903,N_4884);
nor U7837 (N_7837,N_3307,N_3354);
and U7838 (N_7838,N_4138,N_4377);
nand U7839 (N_7839,N_4946,N_4196);
nor U7840 (N_7840,N_5052,N_5618);
or U7841 (N_7841,N_5574,N_5528);
or U7842 (N_7842,N_3424,N_5594);
nand U7843 (N_7843,N_5771,N_3799);
nand U7844 (N_7844,N_6168,N_5053);
xnor U7845 (N_7845,N_3281,N_5047);
xnor U7846 (N_7846,N_3133,N_5453);
and U7847 (N_7847,N_3248,N_5472);
xor U7848 (N_7848,N_6174,N_4782);
and U7849 (N_7849,N_5772,N_5697);
nand U7850 (N_7850,N_5784,N_4182);
or U7851 (N_7851,N_3434,N_4576);
nand U7852 (N_7852,N_4696,N_3868);
nor U7853 (N_7853,N_4174,N_4584);
and U7854 (N_7854,N_5122,N_3635);
or U7855 (N_7855,N_3636,N_4639);
xor U7856 (N_7856,N_4518,N_4057);
nand U7857 (N_7857,N_6183,N_3657);
or U7858 (N_7858,N_6106,N_3331);
nor U7859 (N_7859,N_3853,N_3314);
or U7860 (N_7860,N_5200,N_5126);
and U7861 (N_7861,N_5957,N_6002);
nand U7862 (N_7862,N_3181,N_3324);
and U7863 (N_7863,N_5100,N_3827);
or U7864 (N_7864,N_3599,N_4908);
and U7865 (N_7865,N_6092,N_4908);
or U7866 (N_7866,N_3580,N_3798);
nor U7867 (N_7867,N_4452,N_4142);
nor U7868 (N_7868,N_5172,N_4551);
and U7869 (N_7869,N_4345,N_6203);
and U7870 (N_7870,N_5867,N_6028);
nor U7871 (N_7871,N_3633,N_4759);
nor U7872 (N_7872,N_6249,N_4821);
nor U7873 (N_7873,N_4281,N_5537);
and U7874 (N_7874,N_3931,N_4952);
nor U7875 (N_7875,N_6154,N_4361);
or U7876 (N_7876,N_3632,N_3365);
nor U7877 (N_7877,N_3456,N_6162);
nor U7878 (N_7878,N_5834,N_4605);
or U7879 (N_7879,N_5782,N_4538);
and U7880 (N_7880,N_5359,N_3732);
or U7881 (N_7881,N_4919,N_3755);
and U7882 (N_7882,N_4901,N_3708);
or U7883 (N_7883,N_3166,N_4713);
nor U7884 (N_7884,N_4134,N_4673);
nand U7885 (N_7885,N_5506,N_5742);
and U7886 (N_7886,N_4006,N_4654);
xor U7887 (N_7887,N_3533,N_3951);
or U7888 (N_7888,N_5864,N_3606);
xor U7889 (N_7889,N_4232,N_4533);
and U7890 (N_7890,N_5998,N_4406);
xnor U7891 (N_7891,N_3982,N_3567);
or U7892 (N_7892,N_3863,N_4903);
nor U7893 (N_7893,N_4555,N_5160);
xnor U7894 (N_7894,N_5574,N_5646);
nor U7895 (N_7895,N_4409,N_5391);
nor U7896 (N_7896,N_5472,N_5506);
or U7897 (N_7897,N_6242,N_5852);
nand U7898 (N_7898,N_6014,N_5621);
or U7899 (N_7899,N_5781,N_3545);
or U7900 (N_7900,N_3874,N_6071);
nor U7901 (N_7901,N_3300,N_4301);
or U7902 (N_7902,N_4794,N_3430);
nor U7903 (N_7903,N_4495,N_3269);
or U7904 (N_7904,N_4609,N_3958);
nand U7905 (N_7905,N_4499,N_4257);
or U7906 (N_7906,N_5106,N_3791);
or U7907 (N_7907,N_4553,N_5078);
and U7908 (N_7908,N_3285,N_4978);
nand U7909 (N_7909,N_5667,N_4184);
xnor U7910 (N_7910,N_4458,N_3707);
xor U7911 (N_7911,N_4302,N_3417);
nand U7912 (N_7912,N_4018,N_4546);
or U7913 (N_7913,N_3953,N_3403);
and U7914 (N_7914,N_5412,N_4869);
and U7915 (N_7915,N_3197,N_5116);
nor U7916 (N_7916,N_3142,N_3538);
and U7917 (N_7917,N_6139,N_6038);
nand U7918 (N_7918,N_3533,N_4240);
xor U7919 (N_7919,N_3757,N_3988);
nor U7920 (N_7920,N_4659,N_4987);
or U7921 (N_7921,N_6204,N_5958);
xnor U7922 (N_7922,N_5846,N_3514);
or U7923 (N_7923,N_4420,N_3374);
and U7924 (N_7924,N_4517,N_4874);
xnor U7925 (N_7925,N_5147,N_3226);
nand U7926 (N_7926,N_4158,N_4751);
nand U7927 (N_7927,N_3406,N_4117);
or U7928 (N_7928,N_4803,N_4094);
or U7929 (N_7929,N_6152,N_5179);
nand U7930 (N_7930,N_3196,N_4670);
and U7931 (N_7931,N_5649,N_5330);
nor U7932 (N_7932,N_4321,N_5589);
and U7933 (N_7933,N_4844,N_5746);
nand U7934 (N_7934,N_3980,N_4737);
and U7935 (N_7935,N_5304,N_3329);
nor U7936 (N_7936,N_6054,N_5429);
nand U7937 (N_7937,N_4256,N_5917);
nor U7938 (N_7938,N_4371,N_3185);
and U7939 (N_7939,N_4265,N_4617);
nand U7940 (N_7940,N_5766,N_3802);
and U7941 (N_7941,N_3297,N_6097);
or U7942 (N_7942,N_5329,N_5452);
nand U7943 (N_7943,N_3492,N_5973);
nand U7944 (N_7944,N_4056,N_3384);
or U7945 (N_7945,N_3444,N_5311);
and U7946 (N_7946,N_5435,N_3487);
nor U7947 (N_7947,N_4347,N_5565);
xor U7948 (N_7948,N_4042,N_5920);
nand U7949 (N_7949,N_5662,N_4503);
nand U7950 (N_7950,N_4777,N_5645);
nand U7951 (N_7951,N_3916,N_3315);
nand U7952 (N_7952,N_3515,N_5538);
nor U7953 (N_7953,N_4865,N_4938);
or U7954 (N_7954,N_3811,N_5990);
or U7955 (N_7955,N_4203,N_4548);
nand U7956 (N_7956,N_3899,N_4732);
nor U7957 (N_7957,N_5927,N_3566);
nor U7958 (N_7958,N_4747,N_5017);
nand U7959 (N_7959,N_5376,N_5056);
xnor U7960 (N_7960,N_6167,N_5040);
or U7961 (N_7961,N_3829,N_4636);
or U7962 (N_7962,N_3132,N_5506);
or U7963 (N_7963,N_4123,N_3942);
nor U7964 (N_7964,N_4146,N_3573);
or U7965 (N_7965,N_5390,N_3557);
nand U7966 (N_7966,N_5130,N_5208);
nor U7967 (N_7967,N_4427,N_4646);
nand U7968 (N_7968,N_5316,N_6082);
xor U7969 (N_7969,N_4284,N_5172);
or U7970 (N_7970,N_6219,N_6018);
nand U7971 (N_7971,N_4376,N_4658);
nand U7972 (N_7972,N_5809,N_3726);
or U7973 (N_7973,N_5943,N_4756);
nand U7974 (N_7974,N_5781,N_4486);
or U7975 (N_7975,N_4513,N_5314);
and U7976 (N_7976,N_4137,N_5390);
nor U7977 (N_7977,N_4001,N_5368);
nor U7978 (N_7978,N_3477,N_4646);
or U7979 (N_7979,N_5442,N_5042);
or U7980 (N_7980,N_3216,N_3510);
nor U7981 (N_7981,N_5722,N_6162);
nand U7982 (N_7982,N_5864,N_5166);
nand U7983 (N_7983,N_3473,N_3629);
and U7984 (N_7984,N_3525,N_5330);
or U7985 (N_7985,N_3403,N_5241);
or U7986 (N_7986,N_6232,N_5572);
nor U7987 (N_7987,N_4954,N_6183);
and U7988 (N_7988,N_5144,N_3522);
nor U7989 (N_7989,N_3172,N_6075);
and U7990 (N_7990,N_4929,N_6060);
and U7991 (N_7991,N_3695,N_6216);
and U7992 (N_7992,N_3713,N_6089);
nor U7993 (N_7993,N_4328,N_5894);
xnor U7994 (N_7994,N_5494,N_3673);
nor U7995 (N_7995,N_5551,N_4908);
xor U7996 (N_7996,N_5357,N_4779);
nor U7997 (N_7997,N_5448,N_6020);
and U7998 (N_7998,N_4143,N_5655);
nor U7999 (N_7999,N_3327,N_5989);
nand U8000 (N_8000,N_4326,N_3415);
and U8001 (N_8001,N_3782,N_6022);
nand U8002 (N_8002,N_5939,N_3705);
nor U8003 (N_8003,N_5202,N_4244);
and U8004 (N_8004,N_5419,N_4847);
nor U8005 (N_8005,N_6121,N_5347);
and U8006 (N_8006,N_4985,N_3757);
or U8007 (N_8007,N_3198,N_3622);
nor U8008 (N_8008,N_3424,N_5963);
or U8009 (N_8009,N_3212,N_4963);
and U8010 (N_8010,N_5852,N_3796);
and U8011 (N_8011,N_6046,N_5993);
or U8012 (N_8012,N_4266,N_5671);
and U8013 (N_8013,N_4121,N_3422);
and U8014 (N_8014,N_4749,N_3853);
xor U8015 (N_8015,N_3324,N_5827);
and U8016 (N_8016,N_3568,N_6082);
and U8017 (N_8017,N_5224,N_4500);
or U8018 (N_8018,N_3363,N_5949);
or U8019 (N_8019,N_3971,N_3874);
and U8020 (N_8020,N_3184,N_4999);
nor U8021 (N_8021,N_5661,N_3945);
nor U8022 (N_8022,N_3779,N_5248);
or U8023 (N_8023,N_5091,N_5508);
nor U8024 (N_8024,N_4775,N_4920);
xnor U8025 (N_8025,N_3284,N_5753);
xnor U8026 (N_8026,N_5312,N_4109);
nand U8027 (N_8027,N_5246,N_4276);
or U8028 (N_8028,N_5222,N_5707);
nand U8029 (N_8029,N_4290,N_4895);
nand U8030 (N_8030,N_3777,N_3705);
nor U8031 (N_8031,N_4070,N_5746);
and U8032 (N_8032,N_4411,N_4288);
or U8033 (N_8033,N_4839,N_3507);
nand U8034 (N_8034,N_5208,N_3354);
and U8035 (N_8035,N_4263,N_3606);
xnor U8036 (N_8036,N_5696,N_3497);
nor U8037 (N_8037,N_5566,N_4883);
nor U8038 (N_8038,N_3317,N_6122);
or U8039 (N_8039,N_3420,N_4187);
or U8040 (N_8040,N_4640,N_6068);
nor U8041 (N_8041,N_6238,N_3958);
nand U8042 (N_8042,N_5875,N_4768);
xor U8043 (N_8043,N_3683,N_6209);
nand U8044 (N_8044,N_6121,N_5592);
or U8045 (N_8045,N_6238,N_4453);
nand U8046 (N_8046,N_4832,N_4097);
nand U8047 (N_8047,N_4279,N_4156);
and U8048 (N_8048,N_4509,N_3387);
or U8049 (N_8049,N_5932,N_5679);
xnor U8050 (N_8050,N_5057,N_4956);
nor U8051 (N_8051,N_5526,N_4242);
nor U8052 (N_8052,N_5693,N_4624);
nand U8053 (N_8053,N_3356,N_3312);
xnor U8054 (N_8054,N_5461,N_4512);
and U8055 (N_8055,N_3999,N_4746);
nand U8056 (N_8056,N_4799,N_4269);
nand U8057 (N_8057,N_3466,N_4328);
or U8058 (N_8058,N_5381,N_4315);
and U8059 (N_8059,N_3436,N_4812);
and U8060 (N_8060,N_3345,N_3970);
and U8061 (N_8061,N_6035,N_4916);
xnor U8062 (N_8062,N_4923,N_5239);
and U8063 (N_8063,N_4327,N_4764);
nand U8064 (N_8064,N_4374,N_5791);
xor U8065 (N_8065,N_3592,N_4368);
and U8066 (N_8066,N_4509,N_5210);
or U8067 (N_8067,N_6215,N_5421);
nand U8068 (N_8068,N_3734,N_5293);
and U8069 (N_8069,N_4968,N_3151);
nor U8070 (N_8070,N_4937,N_4089);
and U8071 (N_8071,N_4365,N_5502);
or U8072 (N_8072,N_6099,N_4479);
or U8073 (N_8073,N_5784,N_5483);
nor U8074 (N_8074,N_3866,N_4023);
and U8075 (N_8075,N_3366,N_3956);
nor U8076 (N_8076,N_4901,N_4628);
nand U8077 (N_8077,N_3348,N_6165);
and U8078 (N_8078,N_4112,N_3346);
or U8079 (N_8079,N_5261,N_4631);
nor U8080 (N_8080,N_3339,N_5469);
nor U8081 (N_8081,N_5600,N_5534);
nor U8082 (N_8082,N_3921,N_5590);
and U8083 (N_8083,N_5186,N_3540);
or U8084 (N_8084,N_4308,N_3457);
xnor U8085 (N_8085,N_3748,N_5007);
nand U8086 (N_8086,N_4142,N_4243);
or U8087 (N_8087,N_4021,N_5657);
and U8088 (N_8088,N_4554,N_4089);
and U8089 (N_8089,N_5865,N_5113);
nand U8090 (N_8090,N_5554,N_4417);
nor U8091 (N_8091,N_4731,N_3576);
xnor U8092 (N_8092,N_6016,N_3372);
nand U8093 (N_8093,N_4965,N_5400);
nor U8094 (N_8094,N_4570,N_5258);
and U8095 (N_8095,N_5136,N_4556);
nor U8096 (N_8096,N_4589,N_3425);
nor U8097 (N_8097,N_4660,N_4463);
and U8098 (N_8098,N_3814,N_4553);
nand U8099 (N_8099,N_5259,N_4590);
nand U8100 (N_8100,N_6184,N_4881);
and U8101 (N_8101,N_4766,N_3634);
or U8102 (N_8102,N_5259,N_4747);
nand U8103 (N_8103,N_4857,N_5812);
nand U8104 (N_8104,N_5308,N_4267);
and U8105 (N_8105,N_4011,N_3272);
nor U8106 (N_8106,N_3893,N_3433);
or U8107 (N_8107,N_4745,N_5973);
and U8108 (N_8108,N_5915,N_6208);
nor U8109 (N_8109,N_3240,N_4228);
nor U8110 (N_8110,N_5503,N_4552);
nor U8111 (N_8111,N_4443,N_3207);
nor U8112 (N_8112,N_5119,N_3406);
and U8113 (N_8113,N_4768,N_4630);
or U8114 (N_8114,N_4991,N_3167);
xnor U8115 (N_8115,N_5827,N_5401);
nor U8116 (N_8116,N_6080,N_4308);
nor U8117 (N_8117,N_3180,N_4148);
nor U8118 (N_8118,N_3243,N_5979);
xor U8119 (N_8119,N_4679,N_5767);
or U8120 (N_8120,N_3530,N_6192);
and U8121 (N_8121,N_3976,N_3221);
xnor U8122 (N_8122,N_3290,N_3554);
nor U8123 (N_8123,N_5860,N_5248);
nand U8124 (N_8124,N_6132,N_4561);
and U8125 (N_8125,N_6053,N_3425);
and U8126 (N_8126,N_5410,N_5264);
nand U8127 (N_8127,N_4799,N_3833);
or U8128 (N_8128,N_4832,N_3998);
or U8129 (N_8129,N_5424,N_5991);
nor U8130 (N_8130,N_4218,N_3128);
nor U8131 (N_8131,N_4227,N_5333);
or U8132 (N_8132,N_5099,N_4623);
nand U8133 (N_8133,N_5151,N_5970);
nand U8134 (N_8134,N_5603,N_4323);
xor U8135 (N_8135,N_5395,N_5571);
nand U8136 (N_8136,N_5392,N_3737);
and U8137 (N_8137,N_4737,N_3919);
nor U8138 (N_8138,N_5235,N_5956);
nand U8139 (N_8139,N_3865,N_5190);
nor U8140 (N_8140,N_3194,N_4589);
nor U8141 (N_8141,N_5523,N_5759);
xnor U8142 (N_8142,N_5379,N_6045);
nor U8143 (N_8143,N_3839,N_5220);
xnor U8144 (N_8144,N_4643,N_4208);
or U8145 (N_8145,N_5651,N_4090);
nor U8146 (N_8146,N_5845,N_5889);
nor U8147 (N_8147,N_5055,N_4498);
or U8148 (N_8148,N_5875,N_3279);
nand U8149 (N_8149,N_6131,N_6243);
nand U8150 (N_8150,N_5782,N_3616);
nand U8151 (N_8151,N_3784,N_3399);
or U8152 (N_8152,N_3743,N_5625);
or U8153 (N_8153,N_6199,N_3692);
nand U8154 (N_8154,N_5847,N_3710);
or U8155 (N_8155,N_5723,N_4894);
or U8156 (N_8156,N_3230,N_3971);
or U8157 (N_8157,N_5650,N_3577);
nor U8158 (N_8158,N_4371,N_3845);
and U8159 (N_8159,N_3592,N_4138);
and U8160 (N_8160,N_5324,N_5094);
or U8161 (N_8161,N_5533,N_3536);
and U8162 (N_8162,N_4421,N_3360);
or U8163 (N_8163,N_5335,N_5812);
or U8164 (N_8164,N_3918,N_4715);
nor U8165 (N_8165,N_3725,N_5246);
and U8166 (N_8166,N_4787,N_4986);
or U8167 (N_8167,N_4316,N_4337);
xor U8168 (N_8168,N_4496,N_3752);
nor U8169 (N_8169,N_4857,N_3706);
nor U8170 (N_8170,N_5199,N_5012);
or U8171 (N_8171,N_3774,N_3721);
nor U8172 (N_8172,N_4716,N_5359);
nand U8173 (N_8173,N_5636,N_4946);
nand U8174 (N_8174,N_5555,N_4716);
nand U8175 (N_8175,N_5291,N_5819);
nor U8176 (N_8176,N_4784,N_5016);
nor U8177 (N_8177,N_3570,N_4640);
nand U8178 (N_8178,N_3194,N_4383);
nand U8179 (N_8179,N_4053,N_6224);
or U8180 (N_8180,N_5076,N_5491);
or U8181 (N_8181,N_4736,N_5294);
nor U8182 (N_8182,N_3659,N_5700);
nor U8183 (N_8183,N_5932,N_6054);
nand U8184 (N_8184,N_4295,N_5857);
or U8185 (N_8185,N_3493,N_6117);
and U8186 (N_8186,N_3815,N_4917);
nand U8187 (N_8187,N_5061,N_3163);
and U8188 (N_8188,N_3306,N_5750);
nand U8189 (N_8189,N_4113,N_4591);
nor U8190 (N_8190,N_3920,N_4046);
or U8191 (N_8191,N_4908,N_3885);
nor U8192 (N_8192,N_4654,N_4175);
xnor U8193 (N_8193,N_6074,N_6065);
or U8194 (N_8194,N_3236,N_4383);
nor U8195 (N_8195,N_4919,N_5605);
nand U8196 (N_8196,N_5288,N_5061);
xnor U8197 (N_8197,N_4359,N_3858);
nor U8198 (N_8198,N_5704,N_4823);
or U8199 (N_8199,N_4786,N_5603);
or U8200 (N_8200,N_3833,N_5354);
or U8201 (N_8201,N_5293,N_5880);
and U8202 (N_8202,N_4221,N_4130);
nor U8203 (N_8203,N_4283,N_3333);
or U8204 (N_8204,N_4539,N_5011);
nor U8205 (N_8205,N_4223,N_4429);
or U8206 (N_8206,N_3581,N_3901);
nand U8207 (N_8207,N_3700,N_4512);
nand U8208 (N_8208,N_5595,N_3666);
nor U8209 (N_8209,N_5073,N_5065);
or U8210 (N_8210,N_5779,N_5909);
nand U8211 (N_8211,N_3950,N_5133);
nor U8212 (N_8212,N_4401,N_6014);
nor U8213 (N_8213,N_5031,N_4279);
or U8214 (N_8214,N_4078,N_4867);
nor U8215 (N_8215,N_4557,N_5308);
nand U8216 (N_8216,N_3312,N_5399);
or U8217 (N_8217,N_5227,N_5611);
and U8218 (N_8218,N_3544,N_4652);
or U8219 (N_8219,N_5191,N_5779);
or U8220 (N_8220,N_4284,N_4648);
or U8221 (N_8221,N_5357,N_3260);
and U8222 (N_8222,N_5395,N_5712);
and U8223 (N_8223,N_4843,N_4817);
and U8224 (N_8224,N_4492,N_5124);
or U8225 (N_8225,N_3725,N_6090);
and U8226 (N_8226,N_4344,N_4318);
nor U8227 (N_8227,N_3168,N_5756);
nor U8228 (N_8228,N_6131,N_6154);
and U8229 (N_8229,N_5210,N_4805);
or U8230 (N_8230,N_4518,N_4723);
nor U8231 (N_8231,N_4539,N_5188);
and U8232 (N_8232,N_4745,N_5572);
and U8233 (N_8233,N_3855,N_5745);
and U8234 (N_8234,N_5940,N_5590);
nand U8235 (N_8235,N_6211,N_5041);
and U8236 (N_8236,N_3431,N_4542);
xnor U8237 (N_8237,N_3879,N_5315);
and U8238 (N_8238,N_4084,N_4936);
and U8239 (N_8239,N_3391,N_6147);
nand U8240 (N_8240,N_5133,N_4393);
nor U8241 (N_8241,N_3424,N_5902);
nand U8242 (N_8242,N_3440,N_4389);
and U8243 (N_8243,N_4020,N_4522);
and U8244 (N_8244,N_5529,N_5849);
or U8245 (N_8245,N_6067,N_4643);
and U8246 (N_8246,N_6110,N_4596);
or U8247 (N_8247,N_3762,N_4920);
or U8248 (N_8248,N_4742,N_5300);
nor U8249 (N_8249,N_3875,N_3656);
or U8250 (N_8250,N_4401,N_3797);
or U8251 (N_8251,N_4164,N_4617);
or U8252 (N_8252,N_4150,N_3803);
nor U8253 (N_8253,N_5334,N_5133);
nand U8254 (N_8254,N_5644,N_3314);
and U8255 (N_8255,N_3372,N_4451);
nand U8256 (N_8256,N_5279,N_4905);
nand U8257 (N_8257,N_4741,N_4056);
or U8258 (N_8258,N_4537,N_5266);
nand U8259 (N_8259,N_5174,N_5289);
or U8260 (N_8260,N_3921,N_3802);
nand U8261 (N_8261,N_3187,N_4287);
nor U8262 (N_8262,N_5627,N_3667);
xor U8263 (N_8263,N_4191,N_3780);
nand U8264 (N_8264,N_3497,N_5490);
nor U8265 (N_8265,N_3982,N_5412);
nor U8266 (N_8266,N_5175,N_3695);
and U8267 (N_8267,N_4159,N_5953);
and U8268 (N_8268,N_3164,N_5493);
or U8269 (N_8269,N_3469,N_6027);
nand U8270 (N_8270,N_4030,N_3259);
nor U8271 (N_8271,N_5816,N_3939);
or U8272 (N_8272,N_5137,N_5448);
or U8273 (N_8273,N_3673,N_4634);
or U8274 (N_8274,N_5809,N_3614);
or U8275 (N_8275,N_6053,N_4584);
and U8276 (N_8276,N_4169,N_5119);
and U8277 (N_8277,N_4867,N_4762);
and U8278 (N_8278,N_3905,N_4782);
nand U8279 (N_8279,N_3640,N_4856);
and U8280 (N_8280,N_3253,N_5322);
nor U8281 (N_8281,N_4009,N_5019);
and U8282 (N_8282,N_4324,N_5083);
xor U8283 (N_8283,N_3871,N_5146);
nand U8284 (N_8284,N_5024,N_3666);
or U8285 (N_8285,N_4241,N_4310);
or U8286 (N_8286,N_6225,N_5797);
or U8287 (N_8287,N_5817,N_5745);
or U8288 (N_8288,N_3491,N_4826);
and U8289 (N_8289,N_5989,N_5908);
and U8290 (N_8290,N_5720,N_4711);
nand U8291 (N_8291,N_6166,N_6231);
or U8292 (N_8292,N_6172,N_3995);
and U8293 (N_8293,N_5247,N_5489);
or U8294 (N_8294,N_3176,N_5842);
nor U8295 (N_8295,N_3543,N_4883);
xnor U8296 (N_8296,N_3902,N_3299);
nand U8297 (N_8297,N_5792,N_3474);
nor U8298 (N_8298,N_4778,N_3895);
nor U8299 (N_8299,N_3686,N_3839);
nor U8300 (N_8300,N_4485,N_3858);
nor U8301 (N_8301,N_4640,N_6114);
nor U8302 (N_8302,N_4827,N_4450);
nand U8303 (N_8303,N_4482,N_5474);
and U8304 (N_8304,N_4656,N_4728);
nand U8305 (N_8305,N_5900,N_5658);
or U8306 (N_8306,N_5460,N_5691);
nand U8307 (N_8307,N_5892,N_3616);
nor U8308 (N_8308,N_4534,N_5418);
or U8309 (N_8309,N_5444,N_4723);
nor U8310 (N_8310,N_3769,N_5168);
or U8311 (N_8311,N_5443,N_5521);
or U8312 (N_8312,N_3217,N_4682);
or U8313 (N_8313,N_3208,N_5432);
or U8314 (N_8314,N_4457,N_6076);
nand U8315 (N_8315,N_4138,N_4866);
or U8316 (N_8316,N_3981,N_3337);
and U8317 (N_8317,N_3972,N_5407);
and U8318 (N_8318,N_4774,N_4222);
nor U8319 (N_8319,N_5941,N_3293);
or U8320 (N_8320,N_3554,N_3527);
and U8321 (N_8321,N_3271,N_3439);
nand U8322 (N_8322,N_4793,N_3253);
and U8323 (N_8323,N_3233,N_4035);
or U8324 (N_8324,N_5282,N_4184);
nand U8325 (N_8325,N_5920,N_5244);
nor U8326 (N_8326,N_6050,N_5664);
xor U8327 (N_8327,N_4341,N_3698);
nand U8328 (N_8328,N_3352,N_3448);
and U8329 (N_8329,N_5563,N_3944);
nor U8330 (N_8330,N_3879,N_5363);
nor U8331 (N_8331,N_4712,N_3628);
or U8332 (N_8332,N_4227,N_5491);
and U8333 (N_8333,N_5043,N_5033);
or U8334 (N_8334,N_5913,N_6103);
nor U8335 (N_8335,N_4341,N_5953);
or U8336 (N_8336,N_5328,N_3581);
or U8337 (N_8337,N_5099,N_5898);
nand U8338 (N_8338,N_3792,N_6184);
nor U8339 (N_8339,N_5468,N_4579);
nor U8340 (N_8340,N_5223,N_3844);
or U8341 (N_8341,N_4992,N_3611);
xnor U8342 (N_8342,N_5078,N_4007);
and U8343 (N_8343,N_3768,N_4296);
xor U8344 (N_8344,N_3471,N_5601);
or U8345 (N_8345,N_4595,N_5939);
or U8346 (N_8346,N_3550,N_4237);
or U8347 (N_8347,N_6228,N_3818);
xor U8348 (N_8348,N_3131,N_4023);
or U8349 (N_8349,N_5330,N_5465);
or U8350 (N_8350,N_4207,N_3984);
or U8351 (N_8351,N_4723,N_3596);
or U8352 (N_8352,N_4458,N_3807);
xnor U8353 (N_8353,N_5999,N_4649);
and U8354 (N_8354,N_4507,N_5049);
nand U8355 (N_8355,N_5479,N_4920);
nand U8356 (N_8356,N_5586,N_4660);
xnor U8357 (N_8357,N_3761,N_5773);
or U8358 (N_8358,N_5449,N_4117);
nand U8359 (N_8359,N_6180,N_5719);
nand U8360 (N_8360,N_5975,N_6060);
or U8361 (N_8361,N_5201,N_5673);
or U8362 (N_8362,N_4251,N_3210);
nand U8363 (N_8363,N_5985,N_6065);
or U8364 (N_8364,N_4630,N_4852);
or U8365 (N_8365,N_5607,N_4150);
nand U8366 (N_8366,N_4703,N_3480);
nand U8367 (N_8367,N_5670,N_6201);
nor U8368 (N_8368,N_5816,N_3834);
nor U8369 (N_8369,N_4843,N_6054);
nand U8370 (N_8370,N_5487,N_6176);
nor U8371 (N_8371,N_4227,N_6247);
nand U8372 (N_8372,N_4719,N_5824);
nor U8373 (N_8373,N_4467,N_5425);
xor U8374 (N_8374,N_4022,N_4887);
nor U8375 (N_8375,N_4078,N_4509);
or U8376 (N_8376,N_6182,N_3653);
nor U8377 (N_8377,N_3758,N_5764);
and U8378 (N_8378,N_4477,N_3463);
and U8379 (N_8379,N_5222,N_5855);
nand U8380 (N_8380,N_4657,N_4965);
xor U8381 (N_8381,N_5192,N_5859);
nand U8382 (N_8382,N_5696,N_4244);
xnor U8383 (N_8383,N_5089,N_3461);
nand U8384 (N_8384,N_3589,N_4284);
or U8385 (N_8385,N_5095,N_5613);
nand U8386 (N_8386,N_5429,N_5284);
nor U8387 (N_8387,N_5561,N_4580);
nor U8388 (N_8388,N_5949,N_5188);
and U8389 (N_8389,N_4832,N_4763);
nand U8390 (N_8390,N_5304,N_5020);
and U8391 (N_8391,N_5783,N_3202);
nor U8392 (N_8392,N_6087,N_5113);
and U8393 (N_8393,N_6177,N_5322);
nor U8394 (N_8394,N_5347,N_3330);
and U8395 (N_8395,N_3311,N_4352);
or U8396 (N_8396,N_5375,N_5469);
and U8397 (N_8397,N_3291,N_4745);
nor U8398 (N_8398,N_3362,N_5311);
and U8399 (N_8399,N_4598,N_6133);
xnor U8400 (N_8400,N_4868,N_5083);
and U8401 (N_8401,N_5683,N_4669);
nor U8402 (N_8402,N_4377,N_4307);
nor U8403 (N_8403,N_4777,N_5254);
or U8404 (N_8404,N_4716,N_6130);
and U8405 (N_8405,N_6100,N_4470);
or U8406 (N_8406,N_3572,N_3473);
nand U8407 (N_8407,N_4647,N_4716);
or U8408 (N_8408,N_4913,N_4524);
and U8409 (N_8409,N_3387,N_3797);
and U8410 (N_8410,N_5208,N_5036);
and U8411 (N_8411,N_4202,N_3445);
or U8412 (N_8412,N_3566,N_4635);
and U8413 (N_8413,N_4697,N_5267);
or U8414 (N_8414,N_5330,N_5766);
xor U8415 (N_8415,N_4719,N_3153);
nor U8416 (N_8416,N_4711,N_4490);
nor U8417 (N_8417,N_4356,N_4331);
or U8418 (N_8418,N_5440,N_3226);
and U8419 (N_8419,N_3137,N_4174);
nor U8420 (N_8420,N_5620,N_4794);
xor U8421 (N_8421,N_3295,N_4962);
nand U8422 (N_8422,N_3415,N_5692);
or U8423 (N_8423,N_5151,N_3608);
or U8424 (N_8424,N_6053,N_4676);
or U8425 (N_8425,N_4768,N_3402);
nand U8426 (N_8426,N_5070,N_4426);
nand U8427 (N_8427,N_3748,N_5010);
or U8428 (N_8428,N_4369,N_6106);
and U8429 (N_8429,N_4069,N_3870);
nor U8430 (N_8430,N_4010,N_4764);
nand U8431 (N_8431,N_6213,N_5832);
nor U8432 (N_8432,N_4963,N_3529);
or U8433 (N_8433,N_5333,N_4281);
nand U8434 (N_8434,N_3513,N_3418);
nand U8435 (N_8435,N_5799,N_4218);
or U8436 (N_8436,N_5258,N_5004);
nor U8437 (N_8437,N_3364,N_4576);
nor U8438 (N_8438,N_5310,N_4263);
xor U8439 (N_8439,N_4261,N_3613);
nand U8440 (N_8440,N_4502,N_5641);
xor U8441 (N_8441,N_5844,N_5885);
or U8442 (N_8442,N_6175,N_4667);
nor U8443 (N_8443,N_6134,N_5891);
nor U8444 (N_8444,N_4400,N_4051);
or U8445 (N_8445,N_5184,N_4563);
and U8446 (N_8446,N_5926,N_3924);
and U8447 (N_8447,N_4484,N_3452);
and U8448 (N_8448,N_4016,N_5851);
and U8449 (N_8449,N_4146,N_4977);
and U8450 (N_8450,N_3689,N_4981);
nand U8451 (N_8451,N_5134,N_3967);
nor U8452 (N_8452,N_5240,N_3798);
and U8453 (N_8453,N_4670,N_5544);
nor U8454 (N_8454,N_3693,N_5719);
nand U8455 (N_8455,N_3758,N_3432);
xnor U8456 (N_8456,N_5690,N_5192);
and U8457 (N_8457,N_6049,N_6036);
and U8458 (N_8458,N_5142,N_4569);
xor U8459 (N_8459,N_6115,N_4354);
nor U8460 (N_8460,N_4680,N_3938);
or U8461 (N_8461,N_3147,N_5556);
nor U8462 (N_8462,N_5271,N_5834);
nand U8463 (N_8463,N_6226,N_4065);
xor U8464 (N_8464,N_5447,N_5403);
nor U8465 (N_8465,N_3722,N_4146);
nand U8466 (N_8466,N_3739,N_5377);
or U8467 (N_8467,N_4790,N_5217);
nand U8468 (N_8468,N_5195,N_4997);
nand U8469 (N_8469,N_3215,N_5415);
and U8470 (N_8470,N_3851,N_6053);
nand U8471 (N_8471,N_5863,N_4785);
or U8472 (N_8472,N_3317,N_3981);
or U8473 (N_8473,N_4306,N_4595);
nor U8474 (N_8474,N_5201,N_4667);
nor U8475 (N_8475,N_5673,N_3906);
nand U8476 (N_8476,N_3379,N_5307);
or U8477 (N_8477,N_3780,N_3308);
xor U8478 (N_8478,N_4204,N_3974);
and U8479 (N_8479,N_4851,N_3463);
or U8480 (N_8480,N_4392,N_4755);
nor U8481 (N_8481,N_3332,N_5299);
nor U8482 (N_8482,N_4585,N_3478);
nor U8483 (N_8483,N_3759,N_3153);
and U8484 (N_8484,N_3138,N_5866);
nor U8485 (N_8485,N_5386,N_5750);
nand U8486 (N_8486,N_4558,N_5718);
or U8487 (N_8487,N_5021,N_5212);
and U8488 (N_8488,N_5629,N_4144);
xor U8489 (N_8489,N_5416,N_6014);
nor U8490 (N_8490,N_5199,N_4700);
and U8491 (N_8491,N_4836,N_3588);
nand U8492 (N_8492,N_3308,N_6193);
and U8493 (N_8493,N_4012,N_4837);
or U8494 (N_8494,N_4715,N_5250);
nor U8495 (N_8495,N_3751,N_4816);
and U8496 (N_8496,N_4102,N_4656);
or U8497 (N_8497,N_3248,N_5843);
or U8498 (N_8498,N_6199,N_4312);
or U8499 (N_8499,N_5138,N_4071);
or U8500 (N_8500,N_5949,N_3429);
nand U8501 (N_8501,N_3756,N_3222);
or U8502 (N_8502,N_4201,N_4645);
nand U8503 (N_8503,N_5351,N_3125);
nand U8504 (N_8504,N_3314,N_6029);
nand U8505 (N_8505,N_3285,N_4372);
nand U8506 (N_8506,N_5476,N_4490);
nand U8507 (N_8507,N_5406,N_6224);
or U8508 (N_8508,N_3843,N_5747);
or U8509 (N_8509,N_3192,N_5957);
xnor U8510 (N_8510,N_5271,N_6202);
nor U8511 (N_8511,N_4146,N_5960);
and U8512 (N_8512,N_4182,N_5268);
nand U8513 (N_8513,N_5112,N_3870);
or U8514 (N_8514,N_4759,N_5819);
or U8515 (N_8515,N_4664,N_5046);
and U8516 (N_8516,N_4011,N_3493);
nand U8517 (N_8517,N_4870,N_4942);
nor U8518 (N_8518,N_5991,N_4498);
nor U8519 (N_8519,N_3892,N_5728);
nand U8520 (N_8520,N_4266,N_6207);
or U8521 (N_8521,N_5128,N_5324);
and U8522 (N_8522,N_5428,N_5964);
nand U8523 (N_8523,N_5746,N_4710);
nand U8524 (N_8524,N_6116,N_3195);
and U8525 (N_8525,N_4040,N_5050);
xnor U8526 (N_8526,N_5327,N_3638);
nand U8527 (N_8527,N_4622,N_4481);
or U8528 (N_8528,N_4788,N_3939);
and U8529 (N_8529,N_5496,N_4434);
nor U8530 (N_8530,N_5780,N_3395);
xor U8531 (N_8531,N_3330,N_6159);
and U8532 (N_8532,N_3822,N_5230);
or U8533 (N_8533,N_3647,N_4904);
nand U8534 (N_8534,N_5895,N_4366);
nor U8535 (N_8535,N_5920,N_4495);
and U8536 (N_8536,N_4456,N_6223);
or U8537 (N_8537,N_3926,N_5072);
or U8538 (N_8538,N_3859,N_4457);
nand U8539 (N_8539,N_5670,N_4719);
nor U8540 (N_8540,N_5439,N_4976);
and U8541 (N_8541,N_6118,N_3501);
nor U8542 (N_8542,N_3718,N_5498);
nor U8543 (N_8543,N_3969,N_4330);
nand U8544 (N_8544,N_3928,N_4126);
nand U8545 (N_8545,N_5458,N_6244);
and U8546 (N_8546,N_4706,N_4618);
and U8547 (N_8547,N_5102,N_3806);
nor U8548 (N_8548,N_6103,N_5178);
nor U8549 (N_8549,N_4578,N_5667);
and U8550 (N_8550,N_4174,N_6086);
nand U8551 (N_8551,N_3496,N_3829);
nor U8552 (N_8552,N_4456,N_5264);
or U8553 (N_8553,N_3584,N_6203);
or U8554 (N_8554,N_3320,N_5794);
nand U8555 (N_8555,N_4650,N_4069);
or U8556 (N_8556,N_4265,N_3464);
and U8557 (N_8557,N_5501,N_3405);
and U8558 (N_8558,N_3880,N_4440);
xor U8559 (N_8559,N_4956,N_4578);
or U8560 (N_8560,N_3654,N_4726);
and U8561 (N_8561,N_4825,N_3508);
or U8562 (N_8562,N_3975,N_6037);
nand U8563 (N_8563,N_4191,N_3188);
nand U8564 (N_8564,N_4803,N_3996);
and U8565 (N_8565,N_4348,N_4248);
nor U8566 (N_8566,N_5845,N_6153);
nor U8567 (N_8567,N_4130,N_3572);
nand U8568 (N_8568,N_3183,N_5057);
nand U8569 (N_8569,N_3289,N_5511);
nand U8570 (N_8570,N_5653,N_4971);
and U8571 (N_8571,N_4147,N_3601);
and U8572 (N_8572,N_3407,N_5904);
nand U8573 (N_8573,N_5746,N_4546);
and U8574 (N_8574,N_4072,N_5621);
xor U8575 (N_8575,N_4581,N_5684);
xor U8576 (N_8576,N_6072,N_4383);
nand U8577 (N_8577,N_3921,N_4274);
xnor U8578 (N_8578,N_5554,N_4520);
or U8579 (N_8579,N_4668,N_3520);
or U8580 (N_8580,N_4509,N_4159);
nand U8581 (N_8581,N_5913,N_6214);
or U8582 (N_8582,N_4108,N_5249);
nor U8583 (N_8583,N_5753,N_5805);
or U8584 (N_8584,N_4694,N_4614);
and U8585 (N_8585,N_4260,N_3499);
and U8586 (N_8586,N_4110,N_5800);
nand U8587 (N_8587,N_4198,N_4248);
nor U8588 (N_8588,N_6010,N_6020);
nor U8589 (N_8589,N_4173,N_3595);
nor U8590 (N_8590,N_4172,N_3445);
or U8591 (N_8591,N_5211,N_5372);
xnor U8592 (N_8592,N_6001,N_4288);
nor U8593 (N_8593,N_4397,N_4780);
nand U8594 (N_8594,N_3924,N_4390);
xnor U8595 (N_8595,N_4311,N_6188);
xor U8596 (N_8596,N_4737,N_5470);
and U8597 (N_8597,N_5092,N_4577);
nor U8598 (N_8598,N_3647,N_3817);
xor U8599 (N_8599,N_4104,N_4717);
nand U8600 (N_8600,N_4161,N_4962);
xor U8601 (N_8601,N_3191,N_4852);
nand U8602 (N_8602,N_4950,N_3867);
nor U8603 (N_8603,N_3776,N_3407);
nand U8604 (N_8604,N_4140,N_5306);
or U8605 (N_8605,N_5711,N_5145);
and U8606 (N_8606,N_4081,N_3554);
xnor U8607 (N_8607,N_4472,N_3767);
and U8608 (N_8608,N_3298,N_4808);
and U8609 (N_8609,N_3679,N_3200);
nor U8610 (N_8610,N_4662,N_5431);
and U8611 (N_8611,N_4206,N_4051);
nor U8612 (N_8612,N_5730,N_4374);
xor U8613 (N_8613,N_3840,N_3353);
nand U8614 (N_8614,N_3750,N_5410);
nor U8615 (N_8615,N_3417,N_5132);
nor U8616 (N_8616,N_3647,N_5654);
nor U8617 (N_8617,N_5018,N_6049);
and U8618 (N_8618,N_5713,N_3384);
or U8619 (N_8619,N_5639,N_5445);
or U8620 (N_8620,N_4052,N_3423);
or U8621 (N_8621,N_5426,N_3241);
nand U8622 (N_8622,N_4974,N_5473);
nand U8623 (N_8623,N_6098,N_3292);
and U8624 (N_8624,N_6228,N_4737);
or U8625 (N_8625,N_5454,N_3130);
nor U8626 (N_8626,N_4140,N_3574);
and U8627 (N_8627,N_5210,N_3367);
nor U8628 (N_8628,N_4444,N_5459);
or U8629 (N_8629,N_3627,N_5146);
nand U8630 (N_8630,N_4814,N_4417);
and U8631 (N_8631,N_5493,N_4610);
and U8632 (N_8632,N_5073,N_3154);
or U8633 (N_8633,N_4954,N_4397);
or U8634 (N_8634,N_4233,N_5965);
and U8635 (N_8635,N_3414,N_4555);
and U8636 (N_8636,N_5806,N_4167);
nand U8637 (N_8637,N_5103,N_3933);
nand U8638 (N_8638,N_4931,N_4669);
or U8639 (N_8639,N_3477,N_4185);
and U8640 (N_8640,N_4002,N_3627);
or U8641 (N_8641,N_5404,N_3172);
and U8642 (N_8642,N_3533,N_4083);
nor U8643 (N_8643,N_4732,N_5355);
nor U8644 (N_8644,N_4858,N_4393);
xor U8645 (N_8645,N_3966,N_4584);
nand U8646 (N_8646,N_5852,N_3627);
nand U8647 (N_8647,N_5191,N_4928);
or U8648 (N_8648,N_3547,N_5362);
xor U8649 (N_8649,N_5566,N_5669);
or U8650 (N_8650,N_5755,N_3210);
or U8651 (N_8651,N_3193,N_4388);
nand U8652 (N_8652,N_4340,N_6184);
nor U8653 (N_8653,N_5895,N_6090);
nand U8654 (N_8654,N_5917,N_4560);
or U8655 (N_8655,N_4395,N_5551);
or U8656 (N_8656,N_5750,N_4180);
nor U8657 (N_8657,N_4227,N_4160);
nand U8658 (N_8658,N_5601,N_4014);
or U8659 (N_8659,N_5294,N_3225);
nand U8660 (N_8660,N_3927,N_3200);
nor U8661 (N_8661,N_4485,N_3870);
nor U8662 (N_8662,N_3464,N_3868);
and U8663 (N_8663,N_5392,N_5882);
or U8664 (N_8664,N_4243,N_5413);
nand U8665 (N_8665,N_3651,N_5693);
or U8666 (N_8666,N_4846,N_5296);
or U8667 (N_8667,N_3392,N_4466);
nand U8668 (N_8668,N_3325,N_3201);
and U8669 (N_8669,N_6173,N_5657);
nor U8670 (N_8670,N_5232,N_5637);
nor U8671 (N_8671,N_4091,N_3904);
xor U8672 (N_8672,N_4471,N_3532);
or U8673 (N_8673,N_5620,N_3596);
nor U8674 (N_8674,N_4690,N_4082);
or U8675 (N_8675,N_5250,N_4044);
or U8676 (N_8676,N_3562,N_3744);
nor U8677 (N_8677,N_5854,N_4825);
nor U8678 (N_8678,N_5338,N_3481);
nor U8679 (N_8679,N_3160,N_3888);
or U8680 (N_8680,N_5892,N_4122);
or U8681 (N_8681,N_5054,N_6007);
nand U8682 (N_8682,N_4836,N_5903);
and U8683 (N_8683,N_5927,N_4271);
nand U8684 (N_8684,N_5444,N_5270);
and U8685 (N_8685,N_4388,N_6080);
xnor U8686 (N_8686,N_4515,N_3656);
xnor U8687 (N_8687,N_5087,N_4140);
nand U8688 (N_8688,N_3971,N_3537);
nand U8689 (N_8689,N_3704,N_3960);
nor U8690 (N_8690,N_5772,N_5555);
nand U8691 (N_8691,N_3373,N_3737);
or U8692 (N_8692,N_6183,N_5254);
or U8693 (N_8693,N_6170,N_3893);
xnor U8694 (N_8694,N_5467,N_5390);
nor U8695 (N_8695,N_5835,N_4381);
and U8696 (N_8696,N_5338,N_4905);
and U8697 (N_8697,N_3127,N_4958);
or U8698 (N_8698,N_5086,N_3650);
nand U8699 (N_8699,N_4435,N_3922);
or U8700 (N_8700,N_4235,N_4792);
or U8701 (N_8701,N_5343,N_4543);
nand U8702 (N_8702,N_4980,N_4443);
nand U8703 (N_8703,N_5467,N_5603);
nand U8704 (N_8704,N_5210,N_4088);
or U8705 (N_8705,N_4476,N_4861);
xnor U8706 (N_8706,N_3738,N_5560);
nand U8707 (N_8707,N_6230,N_5949);
or U8708 (N_8708,N_5050,N_5440);
nand U8709 (N_8709,N_3887,N_3648);
nand U8710 (N_8710,N_4410,N_3177);
nor U8711 (N_8711,N_5320,N_5297);
or U8712 (N_8712,N_5276,N_5029);
nand U8713 (N_8713,N_4393,N_4901);
nor U8714 (N_8714,N_5356,N_5042);
nand U8715 (N_8715,N_5480,N_4098);
and U8716 (N_8716,N_4481,N_6106);
nor U8717 (N_8717,N_4433,N_5113);
nor U8718 (N_8718,N_5248,N_6005);
nand U8719 (N_8719,N_3554,N_5453);
and U8720 (N_8720,N_5742,N_3217);
nand U8721 (N_8721,N_3910,N_4576);
xor U8722 (N_8722,N_4548,N_5879);
nand U8723 (N_8723,N_4348,N_3654);
nand U8724 (N_8724,N_3776,N_3300);
and U8725 (N_8725,N_6050,N_3436);
and U8726 (N_8726,N_4481,N_3632);
or U8727 (N_8727,N_5400,N_3914);
xnor U8728 (N_8728,N_4834,N_3355);
and U8729 (N_8729,N_3462,N_4019);
nand U8730 (N_8730,N_5833,N_5309);
or U8731 (N_8731,N_3388,N_5215);
or U8732 (N_8732,N_6070,N_3585);
and U8733 (N_8733,N_4697,N_3416);
nor U8734 (N_8734,N_5668,N_4976);
nor U8735 (N_8735,N_5317,N_5889);
nand U8736 (N_8736,N_5445,N_3341);
nand U8737 (N_8737,N_5485,N_4197);
nor U8738 (N_8738,N_6051,N_4860);
and U8739 (N_8739,N_3301,N_5130);
and U8740 (N_8740,N_3840,N_5535);
and U8741 (N_8741,N_6224,N_3771);
nand U8742 (N_8742,N_3564,N_5517);
xor U8743 (N_8743,N_3597,N_4336);
or U8744 (N_8744,N_5972,N_3190);
or U8745 (N_8745,N_4608,N_4274);
xnor U8746 (N_8746,N_3756,N_3647);
and U8747 (N_8747,N_5345,N_4079);
and U8748 (N_8748,N_4434,N_6090);
xnor U8749 (N_8749,N_5452,N_5204);
nor U8750 (N_8750,N_5600,N_6163);
or U8751 (N_8751,N_4532,N_3565);
nand U8752 (N_8752,N_4367,N_5315);
nand U8753 (N_8753,N_5092,N_5373);
nor U8754 (N_8754,N_5404,N_4042);
and U8755 (N_8755,N_3796,N_5423);
nand U8756 (N_8756,N_4085,N_3924);
nand U8757 (N_8757,N_5450,N_3571);
nor U8758 (N_8758,N_5663,N_5789);
nor U8759 (N_8759,N_5515,N_5544);
and U8760 (N_8760,N_3191,N_5730);
nand U8761 (N_8761,N_3339,N_6068);
nand U8762 (N_8762,N_3638,N_5059);
nor U8763 (N_8763,N_6178,N_3752);
xnor U8764 (N_8764,N_5554,N_4107);
nor U8765 (N_8765,N_5884,N_6217);
nand U8766 (N_8766,N_5633,N_5743);
xnor U8767 (N_8767,N_5783,N_4070);
nand U8768 (N_8768,N_5137,N_5077);
or U8769 (N_8769,N_6179,N_3890);
and U8770 (N_8770,N_4304,N_4025);
and U8771 (N_8771,N_3732,N_4189);
or U8772 (N_8772,N_4510,N_4272);
nand U8773 (N_8773,N_3831,N_4873);
and U8774 (N_8774,N_5439,N_5804);
and U8775 (N_8775,N_4593,N_4496);
and U8776 (N_8776,N_4026,N_6068);
nor U8777 (N_8777,N_5690,N_3215);
and U8778 (N_8778,N_4551,N_4478);
and U8779 (N_8779,N_5467,N_5984);
or U8780 (N_8780,N_3806,N_6051);
xor U8781 (N_8781,N_4918,N_3160);
nor U8782 (N_8782,N_5448,N_4496);
or U8783 (N_8783,N_6220,N_3593);
or U8784 (N_8784,N_4508,N_4454);
and U8785 (N_8785,N_4661,N_6247);
xnor U8786 (N_8786,N_4851,N_4842);
or U8787 (N_8787,N_4015,N_6111);
nor U8788 (N_8788,N_3355,N_5081);
nor U8789 (N_8789,N_5485,N_4927);
nand U8790 (N_8790,N_5300,N_5315);
nor U8791 (N_8791,N_5702,N_5259);
or U8792 (N_8792,N_5434,N_4212);
nand U8793 (N_8793,N_3693,N_5536);
nand U8794 (N_8794,N_5360,N_3149);
nor U8795 (N_8795,N_4254,N_3858);
and U8796 (N_8796,N_4004,N_3973);
nand U8797 (N_8797,N_5494,N_4578);
nand U8798 (N_8798,N_4676,N_4054);
or U8799 (N_8799,N_4292,N_4824);
nor U8800 (N_8800,N_5922,N_3259);
and U8801 (N_8801,N_4700,N_3626);
and U8802 (N_8802,N_4447,N_5594);
nor U8803 (N_8803,N_5163,N_5981);
nand U8804 (N_8804,N_3982,N_4136);
nor U8805 (N_8805,N_4731,N_4831);
nor U8806 (N_8806,N_4126,N_3964);
nor U8807 (N_8807,N_4004,N_3839);
nand U8808 (N_8808,N_4052,N_6007);
nor U8809 (N_8809,N_3231,N_3191);
nand U8810 (N_8810,N_4231,N_3840);
nor U8811 (N_8811,N_6007,N_6197);
and U8812 (N_8812,N_5790,N_5967);
or U8813 (N_8813,N_5305,N_4191);
nor U8814 (N_8814,N_5362,N_5313);
and U8815 (N_8815,N_3750,N_3986);
nor U8816 (N_8816,N_3135,N_6019);
nand U8817 (N_8817,N_3294,N_4437);
or U8818 (N_8818,N_5860,N_6057);
nor U8819 (N_8819,N_4438,N_3853);
nand U8820 (N_8820,N_4243,N_5111);
xnor U8821 (N_8821,N_4356,N_4317);
nor U8822 (N_8822,N_3515,N_3708);
and U8823 (N_8823,N_5617,N_4294);
nor U8824 (N_8824,N_3474,N_5006);
and U8825 (N_8825,N_3161,N_3711);
or U8826 (N_8826,N_3196,N_4949);
nand U8827 (N_8827,N_5698,N_4606);
xnor U8828 (N_8828,N_3482,N_3219);
nor U8829 (N_8829,N_5251,N_3362);
nand U8830 (N_8830,N_3609,N_3182);
nand U8831 (N_8831,N_6102,N_3381);
nand U8832 (N_8832,N_4271,N_4076);
or U8833 (N_8833,N_5037,N_5451);
nor U8834 (N_8834,N_4596,N_5824);
and U8835 (N_8835,N_4696,N_5376);
nand U8836 (N_8836,N_4629,N_6035);
and U8837 (N_8837,N_3158,N_5834);
nand U8838 (N_8838,N_3578,N_4072);
or U8839 (N_8839,N_4715,N_6041);
nand U8840 (N_8840,N_5487,N_4441);
nor U8841 (N_8841,N_3986,N_4781);
nor U8842 (N_8842,N_4049,N_5039);
nor U8843 (N_8843,N_3452,N_3611);
nor U8844 (N_8844,N_4740,N_4176);
xnor U8845 (N_8845,N_5944,N_5257);
or U8846 (N_8846,N_4112,N_3360);
nand U8847 (N_8847,N_5909,N_5485);
and U8848 (N_8848,N_4171,N_4995);
nor U8849 (N_8849,N_3919,N_4999);
nor U8850 (N_8850,N_5920,N_4130);
nor U8851 (N_8851,N_3806,N_5165);
and U8852 (N_8852,N_5386,N_3333);
or U8853 (N_8853,N_5961,N_3503);
nor U8854 (N_8854,N_5700,N_5140);
nor U8855 (N_8855,N_5431,N_4210);
nor U8856 (N_8856,N_5370,N_5019);
nor U8857 (N_8857,N_5506,N_4790);
nor U8858 (N_8858,N_3447,N_5869);
nand U8859 (N_8859,N_5822,N_5532);
or U8860 (N_8860,N_4581,N_5118);
nand U8861 (N_8861,N_3791,N_5251);
nand U8862 (N_8862,N_3574,N_3825);
nand U8863 (N_8863,N_4091,N_5168);
or U8864 (N_8864,N_4714,N_5504);
xnor U8865 (N_8865,N_5154,N_4324);
xor U8866 (N_8866,N_4566,N_5362);
or U8867 (N_8867,N_5732,N_5428);
nand U8868 (N_8868,N_3925,N_6195);
and U8869 (N_8869,N_4767,N_5791);
and U8870 (N_8870,N_5590,N_3868);
nand U8871 (N_8871,N_3223,N_5878);
and U8872 (N_8872,N_5341,N_4024);
xnor U8873 (N_8873,N_3186,N_3541);
nand U8874 (N_8874,N_5815,N_4486);
nor U8875 (N_8875,N_5883,N_3909);
or U8876 (N_8876,N_4927,N_4282);
and U8877 (N_8877,N_4753,N_4933);
and U8878 (N_8878,N_4499,N_5854);
or U8879 (N_8879,N_3477,N_4363);
nand U8880 (N_8880,N_5335,N_3825);
or U8881 (N_8881,N_4392,N_4985);
nor U8882 (N_8882,N_3456,N_5579);
nand U8883 (N_8883,N_4309,N_3995);
and U8884 (N_8884,N_4306,N_5521);
or U8885 (N_8885,N_3427,N_4803);
nand U8886 (N_8886,N_4822,N_3903);
nor U8887 (N_8887,N_4777,N_6158);
and U8888 (N_8888,N_5573,N_5735);
or U8889 (N_8889,N_4202,N_3379);
and U8890 (N_8890,N_4903,N_5600);
or U8891 (N_8891,N_5013,N_4365);
or U8892 (N_8892,N_4149,N_3894);
and U8893 (N_8893,N_4005,N_6004);
and U8894 (N_8894,N_3605,N_6166);
or U8895 (N_8895,N_4344,N_3458);
and U8896 (N_8896,N_5215,N_3801);
nand U8897 (N_8897,N_4916,N_5194);
nand U8898 (N_8898,N_4439,N_3171);
nand U8899 (N_8899,N_5383,N_3969);
xor U8900 (N_8900,N_4339,N_5244);
or U8901 (N_8901,N_5938,N_4847);
or U8902 (N_8902,N_6009,N_5227);
nand U8903 (N_8903,N_5975,N_4224);
and U8904 (N_8904,N_4925,N_5709);
or U8905 (N_8905,N_6139,N_4013);
or U8906 (N_8906,N_3466,N_3594);
or U8907 (N_8907,N_6134,N_6002);
or U8908 (N_8908,N_5768,N_3194);
xnor U8909 (N_8909,N_4847,N_4802);
nand U8910 (N_8910,N_4235,N_5342);
or U8911 (N_8911,N_6049,N_3264);
xnor U8912 (N_8912,N_4030,N_6177);
xor U8913 (N_8913,N_3634,N_3479);
and U8914 (N_8914,N_3823,N_5703);
nand U8915 (N_8915,N_4792,N_3613);
nand U8916 (N_8916,N_6037,N_6016);
nor U8917 (N_8917,N_5171,N_3593);
nor U8918 (N_8918,N_4315,N_5680);
and U8919 (N_8919,N_5426,N_4262);
or U8920 (N_8920,N_3206,N_4913);
nor U8921 (N_8921,N_4638,N_3752);
or U8922 (N_8922,N_4330,N_4767);
and U8923 (N_8923,N_6235,N_5468);
nor U8924 (N_8924,N_4963,N_4242);
nand U8925 (N_8925,N_4740,N_3548);
or U8926 (N_8926,N_4173,N_5681);
or U8927 (N_8927,N_5781,N_5512);
and U8928 (N_8928,N_5191,N_4892);
nor U8929 (N_8929,N_5780,N_5621);
nor U8930 (N_8930,N_4916,N_4392);
nand U8931 (N_8931,N_5367,N_3812);
nand U8932 (N_8932,N_4386,N_4620);
and U8933 (N_8933,N_5320,N_5993);
or U8934 (N_8934,N_3573,N_3138);
nor U8935 (N_8935,N_4489,N_4693);
and U8936 (N_8936,N_5795,N_5466);
nand U8937 (N_8937,N_4759,N_5825);
nor U8938 (N_8938,N_3795,N_4238);
xnor U8939 (N_8939,N_4498,N_5381);
and U8940 (N_8940,N_5767,N_3442);
nand U8941 (N_8941,N_6156,N_4616);
nand U8942 (N_8942,N_3914,N_5907);
nand U8943 (N_8943,N_6187,N_3392);
and U8944 (N_8944,N_4085,N_5716);
nand U8945 (N_8945,N_4024,N_4628);
or U8946 (N_8946,N_3853,N_6052);
or U8947 (N_8947,N_4565,N_5106);
nand U8948 (N_8948,N_3586,N_3286);
and U8949 (N_8949,N_6051,N_4016);
nand U8950 (N_8950,N_5171,N_3126);
nor U8951 (N_8951,N_5015,N_4463);
nor U8952 (N_8952,N_4546,N_4031);
or U8953 (N_8953,N_5884,N_5998);
and U8954 (N_8954,N_3358,N_5405);
xnor U8955 (N_8955,N_3906,N_5758);
or U8956 (N_8956,N_3829,N_3608);
and U8957 (N_8957,N_4392,N_5273);
nor U8958 (N_8958,N_5718,N_5532);
xor U8959 (N_8959,N_3202,N_4425);
and U8960 (N_8960,N_5626,N_3218);
nor U8961 (N_8961,N_3795,N_5377);
or U8962 (N_8962,N_5336,N_4724);
or U8963 (N_8963,N_5331,N_3551);
nand U8964 (N_8964,N_5235,N_3956);
nand U8965 (N_8965,N_5982,N_4105);
nand U8966 (N_8966,N_5243,N_5412);
and U8967 (N_8967,N_4994,N_3365);
xor U8968 (N_8968,N_6152,N_3556);
and U8969 (N_8969,N_4320,N_5294);
or U8970 (N_8970,N_5496,N_3916);
nor U8971 (N_8971,N_5582,N_5075);
nand U8972 (N_8972,N_5375,N_4878);
and U8973 (N_8973,N_5074,N_5022);
or U8974 (N_8974,N_5086,N_4100);
xor U8975 (N_8975,N_5470,N_5780);
nand U8976 (N_8976,N_5021,N_4457);
nor U8977 (N_8977,N_4595,N_5896);
nand U8978 (N_8978,N_6027,N_5909);
xnor U8979 (N_8979,N_5074,N_4006);
and U8980 (N_8980,N_3928,N_3743);
or U8981 (N_8981,N_4527,N_5977);
nor U8982 (N_8982,N_3989,N_3407);
nor U8983 (N_8983,N_3946,N_3372);
and U8984 (N_8984,N_4356,N_3297);
or U8985 (N_8985,N_5758,N_5565);
or U8986 (N_8986,N_6245,N_3997);
nor U8987 (N_8987,N_5097,N_4366);
nor U8988 (N_8988,N_3463,N_3129);
nor U8989 (N_8989,N_4585,N_3941);
and U8990 (N_8990,N_5779,N_5261);
and U8991 (N_8991,N_3501,N_5240);
and U8992 (N_8992,N_4916,N_4470);
or U8993 (N_8993,N_3678,N_3333);
nand U8994 (N_8994,N_3672,N_5184);
and U8995 (N_8995,N_5422,N_3539);
and U8996 (N_8996,N_5171,N_3236);
and U8997 (N_8997,N_5517,N_5765);
xor U8998 (N_8998,N_5503,N_5696);
or U8999 (N_8999,N_4349,N_6180);
nand U9000 (N_9000,N_4074,N_3465);
nor U9001 (N_9001,N_5383,N_5562);
or U9002 (N_9002,N_5314,N_3343);
or U9003 (N_9003,N_3707,N_5391);
nor U9004 (N_9004,N_4985,N_3750);
and U9005 (N_9005,N_3360,N_4721);
or U9006 (N_9006,N_4532,N_4435);
and U9007 (N_9007,N_3485,N_4399);
and U9008 (N_9008,N_5790,N_3162);
xor U9009 (N_9009,N_4986,N_3216);
and U9010 (N_9010,N_4362,N_3678);
or U9011 (N_9011,N_5134,N_5279);
and U9012 (N_9012,N_5063,N_4087);
nand U9013 (N_9013,N_3288,N_4516);
or U9014 (N_9014,N_4845,N_5717);
and U9015 (N_9015,N_3684,N_4167);
xor U9016 (N_9016,N_3882,N_3460);
nand U9017 (N_9017,N_3901,N_5723);
or U9018 (N_9018,N_5883,N_3609);
and U9019 (N_9019,N_4689,N_4057);
nand U9020 (N_9020,N_6136,N_5188);
or U9021 (N_9021,N_3660,N_3694);
or U9022 (N_9022,N_4445,N_5604);
or U9023 (N_9023,N_5743,N_3913);
nand U9024 (N_9024,N_5174,N_5554);
or U9025 (N_9025,N_3924,N_4414);
nor U9026 (N_9026,N_3773,N_5761);
or U9027 (N_9027,N_3822,N_3971);
or U9028 (N_9028,N_6084,N_3498);
and U9029 (N_9029,N_4150,N_3683);
nand U9030 (N_9030,N_4444,N_4087);
or U9031 (N_9031,N_5083,N_6233);
nand U9032 (N_9032,N_3312,N_4652);
nand U9033 (N_9033,N_3582,N_5011);
nand U9034 (N_9034,N_3438,N_6052);
xor U9035 (N_9035,N_5177,N_5212);
or U9036 (N_9036,N_5140,N_3171);
nor U9037 (N_9037,N_4295,N_3297);
and U9038 (N_9038,N_5228,N_4259);
and U9039 (N_9039,N_5972,N_5749);
xnor U9040 (N_9040,N_4768,N_5454);
nand U9041 (N_9041,N_4375,N_3926);
or U9042 (N_9042,N_6187,N_4183);
nor U9043 (N_9043,N_4798,N_5729);
nor U9044 (N_9044,N_5278,N_6173);
nor U9045 (N_9045,N_4388,N_4699);
nand U9046 (N_9046,N_5688,N_5819);
or U9047 (N_9047,N_5276,N_6182);
nand U9048 (N_9048,N_5894,N_5438);
or U9049 (N_9049,N_3483,N_4980);
or U9050 (N_9050,N_5617,N_3230);
nor U9051 (N_9051,N_3942,N_3229);
or U9052 (N_9052,N_5189,N_6186);
nor U9053 (N_9053,N_4743,N_5388);
and U9054 (N_9054,N_3981,N_4952);
or U9055 (N_9055,N_4450,N_5792);
and U9056 (N_9056,N_3535,N_5862);
nor U9057 (N_9057,N_3994,N_3195);
or U9058 (N_9058,N_4037,N_4927);
nor U9059 (N_9059,N_3780,N_4926);
nor U9060 (N_9060,N_5350,N_4625);
nor U9061 (N_9061,N_4067,N_4026);
xor U9062 (N_9062,N_3978,N_5739);
or U9063 (N_9063,N_5696,N_3691);
or U9064 (N_9064,N_6111,N_3737);
or U9065 (N_9065,N_3207,N_5484);
nand U9066 (N_9066,N_5244,N_5313);
and U9067 (N_9067,N_6115,N_5426);
nand U9068 (N_9068,N_5058,N_4009);
nand U9069 (N_9069,N_6014,N_5817);
and U9070 (N_9070,N_5037,N_4517);
or U9071 (N_9071,N_5778,N_3745);
or U9072 (N_9072,N_6000,N_4266);
nor U9073 (N_9073,N_5199,N_5698);
nor U9074 (N_9074,N_3579,N_3652);
or U9075 (N_9075,N_5729,N_5163);
and U9076 (N_9076,N_4184,N_3872);
nand U9077 (N_9077,N_5227,N_4521);
and U9078 (N_9078,N_5452,N_4285);
and U9079 (N_9079,N_5035,N_3899);
and U9080 (N_9080,N_5240,N_4097);
or U9081 (N_9081,N_6195,N_3334);
xnor U9082 (N_9082,N_5668,N_5182);
and U9083 (N_9083,N_4602,N_5385);
nor U9084 (N_9084,N_4655,N_4364);
nand U9085 (N_9085,N_3961,N_4803);
nand U9086 (N_9086,N_3410,N_3499);
or U9087 (N_9087,N_5651,N_5172);
xor U9088 (N_9088,N_3804,N_5054);
or U9089 (N_9089,N_4369,N_4986);
nor U9090 (N_9090,N_5356,N_3689);
or U9091 (N_9091,N_3945,N_3528);
or U9092 (N_9092,N_5008,N_3592);
or U9093 (N_9093,N_5129,N_4731);
xor U9094 (N_9094,N_6178,N_3216);
and U9095 (N_9095,N_4684,N_3646);
and U9096 (N_9096,N_4376,N_4195);
and U9097 (N_9097,N_3399,N_5598);
and U9098 (N_9098,N_4615,N_4557);
and U9099 (N_9099,N_5879,N_5127);
and U9100 (N_9100,N_5051,N_5027);
and U9101 (N_9101,N_5687,N_6181);
and U9102 (N_9102,N_4608,N_4078);
xnor U9103 (N_9103,N_3220,N_3473);
nand U9104 (N_9104,N_4213,N_3191);
nor U9105 (N_9105,N_5447,N_5756);
nand U9106 (N_9106,N_5639,N_5812);
nand U9107 (N_9107,N_4294,N_4647);
or U9108 (N_9108,N_5035,N_4629);
xnor U9109 (N_9109,N_4799,N_5925);
nor U9110 (N_9110,N_4340,N_3619);
or U9111 (N_9111,N_3706,N_5226);
and U9112 (N_9112,N_5571,N_5406);
nand U9113 (N_9113,N_5586,N_5191);
nand U9114 (N_9114,N_5531,N_5953);
and U9115 (N_9115,N_3893,N_4617);
and U9116 (N_9116,N_4261,N_4376);
or U9117 (N_9117,N_3834,N_5744);
nand U9118 (N_9118,N_4277,N_4429);
nor U9119 (N_9119,N_4586,N_4980);
or U9120 (N_9120,N_3466,N_3418);
or U9121 (N_9121,N_3444,N_3503);
and U9122 (N_9122,N_5805,N_6138);
nor U9123 (N_9123,N_4000,N_5963);
or U9124 (N_9124,N_4478,N_6177);
and U9125 (N_9125,N_4440,N_4074);
nand U9126 (N_9126,N_3378,N_3897);
nor U9127 (N_9127,N_5668,N_5629);
and U9128 (N_9128,N_3137,N_3828);
or U9129 (N_9129,N_3130,N_4691);
and U9130 (N_9130,N_3892,N_5460);
nand U9131 (N_9131,N_4793,N_4636);
nor U9132 (N_9132,N_4776,N_3955);
nor U9133 (N_9133,N_5632,N_4682);
nor U9134 (N_9134,N_6204,N_3247);
nor U9135 (N_9135,N_4441,N_6066);
or U9136 (N_9136,N_4748,N_4160);
xnor U9137 (N_9137,N_3358,N_4415);
and U9138 (N_9138,N_5535,N_4599);
nor U9139 (N_9139,N_5534,N_3383);
nor U9140 (N_9140,N_3559,N_5053);
nand U9141 (N_9141,N_3537,N_5225);
nand U9142 (N_9142,N_3977,N_3467);
and U9143 (N_9143,N_4004,N_4781);
or U9144 (N_9144,N_3804,N_4403);
and U9145 (N_9145,N_4507,N_3889);
or U9146 (N_9146,N_3225,N_4738);
and U9147 (N_9147,N_4385,N_4160);
nand U9148 (N_9148,N_6137,N_5219);
and U9149 (N_9149,N_4561,N_5530);
nor U9150 (N_9150,N_4948,N_3339);
nor U9151 (N_9151,N_4118,N_3653);
nand U9152 (N_9152,N_3147,N_5163);
or U9153 (N_9153,N_3620,N_4952);
and U9154 (N_9154,N_4963,N_5244);
nand U9155 (N_9155,N_3749,N_5733);
and U9156 (N_9156,N_5072,N_5557);
or U9157 (N_9157,N_5459,N_6246);
and U9158 (N_9158,N_4374,N_5520);
and U9159 (N_9159,N_5540,N_4924);
nor U9160 (N_9160,N_5445,N_4401);
nand U9161 (N_9161,N_3668,N_3246);
nor U9162 (N_9162,N_3911,N_3311);
and U9163 (N_9163,N_3403,N_5593);
and U9164 (N_9164,N_5389,N_5073);
or U9165 (N_9165,N_3178,N_3412);
and U9166 (N_9166,N_4433,N_3371);
nor U9167 (N_9167,N_3288,N_5937);
or U9168 (N_9168,N_5636,N_6116);
xor U9169 (N_9169,N_5778,N_4269);
nor U9170 (N_9170,N_3697,N_3216);
and U9171 (N_9171,N_4760,N_4240);
xor U9172 (N_9172,N_4549,N_3636);
or U9173 (N_9173,N_5207,N_4506);
and U9174 (N_9174,N_6106,N_4550);
xnor U9175 (N_9175,N_4605,N_3781);
and U9176 (N_9176,N_4474,N_4955);
and U9177 (N_9177,N_3218,N_5535);
nor U9178 (N_9178,N_6150,N_5477);
and U9179 (N_9179,N_4292,N_6046);
nand U9180 (N_9180,N_4022,N_5277);
nor U9181 (N_9181,N_6247,N_6055);
and U9182 (N_9182,N_3615,N_3286);
and U9183 (N_9183,N_5223,N_6248);
xor U9184 (N_9184,N_5215,N_3381);
nor U9185 (N_9185,N_5534,N_5642);
nor U9186 (N_9186,N_3470,N_6088);
xor U9187 (N_9187,N_5703,N_5202);
nand U9188 (N_9188,N_6042,N_3321);
nand U9189 (N_9189,N_5299,N_4559);
and U9190 (N_9190,N_3557,N_3309);
xor U9191 (N_9191,N_3476,N_4817);
nor U9192 (N_9192,N_3303,N_6105);
or U9193 (N_9193,N_4650,N_6162);
nor U9194 (N_9194,N_6195,N_5052);
or U9195 (N_9195,N_5359,N_3888);
and U9196 (N_9196,N_4512,N_4911);
or U9197 (N_9197,N_5157,N_5191);
nand U9198 (N_9198,N_4978,N_5374);
or U9199 (N_9199,N_3281,N_3269);
and U9200 (N_9200,N_5133,N_5154);
and U9201 (N_9201,N_4847,N_4116);
or U9202 (N_9202,N_4354,N_3905);
xnor U9203 (N_9203,N_5248,N_5182);
and U9204 (N_9204,N_4376,N_4486);
and U9205 (N_9205,N_5843,N_5617);
nand U9206 (N_9206,N_5963,N_3271);
and U9207 (N_9207,N_3452,N_4842);
nor U9208 (N_9208,N_4081,N_3787);
nor U9209 (N_9209,N_6079,N_4510);
and U9210 (N_9210,N_3908,N_3481);
and U9211 (N_9211,N_4768,N_3285);
nor U9212 (N_9212,N_4444,N_5656);
and U9213 (N_9213,N_3887,N_3131);
nand U9214 (N_9214,N_3936,N_4016);
or U9215 (N_9215,N_5810,N_5048);
xnor U9216 (N_9216,N_4498,N_5450);
and U9217 (N_9217,N_3397,N_3721);
nand U9218 (N_9218,N_3902,N_3626);
and U9219 (N_9219,N_5333,N_3726);
or U9220 (N_9220,N_3884,N_5043);
nand U9221 (N_9221,N_3137,N_5214);
nor U9222 (N_9222,N_3990,N_5118);
nand U9223 (N_9223,N_5358,N_4402);
nand U9224 (N_9224,N_3245,N_5078);
xor U9225 (N_9225,N_5317,N_4669);
nor U9226 (N_9226,N_3561,N_3993);
nor U9227 (N_9227,N_3239,N_5850);
and U9228 (N_9228,N_5298,N_3921);
nor U9229 (N_9229,N_3517,N_3385);
xor U9230 (N_9230,N_5851,N_3888);
nor U9231 (N_9231,N_4408,N_3655);
and U9232 (N_9232,N_3210,N_6102);
or U9233 (N_9233,N_3940,N_3303);
xor U9234 (N_9234,N_3574,N_3813);
and U9235 (N_9235,N_4712,N_5697);
nand U9236 (N_9236,N_4785,N_4534);
or U9237 (N_9237,N_4165,N_3396);
nor U9238 (N_9238,N_5554,N_4355);
and U9239 (N_9239,N_4767,N_3756);
xor U9240 (N_9240,N_3903,N_5259);
or U9241 (N_9241,N_6106,N_3881);
nor U9242 (N_9242,N_5604,N_5887);
or U9243 (N_9243,N_5395,N_5579);
nor U9244 (N_9244,N_5980,N_4336);
xnor U9245 (N_9245,N_4602,N_3850);
and U9246 (N_9246,N_4684,N_3787);
or U9247 (N_9247,N_5767,N_5577);
nor U9248 (N_9248,N_6069,N_4941);
and U9249 (N_9249,N_5252,N_3320);
nand U9250 (N_9250,N_5592,N_5489);
and U9251 (N_9251,N_4764,N_4605);
and U9252 (N_9252,N_5369,N_3512);
nand U9253 (N_9253,N_4292,N_3412);
nor U9254 (N_9254,N_5140,N_3135);
xor U9255 (N_9255,N_5090,N_5141);
and U9256 (N_9256,N_5887,N_3489);
xor U9257 (N_9257,N_4493,N_3637);
nor U9258 (N_9258,N_6051,N_5153);
and U9259 (N_9259,N_3436,N_5363);
nor U9260 (N_9260,N_5133,N_4717);
or U9261 (N_9261,N_4105,N_5245);
nor U9262 (N_9262,N_4761,N_4581);
nor U9263 (N_9263,N_3527,N_3209);
and U9264 (N_9264,N_4410,N_3652);
or U9265 (N_9265,N_4211,N_4799);
and U9266 (N_9266,N_4915,N_4632);
and U9267 (N_9267,N_4664,N_6032);
nand U9268 (N_9268,N_6007,N_4851);
nor U9269 (N_9269,N_5029,N_4176);
nand U9270 (N_9270,N_6085,N_3949);
nand U9271 (N_9271,N_5875,N_5438);
nor U9272 (N_9272,N_4690,N_3189);
nand U9273 (N_9273,N_5852,N_4643);
nand U9274 (N_9274,N_3676,N_3552);
and U9275 (N_9275,N_5686,N_4603);
nor U9276 (N_9276,N_6139,N_4498);
nor U9277 (N_9277,N_5756,N_4722);
nand U9278 (N_9278,N_4824,N_5158);
nand U9279 (N_9279,N_5059,N_4479);
and U9280 (N_9280,N_5409,N_5025);
or U9281 (N_9281,N_4941,N_3256);
nor U9282 (N_9282,N_6178,N_6203);
nand U9283 (N_9283,N_4697,N_6201);
and U9284 (N_9284,N_3776,N_4131);
nor U9285 (N_9285,N_3178,N_5898);
and U9286 (N_9286,N_5491,N_4753);
nor U9287 (N_9287,N_3607,N_4643);
or U9288 (N_9288,N_4975,N_4913);
nand U9289 (N_9289,N_3323,N_3747);
and U9290 (N_9290,N_3265,N_4347);
and U9291 (N_9291,N_4385,N_4675);
nor U9292 (N_9292,N_3872,N_3575);
nand U9293 (N_9293,N_3942,N_4773);
or U9294 (N_9294,N_3930,N_4342);
and U9295 (N_9295,N_4785,N_3541);
nor U9296 (N_9296,N_3201,N_4192);
nor U9297 (N_9297,N_4856,N_4424);
nor U9298 (N_9298,N_4288,N_3929);
or U9299 (N_9299,N_4710,N_5562);
nand U9300 (N_9300,N_4413,N_4427);
or U9301 (N_9301,N_4258,N_3637);
nand U9302 (N_9302,N_4114,N_5030);
and U9303 (N_9303,N_3612,N_3768);
nand U9304 (N_9304,N_5732,N_3419);
nand U9305 (N_9305,N_5377,N_5527);
nand U9306 (N_9306,N_3969,N_4394);
xor U9307 (N_9307,N_4045,N_4025);
nand U9308 (N_9308,N_3853,N_5245);
or U9309 (N_9309,N_5637,N_5500);
and U9310 (N_9310,N_5632,N_6042);
nor U9311 (N_9311,N_4095,N_3403);
and U9312 (N_9312,N_4521,N_5284);
or U9313 (N_9313,N_4508,N_3539);
xor U9314 (N_9314,N_3470,N_5416);
nor U9315 (N_9315,N_3337,N_4996);
nor U9316 (N_9316,N_6107,N_3872);
and U9317 (N_9317,N_3228,N_3462);
and U9318 (N_9318,N_4537,N_5031);
nand U9319 (N_9319,N_6166,N_4662);
and U9320 (N_9320,N_4514,N_4131);
nand U9321 (N_9321,N_4919,N_4589);
or U9322 (N_9322,N_4614,N_3628);
or U9323 (N_9323,N_5645,N_3612);
nand U9324 (N_9324,N_3286,N_3160);
nor U9325 (N_9325,N_4886,N_4756);
nor U9326 (N_9326,N_4729,N_5184);
and U9327 (N_9327,N_4101,N_4193);
nand U9328 (N_9328,N_5011,N_5843);
or U9329 (N_9329,N_4041,N_5028);
nor U9330 (N_9330,N_3452,N_4457);
nor U9331 (N_9331,N_3896,N_4430);
nand U9332 (N_9332,N_4706,N_5901);
nand U9333 (N_9333,N_4387,N_3613);
and U9334 (N_9334,N_6154,N_3650);
nand U9335 (N_9335,N_4867,N_3416);
or U9336 (N_9336,N_5987,N_5928);
nor U9337 (N_9337,N_3661,N_6174);
or U9338 (N_9338,N_3404,N_4059);
nor U9339 (N_9339,N_5681,N_4920);
nor U9340 (N_9340,N_3514,N_4516);
or U9341 (N_9341,N_4310,N_3556);
xor U9342 (N_9342,N_4602,N_4113);
and U9343 (N_9343,N_5254,N_3698);
nand U9344 (N_9344,N_4800,N_3223);
nand U9345 (N_9345,N_5445,N_5296);
nand U9346 (N_9346,N_5518,N_5668);
and U9347 (N_9347,N_5137,N_3414);
xnor U9348 (N_9348,N_6034,N_4162);
nor U9349 (N_9349,N_4957,N_5472);
nand U9350 (N_9350,N_4313,N_5718);
nor U9351 (N_9351,N_4354,N_4353);
nor U9352 (N_9352,N_4876,N_4302);
xnor U9353 (N_9353,N_4794,N_3260);
or U9354 (N_9354,N_5433,N_4974);
xor U9355 (N_9355,N_3435,N_4273);
nand U9356 (N_9356,N_5186,N_3352);
xnor U9357 (N_9357,N_5911,N_5144);
nand U9358 (N_9358,N_6004,N_4609);
or U9359 (N_9359,N_3827,N_3627);
or U9360 (N_9360,N_6171,N_3761);
or U9361 (N_9361,N_3813,N_5904);
and U9362 (N_9362,N_5383,N_5685);
nor U9363 (N_9363,N_3289,N_5968);
nor U9364 (N_9364,N_4439,N_5895);
and U9365 (N_9365,N_4903,N_3355);
and U9366 (N_9366,N_4518,N_5501);
or U9367 (N_9367,N_5490,N_3987);
and U9368 (N_9368,N_3575,N_4212);
nor U9369 (N_9369,N_5757,N_3958);
nand U9370 (N_9370,N_4870,N_5858);
and U9371 (N_9371,N_4578,N_3526);
or U9372 (N_9372,N_4286,N_4837);
and U9373 (N_9373,N_4237,N_4244);
nand U9374 (N_9374,N_6099,N_6224);
or U9375 (N_9375,N_8457,N_7555);
or U9376 (N_9376,N_8654,N_8005);
or U9377 (N_9377,N_6333,N_6477);
xor U9378 (N_9378,N_7148,N_6361);
nor U9379 (N_9379,N_7389,N_7858);
nor U9380 (N_9380,N_8581,N_8766);
nor U9381 (N_9381,N_7069,N_8161);
or U9382 (N_9382,N_9155,N_7430);
nor U9383 (N_9383,N_7963,N_8349);
xnor U9384 (N_9384,N_8355,N_8783);
nand U9385 (N_9385,N_6984,N_8399);
and U9386 (N_9386,N_8029,N_7848);
nand U9387 (N_9387,N_7526,N_7094);
nor U9388 (N_9388,N_9073,N_7396);
nand U9389 (N_9389,N_8118,N_6359);
and U9390 (N_9390,N_7059,N_6393);
nor U9391 (N_9391,N_8992,N_7382);
nand U9392 (N_9392,N_7826,N_6639);
or U9393 (N_9393,N_8056,N_9242);
nand U9394 (N_9394,N_6924,N_7949);
or U9395 (N_9395,N_7229,N_8590);
and U9396 (N_9396,N_6731,N_6939);
nand U9397 (N_9397,N_8921,N_6257);
xor U9398 (N_9398,N_6672,N_8008);
nor U9399 (N_9399,N_7202,N_6816);
nand U9400 (N_9400,N_8742,N_8153);
nor U9401 (N_9401,N_6349,N_6325);
nor U9402 (N_9402,N_7782,N_6552);
nor U9403 (N_9403,N_8690,N_7985);
or U9404 (N_9404,N_8347,N_8828);
nand U9405 (N_9405,N_7923,N_9257);
nand U9406 (N_9406,N_8064,N_8787);
xor U9407 (N_9407,N_9185,N_8326);
nand U9408 (N_9408,N_7952,N_7019);
and U9409 (N_9409,N_8754,N_7790);
nor U9410 (N_9410,N_9071,N_6296);
xor U9411 (N_9411,N_6466,N_8936);
nor U9412 (N_9412,N_7536,N_9163);
or U9413 (N_9413,N_8557,N_8694);
or U9414 (N_9414,N_7224,N_7279);
nand U9415 (N_9415,N_7958,N_6551);
nor U9416 (N_9416,N_6389,N_7348);
nand U9417 (N_9417,N_7061,N_7617);
nand U9418 (N_9418,N_6809,N_8167);
nor U9419 (N_9419,N_8786,N_7143);
nor U9420 (N_9420,N_7186,N_8856);
nand U9421 (N_9421,N_8362,N_6434);
or U9422 (N_9422,N_6928,N_6829);
and U9423 (N_9423,N_9264,N_7713);
xnor U9424 (N_9424,N_9332,N_9021);
nor U9425 (N_9425,N_9007,N_7503);
or U9426 (N_9426,N_8941,N_6274);
nor U9427 (N_9427,N_8224,N_8375);
nand U9428 (N_9428,N_7475,N_9097);
or U9429 (N_9429,N_6632,N_9126);
and U9430 (N_9430,N_8511,N_6755);
nand U9431 (N_9431,N_8726,N_8894);
and U9432 (N_9432,N_8658,N_8746);
xnor U9433 (N_9433,N_7614,N_6454);
nor U9434 (N_9434,N_8048,N_8427);
nand U9435 (N_9435,N_7932,N_9114);
xnor U9436 (N_9436,N_8981,N_6541);
xnor U9437 (N_9437,N_8236,N_8885);
xnor U9438 (N_9438,N_8736,N_7838);
or U9439 (N_9439,N_6481,N_6375);
nor U9440 (N_9440,N_7683,N_9212);
xnor U9441 (N_9441,N_6726,N_9273);
xor U9442 (N_9442,N_7383,N_9194);
xor U9443 (N_9443,N_6743,N_6366);
nand U9444 (N_9444,N_9127,N_8071);
xor U9445 (N_9445,N_6427,N_9280);
nand U9446 (N_9446,N_6700,N_8961);
nand U9447 (N_9447,N_7337,N_8334);
nand U9448 (N_9448,N_7127,N_6812);
nand U9449 (N_9449,N_8335,N_7048);
nand U9450 (N_9450,N_7257,N_6699);
xnor U9451 (N_9451,N_6528,N_8451);
or U9452 (N_9452,N_8827,N_7737);
or U9453 (N_9453,N_8378,N_6478);
or U9454 (N_9454,N_7761,N_8144);
nor U9455 (N_9455,N_7471,N_7386);
and U9456 (N_9456,N_8262,N_6555);
or U9457 (N_9457,N_6566,N_6640);
nand U9458 (N_9458,N_8614,N_7110);
nor U9459 (N_9459,N_8879,N_9096);
nand U9460 (N_9460,N_6857,N_6740);
and U9461 (N_9461,N_7271,N_8149);
nand U9462 (N_9462,N_8907,N_8088);
nor U9463 (N_9463,N_8040,N_8456);
and U9464 (N_9464,N_7969,N_6608);
and U9465 (N_9465,N_8893,N_8321);
nand U9466 (N_9466,N_7661,N_8779);
nor U9467 (N_9467,N_8434,N_9036);
nor U9468 (N_9468,N_8387,N_7083);
nor U9469 (N_9469,N_8127,N_8775);
nand U9470 (N_9470,N_8583,N_7693);
nor U9471 (N_9471,N_8390,N_7914);
or U9472 (N_9472,N_6383,N_8126);
and U9473 (N_9473,N_9301,N_6429);
and U9474 (N_9474,N_6446,N_8464);
nand U9475 (N_9475,N_7818,N_8668);
xnor U9476 (N_9476,N_9043,N_6706);
nor U9477 (N_9477,N_6490,N_9116);
or U9478 (N_9478,N_7209,N_6884);
xor U9479 (N_9479,N_7967,N_6817);
and U9480 (N_9480,N_7260,N_9058);
and U9481 (N_9481,N_7808,N_7018);
nand U9482 (N_9482,N_8429,N_8163);
and U9483 (N_9483,N_8183,N_8160);
or U9484 (N_9484,N_9230,N_8203);
nand U9485 (N_9485,N_9070,N_7068);
nand U9486 (N_9486,N_9341,N_7791);
xor U9487 (N_9487,N_6854,N_9140);
nor U9488 (N_9488,N_7884,N_7170);
and U9489 (N_9489,N_8195,N_9355);
xnor U9490 (N_9490,N_8274,N_6835);
or U9491 (N_9491,N_8579,N_9111);
or U9492 (N_9492,N_6431,N_7973);
or U9493 (N_9493,N_6694,N_8592);
or U9494 (N_9494,N_6858,N_6982);
nor U9495 (N_9495,N_6293,N_6402);
xnor U9496 (N_9496,N_7243,N_9170);
or U9497 (N_9497,N_9051,N_8510);
or U9498 (N_9498,N_6484,N_8926);
nor U9499 (N_9499,N_6515,N_7623);
nor U9500 (N_9500,N_9271,N_9227);
or U9501 (N_9501,N_8381,N_8312);
nor U9502 (N_9502,N_7219,N_8780);
nand U9503 (N_9503,N_8684,N_7165);
nand U9504 (N_9504,N_8763,N_8735);
nand U9505 (N_9505,N_6272,N_8415);
nor U9506 (N_9506,N_6677,N_8374);
and U9507 (N_9507,N_6533,N_8769);
or U9508 (N_9508,N_6258,N_8458);
nor U9509 (N_9509,N_8608,N_7947);
and U9510 (N_9510,N_7097,N_6462);
nand U9511 (N_9511,N_7040,N_8744);
and U9512 (N_9512,N_8878,N_7763);
nor U9513 (N_9513,N_8616,N_8728);
or U9514 (N_9514,N_6591,N_8793);
or U9515 (N_9515,N_6322,N_7917);
xnor U9516 (N_9516,N_8738,N_8343);
nor U9517 (N_9517,N_7065,N_9309);
and U9518 (N_9518,N_8634,N_7505);
or U9519 (N_9519,N_9358,N_9191);
nor U9520 (N_9520,N_6768,N_9059);
and U9521 (N_9521,N_6653,N_6885);
xnor U9522 (N_9522,N_8846,N_8512);
or U9523 (N_9523,N_8165,N_6949);
nor U9524 (N_9524,N_6705,N_7034);
nor U9525 (N_9525,N_8124,N_8317);
or U9526 (N_9526,N_8023,N_7485);
and U9527 (N_9527,N_7265,N_7298);
nand U9528 (N_9528,N_8782,N_8030);
nor U9529 (N_9529,N_6444,N_7760);
and U9530 (N_9530,N_9228,N_7753);
and U9531 (N_9531,N_6834,N_8376);
xnor U9532 (N_9532,N_8649,N_6983);
nor U9533 (N_9533,N_9158,N_8367);
and U9534 (N_9534,N_8546,N_7494);
nand U9535 (N_9535,N_9334,N_8778);
and U9536 (N_9536,N_7333,N_9243);
nor U9537 (N_9537,N_7128,N_7938);
and U9538 (N_9538,N_6331,N_8282);
xor U9539 (N_9539,N_6804,N_6849);
or U9540 (N_9540,N_7598,N_6558);
xor U9541 (N_9541,N_6752,N_7318);
and U9542 (N_9542,N_8709,N_8465);
nor U9543 (N_9543,N_7570,N_8364);
and U9544 (N_9544,N_7836,N_7664);
nor U9545 (N_9545,N_7984,N_6624);
nand U9546 (N_9546,N_9206,N_8000);
nor U9547 (N_9547,N_9148,N_6489);
nand U9548 (N_9548,N_6407,N_8553);
nand U9549 (N_9549,N_6588,N_6573);
nand U9550 (N_9550,N_8215,N_7246);
nand U9551 (N_9551,N_7255,N_6289);
or U9552 (N_9552,N_7465,N_8929);
xor U9553 (N_9553,N_6439,N_8604);
or U9554 (N_9554,N_8834,N_6832);
or U9555 (N_9555,N_7819,N_7795);
nor U9556 (N_9556,N_6364,N_7037);
or U9557 (N_9557,N_6259,N_6602);
nor U9558 (N_9558,N_7983,N_9052);
nand U9559 (N_9559,N_6674,N_8577);
nor U9560 (N_9560,N_9203,N_7785);
nor U9561 (N_9561,N_7904,N_8997);
and U9562 (N_9562,N_8815,N_9008);
nor U9563 (N_9563,N_8701,N_6783);
and U9564 (N_9564,N_7792,N_6722);
or U9565 (N_9565,N_8999,N_6998);
and U9566 (N_9566,N_6337,N_8586);
and U9567 (N_9567,N_8411,N_7381);
and U9568 (N_9568,N_6356,N_8666);
and U9569 (N_9569,N_6605,N_7432);
nor U9570 (N_9570,N_6719,N_9342);
and U9571 (N_9571,N_8756,N_6796);
or U9572 (N_9572,N_7253,N_9366);
nor U9573 (N_9573,N_7665,N_8781);
or U9574 (N_9574,N_6933,N_8663);
and U9575 (N_9575,N_8304,N_6791);
or U9576 (N_9576,N_8143,N_8811);
nand U9577 (N_9577,N_6955,N_7435);
nor U9578 (N_9578,N_9174,N_8619);
and U9579 (N_9579,N_8896,N_7770);
and U9580 (N_9580,N_7375,N_6584);
nand U9581 (N_9581,N_7748,N_6582);
or U9582 (N_9582,N_8864,N_9083);
nor U9583 (N_9583,N_8015,N_6670);
nor U9584 (N_9584,N_7950,N_7036);
or U9585 (N_9585,N_7953,N_7288);
nor U9586 (N_9586,N_7448,N_6920);
or U9587 (N_9587,N_7680,N_6600);
nand U9588 (N_9588,N_9207,N_9258);
nor U9589 (N_9589,N_6931,N_8814);
and U9590 (N_9590,N_7184,N_6307);
and U9591 (N_9591,N_8212,N_9069);
or U9592 (N_9592,N_6360,N_6543);
or U9593 (N_9593,N_7160,N_8870);
nand U9594 (N_9594,N_8301,N_8617);
xnor U9595 (N_9595,N_7613,N_6893);
nand U9596 (N_9596,N_6990,N_8093);
or U9597 (N_9597,N_6492,N_7362);
or U9598 (N_9598,N_7597,N_8682);
nand U9599 (N_9599,N_7408,N_7264);
nand U9600 (N_9600,N_7134,N_8631);
and U9601 (N_9601,N_6961,N_8998);
or U9602 (N_9602,N_7703,N_6897);
or U9603 (N_9603,N_6362,N_7580);
xor U9604 (N_9604,N_8958,N_7007);
nand U9605 (N_9605,N_8904,N_6286);
or U9606 (N_9606,N_9336,N_9161);
and U9607 (N_9607,N_6271,N_8774);
nand U9608 (N_9608,N_8110,N_8482);
or U9609 (N_9609,N_9371,N_8596);
and U9610 (N_9610,N_7433,N_8012);
or U9611 (N_9611,N_6787,N_7589);
and U9612 (N_9612,N_8141,N_8132);
nand U9613 (N_9613,N_6500,N_9218);
nor U9614 (N_9614,N_6280,N_7604);
and U9615 (N_9615,N_7093,N_8971);
nor U9616 (N_9616,N_8201,N_8761);
or U9617 (N_9617,N_8665,N_8582);
or U9618 (N_9618,N_8425,N_7565);
xnor U9619 (N_9619,N_7890,N_8611);
or U9620 (N_9620,N_7909,N_8599);
nand U9621 (N_9621,N_7974,N_8522);
xnor U9622 (N_9622,N_6807,N_8222);
nor U9623 (N_9623,N_6980,N_7210);
or U9624 (N_9624,N_9178,N_7602);
or U9625 (N_9625,N_8185,N_6475);
xor U9626 (N_9626,N_6610,N_8911);
and U9627 (N_9627,N_8677,N_7687);
and U9628 (N_9628,N_6701,N_8603);
or U9629 (N_9629,N_6493,N_8862);
and U9630 (N_9630,N_8872,N_9356);
or U9631 (N_9631,N_7715,N_8010);
nor U9632 (N_9632,N_7307,N_7530);
nand U9633 (N_9633,N_6305,N_8839);
or U9634 (N_9634,N_8556,N_7029);
nand U9635 (N_9635,N_7894,N_6661);
xnor U9636 (N_9636,N_8851,N_6996);
and U9637 (N_9637,N_8025,N_7457);
and U9638 (N_9638,N_7378,N_8210);
nand U9639 (N_9639,N_8547,N_6499);
xor U9640 (N_9640,N_8257,N_8986);
nor U9641 (N_9641,N_8485,N_9003);
xor U9642 (N_9642,N_6294,N_7496);
and U9643 (N_9643,N_7238,N_6907);
or U9644 (N_9644,N_9035,N_9054);
and U9645 (N_9645,N_9050,N_8752);
nand U9646 (N_9646,N_6277,N_9044);
xor U9647 (N_9647,N_7467,N_7290);
nand U9648 (N_9648,N_6403,N_6748);
xnor U9649 (N_9649,N_9287,N_8174);
nor U9650 (N_9650,N_6775,N_8125);
nor U9651 (N_9651,N_6730,N_8131);
and U9652 (N_9652,N_7400,N_8975);
nor U9653 (N_9653,N_8147,N_6987);
or U9654 (N_9654,N_8108,N_6879);
and U9655 (N_9655,N_7161,N_8285);
nand U9656 (N_9656,N_9020,N_7817);
or U9657 (N_9657,N_8140,N_8247);
and U9658 (N_9658,N_9143,N_7601);
or U9659 (N_9659,N_6875,N_8572);
nor U9660 (N_9660,N_8880,N_7811);
or U9661 (N_9661,N_7393,N_7187);
nand U9662 (N_9662,N_7728,N_8307);
and U9663 (N_9663,N_6510,N_7329);
nand U9664 (N_9664,N_7404,N_6733);
and U9665 (N_9665,N_9339,N_6953);
or U9666 (N_9666,N_6417,N_6391);
and U9667 (N_9667,N_6572,N_8770);
or U9668 (N_9668,N_7341,N_7331);
or U9669 (N_9669,N_8602,N_9082);
and U9670 (N_9670,N_8683,N_7517);
nand U9671 (N_9671,N_8947,N_7146);
nand U9672 (N_9672,N_7373,N_7725);
nor U9673 (N_9673,N_6469,N_8980);
and U9674 (N_9674,N_6902,N_7885);
and U9675 (N_9675,N_7759,N_7873);
or U9676 (N_9676,N_6456,N_7042);
nor U9677 (N_9677,N_8650,N_7572);
nor U9678 (N_9678,N_9214,N_6641);
nand U9679 (N_9679,N_8397,N_8745);
nand U9680 (N_9680,N_8278,N_8768);
or U9681 (N_9681,N_7409,N_7340);
and U9682 (N_9682,N_8609,N_9079);
nor U9683 (N_9683,N_7569,N_6657);
nand U9684 (N_9684,N_8854,N_7274);
nor U9685 (N_9685,N_7273,N_7176);
or U9686 (N_9686,N_9169,N_7289);
or U9687 (N_9687,N_8175,N_8091);
or U9688 (N_9688,N_7643,N_7233);
nand U9689 (N_9689,N_8651,N_8618);
nand U9690 (N_9690,N_8724,N_8509);
or U9691 (N_9691,N_7311,N_8450);
and U9692 (N_9692,N_6916,N_7688);
nor U9693 (N_9693,N_6455,N_6538);
nor U9694 (N_9694,N_8829,N_7853);
nor U9695 (N_9695,N_8876,N_8286);
nor U9696 (N_9696,N_8985,N_8543);
nor U9697 (N_9697,N_9013,N_9254);
nor U9698 (N_9698,N_6662,N_9279);
and U9699 (N_9699,N_7008,N_7232);
nor U9700 (N_9700,N_8657,N_8405);
nor U9701 (N_9701,N_8166,N_6445);
nand U9702 (N_9702,N_8519,N_8914);
and U9703 (N_9703,N_9249,N_8571);
xor U9704 (N_9704,N_7740,N_6581);
or U9705 (N_9705,N_7652,N_8424);
xor U9706 (N_9706,N_7056,N_7312);
nor U9707 (N_9707,N_8594,N_8406);
nor U9708 (N_9708,N_7919,N_8277);
xor U9709 (N_9709,N_6546,N_7085);
and U9710 (N_9710,N_8977,N_6488);
nor U9711 (N_9711,N_7431,N_8216);
nand U9712 (N_9712,N_6626,N_7175);
or U9713 (N_9713,N_8595,N_8187);
nor U9714 (N_9714,N_8137,N_6665);
nand U9715 (N_9715,N_7698,N_7208);
nor U9716 (N_9716,N_8803,N_6724);
and U9717 (N_9717,N_6498,N_7011);
nor U9718 (N_9718,N_9365,N_7384);
nand U9719 (N_9719,N_8363,N_7564);
nand U9720 (N_9720,N_7699,N_8661);
xor U9721 (N_9721,N_9072,N_7867);
xor U9722 (N_9722,N_8263,N_6374);
nand U9723 (N_9723,N_7892,N_6763);
nand U9724 (N_9724,N_6656,N_8753);
and U9725 (N_9725,N_6378,N_8139);
nand U9726 (N_9726,N_6406,N_8231);
nor U9727 (N_9727,N_7640,N_8830);
or U9728 (N_9728,N_6929,N_8276);
and U9729 (N_9729,N_7320,N_8123);
xor U9730 (N_9730,N_8940,N_9225);
nand U9731 (N_9731,N_6367,N_8520);
or U9732 (N_9732,N_9045,N_8831);
nor U9733 (N_9733,N_6732,N_7689);
nor U9734 (N_9734,N_7482,N_6524);
xnor U9735 (N_9735,N_6516,N_8979);
nand U9736 (N_9736,N_6601,N_7016);
or U9737 (N_9737,N_6749,N_7001);
xor U9738 (N_9738,N_6278,N_6467);
or U9739 (N_9739,N_6901,N_8297);
or U9740 (N_9740,N_8328,N_7140);
nor U9741 (N_9741,N_6663,N_7207);
or U9742 (N_9742,N_7907,N_8965);
and U9743 (N_9743,N_7421,N_8816);
nor U9744 (N_9744,N_7801,N_7814);
nand U9745 (N_9745,N_6465,N_7635);
or U9746 (N_9746,N_7439,N_7600);
and U9747 (N_9747,N_8096,N_6348);
or U9748 (N_9748,N_8935,N_8239);
or U9749 (N_9749,N_8867,N_8102);
nor U9750 (N_9750,N_8492,N_6373);
nand U9751 (N_9751,N_8855,N_8400);
nor U9752 (N_9752,N_6310,N_7755);
nand U9753 (N_9753,N_7310,N_7658);
nand U9754 (N_9754,N_6550,N_7747);
or U9755 (N_9755,N_8499,N_7766);
and U9756 (N_9756,N_7343,N_7092);
nand U9757 (N_9757,N_7354,N_7781);
nand U9758 (N_9758,N_7610,N_8479);
and U9759 (N_9759,N_8063,N_8806);
nor U9760 (N_9760,N_7223,N_6534);
nand U9761 (N_9761,N_8681,N_7488);
or U9762 (N_9762,N_6620,N_7437);
nor U9763 (N_9763,N_6539,N_7788);
nand U9764 (N_9764,N_9293,N_6798);
nor U9765 (N_9765,N_8403,N_7491);
and U9766 (N_9766,N_8845,N_8721);
and U9767 (N_9767,N_7380,N_6934);
or U9768 (N_9768,N_7412,N_9349);
nand U9769 (N_9769,N_6847,N_8497);
or U9770 (N_9770,N_9274,N_6593);
and U9771 (N_9771,N_8478,N_7691);
or U9772 (N_9772,N_7481,N_7213);
and U9773 (N_9773,N_7502,N_6992);
and U9774 (N_9774,N_6269,N_7358);
nand U9775 (N_9775,N_6509,N_8993);
or U9776 (N_9776,N_7401,N_6338);
or U9777 (N_9777,N_8670,N_8438);
nand U9778 (N_9778,N_6567,N_7910);
nand U9779 (N_9779,N_6773,N_9354);
nand U9780 (N_9780,N_7533,N_9047);
nor U9781 (N_9781,N_7840,N_8527);
nor U9782 (N_9782,N_6438,N_6959);
and U9783 (N_9783,N_7228,N_6638);
nor U9784 (N_9784,N_7827,N_9313);
nand U9785 (N_9785,N_8311,N_7684);
and U9786 (N_9786,N_9189,N_8398);
nor U9787 (N_9787,N_8336,N_6579);
nand U9788 (N_9788,N_7178,N_7750);
or U9789 (N_9789,N_6935,N_8849);
nand U9790 (N_9790,N_8275,N_7046);
nand U9791 (N_9791,N_6453,N_8493);
xor U9792 (N_9792,N_8812,N_7735);
nand U9793 (N_9793,N_6972,N_6861);
or U9794 (N_9794,N_8046,N_8338);
or U9795 (N_9795,N_7511,N_7305);
nor U9796 (N_9796,N_8873,N_9039);
or U9797 (N_9797,N_8703,N_8711);
or U9798 (N_9798,N_8962,N_8524);
nor U9799 (N_9799,N_9027,N_6667);
nand U9800 (N_9800,N_6883,N_6721);
and U9801 (N_9801,N_7930,N_8559);
and U9802 (N_9802,N_6472,N_6335);
xnor U9803 (N_9803,N_6530,N_7999);
or U9804 (N_9804,N_6675,N_9157);
or U9805 (N_9805,N_7392,N_8268);
nand U9806 (N_9806,N_7107,N_8838);
or U9807 (N_9807,N_6336,N_7831);
nand U9808 (N_9808,N_7960,N_7774);
or U9809 (N_9809,N_9311,N_8121);
xor U9810 (N_9810,N_8662,N_8453);
and U9811 (N_9811,N_6313,N_7667);
and U9812 (N_9812,N_8169,N_8832);
or U9813 (N_9813,N_6483,N_8018);
xnor U9814 (N_9814,N_6725,N_9066);
nor U9815 (N_9815,N_8009,N_6585);
or U9816 (N_9816,N_6614,N_7144);
or U9817 (N_9817,N_8120,N_9259);
or U9818 (N_9818,N_6922,N_6621);
nor U9819 (N_9819,N_8264,N_6421);
nand U9820 (N_9820,N_9081,N_8075);
xnor U9821 (N_9821,N_6253,N_6770);
nand U9822 (N_9822,N_6894,N_7054);
nand U9823 (N_9823,N_7608,N_7088);
or U9824 (N_9824,N_8542,N_6945);
or U9825 (N_9825,N_7198,N_8928);
and U9826 (N_9826,N_8481,N_8537);
xor U9827 (N_9827,N_6457,N_8908);
nand U9828 (N_9828,N_6905,N_6295);
nand U9829 (N_9829,N_8533,N_6911);
xor U9830 (N_9830,N_7115,N_7131);
and U9831 (N_9831,N_9165,N_7451);
nor U9832 (N_9832,N_8391,N_7897);
or U9833 (N_9833,N_8749,N_7216);
nand U9834 (N_9834,N_8821,N_6944);
and U9835 (N_9835,N_6340,N_9176);
nor U9836 (N_9836,N_6636,N_6320);
or U9837 (N_9837,N_7141,N_7156);
and U9838 (N_9838,N_7368,N_8077);
nand U9839 (N_9839,N_6960,N_6908);
nand U9840 (N_9840,N_8705,N_7136);
nand U9841 (N_9841,N_9133,N_7806);
nor U9842 (N_9842,N_7283,N_8004);
and U9843 (N_9843,N_7916,N_7126);
nand U9844 (N_9844,N_8083,N_7648);
nand U9845 (N_9845,N_7411,N_7032);
or U9846 (N_9846,N_9075,N_9246);
nand U9847 (N_9847,N_7833,N_8932);
nand U9848 (N_9848,N_7444,N_7454);
and U9849 (N_9849,N_7538,N_7057);
or U9850 (N_9850,N_6742,N_6718);
nand U9851 (N_9851,N_7534,N_8296);
nand U9852 (N_9852,N_7366,N_8061);
and U9853 (N_9853,N_6947,N_6737);
nand U9854 (N_9854,N_6413,N_8404);
nand U9855 (N_9855,N_6988,N_8060);
nor U9856 (N_9856,N_6937,N_7676);
or U9857 (N_9857,N_6873,N_7862);
or U9858 (N_9858,N_7636,N_8383);
nor U9859 (N_9859,N_6420,N_9262);
or U9860 (N_9860,N_7347,N_8260);
xor U9861 (N_9861,N_6973,N_6290);
or U9862 (N_9862,N_9115,N_6910);
or U9863 (N_9863,N_6334,N_9321);
nand U9864 (N_9864,N_9312,N_7839);
and U9865 (N_9865,N_7248,N_8190);
nand U9866 (N_9866,N_6542,N_6449);
nor U9867 (N_9867,N_9198,N_8966);
and U9868 (N_9868,N_6781,N_8154);
nand U9869 (N_9869,N_7995,N_8580);
or U9870 (N_9870,N_9106,N_9094);
or U9871 (N_9871,N_7174,N_7630);
nor U9872 (N_9872,N_7943,N_6723);
nor U9873 (N_9873,N_7406,N_6747);
or U9874 (N_9874,N_7686,N_8245);
xor U9875 (N_9875,N_7397,N_7731);
nand U9876 (N_9876,N_6887,N_9305);
or U9877 (N_9877,N_9253,N_6728);
nand U9878 (N_9878,N_7926,N_6447);
or U9879 (N_9879,N_6537,N_9182);
or U9880 (N_9880,N_9346,N_9121);
nor U9881 (N_9881,N_6324,N_7931);
nand U9882 (N_9882,N_7403,N_7588);
or U9883 (N_9883,N_6291,N_8441);
and U9884 (N_9884,N_7155,N_8573);
nand U9885 (N_9885,N_8151,N_8168);
xor U9886 (N_9886,N_9340,N_7863);
or U9887 (N_9887,N_8626,N_7721);
or U9888 (N_9888,N_9272,N_8094);
or U9889 (N_9889,N_6746,N_8486);
xnor U9890 (N_9890,N_7422,N_9360);
and U9891 (N_9891,N_8884,N_7263);
or U9892 (N_9892,N_9278,N_8597);
or U9893 (N_9893,N_7717,N_9186);
and U9894 (N_9894,N_7542,N_9224);
nor U9895 (N_9895,N_6261,N_7937);
xnor U9896 (N_9896,N_9361,N_8198);
nor U9897 (N_9897,N_7402,N_6432);
and U9898 (N_9898,N_7872,N_8765);
xnor U9899 (N_9899,N_7286,N_8696);
and U9900 (N_9900,N_6577,N_8565);
and U9901 (N_9901,N_6766,N_9187);
nand U9902 (N_9902,N_6681,N_6741);
nor U9903 (N_9903,N_9129,N_8462);
nand U9904 (N_9904,N_8648,N_7849);
and U9905 (N_9905,N_7835,N_7417);
and U9906 (N_9906,N_7695,N_8706);
and U9907 (N_9907,N_8211,N_8218);
or U9908 (N_9908,N_7109,N_6711);
xnor U9909 (N_9909,N_6418,N_7951);
and U9910 (N_9910,N_7236,N_7841);
or U9911 (N_9911,N_8490,N_6513);
or U9912 (N_9912,N_6697,N_6881);
nand U9913 (N_9913,N_6655,N_6297);
or U9914 (N_9914,N_7752,N_8685);
and U9915 (N_9915,N_7033,N_8022);
nor U9916 (N_9916,N_9101,N_7642);
and U9917 (N_9917,N_8647,N_8409);
nand U9918 (N_9918,N_6415,N_7754);
and U9919 (N_9919,N_6827,N_6299);
and U9920 (N_9920,N_7436,N_8469);
nand U9921 (N_9921,N_7629,N_7250);
and U9922 (N_9922,N_8632,N_8003);
nor U9923 (N_9923,N_8017,N_6470);
nand U9924 (N_9924,N_9315,N_9018);
nand U9925 (N_9925,N_9011,N_9107);
nor U9926 (N_9926,N_7815,N_7532);
nor U9927 (N_9927,N_6793,N_7888);
or U9928 (N_9928,N_7172,N_7944);
and U9929 (N_9929,N_8922,N_7976);
xor U9930 (N_9930,N_8261,N_9331);
nand U9931 (N_9931,N_6840,N_8316);
nor U9932 (N_9932,N_6339,N_8407);
nor U9933 (N_9933,N_8314,N_8252);
xnor U9934 (N_9934,N_8287,N_6270);
nor U9935 (N_9935,N_7586,N_8348);
or U9936 (N_9936,N_7515,N_8081);
nor U9937 (N_9937,N_6482,N_8785);
and U9938 (N_9938,N_7321,N_8722);
nor U9939 (N_9939,N_6669,N_6501);
and U9940 (N_9940,N_7328,N_6512);
xor U9941 (N_9941,N_8638,N_7039);
nor U9942 (N_9942,N_7965,N_7345);
xor U9943 (N_9943,N_7616,N_7268);
xnor U9944 (N_9944,N_6932,N_9286);
nor U9945 (N_9945,N_8688,N_6658);
nand U9946 (N_9946,N_7129,N_6948);
nor U9947 (N_9947,N_9128,N_9049);
nor U9948 (N_9948,N_6589,N_8636);
nand U9949 (N_9949,N_6634,N_8513);
and U9950 (N_9950,N_6821,N_9117);
nand U9951 (N_9951,N_6586,N_8393);
nand U9952 (N_9952,N_8095,N_6536);
nand U9953 (N_9953,N_8819,N_7296);
xor U9954 (N_9954,N_8548,N_6952);
or U9955 (N_9955,N_6845,N_7991);
and U9956 (N_9956,N_9238,N_7388);
or U9957 (N_9957,N_8114,N_9034);
nor U9958 (N_9958,N_8097,N_7220);
nand U9959 (N_9959,N_9195,N_8418);
and U9960 (N_9960,N_8918,N_9092);
nor U9961 (N_9961,N_8523,N_7718);
or U9962 (N_9962,N_6494,N_8196);
nor U9963 (N_9963,N_6815,N_8477);
xnor U9964 (N_9964,N_7645,N_8633);
and U9965 (N_9965,N_9297,N_7712);
nor U9966 (N_9966,N_8319,N_7045);
nor U9967 (N_9967,N_9098,N_9086);
nand U9968 (N_9968,N_7810,N_8044);
and U9969 (N_9969,N_6250,N_8413);
and U9970 (N_9970,N_6298,N_7751);
nand U9971 (N_9971,N_7185,N_8983);
nor U9972 (N_9972,N_6690,N_8281);
nor U9973 (N_9973,N_8669,N_8531);
nand U9974 (N_9974,N_6264,N_7487);
xor U9975 (N_9975,N_7964,N_7449);
or U9976 (N_9976,N_6956,N_6943);
nand U9977 (N_9977,N_7789,N_9030);
and U9978 (N_9978,N_7968,N_7554);
nand U9979 (N_9979,N_6410,N_6906);
and U9980 (N_9980,N_9374,N_8272);
nor U9981 (N_9981,N_7240,N_8973);
nor U9982 (N_9982,N_6556,N_7527);
xnor U9983 (N_9983,N_6471,N_8600);
or U9984 (N_9984,N_6426,N_8813);
xor U9985 (N_9985,N_7992,N_6603);
and U9986 (N_9986,N_9210,N_9149);
xnor U9987 (N_9987,N_6548,N_9316);
and U9988 (N_9988,N_8041,N_7927);
xnor U9989 (N_9989,N_7342,N_7898);
nand U9990 (N_9990,N_7153,N_7972);
and U9991 (N_9991,N_8345,N_6317);
or U9992 (N_9992,N_8001,N_6321);
and U9993 (N_9993,N_8142,N_8191);
nor U9994 (N_9994,N_6696,N_8708);
or U9995 (N_9995,N_7575,N_8401);
and U9996 (N_9996,N_8228,N_8560);
nor U9997 (N_9997,N_6703,N_6540);
nor U9998 (N_9998,N_6869,N_6400);
or U9999 (N_9999,N_7120,N_8978);
xor U10000 (N_10000,N_9123,N_7679);
xor U10001 (N_10001,N_6760,N_8117);
nand U10002 (N_10002,N_8329,N_8402);
and U10003 (N_10003,N_8273,N_7077);
nor U10004 (N_10004,N_7670,N_6838);
and U10005 (N_10005,N_8920,N_7091);
xnor U10006 (N_10006,N_7860,N_6968);
or U10007 (N_10007,N_9048,N_7845);
and U10008 (N_10008,N_6698,N_9351);
or U10009 (N_10009,N_6693,N_8099);
nand U10010 (N_10010,N_6964,N_8437);
nand U10011 (N_10011,N_7078,N_7272);
and U10012 (N_10012,N_8037,N_7456);
or U10013 (N_10013,N_6437,N_8575);
nand U10014 (N_10014,N_8074,N_8449);
nor U10015 (N_10015,N_9350,N_8972);
nand U10016 (N_10016,N_7631,N_9322);
and U10017 (N_10017,N_7438,N_6315);
xnor U10018 (N_10018,N_8354,N_8795);
xnor U10019 (N_10019,N_7701,N_8235);
and U10020 (N_10020,N_8206,N_8777);
nor U10021 (N_10021,N_7646,N_6527);
or U10022 (N_10022,N_8625,N_6345);
nand U10023 (N_10023,N_8503,N_8408);
and U10024 (N_10024,N_9359,N_6926);
or U10025 (N_10025,N_6326,N_7117);
or U10026 (N_10026,N_7591,N_7479);
or U10027 (N_10027,N_7547,N_6720);
and U10028 (N_10028,N_7428,N_9260);
xnor U10029 (N_10029,N_8416,N_6750);
and U10030 (N_10030,N_8331,N_6596);
nand U10031 (N_10031,N_6583,N_6491);
or U10032 (N_10032,N_6870,N_8963);
or U10033 (N_10033,N_8860,N_6284);
and U10034 (N_10034,N_7986,N_9306);
or U10035 (N_10035,N_7152,N_8325);
xor U10036 (N_10036,N_8698,N_8664);
or U10037 (N_10037,N_8974,N_7151);
nand U10038 (N_10038,N_7627,N_7832);
nor U10039 (N_10039,N_7364,N_7906);
or U10040 (N_10040,N_6754,N_8370);
nor U10041 (N_10041,N_6592,N_7823);
nand U10042 (N_10042,N_8801,N_7300);
or U10043 (N_10043,N_8760,N_6370);
xor U10044 (N_10044,N_7125,N_8554);
nand U10045 (N_10045,N_6381,N_7878);
and U10046 (N_10046,N_8484,N_8208);
and U10047 (N_10047,N_8525,N_7234);
nor U10048 (N_10048,N_9244,N_7621);
and U10049 (N_10049,N_9277,N_6963);
and U10050 (N_10050,N_8414,N_8082);
nand U10051 (N_10051,N_8521,N_8794);
nor U10052 (N_10052,N_6734,N_6859);
or U10053 (N_10053,N_7206,N_9325);
nand U10054 (N_10054,N_6648,N_7908);
nand U10055 (N_10055,N_7800,N_8432);
and U10056 (N_10056,N_7877,N_8797);
nand U10057 (N_10057,N_6890,N_9268);
nand U10058 (N_10058,N_7585,N_8758);
nor U10059 (N_10059,N_6777,N_6476);
or U10060 (N_10060,N_7447,N_7966);
nand U10061 (N_10061,N_8624,N_7540);
nand U10062 (N_10062,N_8322,N_6505);
nor U10063 (N_10063,N_7605,N_9328);
or U10064 (N_10064,N_6575,N_7038);
xnor U10065 (N_10065,N_9310,N_9113);
nand U10066 (N_10066,N_7875,N_8475);
or U10067 (N_10067,N_6281,N_7710);
nor U10068 (N_10068,N_8014,N_6630);
xnor U10069 (N_10069,N_8289,N_6458);
xnor U10070 (N_10070,N_6303,N_7730);
nor U10071 (N_10071,N_6544,N_9183);
or U10072 (N_10072,N_8895,N_7281);
nand U10073 (N_10073,N_7659,N_6918);
or U10074 (N_10074,N_9010,N_9196);
nor U10075 (N_10075,N_7067,N_7881);
nor U10076 (N_10076,N_9167,N_7531);
or U10077 (N_10077,N_6714,N_6958);
and U10078 (N_10078,N_8923,N_6569);
and U10079 (N_10079,N_8253,N_9302);
xnor U10080 (N_10080,N_7537,N_8642);
or U10081 (N_10081,N_7420,N_6598);
and U10082 (N_10082,N_7837,N_9265);
and U10083 (N_10083,N_9006,N_7551);
nand U10084 (N_10084,N_7302,N_7169);
nand U10085 (N_10085,N_9343,N_9367);
and U10086 (N_10086,N_6708,N_6330);
nor U10087 (N_10087,N_7724,N_7799);
or U10088 (N_10088,N_9077,N_7003);
nor U10089 (N_10089,N_6565,N_7168);
nor U10090 (N_10090,N_7106,N_6495);
and U10091 (N_10091,N_7010,N_7112);
nand U10092 (N_10092,N_6580,N_8541);
or U10093 (N_10093,N_9132,N_6917);
xor U10094 (N_10094,N_8606,N_6428);
and U10095 (N_10095,N_9088,N_8858);
nor U10096 (N_10096,N_7734,N_7775);
nand U10097 (N_10097,N_9042,N_9067);
or U10098 (N_10098,N_9292,N_8942);
nor U10099 (N_10099,N_6679,N_8805);
nand U10100 (N_10100,N_8968,N_8494);
or U10101 (N_10101,N_7606,N_9269);
nor U10102 (N_10102,N_8598,N_7859);
nand U10103 (N_10103,N_9209,N_6686);
and U10104 (N_10104,N_6668,N_7119);
nor U10105 (N_10105,N_8070,N_8898);
nor U10106 (N_10106,N_8103,N_8817);
or U10107 (N_10107,N_9041,N_7355);
nand U10108 (N_10108,N_7440,N_7886);
nor U10109 (N_10109,N_7317,N_8578);
and U10110 (N_10110,N_9093,N_6354);
and U10111 (N_10111,N_6398,N_6986);
xor U10112 (N_10112,N_6412,N_7522);
or U10113 (N_10113,N_9255,N_8483);
and U10114 (N_10114,N_8784,N_9208);
nand U10115 (N_10115,N_7702,N_8086);
nor U10116 (N_10116,N_7558,N_7013);
or U10117 (N_10117,N_6507,N_6805);
nor U10118 (N_10118,N_7887,N_6995);
nor U10119 (N_10119,N_8915,N_7314);
and U10120 (N_10120,N_8737,N_7803);
xor U10121 (N_10121,N_6806,N_7609);
and U10122 (N_10122,N_8874,N_7252);
or U10123 (N_10123,N_6764,N_8237);
xor U10124 (N_10124,N_8823,N_6312);
or U10125 (N_10125,N_8035,N_7594);
and U10126 (N_10126,N_7675,N_7469);
nand U10127 (N_10127,N_8847,N_7545);
nand U10128 (N_10128,N_8042,N_6954);
and U10129 (N_10129,N_6622,N_7101);
or U10130 (N_10130,N_7506,N_8087);
and U10131 (N_10131,N_7812,N_7500);
and U10132 (N_10132,N_9124,N_6888);
nor U10133 (N_10133,N_7828,N_7959);
or U10134 (N_10134,N_7864,N_8646);
or U10135 (N_10135,N_6702,N_7834);
nand U10136 (N_10136,N_8280,N_8241);
or U10137 (N_10137,N_6974,N_6419);
or U10138 (N_10138,N_8644,N_8719);
nor U10139 (N_10139,N_8092,N_9308);
or U10140 (N_10140,N_6717,N_9033);
nand U10141 (N_10141,N_6823,N_8269);
nor U10142 (N_10142,N_6707,N_7733);
nand U10143 (N_10143,N_7332,N_8221);
and U10144 (N_10144,N_6343,N_8964);
nand U10145 (N_10145,N_7434,N_6625);
nand U10146 (N_10146,N_8807,N_7749);
xor U10147 (N_10147,N_8065,N_7776);
nor U10148 (N_10148,N_7195,N_6531);
xnor U10149 (N_10149,N_7157,N_9089);
or U10150 (N_10150,N_7478,N_9166);
nor U10151 (N_10151,N_7330,N_8987);
and U10152 (N_10152,N_6440,N_8146);
nor U10153 (N_10153,N_6914,N_7241);
nand U10154 (N_10154,N_8555,N_8748);
nor U10155 (N_10155,N_7295,N_8716);
or U10156 (N_10156,N_9220,N_9215);
nor U10157 (N_10157,N_9233,N_6808);
nand U10158 (N_10158,N_8659,N_7493);
and U10159 (N_10159,N_6399,N_7825);
or U10160 (N_10160,N_8679,N_8534);
and U10161 (N_10161,N_8133,N_8843);
xnor U10162 (N_10162,N_6965,N_8943);
nand U10163 (N_10163,N_6765,N_8323);
and U10164 (N_10164,N_9201,N_6563);
nand U10165 (N_10165,N_7655,N_7935);
nor U10166 (N_10166,N_8995,N_6877);
nor U10167 (N_10167,N_8804,N_7095);
nand U10168 (N_10168,N_7254,N_8176);
or U10169 (N_10169,N_6772,N_6761);
and U10170 (N_10170,N_8240,N_6328);
or U10171 (N_10171,N_7820,N_7546);
and U10172 (N_10172,N_8549,N_7308);
or U10173 (N_10173,N_8574,N_8049);
nor U10174 (N_10174,N_7304,N_7190);
nor U10175 (N_10175,N_9145,N_7556);
nand U10176 (N_10176,N_8967,N_9055);
or U10177 (N_10177,N_7405,N_7626);
nand U10178 (N_10178,N_8991,N_7882);
and U10179 (N_10179,N_8526,N_6784);
nor U10180 (N_10180,N_6751,N_8996);
or U10181 (N_10181,N_8924,N_7979);
or U10182 (N_10182,N_6319,N_7971);
nor U10183 (N_10183,N_7519,N_7706);
nand U10184 (N_10184,N_7736,N_8270);
xor U10185 (N_10185,N_6673,N_9162);
or U10186 (N_10186,N_7159,N_7270);
and U10187 (N_10187,N_7138,N_6497);
and U10188 (N_10188,N_6523,N_7813);
xor U10189 (N_10189,N_6844,N_7259);
nor U10190 (N_10190,N_9326,N_7905);
or U10191 (N_10191,N_6695,N_7231);
and U10192 (N_10192,N_6506,N_8234);
nand U10193 (N_10193,N_6411,N_9303);
and U10194 (N_10194,N_6503,N_9102);
nor U10195 (N_10195,N_9168,N_8776);
nor U10196 (N_10196,N_7235,N_8678);
nor U10197 (N_10197,N_8982,N_7266);
and U10198 (N_10198,N_6651,N_8173);
and U10199 (N_10199,N_8799,N_7453);
nor U10200 (N_10200,N_7495,N_6993);
nand U10201 (N_10201,N_6504,N_6649);
xor U10202 (N_10202,N_7100,N_7921);
nand U10203 (N_10203,N_7946,N_9223);
nor U10204 (N_10204,N_8188,N_8019);
or U10205 (N_10205,N_7891,N_9283);
nor U10206 (N_10206,N_9099,N_7450);
nand U10207 (N_10207,N_7516,N_9216);
nor U10208 (N_10208,N_7990,N_7483);
nor U10209 (N_10209,N_8283,N_6780);
xor U10210 (N_10210,N_8181,N_7672);
nor U10211 (N_10211,N_7720,N_7425);
and U10212 (N_10212,N_8024,N_6570);
and U10213 (N_10213,N_8080,N_7191);
or U10214 (N_10214,N_6547,N_7086);
or U10215 (N_10215,N_7215,N_8692);
or U10216 (N_10216,N_6629,N_6644);
and U10217 (N_10217,N_6275,N_6562);
nor U10218 (N_10218,N_6408,N_6836);
nor U10219 (N_10219,N_8930,N_8473);
or U10220 (N_10220,N_8802,N_7166);
nand U10221 (N_10221,N_7247,N_9078);
and U10222 (N_10222,N_6385,N_8369);
nand U10223 (N_10223,N_7879,N_9295);
xor U10224 (N_10224,N_7084,N_9100);
or U10225 (N_10225,N_6654,N_7783);
nor U10226 (N_10226,N_8300,N_8412);
and U10227 (N_10227,N_8290,N_7346);
nor U10228 (N_10228,N_7568,N_9142);
and U10229 (N_10229,N_7280,N_8223);
or U10230 (N_10230,N_8332,N_7518);
nor U10231 (N_10231,N_8350,N_7486);
nor U10232 (N_10232,N_6756,N_7977);
nor U10233 (N_10233,N_6487,N_8066);
and U10234 (N_10234,N_8372,N_7276);
nand U10235 (N_10235,N_8887,N_8284);
nand U10236 (N_10236,N_6919,N_8279);
or U10237 (N_10237,N_8587,N_7344);
or U10238 (N_10238,N_7954,N_8232);
and U10239 (N_10239,N_7473,N_8431);
nor U10240 (N_10240,N_8810,N_9063);
nor U10241 (N_10241,N_6351,N_6970);
nand U10242 (N_10242,N_7287,N_6981);
nor U10243 (N_10243,N_6831,N_7352);
xor U10244 (N_10244,N_6689,N_7379);
nor U10245 (N_10245,N_6866,N_6617);
nand U10246 (N_10246,N_6574,N_8333);
xnor U10247 (N_10247,N_8330,N_8145);
and U10248 (N_10248,N_6511,N_9076);
nand U10249 (N_10249,N_7205,N_8182);
and U10250 (N_10250,N_7291,N_9357);
and U10251 (N_10251,N_8134,N_8026);
or U10252 (N_10252,N_8733,N_8036);
nand U10253 (N_10253,N_9329,N_7293);
and U10254 (N_10254,N_6473,N_9147);
xor U10255 (N_10255,N_7181,N_7452);
xnor U10256 (N_10256,N_7377,N_8315);
or U10257 (N_10257,N_7360,N_6966);
and U10258 (N_10258,N_9091,N_6464);
nand U10259 (N_10259,N_8034,N_9235);
and U10260 (N_10260,N_7049,N_6913);
and U10261 (N_10261,N_7323,N_8535);
and U10262 (N_10262,N_8925,N_7073);
nor U10263 (N_10263,N_7104,N_7282);
xor U10264 (N_10264,N_6841,N_7162);
nand U10265 (N_10265,N_9304,N_6797);
or U10266 (N_10266,N_8098,N_7855);
nand U10267 (N_10267,N_7997,N_8516);
and U10268 (N_10268,N_8764,N_9112);
and U10269 (N_10269,N_9118,N_7939);
nor U10270 (N_10270,N_7662,N_8889);
or U10271 (N_10271,N_6645,N_7501);
nor U10272 (N_10272,N_6545,N_6903);
and U10273 (N_10273,N_6842,N_7285);
and U10274 (N_10274,N_7726,N_8184);
or U10275 (N_10275,N_9060,N_8905);
or U10276 (N_10276,N_8507,N_7395);
nand U10277 (N_10277,N_6710,N_8150);
nor U10278 (N_10278,N_6683,N_9002);
nor U10279 (N_10279,N_6301,N_7367);
or U10280 (N_10280,N_7957,N_6599);
nor U10281 (N_10281,N_8032,N_7398);
nor U10282 (N_10282,N_6687,N_6369);
nand U10283 (N_10283,N_9261,N_8689);
nand U10284 (N_10284,N_7746,N_7786);
xnor U10285 (N_10285,N_7407,N_8868);
nor U10286 (N_10286,N_7309,N_6950);
nand U10287 (N_10287,N_8504,N_8426);
xor U10288 (N_10288,N_8852,N_7102);
and U10289 (N_10289,N_7226,N_9299);
nor U10290 (N_10290,N_6985,N_8903);
nor U10291 (N_10291,N_7026,N_8382);
nor U10292 (N_10292,N_8192,N_8148);
nor U10293 (N_10293,N_8468,N_9138);
nand U10294 (N_10294,N_8459,N_8073);
nand U10295 (N_10295,N_6300,N_7993);
nand U10296 (N_10296,N_7149,N_6704);
or U10297 (N_10297,N_7987,N_9177);
or U10298 (N_10298,N_9131,N_9040);
nor U10299 (N_10299,N_7306,N_6889);
nand U10300 (N_10300,N_7284,N_9023);
nand U10301 (N_10301,N_6646,N_8428);
and U10302 (N_10302,N_6390,N_8881);
nor U10303 (N_10303,N_8564,N_6397);
nand U10304 (N_10304,N_9337,N_6853);
and U10305 (N_10305,N_8791,N_9144);
or U10306 (N_10306,N_7634,N_7415);
and U10307 (N_10307,N_9229,N_6923);
and U10308 (N_10308,N_8747,N_8447);
nand U10309 (N_10309,N_8444,N_9012);
nand U10310 (N_10310,N_6691,N_8199);
and U10311 (N_10311,N_7043,N_6782);
xor U10312 (N_10312,N_9090,N_7051);
xnor U10313 (N_10313,N_9347,N_7549);
nand U10314 (N_10314,N_6480,N_6810);
nor U10315 (N_10315,N_6938,N_9205);
or U10316 (N_10316,N_7649,N_6535);
and U10317 (N_10317,N_8842,N_6404);
or U10318 (N_10318,N_7064,N_7249);
nand U10319 (N_10319,N_8751,N_9275);
or U10320 (N_10320,N_7574,N_7031);
or U10321 (N_10321,N_6396,N_6789);
xnor U10322 (N_10322,N_8233,N_6549);
or U10323 (N_10323,N_8798,N_7315);
or U10324 (N_10324,N_8956,N_6508);
xor U10325 (N_10325,N_6915,N_6774);
or U10326 (N_10326,N_9104,N_7459);
nand U10327 (N_10327,N_7376,N_6520);
nand U10328 (N_10328,N_6896,N_7861);
or U10329 (N_10329,N_6867,N_7809);
or U10330 (N_10330,N_8529,N_7762);
nand U10331 (N_10331,N_6811,N_9344);
or U10332 (N_10332,N_8254,N_8209);
and U10333 (N_10333,N_8078,N_7299);
nand U10334 (N_10334,N_7303,N_7313);
or U10335 (N_10335,N_6616,N_8439);
nand U10336 (N_10336,N_7476,N_7022);
nand U10337 (N_10337,N_8641,N_9193);
or U10338 (N_10338,N_7895,N_8695);
and U10339 (N_10339,N_7145,N_8360);
and U10340 (N_10340,N_6355,N_6606);
and U10341 (N_10341,N_6671,N_7150);
xor U10342 (N_10342,N_6442,N_8656);
nand U10343 (N_10343,N_8452,N_7113);
and U10344 (N_10344,N_8265,N_7142);
nand U10345 (N_10345,N_7470,N_7685);
and U10346 (N_10346,N_6957,N_8373);
xor U10347 (N_10347,N_7566,N_6409);
nand U10348 (N_10348,N_6898,N_8476);
nand U10349 (N_10349,N_7466,N_7948);
or U10350 (N_10350,N_7122,N_9373);
or U10351 (N_10351,N_7327,N_7829);
nand U10352 (N_10352,N_9016,N_7147);
nand U10353 (N_10353,N_7846,N_7578);
xnor U10354 (N_10354,N_8255,N_8466);
nor U10355 (N_10355,N_7912,N_6401);
nor U10356 (N_10356,N_7114,N_8939);
or U10357 (N_10357,N_6386,N_8551);
nand U10358 (N_10358,N_7525,N_7070);
nor U10359 (N_10359,N_8189,N_8544);
nand U10360 (N_10360,N_9298,N_6514);
or U10361 (N_10361,N_6479,N_6788);
or U10362 (N_10362,N_6578,N_8396);
nor U10363 (N_10363,N_8225,N_8610);
nor U10364 (N_10364,N_6899,N_8865);
or U10365 (N_10365,N_7535,N_9160);
or U10366 (N_10366,N_8366,N_6940);
or U10367 (N_10367,N_7694,N_8027);
or U10368 (N_10368,N_8433,N_6352);
and U10369 (N_10369,N_7075,N_9074);
nor U10370 (N_10370,N_7911,N_7461);
nor U10371 (N_10371,N_7581,N_8818);
and U10372 (N_10372,N_7218,N_7105);
or U10373 (N_10373,N_6450,N_8377);
nor U10374 (N_10374,N_8637,N_8031);
and U10375 (N_10375,N_7893,N_8180);
nor U10376 (N_10376,N_7164,N_6739);
nor U10377 (N_10377,N_8514,N_8623);
and U10378 (N_10378,N_7844,N_7563);
nand U10379 (N_10379,N_6262,N_8100);
or U10380 (N_10380,N_8635,N_7203);
and U10381 (N_10381,N_9330,N_8327);
nor U10382 (N_10382,N_7427,N_8808);
nor U10383 (N_10383,N_6416,N_8357);
nand U10384 (N_10384,N_8299,N_8033);
nand U10385 (N_10385,N_8620,N_8105);
and U10386 (N_10386,N_8732,N_8739);
or U10387 (N_10387,N_8460,N_8888);
nand U10388 (N_10388,N_8435,N_7866);
nor U10389 (N_10389,N_7116,N_6568);
nor U10390 (N_10390,N_7816,N_7692);
and U10391 (N_10391,N_8388,N_8825);
and U10392 (N_10392,N_9263,N_7924);
and U10393 (N_10393,N_7719,N_7765);
and U10394 (N_10394,N_6309,N_8230);
nand U10395 (N_10395,N_8246,N_6273);
or U10396 (N_10396,N_8337,N_7027);
nor U10397 (N_10397,N_6560,N_7183);
and U10398 (N_10398,N_8489,N_8313);
nand U10399 (N_10399,N_8540,N_8960);
xnor U10400 (N_10400,N_8714,N_7656);
or U10401 (N_10401,N_7350,N_6712);
nand U10402 (N_10402,N_6283,N_8365);
or U10403 (N_10403,N_8877,N_8957);
or U10404 (N_10404,N_8970,N_8193);
nor U10405 (N_10405,N_8883,N_7258);
nand U10406 (N_10406,N_9234,N_8931);
or U10407 (N_10407,N_8861,N_6525);
and U10408 (N_10408,N_7653,N_7429);
nor U10409 (N_10409,N_8293,N_6678);
and U10410 (N_10410,N_9175,N_8729);
nand U10411 (N_10411,N_9197,N_8530);
nand U10412 (N_10412,N_8202,N_7154);
nand U10413 (N_10413,N_7696,N_7767);
nand U10414 (N_10414,N_6368,N_6882);
nand U10415 (N_10415,N_9173,N_8059);
and U10416 (N_10416,N_7096,N_6517);
and U10417 (N_10417,N_6795,N_9159);
nand U10418 (N_10418,N_6825,N_6713);
or U10419 (N_10419,N_8790,N_7509);
nand U10420 (N_10420,N_7700,N_7507);
or U10421 (N_10421,N_9068,N_7857);
nand U10422 (N_10422,N_7633,N_6685);
nor U10423 (N_10423,N_7416,N_8501);
nand U10424 (N_10424,N_8558,N_6800);
or U10425 (N_10425,N_7681,N_8443);
xor U10426 (N_10426,N_8906,N_8495);
nor U10427 (N_10427,N_7739,N_6994);
nor U10428 (N_10428,N_7615,N_8699);
and U10429 (N_10429,N_6880,N_8612);
nand U10430 (N_10430,N_8505,N_6628);
nor U10431 (N_10431,N_8591,N_7369);
nor U10432 (N_10432,N_7171,N_9109);
and U10433 (N_10433,N_6826,N_6951);
nand U10434 (N_10434,N_8339,N_9046);
nand U10435 (N_10435,N_7201,N_8900);
and U10436 (N_10436,N_6643,N_8318);
nand U10437 (N_10437,N_8054,N_9080);
nor U10438 (N_10438,N_8353,N_8440);
nand U10439 (N_10439,N_9290,N_7214);
xor U10440 (N_10440,N_7325,N_6347);
or U10441 (N_10441,N_6430,N_9032);
nand U10442 (N_10442,N_7560,N_7256);
nand U10443 (N_10443,N_8076,N_8702);
and U10444 (N_10444,N_7000,N_9317);
nor U10445 (N_10445,N_6292,N_8621);
or U10446 (N_10446,N_7071,N_7876);
nor U10447 (N_10447,N_7550,N_7035);
nand U10448 (N_10448,N_6571,N_8422);
or U10449 (N_10449,N_7014,N_8186);
and U10450 (N_10450,N_8859,N_6892);
nor U10451 (N_10451,N_7851,N_6363);
and U10452 (N_10452,N_7784,N_7669);
or U10453 (N_10453,N_6486,N_7446);
or U10454 (N_10454,N_7852,N_6371);
and U10455 (N_10455,N_7764,N_6967);
and U10456 (N_10456,N_9103,N_8068);
or U10457 (N_10457,N_8038,N_7955);
or U10458 (N_10458,N_7387,N_7592);
nand U10459 (N_10459,N_8423,N_8822);
nand U10460 (N_10460,N_7167,N_6874);
nand U10461 (N_10461,N_8172,N_7607);
and U10462 (N_10462,N_7970,N_7089);
xnor U10463 (N_10463,N_9226,N_8792);
nand U10464 (N_10464,N_7773,N_6618);
and U10465 (N_10465,N_8085,N_6659);
and U10466 (N_10466,N_8179,N_9122);
nor U10467 (N_10467,N_7245,N_7889);
or U10468 (N_10468,N_6843,N_8171);
and U10469 (N_10469,N_6318,N_6304);
nor U10470 (N_10470,N_7796,N_9065);
and U10471 (N_10471,N_6627,N_6828);
or U10472 (N_10472,N_8757,N_8341);
or U10473 (N_10473,N_7871,N_8955);
nand U10474 (N_10474,N_6715,N_8057);
or U10475 (N_10475,N_6676,N_7024);
or U10476 (N_10476,N_6346,N_6921);
or U10477 (N_10477,N_8104,N_7336);
nand U10478 (N_10478,N_8250,N_9345);
nor U10479 (N_10479,N_8244,N_7121);
and U10480 (N_10480,N_7744,N_8016);
xor U10481 (N_10481,N_8809,N_8836);
and U10482 (N_10482,N_7363,N_7798);
or U10483 (N_10483,N_9192,N_7772);
or U10484 (N_10484,N_9000,N_7880);
nor U10485 (N_10485,N_8539,N_9362);
or U10486 (N_10486,N_7941,N_9222);
or U10487 (N_10487,N_8392,N_9288);
and U10488 (N_10488,N_9057,N_7925);
nand U10489 (N_10489,N_7528,N_6819);
and U10490 (N_10490,N_9324,N_7514);
xor U10491 (N_10491,N_8740,N_8448);
or U10492 (N_10492,N_6424,N_9108);
nor U10493 (N_10493,N_8773,N_8109);
xor U10494 (N_10494,N_7199,N_6316);
xor U10495 (N_10495,N_7998,N_9369);
or U10496 (N_10496,N_7787,N_8741);
and U10497 (N_10497,N_9087,N_8566);
nand U10498 (N_10498,N_6260,N_8643);
xnor U10499 (N_10499,N_8417,N_8395);
and U10500 (N_10500,N_8837,N_7850);
or U10501 (N_10501,N_6904,N_8342);
nand U10502 (N_10502,N_8762,N_6590);
nand U10503 (N_10503,N_7618,N_7370);
nor U10504 (N_10504,N_7711,N_6864);
xnor U10505 (N_10505,N_7163,N_8291);
nand U10506 (N_10506,N_6716,N_9085);
and U10507 (N_10507,N_8835,N_7802);
or U10508 (N_10508,N_8006,N_6846);
and U10509 (N_10509,N_8676,N_6553);
nand U10510 (N_10510,N_7484,N_6474);
or U10511 (N_10511,N_8508,N_7704);
nand U10512 (N_10512,N_8420,N_6769);
and U10513 (N_10513,N_6848,N_7874);
or U10514 (N_10514,N_8119,N_6623);
nor U10515 (N_10515,N_6329,N_6762);
or U10516 (N_10516,N_6353,N_8562);
or U10517 (N_10517,N_7455,N_7654);
nor U10518 (N_10518,N_8053,N_7595);
or U10519 (N_10519,N_9095,N_8122);
or U10520 (N_10520,N_8820,N_9291);
nor U10521 (N_10521,N_8352,N_8205);
nand U10522 (N_10522,N_8844,N_8712);
or U10523 (N_10523,N_6441,N_6443);
nand U10524 (N_10524,N_8954,N_7625);
nor U10525 (N_10525,N_7468,N_8214);
and U10526 (N_10526,N_7028,N_6532);
nor U10527 (N_10527,N_9029,N_8652);
nand U10528 (N_10528,N_8324,N_6576);
nor U10529 (N_10529,N_9125,N_9120);
nor U10530 (N_10530,N_7275,N_7124);
and U10531 (N_10531,N_7622,N_8613);
nor U10532 (N_10532,N_6461,N_8912);
or U10533 (N_10533,N_7757,N_7414);
or U10534 (N_10534,N_6863,N_7543);
and U10535 (N_10535,N_7442,N_8948);
xnor U10536 (N_10536,N_8238,N_8707);
nand U10537 (N_10537,N_7189,N_8039);
nand U10538 (N_10538,N_8953,N_9323);
or U10539 (N_10539,N_6266,N_7316);
nand U10540 (N_10540,N_8673,N_9250);
nor U10541 (N_10541,N_7561,N_6365);
or U10542 (N_10542,N_8671,N_6314);
and U10543 (N_10543,N_7472,N_7842);
xnor U10544 (N_10544,N_9245,N_6738);
nor U10545 (N_10545,N_9372,N_7678);
or U10546 (N_10546,N_9370,N_7419);
nand U10547 (N_10547,N_6822,N_8159);
nor U10548 (N_10548,N_6925,N_8653);
nor U10549 (N_10549,N_8891,N_8436);
or U10550 (N_10550,N_8717,N_7620);
or U10551 (N_10551,N_6423,N_9204);
nor U10552 (N_10552,N_7660,N_8136);
and U10553 (N_10553,N_8111,N_8249);
and U10554 (N_10554,N_6794,N_8248);
nand U10555 (N_10555,N_7824,N_6376);
nand U10556 (N_10556,N_6814,N_6855);
or U10557 (N_10557,N_7901,N_7590);
nor U10558 (N_10558,N_9200,N_6824);
or U10559 (N_10559,N_7758,N_7267);
or U10560 (N_10560,N_7552,N_8389);
nor U10561 (N_10561,N_7582,N_7385);
nor U10562 (N_10562,N_8158,N_7204);
and U10563 (N_10563,N_7596,N_9150);
or U10564 (N_10564,N_6975,N_8615);
or U10565 (N_10565,N_8227,N_6529);
and U10566 (N_10566,N_8052,N_7212);
nor U10567 (N_10567,N_6635,N_8500);
nand U10568 (N_10568,N_9019,N_7137);
nand U10569 (N_10569,N_7729,N_8294);
or U10570 (N_10570,N_8951,N_8002);
or U10571 (N_10571,N_7539,N_6856);
and U10572 (N_10572,N_6350,N_6971);
nand U10573 (N_10573,N_7587,N_9267);
nand U10574 (N_10574,N_7903,N_7326);
nand U10575 (N_10575,N_6468,N_7529);
nand U10576 (N_10576,N_8072,N_8628);
and U10577 (N_10577,N_9135,N_8601);
and U10578 (N_10578,N_7929,N_7673);
xnor U10579 (N_10579,N_6323,N_7989);
nor U10580 (N_10580,N_7805,N_7918);
or U10581 (N_10581,N_7576,N_8713);
xor U10582 (N_10582,N_8515,N_6405);
or U10583 (N_10583,N_7769,N_8011);
nor U10584 (N_10584,N_6496,N_7513);
nand U10585 (N_10585,N_8934,N_8857);
nor U10586 (N_10586,N_7936,N_7822);
nor U10587 (N_10587,N_7499,N_7920);
nor U10588 (N_10588,N_6341,N_9181);
nor U10589 (N_10589,N_8043,N_7418);
and U10590 (N_10590,N_9134,N_6380);
nand U10591 (N_10591,N_6886,N_7794);
or U10592 (N_10592,N_7647,N_7577);
or U10593 (N_10593,N_7182,N_7756);
nand U10594 (N_10594,N_7557,N_8200);
or U10595 (N_10595,N_7847,N_6802);
or U10596 (N_10596,N_8047,N_7200);
and U10597 (N_10597,N_8243,N_8567);
nor U10598 (N_10598,N_9320,N_8561);
nor U10599 (N_10599,N_7123,N_7707);
nand U10600 (N_10600,N_7261,N_6978);
or U10601 (N_10601,N_8430,N_9171);
nor U10602 (N_10602,N_7058,N_6991);
nor U10603 (N_10603,N_6604,N_8197);
nor U10604 (N_10604,N_8461,N_8605);
nor U10605 (N_10605,N_7870,N_7804);
and U10606 (N_10606,N_6876,N_9266);
and U10607 (N_10607,N_8622,N_8897);
nand U10608 (N_10608,N_8112,N_7227);
xor U10609 (N_10609,N_6276,N_8177);
xor U10610 (N_10610,N_9119,N_8660);
or U10611 (N_10611,N_7464,N_7544);
and U10612 (N_10612,N_6989,N_9270);
nor U10613 (N_10613,N_7371,N_9110);
nand U10614 (N_10614,N_7262,N_8863);
and U10615 (N_10615,N_8788,N_6459);
nor U10616 (N_10616,N_8135,N_8945);
nor U10617 (N_10617,N_7177,N_8518);
or U10618 (N_10618,N_8156,N_7933);
xor U10619 (N_10619,N_8079,N_8020);
nor U10620 (N_10620,N_7677,N_8220);
nor U10621 (N_10621,N_9139,N_8988);
nand U10622 (N_10622,N_6962,N_8667);
nor U10623 (N_10623,N_6463,N_6631);
or U10624 (N_10624,N_7349,N_6519);
and U10625 (N_10625,N_7194,N_6642);
and U10626 (N_10626,N_8680,N_7135);
and U10627 (N_10627,N_7180,N_7356);
nor U10628 (N_10628,N_6311,N_7322);
xor U10629 (N_10629,N_7541,N_7462);
or U10630 (N_10630,N_7074,N_7410);
or U10631 (N_10631,N_6758,N_7567);
or U10632 (N_10632,N_6801,N_8351);
nand U10633 (N_10633,N_8976,N_6650);
nor U10634 (N_10634,N_6388,N_6872);
nor U10635 (N_10635,N_8258,N_7945);
nand U10636 (N_10636,N_9061,N_8309);
or U10637 (N_10637,N_6709,N_8899);
or U10638 (N_10638,N_8627,N_6771);
nor U10639 (N_10639,N_8734,N_9022);
or U10640 (N_10640,N_7956,N_7732);
or U10641 (N_10641,N_8901,N_6909);
or U10642 (N_10642,N_7573,N_6813);
or U10643 (N_10643,N_6757,N_7489);
nor U10644 (N_10644,N_8550,N_7066);
nand U10645 (N_10645,N_8687,N_6865);
and U10646 (N_10646,N_7657,N_7063);
and U10647 (N_10647,N_8055,N_7738);
nor U10648 (N_10648,N_8138,N_7072);
nand U10649 (N_10649,N_9319,N_8743);
nand U10650 (N_10650,N_9017,N_7017);
xnor U10651 (N_10651,N_7365,N_6744);
or U10652 (N_10652,N_7896,N_6251);
or U10653 (N_10653,N_7723,N_6372);
xor U10654 (N_10654,N_6837,N_7996);
nand U10655 (N_10655,N_9031,N_6433);
nor U10656 (N_10656,N_6613,N_6564);
nor U10657 (N_10657,N_8013,N_9038);
nand U10658 (N_10658,N_9294,N_8421);
nand U10659 (N_10659,N_7301,N_9348);
and U10660 (N_10660,N_7883,N_9353);
nand U10661 (N_10661,N_7521,N_8585);
nand U10662 (N_10662,N_6779,N_8959);
nand U10663 (N_10663,N_6692,N_8630);
nand U10664 (N_10664,N_7869,N_8917);
nor U10665 (N_10665,N_6666,N_7611);
xnor U10666 (N_10666,N_8916,N_6778);
and U10667 (N_10667,N_8919,N_6729);
and U10668 (N_10668,N_8471,N_8170);
nand U10669 (N_10669,N_9221,N_7030);
and U10670 (N_10670,N_7087,N_8487);
nor U10671 (N_10671,N_9368,N_7374);
or U10672 (N_10672,N_7612,N_8204);
and U10673 (N_10673,N_7504,N_7055);
xor U10674 (N_10674,N_8368,N_7480);
nor U10675 (N_10675,N_9213,N_9130);
and U10676 (N_10676,N_8007,N_9296);
nand U10677 (N_10677,N_6302,N_8229);
or U10678 (N_10678,N_8871,N_8394);
or U10679 (N_10679,N_8715,N_8115);
and U10680 (N_10680,N_7445,N_7716);
or U10681 (N_10681,N_6862,N_7297);
nand U10682 (N_10682,N_9001,N_9028);
or U10683 (N_10683,N_8506,N_8552);
and U10684 (N_10684,N_7463,N_8340);
and U10685 (N_10685,N_9256,N_8491);
nand U10686 (N_10686,N_8538,N_9024);
xor U10687 (N_10687,N_8106,N_8944);
and U10688 (N_10688,N_8445,N_8259);
or U10689 (N_10689,N_7361,N_7624);
nor U10690 (N_10690,N_8498,N_7239);
nand U10691 (N_10691,N_8101,N_7173);
xor U10692 (N_10692,N_7682,N_8356);
and U10693 (N_10693,N_6997,N_7179);
xnor U10694 (N_10694,N_6436,N_6930);
nor U10695 (N_10695,N_6979,N_6767);
nor U10696 (N_10696,N_8576,N_6850);
nor U10697 (N_10697,N_8639,N_8882);
nor U10698 (N_10698,N_6833,N_7353);
nor U10699 (N_10699,N_8226,N_9137);
or U10700 (N_10700,N_7047,N_7319);
xor U10701 (N_10701,N_8292,N_9335);
and U10702 (N_10702,N_9281,N_6647);
xor U10703 (N_10703,N_7359,N_6252);
nor U10704 (N_10704,N_9211,N_7498);
nand U10705 (N_10705,N_8213,N_7771);
and U10706 (N_10706,N_7571,N_7391);
nand U10707 (N_10707,N_7663,N_8069);
nand U10708 (N_10708,N_6394,N_9300);
and U10709 (N_10709,N_6306,N_9151);
or U10710 (N_10710,N_6554,N_7981);
nor U10711 (N_10711,N_8853,N_7041);
nor U10712 (N_10712,N_8310,N_7490);
nor U10713 (N_10713,N_7460,N_6377);
and U10714 (N_10714,N_6936,N_8674);
nor U10715 (N_10715,N_7012,N_7900);
nand U10716 (N_10716,N_7324,N_9239);
and U10717 (N_10717,N_8162,N_7242);
nand U10718 (N_10718,N_6448,N_9184);
nor U10719 (N_10719,N_8771,N_6652);
nor U10720 (N_10720,N_7651,N_6255);
nor U10721 (N_10721,N_8990,N_9252);
or U10722 (N_10722,N_7913,N_9219);
and U10723 (N_10723,N_7807,N_8584);
and U10724 (N_10724,N_8593,N_9284);
nor U10725 (N_10725,N_8607,N_7994);
and U10726 (N_10726,N_7108,N_7025);
xnor U10727 (N_10727,N_9231,N_6878);
or U10728 (N_10728,N_6518,N_6557);
xnor U10729 (N_10729,N_7225,N_9338);
nand U10730 (N_10730,N_8128,N_8693);
or U10731 (N_10731,N_7192,N_8454);
or U10732 (N_10732,N_6977,N_8840);
or U10733 (N_10733,N_7868,N_6684);
and U10734 (N_10734,N_8588,N_7132);
nand U10735 (N_10735,N_7523,N_7076);
and U10736 (N_10736,N_7666,N_7292);
nand U10737 (N_10737,N_7009,N_7080);
and U10738 (N_10738,N_7099,N_6425);
xnor U10739 (N_10739,N_6561,N_7978);
nand U10740 (N_10740,N_8361,N_7982);
nor U10741 (N_10741,N_6344,N_9062);
or U10742 (N_10742,N_8410,N_7211);
or U10743 (N_10743,N_8723,N_6254);
or U10744 (N_10744,N_8051,N_6521);
and U10745 (N_10745,N_8568,N_9053);
nor U10746 (N_10746,N_8969,N_6263);
nand U10747 (N_10747,N_9199,N_8130);
nor U10748 (N_10748,N_7443,N_9232);
nand U10749 (N_10749,N_8303,N_8288);
or U10750 (N_10750,N_6664,N_6976);
and U10751 (N_10751,N_6790,N_6753);
xnor U10752 (N_10752,N_7821,N_7520);
or U10753 (N_10753,N_8419,N_7188);
nand U10754 (N_10754,N_6282,N_8545);
xor U10755 (N_10755,N_8267,N_8467);
or U10756 (N_10756,N_6288,N_6818);
nand U10757 (N_10757,N_8704,N_8563);
and U10758 (N_10758,N_9190,N_8084);
nor U10759 (N_10759,N_9009,N_7619);
nor U10760 (N_10760,N_6256,N_6285);
and U10761 (N_10761,N_8730,N_7222);
and U10762 (N_10762,N_8697,N_8886);
or U10763 (N_10763,N_8155,N_7082);
or U10764 (N_10764,N_7650,N_6759);
or U10765 (N_10765,N_7424,N_6615);
or U10766 (N_10766,N_8320,N_7394);
and U10767 (N_10767,N_8385,N_9217);
nand U10768 (N_10768,N_7961,N_7399);
or U10769 (N_10769,N_7708,N_6969);
and U10770 (N_10770,N_8028,N_8686);
nand U10771 (N_10771,N_7928,N_9364);
or U10772 (N_10772,N_6308,N_8536);
or U10773 (N_10773,N_6384,N_7705);
or U10774 (N_10774,N_7741,N_8346);
xnor U10775 (N_10775,N_7641,N_7922);
and U10776 (N_10776,N_7742,N_8178);
nand U10777 (N_10777,N_8909,N_7006);
nand U10778 (N_10778,N_7441,N_8869);
or U10779 (N_10779,N_7727,N_6946);
nand U10780 (N_10780,N_8720,N_8731);
xor U10781 (N_10781,N_9056,N_6688);
or U10782 (N_10782,N_8380,N_6868);
or U10783 (N_10783,N_6526,N_9285);
nor U10784 (N_10784,N_7339,N_6435);
xnor U10785 (N_10785,N_7768,N_8164);
or U10786 (N_10786,N_6612,N_7980);
nor U10787 (N_10787,N_8826,N_7196);
nand U10788 (N_10788,N_8949,N_6860);
and U10789 (N_10789,N_9188,N_8062);
nand U10790 (N_10790,N_7294,N_8570);
xor U10791 (N_10791,N_7899,N_6895);
or U10792 (N_10792,N_8371,N_7492);
nand U10793 (N_10793,N_9014,N_6452);
nor U10794 (N_10794,N_7779,N_7079);
nand U10795 (N_10795,N_6387,N_7278);
nand U10796 (N_10796,N_7593,N_8750);
nand U10797 (N_10797,N_8194,N_8946);
nand U10798 (N_10798,N_8474,N_7021);
or U10799 (N_10799,N_6559,N_9141);
and U10800 (N_10800,N_8927,N_8725);
or U10801 (N_10801,N_7743,N_9237);
nor U10802 (N_10802,N_7745,N_6927);
nand U10803 (N_10803,N_7722,N_8463);
nor U10804 (N_10804,N_6785,N_8890);
or U10805 (N_10805,N_8532,N_9289);
nand U10806 (N_10806,N_8472,N_7111);
or U10807 (N_10807,N_9327,N_8242);
nand U10808 (N_10808,N_7090,N_7915);
xor U10809 (N_10809,N_6279,N_6900);
and U10810 (N_10810,N_8295,N_6830);
nor U10811 (N_10811,N_7778,N_9064);
or U10812 (N_10812,N_9318,N_7553);
or U10813 (N_10813,N_6727,N_7193);
nand U10814 (N_10814,N_8640,N_7060);
or U10815 (N_10815,N_8379,N_7940);
nand U10816 (N_10816,N_7714,N_7133);
nand U10817 (N_10817,N_8219,N_8789);
nand U10818 (N_10818,N_8892,N_7020);
nand U10819 (N_10819,N_8528,N_6342);
or U10820 (N_10820,N_7628,N_6382);
nor U10821 (N_10821,N_9037,N_7237);
nor U10822 (N_10822,N_8021,N_7583);
and U10823 (N_10823,N_7510,N_8113);
nor U10824 (N_10824,N_8850,N_8767);
or U10825 (N_10825,N_9248,N_8217);
xor U10826 (N_10826,N_8824,N_8589);
or U10827 (N_10827,N_6587,N_7524);
nand U10828 (N_10828,N_8089,N_7230);
nor U10829 (N_10829,N_6871,N_8157);
and U10830 (N_10830,N_6327,N_7251);
or U10831 (N_10831,N_7052,N_6597);
xnor U10832 (N_10832,N_7023,N_8645);
and U10833 (N_10833,N_8755,N_7843);
nor U10834 (N_10834,N_7988,N_7217);
and U10835 (N_10835,N_8271,N_7599);
nand U10836 (N_10836,N_6607,N_9314);
or U10837 (N_10837,N_7098,N_9363);
nand U10838 (N_10838,N_8841,N_7474);
or U10839 (N_10839,N_8875,N_8386);
or U10840 (N_10840,N_7103,N_7130);
or U10841 (N_10841,N_9084,N_7050);
nor U10842 (N_10842,N_7671,N_9015);
or U10843 (N_10843,N_6609,N_7644);
xor U10844 (N_10844,N_8045,N_8446);
or U10845 (N_10845,N_6637,N_8866);
and U10846 (N_10846,N_9164,N_8207);
and U10847 (N_10847,N_9241,N_7158);
nand U10848 (N_10848,N_8569,N_7338);
and U10849 (N_10849,N_9276,N_7004);
and U10850 (N_10850,N_6268,N_7390);
or U10851 (N_10851,N_9105,N_9154);
nand U10852 (N_10852,N_6422,N_7335);
nor U10853 (N_10853,N_8691,N_8913);
or U10854 (N_10854,N_8256,N_7244);
nand U10855 (N_10855,N_8800,N_7423);
or U10856 (N_10856,N_8308,N_8833);
nand U10857 (N_10857,N_6839,N_7548);
nor U10858 (N_10858,N_9025,N_7709);
or U10859 (N_10859,N_7934,N_7002);
nand U10860 (N_10860,N_8502,N_7579);
or U10861 (N_10861,N_7508,N_7793);
nor U10862 (N_10862,N_7797,N_8675);
xor U10863 (N_10863,N_8152,N_8902);
and U10864 (N_10864,N_8116,N_6595);
and U10865 (N_10865,N_6392,N_7697);
nor U10866 (N_10866,N_6395,N_8700);
and U10867 (N_10867,N_6502,N_6792);
and U10868 (N_10868,N_7044,N_9172);
xnor U10869 (N_10869,N_6522,N_8496);
or U10870 (N_10870,N_8759,N_8672);
and U10871 (N_10871,N_7334,N_6745);
or U10872 (N_10872,N_7357,N_7081);
nand U10873 (N_10873,N_6803,N_7603);
nand U10874 (N_10874,N_7512,N_6414);
and U10875 (N_10875,N_8984,N_8517);
or U10876 (N_10876,N_7277,N_7413);
or U10877 (N_10877,N_8727,N_7865);
or U10878 (N_10878,N_8050,N_7856);
or U10879 (N_10879,N_8655,N_9026);
xnor U10880 (N_10880,N_6379,N_8470);
xnor U10881 (N_10881,N_9352,N_7902);
or U10882 (N_10882,N_9136,N_7854);
and U10883 (N_10883,N_8848,N_8302);
nor U10884 (N_10884,N_6485,N_7221);
nand U10885 (N_10885,N_6619,N_6358);
nand U10886 (N_10886,N_7269,N_9236);
and U10887 (N_10887,N_7777,N_7942);
and U10888 (N_10888,N_8298,N_9152);
nor U10889 (N_10889,N_8442,N_6357);
and U10890 (N_10890,N_7962,N_7559);
and U10891 (N_10891,N_9251,N_8358);
xor U10892 (N_10892,N_6999,N_7351);
nor U10893 (N_10893,N_7477,N_6611);
or U10894 (N_10894,N_6912,N_7975);
and U10895 (N_10895,N_6852,N_8937);
or U10896 (N_10896,N_9180,N_9156);
or U10897 (N_10897,N_8480,N_8359);
or U10898 (N_10898,N_8718,N_6776);
or U10899 (N_10899,N_6267,N_9005);
or U10900 (N_10900,N_7458,N_7062);
xor U10901 (N_10901,N_7015,N_9179);
and U10902 (N_10902,N_7632,N_8950);
nand U10903 (N_10903,N_7139,N_8266);
nand U10904 (N_10904,N_8306,N_7562);
and U10905 (N_10905,N_9307,N_6820);
nor U10906 (N_10906,N_7497,N_8107);
or U10907 (N_10907,N_8129,N_8058);
nor U10908 (N_10908,N_6594,N_8910);
nand U10909 (N_10909,N_8344,N_7584);
and U10910 (N_10910,N_6332,N_8989);
nand U10911 (N_10911,N_8067,N_8952);
nand U10912 (N_10912,N_7639,N_8455);
or U10913 (N_10913,N_6851,N_8090);
and U10914 (N_10914,N_6786,N_6735);
or U10915 (N_10915,N_8251,N_7005);
nand U10916 (N_10916,N_6942,N_9146);
nor U10917 (N_10917,N_6736,N_6265);
and U10918 (N_10918,N_8772,N_7637);
nand U10919 (N_10919,N_8938,N_6633);
or U10920 (N_10920,N_8305,N_7372);
or U10921 (N_10921,N_7426,N_9240);
or U10922 (N_10922,N_9333,N_8629);
nand U10923 (N_10923,N_9202,N_6799);
and U10924 (N_10924,N_7780,N_6460);
and U10925 (N_10925,N_7830,N_7668);
and U10926 (N_10926,N_6287,N_8710);
or U10927 (N_10927,N_9153,N_7053);
nor U10928 (N_10928,N_7674,N_8994);
nor U10929 (N_10929,N_6660,N_8933);
nor U10930 (N_10930,N_8488,N_6891);
and U10931 (N_10931,N_7638,N_6682);
nor U10932 (N_10932,N_9004,N_8384);
nor U10933 (N_10933,N_6680,N_6941);
xor U10934 (N_10934,N_9282,N_7118);
xnor U10935 (N_10935,N_7197,N_6451);
nand U10936 (N_10936,N_7690,N_9247);
nand U10937 (N_10937,N_8796,N_9180);
or U10938 (N_10938,N_8437,N_7338);
and U10939 (N_10939,N_6262,N_7818);
nand U10940 (N_10940,N_7968,N_8848);
nand U10941 (N_10941,N_8522,N_6643);
nand U10942 (N_10942,N_7624,N_8727);
nor U10943 (N_10943,N_6915,N_7376);
and U10944 (N_10944,N_7594,N_7223);
nand U10945 (N_10945,N_8380,N_7533);
xnor U10946 (N_10946,N_6428,N_6664);
nor U10947 (N_10947,N_6894,N_8871);
and U10948 (N_10948,N_8374,N_7250);
or U10949 (N_10949,N_7269,N_8241);
or U10950 (N_10950,N_6667,N_7088);
nand U10951 (N_10951,N_8780,N_8067);
nand U10952 (N_10952,N_8931,N_6546);
nand U10953 (N_10953,N_8915,N_8244);
or U10954 (N_10954,N_7412,N_8147);
or U10955 (N_10955,N_9176,N_6983);
and U10956 (N_10956,N_8358,N_7762);
or U10957 (N_10957,N_9276,N_6352);
xor U10958 (N_10958,N_7536,N_7660);
nor U10959 (N_10959,N_9316,N_7620);
nor U10960 (N_10960,N_6396,N_6658);
or U10961 (N_10961,N_8666,N_6831);
and U10962 (N_10962,N_8210,N_6349);
nor U10963 (N_10963,N_6408,N_7135);
or U10964 (N_10964,N_7804,N_7810);
and U10965 (N_10965,N_6610,N_7770);
or U10966 (N_10966,N_6318,N_9240);
or U10967 (N_10967,N_8015,N_8788);
nand U10968 (N_10968,N_7483,N_6697);
and U10969 (N_10969,N_9039,N_9129);
nand U10970 (N_10970,N_8213,N_6378);
nand U10971 (N_10971,N_7053,N_8701);
and U10972 (N_10972,N_8514,N_7168);
nor U10973 (N_10973,N_9168,N_6909);
nor U10974 (N_10974,N_7257,N_6523);
nand U10975 (N_10975,N_8393,N_7721);
and U10976 (N_10976,N_7561,N_7118);
and U10977 (N_10977,N_8059,N_8537);
nand U10978 (N_10978,N_6537,N_8917);
nand U10979 (N_10979,N_7794,N_7824);
and U10980 (N_10980,N_7651,N_7925);
and U10981 (N_10981,N_8484,N_9318);
nand U10982 (N_10982,N_8293,N_7205);
or U10983 (N_10983,N_6407,N_8585);
and U10984 (N_10984,N_9074,N_6934);
and U10985 (N_10985,N_6656,N_8290);
xnor U10986 (N_10986,N_9144,N_7560);
and U10987 (N_10987,N_8025,N_8289);
or U10988 (N_10988,N_8849,N_8363);
nand U10989 (N_10989,N_8739,N_8417);
nor U10990 (N_10990,N_8082,N_8811);
nand U10991 (N_10991,N_9050,N_8206);
nor U10992 (N_10992,N_6737,N_6844);
and U10993 (N_10993,N_6279,N_9162);
nand U10994 (N_10994,N_8230,N_8603);
nand U10995 (N_10995,N_6917,N_8562);
and U10996 (N_10996,N_6613,N_7319);
nand U10997 (N_10997,N_9096,N_8919);
or U10998 (N_10998,N_9303,N_9032);
and U10999 (N_10999,N_7490,N_8487);
nand U11000 (N_11000,N_8565,N_9066);
nand U11001 (N_11001,N_9129,N_6257);
nand U11002 (N_11002,N_7059,N_7821);
or U11003 (N_11003,N_7389,N_7946);
and U11004 (N_11004,N_8383,N_6427);
nand U11005 (N_11005,N_6581,N_7477);
or U11006 (N_11006,N_8058,N_6503);
nand U11007 (N_11007,N_9193,N_9358);
or U11008 (N_11008,N_7080,N_8471);
xnor U11009 (N_11009,N_8433,N_8947);
and U11010 (N_11010,N_7236,N_9079);
or U11011 (N_11011,N_8552,N_7534);
and U11012 (N_11012,N_7257,N_8800);
and U11013 (N_11013,N_8609,N_6447);
or U11014 (N_11014,N_8251,N_7073);
nand U11015 (N_11015,N_7313,N_6850);
or U11016 (N_11016,N_7179,N_9335);
and U11017 (N_11017,N_8874,N_7566);
nor U11018 (N_11018,N_9338,N_8055);
nand U11019 (N_11019,N_8388,N_8482);
and U11020 (N_11020,N_6615,N_8189);
nand U11021 (N_11021,N_7564,N_6709);
nor U11022 (N_11022,N_8359,N_6305);
nor U11023 (N_11023,N_8063,N_6470);
and U11024 (N_11024,N_9141,N_6383);
or U11025 (N_11025,N_6496,N_7307);
or U11026 (N_11026,N_6857,N_7894);
or U11027 (N_11027,N_7940,N_8663);
and U11028 (N_11028,N_9339,N_8799);
or U11029 (N_11029,N_6640,N_6265);
nor U11030 (N_11030,N_6896,N_8754);
nor U11031 (N_11031,N_6859,N_6675);
or U11032 (N_11032,N_9326,N_7436);
or U11033 (N_11033,N_7041,N_8640);
and U11034 (N_11034,N_8938,N_7386);
xnor U11035 (N_11035,N_7030,N_6747);
nand U11036 (N_11036,N_7672,N_6513);
or U11037 (N_11037,N_8910,N_6963);
xor U11038 (N_11038,N_7527,N_7957);
nor U11039 (N_11039,N_9073,N_6539);
xnor U11040 (N_11040,N_8623,N_6593);
and U11041 (N_11041,N_9082,N_7643);
nor U11042 (N_11042,N_7784,N_8518);
nand U11043 (N_11043,N_8670,N_7522);
or U11044 (N_11044,N_9373,N_6693);
and U11045 (N_11045,N_6560,N_7313);
xnor U11046 (N_11046,N_7797,N_9165);
nand U11047 (N_11047,N_7062,N_8951);
nand U11048 (N_11048,N_8307,N_8450);
or U11049 (N_11049,N_8340,N_9146);
or U11050 (N_11050,N_8229,N_8224);
nand U11051 (N_11051,N_8148,N_7697);
or U11052 (N_11052,N_6293,N_6584);
nand U11053 (N_11053,N_7857,N_7028);
nor U11054 (N_11054,N_7468,N_9351);
or U11055 (N_11055,N_8290,N_6840);
and U11056 (N_11056,N_8698,N_8707);
or U11057 (N_11057,N_6599,N_9196);
xor U11058 (N_11058,N_6971,N_8313);
nor U11059 (N_11059,N_8003,N_8198);
or U11060 (N_11060,N_6253,N_8040);
nor U11061 (N_11061,N_9031,N_8801);
or U11062 (N_11062,N_7810,N_9043);
or U11063 (N_11063,N_9221,N_8145);
nor U11064 (N_11064,N_6977,N_9164);
nand U11065 (N_11065,N_8897,N_6840);
nor U11066 (N_11066,N_7333,N_7846);
nor U11067 (N_11067,N_8792,N_8161);
or U11068 (N_11068,N_7117,N_9335);
xnor U11069 (N_11069,N_7717,N_7710);
nor U11070 (N_11070,N_8871,N_7779);
and U11071 (N_11071,N_8385,N_8874);
nand U11072 (N_11072,N_6508,N_9272);
and U11073 (N_11073,N_8307,N_7848);
or U11074 (N_11074,N_8190,N_8146);
nand U11075 (N_11075,N_8257,N_8381);
nor U11076 (N_11076,N_7063,N_7507);
nand U11077 (N_11077,N_7468,N_9022);
nor U11078 (N_11078,N_7158,N_6352);
nor U11079 (N_11079,N_9252,N_6978);
or U11080 (N_11080,N_9106,N_8436);
nand U11081 (N_11081,N_7629,N_6385);
nor U11082 (N_11082,N_9119,N_6821);
nand U11083 (N_11083,N_8526,N_6309);
nand U11084 (N_11084,N_8724,N_6773);
or U11085 (N_11085,N_8518,N_9058);
nor U11086 (N_11086,N_8838,N_8431);
nand U11087 (N_11087,N_9117,N_6405);
nand U11088 (N_11088,N_6889,N_6271);
and U11089 (N_11089,N_8686,N_7499);
nor U11090 (N_11090,N_8017,N_8224);
nand U11091 (N_11091,N_8348,N_8340);
or U11092 (N_11092,N_8102,N_7525);
and U11093 (N_11093,N_6834,N_7450);
xnor U11094 (N_11094,N_8119,N_6876);
and U11095 (N_11095,N_8927,N_8970);
and U11096 (N_11096,N_8869,N_7133);
nor U11097 (N_11097,N_7541,N_8062);
xnor U11098 (N_11098,N_8237,N_7328);
or U11099 (N_11099,N_8392,N_7105);
nand U11100 (N_11100,N_7382,N_8778);
nand U11101 (N_11101,N_8895,N_7709);
nor U11102 (N_11102,N_6855,N_8104);
nand U11103 (N_11103,N_6291,N_6825);
and U11104 (N_11104,N_8204,N_6727);
nand U11105 (N_11105,N_9109,N_6871);
and U11106 (N_11106,N_7527,N_8599);
xor U11107 (N_11107,N_6858,N_7079);
nand U11108 (N_11108,N_7359,N_8932);
and U11109 (N_11109,N_6774,N_6692);
nand U11110 (N_11110,N_8021,N_7396);
nor U11111 (N_11111,N_9054,N_6745);
or U11112 (N_11112,N_7775,N_6925);
nor U11113 (N_11113,N_7332,N_8583);
or U11114 (N_11114,N_6808,N_8337);
nand U11115 (N_11115,N_8788,N_6327);
nand U11116 (N_11116,N_8351,N_7970);
nand U11117 (N_11117,N_7520,N_6523);
nand U11118 (N_11118,N_6367,N_7010);
nor U11119 (N_11119,N_8176,N_7324);
and U11120 (N_11120,N_9191,N_7654);
nor U11121 (N_11121,N_7738,N_6696);
nand U11122 (N_11122,N_7837,N_7726);
nor U11123 (N_11123,N_8068,N_8580);
or U11124 (N_11124,N_8192,N_7899);
or U11125 (N_11125,N_7744,N_7042);
nor U11126 (N_11126,N_7210,N_7492);
nand U11127 (N_11127,N_8030,N_6355);
nand U11128 (N_11128,N_8634,N_8588);
and U11129 (N_11129,N_7374,N_7290);
xnor U11130 (N_11130,N_6916,N_9273);
or U11131 (N_11131,N_6516,N_8821);
nand U11132 (N_11132,N_8123,N_6620);
or U11133 (N_11133,N_8765,N_8013);
and U11134 (N_11134,N_7143,N_8932);
or U11135 (N_11135,N_8710,N_9370);
and U11136 (N_11136,N_7832,N_8467);
nor U11137 (N_11137,N_8486,N_9066);
or U11138 (N_11138,N_7432,N_7282);
nand U11139 (N_11139,N_8821,N_8496);
nand U11140 (N_11140,N_8880,N_7480);
nor U11141 (N_11141,N_9360,N_6917);
or U11142 (N_11142,N_8618,N_7346);
and U11143 (N_11143,N_6374,N_8554);
and U11144 (N_11144,N_8141,N_9173);
nor U11145 (N_11145,N_8488,N_9291);
and U11146 (N_11146,N_8633,N_6566);
xnor U11147 (N_11147,N_7192,N_6836);
and U11148 (N_11148,N_8920,N_9314);
nor U11149 (N_11149,N_8853,N_8034);
or U11150 (N_11150,N_6467,N_9181);
xnor U11151 (N_11151,N_6643,N_6348);
nand U11152 (N_11152,N_9326,N_9028);
nor U11153 (N_11153,N_7127,N_7497);
xnor U11154 (N_11154,N_6497,N_8019);
nand U11155 (N_11155,N_6819,N_8436);
nand U11156 (N_11156,N_6710,N_7488);
xor U11157 (N_11157,N_8814,N_7591);
nand U11158 (N_11158,N_9190,N_6432);
xnor U11159 (N_11159,N_7315,N_8080);
or U11160 (N_11160,N_7108,N_6341);
nor U11161 (N_11161,N_7423,N_8005);
nor U11162 (N_11162,N_6377,N_8436);
or U11163 (N_11163,N_7587,N_6977);
or U11164 (N_11164,N_9083,N_7109);
nand U11165 (N_11165,N_7181,N_9156);
or U11166 (N_11166,N_8472,N_8110);
nand U11167 (N_11167,N_8861,N_8748);
nand U11168 (N_11168,N_9045,N_7854);
nand U11169 (N_11169,N_8362,N_6522);
nand U11170 (N_11170,N_6307,N_6304);
and U11171 (N_11171,N_8900,N_7313);
or U11172 (N_11172,N_8375,N_7153);
nand U11173 (N_11173,N_6888,N_9032);
nor U11174 (N_11174,N_7352,N_6547);
or U11175 (N_11175,N_7260,N_6526);
xnor U11176 (N_11176,N_7238,N_6878);
nor U11177 (N_11177,N_6541,N_9343);
nor U11178 (N_11178,N_9156,N_7006);
nand U11179 (N_11179,N_8261,N_9258);
and U11180 (N_11180,N_6429,N_6298);
and U11181 (N_11181,N_6713,N_9342);
and U11182 (N_11182,N_7957,N_7416);
nand U11183 (N_11183,N_9009,N_7479);
or U11184 (N_11184,N_7773,N_7104);
nand U11185 (N_11185,N_7150,N_7060);
nor U11186 (N_11186,N_6963,N_8261);
nand U11187 (N_11187,N_6742,N_6518);
nor U11188 (N_11188,N_7773,N_6495);
nand U11189 (N_11189,N_6633,N_7662);
or U11190 (N_11190,N_8057,N_8490);
nand U11191 (N_11191,N_7387,N_9364);
xnor U11192 (N_11192,N_8819,N_8954);
or U11193 (N_11193,N_7579,N_6971);
or U11194 (N_11194,N_9180,N_8958);
nand U11195 (N_11195,N_8557,N_6990);
or U11196 (N_11196,N_8988,N_9270);
nand U11197 (N_11197,N_7015,N_6822);
nor U11198 (N_11198,N_8496,N_6650);
nor U11199 (N_11199,N_9351,N_9211);
and U11200 (N_11200,N_7758,N_7901);
nand U11201 (N_11201,N_8687,N_6678);
nor U11202 (N_11202,N_6353,N_6590);
and U11203 (N_11203,N_8044,N_7812);
and U11204 (N_11204,N_9360,N_8106);
nand U11205 (N_11205,N_6897,N_8361);
nand U11206 (N_11206,N_6407,N_6809);
xnor U11207 (N_11207,N_8283,N_7381);
nor U11208 (N_11208,N_7274,N_8736);
nand U11209 (N_11209,N_9356,N_6936);
nand U11210 (N_11210,N_7306,N_6501);
and U11211 (N_11211,N_7779,N_7939);
xnor U11212 (N_11212,N_7308,N_6955);
and U11213 (N_11213,N_6481,N_7997);
and U11214 (N_11214,N_8421,N_6713);
or U11215 (N_11215,N_6849,N_8054);
or U11216 (N_11216,N_6266,N_7877);
nor U11217 (N_11217,N_7602,N_7332);
nand U11218 (N_11218,N_8073,N_8266);
or U11219 (N_11219,N_6917,N_9278);
and U11220 (N_11220,N_9000,N_7522);
xnor U11221 (N_11221,N_7923,N_6965);
nand U11222 (N_11222,N_7818,N_6701);
nor U11223 (N_11223,N_6818,N_7401);
or U11224 (N_11224,N_6662,N_7737);
nand U11225 (N_11225,N_9309,N_8102);
xor U11226 (N_11226,N_7169,N_6990);
or U11227 (N_11227,N_6652,N_8967);
xor U11228 (N_11228,N_8053,N_8133);
nand U11229 (N_11229,N_7156,N_6663);
nor U11230 (N_11230,N_7630,N_6909);
xnor U11231 (N_11231,N_8606,N_8482);
xor U11232 (N_11232,N_7720,N_9348);
and U11233 (N_11233,N_9133,N_8750);
and U11234 (N_11234,N_7652,N_8777);
nand U11235 (N_11235,N_7289,N_6335);
nor U11236 (N_11236,N_7928,N_8098);
or U11237 (N_11237,N_6474,N_6725);
xor U11238 (N_11238,N_9087,N_8870);
and U11239 (N_11239,N_7343,N_7118);
xor U11240 (N_11240,N_8065,N_8400);
nor U11241 (N_11241,N_8590,N_6329);
or U11242 (N_11242,N_7347,N_6926);
or U11243 (N_11243,N_9366,N_6586);
or U11244 (N_11244,N_7174,N_7707);
or U11245 (N_11245,N_9076,N_8292);
nand U11246 (N_11246,N_6683,N_8016);
nor U11247 (N_11247,N_8117,N_6735);
or U11248 (N_11248,N_8260,N_7686);
nand U11249 (N_11249,N_7678,N_7847);
xor U11250 (N_11250,N_9096,N_6733);
and U11251 (N_11251,N_7915,N_7776);
nand U11252 (N_11252,N_8728,N_8761);
nand U11253 (N_11253,N_6608,N_6372);
and U11254 (N_11254,N_8927,N_8374);
or U11255 (N_11255,N_8234,N_7319);
and U11256 (N_11256,N_8065,N_8835);
nor U11257 (N_11257,N_6262,N_9311);
and U11258 (N_11258,N_9068,N_6309);
or U11259 (N_11259,N_8631,N_7424);
xor U11260 (N_11260,N_6268,N_9199);
nor U11261 (N_11261,N_6577,N_7101);
xnor U11262 (N_11262,N_6460,N_8871);
nor U11263 (N_11263,N_8857,N_9340);
or U11264 (N_11264,N_7160,N_8323);
nor U11265 (N_11265,N_7192,N_7893);
and U11266 (N_11266,N_9344,N_8979);
nand U11267 (N_11267,N_7053,N_8405);
nand U11268 (N_11268,N_7944,N_8437);
nand U11269 (N_11269,N_7826,N_9331);
or U11270 (N_11270,N_6781,N_6686);
and U11271 (N_11271,N_6425,N_7376);
nor U11272 (N_11272,N_7605,N_8506);
xnor U11273 (N_11273,N_9048,N_6699);
nand U11274 (N_11274,N_9293,N_7441);
nand U11275 (N_11275,N_8016,N_8795);
and U11276 (N_11276,N_6258,N_7764);
nor U11277 (N_11277,N_7642,N_7486);
nand U11278 (N_11278,N_6623,N_7538);
nand U11279 (N_11279,N_6301,N_7227);
xnor U11280 (N_11280,N_8681,N_8648);
and U11281 (N_11281,N_6639,N_6792);
xor U11282 (N_11282,N_6570,N_7925);
or U11283 (N_11283,N_6537,N_8109);
or U11284 (N_11284,N_7837,N_6835);
nor U11285 (N_11285,N_8360,N_7439);
or U11286 (N_11286,N_8081,N_9054);
and U11287 (N_11287,N_6915,N_8371);
nor U11288 (N_11288,N_8828,N_8609);
nor U11289 (N_11289,N_6973,N_7176);
nand U11290 (N_11290,N_9025,N_6724);
or U11291 (N_11291,N_7082,N_6561);
or U11292 (N_11292,N_7866,N_7943);
nor U11293 (N_11293,N_6422,N_6332);
nor U11294 (N_11294,N_8068,N_7743);
nand U11295 (N_11295,N_8774,N_9233);
xnor U11296 (N_11296,N_7607,N_8600);
and U11297 (N_11297,N_7819,N_8212);
and U11298 (N_11298,N_7881,N_9322);
or U11299 (N_11299,N_7279,N_6388);
and U11300 (N_11300,N_7664,N_7418);
nor U11301 (N_11301,N_8796,N_6405);
nor U11302 (N_11302,N_9358,N_9204);
and U11303 (N_11303,N_6621,N_6990);
and U11304 (N_11304,N_8317,N_7209);
nor U11305 (N_11305,N_6393,N_8895);
nand U11306 (N_11306,N_8971,N_7752);
and U11307 (N_11307,N_8601,N_6285);
nand U11308 (N_11308,N_6947,N_6778);
nor U11309 (N_11309,N_6554,N_8349);
nand U11310 (N_11310,N_9282,N_8847);
nor U11311 (N_11311,N_6277,N_7342);
nor U11312 (N_11312,N_7473,N_8610);
nor U11313 (N_11313,N_6833,N_7996);
and U11314 (N_11314,N_7595,N_7801);
nand U11315 (N_11315,N_6781,N_6649);
nor U11316 (N_11316,N_7093,N_8129);
nor U11317 (N_11317,N_7011,N_7373);
nand U11318 (N_11318,N_7581,N_9008);
nor U11319 (N_11319,N_6802,N_7643);
nor U11320 (N_11320,N_7751,N_8728);
or U11321 (N_11321,N_9231,N_8675);
and U11322 (N_11322,N_8637,N_8669);
or U11323 (N_11323,N_6725,N_6479);
and U11324 (N_11324,N_7131,N_8399);
and U11325 (N_11325,N_6529,N_7228);
and U11326 (N_11326,N_8899,N_6897);
nand U11327 (N_11327,N_9343,N_6840);
and U11328 (N_11328,N_9129,N_7667);
or U11329 (N_11329,N_9197,N_6376);
or U11330 (N_11330,N_8295,N_8476);
nand U11331 (N_11331,N_6559,N_7106);
and U11332 (N_11332,N_8629,N_7484);
and U11333 (N_11333,N_6592,N_8905);
nand U11334 (N_11334,N_8135,N_7090);
nand U11335 (N_11335,N_6726,N_7218);
and U11336 (N_11336,N_9169,N_6947);
nand U11337 (N_11337,N_7481,N_9334);
nand U11338 (N_11338,N_7340,N_6619);
nand U11339 (N_11339,N_8225,N_8786);
and U11340 (N_11340,N_7461,N_6710);
nand U11341 (N_11341,N_9334,N_7173);
or U11342 (N_11342,N_8039,N_8250);
and U11343 (N_11343,N_7707,N_8576);
xor U11344 (N_11344,N_6893,N_7835);
nand U11345 (N_11345,N_7357,N_7001);
or U11346 (N_11346,N_8217,N_9183);
or U11347 (N_11347,N_6958,N_7619);
or U11348 (N_11348,N_7000,N_7550);
or U11349 (N_11349,N_8529,N_6860);
xnor U11350 (N_11350,N_9053,N_8914);
or U11351 (N_11351,N_8535,N_7579);
nand U11352 (N_11352,N_7062,N_6578);
and U11353 (N_11353,N_7001,N_6297);
nor U11354 (N_11354,N_8677,N_7440);
nor U11355 (N_11355,N_8416,N_7592);
or U11356 (N_11356,N_8290,N_8743);
or U11357 (N_11357,N_8374,N_8541);
and U11358 (N_11358,N_8951,N_6547);
nand U11359 (N_11359,N_6364,N_8137);
or U11360 (N_11360,N_8309,N_8663);
and U11361 (N_11361,N_8898,N_6388);
xnor U11362 (N_11362,N_9232,N_8911);
and U11363 (N_11363,N_7655,N_8530);
or U11364 (N_11364,N_8640,N_7994);
xor U11365 (N_11365,N_8052,N_6592);
and U11366 (N_11366,N_8451,N_8477);
and U11367 (N_11367,N_9112,N_8972);
and U11368 (N_11368,N_7153,N_7268);
nor U11369 (N_11369,N_6268,N_8541);
nor U11370 (N_11370,N_7640,N_6586);
xnor U11371 (N_11371,N_7064,N_6379);
nand U11372 (N_11372,N_6263,N_9269);
and U11373 (N_11373,N_9368,N_6849);
nand U11374 (N_11374,N_6972,N_7932);
and U11375 (N_11375,N_7962,N_6719);
nor U11376 (N_11376,N_6741,N_8349);
and U11377 (N_11377,N_7072,N_7645);
and U11378 (N_11378,N_6896,N_8992);
and U11379 (N_11379,N_7705,N_6370);
nand U11380 (N_11380,N_7655,N_8790);
and U11381 (N_11381,N_6923,N_7212);
nand U11382 (N_11382,N_7523,N_8587);
nand U11383 (N_11383,N_8299,N_8785);
nand U11384 (N_11384,N_8507,N_8102);
xor U11385 (N_11385,N_8651,N_9258);
or U11386 (N_11386,N_8785,N_6527);
nand U11387 (N_11387,N_6286,N_7977);
and U11388 (N_11388,N_8414,N_9289);
nand U11389 (N_11389,N_9211,N_7215);
or U11390 (N_11390,N_6765,N_6534);
nand U11391 (N_11391,N_7576,N_6262);
and U11392 (N_11392,N_8804,N_8096);
nand U11393 (N_11393,N_8683,N_8419);
nand U11394 (N_11394,N_8512,N_8208);
nand U11395 (N_11395,N_7899,N_7503);
nand U11396 (N_11396,N_8985,N_7146);
xor U11397 (N_11397,N_7165,N_7428);
and U11398 (N_11398,N_6499,N_9215);
nand U11399 (N_11399,N_9163,N_6302);
or U11400 (N_11400,N_7586,N_7241);
nor U11401 (N_11401,N_7502,N_7391);
nand U11402 (N_11402,N_8793,N_8925);
or U11403 (N_11403,N_7370,N_8519);
and U11404 (N_11404,N_6258,N_6708);
nand U11405 (N_11405,N_6744,N_8681);
or U11406 (N_11406,N_8543,N_7036);
nand U11407 (N_11407,N_7911,N_7197);
nand U11408 (N_11408,N_6493,N_7192);
and U11409 (N_11409,N_7575,N_7599);
nor U11410 (N_11410,N_8170,N_9245);
and U11411 (N_11411,N_8866,N_7617);
nand U11412 (N_11412,N_7994,N_8163);
or U11413 (N_11413,N_8011,N_9001);
and U11414 (N_11414,N_9180,N_7349);
or U11415 (N_11415,N_8727,N_7323);
or U11416 (N_11416,N_8905,N_7526);
nor U11417 (N_11417,N_8859,N_7379);
or U11418 (N_11418,N_6490,N_7320);
xor U11419 (N_11419,N_8206,N_8708);
nand U11420 (N_11420,N_9105,N_8635);
and U11421 (N_11421,N_9182,N_7588);
and U11422 (N_11422,N_6987,N_7173);
nand U11423 (N_11423,N_9206,N_8195);
xnor U11424 (N_11424,N_9199,N_8278);
and U11425 (N_11425,N_7526,N_7428);
nor U11426 (N_11426,N_7895,N_6690);
and U11427 (N_11427,N_8140,N_9363);
nor U11428 (N_11428,N_9236,N_7498);
xnor U11429 (N_11429,N_9199,N_8186);
and U11430 (N_11430,N_7526,N_8122);
xor U11431 (N_11431,N_8831,N_7131);
nor U11432 (N_11432,N_7936,N_7123);
nor U11433 (N_11433,N_7563,N_8596);
and U11434 (N_11434,N_8817,N_8808);
nor U11435 (N_11435,N_8219,N_7414);
or U11436 (N_11436,N_7462,N_8927);
and U11437 (N_11437,N_7304,N_6620);
xnor U11438 (N_11438,N_8747,N_7062);
nor U11439 (N_11439,N_8837,N_6749);
nor U11440 (N_11440,N_6600,N_7306);
nand U11441 (N_11441,N_7386,N_9027);
xor U11442 (N_11442,N_7471,N_8985);
nor U11443 (N_11443,N_6688,N_9281);
xor U11444 (N_11444,N_8342,N_7494);
nor U11445 (N_11445,N_8788,N_9247);
nand U11446 (N_11446,N_8768,N_8354);
and U11447 (N_11447,N_8106,N_8358);
xnor U11448 (N_11448,N_7930,N_8675);
and U11449 (N_11449,N_6556,N_8648);
nor U11450 (N_11450,N_6568,N_6267);
and U11451 (N_11451,N_8184,N_9217);
nor U11452 (N_11452,N_7739,N_7459);
and U11453 (N_11453,N_7208,N_6441);
xnor U11454 (N_11454,N_8378,N_8550);
nand U11455 (N_11455,N_8324,N_7027);
or U11456 (N_11456,N_6380,N_8871);
and U11457 (N_11457,N_9267,N_7206);
and U11458 (N_11458,N_7060,N_7088);
and U11459 (N_11459,N_7211,N_7734);
nor U11460 (N_11460,N_6474,N_8413);
nor U11461 (N_11461,N_7953,N_8932);
and U11462 (N_11462,N_7044,N_9367);
and U11463 (N_11463,N_6670,N_9031);
or U11464 (N_11464,N_7774,N_9152);
nand U11465 (N_11465,N_9220,N_9162);
and U11466 (N_11466,N_7791,N_7970);
and U11467 (N_11467,N_7558,N_7036);
or U11468 (N_11468,N_8557,N_9002);
nor U11469 (N_11469,N_6712,N_6296);
and U11470 (N_11470,N_6658,N_9134);
or U11471 (N_11471,N_7748,N_7170);
nor U11472 (N_11472,N_6986,N_6769);
and U11473 (N_11473,N_7701,N_8226);
nor U11474 (N_11474,N_8391,N_7364);
nor U11475 (N_11475,N_9262,N_8424);
or U11476 (N_11476,N_8359,N_8737);
nand U11477 (N_11477,N_7394,N_6414);
nand U11478 (N_11478,N_8689,N_7303);
nor U11479 (N_11479,N_7832,N_6815);
nor U11480 (N_11480,N_6622,N_7569);
nand U11481 (N_11481,N_6792,N_7982);
and U11482 (N_11482,N_7565,N_7607);
nand U11483 (N_11483,N_6706,N_6958);
and U11484 (N_11484,N_7510,N_7410);
xnor U11485 (N_11485,N_7473,N_7603);
or U11486 (N_11486,N_8252,N_6596);
and U11487 (N_11487,N_7631,N_8469);
and U11488 (N_11488,N_6329,N_8691);
and U11489 (N_11489,N_8874,N_7052);
or U11490 (N_11490,N_6685,N_8110);
nor U11491 (N_11491,N_8110,N_7485);
or U11492 (N_11492,N_7878,N_7994);
nand U11493 (N_11493,N_6809,N_8434);
nand U11494 (N_11494,N_9192,N_6987);
nand U11495 (N_11495,N_7330,N_6950);
nor U11496 (N_11496,N_8974,N_7410);
nor U11497 (N_11497,N_8194,N_9127);
and U11498 (N_11498,N_6929,N_8803);
xor U11499 (N_11499,N_8430,N_6929);
or U11500 (N_11500,N_7428,N_7371);
xnor U11501 (N_11501,N_9306,N_8978);
nor U11502 (N_11502,N_8363,N_8205);
nor U11503 (N_11503,N_6864,N_7301);
nor U11504 (N_11504,N_8590,N_8940);
and U11505 (N_11505,N_6488,N_9312);
or U11506 (N_11506,N_7333,N_8873);
or U11507 (N_11507,N_6681,N_7212);
nor U11508 (N_11508,N_7481,N_7800);
nand U11509 (N_11509,N_6272,N_7842);
nor U11510 (N_11510,N_8205,N_7708);
xor U11511 (N_11511,N_7349,N_7908);
and U11512 (N_11512,N_8070,N_8753);
xor U11513 (N_11513,N_8730,N_6472);
nand U11514 (N_11514,N_8295,N_8736);
xnor U11515 (N_11515,N_7588,N_8343);
nor U11516 (N_11516,N_6547,N_7692);
and U11517 (N_11517,N_7504,N_8542);
and U11518 (N_11518,N_9025,N_7012);
or U11519 (N_11519,N_7607,N_7032);
and U11520 (N_11520,N_9273,N_6866);
xnor U11521 (N_11521,N_9316,N_7911);
or U11522 (N_11522,N_8126,N_9282);
xor U11523 (N_11523,N_8613,N_9359);
nand U11524 (N_11524,N_8392,N_9118);
and U11525 (N_11525,N_6879,N_7037);
xor U11526 (N_11526,N_6258,N_7074);
nand U11527 (N_11527,N_7276,N_7846);
and U11528 (N_11528,N_7939,N_6440);
and U11529 (N_11529,N_7479,N_7242);
nand U11530 (N_11530,N_7525,N_6492);
and U11531 (N_11531,N_8681,N_9240);
or U11532 (N_11532,N_9106,N_6299);
and U11533 (N_11533,N_8212,N_8562);
nand U11534 (N_11534,N_8381,N_9280);
and U11535 (N_11535,N_8677,N_6431);
nand U11536 (N_11536,N_6356,N_6440);
nand U11537 (N_11537,N_6669,N_7686);
and U11538 (N_11538,N_8817,N_7587);
nand U11539 (N_11539,N_7299,N_6547);
and U11540 (N_11540,N_8911,N_6568);
nand U11541 (N_11541,N_6454,N_8177);
nor U11542 (N_11542,N_7319,N_8455);
or U11543 (N_11543,N_9262,N_6660);
and U11544 (N_11544,N_7652,N_6577);
or U11545 (N_11545,N_8542,N_8418);
nor U11546 (N_11546,N_8545,N_6651);
and U11547 (N_11547,N_8188,N_7932);
xnor U11548 (N_11548,N_6907,N_6558);
and U11549 (N_11549,N_7298,N_8624);
or U11550 (N_11550,N_6981,N_8837);
and U11551 (N_11551,N_7480,N_9076);
nor U11552 (N_11552,N_8143,N_9048);
nand U11553 (N_11553,N_6548,N_6323);
nand U11554 (N_11554,N_6313,N_7135);
nand U11555 (N_11555,N_8800,N_8220);
or U11556 (N_11556,N_7342,N_6736);
or U11557 (N_11557,N_6268,N_6355);
and U11558 (N_11558,N_8172,N_8688);
nor U11559 (N_11559,N_8497,N_8985);
nand U11560 (N_11560,N_7743,N_6263);
or U11561 (N_11561,N_7200,N_7893);
nor U11562 (N_11562,N_8461,N_7124);
and U11563 (N_11563,N_6252,N_7026);
nand U11564 (N_11564,N_7731,N_8485);
or U11565 (N_11565,N_6380,N_7657);
nand U11566 (N_11566,N_6295,N_9093);
xor U11567 (N_11567,N_8051,N_8033);
nand U11568 (N_11568,N_7206,N_7831);
xor U11569 (N_11569,N_6273,N_8576);
nand U11570 (N_11570,N_8350,N_9231);
nor U11571 (N_11571,N_6710,N_7619);
or U11572 (N_11572,N_7048,N_7020);
nor U11573 (N_11573,N_7271,N_7463);
or U11574 (N_11574,N_9206,N_8156);
or U11575 (N_11575,N_8667,N_7738);
nand U11576 (N_11576,N_8632,N_6943);
nor U11577 (N_11577,N_6465,N_7871);
nand U11578 (N_11578,N_7927,N_8479);
nor U11579 (N_11579,N_9085,N_8451);
or U11580 (N_11580,N_7137,N_7850);
or U11581 (N_11581,N_8730,N_8275);
or U11582 (N_11582,N_9148,N_8146);
and U11583 (N_11583,N_7317,N_7498);
nor U11584 (N_11584,N_9062,N_6351);
and U11585 (N_11585,N_7258,N_7659);
nor U11586 (N_11586,N_7157,N_6461);
or U11587 (N_11587,N_6761,N_7017);
nor U11588 (N_11588,N_9334,N_7630);
and U11589 (N_11589,N_6545,N_7396);
and U11590 (N_11590,N_9256,N_8658);
or U11591 (N_11591,N_6280,N_7479);
and U11592 (N_11592,N_9068,N_7362);
or U11593 (N_11593,N_8386,N_8489);
nor U11594 (N_11594,N_7526,N_6342);
nor U11595 (N_11595,N_7366,N_7750);
and U11596 (N_11596,N_8759,N_7545);
and U11597 (N_11597,N_7956,N_8704);
or U11598 (N_11598,N_8231,N_7849);
or U11599 (N_11599,N_9251,N_9020);
or U11600 (N_11600,N_7651,N_6836);
or U11601 (N_11601,N_8669,N_6542);
or U11602 (N_11602,N_8020,N_6641);
nand U11603 (N_11603,N_8695,N_8542);
nand U11604 (N_11604,N_7952,N_6469);
and U11605 (N_11605,N_6990,N_7304);
and U11606 (N_11606,N_8955,N_7133);
nor U11607 (N_11607,N_6911,N_8134);
and U11608 (N_11608,N_6352,N_7277);
nor U11609 (N_11609,N_6337,N_8757);
nand U11610 (N_11610,N_7722,N_8031);
and U11611 (N_11611,N_6650,N_6516);
or U11612 (N_11612,N_8026,N_6793);
or U11613 (N_11613,N_7677,N_7961);
or U11614 (N_11614,N_7995,N_8515);
nor U11615 (N_11615,N_7503,N_8087);
nor U11616 (N_11616,N_6300,N_9007);
xor U11617 (N_11617,N_8148,N_8211);
nor U11618 (N_11618,N_6627,N_8817);
nor U11619 (N_11619,N_7432,N_6401);
nand U11620 (N_11620,N_8672,N_8106);
or U11621 (N_11621,N_8738,N_9290);
or U11622 (N_11622,N_8053,N_9002);
or U11623 (N_11623,N_9336,N_8222);
nor U11624 (N_11624,N_6659,N_8462);
nand U11625 (N_11625,N_7175,N_8855);
nand U11626 (N_11626,N_9064,N_6335);
nand U11627 (N_11627,N_8556,N_8619);
nand U11628 (N_11628,N_7662,N_8296);
nor U11629 (N_11629,N_9344,N_8844);
and U11630 (N_11630,N_6308,N_6315);
xor U11631 (N_11631,N_9350,N_7506);
or U11632 (N_11632,N_6724,N_8116);
and U11633 (N_11633,N_8611,N_7835);
and U11634 (N_11634,N_8196,N_9099);
nand U11635 (N_11635,N_8792,N_8582);
nor U11636 (N_11636,N_7852,N_8161);
or U11637 (N_11637,N_7383,N_9307);
nand U11638 (N_11638,N_7539,N_8839);
and U11639 (N_11639,N_8407,N_9194);
or U11640 (N_11640,N_7688,N_7954);
or U11641 (N_11641,N_8373,N_6688);
or U11642 (N_11642,N_8276,N_6254);
and U11643 (N_11643,N_8445,N_8120);
nor U11644 (N_11644,N_8570,N_8014);
or U11645 (N_11645,N_6886,N_9046);
nand U11646 (N_11646,N_8655,N_7969);
nor U11647 (N_11647,N_7106,N_6563);
and U11648 (N_11648,N_8260,N_7077);
or U11649 (N_11649,N_8004,N_7255);
or U11650 (N_11650,N_9091,N_7398);
nor U11651 (N_11651,N_8356,N_8406);
xnor U11652 (N_11652,N_8003,N_8817);
xnor U11653 (N_11653,N_8501,N_7464);
nor U11654 (N_11654,N_8051,N_7921);
and U11655 (N_11655,N_6350,N_8939);
or U11656 (N_11656,N_6818,N_9114);
nor U11657 (N_11657,N_7880,N_7638);
nand U11658 (N_11658,N_9361,N_6466);
xnor U11659 (N_11659,N_9321,N_9175);
nor U11660 (N_11660,N_9023,N_8338);
nor U11661 (N_11661,N_7395,N_6754);
or U11662 (N_11662,N_6338,N_6574);
nor U11663 (N_11663,N_6813,N_8066);
nor U11664 (N_11664,N_7317,N_6487);
xnor U11665 (N_11665,N_6806,N_7519);
xor U11666 (N_11666,N_8389,N_8088);
nor U11667 (N_11667,N_7858,N_9181);
and U11668 (N_11668,N_7363,N_7214);
nor U11669 (N_11669,N_6755,N_8824);
or U11670 (N_11670,N_8280,N_7101);
nand U11671 (N_11671,N_7498,N_6804);
and U11672 (N_11672,N_6788,N_7807);
or U11673 (N_11673,N_9064,N_6633);
and U11674 (N_11674,N_6281,N_7056);
and U11675 (N_11675,N_8477,N_6332);
nand U11676 (N_11676,N_7061,N_8616);
nor U11677 (N_11677,N_7428,N_9043);
nand U11678 (N_11678,N_7358,N_9343);
or U11679 (N_11679,N_7452,N_7677);
nor U11680 (N_11680,N_6568,N_7417);
nand U11681 (N_11681,N_8076,N_8137);
or U11682 (N_11682,N_8695,N_7031);
nand U11683 (N_11683,N_7804,N_6605);
nand U11684 (N_11684,N_7934,N_8363);
nor U11685 (N_11685,N_6359,N_6704);
nand U11686 (N_11686,N_6452,N_8874);
or U11687 (N_11687,N_8338,N_7633);
and U11688 (N_11688,N_9371,N_6466);
and U11689 (N_11689,N_9114,N_6661);
or U11690 (N_11690,N_6579,N_7927);
nor U11691 (N_11691,N_6407,N_9006);
or U11692 (N_11692,N_6451,N_7440);
nand U11693 (N_11693,N_9121,N_8535);
xnor U11694 (N_11694,N_6909,N_7966);
xor U11695 (N_11695,N_7245,N_8796);
nor U11696 (N_11696,N_8048,N_6536);
nor U11697 (N_11697,N_7785,N_7769);
nand U11698 (N_11698,N_8912,N_9148);
nand U11699 (N_11699,N_7816,N_7450);
nor U11700 (N_11700,N_7873,N_6634);
xor U11701 (N_11701,N_6417,N_8634);
and U11702 (N_11702,N_8865,N_8986);
and U11703 (N_11703,N_9310,N_8908);
nor U11704 (N_11704,N_7979,N_7023);
nor U11705 (N_11705,N_6847,N_6487);
nor U11706 (N_11706,N_8266,N_7745);
nor U11707 (N_11707,N_8021,N_7462);
nand U11708 (N_11708,N_7591,N_8567);
and U11709 (N_11709,N_7135,N_8462);
nand U11710 (N_11710,N_8567,N_6695);
nor U11711 (N_11711,N_7315,N_8425);
or U11712 (N_11712,N_7168,N_6254);
or U11713 (N_11713,N_8417,N_7702);
xnor U11714 (N_11714,N_8416,N_9217);
xor U11715 (N_11715,N_8129,N_6894);
and U11716 (N_11716,N_7072,N_6876);
or U11717 (N_11717,N_7624,N_6913);
or U11718 (N_11718,N_6791,N_8799);
nor U11719 (N_11719,N_6288,N_7099);
nand U11720 (N_11720,N_6473,N_8720);
nor U11721 (N_11721,N_6547,N_7320);
nand U11722 (N_11722,N_9198,N_6575);
nor U11723 (N_11723,N_7514,N_8503);
and U11724 (N_11724,N_8948,N_6365);
nor U11725 (N_11725,N_7572,N_9141);
nand U11726 (N_11726,N_8300,N_9088);
or U11727 (N_11727,N_8835,N_8609);
nor U11728 (N_11728,N_8631,N_7629);
or U11729 (N_11729,N_8388,N_6990);
nor U11730 (N_11730,N_8314,N_8857);
nor U11731 (N_11731,N_9004,N_6930);
xor U11732 (N_11732,N_8571,N_8944);
nand U11733 (N_11733,N_6456,N_9174);
and U11734 (N_11734,N_6616,N_6344);
nor U11735 (N_11735,N_8846,N_7236);
or U11736 (N_11736,N_8829,N_7071);
nor U11737 (N_11737,N_7967,N_8530);
or U11738 (N_11738,N_8031,N_7893);
or U11739 (N_11739,N_6760,N_7310);
nand U11740 (N_11740,N_6955,N_8396);
nor U11741 (N_11741,N_7939,N_7659);
nor U11742 (N_11742,N_7698,N_8281);
or U11743 (N_11743,N_7333,N_8405);
nor U11744 (N_11744,N_8107,N_7834);
nor U11745 (N_11745,N_7177,N_9007);
and U11746 (N_11746,N_7702,N_8682);
or U11747 (N_11747,N_8709,N_9023);
nor U11748 (N_11748,N_8166,N_6869);
and U11749 (N_11749,N_9344,N_7781);
and U11750 (N_11750,N_6536,N_7734);
or U11751 (N_11751,N_8264,N_8411);
or U11752 (N_11752,N_8314,N_8024);
or U11753 (N_11753,N_7058,N_9265);
nand U11754 (N_11754,N_7503,N_6515);
and U11755 (N_11755,N_9294,N_6988);
or U11756 (N_11756,N_9358,N_8992);
xor U11757 (N_11757,N_9139,N_7431);
or U11758 (N_11758,N_6826,N_7456);
nand U11759 (N_11759,N_8448,N_8342);
nor U11760 (N_11760,N_8913,N_7091);
nand U11761 (N_11761,N_9021,N_7949);
and U11762 (N_11762,N_7259,N_8424);
nor U11763 (N_11763,N_6339,N_6669);
nand U11764 (N_11764,N_7414,N_7137);
or U11765 (N_11765,N_7792,N_6677);
and U11766 (N_11766,N_7339,N_9153);
or U11767 (N_11767,N_7003,N_7553);
nor U11768 (N_11768,N_7843,N_7789);
or U11769 (N_11769,N_8020,N_6571);
nand U11770 (N_11770,N_7569,N_6383);
or U11771 (N_11771,N_6386,N_8276);
nand U11772 (N_11772,N_6257,N_7649);
or U11773 (N_11773,N_7885,N_8220);
or U11774 (N_11774,N_9185,N_7894);
and U11775 (N_11775,N_9253,N_7143);
nor U11776 (N_11776,N_7757,N_7042);
or U11777 (N_11777,N_6941,N_7787);
nor U11778 (N_11778,N_8966,N_8757);
and U11779 (N_11779,N_7050,N_7676);
xor U11780 (N_11780,N_8077,N_7806);
nand U11781 (N_11781,N_8548,N_6842);
and U11782 (N_11782,N_7177,N_9074);
or U11783 (N_11783,N_8949,N_7103);
nand U11784 (N_11784,N_8197,N_6687);
or U11785 (N_11785,N_8649,N_7133);
or U11786 (N_11786,N_8016,N_7310);
and U11787 (N_11787,N_7606,N_6423);
nand U11788 (N_11788,N_8726,N_8943);
and U11789 (N_11789,N_6373,N_8824);
or U11790 (N_11790,N_7913,N_8034);
nand U11791 (N_11791,N_9186,N_7350);
and U11792 (N_11792,N_6356,N_6349);
nand U11793 (N_11793,N_8663,N_6272);
nand U11794 (N_11794,N_7421,N_7096);
xnor U11795 (N_11795,N_8590,N_7375);
and U11796 (N_11796,N_6419,N_7936);
and U11797 (N_11797,N_6312,N_8516);
nand U11798 (N_11798,N_7411,N_9199);
nand U11799 (N_11799,N_7434,N_9238);
nor U11800 (N_11800,N_7234,N_9255);
nand U11801 (N_11801,N_7266,N_9138);
and U11802 (N_11802,N_7542,N_6615);
or U11803 (N_11803,N_8079,N_7638);
nor U11804 (N_11804,N_6400,N_8361);
and U11805 (N_11805,N_6283,N_8392);
and U11806 (N_11806,N_7413,N_7708);
nor U11807 (N_11807,N_6572,N_8639);
and U11808 (N_11808,N_6661,N_6721);
nand U11809 (N_11809,N_7049,N_7782);
nand U11810 (N_11810,N_8913,N_8715);
nor U11811 (N_11811,N_8363,N_7617);
nor U11812 (N_11812,N_6426,N_6982);
nand U11813 (N_11813,N_6999,N_6954);
or U11814 (N_11814,N_6971,N_6667);
xnor U11815 (N_11815,N_9170,N_8801);
nor U11816 (N_11816,N_9233,N_7725);
xnor U11817 (N_11817,N_7651,N_7639);
nand U11818 (N_11818,N_6606,N_6860);
nor U11819 (N_11819,N_7708,N_9187);
and U11820 (N_11820,N_6884,N_6820);
or U11821 (N_11821,N_7508,N_9219);
nand U11822 (N_11822,N_8436,N_6973);
nand U11823 (N_11823,N_8098,N_8337);
nand U11824 (N_11824,N_6566,N_9156);
or U11825 (N_11825,N_6281,N_8608);
nand U11826 (N_11826,N_7236,N_6321);
and U11827 (N_11827,N_7374,N_6637);
nor U11828 (N_11828,N_6794,N_7835);
nor U11829 (N_11829,N_8121,N_6481);
or U11830 (N_11830,N_7402,N_7851);
or U11831 (N_11831,N_9040,N_6521);
or U11832 (N_11832,N_6302,N_8879);
or U11833 (N_11833,N_7147,N_9204);
or U11834 (N_11834,N_8579,N_8155);
and U11835 (N_11835,N_8332,N_8496);
nor U11836 (N_11836,N_9261,N_9023);
xnor U11837 (N_11837,N_7144,N_6616);
nand U11838 (N_11838,N_6973,N_8621);
or U11839 (N_11839,N_7925,N_7433);
or U11840 (N_11840,N_8167,N_9188);
nor U11841 (N_11841,N_7043,N_8504);
xor U11842 (N_11842,N_7263,N_8546);
nor U11843 (N_11843,N_8547,N_8182);
and U11844 (N_11844,N_9034,N_8716);
xnor U11845 (N_11845,N_7819,N_6959);
and U11846 (N_11846,N_7452,N_6858);
and U11847 (N_11847,N_8352,N_7494);
nand U11848 (N_11848,N_7294,N_7795);
nor U11849 (N_11849,N_8065,N_7970);
and U11850 (N_11850,N_9078,N_6955);
and U11851 (N_11851,N_8421,N_6462);
nand U11852 (N_11852,N_6781,N_7136);
nand U11853 (N_11853,N_8874,N_8485);
or U11854 (N_11854,N_8819,N_6268);
or U11855 (N_11855,N_6970,N_9089);
or U11856 (N_11856,N_6337,N_8433);
xor U11857 (N_11857,N_7424,N_8026);
or U11858 (N_11858,N_6789,N_8459);
nand U11859 (N_11859,N_8934,N_7961);
xor U11860 (N_11860,N_6420,N_7261);
nor U11861 (N_11861,N_7774,N_7187);
xor U11862 (N_11862,N_7569,N_7130);
nand U11863 (N_11863,N_8319,N_8361);
xnor U11864 (N_11864,N_7742,N_8067);
nand U11865 (N_11865,N_9165,N_7390);
or U11866 (N_11866,N_6792,N_7321);
xor U11867 (N_11867,N_9223,N_7638);
or U11868 (N_11868,N_8697,N_7294);
nor U11869 (N_11869,N_8818,N_6257);
nand U11870 (N_11870,N_6387,N_6741);
or U11871 (N_11871,N_8130,N_8289);
or U11872 (N_11872,N_7447,N_6813);
and U11873 (N_11873,N_9185,N_6408);
nand U11874 (N_11874,N_7557,N_6298);
or U11875 (N_11875,N_6372,N_8995);
nor U11876 (N_11876,N_6899,N_6971);
or U11877 (N_11877,N_7864,N_8911);
nand U11878 (N_11878,N_8534,N_8207);
nor U11879 (N_11879,N_6608,N_7849);
nand U11880 (N_11880,N_9128,N_8326);
nand U11881 (N_11881,N_6735,N_7194);
and U11882 (N_11882,N_9295,N_8171);
nand U11883 (N_11883,N_8993,N_8063);
or U11884 (N_11884,N_7079,N_7798);
nand U11885 (N_11885,N_6454,N_8436);
and U11886 (N_11886,N_7006,N_6361);
nor U11887 (N_11887,N_6255,N_8938);
nand U11888 (N_11888,N_6527,N_8825);
nor U11889 (N_11889,N_8593,N_7503);
and U11890 (N_11890,N_8208,N_7668);
or U11891 (N_11891,N_8659,N_9100);
and U11892 (N_11892,N_8597,N_7582);
nor U11893 (N_11893,N_6496,N_9370);
and U11894 (N_11894,N_8411,N_8248);
nor U11895 (N_11895,N_8131,N_9244);
and U11896 (N_11896,N_9020,N_8844);
nand U11897 (N_11897,N_7128,N_7344);
or U11898 (N_11898,N_6435,N_7135);
and U11899 (N_11899,N_6447,N_8363);
nand U11900 (N_11900,N_8668,N_9066);
nand U11901 (N_11901,N_7406,N_8164);
xor U11902 (N_11902,N_7304,N_8728);
and U11903 (N_11903,N_7573,N_8750);
and U11904 (N_11904,N_8606,N_8589);
nand U11905 (N_11905,N_6299,N_6880);
xor U11906 (N_11906,N_7778,N_9364);
and U11907 (N_11907,N_7643,N_7503);
nor U11908 (N_11908,N_9339,N_9015);
and U11909 (N_11909,N_8997,N_6438);
nand U11910 (N_11910,N_7565,N_7025);
or U11911 (N_11911,N_9240,N_8069);
nor U11912 (N_11912,N_9247,N_7798);
and U11913 (N_11913,N_6626,N_6996);
nand U11914 (N_11914,N_7531,N_7068);
nand U11915 (N_11915,N_6959,N_6419);
xor U11916 (N_11916,N_8177,N_6509);
xnor U11917 (N_11917,N_7137,N_7829);
and U11918 (N_11918,N_7866,N_9201);
nand U11919 (N_11919,N_8276,N_9037);
nor U11920 (N_11920,N_7470,N_8439);
or U11921 (N_11921,N_9201,N_8992);
and U11922 (N_11922,N_6769,N_8754);
nand U11923 (N_11923,N_8789,N_6663);
or U11924 (N_11924,N_8163,N_8982);
and U11925 (N_11925,N_8285,N_8341);
or U11926 (N_11926,N_8584,N_6680);
nor U11927 (N_11927,N_6851,N_6918);
nor U11928 (N_11928,N_6915,N_6781);
or U11929 (N_11929,N_8681,N_7681);
or U11930 (N_11930,N_7388,N_9053);
xnor U11931 (N_11931,N_7270,N_7132);
or U11932 (N_11932,N_8686,N_6719);
nor U11933 (N_11933,N_9209,N_6668);
and U11934 (N_11934,N_8946,N_7003);
nand U11935 (N_11935,N_6915,N_6260);
nand U11936 (N_11936,N_7864,N_6440);
nor U11937 (N_11937,N_6675,N_7228);
nand U11938 (N_11938,N_8929,N_6414);
and U11939 (N_11939,N_7925,N_6469);
xor U11940 (N_11940,N_6477,N_8287);
and U11941 (N_11941,N_6448,N_6308);
and U11942 (N_11942,N_8204,N_6956);
xnor U11943 (N_11943,N_6309,N_7978);
or U11944 (N_11944,N_8667,N_8118);
nand U11945 (N_11945,N_7278,N_8109);
xnor U11946 (N_11946,N_7282,N_7316);
nand U11947 (N_11947,N_7776,N_8860);
nand U11948 (N_11948,N_7749,N_6812);
xnor U11949 (N_11949,N_8555,N_8129);
xor U11950 (N_11950,N_8678,N_7899);
or U11951 (N_11951,N_8123,N_8725);
and U11952 (N_11952,N_7180,N_9239);
nand U11953 (N_11953,N_8961,N_7758);
nor U11954 (N_11954,N_6593,N_7105);
and U11955 (N_11955,N_8618,N_9201);
or U11956 (N_11956,N_7699,N_9080);
nor U11957 (N_11957,N_7255,N_8160);
or U11958 (N_11958,N_7842,N_8128);
xnor U11959 (N_11959,N_6389,N_6584);
xor U11960 (N_11960,N_8265,N_8856);
and U11961 (N_11961,N_7140,N_7803);
and U11962 (N_11962,N_9130,N_8687);
and U11963 (N_11963,N_6763,N_8546);
or U11964 (N_11964,N_9113,N_6786);
and U11965 (N_11965,N_8333,N_6812);
or U11966 (N_11966,N_9004,N_6860);
nor U11967 (N_11967,N_7451,N_8050);
or U11968 (N_11968,N_8666,N_8852);
and U11969 (N_11969,N_6359,N_7247);
or U11970 (N_11970,N_8373,N_9119);
or U11971 (N_11971,N_9296,N_8236);
and U11972 (N_11972,N_7676,N_6812);
or U11973 (N_11973,N_8180,N_7930);
and U11974 (N_11974,N_7225,N_6641);
nor U11975 (N_11975,N_6891,N_7446);
nand U11976 (N_11976,N_8920,N_7835);
nor U11977 (N_11977,N_8744,N_7452);
and U11978 (N_11978,N_6774,N_7896);
nand U11979 (N_11979,N_9029,N_6610);
xor U11980 (N_11980,N_7983,N_7538);
nor U11981 (N_11981,N_8150,N_8207);
xor U11982 (N_11982,N_6783,N_6584);
and U11983 (N_11983,N_6875,N_6611);
xor U11984 (N_11984,N_8793,N_6376);
or U11985 (N_11985,N_8759,N_7664);
nand U11986 (N_11986,N_6563,N_6617);
or U11987 (N_11987,N_6846,N_8599);
and U11988 (N_11988,N_7040,N_8220);
nor U11989 (N_11989,N_7292,N_6601);
xor U11990 (N_11990,N_7489,N_7695);
nand U11991 (N_11991,N_8233,N_7910);
and U11992 (N_11992,N_7834,N_6410);
nor U11993 (N_11993,N_7106,N_9236);
xor U11994 (N_11994,N_6796,N_6969);
nor U11995 (N_11995,N_6851,N_8361);
nand U11996 (N_11996,N_8795,N_7526);
or U11997 (N_11997,N_8552,N_7691);
and U11998 (N_11998,N_6459,N_8924);
or U11999 (N_11999,N_6926,N_7132);
nand U12000 (N_12000,N_8580,N_8292);
or U12001 (N_12001,N_7721,N_6351);
nor U12002 (N_12002,N_8628,N_7469);
nand U12003 (N_12003,N_6636,N_6594);
nand U12004 (N_12004,N_6466,N_9291);
or U12005 (N_12005,N_9040,N_8939);
nor U12006 (N_12006,N_7588,N_8972);
or U12007 (N_12007,N_7394,N_6439);
or U12008 (N_12008,N_9041,N_7329);
or U12009 (N_12009,N_7940,N_8426);
and U12010 (N_12010,N_8316,N_9344);
nand U12011 (N_12011,N_8913,N_8903);
or U12012 (N_12012,N_7965,N_6321);
and U12013 (N_12013,N_6475,N_8753);
nand U12014 (N_12014,N_7688,N_9253);
nor U12015 (N_12015,N_7431,N_6387);
xor U12016 (N_12016,N_6472,N_8845);
nor U12017 (N_12017,N_7183,N_6390);
and U12018 (N_12018,N_8371,N_6696);
and U12019 (N_12019,N_8007,N_9257);
nor U12020 (N_12020,N_8924,N_8321);
and U12021 (N_12021,N_8223,N_8262);
nor U12022 (N_12022,N_8385,N_8041);
xnor U12023 (N_12023,N_8002,N_6556);
or U12024 (N_12024,N_8145,N_7273);
nor U12025 (N_12025,N_8843,N_6334);
and U12026 (N_12026,N_7499,N_8530);
and U12027 (N_12027,N_8224,N_7540);
or U12028 (N_12028,N_8883,N_8680);
or U12029 (N_12029,N_8522,N_7259);
or U12030 (N_12030,N_6838,N_9135);
nor U12031 (N_12031,N_8943,N_7525);
and U12032 (N_12032,N_8631,N_9337);
nand U12033 (N_12033,N_7589,N_6845);
nor U12034 (N_12034,N_7278,N_9264);
xor U12035 (N_12035,N_9201,N_9284);
nor U12036 (N_12036,N_6414,N_8033);
and U12037 (N_12037,N_6465,N_7333);
and U12038 (N_12038,N_7527,N_8873);
xnor U12039 (N_12039,N_8679,N_9286);
or U12040 (N_12040,N_8672,N_8270);
and U12041 (N_12041,N_8466,N_7541);
or U12042 (N_12042,N_7763,N_8821);
and U12043 (N_12043,N_7622,N_6489);
xor U12044 (N_12044,N_8706,N_8772);
or U12045 (N_12045,N_7358,N_6472);
and U12046 (N_12046,N_6296,N_6510);
or U12047 (N_12047,N_6644,N_8117);
nor U12048 (N_12048,N_6894,N_8519);
and U12049 (N_12049,N_6938,N_8061);
or U12050 (N_12050,N_9240,N_7571);
and U12051 (N_12051,N_7905,N_7422);
nor U12052 (N_12052,N_6365,N_7438);
and U12053 (N_12053,N_7243,N_7360);
nor U12054 (N_12054,N_7897,N_6485);
or U12055 (N_12055,N_9166,N_6681);
xnor U12056 (N_12056,N_6287,N_6426);
and U12057 (N_12057,N_7526,N_7770);
or U12058 (N_12058,N_7756,N_7619);
nand U12059 (N_12059,N_7581,N_7615);
and U12060 (N_12060,N_9206,N_8180);
and U12061 (N_12061,N_8286,N_7638);
nand U12062 (N_12062,N_6887,N_7153);
or U12063 (N_12063,N_8583,N_6656);
and U12064 (N_12064,N_6401,N_7398);
nor U12065 (N_12065,N_8191,N_8223);
or U12066 (N_12066,N_8644,N_8633);
or U12067 (N_12067,N_7841,N_8317);
nand U12068 (N_12068,N_7301,N_6274);
or U12069 (N_12069,N_6589,N_8498);
or U12070 (N_12070,N_7961,N_6461);
nor U12071 (N_12071,N_8778,N_8437);
nand U12072 (N_12072,N_6587,N_7862);
or U12073 (N_12073,N_8795,N_7952);
nand U12074 (N_12074,N_9200,N_7496);
nand U12075 (N_12075,N_9097,N_7027);
or U12076 (N_12076,N_9132,N_6975);
nor U12077 (N_12077,N_7311,N_6788);
nor U12078 (N_12078,N_7313,N_7987);
or U12079 (N_12079,N_7190,N_9090);
and U12080 (N_12080,N_7307,N_7001);
nor U12081 (N_12081,N_8027,N_7394);
and U12082 (N_12082,N_7171,N_7907);
or U12083 (N_12083,N_6817,N_8604);
or U12084 (N_12084,N_7641,N_8365);
xnor U12085 (N_12085,N_9044,N_7268);
nor U12086 (N_12086,N_8988,N_7009);
nor U12087 (N_12087,N_6532,N_8763);
nor U12088 (N_12088,N_9284,N_6275);
and U12089 (N_12089,N_7090,N_8937);
nand U12090 (N_12090,N_8953,N_7768);
or U12091 (N_12091,N_7032,N_9110);
xor U12092 (N_12092,N_8803,N_6769);
or U12093 (N_12093,N_8809,N_8561);
and U12094 (N_12094,N_6436,N_7571);
or U12095 (N_12095,N_8360,N_9141);
and U12096 (N_12096,N_9074,N_7189);
nor U12097 (N_12097,N_9230,N_7193);
nand U12098 (N_12098,N_9079,N_7076);
or U12099 (N_12099,N_7048,N_7607);
nand U12100 (N_12100,N_7141,N_8657);
nor U12101 (N_12101,N_9230,N_8202);
nor U12102 (N_12102,N_8965,N_6338);
nand U12103 (N_12103,N_6333,N_7162);
nand U12104 (N_12104,N_7954,N_6909);
and U12105 (N_12105,N_7322,N_6259);
or U12106 (N_12106,N_7890,N_9076);
nand U12107 (N_12107,N_8795,N_6798);
or U12108 (N_12108,N_6329,N_7040);
and U12109 (N_12109,N_7183,N_8500);
nor U12110 (N_12110,N_9298,N_8324);
and U12111 (N_12111,N_7332,N_7735);
and U12112 (N_12112,N_9149,N_8278);
nand U12113 (N_12113,N_8066,N_7290);
and U12114 (N_12114,N_7136,N_7864);
and U12115 (N_12115,N_6412,N_9240);
xnor U12116 (N_12116,N_9034,N_7533);
nor U12117 (N_12117,N_9151,N_7628);
and U12118 (N_12118,N_9006,N_6517);
nor U12119 (N_12119,N_9173,N_8522);
and U12120 (N_12120,N_6515,N_6770);
and U12121 (N_12121,N_6696,N_7977);
nor U12122 (N_12122,N_8431,N_7368);
and U12123 (N_12123,N_9106,N_7697);
and U12124 (N_12124,N_8206,N_8100);
nor U12125 (N_12125,N_7299,N_9004);
or U12126 (N_12126,N_6276,N_9354);
nor U12127 (N_12127,N_6687,N_8811);
nor U12128 (N_12128,N_7761,N_7196);
xnor U12129 (N_12129,N_7712,N_6747);
nand U12130 (N_12130,N_8252,N_8329);
nand U12131 (N_12131,N_6797,N_7498);
or U12132 (N_12132,N_9027,N_6597);
and U12133 (N_12133,N_6395,N_6250);
and U12134 (N_12134,N_7025,N_7801);
nand U12135 (N_12135,N_7802,N_6435);
or U12136 (N_12136,N_8573,N_7569);
and U12137 (N_12137,N_8414,N_8851);
and U12138 (N_12138,N_7211,N_7297);
nand U12139 (N_12139,N_8035,N_6389);
and U12140 (N_12140,N_7273,N_9244);
nor U12141 (N_12141,N_6990,N_8126);
nand U12142 (N_12142,N_8203,N_6803);
nor U12143 (N_12143,N_8563,N_6968);
xnor U12144 (N_12144,N_6826,N_6724);
or U12145 (N_12145,N_6866,N_7341);
nand U12146 (N_12146,N_7735,N_7676);
nand U12147 (N_12147,N_6546,N_8164);
nand U12148 (N_12148,N_9015,N_8344);
and U12149 (N_12149,N_8443,N_6492);
and U12150 (N_12150,N_6664,N_7369);
and U12151 (N_12151,N_8520,N_6684);
xnor U12152 (N_12152,N_7597,N_6570);
and U12153 (N_12153,N_7612,N_7647);
or U12154 (N_12154,N_8823,N_8536);
nor U12155 (N_12155,N_7038,N_7674);
or U12156 (N_12156,N_7415,N_7965);
nand U12157 (N_12157,N_8944,N_9032);
or U12158 (N_12158,N_6903,N_7512);
nor U12159 (N_12159,N_8023,N_8176);
and U12160 (N_12160,N_7347,N_6936);
and U12161 (N_12161,N_8271,N_8448);
nor U12162 (N_12162,N_7637,N_9362);
nor U12163 (N_12163,N_8666,N_9217);
nor U12164 (N_12164,N_7963,N_8618);
and U12165 (N_12165,N_6286,N_6780);
and U12166 (N_12166,N_8304,N_8875);
xnor U12167 (N_12167,N_6325,N_7283);
or U12168 (N_12168,N_6441,N_7434);
nand U12169 (N_12169,N_7318,N_7746);
and U12170 (N_12170,N_8628,N_8111);
or U12171 (N_12171,N_9264,N_7627);
xnor U12172 (N_12172,N_7111,N_9012);
or U12173 (N_12173,N_8578,N_7001);
nand U12174 (N_12174,N_8293,N_7518);
nor U12175 (N_12175,N_7707,N_8470);
and U12176 (N_12176,N_8328,N_7318);
nand U12177 (N_12177,N_9360,N_8278);
nor U12178 (N_12178,N_7589,N_7164);
nand U12179 (N_12179,N_8499,N_7491);
or U12180 (N_12180,N_6390,N_6338);
and U12181 (N_12181,N_9139,N_6437);
xnor U12182 (N_12182,N_6488,N_8464);
nand U12183 (N_12183,N_7098,N_7733);
nor U12184 (N_12184,N_7444,N_6899);
nor U12185 (N_12185,N_8539,N_7889);
or U12186 (N_12186,N_8649,N_7301);
nor U12187 (N_12187,N_8065,N_9069);
nor U12188 (N_12188,N_6862,N_7899);
or U12189 (N_12189,N_9192,N_8445);
nor U12190 (N_12190,N_8122,N_6662);
or U12191 (N_12191,N_7170,N_7790);
nand U12192 (N_12192,N_6891,N_6551);
and U12193 (N_12193,N_6951,N_6988);
or U12194 (N_12194,N_8207,N_7414);
or U12195 (N_12195,N_8759,N_8491);
nand U12196 (N_12196,N_9013,N_8435);
or U12197 (N_12197,N_6718,N_8418);
nand U12198 (N_12198,N_8715,N_8142);
nor U12199 (N_12199,N_8055,N_9273);
and U12200 (N_12200,N_9100,N_8436);
and U12201 (N_12201,N_7680,N_6691);
nand U12202 (N_12202,N_9262,N_8508);
and U12203 (N_12203,N_7847,N_8426);
and U12204 (N_12204,N_7248,N_6748);
or U12205 (N_12205,N_6342,N_7826);
xnor U12206 (N_12206,N_7604,N_6314);
and U12207 (N_12207,N_8127,N_9168);
nor U12208 (N_12208,N_7661,N_9277);
or U12209 (N_12209,N_6902,N_6538);
nand U12210 (N_12210,N_8018,N_6877);
and U12211 (N_12211,N_9079,N_6991);
or U12212 (N_12212,N_6665,N_7517);
nor U12213 (N_12213,N_7939,N_7037);
and U12214 (N_12214,N_7553,N_8055);
nand U12215 (N_12215,N_8063,N_7862);
xnor U12216 (N_12216,N_8317,N_8185);
nor U12217 (N_12217,N_7229,N_8649);
nand U12218 (N_12218,N_9091,N_8303);
or U12219 (N_12219,N_9263,N_9243);
nor U12220 (N_12220,N_7071,N_7087);
nand U12221 (N_12221,N_7317,N_7334);
nand U12222 (N_12222,N_9209,N_6756);
or U12223 (N_12223,N_7677,N_7288);
and U12224 (N_12224,N_7836,N_7591);
or U12225 (N_12225,N_8331,N_7734);
and U12226 (N_12226,N_8326,N_7857);
nand U12227 (N_12227,N_6921,N_6509);
nand U12228 (N_12228,N_9359,N_6718);
nor U12229 (N_12229,N_7064,N_6793);
or U12230 (N_12230,N_9248,N_8283);
nand U12231 (N_12231,N_7256,N_6501);
or U12232 (N_12232,N_6713,N_7010);
nand U12233 (N_12233,N_7435,N_7921);
nor U12234 (N_12234,N_6347,N_9229);
nand U12235 (N_12235,N_8069,N_9042);
nor U12236 (N_12236,N_7351,N_7100);
nand U12237 (N_12237,N_8756,N_8225);
nor U12238 (N_12238,N_8187,N_8126);
or U12239 (N_12239,N_7730,N_8176);
nand U12240 (N_12240,N_6604,N_9173);
nor U12241 (N_12241,N_8436,N_7713);
or U12242 (N_12242,N_6928,N_9079);
and U12243 (N_12243,N_6537,N_7209);
nand U12244 (N_12244,N_8858,N_7041);
and U12245 (N_12245,N_6748,N_8266);
nor U12246 (N_12246,N_8974,N_6915);
and U12247 (N_12247,N_7499,N_7724);
and U12248 (N_12248,N_7837,N_8198);
nor U12249 (N_12249,N_7853,N_6269);
nor U12250 (N_12250,N_6604,N_9096);
nand U12251 (N_12251,N_8815,N_7210);
nand U12252 (N_12252,N_7623,N_6448);
nand U12253 (N_12253,N_7522,N_6425);
xnor U12254 (N_12254,N_6594,N_9250);
or U12255 (N_12255,N_9152,N_8533);
or U12256 (N_12256,N_6436,N_8030);
nand U12257 (N_12257,N_6952,N_6306);
or U12258 (N_12258,N_8433,N_9252);
xnor U12259 (N_12259,N_7021,N_6739);
or U12260 (N_12260,N_6447,N_8221);
or U12261 (N_12261,N_7101,N_6608);
nand U12262 (N_12262,N_8388,N_8270);
or U12263 (N_12263,N_7905,N_7854);
or U12264 (N_12264,N_7885,N_7700);
nor U12265 (N_12265,N_6835,N_6693);
or U12266 (N_12266,N_7701,N_8351);
nand U12267 (N_12267,N_8760,N_8614);
or U12268 (N_12268,N_6398,N_8810);
and U12269 (N_12269,N_8381,N_8135);
or U12270 (N_12270,N_8016,N_7363);
nand U12271 (N_12271,N_7854,N_7427);
or U12272 (N_12272,N_6286,N_8633);
or U12273 (N_12273,N_9222,N_7265);
and U12274 (N_12274,N_8594,N_9312);
nand U12275 (N_12275,N_7532,N_7356);
or U12276 (N_12276,N_7956,N_7008);
and U12277 (N_12277,N_9154,N_9265);
or U12278 (N_12278,N_7062,N_7004);
nor U12279 (N_12279,N_7818,N_8065);
nor U12280 (N_12280,N_7481,N_7447);
xor U12281 (N_12281,N_6561,N_8850);
or U12282 (N_12282,N_8437,N_7098);
nand U12283 (N_12283,N_8421,N_7544);
and U12284 (N_12284,N_7530,N_8482);
or U12285 (N_12285,N_8965,N_8256);
nor U12286 (N_12286,N_8082,N_6970);
nor U12287 (N_12287,N_7345,N_8670);
or U12288 (N_12288,N_7828,N_7218);
or U12289 (N_12289,N_6843,N_8647);
nand U12290 (N_12290,N_6688,N_6746);
nand U12291 (N_12291,N_6411,N_7166);
nand U12292 (N_12292,N_6923,N_8818);
nand U12293 (N_12293,N_8328,N_7024);
and U12294 (N_12294,N_6258,N_7933);
nor U12295 (N_12295,N_7931,N_9247);
or U12296 (N_12296,N_7192,N_6725);
or U12297 (N_12297,N_6902,N_7321);
or U12298 (N_12298,N_9308,N_7015);
nor U12299 (N_12299,N_6534,N_6395);
or U12300 (N_12300,N_7376,N_7558);
or U12301 (N_12301,N_6483,N_8594);
nor U12302 (N_12302,N_9165,N_7746);
xnor U12303 (N_12303,N_9272,N_6781);
and U12304 (N_12304,N_6526,N_8045);
or U12305 (N_12305,N_8341,N_9211);
and U12306 (N_12306,N_9113,N_7759);
nor U12307 (N_12307,N_7815,N_7749);
xnor U12308 (N_12308,N_6409,N_7933);
nand U12309 (N_12309,N_8710,N_8492);
and U12310 (N_12310,N_6360,N_7625);
nand U12311 (N_12311,N_8001,N_8190);
or U12312 (N_12312,N_7297,N_8343);
nand U12313 (N_12313,N_8073,N_7374);
or U12314 (N_12314,N_8878,N_7653);
and U12315 (N_12315,N_6881,N_8465);
or U12316 (N_12316,N_9342,N_7786);
nor U12317 (N_12317,N_8302,N_6265);
or U12318 (N_12318,N_7520,N_9020);
nor U12319 (N_12319,N_8800,N_8746);
and U12320 (N_12320,N_6837,N_6879);
or U12321 (N_12321,N_6986,N_7650);
or U12322 (N_12322,N_7555,N_8778);
nand U12323 (N_12323,N_8649,N_7923);
and U12324 (N_12324,N_6914,N_8540);
nand U12325 (N_12325,N_7958,N_7480);
or U12326 (N_12326,N_7940,N_9187);
nor U12327 (N_12327,N_9322,N_6942);
or U12328 (N_12328,N_8939,N_8021);
nor U12329 (N_12329,N_8821,N_9105);
and U12330 (N_12330,N_6711,N_7906);
nand U12331 (N_12331,N_8130,N_9021);
and U12332 (N_12332,N_7943,N_8247);
or U12333 (N_12333,N_7196,N_7633);
and U12334 (N_12334,N_7680,N_8239);
nand U12335 (N_12335,N_8147,N_8808);
and U12336 (N_12336,N_8186,N_6917);
xor U12337 (N_12337,N_7799,N_8095);
and U12338 (N_12338,N_7540,N_6353);
and U12339 (N_12339,N_8271,N_7923);
or U12340 (N_12340,N_8634,N_8458);
or U12341 (N_12341,N_8760,N_7072);
nor U12342 (N_12342,N_6315,N_7554);
or U12343 (N_12343,N_9067,N_8009);
nand U12344 (N_12344,N_6914,N_6305);
nor U12345 (N_12345,N_8138,N_6795);
nor U12346 (N_12346,N_7242,N_6479);
and U12347 (N_12347,N_7640,N_8978);
nor U12348 (N_12348,N_6616,N_9040);
nand U12349 (N_12349,N_8835,N_8724);
nor U12350 (N_12350,N_8023,N_7808);
xor U12351 (N_12351,N_8005,N_8207);
or U12352 (N_12352,N_8981,N_6756);
nand U12353 (N_12353,N_6271,N_7949);
xnor U12354 (N_12354,N_7870,N_7589);
nor U12355 (N_12355,N_7745,N_8793);
nor U12356 (N_12356,N_9027,N_7276);
nand U12357 (N_12357,N_6629,N_6606);
or U12358 (N_12358,N_7008,N_9295);
nand U12359 (N_12359,N_7925,N_7823);
nand U12360 (N_12360,N_6795,N_7825);
xor U12361 (N_12361,N_7287,N_8128);
nor U12362 (N_12362,N_6989,N_8397);
and U12363 (N_12363,N_6936,N_6356);
nor U12364 (N_12364,N_8792,N_8021);
and U12365 (N_12365,N_6507,N_8493);
nor U12366 (N_12366,N_8205,N_8117);
and U12367 (N_12367,N_7453,N_9047);
and U12368 (N_12368,N_6655,N_7426);
nor U12369 (N_12369,N_8266,N_8519);
nand U12370 (N_12370,N_8462,N_7804);
or U12371 (N_12371,N_8486,N_8395);
or U12372 (N_12372,N_7334,N_8010);
nor U12373 (N_12373,N_7135,N_6570);
and U12374 (N_12374,N_6601,N_7112);
nand U12375 (N_12375,N_6616,N_6348);
or U12376 (N_12376,N_9308,N_6856);
and U12377 (N_12377,N_8911,N_7988);
and U12378 (N_12378,N_7069,N_8386);
nand U12379 (N_12379,N_6891,N_9333);
or U12380 (N_12380,N_8400,N_8736);
nor U12381 (N_12381,N_7710,N_8067);
nand U12382 (N_12382,N_7721,N_7627);
nor U12383 (N_12383,N_8793,N_9093);
nand U12384 (N_12384,N_9181,N_7760);
or U12385 (N_12385,N_7462,N_8003);
xnor U12386 (N_12386,N_7793,N_8632);
nand U12387 (N_12387,N_7730,N_8611);
or U12388 (N_12388,N_8036,N_7351);
xor U12389 (N_12389,N_6520,N_7761);
and U12390 (N_12390,N_7800,N_8989);
and U12391 (N_12391,N_6593,N_9247);
nand U12392 (N_12392,N_9315,N_7790);
xnor U12393 (N_12393,N_9043,N_6485);
or U12394 (N_12394,N_7286,N_7120);
nand U12395 (N_12395,N_7120,N_7878);
nor U12396 (N_12396,N_8023,N_7478);
nor U12397 (N_12397,N_8296,N_7356);
nand U12398 (N_12398,N_8273,N_8582);
and U12399 (N_12399,N_8713,N_6854);
nand U12400 (N_12400,N_6434,N_6629);
nor U12401 (N_12401,N_8933,N_7382);
and U12402 (N_12402,N_6302,N_7527);
or U12403 (N_12403,N_7252,N_7532);
or U12404 (N_12404,N_7317,N_9359);
or U12405 (N_12405,N_6722,N_6770);
or U12406 (N_12406,N_6793,N_8517);
and U12407 (N_12407,N_8477,N_9260);
xnor U12408 (N_12408,N_8308,N_9020);
xor U12409 (N_12409,N_8126,N_8477);
nand U12410 (N_12410,N_8672,N_7693);
nand U12411 (N_12411,N_6772,N_7736);
and U12412 (N_12412,N_6991,N_6968);
xor U12413 (N_12413,N_6881,N_6819);
or U12414 (N_12414,N_6332,N_6712);
and U12415 (N_12415,N_7472,N_6651);
xor U12416 (N_12416,N_9278,N_9031);
or U12417 (N_12417,N_7217,N_7238);
or U12418 (N_12418,N_6998,N_8056);
xor U12419 (N_12419,N_7307,N_9085);
nor U12420 (N_12420,N_6687,N_7084);
and U12421 (N_12421,N_8769,N_6513);
nor U12422 (N_12422,N_6323,N_7746);
nand U12423 (N_12423,N_9341,N_7429);
or U12424 (N_12424,N_8041,N_7294);
nand U12425 (N_12425,N_6642,N_8295);
nor U12426 (N_12426,N_7715,N_7582);
and U12427 (N_12427,N_8077,N_8684);
nor U12428 (N_12428,N_9165,N_6479);
and U12429 (N_12429,N_7390,N_7494);
nand U12430 (N_12430,N_6264,N_7211);
nand U12431 (N_12431,N_8401,N_9011);
or U12432 (N_12432,N_6517,N_6796);
and U12433 (N_12433,N_8462,N_8504);
nand U12434 (N_12434,N_7256,N_7831);
or U12435 (N_12435,N_9066,N_8773);
or U12436 (N_12436,N_7300,N_6827);
or U12437 (N_12437,N_7478,N_7535);
nor U12438 (N_12438,N_8223,N_8288);
and U12439 (N_12439,N_7552,N_6330);
nand U12440 (N_12440,N_8086,N_7985);
or U12441 (N_12441,N_8567,N_9368);
or U12442 (N_12442,N_8117,N_6769);
nand U12443 (N_12443,N_7331,N_6593);
and U12444 (N_12444,N_8276,N_8138);
and U12445 (N_12445,N_6393,N_6811);
and U12446 (N_12446,N_8407,N_7256);
or U12447 (N_12447,N_6687,N_8789);
and U12448 (N_12448,N_6532,N_6319);
nand U12449 (N_12449,N_6450,N_6365);
and U12450 (N_12450,N_8725,N_6723);
nand U12451 (N_12451,N_8906,N_8165);
xor U12452 (N_12452,N_6418,N_8776);
xor U12453 (N_12453,N_7253,N_7225);
and U12454 (N_12454,N_8465,N_8238);
nand U12455 (N_12455,N_8167,N_9355);
nand U12456 (N_12456,N_6565,N_8886);
nor U12457 (N_12457,N_7698,N_6831);
nand U12458 (N_12458,N_8352,N_8698);
nor U12459 (N_12459,N_9358,N_8391);
nand U12460 (N_12460,N_9165,N_6836);
and U12461 (N_12461,N_8996,N_8402);
nand U12462 (N_12462,N_6370,N_9057);
xnor U12463 (N_12463,N_8610,N_6346);
nand U12464 (N_12464,N_7561,N_8553);
and U12465 (N_12465,N_7055,N_8929);
and U12466 (N_12466,N_7364,N_9183);
and U12467 (N_12467,N_8123,N_8571);
or U12468 (N_12468,N_9232,N_6813);
and U12469 (N_12469,N_8060,N_7083);
or U12470 (N_12470,N_7166,N_7876);
nor U12471 (N_12471,N_8203,N_8072);
or U12472 (N_12472,N_7862,N_7354);
nand U12473 (N_12473,N_7767,N_9009);
nor U12474 (N_12474,N_7470,N_6991);
or U12475 (N_12475,N_8181,N_7675);
nand U12476 (N_12476,N_9291,N_8811);
and U12477 (N_12477,N_7565,N_7194);
or U12478 (N_12478,N_8476,N_6436);
or U12479 (N_12479,N_6903,N_7415);
nor U12480 (N_12480,N_8004,N_6377);
nand U12481 (N_12481,N_8844,N_9087);
and U12482 (N_12482,N_7975,N_7471);
nand U12483 (N_12483,N_7181,N_7145);
or U12484 (N_12484,N_8999,N_8051);
nor U12485 (N_12485,N_8839,N_8714);
and U12486 (N_12486,N_9138,N_6571);
or U12487 (N_12487,N_6756,N_6937);
xor U12488 (N_12488,N_8031,N_8173);
or U12489 (N_12489,N_8677,N_8931);
and U12490 (N_12490,N_8501,N_9323);
xor U12491 (N_12491,N_8026,N_8731);
xor U12492 (N_12492,N_8272,N_6267);
nor U12493 (N_12493,N_6330,N_6286);
nand U12494 (N_12494,N_6674,N_7400);
xnor U12495 (N_12495,N_7501,N_8198);
or U12496 (N_12496,N_6481,N_8138);
nand U12497 (N_12497,N_8504,N_6715);
nand U12498 (N_12498,N_7067,N_6732);
nand U12499 (N_12499,N_8754,N_8482);
and U12500 (N_12500,N_9410,N_10293);
nor U12501 (N_12501,N_12118,N_9542);
and U12502 (N_12502,N_10579,N_11611);
nand U12503 (N_12503,N_11959,N_9898);
nor U12504 (N_12504,N_11974,N_12413);
nor U12505 (N_12505,N_9647,N_11324);
nor U12506 (N_12506,N_9727,N_12164);
nor U12507 (N_12507,N_9512,N_11049);
nand U12508 (N_12508,N_11635,N_9871);
xor U12509 (N_12509,N_11864,N_10511);
or U12510 (N_12510,N_9841,N_11646);
or U12511 (N_12511,N_10074,N_9428);
or U12512 (N_12512,N_12080,N_10157);
or U12513 (N_12513,N_11528,N_11020);
nor U12514 (N_12514,N_11856,N_11709);
or U12515 (N_12515,N_10323,N_10077);
or U12516 (N_12516,N_9847,N_9579);
or U12517 (N_12517,N_10936,N_12354);
or U12518 (N_12518,N_11209,N_10634);
and U12519 (N_12519,N_10126,N_9897);
and U12520 (N_12520,N_11792,N_10431);
nor U12521 (N_12521,N_10999,N_12220);
nor U12522 (N_12522,N_11417,N_10558);
nor U12523 (N_12523,N_9610,N_11796);
or U12524 (N_12524,N_9786,N_9617);
nand U12525 (N_12525,N_12036,N_9738);
or U12526 (N_12526,N_10757,N_9588);
nand U12527 (N_12527,N_12204,N_11907);
nand U12528 (N_12528,N_11036,N_9524);
or U12529 (N_12529,N_11352,N_10636);
nand U12530 (N_12530,N_12134,N_10540);
and U12531 (N_12531,N_11575,N_11519);
xor U12532 (N_12532,N_11463,N_9711);
and U12533 (N_12533,N_9824,N_9714);
or U12534 (N_12534,N_10422,N_11403);
or U12535 (N_12535,N_11906,N_12451);
nor U12536 (N_12536,N_11683,N_10115);
or U12537 (N_12537,N_10060,N_9555);
or U12538 (N_12538,N_12205,N_12092);
nor U12539 (N_12539,N_12446,N_10080);
and U12540 (N_12540,N_9845,N_11250);
and U12541 (N_12541,N_12210,N_10568);
or U12542 (N_12542,N_11424,N_11069);
or U12543 (N_12543,N_12287,N_12110);
nand U12544 (N_12544,N_10976,N_10038);
or U12545 (N_12545,N_10406,N_12291);
nand U12546 (N_12546,N_9816,N_12111);
nor U12547 (N_12547,N_11487,N_11929);
and U12548 (N_12548,N_11775,N_12388);
and U12549 (N_12549,N_10905,N_11493);
nand U12550 (N_12550,N_11068,N_10090);
nand U12551 (N_12551,N_11261,N_10529);
or U12552 (N_12552,N_12441,N_11938);
nand U12553 (N_12553,N_12131,N_11479);
xor U12554 (N_12554,N_11602,N_10466);
and U12555 (N_12555,N_12012,N_9820);
nor U12556 (N_12556,N_11383,N_12297);
nand U12557 (N_12557,N_11599,N_12495);
nand U12558 (N_12558,N_11946,N_10029);
and U12559 (N_12559,N_10191,N_10164);
and U12560 (N_12560,N_11283,N_11983);
xnor U12561 (N_12561,N_11244,N_11146);
nor U12562 (N_12562,N_10792,N_10723);
nor U12563 (N_12563,N_12145,N_9656);
nand U12564 (N_12564,N_10276,N_9537);
or U12565 (N_12565,N_11445,N_11640);
nor U12566 (N_12566,N_12469,N_9722);
or U12567 (N_12567,N_10174,N_10317);
nor U12568 (N_12568,N_9913,N_11208);
and U12569 (N_12569,N_12307,N_9511);
nand U12570 (N_12570,N_9639,N_10853);
nand U12571 (N_12571,N_12417,N_12265);
or U12572 (N_12572,N_12169,N_11106);
nor U12573 (N_12573,N_10530,N_10050);
nand U12574 (N_12574,N_11287,N_9960);
and U12575 (N_12575,N_11758,N_12168);
and U12576 (N_12576,N_10461,N_11960);
and U12577 (N_12577,N_11355,N_11369);
nand U12578 (N_12578,N_12112,N_10374);
nor U12579 (N_12579,N_10385,N_11260);
and U12580 (N_12580,N_12200,N_11667);
nand U12581 (N_12581,N_11211,N_9403);
or U12582 (N_12582,N_11668,N_12207);
xnor U12583 (N_12583,N_10852,N_10479);
and U12584 (N_12584,N_11399,N_9645);
and U12585 (N_12585,N_9809,N_12258);
nand U12586 (N_12586,N_11894,N_9783);
nor U12587 (N_12587,N_9942,N_11536);
xnor U12588 (N_12588,N_11892,N_11913);
nand U12589 (N_12589,N_12459,N_9605);
and U12590 (N_12590,N_11825,N_9583);
xor U12591 (N_12591,N_9706,N_10549);
and U12592 (N_12592,N_12418,N_11924);
nor U12593 (N_12593,N_10205,N_12453);
or U12594 (N_12594,N_11300,N_12242);
and U12595 (N_12595,N_11844,N_11425);
and U12596 (N_12596,N_10279,N_10150);
or U12597 (N_12597,N_10575,N_10800);
and U12598 (N_12598,N_9975,N_10469);
nor U12599 (N_12599,N_10261,N_12032);
nor U12600 (N_12600,N_12030,N_11060);
or U12601 (N_12601,N_10761,N_11077);
or U12602 (N_12602,N_11502,N_9859);
and U12603 (N_12603,N_12487,N_9480);
or U12604 (N_12604,N_12363,N_11473);
nor U12605 (N_12605,N_10501,N_12248);
nor U12606 (N_12606,N_11524,N_10448);
or U12607 (N_12607,N_9996,N_10547);
nand U12608 (N_12608,N_12055,N_11948);
or U12609 (N_12609,N_10860,N_10127);
and U12610 (N_12610,N_9799,N_11172);
nand U12611 (N_12611,N_11375,N_11347);
or U12612 (N_12612,N_12481,N_11409);
or U12613 (N_12613,N_10352,N_9528);
nor U12614 (N_12614,N_12311,N_10232);
or U12615 (N_12615,N_9762,N_11663);
or U12616 (N_12616,N_11122,N_11632);
xor U12617 (N_12617,N_12347,N_11530);
and U12618 (N_12618,N_9592,N_10846);
xor U12619 (N_12619,N_12235,N_11510);
and U12620 (N_12620,N_10697,N_9586);
or U12621 (N_12621,N_11943,N_11870);
or U12622 (N_12622,N_11291,N_11500);
xor U12623 (N_12623,N_12218,N_10245);
or U12624 (N_12624,N_9467,N_11328);
or U12625 (N_12625,N_12485,N_11379);
and U12626 (N_12626,N_10661,N_9736);
and U12627 (N_12627,N_10780,N_11017);
nor U12628 (N_12628,N_10503,N_11206);
and U12629 (N_12629,N_11645,N_10553);
and U12630 (N_12630,N_10649,N_10361);
nor U12631 (N_12631,N_11176,N_10358);
nor U12632 (N_12632,N_9676,N_10236);
nand U12633 (N_12633,N_10504,N_9958);
nand U12634 (N_12634,N_11367,N_10766);
nor U12635 (N_12635,N_11885,N_9563);
and U12636 (N_12636,N_10637,N_10909);
nand U12637 (N_12637,N_11656,N_10414);
xor U12638 (N_12638,N_10024,N_9657);
nor U12639 (N_12639,N_12249,N_9532);
or U12640 (N_12640,N_9462,N_12183);
xnor U12641 (N_12641,N_10147,N_10367);
and U12642 (N_12642,N_12197,N_10769);
or U12643 (N_12643,N_9981,N_11295);
and U12644 (N_12644,N_10326,N_11790);
or U12645 (N_12645,N_11034,N_10110);
or U12646 (N_12646,N_11489,N_9490);
or U12647 (N_12647,N_10678,N_11609);
nor U12648 (N_12648,N_10179,N_10258);
nor U12649 (N_12649,N_11769,N_10671);
nor U12650 (N_12650,N_9572,N_9417);
or U12651 (N_12651,N_9827,N_11135);
xnor U12652 (N_12652,N_9858,N_11706);
or U12653 (N_12653,N_11033,N_11224);
nor U12654 (N_12654,N_11939,N_10295);
and U12655 (N_12655,N_9932,N_11021);
or U12656 (N_12656,N_9911,N_9468);
nor U12657 (N_12657,N_10880,N_10351);
xor U12658 (N_12658,N_10460,N_12040);
or U12659 (N_12659,N_12116,N_10524);
and U12660 (N_12660,N_11361,N_11827);
and U12661 (N_12661,N_10019,N_9589);
nand U12662 (N_12662,N_9398,N_10322);
or U12663 (N_12663,N_11980,N_10305);
and U12664 (N_12664,N_12463,N_12185);
nand U12665 (N_12665,N_12011,N_10920);
or U12666 (N_12666,N_12295,N_10531);
xnor U12667 (N_12667,N_10874,N_10794);
nor U12668 (N_12668,N_9479,N_10864);
nand U12669 (N_12669,N_10255,N_10263);
nor U12670 (N_12670,N_10200,N_11183);
nor U12671 (N_12671,N_10394,N_12428);
and U12672 (N_12672,N_11171,N_10892);
or U12673 (N_12673,N_12091,N_9392);
or U12674 (N_12674,N_11826,N_9884);
nor U12675 (N_12675,N_9716,N_10573);
xor U12676 (N_12676,N_9574,N_12304);
or U12677 (N_12677,N_9650,N_10949);
and U12678 (N_12678,N_10228,N_10078);
nand U12679 (N_12679,N_9654,N_11065);
nand U12680 (N_12680,N_10546,N_11610);
and U12681 (N_12681,N_12315,N_10337);
nor U12682 (N_12682,N_10230,N_11574);
nand U12683 (N_12683,N_10243,N_9535);
or U12684 (N_12684,N_10881,N_10885);
and U12685 (N_12685,N_10362,N_9581);
nand U12686 (N_12686,N_10740,N_10070);
nor U12687 (N_12687,N_10388,N_12351);
nand U12688 (N_12688,N_10452,N_11623);
nand U12689 (N_12689,N_11321,N_9876);
or U12690 (N_12690,N_12400,N_11761);
nand U12691 (N_12691,N_11071,N_10590);
nor U12692 (N_12692,N_9780,N_9988);
and U12693 (N_12693,N_10870,N_12152);
or U12694 (N_12694,N_9702,N_11903);
xnor U12695 (N_12695,N_10162,N_12419);
nor U12696 (N_12696,N_11562,N_10459);
and U12697 (N_12697,N_11338,N_11062);
or U12698 (N_12698,N_10600,N_12216);
nand U12699 (N_12699,N_11205,N_11670);
and U12700 (N_12700,N_10525,N_10589);
nor U12701 (N_12701,N_10248,N_12394);
or U12702 (N_12702,N_12370,N_11253);
and U12703 (N_12703,N_12102,N_9851);
nand U12704 (N_12704,N_10030,N_11415);
or U12705 (N_12705,N_10328,N_10188);
nor U12706 (N_12706,N_10972,N_11503);
nor U12707 (N_12707,N_11927,N_11978);
and U12708 (N_12708,N_12461,N_11764);
nor U12709 (N_12709,N_9466,N_9606);
or U12710 (N_12710,N_11525,N_10166);
xor U12711 (N_12711,N_10533,N_12027);
and U12712 (N_12712,N_11850,N_10165);
and U12713 (N_12713,N_11830,N_10012);
nand U12714 (N_12714,N_10197,N_9611);
and U12715 (N_12715,N_10993,N_9566);
or U12716 (N_12716,N_10994,N_11437);
xnor U12717 (N_12717,N_11160,N_11809);
nand U12718 (N_12718,N_10873,N_11564);
or U12719 (N_12719,N_11351,N_10052);
and U12720 (N_12720,N_10268,N_11474);
and U12721 (N_12721,N_10376,N_9424);
xor U12722 (N_12722,N_10919,N_10576);
nand U12723 (N_12723,N_9507,N_12335);
or U12724 (N_12724,N_9927,N_9878);
xor U12725 (N_12725,N_10768,N_12142);
or U12726 (N_12726,N_11837,N_9472);
xor U12727 (N_12727,N_10064,N_12088);
or U12728 (N_12728,N_9798,N_11847);
and U12729 (N_12729,N_9698,N_12090);
and U12730 (N_12730,N_12044,N_11700);
nor U12731 (N_12731,N_9947,N_10476);
nor U12732 (N_12732,N_9890,N_10513);
or U12733 (N_12733,N_10206,N_10310);
xor U12734 (N_12734,N_11398,N_11451);
xor U12735 (N_12735,N_12137,N_9747);
nor U12736 (N_12736,N_11265,N_11123);
and U12737 (N_12737,N_11685,N_10798);
and U12738 (N_12738,N_12189,N_10101);
and U12739 (N_12739,N_10221,N_12293);
and U12740 (N_12740,N_12028,N_12380);
nor U12741 (N_12741,N_11374,N_11388);
nor U12742 (N_12742,N_11155,N_9648);
xnor U12743 (N_12743,N_9997,N_11391);
nor U12744 (N_12744,N_12119,N_11288);
nor U12745 (N_12745,N_9935,N_10325);
or U12746 (N_12746,N_11157,N_10336);
nor U12747 (N_12747,N_10446,N_12299);
nand U12748 (N_12748,N_11711,N_9561);
and U12749 (N_12749,N_11325,N_10789);
nor U12750 (N_12750,N_9458,N_12136);
or U12751 (N_12751,N_10148,N_10534);
or U12752 (N_12752,N_10722,N_12113);
and U12753 (N_12753,N_9705,N_11832);
or U12754 (N_12754,N_10105,N_12155);
and U12755 (N_12755,N_11026,N_12224);
and U12756 (N_12756,N_9986,N_12236);
nor U12757 (N_12757,N_11133,N_10537);
and U12758 (N_12758,N_10380,N_9642);
or U12759 (N_12759,N_10063,N_10630);
or U12760 (N_12760,N_11006,N_10833);
or U12761 (N_12761,N_11705,N_10495);
or U12762 (N_12762,N_11882,N_10283);
nand U12763 (N_12763,N_11795,N_11412);
nand U12764 (N_12764,N_9517,N_10492);
nand U12765 (N_12765,N_9644,N_10721);
or U12766 (N_12766,N_11331,N_9452);
nor U12767 (N_12767,N_11613,N_10412);
nand U12768 (N_12768,N_9630,N_10507);
nor U12769 (N_12769,N_9697,N_11266);
and U12770 (N_12770,N_10342,N_12029);
or U12771 (N_12771,N_10658,N_12460);
nand U12772 (N_12772,N_10175,N_11993);
xnor U12773 (N_12773,N_10932,N_9487);
nor U12774 (N_12774,N_12156,N_11967);
nand U12775 (N_12775,N_12133,N_12383);
nor U12776 (N_12776,N_12273,N_10552);
or U12777 (N_12777,N_11109,N_10208);
or U12778 (N_12778,N_10314,N_10582);
xnor U12779 (N_12779,N_11087,N_10257);
xnor U12780 (N_12780,N_11693,N_9513);
nand U12781 (N_12781,N_10122,N_9712);
and U12782 (N_12782,N_12252,N_10081);
xnor U12783 (N_12783,N_10004,N_11333);
and U12784 (N_12784,N_9916,N_9771);
nor U12785 (N_12785,N_10650,N_11053);
and U12786 (N_12786,N_11050,N_11431);
xnor U12787 (N_12787,N_10787,N_10424);
xnor U12788 (N_12788,N_9476,N_10333);
nor U12789 (N_12789,N_12073,N_10981);
nand U12790 (N_12790,N_12060,N_10581);
or U12791 (N_12791,N_12081,N_10320);
nor U12792 (N_12792,N_10416,N_12026);
nor U12793 (N_12793,N_11469,N_9545);
or U12794 (N_12794,N_9800,N_9971);
or U12795 (N_12795,N_11996,N_9686);
nand U12796 (N_12796,N_10031,N_11861);
or U12797 (N_12797,N_11901,N_10539);
or U12798 (N_12798,N_11440,N_12117);
nand U12799 (N_12799,N_12476,N_10714);
and U12800 (N_12800,N_10491,N_12283);
nand U12801 (N_12801,N_10824,N_9883);
and U12802 (N_12802,N_11771,N_9879);
nand U12803 (N_12803,N_10015,N_11900);
and U12804 (N_12804,N_9594,N_12284);
nor U12805 (N_12805,N_9618,N_11012);
nand U12806 (N_12806,N_9602,N_10938);
or U12807 (N_12807,N_10808,N_10904);
nand U12808 (N_12808,N_9739,N_9431);
or U12809 (N_12809,N_9502,N_11660);
and U12810 (N_12810,N_10494,N_10002);
or U12811 (N_12811,N_10851,N_10040);
or U12812 (N_12812,N_11499,N_10974);
nor U12813 (N_12813,N_11986,N_11047);
or U12814 (N_12814,N_10089,N_11849);
nand U12815 (N_12815,N_10251,N_11201);
or U12816 (N_12816,N_11551,N_12390);
and U12817 (N_12817,N_10646,N_11189);
nand U12818 (N_12818,N_10269,N_10401);
nor U12819 (N_12819,N_10304,N_11416);
nor U12820 (N_12820,N_11101,N_12456);
nor U12821 (N_12821,N_11975,N_9519);
nor U12822 (N_12822,N_12101,N_10644);
nor U12823 (N_12823,N_9673,N_9781);
or U12824 (N_12824,N_10975,N_10464);
and U12825 (N_12825,N_9941,N_11345);
and U12826 (N_12826,N_10706,N_9983);
or U12827 (N_12827,N_10350,N_11460);
nand U12828 (N_12828,N_12472,N_12322);
and U12829 (N_12829,N_9896,N_10729);
nor U12830 (N_12830,N_10843,N_11526);
and U12831 (N_12831,N_11905,N_9886);
or U12832 (N_12832,N_11968,N_11052);
or U12833 (N_12833,N_9386,N_9470);
and U12834 (N_12834,N_12443,N_9628);
nand U12835 (N_12835,N_10871,N_11937);
or U12836 (N_12836,N_9842,N_11802);
nand U12837 (N_12837,N_10161,N_11197);
xor U12838 (N_12838,N_10108,N_10502);
nand U12839 (N_12839,N_11397,N_10914);
xor U12840 (N_12840,N_12286,N_10647);
and U12841 (N_12841,N_11869,N_10397);
xor U12842 (N_12842,N_9929,N_11535);
nand U12843 (N_12843,N_10759,N_9797);
and U12844 (N_12844,N_11971,N_11357);
and U12845 (N_12845,N_12330,N_11322);
nor U12846 (N_12846,N_10596,N_9779);
or U12847 (N_12847,N_11027,N_12493);
or U12848 (N_12848,N_9742,N_10434);
nand U12849 (N_12849,N_11738,N_10672);
xor U12850 (N_12850,N_9641,N_12368);
nand U12851 (N_12851,N_9707,N_9668);
nor U12852 (N_12852,N_12176,N_11175);
nor U12853 (N_12853,N_9433,N_10519);
and U12854 (N_12854,N_10087,N_9399);
nand U12855 (N_12855,N_12375,N_10820);
and U12856 (N_12856,N_11079,N_10143);
nand U12857 (N_12857,N_11497,N_10942);
xnor U12858 (N_12858,N_11520,N_12182);
and U12859 (N_12859,N_9904,N_10447);
nand U12860 (N_12860,N_11957,N_12072);
nor U12861 (N_12861,N_10468,N_9378);
xor U12862 (N_12862,N_12320,N_9536);
nand U12863 (N_12863,N_11605,N_10571);
nand U12864 (N_12864,N_9471,N_11751);
nand U12865 (N_12865,N_10802,N_10605);
and U12866 (N_12866,N_12075,N_11787);
and U12867 (N_12867,N_12350,N_10347);
nor U12868 (N_12868,N_11332,N_10897);
xor U12869 (N_12869,N_10169,N_12396);
xnor U12870 (N_12870,N_9494,N_9939);
nor U12871 (N_12871,N_12438,N_11414);
and U12872 (N_12872,N_9732,N_11543);
or U12873 (N_12873,N_9749,N_11899);
or U12874 (N_12874,N_9559,N_9531);
nor U12875 (N_12875,N_9836,N_12229);
nor U12876 (N_12876,N_12243,N_12431);
xnor U12877 (N_12877,N_11945,N_11597);
or U12878 (N_12878,N_11498,N_9670);
or U12879 (N_12879,N_11982,N_10793);
nor U12880 (N_12880,N_12381,N_10044);
or U12881 (N_12881,N_10704,N_12093);
or U12882 (N_12882,N_11890,N_12361);
or U12883 (N_12883,N_12256,N_11721);
and U12884 (N_12884,N_10027,N_9597);
nor U12885 (N_12885,N_11363,N_12292);
nor U12886 (N_12886,N_9978,N_12069);
and U12887 (N_12887,N_12174,N_10804);
and U12888 (N_12888,N_11868,N_10713);
xnor U12889 (N_12889,N_10771,N_11167);
and U12890 (N_12890,N_10173,N_12192);
nor U12891 (N_12891,N_11581,N_10253);
nand U12892 (N_12892,N_12379,N_10371);
and U12893 (N_12893,N_10407,N_9867);
nand U12894 (N_12894,N_11539,N_11102);
nand U12895 (N_12895,N_9846,N_10739);
or U12896 (N_12896,N_9478,N_9539);
nand U12897 (N_12897,N_10982,N_10986);
nor U12898 (N_12898,N_12278,N_11675);
nand U12899 (N_12899,N_12349,N_11225);
nor U12900 (N_12900,N_9992,N_10271);
nor U12901 (N_12901,N_11478,N_11703);
nor U12902 (N_12902,N_10445,N_10086);
or U12903 (N_12903,N_10701,N_10542);
or U12904 (N_12904,N_10062,N_11521);
nand U12905 (N_12905,N_11243,N_9785);
or U12906 (N_12906,N_9773,N_10061);
nor U12907 (N_12907,N_10617,N_11271);
and U12908 (N_12908,N_11022,N_10439);
nor U12909 (N_12909,N_12448,N_9873);
and U12910 (N_12910,N_12475,N_12042);
xor U12911 (N_12911,N_9987,N_11737);
or U12912 (N_12912,N_9765,N_11335);
nand U12913 (N_12913,N_12314,N_11532);
or U12914 (N_12914,N_11296,N_11138);
nor U12915 (N_12915,N_10692,N_9903);
nor U12916 (N_12916,N_11215,N_12412);
xnor U12917 (N_12917,N_9991,N_10129);
or U12918 (N_12918,N_12313,N_10125);
or U12919 (N_12919,N_9989,N_10256);
nand U12920 (N_12920,N_12442,N_12135);
and U12921 (N_12921,N_9685,N_10487);
and U12922 (N_12922,N_9623,N_10598);
or U12923 (N_12923,N_10277,N_10896);
and U12924 (N_12924,N_10001,N_12035);
and U12925 (N_12925,N_11184,N_11672);
and U12926 (N_12926,N_10133,N_11916);
nand U12927 (N_12927,N_10396,N_10618);
and U12928 (N_12928,N_10807,N_11637);
xor U12929 (N_12929,N_12046,N_11237);
xnor U12930 (N_12930,N_9664,N_11435);
and U12931 (N_12931,N_9534,N_9844);
nor U12932 (N_12932,N_9681,N_9460);
and U12933 (N_12933,N_11105,N_9906);
nor U12934 (N_12934,N_11084,N_9750);
nand U12935 (N_12935,N_11893,N_9582);
nor U12936 (N_12936,N_9743,N_10267);
and U12937 (N_12937,N_11631,N_9769);
and U12938 (N_12938,N_9968,N_10033);
nand U12939 (N_12939,N_11098,N_9701);
xor U12940 (N_12940,N_12470,N_11279);
nand U12941 (N_12941,N_10883,N_10578);
and U12942 (N_12942,N_9447,N_11307);
and U12943 (N_12943,N_12408,N_12167);
nand U12944 (N_12944,N_11748,N_11720);
or U12945 (N_12945,N_10801,N_12141);
nor U12946 (N_12946,N_11633,N_10136);
xnor U12947 (N_12947,N_11236,N_12332);
nand U12948 (N_12948,N_9834,N_9729);
nor U12949 (N_12949,N_12409,N_11136);
xor U12950 (N_12950,N_12411,N_10130);
nor U12951 (N_12951,N_11152,N_9949);
nand U12952 (N_12952,N_10065,N_11545);
nor U12953 (N_12953,N_11185,N_11747);
nand U12954 (N_12954,N_12261,N_11559);
nor U12955 (N_12955,N_9857,N_9680);
or U12956 (N_12956,N_10499,N_9390);
and U12957 (N_12957,N_11652,N_9544);
or U12958 (N_12958,N_10670,N_11150);
and U12959 (N_12959,N_11954,N_9434);
or U12960 (N_12960,N_11746,N_10234);
nand U12961 (N_12961,N_12467,N_12397);
xnor U12962 (N_12962,N_10850,N_11895);
and U12963 (N_12963,N_12103,N_11735);
and U12964 (N_12964,N_11782,N_11380);
nor U12965 (N_12965,N_12083,N_11423);
or U12966 (N_12966,N_9870,N_11264);
and U12967 (N_12967,N_10049,N_10677);
and U12968 (N_12968,N_9416,N_12146);
nand U12969 (N_12969,N_10763,N_11793);
or U12970 (N_12970,N_11108,N_11577);
and U12971 (N_12971,N_11518,N_9877);
and U12972 (N_12972,N_10685,N_10470);
nor U12973 (N_12973,N_10222,N_11984);
nor U12974 (N_12974,N_9833,N_10948);
and U12975 (N_12975,N_9792,N_11411);
and U12976 (N_12976,N_12017,N_11789);
xnor U12977 (N_12977,N_11259,N_11915);
xnor U12978 (N_12978,N_9848,N_9804);
and U12979 (N_12979,N_10574,N_11396);
or U12980 (N_12980,N_11025,N_11294);
and U12981 (N_12981,N_11854,N_10676);
or U12982 (N_12982,N_9500,N_11289);
or U12983 (N_12983,N_12430,N_12318);
nand U12984 (N_12984,N_11750,N_9984);
or U12985 (N_12985,N_10569,N_10831);
and U12986 (N_12986,N_9880,N_11443);
nand U12987 (N_12987,N_10076,N_12422);
or U12988 (N_12988,N_11015,N_10508);
and U12989 (N_12989,N_10592,N_10048);
xor U12990 (N_12990,N_10930,N_11420);
and U12991 (N_12991,N_12432,N_11239);
nor U12992 (N_12992,N_12059,N_12108);
nand U12993 (N_12993,N_11884,N_10746);
or U12994 (N_12994,N_9520,N_9415);
xnor U12995 (N_12995,N_10716,N_12263);
nor U12996 (N_12996,N_10318,N_11565);
nand U12997 (N_12997,N_11908,N_11276);
or U12998 (N_12998,N_9455,N_12391);
and U12999 (N_12999,N_12198,N_10991);
or U13000 (N_13000,N_11607,N_11919);
xnor U13001 (N_13001,N_10390,N_10584);
or U13002 (N_13002,N_10192,N_9724);
nand U13003 (N_13003,N_10493,N_11014);
nor U13004 (N_13004,N_10292,N_9881);
or U13005 (N_13005,N_9819,N_10583);
nand U13006 (N_13006,N_12228,N_10538);
or U13007 (N_13007,N_10707,N_11767);
nor U13008 (N_13008,N_9856,N_11533);
or U13009 (N_13009,N_12395,N_11754);
xor U13010 (N_13010,N_12097,N_10429);
nor U13011 (N_13011,N_10684,N_11426);
or U13012 (N_13012,N_10674,N_11129);
nor U13013 (N_13013,N_11877,N_12226);
and U13014 (N_13014,N_9715,N_9772);
and U13015 (N_13015,N_11654,N_10641);
nand U13016 (N_13016,N_10543,N_11863);
xor U13017 (N_13017,N_12144,N_11622);
or U13018 (N_13018,N_11853,N_12045);
or U13019 (N_13019,N_11267,N_12499);
nor U13020 (N_13020,N_10409,N_10381);
nor U13021 (N_13021,N_12180,N_10072);
nand U13022 (N_13022,N_10327,N_10152);
or U13023 (N_13023,N_9485,N_12123);
or U13024 (N_13024,N_11958,N_12085);
and U13025 (N_13025,N_10805,N_10554);
xnor U13026 (N_13026,N_11953,N_9901);
or U13027 (N_13027,N_11188,N_12290);
nor U13028 (N_13028,N_12037,N_11690);
xor U13029 (N_13029,N_10051,N_9631);
nand U13030 (N_13030,N_12121,N_9601);
or U13031 (N_13031,N_10772,N_10541);
nor U13032 (N_13032,N_10456,N_12288);
nand U13033 (N_13033,N_9571,N_12367);
or U13034 (N_13034,N_10481,N_12105);
nor U13035 (N_13035,N_11130,N_9734);
nor U13036 (N_13036,N_11742,N_11207);
nand U13037 (N_13037,N_10809,N_11820);
or U13038 (N_13038,N_12244,N_9832);
nor U13039 (N_13039,N_9759,N_9860);
nor U13040 (N_13040,N_9385,N_9666);
and U13041 (N_13041,N_12053,N_11297);
nand U13042 (N_13042,N_12107,N_12452);
or U13043 (N_13043,N_9393,N_10473);
xor U13044 (N_13044,N_9674,N_9720);
nor U13045 (N_13045,N_12148,N_12393);
nand U13046 (N_13046,N_12484,N_11995);
nand U13047 (N_13047,N_11676,N_11669);
nand U13048 (N_13048,N_11584,N_10566);
xor U13049 (N_13049,N_9704,N_10917);
or U13050 (N_13050,N_9835,N_10821);
nor U13051 (N_13051,N_10021,N_11928);
xor U13052 (N_13052,N_11579,N_12309);
or U13053 (N_13053,N_10425,N_11427);
nand U13054 (N_13054,N_10778,N_9506);
and U13055 (N_13055,N_11603,N_11377);
xor U13056 (N_13056,N_11281,N_11998);
nor U13057 (N_13057,N_10141,N_11647);
and U13058 (N_13058,N_12066,N_10946);
nand U13059 (N_13059,N_10168,N_11240);
or U13060 (N_13060,N_11834,N_10023);
nor U13061 (N_13061,N_11381,N_11151);
nor U13062 (N_13062,N_11097,N_10307);
nor U13063 (N_13063,N_10054,N_11529);
or U13064 (N_13064,N_10372,N_11282);
or U13065 (N_13065,N_12280,N_11000);
nand U13066 (N_13066,N_9853,N_9636);
nor U13067 (N_13067,N_11587,N_10705);
nor U13068 (N_13068,N_10096,N_12373);
xor U13069 (N_13069,N_9510,N_10014);
and U13070 (N_13070,N_10217,N_10008);
nand U13071 (N_13071,N_11482,N_11638);
nor U13072 (N_13072,N_10196,N_11618);
xnor U13073 (N_13073,N_9755,N_10865);
nor U13074 (N_13074,N_9687,N_11848);
nand U13075 (N_13075,N_11572,N_11413);
nor U13076 (N_13076,N_10625,N_9527);
or U13077 (N_13077,N_9613,N_12139);
nand U13078 (N_13078,N_10199,N_12048);
nand U13079 (N_13079,N_11406,N_10709);
or U13080 (N_13080,N_11100,N_10829);
xor U13081 (N_13081,N_11665,N_10335);
or U13082 (N_13082,N_9710,N_11304);
nor U13083 (N_13083,N_12489,N_10321);
or U13084 (N_13084,N_9522,N_11568);
nand U13085 (N_13085,N_11382,N_11544);
nand U13086 (N_13086,N_12281,N_11329);
nand U13087 (N_13087,N_10536,N_10404);
nand U13088 (N_13088,N_10648,N_12316);
and U13089 (N_13089,N_10075,N_10088);
nor U13090 (N_13090,N_9451,N_9445);
and U13091 (N_13091,N_10696,N_12114);
or U13092 (N_13092,N_10621,N_10731);
or U13093 (N_13093,N_10638,N_11932);
nand U13094 (N_13094,N_10653,N_10158);
xnor U13095 (N_13095,N_9616,N_11979);
and U13096 (N_13096,N_12491,N_10998);
or U13097 (N_13097,N_10099,N_9554);
nand U13098 (N_13098,N_11298,N_9726);
nor U13099 (N_13099,N_9757,N_11736);
or U13100 (N_13100,N_11143,N_9627);
nor U13101 (N_13101,N_12201,N_11955);
or U13102 (N_13102,N_10420,N_9963);
nor U13103 (N_13103,N_10899,N_10748);
and U13104 (N_13104,N_10688,N_11317);
nand U13105 (N_13105,N_10668,N_9625);
nand U13106 (N_13106,N_10760,N_9573);
or U13107 (N_13107,N_10005,N_11909);
nand U13108 (N_13108,N_10725,N_11232);
nor U13109 (N_13109,N_9993,N_10597);
nor U13110 (N_13110,N_10442,N_9994);
nor U13111 (N_13111,N_10344,N_11139);
nand U13112 (N_13112,N_9683,N_10259);
nand U13113 (N_13113,N_9910,N_11936);
nor U13114 (N_13114,N_11756,N_10387);
or U13115 (N_13115,N_9660,N_11013);
and U13116 (N_13116,N_9493,N_9882);
nor U13117 (N_13117,N_11064,N_11039);
nand U13118 (N_13118,N_11896,N_11318);
and U13119 (N_13119,N_11776,N_12454);
and U13120 (N_13120,N_10091,N_10022);
or U13121 (N_13121,N_12301,N_11866);
nor U13122 (N_13122,N_9790,N_10107);
and U13123 (N_13123,N_10116,N_12341);
and U13124 (N_13124,N_9492,N_10043);
and U13125 (N_13125,N_10639,N_11734);
and U13126 (N_13126,N_11055,N_9954);
and U13127 (N_13127,N_10455,N_10884);
xnor U13128 (N_13128,N_10689,N_12276);
and U13129 (N_13129,N_10878,N_11745);
or U13130 (N_13130,N_11394,N_10774);
or U13131 (N_13131,N_11459,N_9751);
nand U13132 (N_13132,N_11547,N_10931);
nand U13133 (N_13133,N_9967,N_12337);
nor U13134 (N_13134,N_10995,N_11590);
or U13135 (N_13135,N_10916,N_12348);
xor U13136 (N_13136,N_10329,N_10908);
xor U13137 (N_13137,N_12433,N_9782);
or U13138 (N_13138,N_10925,N_10159);
nor U13139 (N_13139,N_9700,N_10749);
nand U13140 (N_13140,N_9540,N_11888);
and U13141 (N_13141,N_10580,N_10209);
nand U13142 (N_13142,N_10564,N_10888);
and U13143 (N_13143,N_10823,N_9603);
or U13144 (N_13144,N_11912,N_10124);
nor U13145 (N_13145,N_12331,N_10743);
nand U13146 (N_13146,N_10655,N_10506);
xor U13147 (N_13147,N_12234,N_11408);
or U13148 (N_13148,N_9427,N_10979);
or U13149 (N_13149,N_12264,N_10007);
nor U13150 (N_13150,N_11041,N_11278);
and U13151 (N_13151,N_9671,N_12171);
and U13152 (N_13152,N_10900,N_10118);
and U13153 (N_13153,N_10405,N_10120);
nand U13154 (N_13154,N_9754,N_10366);
nor U13155 (N_13155,N_12272,N_10303);
xor U13156 (N_13156,N_10368,N_10693);
nor U13157 (N_13157,N_11046,N_12140);
xnor U13158 (N_13158,N_11434,N_10953);
nand U13159 (N_13159,N_11089,N_11949);
nor U13160 (N_13160,N_10711,N_10128);
and U13161 (N_13161,N_12099,N_11989);
or U13162 (N_13162,N_9637,N_10847);
nor U13163 (N_13163,N_11040,N_10095);
nand U13164 (N_13164,N_10866,N_11273);
and U13165 (N_13165,N_12294,N_12149);
nand U13166 (N_13166,N_11174,N_12000);
nor U13167 (N_13167,N_11962,N_10901);
nor U13168 (N_13168,N_10458,N_9541);
xnor U13169 (N_13169,N_11384,N_11358);
and U13170 (N_13170,N_10483,N_11270);
nor U13171 (N_13171,N_10736,N_11878);
xnor U13172 (N_13172,N_9825,N_10463);
and U13173 (N_13173,N_10790,N_11066);
nor U13174 (N_13174,N_10755,N_12120);
nand U13175 (N_13175,N_9930,N_9926);
or U13176 (N_13176,N_9761,N_11447);
nand U13177 (N_13177,N_9950,N_10822);
and U13178 (N_13178,N_9595,N_10242);
and U13179 (N_13179,N_9619,N_10083);
xnor U13180 (N_13180,N_11343,N_11846);
and U13181 (N_13181,N_9640,N_12359);
or U13182 (N_13182,N_10382,N_11362);
xor U13183 (N_13183,N_10795,N_9925);
and U13184 (N_13184,N_11076,N_11492);
nand U13185 (N_13185,N_10521,N_11003);
and U13186 (N_13186,N_10608,N_11070);
nor U13187 (N_13187,N_11016,N_9388);
nand U13188 (N_13188,N_11682,N_10837);
or U13189 (N_13189,N_11865,N_12033);
xor U13190 (N_13190,N_11722,N_11428);
nand U13191 (N_13191,N_10518,N_11285);
and U13192 (N_13192,N_11218,N_9651);
and U13193 (N_13193,N_12282,N_10100);
nor U13194 (N_13194,N_10950,N_10264);
nand U13195 (N_13195,N_11299,N_10238);
and U13196 (N_13196,N_10732,N_11807);
or U13197 (N_13197,N_10426,N_11051);
nor U13198 (N_13198,N_11788,N_12345);
nand U13199 (N_13199,N_11553,N_9423);
or U13200 (N_13200,N_12392,N_10839);
nand U13201 (N_13201,N_11509,N_9591);
xor U13202 (N_13202,N_10703,N_9945);
nor U13203 (N_13203,N_12334,N_11630);
or U13204 (N_13204,N_10403,N_11030);
nand U13205 (N_13205,N_10815,N_11088);
nor U13206 (N_13206,N_10170,N_12371);
nand U13207 (N_13207,N_11583,N_11774);
nor U13208 (N_13208,N_9587,N_12147);
nor U13209 (N_13209,N_11887,N_11766);
or U13210 (N_13210,N_9665,N_11659);
and U13211 (N_13211,N_10640,N_10747);
nor U13212 (N_13212,N_11162,N_11350);
nand U13213 (N_13213,N_10838,N_10254);
or U13214 (N_13214,N_9454,N_12425);
or U13215 (N_13215,N_9948,N_9565);
and U13216 (N_13216,N_11719,N_9719);
and U13217 (N_13217,N_11550,N_9420);
or U13218 (N_13218,N_11950,N_9943);
nor U13219 (N_13219,N_9379,N_11485);
nand U13220 (N_13220,N_11319,N_10109);
nand U13221 (N_13221,N_12022,N_10441);
nand U13222 (N_13222,N_10204,N_10710);
xor U13223 (N_13223,N_12172,N_10962);
or U13224 (N_13224,N_11165,N_12034);
xor U13225 (N_13225,N_9895,N_10570);
xor U13226 (N_13226,N_9914,N_9843);
and U13227 (N_13227,N_11641,N_12296);
and U13228 (N_13228,N_11836,N_11765);
nor U13229 (N_13229,N_10246,N_10233);
nand U13230 (N_13230,N_10467,N_9662);
nor U13231 (N_13231,N_9558,N_10862);
nor U13232 (N_13232,N_11245,N_11198);
and U13233 (N_13233,N_9814,N_9956);
nor U13234 (N_13234,N_9934,N_10783);
xor U13235 (N_13235,N_12241,N_9376);
nand U13236 (N_13236,N_11045,N_10391);
or U13237 (N_13237,N_9999,N_11558);
and U13238 (N_13238,N_11368,N_12078);
and U13239 (N_13239,N_10036,N_10734);
nor U13240 (N_13240,N_11592,N_10231);
and U13241 (N_13241,N_11246,N_10679);
and U13242 (N_13242,N_10316,N_11952);
nor U13243 (N_13243,N_12132,N_11803);
or U13244 (N_13244,N_12094,N_12404);
or U13245 (N_13245,N_9564,N_9419);
nor U13246 (N_13246,N_10827,N_10659);
nand U13247 (N_13247,N_11935,N_11823);
nand U13248 (N_13248,N_10332,N_9529);
and U13249 (N_13249,N_10389,N_10762);
nor U13250 (N_13250,N_11092,N_10891);
and U13251 (N_13251,N_11115,N_10796);
or U13252 (N_13252,N_11505,N_10586);
and U13253 (N_13253,N_10379,N_12008);
or U13254 (N_13254,N_12328,N_10067);
nor U13255 (N_13255,N_10698,N_12420);
and U13256 (N_13256,N_9938,N_9383);
or U13257 (N_13257,N_11999,N_10430);
or U13258 (N_13258,N_11449,N_11169);
nand U13259 (N_13259,N_10959,N_9547);
or U13260 (N_13260,N_11555,N_11627);
or U13261 (N_13261,N_10682,N_10395);
nor U13262 (N_13262,N_9652,N_10119);
xor U13263 (N_13263,N_11063,N_12052);
and U13264 (N_13264,N_9692,N_10830);
and U13265 (N_13265,N_12095,N_10985);
nor U13266 (N_13266,N_11483,N_10000);
and U13267 (N_13267,N_11094,N_11372);
and U13268 (N_13268,N_11334,N_9728);
nor U13269 (N_13269,N_10334,N_9760);
nor U13270 (N_13270,N_9523,N_12219);
and U13271 (N_13271,N_10907,N_9990);
or U13272 (N_13272,N_11132,N_9917);
nand U13273 (N_13273,N_10457,N_9875);
nor U13274 (N_13274,N_10978,N_9789);
and U13275 (N_13275,N_11404,N_11811);
nand U13276 (N_13276,N_12246,N_11390);
nor U13277 (N_13277,N_10482,N_12352);
nor U13278 (N_13278,N_10859,N_11241);
nand U13279 (N_13279,N_11930,N_12071);
or U13280 (N_13280,N_9380,N_10111);
and U13281 (N_13281,N_10910,N_9624);
nor U13282 (N_13282,N_10500,N_10872);
nor U13283 (N_13283,N_10960,N_10138);
and U13284 (N_13284,N_11438,N_11557);
or U13285 (N_13285,N_10094,N_12047);
nand U13286 (N_13286,N_10121,N_11356);
nand U13287 (N_13287,N_11359,N_9937);
xor U13288 (N_13288,N_9752,N_10477);
and U13289 (N_13289,N_11309,N_12262);
xor U13290 (N_13290,N_9940,N_10423);
nand U13291 (N_13291,N_10046,N_11858);
and U13292 (N_13292,N_11346,N_11407);
and U13293 (N_13293,N_10612,N_11598);
xnor U13294 (N_13294,N_11354,N_9446);
or U13295 (N_13295,N_10810,N_11730);
nand U13296 (N_13296,N_9508,N_12466);
xnor U13297 (N_13297,N_10386,N_11490);
nand U13298 (N_13298,N_9868,N_11511);
nor U13299 (N_13299,N_9746,N_11154);
or U13300 (N_13300,N_9659,N_11007);
or U13301 (N_13301,N_11217,N_10353);
and U13302 (N_13302,N_10343,N_12233);
and U13303 (N_13303,N_11513,N_12308);
nand U13304 (N_13304,N_11762,N_12068);
nand U13305 (N_13305,N_10171,N_10486);
xor U13306 (N_13306,N_12003,N_10471);
and U13307 (N_13307,N_11871,N_10082);
nor U13308 (N_13308,N_9516,N_11159);
nor U13309 (N_13309,N_11272,N_9801);
or U13310 (N_13310,N_9708,N_11186);
or U13311 (N_13311,N_9822,N_11491);
nand U13312 (N_13312,N_10735,N_11914);
xnor U13313 (N_13313,N_9788,N_9677);
nand U13314 (N_13314,N_11933,N_11537);
nor U13315 (N_13315,N_9560,N_12163);
and U13316 (N_13316,N_11963,N_10879);
and U13317 (N_13317,N_11148,N_10727);
and U13318 (N_13318,N_11576,N_9946);
nor U13319 (N_13319,N_10073,N_11233);
nand U13320 (N_13320,N_11512,N_12365);
and U13321 (N_13321,N_10400,N_11522);
or U13322 (N_13322,N_9764,N_9885);
nand U13323 (N_13323,N_11600,N_9823);
or U13324 (N_13324,N_12342,N_11158);
nor U13325 (N_13325,N_11886,N_10591);
or U13326 (N_13326,N_9382,N_10025);
nor U13327 (N_13327,N_12196,N_12490);
nand U13328 (N_13328,N_12494,N_12206);
or U13329 (N_13329,N_10104,N_9756);
nor U13330 (N_13330,N_9900,N_10599);
or U13331 (N_13331,N_9633,N_10961);
xor U13332 (N_13332,N_11806,N_10454);
or U13333 (N_13333,N_12231,N_11552);
xnor U13334 (N_13334,N_11580,N_11323);
nor U13335 (N_13335,N_11400,N_10894);
nand U13336 (N_13336,N_10378,N_10226);
nor U13337 (N_13337,N_10045,N_9891);
or U13338 (N_13338,N_10912,N_9852);
and U13339 (N_13339,N_12070,N_10319);
nand U13340 (N_13340,N_11134,N_10515);
and U13341 (N_13341,N_10224,N_10496);
or U13342 (N_13342,N_12064,N_9955);
nor U13343 (N_13343,N_9970,N_10275);
xnor U13344 (N_13344,N_12324,N_11540);
nand U13345 (N_13345,N_10011,N_9972);
or U13346 (N_13346,N_12356,N_11032);
and U13347 (N_13347,N_9568,N_10841);
xor U13348 (N_13348,N_11419,N_12193);
and U13349 (N_13349,N_11495,N_12039);
or U13350 (N_13350,N_9632,N_12162);
nor U13351 (N_13351,N_10377,N_11432);
nand U13352 (N_13352,N_12175,N_10606);
and U13353 (N_13353,N_12013,N_11095);
nor U13354 (N_13354,N_12372,N_11925);
nand U13355 (N_13355,N_11680,N_9725);
nand U13356 (N_13356,N_9590,N_9486);
xor U13357 (N_13357,N_10610,N_10132);
nand U13358 (N_13358,N_11517,N_10855);
nand U13359 (N_13359,N_11405,N_10882);
and U13360 (N_13360,N_9538,N_9831);
xor U13361 (N_13361,N_10184,N_11195);
and U13362 (N_13362,N_11686,N_10028);
nor U13363 (N_13363,N_10215,N_10895);
or U13364 (N_13364,N_12358,N_10664);
and U13365 (N_13365,N_10750,N_11857);
or U13366 (N_13366,N_11118,N_11918);
nand U13367 (N_13367,N_11316,N_11538);
or U13368 (N_13368,N_9969,N_11149);
nand U13369 (N_13369,N_9504,N_10758);
nand U13370 (N_13370,N_9695,N_10298);
nand U13371 (N_13371,N_11385,N_10180);
nand U13372 (N_13372,N_12421,N_11290);
and U13373 (N_13373,N_11818,N_10399);
nand U13374 (N_13374,N_10240,N_10814);
nor U13375 (N_13375,N_12245,N_10252);
xnor U13376 (N_13376,N_10965,N_11595);
and U13377 (N_13377,N_10977,N_10098);
or U13378 (N_13378,N_12232,N_12464);
nor U13379 (N_13379,N_11376,N_11586);
and U13380 (N_13380,N_11688,N_10663);
or U13381 (N_13381,N_11920,N_12435);
nor U13382 (N_13382,N_11306,N_9672);
and U13383 (N_13383,N_11571,N_11389);
and U13384 (N_13384,N_10927,N_11843);
xor U13385 (N_13385,N_9795,N_10635);
nor U13386 (N_13386,N_11727,N_11697);
xnor U13387 (N_13387,N_12181,N_12143);
and U13388 (N_13388,N_9899,N_10858);
or U13389 (N_13389,N_12153,N_9723);
nor U13390 (N_13390,N_9667,N_9482);
or U13391 (N_13391,N_11341,N_11019);
nand U13392 (N_13392,N_11718,N_10545);
nor U13393 (N_13393,N_11057,N_10437);
nand U13394 (N_13394,N_9753,N_11330);
nand U13395 (N_13395,N_10291,N_9552);
nor U13396 (N_13396,N_9959,N_9549);
nor U13397 (N_13397,N_11514,N_10844);
and U13398 (N_13398,N_12221,N_9491);
xor U13399 (N_13399,N_11182,N_11985);
or U13400 (N_13400,N_12230,N_12208);
and U13401 (N_13401,N_10987,N_9889);
and U13402 (N_13402,N_11477,N_11749);
or U13403 (N_13403,N_11814,N_12203);
nor U13404 (N_13404,N_10826,N_10364);
nor U13405 (N_13405,N_12128,N_10237);
nand U13406 (N_13406,N_9919,N_10278);
nand U13407 (N_13407,N_11621,N_10773);
or U13408 (N_13408,N_11726,N_11035);
xnor U13409 (N_13409,N_11657,N_11219);
nand U13410 (N_13410,N_9436,N_11990);
nand U13411 (N_13411,N_12402,N_11433);
nand U13412 (N_13412,N_12015,N_11141);
nand U13413 (N_13413,N_9961,N_12251);
nand U13414 (N_13414,N_10037,N_10016);
nor U13415 (N_13415,N_9866,N_10013);
nand U13416 (N_13416,N_11348,N_9957);
or U13417 (N_13417,N_11494,N_9920);
nor U13418 (N_13418,N_11249,N_9874);
or U13419 (N_13419,N_10032,N_12138);
and U13420 (N_13420,N_11131,N_11116);
or U13421 (N_13421,N_10296,N_11714);
nor U13422 (N_13422,N_11923,N_11966);
or U13423 (N_13423,N_10489,N_9629);
xnor U13424 (N_13424,N_11301,N_11256);
and U13425 (N_13425,N_10886,N_11773);
and U13426 (N_13426,N_11200,N_11484);
nand U13427 (N_13427,N_12471,N_9614);
nand U13428 (N_13428,N_10622,N_10517);
or U13429 (N_13429,N_11326,N_10863);
xnor U13430 (N_13430,N_10913,N_12157);
xor U13431 (N_13431,N_11817,N_11608);
and U13432 (N_13432,N_12043,N_11086);
or U13433 (N_13433,N_9578,N_10523);
xor U13434 (N_13434,N_9509,N_11694);
or U13435 (N_13435,N_10786,N_11125);
or U13436 (N_13436,N_10937,N_11336);
xor U13437 (N_13437,N_10572,N_12223);
or U13438 (N_13438,N_9730,N_11173);
xor U13439 (N_13439,N_10465,N_10903);
and U13440 (N_13440,N_10421,N_11981);
nor U13441 (N_13441,N_11472,N_11268);
xor U13442 (N_13442,N_10654,N_11601);
xor U13443 (N_13443,N_10941,N_12006);
nor U13444 (N_13444,N_12440,N_10114);
or U13445 (N_13445,N_9811,N_11678);
nand U13446 (N_13446,N_9604,N_9426);
and U13447 (N_13447,N_12268,N_11103);
xnor U13448 (N_13448,N_9557,N_12384);
nor U13449 (N_13449,N_12382,N_12215);
nand U13450 (N_13450,N_11054,N_11313);
nand U13451 (N_13451,N_12403,N_11366);
and U13452 (N_13452,N_12247,N_12023);
or U13453 (N_13453,N_11111,N_11280);
nand U13454 (N_13454,N_10185,N_10733);
nor U13455 (N_13455,N_11760,N_11642);
nand U13456 (N_13456,N_12025,N_12202);
xnor U13457 (N_13457,N_10560,N_10902);
or U13458 (N_13458,N_10360,N_9849);
or U13459 (N_13459,N_12285,N_10911);
or U13460 (N_13460,N_11876,N_11327);
nor U13461 (N_13461,N_11204,N_11994);
nor U13462 (N_13462,N_9449,N_11554);
or U13463 (N_13463,N_9717,N_10153);
nand U13464 (N_13464,N_10980,N_11596);
nor U13465 (N_13465,N_9429,N_12423);
or U13466 (N_13466,N_11373,N_10490);
nor U13467 (N_13467,N_12179,N_9813);
and U13468 (N_13468,N_10058,N_10287);
nor U13469 (N_13469,N_11813,N_12369);
nand U13470 (N_13470,N_12270,N_10195);
nor U13471 (N_13471,N_10149,N_11370);
and U13472 (N_13472,N_9643,N_11614);
and U13473 (N_13473,N_9775,N_11992);
nand U13474 (N_13474,N_9922,N_11190);
nor U13475 (N_13475,N_11191,N_12005);
or U13476 (N_13476,N_9830,N_12125);
xnor U13477 (N_13477,N_10848,N_10867);
or U13478 (N_13478,N_11457,N_10160);
nand U13479 (N_13479,N_12170,N_9397);
xnor U13480 (N_13480,N_9553,N_12414);
nor U13481 (N_13481,N_11692,N_10939);
and U13482 (N_13482,N_9577,N_10777);
or U13483 (N_13483,N_9995,N_10472);
nor U13484 (N_13484,N_12298,N_11242);
or U13485 (N_13485,N_10181,N_10765);
and U13486 (N_13486,N_11465,N_10163);
and U13487 (N_13487,N_11941,N_9477);
xor U13488 (N_13488,N_10741,N_11506);
xnor U13489 (N_13489,N_12339,N_11801);
nor U13490 (N_13490,N_11193,N_11701);
or U13491 (N_13491,N_11833,N_10384);
and U13492 (N_13492,N_11588,N_10595);
and U13493 (N_13493,N_10436,N_11852);
or U13494 (N_13494,N_10010,N_12357);
or U13495 (N_13495,N_9580,N_10784);
nand U13496 (N_13496,N_11947,N_12130);
nor U13497 (N_13497,N_9837,N_12277);
nand U13498 (N_13498,N_10645,N_10433);
xnor U13499 (N_13499,N_10616,N_12237);
or U13500 (N_13500,N_10745,N_10418);
xnor U13501 (N_13501,N_10041,N_12199);
nand U13502 (N_13502,N_9439,N_11940);
or U13503 (N_13503,N_11442,N_9550);
and U13504 (N_13504,N_11723,N_12054);
nand U13505 (N_13505,N_10719,N_10700);
xnor U13506 (N_13506,N_12049,N_10042);
and U13507 (N_13507,N_9808,N_12214);
or U13508 (N_13508,N_11716,N_12191);
and U13509 (N_13509,N_12355,N_11713);
and U13510 (N_13510,N_10177,N_12115);
nand U13511 (N_13511,N_10926,N_12346);
nor U13512 (N_13512,N_10239,N_11410);
nand U13513 (N_13513,N_11702,N_10144);
nand U13514 (N_13514,N_10781,N_9855);
and U13515 (N_13515,N_11126,N_9768);
nand U13516 (N_13516,N_9556,N_12478);
nand U13517 (N_13517,N_11880,N_10297);
nand U13518 (N_13518,N_12106,N_10415);
nor U13519 (N_13519,N_11977,N_11470);
xor U13520 (N_13520,N_11542,N_10068);
nand U13521 (N_13521,N_9475,N_12031);
nor U13522 (N_13522,N_9441,N_11922);
or U13523 (N_13523,N_12488,N_10651);
or U13524 (N_13524,N_12480,N_11921);
nand U13525 (N_13525,N_11202,N_11471);
or U13526 (N_13526,N_10680,N_9607);
or U13527 (N_13527,N_11144,N_12194);
nand U13528 (N_13528,N_11560,N_10681);
nor U13529 (N_13529,N_9977,N_11951);
or U13530 (N_13530,N_10799,N_11778);
nor U13531 (N_13531,N_10955,N_12455);
and U13532 (N_13532,N_9653,N_12340);
nand U13533 (N_13533,N_10281,N_11679);
and U13534 (N_13534,N_11573,N_12325);
and U13535 (N_13535,N_11074,N_12165);
or U13536 (N_13536,N_10988,N_9952);
nor U13537 (N_13537,N_9893,N_12238);
nand U13538 (N_13538,N_9731,N_10172);
and U13539 (N_13539,N_9461,N_10997);
xor U13540 (N_13540,N_10675,N_10849);
nand U13541 (N_13541,N_11725,N_12474);
or U13542 (N_13542,N_10782,N_10102);
nor U13543 (N_13543,N_12122,N_10355);
and U13544 (N_13544,N_10775,N_10924);
xor U13545 (N_13545,N_10017,N_9675);
nand U13546 (N_13546,N_9682,N_12496);
nand U13547 (N_13547,N_11815,N_10285);
nor U13548 (N_13548,N_9815,N_9805);
nand U13549 (N_13549,N_10053,N_12336);
or U13550 (N_13550,N_10309,N_9912);
nand U13551 (N_13551,N_9593,N_9684);
nand U13552 (N_13552,N_10066,N_9435);
nor U13553 (N_13553,N_11314,N_11724);
nor U13554 (N_13554,N_11879,N_10272);
nor U13555 (N_13555,N_11274,N_11112);
and U13556 (N_13556,N_10601,N_12429);
xor U13557 (N_13557,N_11456,N_10708);
nor U13558 (N_13558,N_11418,N_9496);
nand U13559 (N_13559,N_9465,N_10139);
and U13560 (N_13560,N_9740,N_10216);
or U13561 (N_13561,N_11504,N_9396);
or U13562 (N_13562,N_11976,N_11166);
and U13563 (N_13563,N_10660,N_12259);
nor U13564 (N_13564,N_10857,N_11421);
or U13565 (N_13565,N_12079,N_10250);
xor U13566 (N_13566,N_10989,N_10194);
nand U13567 (N_13567,N_11004,N_12127);
and U13568 (N_13568,N_12004,N_9869);
nor U13569 (N_13569,N_11673,N_10889);
and U13570 (N_13570,N_11757,N_9696);
or U13571 (N_13571,N_12050,N_11360);
or U13572 (N_13572,N_11578,N_11439);
and U13573 (N_13573,N_11628,N_9375);
and U13574 (N_13574,N_9612,N_10834);
nor U13575 (N_13575,N_11048,N_10738);
or U13576 (N_13576,N_11859,N_10791);
and U13577 (N_13577,N_10528,N_9817);
and U13578 (N_13578,N_10922,N_10059);
or U13579 (N_13579,N_9905,N_11768);
and U13580 (N_13580,N_9448,N_12098);
and U13581 (N_13581,N_11228,N_12188);
nand U13582 (N_13582,N_10190,N_11875);
nand U13583 (N_13583,N_11371,N_9807);
nand U13584 (N_13584,N_11468,N_12253);
nand U13585 (N_13585,N_10413,N_10945);
and U13586 (N_13586,N_11728,N_10906);
nor U13587 (N_13587,N_11164,N_9689);
nor U13588 (N_13588,N_10112,N_10056);
nor U13589 (N_13589,N_10933,N_11658);
and U13590 (N_13590,N_11147,N_10555);
nand U13591 (N_13591,N_11970,N_9924);
nand U13592 (N_13592,N_12056,N_10375);
xnor U13593 (N_13593,N_10146,N_9661);
xnor U13594 (N_13594,N_11783,N_10009);
or U13595 (N_13595,N_9635,N_10392);
or U13596 (N_13596,N_12479,N_12222);
and U13597 (N_13597,N_9909,N_9806);
and U13598 (N_13598,N_9915,N_10923);
nor U13599 (N_13599,N_10308,N_9862);
xor U13600 (N_13600,N_9515,N_12344);
nand U13601 (N_13601,N_11402,N_10428);
nand U13602 (N_13602,N_9430,N_9404);
or U13603 (N_13603,N_12434,N_11810);
xnor U13604 (N_13604,N_10117,N_11548);
nand U13605 (N_13605,N_11698,N_10764);
or U13606 (N_13606,N_12426,N_11113);
or U13607 (N_13607,N_10984,N_11028);
and U13608 (N_13608,N_9965,N_11636);
or U13609 (N_13609,N_12329,N_10393);
nand U13610 (N_13610,N_12058,N_11080);
or U13611 (N_13611,N_11342,N_11061);
nor U13612 (N_13612,N_12449,N_12427);
or U13613 (N_13613,N_9484,N_9828);
and U13614 (N_13614,N_9663,N_11687);
nor U13615 (N_13615,N_9778,N_9974);
nand U13616 (N_13616,N_11078,N_11987);
nand U13617 (N_13617,N_11515,N_12184);
nand U13618 (N_13618,N_12497,N_11589);
nand U13619 (N_13619,N_12398,N_10614);
or U13620 (N_13620,N_11689,N_11312);
or U13621 (N_13621,N_10410,N_12300);
nor U13622 (N_13622,N_11777,N_10176);
or U13623 (N_13623,N_11794,N_9400);
nand U13624 (N_13624,N_9733,N_10898);
nor U13625 (N_13625,N_10756,N_9907);
nand U13626 (N_13626,N_11349,N_12333);
nand U13627 (N_13627,N_9976,N_10603);
and U13628 (N_13628,N_11770,N_10106);
nor U13629 (N_13629,N_11010,N_9861);
or U13630 (N_13630,N_11458,N_9576);
nand U13631 (N_13631,N_11615,N_10921);
or U13632 (N_13632,N_10324,N_10103);
nor U13633 (N_13633,N_10057,N_9964);
and U13634 (N_13634,N_11911,N_11177);
or U13635 (N_13635,N_10940,N_10754);
xnor U13636 (N_13636,N_12019,N_10348);
and U13637 (N_13637,N_9453,N_12405);
and U13638 (N_13638,N_10207,N_12104);
and U13639 (N_13639,N_10797,N_9473);
nand U13640 (N_13640,N_10631,N_11043);
or U13641 (N_13641,N_9777,N_12410);
nor U13642 (N_13642,N_9953,N_10915);
nand U13643 (N_13643,N_9973,N_12077);
nand U13644 (N_13644,N_11235,N_10806);
and U13645 (N_13645,N_10963,N_11257);
nor U13646 (N_13646,N_12020,N_11534);
or U13647 (N_13647,N_10035,N_11067);
xor U13648 (N_13648,N_10996,N_10363);
or U13649 (N_13649,N_11226,N_10453);
or U13650 (N_13650,N_11828,N_12211);
and U13651 (N_13651,N_9450,N_9495);
xnor U13652 (N_13652,N_10753,N_9600);
nor U13653 (N_13653,N_11991,N_10370);
nand U13654 (N_13654,N_10438,N_12477);
nand U13655 (N_13655,N_9499,N_9918);
and U13656 (N_13656,N_10726,N_12260);
nand U13657 (N_13657,N_10785,N_9384);
nor U13658 (N_13658,N_9422,N_9854);
or U13659 (N_13659,N_11786,N_11784);
and U13660 (N_13660,N_10819,N_10274);
nor U13661 (N_13661,N_11227,N_12279);
or U13662 (N_13662,N_10229,N_10330);
or U13663 (N_13663,N_11179,N_12444);
nor U13664 (N_13664,N_11082,N_11436);
nand U13665 (N_13665,N_10667,N_10113);
nor U13666 (N_13666,N_11140,N_10339);
and U13667 (N_13667,N_12376,N_12212);
or U13668 (N_13668,N_9721,N_9766);
nand U13669 (N_13669,N_9501,N_11808);
xnor U13670 (N_13670,N_9691,N_11277);
nor U13671 (N_13671,N_10532,N_9693);
and U13672 (N_13672,N_9608,N_10840);
xor U13673 (N_13673,N_10193,N_9803);
and U13674 (N_13674,N_9546,N_10577);
or U13675 (N_13675,N_11378,N_11303);
nand U13676 (N_13676,N_10093,N_11838);
or U13677 (N_13677,N_11073,N_11422);
nor U13678 (N_13678,N_11740,N_11626);
nand U13679 (N_13679,N_11629,N_9394);
nor U13680 (N_13680,N_11812,N_9474);
nand U13681 (N_13681,N_9551,N_9567);
nor U13682 (N_13682,N_10262,N_11163);
nand U13683 (N_13683,N_10854,N_12274);
nor U13684 (N_13684,N_9709,N_12386);
and U13685 (N_13685,N_10832,N_11029);
nand U13686 (N_13686,N_9810,N_10480);
and U13687 (N_13687,N_11729,N_10282);
xor U13688 (N_13688,N_9744,N_10265);
or U13689 (N_13689,N_12024,N_10565);
and U13690 (N_13690,N_11655,N_12126);
or U13691 (N_13691,N_9389,N_11835);
and U13692 (N_13692,N_9735,N_10526);
or U13693 (N_13693,N_11212,N_10520);
nand U13694 (N_13694,N_11816,N_11455);
nor U13695 (N_13695,N_11429,N_9821);
nor U13696 (N_13696,N_9411,N_11797);
nand U13697 (N_13697,N_10218,N_9596);
or U13698 (N_13698,N_10788,N_11606);
and U13699 (N_13699,N_11874,N_11855);
or U13700 (N_13700,N_10673,N_10155);
xnor U13701 (N_13701,N_10411,N_10443);
and U13702 (N_13702,N_12151,N_12302);
and U13703 (N_13703,N_9678,N_12271);
nand U13704 (N_13704,N_9421,N_11699);
nor U13705 (N_13705,N_10973,N_9585);
nor U13706 (N_13706,N_11466,N_11305);
nand U13707 (N_13707,N_10957,N_11860);
nand U13708 (N_13708,N_10767,N_9850);
or U13709 (N_13709,N_12360,N_10026);
and U13710 (N_13710,N_12257,N_12178);
and U13711 (N_13711,N_10952,N_9894);
nor U13712 (N_13712,N_10557,N_9826);
and U13713 (N_13713,N_10544,N_12187);
xor U13714 (N_13714,N_9620,N_11569);
nand U13715 (N_13715,N_10956,N_12166);
nor U13716 (N_13716,N_9440,N_9865);
nand U13717 (N_13717,N_10249,N_11231);
nor U13718 (N_13718,N_9658,N_10742);
nand U13719 (N_13719,N_11199,N_10223);
nand U13720 (N_13720,N_11444,N_10516);
nor U13721 (N_13721,N_10699,N_10123);
or U13722 (N_13722,N_11684,N_11872);
or U13723 (N_13723,N_11942,N_12437);
or U13724 (N_13724,N_10812,N_11897);
nor U13725 (N_13725,N_11799,N_9599);
nor U13726 (N_13726,N_9414,N_10562);
and U13727 (N_13727,N_11546,N_10825);
and U13728 (N_13728,N_11840,N_11594);
nor U13729 (N_13729,N_11156,N_10643);
or U13730 (N_13730,N_10450,N_10341);
xnor U13731 (N_13731,N_9525,N_10752);
nor U13732 (N_13732,N_11707,N_9488);
nor U13733 (N_13733,N_11961,N_12038);
and U13734 (N_13734,N_11666,N_12051);
nor U13735 (N_13735,N_9763,N_10687);
nand U13736 (N_13736,N_9464,N_10611);
nor U13737 (N_13737,N_10951,N_10856);
xor U13738 (N_13738,N_10003,N_12343);
and U13739 (N_13739,N_10167,N_10444);
nand U13740 (N_13740,N_10944,N_10585);
or U13741 (N_13741,N_11223,N_9758);
nor U13742 (N_13742,N_9690,N_9442);
and U13743 (N_13743,N_10875,N_11541);
xnor U13744 (N_13744,N_11258,N_9902);
and U13745 (N_13745,N_9694,N_11467);
and U13746 (N_13746,N_11804,N_9791);
xor U13747 (N_13747,N_10629,N_9796);
nor U13748 (N_13748,N_10509,N_12269);
nor U13749 (N_13749,N_11973,N_10210);
and U13750 (N_13750,N_12378,N_11881);
xnor U13751 (N_13751,N_11805,N_11192);
nor U13752 (N_13752,N_11527,N_10178);
nand U13753 (N_13753,N_10861,N_9413);
or U13754 (N_13754,N_10869,N_10312);
or U13755 (N_13755,N_10548,N_12445);
nand U13756 (N_13756,N_11269,N_12310);
and U13757 (N_13757,N_12407,N_9774);
and U13758 (N_13758,N_12074,N_11715);
and U13759 (N_13759,N_11096,N_12462);
or U13760 (N_13760,N_11624,N_9425);
and U13761 (N_13761,N_12100,N_12364);
nand U13762 (N_13762,N_12415,N_11619);
nor U13763 (N_13763,N_12267,N_10970);
nand U13764 (N_13764,N_10968,N_9767);
nor U13765 (N_13765,N_11956,N_10770);
nand U13766 (N_13766,N_10039,N_11964);
nand U13767 (N_13767,N_12317,N_11461);
nand U13768 (N_13768,N_9481,N_9839);
nor U13769 (N_13769,N_11741,N_11221);
nor U13770 (N_13770,N_9794,N_9787);
and U13771 (N_13771,N_12195,N_10510);
and U13772 (N_13772,N_12217,N_12275);
or U13773 (N_13773,N_11056,N_11910);
xnor U13774 (N_13774,N_9548,N_10876);
and U13775 (N_13775,N_12387,N_10992);
and U13776 (N_13776,N_11234,N_12323);
or U13777 (N_13777,N_11114,N_9405);
xor U13778 (N_13778,N_11145,N_11137);
and U13779 (N_13779,N_11386,N_10427);
nand U13780 (N_13780,N_9626,N_11585);
and U13781 (N_13781,N_10201,N_12009);
or U13782 (N_13782,N_10642,N_10662);
nand U13783 (N_13783,N_11364,N_10990);
nor U13784 (N_13784,N_12447,N_11523);
nor U13785 (N_13785,N_11531,N_12492);
and U13786 (N_13786,N_10813,N_9646);
and U13787 (N_13787,N_10527,N_9418);
nor U13788 (N_13788,N_11085,N_11058);
or U13789 (N_13789,N_10135,N_10092);
nand U13790 (N_13790,N_12326,N_9888);
or U13791 (N_13791,N_12353,N_10751);
nor U13792 (N_13792,N_11441,N_11695);
xor U13793 (N_13793,N_10069,N_11845);
nand U13794 (N_13794,N_11194,N_10969);
xnor U13795 (N_13795,N_10145,N_11127);
nand U13796 (N_13796,N_11561,N_9931);
nor U13797 (N_13797,N_9569,N_10818);
or U13798 (N_13798,N_10071,N_10803);
or U13799 (N_13799,N_10928,N_12486);
nand U13800 (N_13800,N_9444,N_11251);
and U13801 (N_13801,N_11625,N_10628);
and U13802 (N_13802,N_11252,N_10842);
xnor U13803 (N_13803,N_10744,N_9489);
nor U13804 (N_13804,N_9770,N_11453);
and U13805 (N_13805,N_9998,N_11819);
and U13806 (N_13806,N_11247,N_10085);
xnor U13807 (N_13807,N_9463,N_10624);
xnor U13808 (N_13808,N_10811,N_12001);
nand U13809 (N_13809,N_10478,N_11220);
nand U13810 (N_13810,N_12458,N_10620);
and U13811 (N_13811,N_10311,N_10632);
nor U13812 (N_13812,N_12424,N_9443);
and U13813 (N_13813,N_11965,N_10720);
nor U13814 (N_13814,N_10301,N_11320);
nand U13815 (N_13815,N_11753,N_10211);
and U13816 (N_13816,N_11785,N_10340);
nand U13817 (N_13817,N_10607,N_11011);
xor U13818 (N_13818,N_9408,N_10440);
and U13819 (N_13819,N_12338,N_10235);
nand U13820 (N_13820,N_10198,N_12159);
or U13821 (N_13821,N_10943,N_11653);
nor U13822 (N_13822,N_9503,N_12406);
nor U13823 (N_13823,N_10354,N_10724);
nand U13824 (N_13824,N_9407,N_10203);
or U13825 (N_13825,N_10417,N_9812);
nand U13826 (N_13826,N_11075,N_9622);
and U13827 (N_13827,N_10346,N_10934);
and U13828 (N_13828,N_10294,N_10877);
or U13829 (N_13829,N_10633,N_11677);
nand U13830 (N_13830,N_12225,N_9669);
and U13831 (N_13831,N_11044,N_10034);
or U13832 (N_13832,N_10828,N_9829);
and U13833 (N_13833,N_10006,N_11508);
xor U13834 (N_13834,N_12436,N_10302);
nor U13835 (N_13835,N_10929,N_10131);
nor U13836 (N_13836,N_11262,N_11563);
nand U13837 (N_13837,N_11475,N_10623);
xor U13838 (N_13838,N_9840,N_12213);
and U13839 (N_13839,N_9864,N_9979);
nor U13840 (N_13840,N_9459,N_10313);
nor U13841 (N_13841,N_10657,N_10593);
and U13842 (N_13842,N_10563,N_9872);
and U13843 (N_13843,N_12374,N_11779);
xor U13844 (N_13844,N_11120,N_10284);
nand U13845 (N_13845,N_11744,N_12014);
and U13846 (N_13846,N_11842,N_11763);
or U13847 (N_13847,N_11170,N_10561);
nand U13848 (N_13848,N_9985,N_12457);
nor U13849 (N_13849,N_11476,N_10498);
nand U13850 (N_13850,N_9921,N_9908);
nand U13851 (N_13851,N_12498,N_10550);
nand U13852 (N_13852,N_10359,N_9718);
xor U13853 (N_13853,N_11674,N_11099);
nand U13854 (N_13854,N_10349,N_10776);
and U13855 (N_13855,N_11824,N_10398);
xor U13856 (N_13856,N_10331,N_11643);
and U13857 (N_13857,N_11214,N_11229);
and U13858 (N_13858,N_10613,N_11187);
nor U13859 (N_13859,N_9980,N_11781);
nand U13860 (N_13860,N_11620,N_11365);
and U13861 (N_13861,N_9543,N_10712);
xor U13862 (N_13862,N_11091,N_10018);
nand U13863 (N_13863,N_10512,N_11988);
nand U13864 (N_13864,N_10357,N_12124);
nand U13865 (N_13865,N_11496,N_12303);
or U13866 (N_13866,N_9406,N_12065);
nand U13867 (N_13867,N_9437,N_10556);
nor U13868 (N_13868,N_10435,N_10306);
or U13869 (N_13869,N_10715,N_12007);
or U13870 (N_13870,N_12021,N_9713);
nand U13871 (N_13871,N_12312,N_11395);
or U13872 (N_13872,N_9655,N_10816);
or U13873 (N_13873,N_9748,N_9498);
and U13874 (N_13874,N_11691,N_9391);
nor U13875 (N_13875,N_10594,N_11883);
and U13876 (N_13876,N_9982,N_11582);
nor U13877 (N_13877,N_11117,N_11081);
and U13878 (N_13878,N_11337,N_12401);
and U13879 (N_13879,N_12266,N_12150);
nor U13880 (N_13880,N_11501,N_10142);
nor U13881 (N_13881,N_12482,N_10947);
nand U13882 (N_13882,N_12439,N_10402);
nand U13883 (N_13883,N_11839,N_9526);
and U13884 (N_13884,N_10451,N_12377);
and U13885 (N_13885,N_11210,N_11450);
nor U13886 (N_13886,N_10186,N_9892);
and U13887 (N_13887,N_12468,N_11969);
and U13888 (N_13888,N_10588,N_10365);
nand U13889 (N_13889,N_10737,N_12416);
nor U13890 (N_13890,N_12057,N_9598);
nor U13891 (N_13891,N_10079,N_12240);
or U13892 (N_13892,N_11772,N_10652);
and U13893 (N_13893,N_11612,N_9518);
nand U13894 (N_13894,N_11704,N_10383);
xor U13895 (N_13895,N_9533,N_11339);
nand U13896 (N_13896,N_11661,N_11263);
xnor U13897 (N_13897,N_10338,N_11851);
nor U13898 (N_13898,N_11549,N_9521);
xor U13899 (N_13899,N_12306,N_10183);
nand U13900 (N_13900,N_12209,N_12086);
nor U13901 (N_13901,N_10241,N_11124);
nor U13902 (N_13902,N_11696,N_10779);
and U13903 (N_13903,N_10683,N_11392);
or U13904 (N_13904,N_11889,N_10137);
and U13905 (N_13905,N_12076,N_11387);
xnor U13906 (N_13906,N_11119,N_11567);
and U13907 (N_13907,N_9741,N_10227);
and U13908 (N_13908,N_10047,N_9584);
xor U13909 (N_13909,N_10615,N_11059);
and U13910 (N_13910,N_9962,N_9412);
and U13911 (N_13911,N_11254,N_12002);
nor U13912 (N_13912,N_9649,N_10535);
nor U13913 (N_13913,N_11128,N_10369);
nand U13914 (N_13914,N_11904,N_11031);
and U13915 (N_13915,N_11311,N_10686);
nand U13916 (N_13916,N_10691,N_10728);
or U13917 (N_13917,N_11093,N_9737);
nor U13918 (N_13918,N_10300,N_10097);
nand U13919 (N_13919,N_11732,N_11001);
or U13920 (N_13920,N_11648,N_11649);
and U13921 (N_13921,N_9483,N_11566);
nor U13922 (N_13922,N_12254,N_9401);
or U13923 (N_13923,N_11308,N_11712);
xor U13924 (N_13924,N_11153,N_10485);
and U13925 (N_13925,N_9514,N_9638);
and U13926 (N_13926,N_10154,N_11841);
or U13927 (N_13927,N_10189,N_11446);
or U13928 (N_13928,N_10202,N_11944);
xnor U13929 (N_13929,N_9469,N_10497);
nor U13930 (N_13930,N_12289,N_10214);
or U13931 (N_13931,N_9923,N_9703);
nand U13932 (N_13932,N_11731,N_10488);
nand U13933 (N_13933,N_12227,N_10559);
or U13934 (N_13934,N_10449,N_11344);
nand U13935 (N_13935,N_11005,N_9615);
nor U13936 (N_13936,N_12010,N_11917);
or U13937 (N_13937,N_11222,N_9793);
or U13938 (N_13938,N_10665,N_12161);
or U13939 (N_13939,N_11315,N_10244);
nand U13940 (N_13940,N_11037,N_9944);
and U13941 (N_13941,N_11972,N_9381);
nor U13942 (N_13942,N_9377,N_10475);
nor U13943 (N_13943,N_11293,N_11488);
nor U13944 (N_13944,N_11516,N_9928);
and U13945 (N_13945,N_10345,N_12450);
and U13946 (N_13946,N_10484,N_11681);
nand U13947 (N_13947,N_9784,N_12089);
nand U13948 (N_13948,N_10187,N_11822);
nor U13949 (N_13949,N_11800,N_12305);
nor U13950 (N_13950,N_9818,N_11310);
nand U13951 (N_13951,N_10836,N_11009);
nand U13952 (N_13952,N_11798,N_10055);
nor U13953 (N_13953,N_11018,N_10134);
nor U13954 (N_13954,N_11072,N_12319);
nand U13955 (N_13955,N_10690,N_12063);
nor U13956 (N_13956,N_12016,N_11480);
nor U13957 (N_13957,N_12041,N_9497);
or U13958 (N_13958,N_11755,N_11038);
nor U13959 (N_13959,N_11862,N_11023);
and U13960 (N_13960,N_11121,N_9679);
or U13961 (N_13961,N_9621,N_9802);
nor U13962 (N_13962,N_11570,N_12255);
nand U13963 (N_13963,N_12465,N_10604);
and U13964 (N_13964,N_11780,N_12190);
nor U13965 (N_13965,N_12061,N_12366);
or U13966 (N_13966,N_11639,N_12082);
nand U13967 (N_13967,N_10247,N_9438);
and U13968 (N_13968,N_11708,N_11178);
and U13969 (N_13969,N_10462,N_9933);
and U13970 (N_13970,N_9395,N_10890);
nand U13971 (N_13971,N_11902,N_11340);
nand U13972 (N_13972,N_11203,N_9745);
xor U13973 (N_13973,N_12399,N_10551);
or U13974 (N_13974,N_12067,N_10694);
or U13975 (N_13975,N_10695,N_11255);
nor U13976 (N_13976,N_11616,N_10419);
nor U13977 (N_13977,N_11644,N_11593);
nand U13978 (N_13978,N_11454,N_11302);
and U13979 (N_13979,N_10887,N_12087);
nand U13980 (N_13980,N_10220,N_10967);
nand U13981 (N_13981,N_10273,N_11481);
nand U13982 (N_13982,N_10432,N_11486);
nand U13983 (N_13983,N_10140,N_11090);
and U13984 (N_13984,N_10656,N_12321);
nor U13985 (N_13985,N_11743,N_11662);
nor U13986 (N_13986,N_9570,N_9951);
nand U13987 (N_13987,N_11042,N_11997);
nand U13988 (N_13988,N_10225,N_11752);
xnor U13989 (N_13989,N_12129,N_12473);
nand U13990 (N_13990,N_11464,N_11591);
or U13991 (N_13991,N_11161,N_11821);
or U13992 (N_13992,N_10918,N_11292);
xnor U13993 (N_13993,N_11008,N_11142);
and U13994 (N_13994,N_10286,N_10280);
nand U13995 (N_13995,N_10966,N_11275);
or U13996 (N_13996,N_10514,N_9409);
and U13997 (N_13997,N_11401,N_9609);
and U13998 (N_13998,N_11104,N_12158);
nor U13999 (N_13999,N_9887,N_11634);
nor U14000 (N_14000,N_10299,N_11617);
and U14001 (N_14001,N_10845,N_9688);
or U14002 (N_14002,N_11873,N_11181);
nand U14003 (N_14003,N_11829,N_11759);
and U14004 (N_14004,N_12154,N_10315);
nor U14005 (N_14005,N_10954,N_9562);
or U14006 (N_14006,N_11180,N_10602);
xor U14007 (N_14007,N_12062,N_11448);
nand U14008 (N_14008,N_9457,N_10151);
nand U14009 (N_14009,N_11664,N_10983);
and U14010 (N_14010,N_10020,N_10702);
nor U14011 (N_14011,N_10609,N_10156);
xor U14012 (N_14012,N_11002,N_12173);
nand U14013 (N_14013,N_9966,N_10212);
and U14014 (N_14014,N_11650,N_10619);
and U14015 (N_14015,N_12385,N_10868);
nand U14016 (N_14016,N_10289,N_11671);
or U14017 (N_14017,N_10717,N_10408);
nand U14018 (N_14018,N_10219,N_11556);
or U14019 (N_14019,N_10718,N_10893);
nand U14020 (N_14020,N_9530,N_12160);
nor U14021 (N_14021,N_10356,N_11353);
nand U14022 (N_14022,N_11926,N_11934);
nand U14023 (N_14023,N_11739,N_10270);
nand U14024 (N_14024,N_12389,N_10567);
and U14025 (N_14025,N_11507,N_10666);
or U14026 (N_14026,N_10505,N_11107);
xnor U14027 (N_14027,N_11230,N_12084);
nand U14028 (N_14028,N_9456,N_12250);
or U14029 (N_14029,N_11248,N_11867);
nand U14030 (N_14030,N_10373,N_10626);
nand U14031 (N_14031,N_10587,N_10935);
and U14032 (N_14032,N_11462,N_10971);
and U14033 (N_14033,N_11196,N_12327);
nand U14034 (N_14034,N_12483,N_12109);
or U14035 (N_14035,N_11891,N_12362);
nand U14036 (N_14036,N_11284,N_10627);
nor U14037 (N_14037,N_10290,N_10669);
nor U14038 (N_14038,N_10260,N_11238);
and U14039 (N_14039,N_10817,N_9634);
or U14040 (N_14040,N_10958,N_11430);
or U14041 (N_14041,N_9699,N_9575);
nor U14042 (N_14042,N_11604,N_10213);
and U14043 (N_14043,N_10182,N_10730);
nand U14044 (N_14044,N_11083,N_9505);
or U14045 (N_14045,N_12096,N_12018);
nand U14046 (N_14046,N_11213,N_9432);
nand U14047 (N_14047,N_11216,N_11831);
xor U14048 (N_14048,N_10835,N_9776);
nor U14049 (N_14049,N_10522,N_10288);
and U14050 (N_14050,N_11286,N_11452);
nand U14051 (N_14051,N_10474,N_11733);
nand U14052 (N_14052,N_9387,N_11898);
or U14053 (N_14053,N_11791,N_11168);
xor U14054 (N_14054,N_9863,N_9936);
or U14055 (N_14055,N_11651,N_10084);
or U14056 (N_14056,N_11717,N_11710);
nand U14057 (N_14057,N_12186,N_11024);
or U14058 (N_14058,N_11110,N_9402);
xnor U14059 (N_14059,N_11393,N_10266);
or U14060 (N_14060,N_12239,N_9838);
nand U14061 (N_14061,N_11931,N_12177);
and U14062 (N_14062,N_10964,N_12035);
nand U14063 (N_14063,N_10933,N_10272);
or U14064 (N_14064,N_10604,N_12040);
nor U14065 (N_14065,N_12247,N_12387);
xnor U14066 (N_14066,N_10298,N_9536);
nor U14067 (N_14067,N_9499,N_10788);
nand U14068 (N_14068,N_10092,N_11319);
and U14069 (N_14069,N_11240,N_9562);
and U14070 (N_14070,N_11574,N_9700);
nand U14071 (N_14071,N_10494,N_9389);
or U14072 (N_14072,N_10941,N_12419);
and U14073 (N_14073,N_9828,N_11919);
nand U14074 (N_14074,N_11887,N_12237);
nor U14075 (N_14075,N_10440,N_12140);
nand U14076 (N_14076,N_11649,N_11737);
nor U14077 (N_14077,N_12035,N_10055);
or U14078 (N_14078,N_12131,N_11953);
nand U14079 (N_14079,N_10972,N_10664);
or U14080 (N_14080,N_11377,N_11215);
or U14081 (N_14081,N_9657,N_12324);
and U14082 (N_14082,N_9672,N_12034);
or U14083 (N_14083,N_11652,N_12164);
or U14084 (N_14084,N_12438,N_12354);
nand U14085 (N_14085,N_9924,N_11329);
or U14086 (N_14086,N_10097,N_11327);
nand U14087 (N_14087,N_9383,N_11276);
and U14088 (N_14088,N_12444,N_12211);
nor U14089 (N_14089,N_10971,N_9636);
nand U14090 (N_14090,N_9440,N_11813);
and U14091 (N_14091,N_10491,N_10899);
or U14092 (N_14092,N_11655,N_11660);
nor U14093 (N_14093,N_9772,N_11510);
nor U14094 (N_14094,N_11434,N_10116);
or U14095 (N_14095,N_10040,N_9779);
and U14096 (N_14096,N_10421,N_10497);
and U14097 (N_14097,N_10907,N_10031);
nand U14098 (N_14098,N_9472,N_10961);
xnor U14099 (N_14099,N_11978,N_10817);
and U14100 (N_14100,N_12440,N_10746);
nor U14101 (N_14101,N_9866,N_11444);
nor U14102 (N_14102,N_10034,N_10399);
nor U14103 (N_14103,N_12274,N_11704);
and U14104 (N_14104,N_11890,N_11861);
and U14105 (N_14105,N_10218,N_9769);
or U14106 (N_14106,N_10572,N_12151);
nor U14107 (N_14107,N_12164,N_9558);
and U14108 (N_14108,N_12087,N_9985);
and U14109 (N_14109,N_9804,N_9793);
nand U14110 (N_14110,N_10898,N_11210);
and U14111 (N_14111,N_10546,N_12273);
and U14112 (N_14112,N_11146,N_11732);
xnor U14113 (N_14113,N_10444,N_9913);
and U14114 (N_14114,N_10010,N_11759);
nand U14115 (N_14115,N_11985,N_10925);
and U14116 (N_14116,N_11146,N_11488);
xor U14117 (N_14117,N_9403,N_11775);
or U14118 (N_14118,N_9514,N_11117);
and U14119 (N_14119,N_11029,N_9442);
or U14120 (N_14120,N_9456,N_10641);
nor U14121 (N_14121,N_11974,N_10092);
or U14122 (N_14122,N_11258,N_11159);
and U14123 (N_14123,N_9609,N_12377);
and U14124 (N_14124,N_12098,N_11929);
and U14125 (N_14125,N_12469,N_10991);
nand U14126 (N_14126,N_9654,N_10475);
and U14127 (N_14127,N_10713,N_11254);
and U14128 (N_14128,N_10226,N_10324);
or U14129 (N_14129,N_10705,N_11452);
xor U14130 (N_14130,N_9850,N_11623);
xnor U14131 (N_14131,N_10344,N_11565);
or U14132 (N_14132,N_12415,N_12248);
and U14133 (N_14133,N_11264,N_9889);
xnor U14134 (N_14134,N_12233,N_10654);
nand U14135 (N_14135,N_10273,N_10943);
or U14136 (N_14136,N_10876,N_10707);
or U14137 (N_14137,N_9956,N_9890);
nor U14138 (N_14138,N_11329,N_11560);
nand U14139 (N_14139,N_11902,N_12217);
nand U14140 (N_14140,N_11711,N_9661);
nor U14141 (N_14141,N_10394,N_10223);
nor U14142 (N_14142,N_9482,N_10679);
nand U14143 (N_14143,N_11491,N_10102);
xor U14144 (N_14144,N_11955,N_12128);
nand U14145 (N_14145,N_9601,N_11761);
nand U14146 (N_14146,N_11886,N_11974);
nor U14147 (N_14147,N_9519,N_10182);
nor U14148 (N_14148,N_12067,N_9567);
nand U14149 (N_14149,N_11305,N_9393);
and U14150 (N_14150,N_11128,N_12465);
or U14151 (N_14151,N_11906,N_11898);
or U14152 (N_14152,N_10989,N_9816);
or U14153 (N_14153,N_12379,N_11210);
or U14154 (N_14154,N_9951,N_11621);
and U14155 (N_14155,N_10678,N_11419);
nand U14156 (N_14156,N_12476,N_9600);
nand U14157 (N_14157,N_9996,N_12188);
or U14158 (N_14158,N_10375,N_10595);
nor U14159 (N_14159,N_11649,N_12490);
xnor U14160 (N_14160,N_10825,N_11057);
nand U14161 (N_14161,N_10566,N_11856);
nand U14162 (N_14162,N_10311,N_10139);
nand U14163 (N_14163,N_9520,N_11674);
and U14164 (N_14164,N_11643,N_11238);
xnor U14165 (N_14165,N_11070,N_10231);
or U14166 (N_14166,N_9802,N_11788);
nand U14167 (N_14167,N_9683,N_11080);
or U14168 (N_14168,N_10211,N_11936);
nand U14169 (N_14169,N_10267,N_11098);
or U14170 (N_14170,N_12391,N_12243);
xnor U14171 (N_14171,N_12118,N_9802);
or U14172 (N_14172,N_11300,N_9919);
xnor U14173 (N_14173,N_11300,N_9958);
and U14174 (N_14174,N_9936,N_11258);
or U14175 (N_14175,N_11753,N_9888);
xor U14176 (N_14176,N_11116,N_9665);
and U14177 (N_14177,N_11625,N_11512);
or U14178 (N_14178,N_12263,N_10510);
and U14179 (N_14179,N_11118,N_10401);
and U14180 (N_14180,N_9516,N_12290);
or U14181 (N_14181,N_11324,N_10760);
nor U14182 (N_14182,N_12486,N_12253);
nor U14183 (N_14183,N_10761,N_10044);
nand U14184 (N_14184,N_11172,N_10838);
or U14185 (N_14185,N_10914,N_10142);
nor U14186 (N_14186,N_10997,N_11855);
and U14187 (N_14187,N_11068,N_10307);
or U14188 (N_14188,N_12207,N_11224);
or U14189 (N_14189,N_12222,N_10511);
and U14190 (N_14190,N_9396,N_9612);
and U14191 (N_14191,N_9820,N_11426);
nor U14192 (N_14192,N_10559,N_9740);
and U14193 (N_14193,N_9765,N_10064);
and U14194 (N_14194,N_12051,N_9607);
nand U14195 (N_14195,N_10989,N_10993);
xor U14196 (N_14196,N_10919,N_10393);
and U14197 (N_14197,N_9524,N_10108);
xor U14198 (N_14198,N_10330,N_11929);
and U14199 (N_14199,N_11150,N_11759);
xnor U14200 (N_14200,N_12389,N_11458);
or U14201 (N_14201,N_11697,N_10515);
nor U14202 (N_14202,N_12321,N_10393);
nor U14203 (N_14203,N_10678,N_9451);
nand U14204 (N_14204,N_11866,N_9615);
or U14205 (N_14205,N_10753,N_10235);
or U14206 (N_14206,N_10914,N_11026);
nand U14207 (N_14207,N_10275,N_11390);
and U14208 (N_14208,N_12207,N_10880);
or U14209 (N_14209,N_12289,N_11010);
nand U14210 (N_14210,N_11374,N_10460);
or U14211 (N_14211,N_11875,N_10057);
or U14212 (N_14212,N_10646,N_11007);
and U14213 (N_14213,N_11507,N_10436);
and U14214 (N_14214,N_9968,N_10463);
nor U14215 (N_14215,N_9654,N_9634);
nand U14216 (N_14216,N_11869,N_9514);
nor U14217 (N_14217,N_11883,N_12281);
nand U14218 (N_14218,N_9677,N_9724);
or U14219 (N_14219,N_9959,N_9659);
or U14220 (N_14220,N_10126,N_10254);
xnor U14221 (N_14221,N_10413,N_11729);
and U14222 (N_14222,N_11425,N_11126);
and U14223 (N_14223,N_10021,N_10128);
xor U14224 (N_14224,N_12277,N_11836);
and U14225 (N_14225,N_10864,N_10876);
and U14226 (N_14226,N_10460,N_10159);
nor U14227 (N_14227,N_10215,N_10528);
nand U14228 (N_14228,N_11058,N_9659);
or U14229 (N_14229,N_10586,N_12019);
nand U14230 (N_14230,N_11239,N_10092);
nand U14231 (N_14231,N_10512,N_11403);
nor U14232 (N_14232,N_12096,N_11596);
nand U14233 (N_14233,N_11892,N_12021);
nand U14234 (N_14234,N_10877,N_11754);
and U14235 (N_14235,N_11986,N_9442);
nor U14236 (N_14236,N_12323,N_9479);
nand U14237 (N_14237,N_11960,N_10462);
nand U14238 (N_14238,N_11208,N_11027);
and U14239 (N_14239,N_10268,N_10004);
nor U14240 (N_14240,N_11569,N_9967);
xor U14241 (N_14241,N_10546,N_10626);
nor U14242 (N_14242,N_10621,N_11827);
nand U14243 (N_14243,N_10838,N_9960);
and U14244 (N_14244,N_11605,N_10121);
and U14245 (N_14245,N_11619,N_11165);
nor U14246 (N_14246,N_11177,N_11568);
or U14247 (N_14247,N_9738,N_9760);
and U14248 (N_14248,N_12445,N_10836);
nor U14249 (N_14249,N_10548,N_10973);
or U14250 (N_14250,N_12229,N_11647);
or U14251 (N_14251,N_12307,N_9472);
nand U14252 (N_14252,N_11035,N_11147);
and U14253 (N_14253,N_10621,N_10869);
and U14254 (N_14254,N_11082,N_10092);
xnor U14255 (N_14255,N_10746,N_10996);
xnor U14256 (N_14256,N_9409,N_12334);
nand U14257 (N_14257,N_9810,N_11781);
or U14258 (N_14258,N_10852,N_11128);
xor U14259 (N_14259,N_9524,N_10629);
or U14260 (N_14260,N_12308,N_10499);
xor U14261 (N_14261,N_11108,N_10624);
or U14262 (N_14262,N_10680,N_11386);
and U14263 (N_14263,N_9980,N_10736);
xnor U14264 (N_14264,N_11099,N_10996);
and U14265 (N_14265,N_10231,N_12069);
nor U14266 (N_14266,N_9791,N_10603);
or U14267 (N_14267,N_11978,N_12448);
nor U14268 (N_14268,N_12116,N_12288);
and U14269 (N_14269,N_11757,N_11228);
or U14270 (N_14270,N_10856,N_11533);
and U14271 (N_14271,N_11383,N_11134);
nor U14272 (N_14272,N_12262,N_9745);
nor U14273 (N_14273,N_10576,N_11806);
nand U14274 (N_14274,N_11277,N_9789);
or U14275 (N_14275,N_12063,N_12470);
xor U14276 (N_14276,N_11858,N_10256);
or U14277 (N_14277,N_11170,N_11834);
nand U14278 (N_14278,N_12018,N_12373);
and U14279 (N_14279,N_11049,N_11132);
and U14280 (N_14280,N_11298,N_12412);
or U14281 (N_14281,N_9552,N_11448);
and U14282 (N_14282,N_10272,N_11401);
and U14283 (N_14283,N_11454,N_9731);
nand U14284 (N_14284,N_11068,N_10864);
nand U14285 (N_14285,N_12108,N_10049);
and U14286 (N_14286,N_12084,N_10405);
nand U14287 (N_14287,N_10779,N_11380);
or U14288 (N_14288,N_11667,N_11416);
nor U14289 (N_14289,N_10978,N_12000);
nand U14290 (N_14290,N_9683,N_10798);
nand U14291 (N_14291,N_9664,N_10658);
nand U14292 (N_14292,N_10542,N_11785);
nor U14293 (N_14293,N_10652,N_9597);
or U14294 (N_14294,N_9776,N_9603);
and U14295 (N_14295,N_12293,N_10994);
nor U14296 (N_14296,N_11158,N_10235);
xor U14297 (N_14297,N_11657,N_10210);
nand U14298 (N_14298,N_11613,N_12481);
and U14299 (N_14299,N_11733,N_12265);
nand U14300 (N_14300,N_10028,N_11907);
and U14301 (N_14301,N_11950,N_10607);
and U14302 (N_14302,N_9745,N_11601);
or U14303 (N_14303,N_12301,N_12336);
nand U14304 (N_14304,N_11050,N_11945);
nor U14305 (N_14305,N_10095,N_11585);
xnor U14306 (N_14306,N_12398,N_10440);
nand U14307 (N_14307,N_10986,N_9493);
nand U14308 (N_14308,N_11649,N_9781);
or U14309 (N_14309,N_11653,N_11375);
and U14310 (N_14310,N_11798,N_9408);
and U14311 (N_14311,N_11588,N_9934);
nor U14312 (N_14312,N_9552,N_11364);
or U14313 (N_14313,N_9627,N_11853);
and U14314 (N_14314,N_11527,N_10853);
xor U14315 (N_14315,N_11464,N_9799);
nand U14316 (N_14316,N_11989,N_9935);
and U14317 (N_14317,N_10294,N_10223);
and U14318 (N_14318,N_11384,N_11172);
or U14319 (N_14319,N_11480,N_12427);
nor U14320 (N_14320,N_10456,N_12269);
nor U14321 (N_14321,N_10118,N_9901);
nor U14322 (N_14322,N_10075,N_11678);
and U14323 (N_14323,N_12475,N_11713);
or U14324 (N_14324,N_11185,N_10913);
nand U14325 (N_14325,N_11025,N_10116);
nand U14326 (N_14326,N_9890,N_9792);
or U14327 (N_14327,N_12133,N_11862);
or U14328 (N_14328,N_10987,N_11898);
nor U14329 (N_14329,N_9574,N_10730);
and U14330 (N_14330,N_11730,N_11130);
nor U14331 (N_14331,N_10770,N_9652);
and U14332 (N_14332,N_9880,N_11100);
nor U14333 (N_14333,N_11649,N_10202);
nor U14334 (N_14334,N_11902,N_10051);
nand U14335 (N_14335,N_11622,N_9899);
xor U14336 (N_14336,N_12323,N_10903);
xor U14337 (N_14337,N_11864,N_11647);
or U14338 (N_14338,N_11313,N_12130);
or U14339 (N_14339,N_11928,N_11910);
or U14340 (N_14340,N_10767,N_9965);
nand U14341 (N_14341,N_10652,N_11162);
nor U14342 (N_14342,N_10145,N_10208);
nor U14343 (N_14343,N_10492,N_11624);
xnor U14344 (N_14344,N_11123,N_11696);
or U14345 (N_14345,N_11866,N_9769);
nor U14346 (N_14346,N_11087,N_10056);
nand U14347 (N_14347,N_11496,N_12404);
nor U14348 (N_14348,N_11770,N_9439);
nor U14349 (N_14349,N_10159,N_10369);
or U14350 (N_14350,N_11993,N_10629);
or U14351 (N_14351,N_11464,N_11055);
nand U14352 (N_14352,N_12279,N_10707);
or U14353 (N_14353,N_10286,N_9410);
nor U14354 (N_14354,N_12228,N_12114);
nand U14355 (N_14355,N_10472,N_11890);
and U14356 (N_14356,N_9409,N_12080);
nand U14357 (N_14357,N_9422,N_10584);
nand U14358 (N_14358,N_9422,N_10262);
and U14359 (N_14359,N_11597,N_12424);
nor U14360 (N_14360,N_12268,N_12071);
nor U14361 (N_14361,N_12015,N_12056);
and U14362 (N_14362,N_11611,N_10418);
xnor U14363 (N_14363,N_10572,N_9608);
and U14364 (N_14364,N_9671,N_11579);
or U14365 (N_14365,N_9805,N_9944);
xnor U14366 (N_14366,N_12151,N_12294);
and U14367 (N_14367,N_10311,N_10010);
or U14368 (N_14368,N_11923,N_10873);
nand U14369 (N_14369,N_12267,N_10576);
nor U14370 (N_14370,N_10331,N_10060);
or U14371 (N_14371,N_10610,N_11259);
or U14372 (N_14372,N_10361,N_12076);
nand U14373 (N_14373,N_11617,N_10226);
nand U14374 (N_14374,N_11377,N_9953);
nand U14375 (N_14375,N_11927,N_10460);
or U14376 (N_14376,N_10081,N_12067);
xnor U14377 (N_14377,N_10942,N_11544);
or U14378 (N_14378,N_10224,N_9490);
xor U14379 (N_14379,N_9482,N_11273);
nor U14380 (N_14380,N_11508,N_9932);
and U14381 (N_14381,N_11874,N_11082);
or U14382 (N_14382,N_12051,N_12246);
nand U14383 (N_14383,N_10519,N_12142);
or U14384 (N_14384,N_12409,N_9458);
or U14385 (N_14385,N_10623,N_10463);
xor U14386 (N_14386,N_10762,N_11757);
or U14387 (N_14387,N_10657,N_10255);
or U14388 (N_14388,N_10399,N_10099);
nand U14389 (N_14389,N_10713,N_10872);
or U14390 (N_14390,N_12292,N_10295);
and U14391 (N_14391,N_9589,N_12288);
and U14392 (N_14392,N_9641,N_12497);
and U14393 (N_14393,N_12005,N_10130);
nand U14394 (N_14394,N_9736,N_10261);
or U14395 (N_14395,N_11772,N_11929);
nor U14396 (N_14396,N_10229,N_9420);
xor U14397 (N_14397,N_9410,N_11673);
nor U14398 (N_14398,N_10219,N_11010);
and U14399 (N_14399,N_11495,N_10500);
nand U14400 (N_14400,N_11101,N_11022);
or U14401 (N_14401,N_11178,N_10308);
and U14402 (N_14402,N_9600,N_10285);
nand U14403 (N_14403,N_9660,N_11913);
or U14404 (N_14404,N_10113,N_12440);
nor U14405 (N_14405,N_11826,N_11127);
nor U14406 (N_14406,N_11914,N_12126);
xor U14407 (N_14407,N_12004,N_9681);
nor U14408 (N_14408,N_9428,N_11858);
and U14409 (N_14409,N_10601,N_12320);
or U14410 (N_14410,N_9491,N_10150);
nor U14411 (N_14411,N_10171,N_11762);
or U14412 (N_14412,N_9445,N_11613);
and U14413 (N_14413,N_9757,N_10098);
and U14414 (N_14414,N_10412,N_9961);
or U14415 (N_14415,N_10646,N_11713);
nor U14416 (N_14416,N_11478,N_11309);
nor U14417 (N_14417,N_12199,N_11499);
or U14418 (N_14418,N_10311,N_11840);
nand U14419 (N_14419,N_10613,N_12179);
or U14420 (N_14420,N_11232,N_11587);
and U14421 (N_14421,N_9598,N_9941);
nand U14422 (N_14422,N_10686,N_11177);
nand U14423 (N_14423,N_11967,N_10697);
or U14424 (N_14424,N_12379,N_10663);
and U14425 (N_14425,N_11247,N_11292);
xor U14426 (N_14426,N_11049,N_12384);
nand U14427 (N_14427,N_10089,N_9718);
and U14428 (N_14428,N_11488,N_12436);
and U14429 (N_14429,N_10274,N_11694);
nor U14430 (N_14430,N_10687,N_10705);
and U14431 (N_14431,N_11362,N_12176);
xnor U14432 (N_14432,N_12350,N_12385);
xnor U14433 (N_14433,N_9605,N_11099);
xnor U14434 (N_14434,N_12315,N_11610);
or U14435 (N_14435,N_11818,N_9538);
nor U14436 (N_14436,N_11525,N_11211);
xnor U14437 (N_14437,N_11376,N_11689);
and U14438 (N_14438,N_11044,N_10726);
nand U14439 (N_14439,N_9580,N_11949);
nand U14440 (N_14440,N_10501,N_11491);
or U14441 (N_14441,N_11585,N_11800);
nor U14442 (N_14442,N_9456,N_11048);
nand U14443 (N_14443,N_10257,N_10148);
nor U14444 (N_14444,N_10675,N_11609);
xor U14445 (N_14445,N_10882,N_11501);
nand U14446 (N_14446,N_11207,N_11834);
or U14447 (N_14447,N_10002,N_9946);
nand U14448 (N_14448,N_9808,N_11478);
nor U14449 (N_14449,N_12391,N_11777);
nand U14450 (N_14450,N_12359,N_11257);
nor U14451 (N_14451,N_9798,N_11906);
nor U14452 (N_14452,N_11016,N_11831);
xnor U14453 (N_14453,N_10528,N_11651);
or U14454 (N_14454,N_10700,N_10390);
or U14455 (N_14455,N_11617,N_9779);
or U14456 (N_14456,N_9781,N_10588);
or U14457 (N_14457,N_11397,N_12445);
nand U14458 (N_14458,N_9617,N_10188);
nor U14459 (N_14459,N_11181,N_11717);
nor U14460 (N_14460,N_11061,N_11569);
nand U14461 (N_14461,N_10218,N_9812);
nand U14462 (N_14462,N_11273,N_10386);
and U14463 (N_14463,N_11224,N_11257);
nand U14464 (N_14464,N_12488,N_11550);
and U14465 (N_14465,N_10176,N_12266);
or U14466 (N_14466,N_11594,N_10155);
nand U14467 (N_14467,N_12462,N_12466);
xor U14468 (N_14468,N_9465,N_9533);
and U14469 (N_14469,N_11571,N_11790);
or U14470 (N_14470,N_11498,N_11529);
nor U14471 (N_14471,N_11902,N_11067);
xor U14472 (N_14472,N_9816,N_10637);
xnor U14473 (N_14473,N_11397,N_10293);
and U14474 (N_14474,N_12109,N_9973);
and U14475 (N_14475,N_11810,N_12396);
nand U14476 (N_14476,N_12212,N_10673);
nor U14477 (N_14477,N_11960,N_10956);
nor U14478 (N_14478,N_11883,N_10984);
xnor U14479 (N_14479,N_12121,N_11818);
nor U14480 (N_14480,N_11278,N_9502);
nand U14481 (N_14481,N_10703,N_10760);
nor U14482 (N_14482,N_10221,N_10083);
or U14483 (N_14483,N_12396,N_10780);
nand U14484 (N_14484,N_12409,N_12227);
nor U14485 (N_14485,N_9793,N_9745);
xnor U14486 (N_14486,N_12099,N_11387);
and U14487 (N_14487,N_10391,N_10097);
and U14488 (N_14488,N_10744,N_11532);
xor U14489 (N_14489,N_12117,N_11549);
nand U14490 (N_14490,N_9573,N_11418);
nand U14491 (N_14491,N_11613,N_9932);
nand U14492 (N_14492,N_10189,N_10860);
xor U14493 (N_14493,N_10330,N_11014);
xnor U14494 (N_14494,N_11052,N_11075);
nand U14495 (N_14495,N_10266,N_11396);
and U14496 (N_14496,N_10875,N_10776);
or U14497 (N_14497,N_9819,N_12337);
nor U14498 (N_14498,N_12323,N_10171);
and U14499 (N_14499,N_10152,N_10112);
nand U14500 (N_14500,N_12319,N_11870);
or U14501 (N_14501,N_10378,N_10668);
or U14502 (N_14502,N_11272,N_11253);
and U14503 (N_14503,N_10070,N_9997);
and U14504 (N_14504,N_9626,N_11014);
nor U14505 (N_14505,N_11430,N_12010);
nand U14506 (N_14506,N_11632,N_12077);
nor U14507 (N_14507,N_11406,N_10211);
and U14508 (N_14508,N_10319,N_12098);
or U14509 (N_14509,N_10978,N_10458);
xor U14510 (N_14510,N_12193,N_11584);
and U14511 (N_14511,N_10048,N_10755);
or U14512 (N_14512,N_11779,N_11428);
and U14513 (N_14513,N_11455,N_11184);
xnor U14514 (N_14514,N_11461,N_12023);
or U14515 (N_14515,N_10662,N_11586);
or U14516 (N_14516,N_10252,N_9650);
nand U14517 (N_14517,N_11512,N_12073);
nor U14518 (N_14518,N_12096,N_9770);
nor U14519 (N_14519,N_10894,N_10427);
or U14520 (N_14520,N_10281,N_10769);
or U14521 (N_14521,N_11066,N_12492);
or U14522 (N_14522,N_10734,N_12219);
nand U14523 (N_14523,N_12474,N_10211);
nor U14524 (N_14524,N_10280,N_12278);
or U14525 (N_14525,N_11225,N_9382);
or U14526 (N_14526,N_9486,N_11114);
or U14527 (N_14527,N_11258,N_12025);
and U14528 (N_14528,N_9595,N_11023);
and U14529 (N_14529,N_10452,N_9792);
nor U14530 (N_14530,N_12037,N_10746);
and U14531 (N_14531,N_11392,N_10931);
xnor U14532 (N_14532,N_10337,N_9628);
nand U14533 (N_14533,N_11314,N_12295);
nand U14534 (N_14534,N_11002,N_10686);
or U14535 (N_14535,N_9425,N_10255);
nor U14536 (N_14536,N_12389,N_12101);
xnor U14537 (N_14537,N_9592,N_10725);
or U14538 (N_14538,N_10185,N_11284);
xor U14539 (N_14539,N_12289,N_11213);
and U14540 (N_14540,N_11422,N_9963);
nor U14541 (N_14541,N_11761,N_11396);
or U14542 (N_14542,N_11720,N_10936);
and U14543 (N_14543,N_9771,N_11141);
or U14544 (N_14544,N_10687,N_10220);
nor U14545 (N_14545,N_10286,N_9814);
nor U14546 (N_14546,N_12283,N_9535);
nand U14547 (N_14547,N_9922,N_11025);
nor U14548 (N_14548,N_11545,N_9936);
or U14549 (N_14549,N_9989,N_10379);
nand U14550 (N_14550,N_11954,N_12401);
or U14551 (N_14551,N_11057,N_9709);
nor U14552 (N_14552,N_12401,N_10095);
xnor U14553 (N_14553,N_9470,N_10242);
xor U14554 (N_14554,N_10547,N_10739);
nand U14555 (N_14555,N_12323,N_11142);
nor U14556 (N_14556,N_11687,N_11174);
nor U14557 (N_14557,N_10160,N_9431);
nand U14558 (N_14558,N_10506,N_10520);
or U14559 (N_14559,N_9957,N_11177);
and U14560 (N_14560,N_9737,N_11135);
nand U14561 (N_14561,N_11249,N_12003);
nand U14562 (N_14562,N_11801,N_11535);
and U14563 (N_14563,N_10647,N_11576);
nand U14564 (N_14564,N_9864,N_10380);
nand U14565 (N_14565,N_9443,N_11494);
and U14566 (N_14566,N_10593,N_12408);
or U14567 (N_14567,N_10476,N_11173);
xnor U14568 (N_14568,N_10610,N_11160);
nand U14569 (N_14569,N_10759,N_9957);
nand U14570 (N_14570,N_10573,N_9438);
or U14571 (N_14571,N_11893,N_10801);
and U14572 (N_14572,N_9630,N_11331);
or U14573 (N_14573,N_9534,N_12335);
nor U14574 (N_14574,N_10943,N_9908);
or U14575 (N_14575,N_9707,N_10458);
nor U14576 (N_14576,N_9877,N_12369);
nand U14577 (N_14577,N_12011,N_12399);
nor U14578 (N_14578,N_12001,N_11338);
nor U14579 (N_14579,N_12153,N_9650);
or U14580 (N_14580,N_11179,N_11040);
xnor U14581 (N_14581,N_9807,N_11520);
and U14582 (N_14582,N_10638,N_9499);
or U14583 (N_14583,N_9665,N_10790);
nand U14584 (N_14584,N_10816,N_9912);
nand U14585 (N_14585,N_10591,N_9955);
or U14586 (N_14586,N_12005,N_11790);
nand U14587 (N_14587,N_9910,N_11760);
xor U14588 (N_14588,N_11871,N_12319);
xor U14589 (N_14589,N_12390,N_10151);
nor U14590 (N_14590,N_12293,N_9689);
or U14591 (N_14591,N_9392,N_10045);
nor U14592 (N_14592,N_9531,N_11689);
and U14593 (N_14593,N_11584,N_11110);
xnor U14594 (N_14594,N_9785,N_10697);
or U14595 (N_14595,N_12362,N_9620);
nor U14596 (N_14596,N_11228,N_9491);
or U14597 (N_14597,N_12441,N_10525);
xor U14598 (N_14598,N_10121,N_11779);
nor U14599 (N_14599,N_9716,N_11922);
or U14600 (N_14600,N_11206,N_11082);
and U14601 (N_14601,N_9505,N_10457);
nand U14602 (N_14602,N_12485,N_11037);
nor U14603 (N_14603,N_10956,N_11503);
and U14604 (N_14604,N_10779,N_10388);
xnor U14605 (N_14605,N_10709,N_11820);
or U14606 (N_14606,N_10078,N_12130);
or U14607 (N_14607,N_9573,N_10882);
xor U14608 (N_14608,N_11554,N_11679);
nor U14609 (N_14609,N_11379,N_10295);
or U14610 (N_14610,N_9920,N_10609);
and U14611 (N_14611,N_9944,N_10851);
xor U14612 (N_14612,N_12201,N_12048);
nor U14613 (N_14613,N_10490,N_10105);
xnor U14614 (N_14614,N_11157,N_9695);
nand U14615 (N_14615,N_11128,N_10870);
and U14616 (N_14616,N_9515,N_11628);
nand U14617 (N_14617,N_10023,N_9422);
or U14618 (N_14618,N_9442,N_11669);
nand U14619 (N_14619,N_10887,N_12276);
nor U14620 (N_14620,N_9737,N_11121);
xor U14621 (N_14621,N_10501,N_11810);
xnor U14622 (N_14622,N_11003,N_9616);
nand U14623 (N_14623,N_11135,N_11270);
xnor U14624 (N_14624,N_12472,N_10850);
nand U14625 (N_14625,N_12439,N_11556);
and U14626 (N_14626,N_11094,N_10026);
nand U14627 (N_14627,N_12117,N_11494);
and U14628 (N_14628,N_11319,N_9784);
and U14629 (N_14629,N_10561,N_11041);
or U14630 (N_14630,N_10860,N_11739);
and U14631 (N_14631,N_9381,N_10970);
nand U14632 (N_14632,N_11909,N_9687);
nor U14633 (N_14633,N_10584,N_10565);
and U14634 (N_14634,N_9902,N_12410);
or U14635 (N_14635,N_12128,N_11284);
nand U14636 (N_14636,N_10856,N_11821);
nor U14637 (N_14637,N_9411,N_12023);
xnor U14638 (N_14638,N_11030,N_9793);
and U14639 (N_14639,N_10333,N_11793);
xnor U14640 (N_14640,N_10426,N_9956);
and U14641 (N_14641,N_9383,N_11865);
and U14642 (N_14642,N_10166,N_11625);
nor U14643 (N_14643,N_11341,N_11762);
nand U14644 (N_14644,N_11496,N_11568);
xor U14645 (N_14645,N_11520,N_11772);
nand U14646 (N_14646,N_9990,N_11590);
nand U14647 (N_14647,N_10396,N_10671);
and U14648 (N_14648,N_10026,N_11080);
nand U14649 (N_14649,N_12113,N_10758);
nand U14650 (N_14650,N_10359,N_11253);
nand U14651 (N_14651,N_10078,N_11954);
nand U14652 (N_14652,N_9529,N_9513);
and U14653 (N_14653,N_11062,N_11364);
nor U14654 (N_14654,N_10739,N_12269);
and U14655 (N_14655,N_12393,N_12343);
nor U14656 (N_14656,N_10040,N_9600);
nor U14657 (N_14657,N_11452,N_10024);
nand U14658 (N_14658,N_10526,N_9586);
nor U14659 (N_14659,N_10460,N_9581);
nand U14660 (N_14660,N_12143,N_9779);
nand U14661 (N_14661,N_10007,N_9717);
xnor U14662 (N_14662,N_12006,N_9398);
and U14663 (N_14663,N_10962,N_10372);
or U14664 (N_14664,N_9620,N_12143);
nand U14665 (N_14665,N_9903,N_11267);
and U14666 (N_14666,N_10842,N_10286);
xnor U14667 (N_14667,N_10965,N_11771);
and U14668 (N_14668,N_10062,N_11853);
nor U14669 (N_14669,N_12094,N_11775);
and U14670 (N_14670,N_10236,N_12026);
or U14671 (N_14671,N_10962,N_12245);
nor U14672 (N_14672,N_11351,N_9747);
xnor U14673 (N_14673,N_11338,N_11277);
xor U14674 (N_14674,N_11700,N_10770);
and U14675 (N_14675,N_12109,N_12284);
nand U14676 (N_14676,N_11691,N_11513);
and U14677 (N_14677,N_10031,N_12013);
nor U14678 (N_14678,N_10499,N_11255);
or U14679 (N_14679,N_12212,N_11028);
nor U14680 (N_14680,N_11071,N_10321);
or U14681 (N_14681,N_11594,N_11308);
nand U14682 (N_14682,N_9629,N_9525);
and U14683 (N_14683,N_9544,N_11021);
and U14684 (N_14684,N_11948,N_9811);
nor U14685 (N_14685,N_9381,N_11103);
nand U14686 (N_14686,N_10771,N_9679);
nand U14687 (N_14687,N_9635,N_9930);
xor U14688 (N_14688,N_10988,N_9938);
nand U14689 (N_14689,N_9979,N_10961);
or U14690 (N_14690,N_11782,N_11479);
or U14691 (N_14691,N_12433,N_9601);
and U14692 (N_14692,N_10226,N_11394);
and U14693 (N_14693,N_10035,N_10501);
xnor U14694 (N_14694,N_11260,N_10313);
and U14695 (N_14695,N_9956,N_12463);
or U14696 (N_14696,N_9640,N_12179);
nand U14697 (N_14697,N_11432,N_10376);
nand U14698 (N_14698,N_9429,N_9449);
nor U14699 (N_14699,N_11370,N_11941);
or U14700 (N_14700,N_12392,N_9497);
nand U14701 (N_14701,N_10673,N_11884);
nand U14702 (N_14702,N_10969,N_10770);
nand U14703 (N_14703,N_9581,N_11312);
and U14704 (N_14704,N_9712,N_12304);
nor U14705 (N_14705,N_9389,N_10747);
and U14706 (N_14706,N_11664,N_10165);
nand U14707 (N_14707,N_12209,N_11653);
nand U14708 (N_14708,N_11435,N_11116);
or U14709 (N_14709,N_12488,N_10303);
xnor U14710 (N_14710,N_11151,N_9672);
or U14711 (N_14711,N_10280,N_9959);
or U14712 (N_14712,N_9415,N_11103);
nand U14713 (N_14713,N_12003,N_12393);
or U14714 (N_14714,N_11124,N_12152);
or U14715 (N_14715,N_10449,N_11798);
or U14716 (N_14716,N_11817,N_10584);
or U14717 (N_14717,N_12374,N_11589);
and U14718 (N_14718,N_10830,N_11716);
nor U14719 (N_14719,N_9748,N_9728);
or U14720 (N_14720,N_10353,N_9784);
or U14721 (N_14721,N_10081,N_9483);
or U14722 (N_14722,N_12288,N_9798);
nor U14723 (N_14723,N_10792,N_9614);
and U14724 (N_14724,N_11808,N_10622);
nand U14725 (N_14725,N_11109,N_9693);
nor U14726 (N_14726,N_9839,N_11703);
or U14727 (N_14727,N_10263,N_10432);
nor U14728 (N_14728,N_9517,N_10483);
and U14729 (N_14729,N_9429,N_10698);
and U14730 (N_14730,N_10998,N_11918);
and U14731 (N_14731,N_11030,N_11100);
nand U14732 (N_14732,N_9866,N_9950);
nor U14733 (N_14733,N_9809,N_12358);
and U14734 (N_14734,N_12475,N_10224);
and U14735 (N_14735,N_12339,N_11563);
nand U14736 (N_14736,N_9946,N_11041);
xnor U14737 (N_14737,N_12483,N_11541);
nor U14738 (N_14738,N_12305,N_10376);
and U14739 (N_14739,N_10862,N_10561);
nand U14740 (N_14740,N_12355,N_10928);
or U14741 (N_14741,N_9969,N_12390);
or U14742 (N_14742,N_11759,N_11458);
nor U14743 (N_14743,N_10706,N_9880);
and U14744 (N_14744,N_10256,N_10667);
and U14745 (N_14745,N_11233,N_11846);
nand U14746 (N_14746,N_10812,N_10491);
nor U14747 (N_14747,N_9867,N_10887);
and U14748 (N_14748,N_10606,N_11969);
nand U14749 (N_14749,N_9821,N_12055);
xor U14750 (N_14750,N_10005,N_12382);
nor U14751 (N_14751,N_12045,N_10427);
nor U14752 (N_14752,N_10361,N_12439);
nor U14753 (N_14753,N_11085,N_10314);
xor U14754 (N_14754,N_12316,N_9440);
or U14755 (N_14755,N_10735,N_11231);
xnor U14756 (N_14756,N_12354,N_9610);
or U14757 (N_14757,N_11917,N_12048);
nand U14758 (N_14758,N_10828,N_11879);
nor U14759 (N_14759,N_9650,N_9421);
nor U14760 (N_14760,N_12368,N_11271);
or U14761 (N_14761,N_12045,N_9819);
nand U14762 (N_14762,N_10843,N_11878);
nand U14763 (N_14763,N_12059,N_11364);
or U14764 (N_14764,N_11847,N_9631);
nor U14765 (N_14765,N_10943,N_10611);
nand U14766 (N_14766,N_10552,N_11121);
or U14767 (N_14767,N_12320,N_11421);
nand U14768 (N_14768,N_10290,N_11119);
nor U14769 (N_14769,N_9973,N_10563);
and U14770 (N_14770,N_12042,N_11876);
nor U14771 (N_14771,N_10902,N_11149);
and U14772 (N_14772,N_9957,N_9558);
nand U14773 (N_14773,N_11585,N_9650);
or U14774 (N_14774,N_11495,N_10890);
or U14775 (N_14775,N_9990,N_11163);
nor U14776 (N_14776,N_10126,N_10788);
or U14777 (N_14777,N_9521,N_11706);
nand U14778 (N_14778,N_11119,N_11957);
nand U14779 (N_14779,N_9735,N_10051);
or U14780 (N_14780,N_10471,N_10684);
or U14781 (N_14781,N_9971,N_12214);
or U14782 (N_14782,N_9608,N_11196);
nor U14783 (N_14783,N_9851,N_10056);
nor U14784 (N_14784,N_10910,N_9840);
nand U14785 (N_14785,N_10229,N_10895);
or U14786 (N_14786,N_10901,N_10321);
nand U14787 (N_14787,N_10699,N_9404);
or U14788 (N_14788,N_12493,N_12343);
nand U14789 (N_14789,N_9624,N_10541);
xnor U14790 (N_14790,N_11844,N_9816);
or U14791 (N_14791,N_12377,N_10930);
or U14792 (N_14792,N_12149,N_9814);
nand U14793 (N_14793,N_10135,N_12380);
and U14794 (N_14794,N_11462,N_11961);
nor U14795 (N_14795,N_10312,N_11703);
and U14796 (N_14796,N_12367,N_12466);
nand U14797 (N_14797,N_12174,N_10463);
and U14798 (N_14798,N_9877,N_10982);
or U14799 (N_14799,N_10822,N_11170);
and U14800 (N_14800,N_12088,N_12289);
and U14801 (N_14801,N_9559,N_12321);
nand U14802 (N_14802,N_12079,N_11816);
nor U14803 (N_14803,N_11259,N_11037);
or U14804 (N_14804,N_12231,N_12459);
nand U14805 (N_14805,N_9878,N_10969);
nor U14806 (N_14806,N_9672,N_11047);
nor U14807 (N_14807,N_12366,N_9541);
or U14808 (N_14808,N_10053,N_9839);
nor U14809 (N_14809,N_9538,N_11508);
and U14810 (N_14810,N_11624,N_12373);
or U14811 (N_14811,N_9668,N_10955);
nor U14812 (N_14812,N_10151,N_10094);
nor U14813 (N_14813,N_11715,N_11442);
nor U14814 (N_14814,N_10577,N_10159);
and U14815 (N_14815,N_11540,N_11743);
or U14816 (N_14816,N_11937,N_10940);
nor U14817 (N_14817,N_10203,N_12248);
and U14818 (N_14818,N_10650,N_9911);
nand U14819 (N_14819,N_11350,N_11243);
xor U14820 (N_14820,N_10797,N_12428);
and U14821 (N_14821,N_9478,N_10148);
or U14822 (N_14822,N_12220,N_11140);
nor U14823 (N_14823,N_9607,N_9952);
nand U14824 (N_14824,N_11464,N_9969);
nand U14825 (N_14825,N_10849,N_12324);
xor U14826 (N_14826,N_10243,N_9437);
nand U14827 (N_14827,N_11598,N_11480);
nor U14828 (N_14828,N_9799,N_11807);
nor U14829 (N_14829,N_12453,N_11065);
nor U14830 (N_14830,N_9583,N_9755);
or U14831 (N_14831,N_12370,N_11842);
xnor U14832 (N_14832,N_11789,N_11000);
and U14833 (N_14833,N_9471,N_10822);
nand U14834 (N_14834,N_12325,N_11236);
and U14835 (N_14835,N_11954,N_12407);
nor U14836 (N_14836,N_10265,N_10721);
nor U14837 (N_14837,N_9500,N_11005);
or U14838 (N_14838,N_9886,N_9800);
or U14839 (N_14839,N_11050,N_10278);
nor U14840 (N_14840,N_9861,N_11708);
and U14841 (N_14841,N_10386,N_11336);
nor U14842 (N_14842,N_11290,N_11477);
and U14843 (N_14843,N_10183,N_11995);
and U14844 (N_14844,N_9383,N_11158);
and U14845 (N_14845,N_11392,N_11853);
nand U14846 (N_14846,N_10731,N_9915);
nor U14847 (N_14847,N_11373,N_12378);
nand U14848 (N_14848,N_10641,N_9429);
nand U14849 (N_14849,N_12408,N_10107);
or U14850 (N_14850,N_10221,N_9816);
nand U14851 (N_14851,N_10078,N_12336);
nand U14852 (N_14852,N_12041,N_10214);
and U14853 (N_14853,N_12077,N_9922);
xnor U14854 (N_14854,N_11829,N_12318);
nand U14855 (N_14855,N_9947,N_9593);
nor U14856 (N_14856,N_12309,N_12270);
xnor U14857 (N_14857,N_12044,N_9667);
xor U14858 (N_14858,N_10684,N_12292);
nor U14859 (N_14859,N_10322,N_11704);
or U14860 (N_14860,N_9423,N_9828);
and U14861 (N_14861,N_11412,N_11279);
or U14862 (N_14862,N_9744,N_11081);
nor U14863 (N_14863,N_11479,N_11887);
xnor U14864 (N_14864,N_11015,N_11101);
and U14865 (N_14865,N_11893,N_11648);
or U14866 (N_14866,N_9751,N_9550);
nor U14867 (N_14867,N_9966,N_10935);
xor U14868 (N_14868,N_10166,N_10301);
nor U14869 (N_14869,N_12145,N_10136);
and U14870 (N_14870,N_11354,N_9482);
nor U14871 (N_14871,N_9787,N_9914);
and U14872 (N_14872,N_10101,N_11824);
and U14873 (N_14873,N_12057,N_11673);
or U14874 (N_14874,N_11565,N_12154);
nor U14875 (N_14875,N_9706,N_11437);
nor U14876 (N_14876,N_11768,N_11754);
xnor U14877 (N_14877,N_11728,N_11680);
nand U14878 (N_14878,N_11816,N_9387);
or U14879 (N_14879,N_12376,N_10912);
and U14880 (N_14880,N_12204,N_9400);
nor U14881 (N_14881,N_10455,N_11347);
or U14882 (N_14882,N_10654,N_12364);
xor U14883 (N_14883,N_10255,N_11992);
or U14884 (N_14884,N_10622,N_10645);
and U14885 (N_14885,N_11486,N_10171);
and U14886 (N_14886,N_11174,N_11570);
xnor U14887 (N_14887,N_11866,N_11830);
and U14888 (N_14888,N_11595,N_11456);
nor U14889 (N_14889,N_9497,N_10019);
or U14890 (N_14890,N_12274,N_10817);
nor U14891 (N_14891,N_11066,N_10427);
and U14892 (N_14892,N_10201,N_11097);
nor U14893 (N_14893,N_10481,N_10668);
nor U14894 (N_14894,N_12262,N_12435);
xor U14895 (N_14895,N_11902,N_10698);
or U14896 (N_14896,N_9934,N_9606);
or U14897 (N_14897,N_10156,N_12294);
or U14898 (N_14898,N_12146,N_9877);
or U14899 (N_14899,N_11709,N_10189);
or U14900 (N_14900,N_9776,N_10763);
nor U14901 (N_14901,N_10630,N_10579);
or U14902 (N_14902,N_11080,N_9625);
nand U14903 (N_14903,N_9576,N_10195);
xnor U14904 (N_14904,N_9453,N_9985);
and U14905 (N_14905,N_11714,N_9426);
nor U14906 (N_14906,N_9840,N_10887);
and U14907 (N_14907,N_10735,N_11130);
and U14908 (N_14908,N_10916,N_10471);
nand U14909 (N_14909,N_10580,N_11785);
nand U14910 (N_14910,N_11570,N_9942);
nor U14911 (N_14911,N_11568,N_10269);
and U14912 (N_14912,N_11557,N_11222);
nor U14913 (N_14913,N_12308,N_12043);
or U14914 (N_14914,N_10785,N_11250);
and U14915 (N_14915,N_11347,N_12208);
nand U14916 (N_14916,N_10205,N_11988);
or U14917 (N_14917,N_11453,N_9612);
and U14918 (N_14918,N_11387,N_10235);
xor U14919 (N_14919,N_11212,N_11521);
xor U14920 (N_14920,N_10693,N_9950);
and U14921 (N_14921,N_11888,N_10003);
or U14922 (N_14922,N_9468,N_9981);
and U14923 (N_14923,N_12304,N_9932);
nor U14924 (N_14924,N_11716,N_12074);
and U14925 (N_14925,N_10672,N_9631);
and U14926 (N_14926,N_12361,N_11238);
or U14927 (N_14927,N_9801,N_9706);
nand U14928 (N_14928,N_12288,N_9567);
nor U14929 (N_14929,N_10514,N_12416);
and U14930 (N_14930,N_12440,N_9412);
and U14931 (N_14931,N_11994,N_10076);
nor U14932 (N_14932,N_11720,N_11019);
nand U14933 (N_14933,N_11485,N_11633);
nor U14934 (N_14934,N_10824,N_9506);
and U14935 (N_14935,N_9448,N_11353);
xnor U14936 (N_14936,N_9969,N_11099);
and U14937 (N_14937,N_9874,N_11671);
nor U14938 (N_14938,N_11905,N_10800);
or U14939 (N_14939,N_10204,N_12284);
nor U14940 (N_14940,N_9803,N_11115);
or U14941 (N_14941,N_10322,N_12163);
and U14942 (N_14942,N_12135,N_11742);
or U14943 (N_14943,N_12205,N_12240);
or U14944 (N_14944,N_9461,N_11511);
or U14945 (N_14945,N_10899,N_12380);
and U14946 (N_14946,N_10825,N_10568);
and U14947 (N_14947,N_12483,N_11229);
xor U14948 (N_14948,N_10023,N_11741);
xnor U14949 (N_14949,N_10695,N_11834);
nor U14950 (N_14950,N_12294,N_9524);
and U14951 (N_14951,N_9844,N_10423);
nand U14952 (N_14952,N_9738,N_10574);
and U14953 (N_14953,N_11694,N_10549);
nor U14954 (N_14954,N_10881,N_11322);
nand U14955 (N_14955,N_12441,N_9887);
and U14956 (N_14956,N_11207,N_10665);
xor U14957 (N_14957,N_9636,N_11322);
and U14958 (N_14958,N_11931,N_9397);
nand U14959 (N_14959,N_10698,N_9584);
nor U14960 (N_14960,N_11090,N_10812);
or U14961 (N_14961,N_9781,N_11070);
nand U14962 (N_14962,N_10649,N_11557);
or U14963 (N_14963,N_12447,N_10044);
or U14964 (N_14964,N_10754,N_12252);
nand U14965 (N_14965,N_9898,N_12058);
nor U14966 (N_14966,N_10274,N_11909);
or U14967 (N_14967,N_9839,N_9498);
and U14968 (N_14968,N_10122,N_11880);
or U14969 (N_14969,N_11691,N_9509);
nor U14970 (N_14970,N_11910,N_12061);
or U14971 (N_14971,N_11702,N_9804);
or U14972 (N_14972,N_10166,N_11002);
xor U14973 (N_14973,N_10608,N_10834);
and U14974 (N_14974,N_9613,N_10893);
and U14975 (N_14975,N_11759,N_11062);
nor U14976 (N_14976,N_12412,N_10587);
nand U14977 (N_14977,N_12422,N_9877);
nor U14978 (N_14978,N_10702,N_10292);
nand U14979 (N_14979,N_9504,N_10938);
and U14980 (N_14980,N_11481,N_11469);
nand U14981 (N_14981,N_10960,N_10253);
xor U14982 (N_14982,N_10478,N_11953);
and U14983 (N_14983,N_11174,N_11341);
nor U14984 (N_14984,N_10109,N_11346);
nor U14985 (N_14985,N_9722,N_9939);
and U14986 (N_14986,N_9454,N_10662);
or U14987 (N_14987,N_12304,N_12282);
or U14988 (N_14988,N_10532,N_11107);
nor U14989 (N_14989,N_12358,N_12414);
or U14990 (N_14990,N_11883,N_12300);
nor U14991 (N_14991,N_11950,N_11645);
nand U14992 (N_14992,N_11147,N_11713);
nand U14993 (N_14993,N_11216,N_9934);
nand U14994 (N_14994,N_11450,N_11205);
nor U14995 (N_14995,N_11619,N_10655);
xnor U14996 (N_14996,N_10496,N_11100);
nand U14997 (N_14997,N_9614,N_10392);
nand U14998 (N_14998,N_11825,N_10779);
and U14999 (N_14999,N_10083,N_10149);
and U15000 (N_15000,N_10179,N_10272);
nor U15001 (N_15001,N_9626,N_11197);
nand U15002 (N_15002,N_9729,N_11967);
nor U15003 (N_15003,N_9568,N_10042);
nor U15004 (N_15004,N_10178,N_9932);
and U15005 (N_15005,N_12025,N_9997);
nand U15006 (N_15006,N_9924,N_12123);
nor U15007 (N_15007,N_9866,N_12171);
or U15008 (N_15008,N_10736,N_11646);
nand U15009 (N_15009,N_12020,N_10120);
and U15010 (N_15010,N_10855,N_10896);
and U15011 (N_15011,N_11268,N_11383);
and U15012 (N_15012,N_12213,N_11607);
nand U15013 (N_15013,N_11282,N_11237);
and U15014 (N_15014,N_11978,N_10613);
and U15015 (N_15015,N_10046,N_10789);
nand U15016 (N_15016,N_12497,N_9622);
or U15017 (N_15017,N_9684,N_11656);
nor U15018 (N_15018,N_11566,N_10722);
xor U15019 (N_15019,N_9733,N_10430);
nor U15020 (N_15020,N_11729,N_9787);
and U15021 (N_15021,N_11451,N_11649);
or U15022 (N_15022,N_12447,N_11312);
nor U15023 (N_15023,N_10934,N_9520);
xor U15024 (N_15024,N_10271,N_9959);
and U15025 (N_15025,N_10743,N_9498);
and U15026 (N_15026,N_9670,N_11179);
nor U15027 (N_15027,N_11060,N_10607);
or U15028 (N_15028,N_9899,N_10648);
nor U15029 (N_15029,N_11018,N_10700);
and U15030 (N_15030,N_9937,N_11505);
nand U15031 (N_15031,N_11665,N_10537);
nor U15032 (N_15032,N_10359,N_10797);
nand U15033 (N_15033,N_9481,N_12199);
nor U15034 (N_15034,N_11424,N_12166);
xor U15035 (N_15035,N_12421,N_10600);
and U15036 (N_15036,N_12009,N_11474);
nand U15037 (N_15037,N_10988,N_11636);
nor U15038 (N_15038,N_9750,N_12222);
nor U15039 (N_15039,N_10537,N_11663);
or U15040 (N_15040,N_10530,N_11142);
nor U15041 (N_15041,N_10016,N_10689);
and U15042 (N_15042,N_11097,N_10931);
and U15043 (N_15043,N_11619,N_11337);
and U15044 (N_15044,N_12331,N_11896);
nor U15045 (N_15045,N_11190,N_10452);
or U15046 (N_15046,N_9609,N_11132);
nor U15047 (N_15047,N_12395,N_12426);
and U15048 (N_15048,N_11750,N_10813);
nand U15049 (N_15049,N_11251,N_9995);
nor U15050 (N_15050,N_11048,N_10784);
or U15051 (N_15051,N_11337,N_9938);
nand U15052 (N_15052,N_11861,N_9672);
nor U15053 (N_15053,N_10992,N_11106);
or U15054 (N_15054,N_10204,N_10793);
or U15055 (N_15055,N_9987,N_9725);
nand U15056 (N_15056,N_10789,N_12308);
and U15057 (N_15057,N_9509,N_12017);
nand U15058 (N_15058,N_11839,N_11971);
nand U15059 (N_15059,N_9547,N_11463);
or U15060 (N_15060,N_11512,N_10176);
nand U15061 (N_15061,N_10483,N_12369);
nor U15062 (N_15062,N_11375,N_11508);
nand U15063 (N_15063,N_10827,N_10409);
nor U15064 (N_15064,N_9400,N_11629);
xor U15065 (N_15065,N_10949,N_9743);
or U15066 (N_15066,N_12424,N_10276);
nand U15067 (N_15067,N_9723,N_11226);
and U15068 (N_15068,N_11700,N_10789);
nor U15069 (N_15069,N_11215,N_10352);
and U15070 (N_15070,N_10106,N_12274);
nor U15071 (N_15071,N_12141,N_11441);
xor U15072 (N_15072,N_12445,N_9893);
nand U15073 (N_15073,N_12124,N_9442);
nand U15074 (N_15074,N_11488,N_9684);
nand U15075 (N_15075,N_10591,N_12027);
xor U15076 (N_15076,N_11625,N_10849);
and U15077 (N_15077,N_10142,N_10687);
or U15078 (N_15078,N_11353,N_10570);
or U15079 (N_15079,N_11036,N_10975);
or U15080 (N_15080,N_11580,N_10036);
nand U15081 (N_15081,N_12071,N_9504);
xnor U15082 (N_15082,N_11868,N_10853);
nand U15083 (N_15083,N_10936,N_10424);
and U15084 (N_15084,N_12265,N_12224);
nand U15085 (N_15085,N_10851,N_11373);
and U15086 (N_15086,N_10255,N_11718);
and U15087 (N_15087,N_9888,N_9622);
and U15088 (N_15088,N_12493,N_12020);
nand U15089 (N_15089,N_10817,N_10853);
or U15090 (N_15090,N_12371,N_10910);
nand U15091 (N_15091,N_9926,N_11884);
xnor U15092 (N_15092,N_11283,N_12489);
nand U15093 (N_15093,N_12096,N_11618);
nor U15094 (N_15094,N_12116,N_10342);
xor U15095 (N_15095,N_12453,N_10867);
or U15096 (N_15096,N_9435,N_10597);
and U15097 (N_15097,N_9665,N_11862);
or U15098 (N_15098,N_10139,N_11159);
nor U15099 (N_15099,N_11048,N_12118);
nor U15100 (N_15100,N_10032,N_12243);
nand U15101 (N_15101,N_11259,N_11564);
nor U15102 (N_15102,N_11235,N_10107);
nor U15103 (N_15103,N_11222,N_12468);
nor U15104 (N_15104,N_10826,N_12203);
nor U15105 (N_15105,N_11680,N_10586);
xnor U15106 (N_15106,N_12035,N_12342);
xnor U15107 (N_15107,N_11748,N_12307);
and U15108 (N_15108,N_9821,N_10567);
and U15109 (N_15109,N_12085,N_10644);
nor U15110 (N_15110,N_10738,N_9594);
nand U15111 (N_15111,N_11095,N_9960);
nor U15112 (N_15112,N_11053,N_9476);
xnor U15113 (N_15113,N_10464,N_11533);
nor U15114 (N_15114,N_12408,N_9622);
or U15115 (N_15115,N_9412,N_11318);
and U15116 (N_15116,N_11856,N_10960);
nor U15117 (N_15117,N_12446,N_11760);
nor U15118 (N_15118,N_11524,N_9498);
nand U15119 (N_15119,N_10332,N_9935);
xnor U15120 (N_15120,N_9769,N_10339);
nor U15121 (N_15121,N_12014,N_11312);
nand U15122 (N_15122,N_11437,N_10160);
xor U15123 (N_15123,N_10641,N_11177);
xnor U15124 (N_15124,N_9453,N_11835);
or U15125 (N_15125,N_12408,N_12241);
nor U15126 (N_15126,N_11837,N_10361);
nor U15127 (N_15127,N_10783,N_10366);
nor U15128 (N_15128,N_10021,N_10432);
and U15129 (N_15129,N_10174,N_10393);
nor U15130 (N_15130,N_9907,N_12196);
or U15131 (N_15131,N_11371,N_11019);
and U15132 (N_15132,N_11501,N_9568);
nand U15133 (N_15133,N_10650,N_10900);
and U15134 (N_15134,N_10737,N_12135);
or U15135 (N_15135,N_11266,N_10553);
nand U15136 (N_15136,N_11617,N_12217);
xnor U15137 (N_15137,N_10835,N_11716);
xnor U15138 (N_15138,N_11398,N_11916);
or U15139 (N_15139,N_10267,N_11985);
and U15140 (N_15140,N_11062,N_10429);
nor U15141 (N_15141,N_9644,N_12045);
or U15142 (N_15142,N_9943,N_10119);
and U15143 (N_15143,N_11751,N_12169);
nand U15144 (N_15144,N_9543,N_11230);
nand U15145 (N_15145,N_10717,N_11480);
and U15146 (N_15146,N_11846,N_11757);
nand U15147 (N_15147,N_10950,N_12066);
nor U15148 (N_15148,N_11088,N_10504);
and U15149 (N_15149,N_10688,N_9829);
and U15150 (N_15150,N_10570,N_10235);
and U15151 (N_15151,N_9662,N_10783);
or U15152 (N_15152,N_12132,N_12329);
nand U15153 (N_15153,N_10912,N_9802);
nor U15154 (N_15154,N_10839,N_11042);
or U15155 (N_15155,N_11897,N_11492);
nor U15156 (N_15156,N_12420,N_11141);
xor U15157 (N_15157,N_12320,N_11024);
and U15158 (N_15158,N_9872,N_10894);
nand U15159 (N_15159,N_12054,N_9706);
xnor U15160 (N_15160,N_12491,N_11942);
and U15161 (N_15161,N_12457,N_11064);
nor U15162 (N_15162,N_11286,N_12151);
and U15163 (N_15163,N_9721,N_11381);
nand U15164 (N_15164,N_9503,N_12275);
or U15165 (N_15165,N_10202,N_11361);
nor U15166 (N_15166,N_10242,N_9619);
nor U15167 (N_15167,N_10791,N_9496);
nor U15168 (N_15168,N_9828,N_10872);
nor U15169 (N_15169,N_9653,N_12093);
xnor U15170 (N_15170,N_10061,N_9530);
nor U15171 (N_15171,N_11456,N_12286);
or U15172 (N_15172,N_11931,N_11388);
nand U15173 (N_15173,N_12281,N_9717);
nand U15174 (N_15174,N_11060,N_9494);
nor U15175 (N_15175,N_10880,N_11263);
nand U15176 (N_15176,N_12092,N_11531);
nor U15177 (N_15177,N_12470,N_11545);
nand U15178 (N_15178,N_10251,N_10606);
and U15179 (N_15179,N_12037,N_10222);
nor U15180 (N_15180,N_12202,N_9510);
or U15181 (N_15181,N_9879,N_10051);
or U15182 (N_15182,N_9891,N_11762);
and U15183 (N_15183,N_9782,N_9755);
and U15184 (N_15184,N_11527,N_9546);
xor U15185 (N_15185,N_9516,N_12261);
xnor U15186 (N_15186,N_10675,N_12215);
xnor U15187 (N_15187,N_11613,N_10695);
xnor U15188 (N_15188,N_11923,N_12037);
and U15189 (N_15189,N_10622,N_10337);
and U15190 (N_15190,N_10616,N_10421);
and U15191 (N_15191,N_9585,N_12350);
or U15192 (N_15192,N_9768,N_10930);
or U15193 (N_15193,N_12213,N_10717);
and U15194 (N_15194,N_10307,N_12302);
nand U15195 (N_15195,N_9890,N_11282);
nand U15196 (N_15196,N_11075,N_12428);
nand U15197 (N_15197,N_11655,N_12451);
and U15198 (N_15198,N_11482,N_9823);
and U15199 (N_15199,N_11632,N_9567);
nor U15200 (N_15200,N_11906,N_10442);
and U15201 (N_15201,N_9807,N_9480);
and U15202 (N_15202,N_11213,N_11649);
nand U15203 (N_15203,N_10518,N_10335);
and U15204 (N_15204,N_11055,N_11429);
and U15205 (N_15205,N_12223,N_11284);
and U15206 (N_15206,N_10437,N_9536);
and U15207 (N_15207,N_11500,N_10006);
and U15208 (N_15208,N_12039,N_12135);
and U15209 (N_15209,N_11366,N_10691);
or U15210 (N_15210,N_12039,N_11479);
and U15211 (N_15211,N_9621,N_12299);
or U15212 (N_15212,N_10836,N_10587);
or U15213 (N_15213,N_9442,N_11693);
or U15214 (N_15214,N_10616,N_10765);
xnor U15215 (N_15215,N_10865,N_10146);
nand U15216 (N_15216,N_10782,N_10596);
or U15217 (N_15217,N_9624,N_10098);
or U15218 (N_15218,N_10174,N_10436);
nor U15219 (N_15219,N_11241,N_9545);
nand U15220 (N_15220,N_9973,N_10456);
nand U15221 (N_15221,N_11990,N_11667);
nand U15222 (N_15222,N_9993,N_12467);
and U15223 (N_15223,N_11857,N_11200);
or U15224 (N_15224,N_10952,N_9603);
nand U15225 (N_15225,N_12217,N_10717);
and U15226 (N_15226,N_12186,N_10915);
nor U15227 (N_15227,N_11743,N_10339);
or U15228 (N_15228,N_10822,N_10709);
and U15229 (N_15229,N_11510,N_11757);
or U15230 (N_15230,N_11760,N_11676);
nor U15231 (N_15231,N_12105,N_11983);
nand U15232 (N_15232,N_11784,N_12473);
and U15233 (N_15233,N_11077,N_12146);
nand U15234 (N_15234,N_10953,N_11589);
nand U15235 (N_15235,N_11533,N_10692);
and U15236 (N_15236,N_12262,N_11387);
nand U15237 (N_15237,N_10379,N_11681);
nand U15238 (N_15238,N_11198,N_10121);
nand U15239 (N_15239,N_10110,N_11139);
or U15240 (N_15240,N_11030,N_9945);
nand U15241 (N_15241,N_11394,N_9411);
nor U15242 (N_15242,N_12240,N_9676);
nor U15243 (N_15243,N_10530,N_11576);
nor U15244 (N_15244,N_9709,N_9385);
or U15245 (N_15245,N_9634,N_12448);
nor U15246 (N_15246,N_11739,N_12266);
or U15247 (N_15247,N_11116,N_11818);
and U15248 (N_15248,N_12031,N_11601);
nand U15249 (N_15249,N_11441,N_10945);
and U15250 (N_15250,N_10726,N_10356);
or U15251 (N_15251,N_9577,N_11089);
nor U15252 (N_15252,N_11616,N_12241);
or U15253 (N_15253,N_11698,N_9486);
and U15254 (N_15254,N_12270,N_10261);
nor U15255 (N_15255,N_11211,N_9867);
nor U15256 (N_15256,N_11416,N_11223);
and U15257 (N_15257,N_9469,N_10531);
nor U15258 (N_15258,N_11704,N_11306);
nor U15259 (N_15259,N_12248,N_11759);
nor U15260 (N_15260,N_11944,N_10586);
nor U15261 (N_15261,N_10662,N_9499);
or U15262 (N_15262,N_11508,N_11722);
nand U15263 (N_15263,N_11581,N_10581);
nand U15264 (N_15264,N_11757,N_9928);
nand U15265 (N_15265,N_11948,N_9493);
nor U15266 (N_15266,N_10349,N_10134);
and U15267 (N_15267,N_9969,N_10190);
and U15268 (N_15268,N_12046,N_12045);
and U15269 (N_15269,N_10184,N_11129);
nand U15270 (N_15270,N_11779,N_10249);
and U15271 (N_15271,N_10200,N_12439);
and U15272 (N_15272,N_10691,N_9674);
or U15273 (N_15273,N_11768,N_10917);
xnor U15274 (N_15274,N_12069,N_10399);
xnor U15275 (N_15275,N_9399,N_12444);
xnor U15276 (N_15276,N_11290,N_9683);
or U15277 (N_15277,N_10862,N_11482);
and U15278 (N_15278,N_10629,N_11482);
nor U15279 (N_15279,N_9476,N_10431);
nor U15280 (N_15280,N_9988,N_11777);
nor U15281 (N_15281,N_10630,N_10798);
nor U15282 (N_15282,N_12326,N_11924);
xnor U15283 (N_15283,N_9729,N_11960);
or U15284 (N_15284,N_11035,N_11963);
nor U15285 (N_15285,N_10187,N_11115);
or U15286 (N_15286,N_10106,N_9889);
and U15287 (N_15287,N_11005,N_9959);
and U15288 (N_15288,N_10609,N_10847);
nand U15289 (N_15289,N_12465,N_9389);
nand U15290 (N_15290,N_10351,N_11743);
nand U15291 (N_15291,N_10483,N_10216);
nor U15292 (N_15292,N_9896,N_10123);
and U15293 (N_15293,N_10062,N_9413);
or U15294 (N_15294,N_9502,N_11401);
or U15295 (N_15295,N_10863,N_12453);
and U15296 (N_15296,N_11462,N_10232);
and U15297 (N_15297,N_9498,N_10332);
nand U15298 (N_15298,N_11091,N_10280);
and U15299 (N_15299,N_12002,N_11181);
nand U15300 (N_15300,N_11248,N_11773);
or U15301 (N_15301,N_11590,N_9746);
nor U15302 (N_15302,N_11489,N_10863);
xnor U15303 (N_15303,N_11538,N_11336);
or U15304 (N_15304,N_11139,N_11204);
nand U15305 (N_15305,N_10307,N_9770);
and U15306 (N_15306,N_12250,N_10202);
or U15307 (N_15307,N_10953,N_9698);
or U15308 (N_15308,N_10676,N_12290);
nor U15309 (N_15309,N_10170,N_10993);
nor U15310 (N_15310,N_10123,N_12393);
nand U15311 (N_15311,N_9918,N_11402);
nor U15312 (N_15312,N_9376,N_10459);
and U15313 (N_15313,N_10190,N_12122);
nor U15314 (N_15314,N_10487,N_11962);
nor U15315 (N_15315,N_11657,N_12353);
nor U15316 (N_15316,N_10479,N_10243);
nand U15317 (N_15317,N_11154,N_12109);
or U15318 (N_15318,N_10716,N_10000);
or U15319 (N_15319,N_10560,N_11442);
nand U15320 (N_15320,N_9718,N_12236);
xor U15321 (N_15321,N_11049,N_11537);
nand U15322 (N_15322,N_10505,N_10347);
nand U15323 (N_15323,N_10884,N_11087);
or U15324 (N_15324,N_11732,N_12070);
nor U15325 (N_15325,N_11934,N_9943);
or U15326 (N_15326,N_10635,N_9434);
nand U15327 (N_15327,N_11711,N_9874);
or U15328 (N_15328,N_11268,N_11214);
nand U15329 (N_15329,N_10444,N_11704);
or U15330 (N_15330,N_10060,N_9425);
nor U15331 (N_15331,N_9728,N_12063);
and U15332 (N_15332,N_9976,N_11705);
and U15333 (N_15333,N_10542,N_10381);
and U15334 (N_15334,N_10040,N_11058);
or U15335 (N_15335,N_10266,N_12283);
nand U15336 (N_15336,N_11647,N_10273);
xnor U15337 (N_15337,N_11954,N_10247);
nand U15338 (N_15338,N_10216,N_12427);
xnor U15339 (N_15339,N_9552,N_10296);
and U15340 (N_15340,N_11816,N_9746);
or U15341 (N_15341,N_10937,N_9636);
and U15342 (N_15342,N_12420,N_10138);
nor U15343 (N_15343,N_12310,N_10489);
nor U15344 (N_15344,N_10896,N_11474);
or U15345 (N_15345,N_11319,N_11140);
and U15346 (N_15346,N_9905,N_10672);
and U15347 (N_15347,N_11795,N_9602);
nor U15348 (N_15348,N_11666,N_12360);
nor U15349 (N_15349,N_10772,N_9814);
and U15350 (N_15350,N_11775,N_11755);
nand U15351 (N_15351,N_11224,N_9962);
and U15352 (N_15352,N_9526,N_10015);
nor U15353 (N_15353,N_12339,N_12492);
nand U15354 (N_15354,N_9435,N_9758);
or U15355 (N_15355,N_9666,N_12482);
nor U15356 (N_15356,N_10897,N_11733);
and U15357 (N_15357,N_11438,N_10093);
and U15358 (N_15358,N_11640,N_10833);
and U15359 (N_15359,N_12485,N_11041);
nand U15360 (N_15360,N_11538,N_11058);
nand U15361 (N_15361,N_11847,N_11082);
and U15362 (N_15362,N_9940,N_10742);
nand U15363 (N_15363,N_9625,N_9749);
and U15364 (N_15364,N_11213,N_10005);
nand U15365 (N_15365,N_10683,N_11950);
and U15366 (N_15366,N_11460,N_12479);
or U15367 (N_15367,N_9670,N_11907);
nor U15368 (N_15368,N_10192,N_11469);
and U15369 (N_15369,N_11818,N_9726);
nor U15370 (N_15370,N_11420,N_9985);
nor U15371 (N_15371,N_12377,N_12141);
nor U15372 (N_15372,N_12440,N_9743);
or U15373 (N_15373,N_12077,N_11361);
or U15374 (N_15374,N_10551,N_11061);
and U15375 (N_15375,N_9716,N_9463);
or U15376 (N_15376,N_10671,N_10093);
nand U15377 (N_15377,N_11393,N_10309);
xnor U15378 (N_15378,N_11354,N_10702);
or U15379 (N_15379,N_12059,N_12225);
nor U15380 (N_15380,N_10900,N_9382);
nand U15381 (N_15381,N_12115,N_10264);
and U15382 (N_15382,N_11103,N_11876);
nor U15383 (N_15383,N_9788,N_11045);
and U15384 (N_15384,N_12315,N_10829);
and U15385 (N_15385,N_10212,N_12133);
nand U15386 (N_15386,N_11951,N_10905);
nand U15387 (N_15387,N_9506,N_10071);
nor U15388 (N_15388,N_10866,N_10580);
and U15389 (N_15389,N_11183,N_11610);
and U15390 (N_15390,N_9923,N_9752);
nand U15391 (N_15391,N_12467,N_11030);
and U15392 (N_15392,N_11654,N_11586);
and U15393 (N_15393,N_12199,N_10895);
xor U15394 (N_15394,N_12369,N_12305);
or U15395 (N_15395,N_9782,N_10248);
and U15396 (N_15396,N_10095,N_11846);
xnor U15397 (N_15397,N_9886,N_12232);
nor U15398 (N_15398,N_11514,N_9832);
nand U15399 (N_15399,N_11076,N_10253);
xnor U15400 (N_15400,N_11372,N_11009);
or U15401 (N_15401,N_10200,N_12394);
nor U15402 (N_15402,N_12207,N_11091);
or U15403 (N_15403,N_10758,N_11451);
nand U15404 (N_15404,N_10746,N_11063);
or U15405 (N_15405,N_10169,N_10825);
nor U15406 (N_15406,N_11149,N_11954);
nand U15407 (N_15407,N_10969,N_10930);
xor U15408 (N_15408,N_9468,N_11041);
xor U15409 (N_15409,N_11249,N_12093);
nor U15410 (N_15410,N_11262,N_10005);
nand U15411 (N_15411,N_9565,N_9870);
and U15412 (N_15412,N_10892,N_11641);
nor U15413 (N_15413,N_12218,N_10456);
xor U15414 (N_15414,N_11980,N_11599);
nor U15415 (N_15415,N_11508,N_12331);
and U15416 (N_15416,N_10333,N_12081);
or U15417 (N_15417,N_10783,N_10761);
and U15418 (N_15418,N_10528,N_11306);
nor U15419 (N_15419,N_9393,N_10906);
and U15420 (N_15420,N_11728,N_9823);
and U15421 (N_15421,N_11152,N_11463);
xor U15422 (N_15422,N_11377,N_9762);
nand U15423 (N_15423,N_11519,N_10765);
or U15424 (N_15424,N_12485,N_9955);
nor U15425 (N_15425,N_12050,N_9475);
and U15426 (N_15426,N_10541,N_9580);
and U15427 (N_15427,N_11642,N_10247);
nor U15428 (N_15428,N_10627,N_11569);
nand U15429 (N_15429,N_11625,N_9377);
or U15430 (N_15430,N_9573,N_11529);
or U15431 (N_15431,N_9963,N_10945);
nor U15432 (N_15432,N_12293,N_10708);
nor U15433 (N_15433,N_11661,N_11515);
nand U15434 (N_15434,N_12306,N_11576);
or U15435 (N_15435,N_12043,N_12136);
or U15436 (N_15436,N_10617,N_10541);
nor U15437 (N_15437,N_9626,N_11580);
nand U15438 (N_15438,N_11661,N_11357);
nor U15439 (N_15439,N_11394,N_11282);
nand U15440 (N_15440,N_9869,N_10203);
nand U15441 (N_15441,N_9403,N_11087);
nand U15442 (N_15442,N_10858,N_11038);
or U15443 (N_15443,N_10492,N_11889);
or U15444 (N_15444,N_9563,N_10582);
nor U15445 (N_15445,N_10283,N_10469);
and U15446 (N_15446,N_11265,N_11006);
nand U15447 (N_15447,N_10580,N_11435);
and U15448 (N_15448,N_10272,N_10871);
nor U15449 (N_15449,N_11663,N_11312);
and U15450 (N_15450,N_10965,N_10422);
or U15451 (N_15451,N_11253,N_11700);
or U15452 (N_15452,N_10817,N_10419);
nand U15453 (N_15453,N_11594,N_11221);
and U15454 (N_15454,N_10751,N_12223);
xor U15455 (N_15455,N_9463,N_11298);
xor U15456 (N_15456,N_10135,N_12206);
xor U15457 (N_15457,N_12303,N_12167);
and U15458 (N_15458,N_11114,N_10699);
xor U15459 (N_15459,N_9622,N_10944);
and U15460 (N_15460,N_9606,N_11714);
and U15461 (N_15461,N_9863,N_9488);
nand U15462 (N_15462,N_9995,N_9720);
nand U15463 (N_15463,N_11823,N_10246);
nand U15464 (N_15464,N_12229,N_9997);
nand U15465 (N_15465,N_10781,N_10504);
or U15466 (N_15466,N_11069,N_12077);
nor U15467 (N_15467,N_10836,N_11132);
nand U15468 (N_15468,N_10083,N_11634);
or U15469 (N_15469,N_12273,N_10792);
or U15470 (N_15470,N_9804,N_11824);
and U15471 (N_15471,N_9889,N_11647);
nor U15472 (N_15472,N_11360,N_11182);
xnor U15473 (N_15473,N_12223,N_11144);
xor U15474 (N_15474,N_11542,N_9572);
or U15475 (N_15475,N_12059,N_10626);
nor U15476 (N_15476,N_12007,N_10935);
nor U15477 (N_15477,N_10734,N_12164);
nand U15478 (N_15478,N_11318,N_11571);
xnor U15479 (N_15479,N_12310,N_10460);
and U15480 (N_15480,N_10285,N_10517);
or U15481 (N_15481,N_10826,N_12214);
nor U15482 (N_15482,N_10618,N_11903);
or U15483 (N_15483,N_11017,N_11656);
and U15484 (N_15484,N_10084,N_11483);
nand U15485 (N_15485,N_10615,N_10357);
or U15486 (N_15486,N_10928,N_10755);
nand U15487 (N_15487,N_11113,N_11202);
or U15488 (N_15488,N_10965,N_10944);
nand U15489 (N_15489,N_11798,N_11638);
nand U15490 (N_15490,N_12142,N_10837);
nand U15491 (N_15491,N_12021,N_11338);
and U15492 (N_15492,N_12055,N_9526);
nand U15493 (N_15493,N_12317,N_11746);
nand U15494 (N_15494,N_12380,N_9917);
nor U15495 (N_15495,N_11042,N_10536);
xor U15496 (N_15496,N_9710,N_9511);
nor U15497 (N_15497,N_9862,N_10552);
and U15498 (N_15498,N_10652,N_10584);
nor U15499 (N_15499,N_10664,N_12106);
nand U15500 (N_15500,N_9735,N_10965);
nor U15501 (N_15501,N_9869,N_11556);
nand U15502 (N_15502,N_12093,N_12217);
or U15503 (N_15503,N_9625,N_11458);
or U15504 (N_15504,N_12360,N_11797);
nor U15505 (N_15505,N_10488,N_9666);
nand U15506 (N_15506,N_12119,N_9932);
nand U15507 (N_15507,N_11183,N_11889);
nor U15508 (N_15508,N_11445,N_9580);
or U15509 (N_15509,N_10597,N_12111);
or U15510 (N_15510,N_12429,N_10702);
or U15511 (N_15511,N_10065,N_10227);
or U15512 (N_15512,N_11754,N_11671);
xor U15513 (N_15513,N_10569,N_11829);
or U15514 (N_15514,N_11292,N_9534);
nor U15515 (N_15515,N_10083,N_12118);
or U15516 (N_15516,N_11519,N_10696);
and U15517 (N_15517,N_9869,N_11791);
and U15518 (N_15518,N_11880,N_10974);
or U15519 (N_15519,N_12137,N_9715);
nor U15520 (N_15520,N_11499,N_9537);
and U15521 (N_15521,N_9562,N_9887);
nand U15522 (N_15522,N_11754,N_10133);
nand U15523 (N_15523,N_12287,N_10799);
or U15524 (N_15524,N_11404,N_10737);
and U15525 (N_15525,N_11265,N_10212);
nand U15526 (N_15526,N_9503,N_9420);
and U15527 (N_15527,N_10887,N_11306);
and U15528 (N_15528,N_10550,N_11593);
nand U15529 (N_15529,N_11216,N_10889);
xnor U15530 (N_15530,N_9788,N_11478);
nand U15531 (N_15531,N_10073,N_12053);
and U15532 (N_15532,N_10792,N_9927);
nand U15533 (N_15533,N_12096,N_11603);
or U15534 (N_15534,N_10971,N_12369);
xnor U15535 (N_15535,N_11696,N_11036);
nor U15536 (N_15536,N_12133,N_12186);
nand U15537 (N_15537,N_10253,N_12270);
nor U15538 (N_15538,N_10628,N_10820);
xnor U15539 (N_15539,N_11623,N_11126);
nand U15540 (N_15540,N_10143,N_10572);
nand U15541 (N_15541,N_11953,N_10813);
or U15542 (N_15542,N_10170,N_10291);
xnor U15543 (N_15543,N_9408,N_10497);
and U15544 (N_15544,N_10210,N_11902);
or U15545 (N_15545,N_12071,N_10108);
nor U15546 (N_15546,N_10961,N_10411);
nand U15547 (N_15547,N_12203,N_11496);
nor U15548 (N_15548,N_11561,N_11545);
and U15549 (N_15549,N_10856,N_11197);
or U15550 (N_15550,N_11381,N_10154);
xor U15551 (N_15551,N_9410,N_10328);
nor U15552 (N_15552,N_11561,N_11568);
nand U15553 (N_15553,N_11463,N_11311);
or U15554 (N_15554,N_9594,N_10381);
nand U15555 (N_15555,N_11179,N_11898);
nor U15556 (N_15556,N_9821,N_12126);
nor U15557 (N_15557,N_11956,N_12051);
nand U15558 (N_15558,N_10424,N_9869);
or U15559 (N_15559,N_10755,N_12487);
nor U15560 (N_15560,N_11931,N_9585);
nor U15561 (N_15561,N_11242,N_9379);
or U15562 (N_15562,N_11947,N_10384);
and U15563 (N_15563,N_9612,N_12251);
and U15564 (N_15564,N_11359,N_10187);
or U15565 (N_15565,N_9864,N_10127);
xnor U15566 (N_15566,N_9853,N_10765);
nor U15567 (N_15567,N_11128,N_9426);
or U15568 (N_15568,N_11592,N_11829);
and U15569 (N_15569,N_12249,N_11609);
xor U15570 (N_15570,N_10345,N_11647);
nand U15571 (N_15571,N_11340,N_9997);
nor U15572 (N_15572,N_10759,N_10376);
nor U15573 (N_15573,N_10599,N_11293);
xnor U15574 (N_15574,N_11883,N_9766);
and U15575 (N_15575,N_9846,N_12411);
nor U15576 (N_15576,N_12366,N_11848);
nor U15577 (N_15577,N_10310,N_10041);
or U15578 (N_15578,N_10057,N_9425);
xnor U15579 (N_15579,N_12338,N_9575);
and U15580 (N_15580,N_9579,N_11889);
xnor U15581 (N_15581,N_9597,N_11677);
xor U15582 (N_15582,N_11136,N_11124);
nor U15583 (N_15583,N_11945,N_11704);
nand U15584 (N_15584,N_11415,N_10116);
and U15585 (N_15585,N_9605,N_10158);
or U15586 (N_15586,N_12470,N_10284);
xor U15587 (N_15587,N_12138,N_10261);
nor U15588 (N_15588,N_12069,N_10416);
nand U15589 (N_15589,N_10079,N_11162);
xnor U15590 (N_15590,N_9835,N_10572);
or U15591 (N_15591,N_9399,N_10109);
nand U15592 (N_15592,N_11690,N_11327);
nor U15593 (N_15593,N_10136,N_11161);
nor U15594 (N_15594,N_11474,N_12067);
or U15595 (N_15595,N_10489,N_11664);
nor U15596 (N_15596,N_10528,N_11646);
nand U15597 (N_15597,N_11915,N_11751);
or U15598 (N_15598,N_9526,N_10084);
nand U15599 (N_15599,N_11307,N_9645);
xor U15600 (N_15600,N_9451,N_11863);
nor U15601 (N_15601,N_10922,N_9995);
and U15602 (N_15602,N_9869,N_11376);
xor U15603 (N_15603,N_10064,N_10016);
and U15604 (N_15604,N_11632,N_12302);
and U15605 (N_15605,N_10919,N_10008);
nor U15606 (N_15606,N_11034,N_11754);
nor U15607 (N_15607,N_10219,N_12441);
nor U15608 (N_15608,N_12083,N_10825);
or U15609 (N_15609,N_9459,N_11682);
or U15610 (N_15610,N_10275,N_10416);
nand U15611 (N_15611,N_12193,N_9774);
or U15612 (N_15612,N_10295,N_10159);
nand U15613 (N_15613,N_10265,N_12359);
xor U15614 (N_15614,N_10624,N_9601);
xnor U15615 (N_15615,N_10252,N_9520);
or U15616 (N_15616,N_12270,N_10815);
or U15617 (N_15617,N_9945,N_9927);
and U15618 (N_15618,N_10087,N_11981);
nor U15619 (N_15619,N_12051,N_12386);
and U15620 (N_15620,N_10406,N_10915);
nand U15621 (N_15621,N_11343,N_10171);
or U15622 (N_15622,N_11795,N_12293);
and U15623 (N_15623,N_9721,N_11052);
nand U15624 (N_15624,N_9725,N_11733);
or U15625 (N_15625,N_13926,N_13937);
and U15626 (N_15626,N_13619,N_13305);
nand U15627 (N_15627,N_13229,N_13100);
and U15628 (N_15628,N_15282,N_12917);
nand U15629 (N_15629,N_14116,N_15201);
nor U15630 (N_15630,N_15147,N_14861);
and U15631 (N_15631,N_12553,N_12713);
and U15632 (N_15632,N_15474,N_13717);
and U15633 (N_15633,N_12981,N_14311);
nor U15634 (N_15634,N_15013,N_12655);
nand U15635 (N_15635,N_14415,N_15274);
xor U15636 (N_15636,N_14409,N_15601);
xor U15637 (N_15637,N_14993,N_13047);
xnor U15638 (N_15638,N_14045,N_14199);
and U15639 (N_15639,N_15249,N_12963);
or U15640 (N_15640,N_12872,N_14060);
nand U15641 (N_15641,N_15310,N_13409);
nor U15642 (N_15642,N_14112,N_13623);
nor U15643 (N_15643,N_14516,N_14456);
and U15644 (N_15644,N_13613,N_13219);
nor U15645 (N_15645,N_13133,N_12833);
nor U15646 (N_15646,N_13686,N_14690);
nand U15647 (N_15647,N_14169,N_14617);
and U15648 (N_15648,N_13343,N_15146);
and U15649 (N_15649,N_14852,N_14417);
or U15650 (N_15650,N_15520,N_14575);
xnor U15651 (N_15651,N_13429,N_15382);
and U15652 (N_15652,N_15069,N_13073);
or U15653 (N_15653,N_14623,N_15402);
and U15654 (N_15654,N_13145,N_15361);
and U15655 (N_15655,N_14356,N_14096);
nand U15656 (N_15656,N_14384,N_14020);
and U15657 (N_15657,N_12686,N_14142);
and U15658 (N_15658,N_14372,N_12716);
or U15659 (N_15659,N_12809,N_13199);
and U15660 (N_15660,N_14909,N_14598);
nor U15661 (N_15661,N_14192,N_12783);
xor U15662 (N_15662,N_15546,N_13163);
and U15663 (N_15663,N_12982,N_13706);
and U15664 (N_15664,N_12871,N_13584);
nor U15665 (N_15665,N_13443,N_15371);
nor U15666 (N_15666,N_15124,N_15059);
nor U15667 (N_15667,N_12508,N_13468);
nand U15668 (N_15668,N_13304,N_12988);
or U15669 (N_15669,N_14407,N_13827);
or U15670 (N_15670,N_13460,N_12543);
and U15671 (N_15671,N_14362,N_13854);
nor U15672 (N_15672,N_14021,N_15264);
nor U15673 (N_15673,N_13770,N_13734);
or U15674 (N_15674,N_14803,N_15503);
or U15675 (N_15675,N_13867,N_14237);
and U15676 (N_15676,N_14238,N_12885);
and U15677 (N_15677,N_13215,N_15624);
nand U15678 (N_15678,N_13297,N_12693);
xor U15679 (N_15679,N_14405,N_12751);
and U15680 (N_15680,N_13438,N_13766);
and U15681 (N_15681,N_14500,N_15522);
nor U15682 (N_15682,N_12940,N_14908);
xor U15683 (N_15683,N_14161,N_15394);
nor U15684 (N_15684,N_15058,N_14596);
nand U15685 (N_15685,N_14485,N_14375);
nand U15686 (N_15686,N_14581,N_15528);
or U15687 (N_15687,N_12594,N_14642);
and U15688 (N_15688,N_13490,N_15428);
xnor U15689 (N_15689,N_13108,N_13467);
nand U15690 (N_15690,N_13448,N_14501);
nand U15691 (N_15691,N_15134,N_14432);
and U15692 (N_15692,N_14184,N_13319);
and U15693 (N_15693,N_12608,N_13576);
and U15694 (N_15694,N_15262,N_13189);
and U15695 (N_15695,N_13381,N_13990);
or U15696 (N_15696,N_12670,N_14573);
or U15697 (N_15697,N_14895,N_13124);
nor U15698 (N_15698,N_15043,N_13664);
or U15699 (N_15699,N_15063,N_15468);
nand U15700 (N_15700,N_13037,N_12818);
nand U15701 (N_15701,N_15494,N_13682);
or U15702 (N_15702,N_13066,N_12763);
nand U15703 (N_15703,N_14555,N_14350);
nand U15704 (N_15704,N_13668,N_12630);
nor U15705 (N_15705,N_15238,N_14657);
xor U15706 (N_15706,N_14484,N_13691);
or U15707 (N_15707,N_12537,N_14232);
nand U15708 (N_15708,N_15560,N_14549);
or U15709 (N_15709,N_12626,N_13228);
or U15710 (N_15710,N_14593,N_13893);
nor U15711 (N_15711,N_15595,N_14578);
and U15712 (N_15712,N_15006,N_13555);
xnor U15713 (N_15713,N_15539,N_14980);
and U15714 (N_15714,N_13981,N_14547);
nor U15715 (N_15715,N_15532,N_14208);
or U15716 (N_15716,N_14209,N_12647);
or U15717 (N_15717,N_15159,N_13747);
and U15718 (N_15718,N_14807,N_14651);
xor U15719 (N_15719,N_13337,N_13850);
nor U15720 (N_15720,N_15442,N_13362);
and U15721 (N_15721,N_15504,N_15187);
nor U15722 (N_15722,N_14509,N_14014);
nor U15723 (N_15723,N_14486,N_12549);
and U15724 (N_15724,N_13900,N_15161);
nor U15725 (N_15725,N_13978,N_15047);
and U15726 (N_15726,N_13763,N_13147);
or U15727 (N_15727,N_13864,N_12855);
nor U15728 (N_15728,N_13670,N_13294);
or U15729 (N_15729,N_13692,N_15505);
and U15730 (N_15730,N_14393,N_13107);
or U15731 (N_15731,N_13431,N_12867);
and U15732 (N_15732,N_14505,N_12683);
or U15733 (N_15733,N_13223,N_12901);
or U15734 (N_15734,N_13799,N_15457);
nand U15735 (N_15735,N_12789,N_14317);
and U15736 (N_15736,N_14524,N_12910);
and U15737 (N_15737,N_14172,N_15220);
nand U15738 (N_15738,N_13702,N_15436);
and U15739 (N_15739,N_15343,N_15455);
and U15740 (N_15740,N_12709,N_14226);
or U15741 (N_15741,N_13502,N_14977);
nor U15742 (N_15742,N_14273,N_14211);
and U15743 (N_15743,N_12842,N_15353);
or U15744 (N_15744,N_14214,N_14247);
or U15745 (N_15745,N_13583,N_13793);
or U15746 (N_15746,N_13602,N_13835);
or U15747 (N_15747,N_14075,N_15111);
xor U15748 (N_15748,N_14278,N_13138);
nand U15749 (N_15749,N_14042,N_12820);
nor U15750 (N_15750,N_14202,N_14864);
nor U15751 (N_15751,N_13608,N_14682);
or U15752 (N_15752,N_13440,N_14248);
nor U15753 (N_15753,N_13144,N_14183);
and U15754 (N_15754,N_13512,N_12769);
and U15755 (N_15755,N_14560,N_15385);
nor U15756 (N_15756,N_13915,N_14093);
nand U15757 (N_15757,N_15255,N_12996);
nand U15758 (N_15758,N_14207,N_13063);
and U15759 (N_15759,N_15070,N_14867);
nand U15760 (N_15760,N_13984,N_14676);
or U15761 (N_15761,N_14600,N_13573);
and U15762 (N_15762,N_13323,N_14512);
nand U15763 (N_15763,N_14503,N_12924);
and U15764 (N_15764,N_12504,N_12653);
xor U15765 (N_15765,N_15475,N_15233);
or U15766 (N_15766,N_14240,N_15496);
or U15767 (N_15767,N_12581,N_12663);
nand U15768 (N_15768,N_14707,N_14167);
xor U15769 (N_15769,N_12754,N_14791);
and U15770 (N_15770,N_13476,N_15037);
nor U15771 (N_15771,N_15533,N_14638);
nor U15772 (N_15772,N_15443,N_14588);
and U15773 (N_15773,N_15091,N_14328);
xnor U15774 (N_15774,N_14308,N_13836);
nor U15775 (N_15775,N_15359,N_13164);
nand U15776 (N_15776,N_15568,N_14586);
or U15777 (N_15777,N_13139,N_14648);
nor U15778 (N_15778,N_14507,N_13407);
and U15779 (N_15779,N_13852,N_14126);
or U15780 (N_15780,N_13296,N_14763);
nand U15781 (N_15781,N_14611,N_13814);
nor U15782 (N_15782,N_14844,N_14010);
nand U15783 (N_15783,N_14866,N_13284);
or U15784 (N_15784,N_13588,N_13665);
xnor U15785 (N_15785,N_13374,N_14963);
or U15786 (N_15786,N_12680,N_13239);
nand U15787 (N_15787,N_13051,N_15529);
xor U15788 (N_15788,N_15270,N_14544);
nor U15789 (N_15789,N_13534,N_14065);
nand U15790 (N_15790,N_14039,N_15622);
or U15791 (N_15791,N_14241,N_12619);
xor U15792 (N_15792,N_13444,N_14145);
and U15793 (N_15793,N_14664,N_13846);
nor U15794 (N_15794,N_15400,N_12986);
nor U15795 (N_15795,N_14222,N_13539);
or U15796 (N_15796,N_13020,N_13012);
and U15797 (N_15797,N_12919,N_13211);
nand U15798 (N_15798,N_13976,N_14421);
and U15799 (N_15799,N_14494,N_13265);
and U15800 (N_15800,N_13038,N_14258);
nand U15801 (N_15801,N_12736,N_12827);
or U15802 (N_15802,N_14164,N_14146);
and U15803 (N_15803,N_13470,N_12638);
or U15804 (N_15804,N_13868,N_13029);
nor U15805 (N_15805,N_12743,N_14787);
and U15806 (N_15806,N_14334,N_13271);
nor U15807 (N_15807,N_15180,N_15362);
nor U15808 (N_15808,N_13141,N_14858);
nor U15809 (N_15809,N_15133,N_14860);
or U15810 (N_15810,N_14002,N_14534);
or U15811 (N_15811,N_14103,N_14661);
nor U15812 (N_15812,N_13987,N_12556);
nand U15813 (N_15813,N_13866,N_14027);
xor U15814 (N_15814,N_13414,N_15525);
or U15815 (N_15815,N_14819,N_13459);
xor U15816 (N_15816,N_14059,N_15322);
nand U15817 (N_15817,N_12891,N_14967);
nor U15818 (N_15818,N_12899,N_13955);
xor U15819 (N_15819,N_14277,N_14413);
nor U15820 (N_15820,N_13559,N_13340);
nor U15821 (N_15821,N_14605,N_12757);
nor U15822 (N_15822,N_14660,N_13166);
nand U15823 (N_15823,N_14905,N_15089);
or U15824 (N_15824,N_13259,N_14764);
and U15825 (N_15825,N_15352,N_14902);
nor U15826 (N_15826,N_12548,N_12731);
or U15827 (N_15827,N_12816,N_15257);
nand U15828 (N_15828,N_13090,N_14430);
and U15829 (N_15829,N_15464,N_14904);
nor U15830 (N_15830,N_13365,N_13533);
nand U15831 (N_15831,N_14058,N_15421);
nor U15832 (N_15832,N_15182,N_13572);
xnor U15833 (N_15833,N_14284,N_14310);
xor U15834 (N_15834,N_14446,N_15398);
or U15835 (N_15835,N_12603,N_13195);
and U15836 (N_15836,N_14677,N_14538);
and U15837 (N_15837,N_15116,N_13397);
nor U15838 (N_15838,N_13498,N_13030);
or U15839 (N_15839,N_13153,N_14156);
and U15840 (N_15840,N_14491,N_14041);
or U15841 (N_15841,N_13201,N_15409);
nand U15842 (N_15842,N_15196,N_15336);
nor U15843 (N_15843,N_12667,N_14359);
or U15844 (N_15844,N_15597,N_15125);
and U15845 (N_15845,N_12977,N_15387);
nor U15846 (N_15846,N_13146,N_14134);
nor U15847 (N_15847,N_14121,N_14071);
nor U15848 (N_15848,N_12799,N_12925);
xor U15849 (N_15849,N_13525,N_14466);
and U15850 (N_15850,N_14386,N_13917);
nor U15851 (N_15851,N_13805,N_14804);
nor U15852 (N_15852,N_14685,N_15507);
and U15853 (N_15853,N_14400,N_12620);
and U15854 (N_15854,N_13352,N_13825);
and U15855 (N_15855,N_15330,N_14784);
and U15856 (N_15856,N_14644,N_14865);
and U15857 (N_15857,N_15498,N_14290);
nor U15858 (N_15858,N_14283,N_13336);
or U15859 (N_15859,N_14450,N_15115);
or U15860 (N_15860,N_13168,N_12729);
or U15861 (N_15861,N_14857,N_13118);
and U15862 (N_15862,N_15315,N_15388);
or U15863 (N_15863,N_13688,N_12826);
and U15864 (N_15864,N_14343,N_15338);
or U15865 (N_15865,N_12691,N_15407);
xor U15866 (N_15866,N_13359,N_13819);
nand U15867 (N_15867,N_14173,N_12895);
and U15868 (N_15868,N_14155,N_14254);
and U15869 (N_15869,N_15127,N_12905);
and U15870 (N_15870,N_13536,N_12926);
and U15871 (N_15871,N_13878,N_14987);
or U15872 (N_15872,N_12633,N_13735);
nand U15873 (N_15873,N_14540,N_13300);
nor U15874 (N_15874,N_12983,N_14584);
nor U15875 (N_15875,N_13475,N_14726);
or U15876 (N_15876,N_13941,N_13425);
nand U15877 (N_15877,N_14341,N_13785);
nand U15878 (N_15878,N_15437,N_14216);
and U15879 (N_15879,N_15547,N_13916);
or U15880 (N_15880,N_15450,N_14650);
nor U15881 (N_15881,N_15185,N_13391);
nor U15882 (N_15882,N_13413,N_13485);
and U15883 (N_15883,N_15216,N_13140);
nand U15884 (N_15884,N_14365,N_12949);
nand U15885 (N_15885,N_14796,N_13094);
nand U15886 (N_15886,N_15379,N_15082);
xor U15887 (N_15887,N_13254,N_15042);
nor U15888 (N_15888,N_15175,N_15405);
nand U15889 (N_15889,N_13574,N_15084);
and U15890 (N_15890,N_14451,N_12672);
nand U15891 (N_15891,N_14468,N_15317);
and U15892 (N_15892,N_14576,N_14887);
nor U15893 (N_15893,N_12806,N_15273);
xor U15894 (N_15894,N_12834,N_15303);
or U15895 (N_15895,N_14378,N_13594);
and U15896 (N_15896,N_13237,N_15383);
nor U15897 (N_15897,N_13895,N_15429);
or U15898 (N_15898,N_15411,N_15575);
xor U15899 (N_15899,N_14734,N_14064);
or U15900 (N_15900,N_13729,N_14281);
nand U15901 (N_15901,N_14038,N_13604);
or U15902 (N_15902,N_14633,N_12717);
or U15903 (N_15903,N_14831,N_15325);
nand U15904 (N_15904,N_13791,N_15583);
or U15905 (N_15905,N_13357,N_12930);
and U15906 (N_15906,N_13378,N_13416);
nor U15907 (N_15907,N_14000,N_14130);
or U15908 (N_15908,N_15151,N_12900);
nand U15909 (N_15909,N_14785,N_13714);
or U15910 (N_15910,N_15252,N_13642);
and U15911 (N_15911,N_14178,N_15004);
or U15912 (N_15912,N_15256,N_13629);
nand U15913 (N_15913,N_15408,N_13358);
or U15914 (N_15914,N_12712,N_15572);
and U15915 (N_15915,N_14652,N_12547);
nor U15916 (N_15916,N_14536,N_12501);
and U15917 (N_15917,N_14185,N_12705);
xnor U15918 (N_15918,N_14300,N_15549);
xnor U15919 (N_15919,N_13447,N_14649);
nand U15920 (N_15920,N_15452,N_13433);
and U15921 (N_15921,N_14402,N_13392);
or U15922 (N_15922,N_12909,N_13932);
nand U15923 (N_15923,N_14572,N_14473);
xnor U15924 (N_15924,N_12824,N_14622);
nand U15925 (N_15925,N_14129,N_13759);
xor U15926 (N_15926,N_15565,N_13293);
and U15927 (N_15927,N_12708,N_15491);
nand U15928 (N_15928,N_12894,N_12839);
or U15929 (N_15929,N_14691,N_12918);
nor U15930 (N_15930,N_14424,N_12529);
nand U15931 (N_15931,N_14429,N_12516);
or U15932 (N_15932,N_14715,N_14698);
and U15933 (N_15933,N_13449,N_12665);
or U15934 (N_15934,N_13491,N_14686);
nand U15935 (N_15935,N_14983,N_13494);
nor U15936 (N_15936,N_13657,N_15612);
nand U15937 (N_15937,N_15399,N_14986);
and U15938 (N_15938,N_13858,N_14625);
xnor U15939 (N_15939,N_12844,N_13541);
and U15940 (N_15940,N_14464,N_13411);
or U15941 (N_15941,N_15316,N_12800);
or U15942 (N_15942,N_15214,N_15422);
nand U15943 (N_15943,N_12539,N_13748);
and U15944 (N_15944,N_13615,N_13400);
xor U15945 (N_15945,N_15259,N_14321);
or U15946 (N_15946,N_15426,N_13285);
nor U15947 (N_15947,N_13312,N_13267);
or U15948 (N_15948,N_12830,N_14062);
nor U15949 (N_15949,N_13731,N_15613);
nor U15950 (N_15950,N_13303,N_13730);
or U15951 (N_15951,N_13804,N_15113);
or U15952 (N_15952,N_14256,N_13205);
or U15953 (N_15953,N_12759,N_12921);
nand U15954 (N_15954,N_14774,N_13010);
nand U15955 (N_15955,N_14898,N_13098);
or U15956 (N_15956,N_12681,N_15363);
nor U15957 (N_15957,N_13174,N_13953);
or U15958 (N_15958,N_14104,N_12942);
and U15959 (N_15959,N_13698,N_14636);
and U15960 (N_15960,N_14641,N_13531);
and U15961 (N_15961,N_15438,N_15615);
nor U15962 (N_15962,N_14699,N_13086);
nor U15963 (N_15963,N_14084,N_14320);
nand U15964 (N_15964,N_14376,N_13130);
xnor U15965 (N_15965,N_14981,N_12528);
or U15966 (N_15966,N_15354,N_12902);
or U15967 (N_15967,N_14243,N_15204);
or U15968 (N_15968,N_14833,N_14032);
nor U15969 (N_15969,N_13207,N_15356);
or U15970 (N_15970,N_15278,N_13085);
or U15971 (N_15971,N_13519,N_14478);
nand U15972 (N_15972,N_12884,N_15415);
nand U15973 (N_15973,N_13694,N_14125);
or U15974 (N_15974,N_13666,N_12511);
and U15975 (N_15975,N_12632,N_13457);
or U15976 (N_15976,N_13538,N_14031);
xnor U15977 (N_15977,N_14949,N_14011);
nor U15978 (N_15978,N_13996,N_13870);
xor U15979 (N_15979,N_14219,N_13812);
or U15980 (N_15980,N_14890,N_15319);
nor U15981 (N_15981,N_15229,N_14761);
nor U15982 (N_15982,N_14825,N_13757);
or U15983 (N_15983,N_15164,N_15098);
nand U15984 (N_15984,N_12676,N_13771);
or U15985 (N_15985,N_13226,N_12878);
nand U15986 (N_15986,N_12675,N_14186);
nand U15987 (N_15987,N_13807,N_14618);
nor U15988 (N_15988,N_13127,N_13241);
nand U15989 (N_15989,N_14316,N_15594);
or U15990 (N_15990,N_12810,N_15244);
nor U15991 (N_15991,N_15100,N_14452);
nand U15992 (N_15992,N_13767,N_14862);
xor U15993 (N_15993,N_12542,N_15493);
nand U15994 (N_15994,N_13695,N_14810);
and U15995 (N_15995,N_15258,N_13869);
nand U15996 (N_15996,N_14742,N_12588);
or U15997 (N_15997,N_13843,N_12568);
nor U15998 (N_15998,N_15205,N_14204);
and U15999 (N_15999,N_15564,N_14251);
nor U16000 (N_16000,N_13660,N_15368);
nor U16001 (N_16001,N_15534,N_12641);
and U16002 (N_16002,N_13109,N_12658);
nand U16003 (N_16003,N_15049,N_15620);
and U16004 (N_16004,N_15555,N_14197);
nor U16005 (N_16005,N_15040,N_15413);
or U16006 (N_16006,N_15334,N_14680);
nand U16007 (N_16007,N_14885,N_14974);
nor U16008 (N_16008,N_15588,N_12808);
nand U16009 (N_16009,N_12503,N_14643);
nand U16010 (N_16010,N_12879,N_15190);
nand U16011 (N_16011,N_13579,N_14510);
and U16012 (N_16012,N_13535,N_13755);
and U16013 (N_16013,N_13997,N_12703);
nor U16014 (N_16014,N_15032,N_14561);
or U16015 (N_16015,N_15033,N_12929);
nand U16016 (N_16016,N_12642,N_14245);
nor U16017 (N_16017,N_15126,N_13966);
nand U16018 (N_16018,N_15251,N_13257);
nor U16019 (N_16019,N_15531,N_13458);
xor U16020 (N_16020,N_14855,N_12598);
nand U16021 (N_16021,N_15418,N_13057);
nor U16022 (N_16022,N_12805,N_14521);
nand U16023 (N_16023,N_14353,N_14765);
and U16024 (N_16024,N_14305,N_13669);
and U16025 (N_16025,N_14778,N_14639);
or U16026 (N_16026,N_14782,N_14048);
and U16027 (N_16027,N_13513,N_13592);
and U16028 (N_16028,N_14115,N_12835);
nor U16029 (N_16029,N_15292,N_12892);
or U16030 (N_16030,N_14995,N_14271);
and U16031 (N_16031,N_14026,N_14291);
and U16032 (N_16032,N_13879,N_13739);
nor U16033 (N_16033,N_15170,N_12999);
or U16034 (N_16034,N_13192,N_14013);
nor U16035 (N_16035,N_14552,N_15005);
and U16036 (N_16036,N_13039,N_14231);
or U16037 (N_16037,N_13992,N_14612);
nand U16038 (N_16038,N_15154,N_14325);
and U16039 (N_16039,N_13453,N_12613);
nor U16040 (N_16040,N_13123,N_14459);
or U16041 (N_16041,N_15536,N_14871);
nor U16042 (N_16042,N_13764,N_12972);
or U16043 (N_16043,N_13423,N_13761);
and U16044 (N_16044,N_15608,N_13872);
and U16045 (N_16045,N_13261,N_13684);
nand U16046 (N_16046,N_12610,N_12564);
nand U16047 (N_16047,N_13591,N_14480);
and U16048 (N_16048,N_15038,N_14921);
nor U16049 (N_16049,N_14492,N_15423);
and U16050 (N_16050,N_13246,N_14659);
or U16051 (N_16051,N_13441,N_12728);
and U16052 (N_16052,N_12943,N_13269);
nand U16053 (N_16053,N_12531,N_13222);
nor U16054 (N_16054,N_13577,N_15088);
nor U16055 (N_16055,N_13558,N_14854);
xor U16056 (N_16056,N_14700,N_14813);
nor U16057 (N_16057,N_12749,N_12995);
nand U16058 (N_16058,N_12941,N_13311);
nor U16059 (N_16059,N_12825,N_15136);
or U16060 (N_16060,N_13874,N_14263);
nor U16061 (N_16061,N_13213,N_14880);
nand U16062 (N_16062,N_14889,N_14055);
xnor U16063 (N_16063,N_12848,N_14297);
or U16064 (N_16064,N_14727,N_13469);
nor U16065 (N_16065,N_14792,N_15537);
or U16066 (N_16066,N_12687,N_13417);
nor U16067 (N_16067,N_13609,N_13821);
nor U16068 (N_16068,N_14523,N_14171);
xnor U16069 (N_16069,N_14483,N_12938);
nor U16070 (N_16070,N_14106,N_15559);
or U16071 (N_16071,N_13489,N_14498);
nor U16072 (N_16072,N_15318,N_12804);
nor U16073 (N_16073,N_14379,N_14693);
nor U16074 (N_16074,N_15489,N_14092);
nand U16075 (N_16075,N_13104,N_15460);
or U16076 (N_16076,N_13351,N_14016);
nand U16077 (N_16077,N_13083,N_15576);
nor U16078 (N_16078,N_15002,N_14314);
nand U16079 (N_16079,N_13170,N_14809);
or U16080 (N_16080,N_12742,N_12968);
xnor U16081 (N_16081,N_13775,N_14443);
nand U16082 (N_16082,N_14800,N_14174);
and U16083 (N_16083,N_15162,N_13749);
and U16084 (N_16084,N_13969,N_14745);
and U16085 (N_16085,N_15206,N_13169);
nand U16086 (N_16086,N_15465,N_12518);
nand U16087 (N_16087,N_12822,N_15028);
nor U16088 (N_16088,N_13214,N_13593);
xor U16089 (N_16089,N_15189,N_13601);
nor U16090 (N_16090,N_15131,N_12959);
nand U16091 (N_16091,N_14098,N_15376);
or U16092 (N_16092,N_12797,N_15604);
or U16093 (N_16093,N_13782,N_14626);
xor U16094 (N_16094,N_14182,N_13910);
nand U16095 (N_16095,N_13885,N_13951);
nor U16096 (N_16096,N_13283,N_15476);
or U16097 (N_16097,N_14559,N_14044);
or U16098 (N_16098,N_14603,N_12519);
nor U16099 (N_16099,N_13795,N_15578);
or U16100 (N_16100,N_13837,N_13291);
and U16101 (N_16101,N_12533,N_14170);
nand U16102 (N_16102,N_12690,N_13005);
and U16103 (N_16103,N_14229,N_13310);
xnor U16104 (N_16104,N_13553,N_13645);
or U16105 (N_16105,N_13473,N_15449);
nand U16106 (N_16106,N_12868,N_13673);
nor U16107 (N_16107,N_15332,N_14015);
nand U16108 (N_16108,N_14750,N_12637);
and U16109 (N_16109,N_12677,N_12954);
and U16110 (N_16110,N_12984,N_14574);
nor U16111 (N_16111,N_15511,N_13662);
nor U16112 (N_16112,N_12513,N_12506);
nor U16113 (N_16113,N_14845,N_13683);
and U16114 (N_16114,N_13523,N_14733);
xnor U16115 (N_16115,N_14760,N_14797);
nand U16116 (N_16116,N_13882,N_14108);
nand U16117 (N_16117,N_13251,N_14812);
or U16118 (N_16118,N_12560,N_14465);
and U16119 (N_16119,N_13824,N_12790);
xor U16120 (N_16120,N_13656,N_14775);
or U16121 (N_16121,N_14566,N_13798);
or U16122 (N_16122,N_15545,N_14153);
nor U16123 (N_16123,N_15571,N_15110);
nor U16124 (N_16124,N_13128,N_14928);
or U16125 (N_16125,N_13789,N_12890);
nand U16126 (N_16126,N_15160,N_14074);
nand U16127 (N_16127,N_14728,N_13445);
xnor U16128 (N_16128,N_13725,N_14076);
nand U16129 (N_16129,N_14755,N_15261);
and U16130 (N_16130,N_13484,N_12947);
and U16131 (N_16131,N_14960,N_13888);
xnor U16132 (N_16132,N_13274,N_13650);
nand U16133 (N_16133,N_14590,N_13550);
nand U16134 (N_16134,N_13218,N_15552);
nor U16135 (N_16135,N_13671,N_14925);
and U16136 (N_16136,N_13635,N_14533);
or U16137 (N_16137,N_14786,N_13021);
nor U16138 (N_16138,N_13394,N_14528);
nand U16139 (N_16139,N_13743,N_14445);
nor U16140 (N_16140,N_13845,N_14771);
and U16141 (N_16141,N_12573,N_14139);
nand U16142 (N_16142,N_13646,N_13089);
nor U16143 (N_16143,N_14383,N_13902);
nand U16144 (N_16144,N_15462,N_13058);
or U16145 (N_16145,N_14228,N_15535);
and U16146 (N_16146,N_14920,N_14915);
nor U16147 (N_16147,N_15427,N_12862);
and U16148 (N_16148,N_14522,N_15526);
or U16149 (N_16149,N_12812,N_12913);
and U16150 (N_16150,N_12796,N_14454);
xnor U16151 (N_16151,N_15439,N_14005);
or U16152 (N_16152,N_14081,N_14099);
or U16153 (N_16153,N_13705,N_14768);
or U16154 (N_16154,N_15308,N_13560);
and U16155 (N_16155,N_13321,N_15285);
nand U16156 (N_16156,N_15466,N_14970);
nand U16157 (N_16157,N_14955,N_12980);
and U16158 (N_16158,N_12753,N_13647);
and U16159 (N_16159,N_12741,N_14295);
or U16160 (N_16160,N_12911,N_13270);
or U16161 (N_16161,N_14336,N_12865);
or U16162 (N_16162,N_13703,N_13675);
xor U16163 (N_16163,N_14922,N_13156);
and U16164 (N_16164,N_12933,N_14435);
nor U16165 (N_16165,N_15232,N_13111);
or U16166 (N_16166,N_14090,N_14165);
and U16167 (N_16167,N_15510,N_14720);
nor U16168 (N_16168,N_13971,N_13876);
nand U16169 (N_16169,N_15306,N_13115);
xnor U16170 (N_16170,N_14712,N_14412);
nor U16171 (N_16171,N_14461,N_12960);
nor U16172 (N_16172,N_14711,N_12976);
xnor U16173 (N_16173,N_14539,N_14499);
or U16174 (N_16174,N_13125,N_14077);
nor U16175 (N_16175,N_13154,N_14799);
nor U16176 (N_16176,N_14488,N_14319);
nor U16177 (N_16177,N_14063,N_14416);
nor U16178 (N_16178,N_14748,N_14458);
and U16179 (N_16179,N_14828,N_13778);
nor U16180 (N_16180,N_13811,N_12585);
or U16181 (N_16181,N_14990,N_12766);
nor U16182 (N_16182,N_15485,N_15265);
and U16183 (N_16183,N_13603,N_12600);
or U16184 (N_16184,N_14996,N_14436);
or U16185 (N_16185,N_14340,N_14708);
and U16186 (N_16186,N_12517,N_12609);
nand U16187 (N_16187,N_13653,N_15523);
nor U16188 (N_16188,N_13442,N_15101);
nor U16189 (N_16189,N_13325,N_12792);
nor U16190 (N_16190,N_14147,N_13395);
and U16191 (N_16191,N_12979,N_14244);
or U16192 (N_16192,N_13752,N_14293);
nor U16193 (N_16193,N_15433,N_14043);
and U16194 (N_16194,N_14023,N_14795);
or U16195 (N_16195,N_14040,N_14631);
or U16196 (N_16196,N_14609,N_13408);
nor U16197 (N_16197,N_12778,N_12761);
or U16198 (N_16198,N_14875,N_14347);
or U16199 (N_16199,N_14692,N_13344);
xnor U16200 (N_16200,N_12893,N_14150);
or U16201 (N_16201,N_15172,N_15242);
or U16202 (N_16202,N_14729,N_13081);
nor U16203 (N_16203,N_13151,N_14057);
nand U16204 (N_16204,N_14526,N_13787);
nor U16205 (N_16205,N_13758,N_14382);
and U16206 (N_16206,N_14180,N_12927);
and U16207 (N_16207,N_12837,N_13119);
nand U16208 (N_16208,N_14817,N_13540);
or U16209 (N_16209,N_13193,N_15077);
or U16210 (N_16210,N_12768,N_13639);
or U16211 (N_16211,N_14517,N_12545);
nor U16212 (N_16212,N_14621,N_13911);
and U16213 (N_16213,N_14054,N_12953);
nor U16214 (N_16214,N_13815,N_12565);
and U16215 (N_16215,N_13187,N_14834);
and U16216 (N_16216,N_13920,N_15060);
and U16217 (N_16217,N_14881,N_12849);
nand U16218 (N_16218,N_13620,N_12993);
or U16219 (N_16219,N_13018,N_14212);
or U16220 (N_16220,N_14941,N_14916);
or U16221 (N_16221,N_14056,N_12908);
and U16222 (N_16222,N_14506,N_14531);
nand U16223 (N_16223,N_15313,N_15530);
nand U16224 (N_16224,N_12607,N_13707);
nor U16225 (N_16225,N_13177,N_13216);
and U16226 (N_16226,N_14475,N_12719);
xor U16227 (N_16227,N_13045,N_14689);
nand U16228 (N_16228,N_13256,N_15079);
and U16229 (N_16229,N_12701,N_14658);
nand U16230 (N_16230,N_14166,N_12692);
and U16231 (N_16231,N_13366,N_14061);
nand U16232 (N_16232,N_14377,N_13499);
or U16233 (N_16233,N_15484,N_14111);
nand U16234 (N_16234,N_15590,N_13117);
nor U16235 (N_16235,N_13570,N_13235);
nand U16236 (N_16236,N_14847,N_15592);
and U16237 (N_16237,N_14645,N_14718);
or U16238 (N_16238,N_13329,N_13482);
nand U16239 (N_16239,N_13339,N_13960);
and U16240 (N_16240,N_15556,N_14926);
nand U16241 (N_16241,N_13715,N_13908);
xnor U16242 (N_16242,N_13288,N_12869);
xor U16243 (N_16243,N_14710,N_13353);
nor U16244 (N_16244,N_12557,N_14972);
nor U16245 (N_16245,N_14762,N_14148);
and U16246 (N_16246,N_13649,N_12525);
or U16247 (N_16247,N_12813,N_14276);
nand U16248 (N_16248,N_13188,N_14373);
and U16249 (N_16249,N_15367,N_13132);
or U16250 (N_16250,N_15072,N_13227);
nand U16251 (N_16251,N_14789,N_14897);
nor U16252 (N_16252,N_13659,N_14620);
nor U16253 (N_16253,N_14482,N_14550);
nor U16254 (N_16254,N_15384,N_15081);
xnor U16255 (N_16255,N_13097,N_14628);
xor U16256 (N_16256,N_12904,N_14681);
or U16257 (N_16257,N_13074,N_14345);
or U16258 (N_16258,N_13070,N_14556);
and U16259 (N_16259,N_12684,N_15424);
nand U16260 (N_16260,N_15499,N_13415);
or U16261 (N_16261,N_13999,N_13446);
or U16262 (N_16262,N_15623,N_12775);
and U16263 (N_16263,N_13809,N_15614);
or U16264 (N_16264,N_15454,N_12916);
and U16265 (N_16265,N_12762,N_14200);
nand U16266 (N_16266,N_15288,N_14236);
or U16267 (N_16267,N_14469,N_14903);
nand U16268 (N_16268,N_14548,N_12780);
or U16269 (N_16269,N_15171,N_15337);
nand U16270 (N_16270,N_15611,N_12596);
nand U16271 (N_16271,N_14337,N_13194);
and U16272 (N_16272,N_15035,N_14579);
or U16273 (N_16273,N_13736,N_15297);
or U16274 (N_16274,N_13622,N_14508);
and U16275 (N_16275,N_14994,N_14034);
nor U16276 (N_16276,N_15351,N_15192);
nor U16277 (N_16277,N_14798,N_14545);
nand U16278 (N_16278,N_12714,N_14137);
nor U16279 (N_16279,N_14943,N_14355);
nor U16280 (N_16280,N_14543,N_12866);
or U16281 (N_16281,N_15152,N_13210);
xnor U16282 (N_16282,N_13982,N_15248);
and U16283 (N_16283,N_15074,N_14280);
and U16284 (N_16284,N_14532,N_13309);
and U16285 (N_16285,N_14224,N_15203);
nor U16286 (N_16286,N_14849,N_14730);
nor U16287 (N_16287,N_13520,N_13061);
or U16288 (N_16288,N_13676,N_14423);
or U16289 (N_16289,N_12661,N_15355);
nor U16290 (N_16290,N_13387,N_14460);
nor U16291 (N_16291,N_14331,N_15050);
nor U16292 (N_16292,N_13456,N_13500);
and U16293 (N_16293,N_13532,N_14719);
and U16294 (N_16294,N_15544,N_15558);
nor U16295 (N_16295,N_13055,N_12937);
nand U16296 (N_16296,N_14694,N_13451);
or U16297 (N_16297,N_14739,N_15018);
and U16298 (N_16298,N_13003,N_14360);
and U16299 (N_16299,N_13430,N_13741);
and U16300 (N_16300,N_12785,N_15481);
and U16301 (N_16301,N_13784,N_12952);
nor U16302 (N_16302,N_13595,N_13527);
and U16303 (N_16303,N_13292,N_12821);
nor U16304 (N_16304,N_13396,N_15419);
xnor U16305 (N_16305,N_15017,N_13173);
xor U16306 (N_16306,N_14562,N_14357);
xnor U16307 (N_16307,N_13105,N_12987);
and U16308 (N_16308,N_14953,N_14839);
and U16309 (N_16309,N_13247,N_14741);
nand U16310 (N_16310,N_15506,N_15543);
and U16311 (N_16311,N_13517,N_15518);
nand U16312 (N_16312,N_12592,N_14840);
or U16313 (N_16313,N_15057,N_14836);
or U16314 (N_16314,N_13313,N_14470);
nor U16315 (N_16315,N_14665,N_12589);
nor U16316 (N_16316,N_13080,N_15140);
and U16317 (N_16317,N_14262,N_14978);
and U16318 (N_16318,N_14961,N_14036);
or U16319 (N_16319,N_14717,N_13483);
nand U16320 (N_16320,N_15551,N_13582);
nand U16321 (N_16321,N_13972,N_14891);
or U16322 (N_16322,N_12748,N_14419);
or U16323 (N_16323,N_13149,N_13983);
and U16324 (N_16324,N_13658,N_14037);
nand U16325 (N_16325,N_13160,N_15281);
nand U16326 (N_16326,N_14050,N_12510);
xor U16327 (N_16327,N_15269,N_14292);
nand U16328 (N_16328,N_13137,N_12656);
or U16329 (N_16329,N_12724,N_13348);
and U16330 (N_16330,N_13633,N_13648);
nor U16331 (N_16331,N_13019,N_15584);
or U16332 (N_16332,N_13680,N_13762);
and U16333 (N_16333,N_14723,N_12552);
nor U16334 (N_16334,N_12536,N_15108);
and U16335 (N_16335,N_12599,N_13101);
or U16336 (N_16336,N_15055,N_12730);
nor U16337 (N_16337,N_15567,N_14051);
or U16338 (N_16338,N_15328,N_14666);
nand U16339 (N_16339,N_13054,N_14838);
and U16340 (N_16340,N_13286,N_15107);
nand U16341 (N_16341,N_14333,N_13853);
nand U16342 (N_16342,N_15609,N_13977);
xnor U16343 (N_16343,N_12591,N_13959);
nor U16344 (N_16344,N_13224,N_12814);
nand U16345 (N_16345,N_15150,N_13114);
or U16346 (N_16346,N_13654,N_12650);
nand U16347 (N_16347,N_14018,N_13373);
nor U16348 (N_16348,N_14756,N_15174);
nor U16349 (N_16349,N_14107,N_13155);
nand U16350 (N_16350,N_14873,N_15141);
or U16351 (N_16351,N_14779,N_15104);
xor U16352 (N_16352,N_15486,N_15046);
nor U16353 (N_16353,N_13266,N_15221);
nand U16354 (N_16354,N_13985,N_13851);
nand U16355 (N_16355,N_15041,N_15219);
and U16356 (N_16356,N_15286,N_13143);
and U16357 (N_16357,N_15284,N_12779);
nor U16358 (N_16358,N_13515,N_15482);
or U16359 (N_16359,N_13260,N_15347);
nor U16360 (N_16360,N_14951,N_14175);
or U16361 (N_16361,N_15234,N_14997);
or U16362 (N_16362,N_13120,N_14420);
and U16363 (N_16363,N_13564,N_15036);
and U16364 (N_16364,N_13901,N_13914);
and U16365 (N_16365,N_14684,N_14781);
nand U16366 (N_16366,N_15092,N_14426);
nor U16367 (N_16367,N_15309,N_13892);
nand U16368 (N_16368,N_12502,N_14288);
nand U16369 (N_16369,N_15128,N_15414);
nand U16370 (N_16370,N_15235,N_14546);
and U16371 (N_16371,N_14003,N_15326);
and U16372 (N_16372,N_12786,N_14234);
nand U16373 (N_16373,N_14514,N_14675);
and U16374 (N_16374,N_14346,N_15307);
nand U16375 (N_16375,N_15025,N_13979);
nand U16376 (N_16376,N_14959,N_14195);
or U16377 (N_16377,N_13575,N_13719);
or U16378 (N_16378,N_13848,N_12997);
or U16379 (N_16379,N_13369,N_13307);
nand U16380 (N_16380,N_14646,N_13161);
xnor U16381 (N_16381,N_15135,N_15618);
nand U16382 (N_16382,N_13724,N_14876);
nor U16383 (N_16383,N_12645,N_12688);
and U16384 (N_16384,N_14604,N_14518);
nor U16385 (N_16385,N_14577,N_12735);
xor U16386 (N_16386,N_13726,N_14906);
xor U16387 (N_16387,N_14667,N_13095);
or U16388 (N_16388,N_14900,N_12590);
nor U16389 (N_16389,N_12574,N_12711);
nor U16390 (N_16390,N_13930,N_13863);
nand U16391 (N_16391,N_13643,N_14802);
and U16392 (N_16392,N_14969,N_15617);
xnor U16393 (N_16393,N_13501,N_14725);
nor U16394 (N_16394,N_12720,N_14671);
or U16395 (N_16395,N_13514,N_15197);
or U16396 (N_16396,N_15497,N_14073);
or U16397 (N_16397,N_13701,N_13644);
xor U16398 (N_16398,N_14131,N_14910);
or U16399 (N_16399,N_14127,N_13847);
and U16400 (N_16400,N_13956,N_13186);
or U16401 (N_16401,N_13607,N_14264);
nor U16402 (N_16402,N_12795,N_12773);
nand U16403 (N_16403,N_12644,N_14088);
nand U16404 (N_16404,N_13480,N_13923);
or U16405 (N_16405,N_12955,N_12782);
and U16406 (N_16406,N_15420,N_12554);
or U16407 (N_16407,N_14406,N_12992);
nand U16408 (N_16408,N_12758,N_12882);
nand U16409 (N_16409,N_12831,N_14006);
nor U16410 (N_16410,N_15243,N_12583);
and U16411 (N_16411,N_13652,N_15066);
and U16412 (N_16412,N_13371,N_14892);
and U16413 (N_16413,N_13099,N_13203);
nand U16414 (N_16414,N_13342,N_12704);
nand U16415 (N_16415,N_14287,N_14428);
nor U16416 (N_16416,N_13001,N_13406);
nor U16417 (N_16417,N_13040,N_14701);
nand U16418 (N_16418,N_14403,N_15268);
and U16419 (N_16419,N_13043,N_13014);
nand U16420 (N_16420,N_13315,N_14004);
nor U16421 (N_16421,N_15153,N_13786);
nand U16422 (N_16422,N_13404,N_14738);
nor U16423 (N_16423,N_13506,N_15193);
nand U16424 (N_16424,N_13891,N_14998);
and U16425 (N_16425,N_15254,N_13042);
or U16426 (N_16426,N_13968,N_13421);
nand U16427 (N_16427,N_14884,N_13949);
xnor U16428 (N_16428,N_14835,N_13474);
nand U16429 (N_16429,N_14210,N_12601);
xnor U16430 (N_16430,N_14743,N_15432);
and U16431 (N_16431,N_13253,N_15073);
and U16432 (N_16432,N_15165,N_14747);
nor U16433 (N_16433,N_14770,N_12602);
nor U16434 (N_16434,N_12734,N_12843);
xor U16435 (N_16435,N_14444,N_13036);
and U16436 (N_16436,N_13690,N_13697);
and U16437 (N_16437,N_15300,N_15440);
nor U16438 (N_16438,N_13964,N_15211);
and U16439 (N_16439,N_15155,N_14947);
nor U16440 (N_16440,N_15138,N_13865);
or U16441 (N_16441,N_15026,N_14640);
nor U16442 (N_16442,N_12934,N_13565);
or U16443 (N_16443,N_12535,N_14613);
xor U16444 (N_16444,N_14793,N_13190);
or U16445 (N_16445,N_15022,N_13463);
nand U16446 (N_16446,N_13810,N_13208);
nand U16447 (N_16447,N_14440,N_13817);
xnor U16448 (N_16448,N_12876,N_14917);
or U16449 (N_16449,N_13065,N_14358);
and U16450 (N_16450,N_14911,N_14431);
nand U16451 (N_16451,N_15598,N_13103);
and U16452 (N_16452,N_13826,N_12970);
or U16453 (N_16453,N_15121,N_13011);
and U16454 (N_16454,N_12973,N_13410);
xnor U16455 (N_16455,N_12700,N_15020);
nand U16456 (N_16456,N_12669,N_15451);
xnor U16457 (N_16457,N_14989,N_13828);
xnor U16458 (N_16458,N_12551,N_12875);
nand U16459 (N_16459,N_15301,N_12595);
or U16460 (N_16460,N_13158,N_14285);
nor U16461 (N_16461,N_12507,N_14607);
nor U16462 (N_16462,N_13549,N_12912);
nand U16463 (N_16463,N_12678,N_13510);
or U16464 (N_16464,N_14958,N_13242);
and U16465 (N_16465,N_13578,N_13262);
and U16466 (N_16466,N_12881,N_14176);
and U16467 (N_16467,N_14629,N_12569);
or U16468 (N_16468,N_14397,N_13750);
nor U16469 (N_16469,N_14286,N_15178);
and U16470 (N_16470,N_14030,N_15396);
nor U16471 (N_16471,N_15327,N_14851);
xor U16472 (N_16472,N_15030,N_13861);
nor U16473 (N_16473,N_15053,N_12732);
nand U16474 (N_16474,N_14616,N_12612);
nor U16475 (N_16475,N_13708,N_12967);
or U16476 (N_16476,N_14474,N_14307);
nor U16477 (N_16477,N_14826,N_13945);
xor U16478 (N_16478,N_13605,N_13361);
nor U16479 (N_16479,N_13711,N_14624);
or U16480 (N_16480,N_14594,N_13877);
and U16481 (N_16481,N_13221,N_12580);
xnor U16482 (N_16482,N_15094,N_13581);
and U16483 (N_16483,N_12828,N_15410);
and U16484 (N_16484,N_13922,N_14850);
nor U16485 (N_16485,N_13716,N_14313);
nand U16486 (N_16486,N_13924,N_12571);
xor U16487 (N_16487,N_14289,N_13320);
xnor U16488 (N_16488,N_14367,N_13035);
nor U16489 (N_16489,N_14557,N_13834);
or U16490 (N_16490,N_14587,N_14919);
nor U16491 (N_16491,N_15391,N_14602);
or U16492 (N_16492,N_14122,N_13112);
or U16493 (N_16493,N_12961,N_14933);
nor U16494 (N_16494,N_13487,N_15444);
or U16495 (N_16495,N_13563,N_14193);
or U16496 (N_16496,N_14268,N_14656);
and U16497 (N_16497,N_14954,N_13599);
xnor U16498 (N_16498,N_13232,N_12801);
or U16499 (N_16499,N_15076,N_13196);
nor U16500 (N_16500,N_14842,N_14554);
xor U16501 (N_16501,N_15323,N_14886);
and U16502 (N_16502,N_14722,N_15200);
nor U16503 (N_16503,N_13071,N_13589);
nand U16504 (N_16504,N_15458,N_12861);
and U16505 (N_16505,N_12636,N_13258);
nand U16506 (N_16506,N_12558,N_13280);
and U16507 (N_16507,N_15007,N_13681);
and U16508 (N_16508,N_13880,N_14132);
nand U16509 (N_16509,N_13078,N_13420);
nand U16510 (N_16510,N_15561,N_15566);
xor U16511 (N_16511,N_15348,N_15226);
nand U16512 (N_16512,N_15477,N_14462);
and U16513 (N_16513,N_14140,N_14737);
and U16514 (N_16514,N_15105,N_14028);
xor U16515 (N_16515,N_15225,N_13167);
nand U16516 (N_16516,N_12974,N_14354);
xor U16517 (N_16517,N_15132,N_13634);
and U16518 (N_16518,N_15239,N_14703);
xnor U16519 (N_16519,N_13060,N_13263);
and U16520 (N_16520,N_14918,N_15619);
nor U16521 (N_16521,N_14230,N_12514);
and U16522 (N_16522,N_15202,N_14249);
and U16523 (N_16523,N_14740,N_13840);
or U16524 (N_16524,N_14124,N_14008);
or U16525 (N_16525,N_13503,N_13556);
nand U16526 (N_16526,N_15056,N_14323);
nand U16527 (N_16527,N_15168,N_14252);
nand U16528 (N_16528,N_13052,N_15456);
nand U16529 (N_16529,N_12851,N_15412);
nor U16530 (N_16530,N_13505,N_14190);
nor U16531 (N_16531,N_14655,N_13511);
xor U16532 (N_16532,N_12532,N_13209);
nand U16533 (N_16533,N_14869,N_13068);
and U16534 (N_16534,N_15401,N_14441);
and U16535 (N_16535,N_13180,N_13733);
nor U16536 (N_16536,N_13944,N_14344);
nor U16537 (N_16537,N_14221,N_13661);
nand U16538 (N_16538,N_15003,N_13830);
nand U16539 (N_16539,N_15448,N_12500);
and U16540 (N_16540,N_14437,N_12685);
nor U16541 (N_16541,N_13370,N_13773);
xnor U16542 (N_16542,N_13543,N_13769);
or U16543 (N_16543,N_12978,N_12907);
or U16544 (N_16544,N_15031,N_12526);
xnor U16545 (N_16545,N_12745,N_15459);
xnor U16546 (N_16546,N_13466,N_14999);
or U16547 (N_16547,N_13710,N_14194);
and U16548 (N_16548,N_13148,N_14716);
nand U16549 (N_16549,N_14422,N_15065);
and U16550 (N_16550,N_14322,N_15195);
nor U16551 (N_16551,N_13606,N_12530);
nand U16552 (N_16552,N_12852,N_14599);
and U16553 (N_16553,N_14815,N_14425);
and U16554 (N_16554,N_15579,N_13116);
nand U16555 (N_16555,N_13322,N_13008);
or U16556 (N_16556,N_15169,N_13172);
nand U16557 (N_16557,N_14769,N_13110);
and U16558 (N_16558,N_12622,N_15553);
or U16559 (N_16559,N_14511,N_13053);
nand U16560 (N_16560,N_12584,N_13079);
and U16561 (N_16561,N_14615,N_15339);
nand U16562 (N_16562,N_14338,N_13426);
xor U16563 (N_16563,N_12652,N_13742);
nor U16564 (N_16564,N_14670,N_13376);
nand U16565 (N_16565,N_13897,N_13768);
nand U16566 (N_16566,N_14759,N_14033);
and U16567 (N_16567,N_14189,N_12856);
nand U16568 (N_16568,N_13248,N_13772);
or U16569 (N_16569,N_13087,N_12505);
nor U16570 (N_16570,N_13162,N_14066);
and U16571 (N_16571,N_14752,N_14777);
nand U16572 (N_16572,N_13728,N_12682);
nor U16573 (N_16573,N_12746,N_12555);
nand U16574 (N_16574,N_14870,N_15212);
nand U16575 (N_16575,N_15302,N_14635);
or U16576 (N_16576,N_12945,N_15557);
and U16577 (N_16577,N_14713,N_13839);
xnor U16578 (N_16578,N_13598,N_15118);
and U16579 (N_16579,N_12920,N_12935);
or U16580 (N_16580,N_15463,N_13871);
nor U16581 (N_16581,N_13890,N_15215);
nand U16582 (N_16582,N_13142,N_15607);
xnor U16583 (N_16583,N_14706,N_13062);
and U16584 (N_16584,N_14823,N_15023);
nand U16585 (N_16585,N_13689,N_12567);
or U16586 (N_16586,N_12776,N_13672);
nand U16587 (N_16587,N_15375,N_14332);
nand U16588 (N_16588,N_15109,N_13025);
nand U16589 (N_16589,N_14520,N_13894);
or U16590 (N_16590,N_12847,N_14114);
nor U16591 (N_16591,N_12702,N_12509);
or U16592 (N_16592,N_15240,N_13024);
xor U16593 (N_16593,N_14133,N_12994);
xor U16594 (N_16594,N_14551,N_15335);
and U16595 (N_16595,N_13185,N_12586);
and U16596 (N_16596,N_13200,N_13522);
xnor U16597 (N_16597,N_12863,N_12765);
or U16598 (N_16598,N_13380,N_12777);
nor U16599 (N_16599,N_14965,N_13732);
or U16600 (N_16600,N_13571,N_13638);
or U16601 (N_16601,N_12914,N_13379);
or U16602 (N_16602,N_14940,N_13282);
and U16603 (N_16603,N_13720,N_14110);
and U16604 (N_16604,N_14942,N_15341);
and U16605 (N_16605,N_13838,N_14370);
nor U16606 (N_16606,N_13860,N_14683);
and U16607 (N_16607,N_14872,N_12752);
nand U16608 (N_16608,N_15096,N_12639);
nor U16609 (N_16609,N_13547,N_12737);
xnor U16610 (N_16610,N_14893,N_15021);
and U16611 (N_16611,N_14119,N_15250);
and U16612 (N_16612,N_15577,N_14120);
nor U16613 (N_16613,N_13106,N_13943);
and U16614 (N_16614,N_14363,N_15207);
nor U16615 (N_16615,N_13077,N_13611);
and U16616 (N_16616,N_13562,N_12932);
nor U16617 (N_16617,N_13674,N_14589);
and U16618 (N_16618,N_14962,N_13092);
or U16619 (N_16619,N_14991,N_13760);
xor U16620 (N_16620,N_14816,N_13687);
and U16621 (N_16621,N_14086,N_13435);
and U16622 (N_16622,N_14017,N_13277);
nor U16623 (N_16623,N_15593,N_13461);
nand U16624 (N_16624,N_12815,N_13402);
xnor U16625 (N_16625,N_15034,N_14012);
xnor U16626 (N_16626,N_13013,N_12521);
and U16627 (N_16627,N_15490,N_13134);
nand U16628 (N_16628,N_13341,N_14569);
nor U16629 (N_16629,N_15158,N_13316);
or U16630 (N_16630,N_13954,N_12870);
nand U16631 (N_16631,N_14950,N_13075);
and U16632 (N_16632,N_14790,N_15369);
or U16633 (N_16633,N_15078,N_14564);
nor U16634 (N_16634,N_15014,N_14246);
nand U16635 (N_16635,N_14496,N_13857);
or U16636 (N_16636,N_12627,N_13942);
or U16637 (N_16637,N_13746,N_12623);
and U16638 (N_16638,N_14046,N_13368);
nor U16639 (N_16639,N_14934,N_14198);
xor U16640 (N_16640,N_13129,N_14215);
nand U16641 (N_16641,N_13434,N_13931);
or U16642 (N_16642,N_15009,N_12750);
xnor U16643 (N_16643,N_15587,N_13306);
and U16644 (N_16644,N_13841,N_13630);
nand U16645 (N_16645,N_14731,N_13198);
and U16646 (N_16646,N_15106,N_13452);
nand U16647 (N_16647,N_13126,N_14094);
and U16648 (N_16648,N_13529,N_14766);
or U16649 (N_16649,N_14151,N_15194);
nand U16650 (N_16650,N_14136,N_13450);
nand U16651 (N_16651,N_12944,N_13849);
nor U16652 (N_16652,N_12858,N_13472);
nor U16653 (N_16653,N_14392,N_14388);
nor U16654 (N_16654,N_15538,N_15461);
or U16655 (N_16655,N_12764,N_14079);
and U16656 (N_16656,N_14824,N_14438);
nand U16657 (N_16657,N_13165,N_13388);
nor U16658 (N_16658,N_13833,N_13082);
and U16659 (N_16659,N_12877,N_15389);
or U16660 (N_16660,N_15610,N_13428);
nor U16661 (N_16661,N_13947,N_12738);
or U16662 (N_16662,N_14901,N_14601);
nor U16663 (N_16663,N_12971,N_13738);
or U16664 (N_16664,N_14515,N_15582);
and U16665 (N_16665,N_13829,N_14025);
nand U16666 (N_16666,N_14827,N_14160);
nor U16667 (N_16667,N_14203,N_13567);
nor U16668 (N_16668,N_14303,N_13754);
nand U16669 (N_16669,N_13756,N_15374);
nand U16670 (N_16670,N_14976,N_14829);
nand U16671 (N_16671,N_15512,N_14477);
nor U16672 (N_16672,N_14396,N_14754);
or U16673 (N_16673,N_14163,N_15377);
and U16674 (N_16674,N_14113,N_12695);
or U16675 (N_16675,N_13252,N_13135);
nand U16676 (N_16676,N_15198,N_12706);
nor U16677 (N_16677,N_13245,N_14398);
and U16678 (N_16678,N_13422,N_15290);
nor U16679 (N_16679,N_13345,N_15487);
or U16680 (N_16680,N_14758,N_13561);
and U16681 (N_16681,N_13967,N_13667);
nor U16682 (N_16682,N_14753,N_15173);
nor U16683 (N_16683,N_15142,N_15469);
nand U16684 (N_16684,N_12975,N_13243);
nand U16685 (N_16685,N_13419,N_12854);
xnor U16686 (N_16686,N_14007,N_13859);
nor U16687 (N_16687,N_14408,N_14806);
or U16688 (N_16688,N_15516,N_14266);
and U16689 (N_16689,N_15188,N_15117);
nor U16690 (N_16690,N_12860,N_13918);
nand U16691 (N_16691,N_14149,N_14582);
or U16692 (N_16692,N_15470,N_14966);
nor U16693 (N_16693,N_13929,N_15130);
or U16694 (N_16694,N_13718,N_15378);
xnor U16695 (N_16695,N_13067,N_12906);
and U16696 (N_16696,N_15483,N_14929);
and U16697 (N_16697,N_14411,N_14964);
nand U16698 (N_16698,N_14082,N_13206);
and U16699 (N_16699,N_14265,N_15054);
nor U16700 (N_16700,N_13781,N_14924);
nand U16701 (N_16701,N_12922,N_13600);
and U16702 (N_16702,N_15166,N_12615);
nor U16703 (N_16703,N_14335,N_15550);
nor U16704 (N_16704,N_13957,N_14434);
nand U16705 (N_16705,N_12725,N_15380);
nand U16706 (N_16706,N_13528,N_13526);
nor U16707 (N_16707,N_13948,N_14223);
nor U16708 (N_16708,N_14668,N_12727);
nand U16709 (N_16709,N_15011,N_13276);
nor U16710 (N_16710,N_14567,N_14856);
and U16711 (N_16711,N_12991,N_13338);
and U16712 (N_16712,N_14818,N_13844);
or U16713 (N_16713,N_15447,N_13326);
and U16714 (N_16714,N_13504,N_12699);
and U16715 (N_16715,N_14529,N_12546);
nor U16716 (N_16716,N_14371,N_12563);
nor U16717 (N_16717,N_12985,N_12648);
and U16718 (N_16718,N_13016,N_15581);
xor U16719 (N_16719,N_13217,N_13088);
nand U16720 (N_16720,N_13382,N_15000);
nand U16721 (N_16721,N_13632,N_13566);
and U16722 (N_16722,N_14788,N_12643);
or U16723 (N_16723,N_13516,N_14863);
and U16724 (N_16724,N_12540,N_12624);
nor U16725 (N_16725,N_12807,N_13580);
and U16726 (N_16726,N_15016,N_14931);
nand U16727 (N_16727,N_14647,N_15333);
and U16728 (N_16728,N_12631,N_15231);
and U16729 (N_16729,N_15514,N_15294);
or U16730 (N_16730,N_12651,N_14776);
and U16731 (N_16731,N_14674,N_12659);
or U16732 (N_16732,N_13801,N_14206);
or U16733 (N_16733,N_15344,N_13279);
xnor U16734 (N_16734,N_14580,N_13439);
nand U16735 (N_16735,N_15271,N_12625);
nor U16736 (N_16736,N_14364,N_15589);
and U16737 (N_16737,N_14843,N_15295);
nor U16738 (N_16738,N_12886,N_12689);
nand U16739 (N_16739,N_13034,N_12629);
or U16740 (N_16740,N_15227,N_15097);
or U16741 (N_16741,N_15027,N_13796);
or U16742 (N_16742,N_15321,N_12874);
nor U16743 (N_16743,N_12965,N_13928);
and U16744 (N_16744,N_15276,N_12957);
nand U16745 (N_16745,N_14820,N_15509);
nor U16746 (N_16746,N_14233,N_13938);
and U16747 (N_16747,N_13808,N_15280);
xnor U16748 (N_16748,N_15157,N_13780);
and U16749 (N_16749,N_15163,N_15015);
and U16750 (N_16750,N_15541,N_13102);
xor U16751 (N_16751,N_13462,N_15548);
nand U16752 (N_16752,N_13327,N_14078);
nor U16753 (N_16753,N_12559,N_14349);
or U16754 (N_16754,N_14808,N_13331);
and U16755 (N_16755,N_13176,N_13069);
and U16756 (N_16756,N_15099,N_15305);
or U16757 (N_16757,N_14118,N_14101);
nor U16758 (N_16758,N_13486,N_15508);
nor U16759 (N_16759,N_14654,N_13290);
xor U16760 (N_16760,N_15320,N_13788);
nand U16761 (N_16761,N_13641,N_12817);
and U16762 (N_16762,N_13899,N_13862);
nor U16763 (N_16763,N_12898,N_14487);
and U16764 (N_16764,N_15585,N_13072);
and U16765 (N_16765,N_13383,N_13424);
nand U16766 (N_16766,N_13318,N_14565);
nor U16767 (N_16767,N_15010,N_14351);
and U16768 (N_16768,N_15029,N_13980);
and U16769 (N_16769,N_14936,N_15395);
nand U16770 (N_16770,N_13171,N_13268);
xnor U16771 (N_16771,N_15430,N_13377);
or U16772 (N_16772,N_13740,N_15080);
or U16773 (N_16773,N_14009,N_12756);
and U16774 (N_16774,N_14695,N_14070);
xor U16775 (N_16775,N_14399,N_14927);
or U16776 (N_16776,N_14168,N_15217);
nand U16777 (N_16777,N_14971,N_13432);
or U16778 (N_16778,N_13776,N_15342);
or U16779 (N_16779,N_13418,N_15184);
and U16780 (N_16780,N_13046,N_13989);
or U16781 (N_16781,N_13385,N_13751);
or U16782 (N_16782,N_15404,N_14227);
and U16783 (N_16783,N_12561,N_15087);
and U16784 (N_16784,N_13816,N_12544);
or U16785 (N_16785,N_13896,N_13823);
or U16786 (N_16786,N_13548,N_14410);
or U16787 (N_16787,N_14982,N_14394);
nor U16788 (N_16788,N_15350,N_13934);
or U16789 (N_16789,N_13384,N_15393);
and U16790 (N_16790,N_12722,N_13590);
or U16791 (N_16791,N_14899,N_12962);
nand U16792 (N_16792,N_15103,N_14401);
nor U16793 (N_16793,N_12793,N_15479);
nand U16794 (N_16794,N_15102,N_12887);
and U16795 (N_16795,N_13250,N_12772);
nor U16796 (N_16796,N_15364,N_14882);
and U16797 (N_16797,N_13028,N_12527);
nor U16798 (N_16798,N_12635,N_15502);
nand U16799 (N_16799,N_14878,N_13906);
nor U16800 (N_16800,N_13122,N_13479);
or U16801 (N_16801,N_13919,N_13624);
xor U16802 (N_16802,N_15602,N_12616);
or U16803 (N_16803,N_13699,N_13637);
nor U16804 (N_16804,N_14463,N_15048);
nor U16805 (N_16805,N_12990,N_15513);
and U16806 (N_16806,N_13904,N_15580);
and U16807 (N_16807,N_13405,N_15001);
xnor U16808 (N_16808,N_14476,N_14744);
or U16809 (N_16809,N_14162,N_13299);
nand U16810 (N_16810,N_15329,N_15563);
nor U16811 (N_16811,N_14563,N_14085);
or U16812 (N_16812,N_14158,N_12948);
or U16813 (N_16813,N_14896,N_13264);
or U16814 (N_16814,N_14279,N_12524);
nor U16815 (N_16815,N_13970,N_14100);
or U16816 (N_16816,N_14138,N_14324);
nand U16817 (N_16817,N_12605,N_15472);
and U16818 (N_16818,N_13183,N_13616);
and U16819 (N_16819,N_14805,N_12566);
nand U16820 (N_16820,N_13530,N_14312);
nor U16821 (N_16821,N_13212,N_14022);
or U16822 (N_16822,N_12696,N_13818);
and U16823 (N_16823,N_13508,N_13360);
and U16824 (N_16824,N_14883,N_15311);
and U16825 (N_16825,N_15123,N_15236);
and U16826 (N_16826,N_14442,N_15570);
or U16827 (N_16827,N_15397,N_14705);
nand U16828 (N_16828,N_13393,N_15149);
or U16829 (N_16829,N_15291,N_14091);
nor U16830 (N_16830,N_15246,N_12604);
or U16831 (N_16831,N_13349,N_14052);
or U16832 (N_16832,N_15277,N_13492);
nor U16833 (N_16833,N_13093,N_13973);
nand U16834 (N_16834,N_12950,N_13178);
nor U16835 (N_16835,N_13700,N_13015);
nor U16836 (N_16836,N_15061,N_15119);
nand U16837 (N_16837,N_14260,N_13797);
and U16838 (N_16838,N_13356,N_14298);
nand U16839 (N_16839,N_13524,N_14269);
nor U16840 (N_16840,N_14568,N_13006);
or U16841 (N_16841,N_15478,N_13455);
or U16842 (N_16842,N_15230,N_12710);
nand U16843 (N_16843,N_13794,N_13544);
or U16844 (N_16844,N_12606,N_15218);
nor U16845 (N_16845,N_13610,N_15143);
xor U16846 (N_16846,N_14457,N_15392);
and U16847 (N_16847,N_12614,N_15358);
nand U16848 (N_16848,N_15179,N_13883);
or U16849 (N_16849,N_12838,N_13230);
xor U16850 (N_16850,N_12755,N_13017);
or U16851 (N_16851,N_14669,N_13375);
nand U16852 (N_16852,N_14746,N_14001);
and U16853 (N_16853,N_12923,N_14973);
nor U16854 (N_16854,N_15208,N_12666);
and U16855 (N_16855,N_13249,N_14497);
and U16856 (N_16856,N_14985,N_13679);
nor U16857 (N_16857,N_14939,N_14144);
nor U16858 (N_16858,N_13273,N_14678);
and U16859 (N_16859,N_13806,N_15304);
nand U16860 (N_16860,N_13995,N_14992);
xor U16861 (N_16861,N_13295,N_13220);
and U16862 (N_16862,N_13820,N_15435);
nor U16863 (N_16863,N_14830,N_15331);
nand U16864 (N_16864,N_13048,N_14945);
xnor U16865 (N_16865,N_14541,N_12969);
and U16866 (N_16866,N_12572,N_15501);
nor U16867 (N_16867,N_13233,N_13096);
nor U16868 (N_16868,N_12575,N_13903);
nor U16869 (N_16869,N_13712,N_14495);
or U16870 (N_16870,N_15299,N_13713);
nand U16871 (N_16871,N_15181,N_13962);
or U16872 (N_16872,N_14608,N_13554);
or U16873 (N_16873,N_14938,N_12562);
nor U16874 (N_16874,N_14571,N_15540);
nand U16875 (N_16875,N_14591,N_14627);
nor U16876 (N_16876,N_14935,N_13569);
nor U16877 (N_16877,N_14117,N_14944);
nand U16878 (N_16878,N_13790,N_14570);
nor U16879 (N_16879,N_15519,N_13744);
nor U16880 (N_16880,N_12570,N_12857);
and U16881 (N_16881,N_13302,N_13272);
nand U16882 (N_16882,N_13033,N_15349);
nor U16883 (N_16883,N_15137,N_15390);
nor U16884 (N_16884,N_14361,N_13685);
nor U16885 (N_16885,N_13113,N_15177);
or U16886 (N_16886,N_13179,N_14448);
or U16887 (N_16887,N_15044,N_14217);
xor U16888 (N_16888,N_14868,N_14447);
nand U16889 (N_16889,N_13471,N_13950);
nand U16890 (N_16890,N_14366,N_15467);
nand U16891 (N_16891,N_14874,N_13546);
or U16892 (N_16892,N_14089,N_15183);
xor U16893 (N_16893,N_14455,N_13696);
nor U16894 (N_16894,N_14387,N_15148);
or U16895 (N_16895,N_13493,N_13986);
or U16896 (N_16896,N_15573,N_13287);
and U16897 (N_16897,N_12654,N_13881);
and U16898 (N_16898,N_13614,N_15569);
nor U16899 (N_16899,N_12832,N_15340);
and U16900 (N_16900,N_12787,N_13912);
and U16901 (N_16901,N_14205,N_13152);
nand U16902 (N_16902,N_13585,N_15289);
nor U16903 (N_16903,N_12936,N_14374);
or U16904 (N_16904,N_14047,N_15365);
nand U16905 (N_16905,N_14968,N_13334);
xor U16906 (N_16906,N_14369,N_15370);
nor U16907 (N_16907,N_15019,N_14542);
and U16908 (N_16908,N_15298,N_13783);
nor U16909 (N_16909,N_13159,N_15406);
nor U16910 (N_16910,N_15279,N_15431);
nor U16911 (N_16911,N_13993,N_13774);
and U16912 (N_16912,N_12896,N_12715);
or U16913 (N_16913,N_15596,N_13478);
xnor U16914 (N_16914,N_14525,N_12657);
xnor U16915 (N_16915,N_13027,N_13401);
nor U16916 (N_16916,N_14736,N_14213);
nand U16917 (N_16917,N_15112,N_14097);
nor U16918 (N_16918,N_13994,N_14095);
nand U16919 (N_16919,N_14390,N_13921);
nor U16920 (N_16920,N_13150,N_15008);
xor U16921 (N_16921,N_14087,N_14772);
and U16922 (N_16922,N_15471,N_13958);
nand U16923 (N_16923,N_14453,N_15345);
nor U16924 (N_16924,N_13026,N_14519);
nand U16925 (N_16925,N_14606,N_13963);
nor U16926 (N_16926,N_15222,N_15263);
and U16927 (N_16927,N_13275,N_13389);
nand U16928 (N_16928,N_14080,N_14250);
and U16929 (N_16929,N_15052,N_14932);
nand U16930 (N_16930,N_13832,N_14732);
and U16931 (N_16931,N_12883,N_14024);
or U16932 (N_16932,N_13765,N_12726);
nor U16933 (N_16933,N_14329,N_15039);
and U16934 (N_16934,N_13856,N_13050);
nor U16935 (N_16935,N_15542,N_13289);
and U16936 (N_16936,N_12640,N_13032);
nand U16937 (N_16937,N_13332,N_14535);
or U16938 (N_16938,N_13779,N_12903);
or U16939 (N_16939,N_14467,N_13076);
and U16940 (N_16940,N_12747,N_13507);
nand U16941 (N_16941,N_13488,N_15488);
and U16942 (N_16942,N_15075,N_14673);
nand U16943 (N_16943,N_14979,N_12721);
nor U16944 (N_16944,N_13557,N_13988);
nor U16945 (N_16945,N_14220,N_12989);
nand U16946 (N_16946,N_13621,N_13913);
and U16947 (N_16947,N_12723,N_15312);
nand U16948 (N_16948,N_15067,N_15416);
nand U16949 (N_16949,N_15603,N_13521);
and U16950 (N_16950,N_15051,N_14427);
nor U16951 (N_16951,N_13136,N_13933);
nor U16952 (N_16952,N_14696,N_12694);
nand U16953 (N_16953,N_14984,N_14109);
and U16954 (N_16954,N_14877,N_13347);
and U16955 (N_16955,N_13909,N_12649);
nand U16956 (N_16956,N_12673,N_13842);
nor U16957 (N_16957,N_13722,N_12897);
and U16958 (N_16958,N_12739,N_14783);
and U16959 (N_16959,N_15223,N_13031);
or U16960 (N_16960,N_12550,N_15366);
or U16961 (N_16961,N_12597,N_14135);
or U16962 (N_16962,N_15473,N_14181);
nor U16963 (N_16963,N_13792,N_12873);
nor U16964 (N_16964,N_13946,N_13372);
or U16965 (N_16965,N_12880,N_14342);
and U16966 (N_16966,N_15283,N_14481);
nand U16967 (N_16967,N_14553,N_13056);
and U16968 (N_16968,N_12850,N_14822);
nor U16969 (N_16969,N_12611,N_14261);
xor U16970 (N_16970,N_14894,N_12522);
nand U16971 (N_16971,N_12840,N_13004);
nor U16972 (N_16972,N_14988,N_14757);
nor U16973 (N_16973,N_15266,N_14749);
and U16974 (N_16974,N_13022,N_14634);
xnor U16975 (N_16975,N_14274,N_15224);
or U16976 (N_16976,N_12802,N_13314);
nand U16977 (N_16977,N_15267,N_14301);
nand U16978 (N_16978,N_12534,N_12576);
nor U16979 (N_16979,N_15606,N_13477);
nand U16980 (N_16980,N_13328,N_13234);
or U16981 (N_16981,N_13802,N_14242);
nand U16982 (N_16982,N_14610,N_14801);
nand U16983 (N_16983,N_12662,N_15272);
and U16984 (N_16984,N_13002,N_14662);
and U16985 (N_16985,N_14530,N_14391);
nor U16986 (N_16986,N_13537,N_13301);
or U16987 (N_16987,N_13427,N_12788);
nor U16988 (N_16988,N_13317,N_13612);
nand U16989 (N_16989,N_12628,N_15139);
and U16990 (N_16990,N_13803,N_13244);
nor U16991 (N_16991,N_14225,N_14253);
nor U16992 (N_16992,N_15260,N_12523);
nor U16993 (N_16993,N_12733,N_13618);
nand U16994 (N_16994,N_13628,N_14773);
and U16995 (N_16995,N_13631,N_13350);
nand U16996 (N_16996,N_14583,N_12928);
nand U16997 (N_16997,N_13813,N_15045);
nor U16998 (N_16998,N_13961,N_15209);
or U16999 (N_16999,N_12707,N_13281);
nor U17000 (N_17000,N_12668,N_12679);
and U17001 (N_17001,N_15156,N_15241);
nand U17002 (N_17002,N_13131,N_14143);
or U17003 (N_17003,N_14811,N_15360);
nor U17004 (N_17004,N_13636,N_14490);
nand U17005 (N_17005,N_13403,N_13777);
and U17006 (N_17006,N_14201,N_14888);
nand U17007 (N_17007,N_14177,N_14069);
nand U17008 (N_17008,N_14389,N_15144);
nand U17009 (N_17009,N_12859,N_13091);
or U17010 (N_17010,N_14527,N_14053);
or U17011 (N_17011,N_15122,N_13197);
or U17012 (N_17012,N_13240,N_14471);
nand U17013 (N_17013,N_14272,N_13324);
nor U17014 (N_17014,N_12791,N_14304);
or U17015 (N_17015,N_14348,N_12718);
or U17016 (N_17016,N_14952,N_15446);
and U17017 (N_17017,N_14141,N_13727);
or U17018 (N_17018,N_15062,N_12618);
or U17019 (N_17019,N_12740,N_15191);
nor U17020 (N_17020,N_13737,N_14537);
or U17021 (N_17021,N_13651,N_12520);
and U17022 (N_17022,N_13974,N_13335);
or U17023 (N_17023,N_14687,N_12577);
nand U17024 (N_17024,N_15093,N_14072);
nand U17025 (N_17025,N_14592,N_14306);
nand U17026 (N_17026,N_14267,N_13721);
nand U17027 (N_17027,N_15574,N_13655);
nand U17028 (N_17028,N_15237,N_13678);
nor U17029 (N_17029,N_14296,N_13182);
and U17030 (N_17030,N_13800,N_15554);
and U17031 (N_17031,N_14404,N_14105);
xor U17032 (N_17032,N_14479,N_13386);
or U17033 (N_17033,N_14688,N_13465);
and U17034 (N_17034,N_13157,N_15085);
or U17035 (N_17035,N_12958,N_15495);
or U17036 (N_17036,N_13399,N_14585);
nand U17037 (N_17037,N_13049,N_13887);
or U17038 (N_17038,N_13497,N_15403);
and U17039 (N_17039,N_14102,N_13481);
nand U17040 (N_17040,N_13905,N_14767);
nand U17041 (N_17041,N_13626,N_15599);
or U17042 (N_17042,N_14975,N_13346);
and U17043 (N_17043,N_15324,N_13884);
or U17044 (N_17044,N_14302,N_13693);
nand U17045 (N_17045,N_13398,N_13184);
nand U17046 (N_17046,N_13175,N_15453);
and U17047 (N_17047,N_14619,N_14083);
or U17048 (N_17048,N_13255,N_12646);
nand U17049 (N_17049,N_14275,N_12931);
nor U17050 (N_17050,N_14067,N_13677);
or U17051 (N_17051,N_14914,N_14395);
xnor U17052 (N_17052,N_13939,N_14068);
and U17053 (N_17053,N_12760,N_13023);
nand U17054 (N_17054,N_15480,N_15167);
nor U17055 (N_17055,N_15145,N_15186);
and U17056 (N_17056,N_13181,N_14330);
xor U17057 (N_17057,N_13298,N_14672);
and U17058 (N_17058,N_15357,N_14179);
xor U17059 (N_17059,N_14913,N_15120);
xor U17060 (N_17060,N_15500,N_13509);
and U17061 (N_17061,N_13084,N_12617);
or U17062 (N_17062,N_13454,N_14597);
or U17063 (N_17063,N_12781,N_15213);
nand U17064 (N_17064,N_12634,N_12829);
or U17065 (N_17065,N_15434,N_12846);
nor U17066 (N_17066,N_13586,N_14513);
nor U17067 (N_17067,N_12811,N_14923);
and U17068 (N_17068,N_12579,N_12823);
or U17069 (N_17069,N_13965,N_14697);
nand U17070 (N_17070,N_14637,N_14502);
nand U17071 (N_17071,N_15524,N_15527);
and U17072 (N_17072,N_13925,N_14282);
nor U17073 (N_17073,N_14239,N_12966);
nand U17074 (N_17074,N_13822,N_13436);
xor U17075 (N_17075,N_15441,N_12578);
or U17076 (N_17076,N_12803,N_13998);
or U17077 (N_17077,N_12593,N_14751);
and U17078 (N_17078,N_14385,N_12582);
or U17079 (N_17079,N_14218,N_13044);
and U17080 (N_17080,N_12774,N_14029);
nand U17081 (N_17081,N_12888,N_15417);
nand U17082 (N_17082,N_13236,N_13278);
or U17083 (N_17083,N_15562,N_14702);
or U17084 (N_17084,N_13191,N_14294);
or U17085 (N_17085,N_14315,N_15515);
nand U17086 (N_17086,N_13596,N_14380);
nor U17087 (N_17087,N_15253,N_14196);
nand U17088 (N_17088,N_13367,N_14721);
nand U17089 (N_17089,N_14821,N_12951);
and U17090 (N_17090,N_15314,N_14414);
or U17091 (N_17091,N_14327,N_13907);
and U17092 (N_17092,N_15024,N_12841);
nand U17093 (N_17093,N_15372,N_15591);
nand U17094 (N_17094,N_13627,N_13009);
nand U17095 (N_17095,N_14846,N_13935);
nand U17096 (N_17096,N_14841,N_12864);
nand U17097 (N_17097,N_15517,N_15275);
nor U17098 (N_17098,N_14614,N_14188);
nor U17099 (N_17099,N_12697,N_14326);
or U17100 (N_17100,N_14339,N_14309);
and U17101 (N_17101,N_13551,N_15129);
nor U17102 (N_17102,N_15605,N_13354);
nand U17103 (N_17103,N_15176,N_14299);
nor U17104 (N_17104,N_12515,N_15492);
nor U17105 (N_17105,N_15210,N_13640);
and U17106 (N_17106,N_12946,N_13991);
nor U17107 (N_17107,N_13231,N_13333);
nand U17108 (N_17108,N_13831,N_13202);
or U17109 (N_17109,N_13363,N_13121);
and U17110 (N_17110,N_15083,N_14709);
or U17111 (N_17111,N_15086,N_15386);
and U17112 (N_17112,N_15114,N_13663);
and U17113 (N_17113,N_14848,N_14879);
or U17114 (N_17114,N_14152,N_14853);
nor U17115 (N_17115,N_14679,N_12767);
or U17116 (N_17116,N_14352,N_14381);
and U17117 (N_17117,N_15346,N_14257);
and U17118 (N_17118,N_13064,N_12698);
xor U17119 (N_17119,N_14735,N_13204);
or U17120 (N_17120,N_13704,N_15616);
nor U17121 (N_17121,N_14558,N_13568);
nand U17122 (N_17122,N_14049,N_15296);
nand U17123 (N_17123,N_14472,N_15064);
nand U17124 (N_17124,N_13041,N_15373);
or U17125 (N_17125,N_15071,N_13238);
and U17126 (N_17126,N_14270,N_14714);
and U17127 (N_17127,N_13745,N_14128);
nand U17128 (N_17128,N_14957,N_12771);
or U17129 (N_17129,N_14907,N_14449);
and U17130 (N_17130,N_12674,N_14123);
or U17131 (N_17131,N_15521,N_14489);
nor U17132 (N_17132,N_15600,N_13617);
nand U17133 (N_17133,N_13007,N_14653);
nor U17134 (N_17134,N_14255,N_14235);
or U17135 (N_17135,N_14859,N_12915);
nand U17136 (N_17136,N_13889,N_15245);
nor U17137 (N_17137,N_15228,N_15012);
or U17138 (N_17138,N_13936,N_12671);
xor U17139 (N_17139,N_13495,N_13875);
xnor U17140 (N_17140,N_13464,N_14946);
and U17141 (N_17141,N_14418,N_15199);
and U17142 (N_17142,N_13542,N_14259);
or U17143 (N_17143,N_13587,N_13873);
or U17144 (N_17144,N_12964,N_14630);
or U17145 (N_17145,N_13855,N_14663);
nor U17146 (N_17146,N_14504,N_14439);
nand U17147 (N_17147,N_14154,N_15090);
and U17148 (N_17148,N_14956,N_13552);
xor U17149 (N_17149,N_14157,N_15287);
nand U17150 (N_17150,N_13753,N_15586);
or U17151 (N_17151,N_12956,N_12770);
or U17152 (N_17152,N_12541,N_12664);
or U17153 (N_17153,N_14930,N_13927);
xnor U17154 (N_17154,N_13225,N_12853);
nor U17155 (N_17155,N_13898,N_12998);
or U17156 (N_17156,N_15621,N_15293);
nand U17157 (N_17157,N_14433,N_13723);
nand U17158 (N_17158,N_13952,N_13518);
or U17159 (N_17159,N_12744,N_12889);
nand U17160 (N_17160,N_14794,N_14832);
or U17161 (N_17161,N_14704,N_14318);
and U17162 (N_17162,N_12621,N_14937);
or U17163 (N_17163,N_12794,N_15247);
or U17164 (N_17164,N_14780,N_15381);
and U17165 (N_17165,N_14948,N_12836);
and U17166 (N_17166,N_14837,N_12939);
or U17167 (N_17167,N_13975,N_13709);
or U17168 (N_17168,N_13412,N_12512);
nand U17169 (N_17169,N_13308,N_12538);
nor U17170 (N_17170,N_14191,N_14187);
nor U17171 (N_17171,N_12784,N_14035);
nor U17172 (N_17172,N_14019,N_13364);
nand U17173 (N_17173,N_13496,N_13437);
and U17174 (N_17174,N_14368,N_12660);
nor U17175 (N_17175,N_14493,N_15068);
or U17176 (N_17176,N_15445,N_12845);
or U17177 (N_17177,N_13940,N_12587);
nand U17178 (N_17178,N_14159,N_13059);
nor U17179 (N_17179,N_14814,N_13390);
and U17180 (N_17180,N_15425,N_13625);
and U17181 (N_17181,N_13330,N_12819);
nor U17182 (N_17182,N_13355,N_13886);
or U17183 (N_17183,N_13597,N_14912);
or U17184 (N_17184,N_15095,N_14724);
or U17185 (N_17185,N_12798,N_14595);
and U17186 (N_17186,N_14632,N_13545);
and U17187 (N_17187,N_13000,N_14226);
or U17188 (N_17188,N_12505,N_14403);
or U17189 (N_17189,N_14697,N_13812);
nor U17190 (N_17190,N_15202,N_14084);
xnor U17191 (N_17191,N_13509,N_12504);
or U17192 (N_17192,N_13102,N_14076);
nor U17193 (N_17193,N_13486,N_15373);
nand U17194 (N_17194,N_13964,N_15041);
and U17195 (N_17195,N_13715,N_15340);
nor U17196 (N_17196,N_14353,N_14993);
nand U17197 (N_17197,N_13114,N_12561);
nand U17198 (N_17198,N_14848,N_14419);
and U17199 (N_17199,N_13253,N_14487);
nor U17200 (N_17200,N_13443,N_12817);
nor U17201 (N_17201,N_14316,N_14991);
nand U17202 (N_17202,N_14076,N_13928);
nor U17203 (N_17203,N_12527,N_13791);
xor U17204 (N_17204,N_13617,N_14804);
or U17205 (N_17205,N_14703,N_14793);
nor U17206 (N_17206,N_14301,N_13936);
or U17207 (N_17207,N_15246,N_12928);
xor U17208 (N_17208,N_14122,N_14652);
nand U17209 (N_17209,N_13818,N_13244);
xor U17210 (N_17210,N_14267,N_15285);
nand U17211 (N_17211,N_15507,N_14952);
nor U17212 (N_17212,N_13558,N_14472);
or U17213 (N_17213,N_14884,N_13102);
nand U17214 (N_17214,N_14751,N_12654);
nand U17215 (N_17215,N_13598,N_14479);
nor U17216 (N_17216,N_13721,N_14368);
and U17217 (N_17217,N_14095,N_14570);
nor U17218 (N_17218,N_12639,N_13459);
or U17219 (N_17219,N_13441,N_15395);
or U17220 (N_17220,N_13758,N_13682);
or U17221 (N_17221,N_14998,N_14590);
nand U17222 (N_17222,N_12866,N_14910);
or U17223 (N_17223,N_13416,N_14045);
or U17224 (N_17224,N_14414,N_15290);
or U17225 (N_17225,N_14939,N_15242);
or U17226 (N_17226,N_15334,N_13229);
and U17227 (N_17227,N_15528,N_15118);
or U17228 (N_17228,N_14268,N_13873);
xnor U17229 (N_17229,N_15425,N_13979);
nor U17230 (N_17230,N_12907,N_13853);
and U17231 (N_17231,N_14868,N_15242);
nand U17232 (N_17232,N_13050,N_13697);
and U17233 (N_17233,N_13954,N_14738);
nor U17234 (N_17234,N_13000,N_14709);
nor U17235 (N_17235,N_15194,N_13992);
or U17236 (N_17236,N_12907,N_12889);
nand U17237 (N_17237,N_14722,N_14877);
nor U17238 (N_17238,N_13320,N_15347);
nand U17239 (N_17239,N_14233,N_15142);
nand U17240 (N_17240,N_13936,N_13297);
nand U17241 (N_17241,N_14314,N_12659);
or U17242 (N_17242,N_15046,N_15319);
and U17243 (N_17243,N_14919,N_14178);
or U17244 (N_17244,N_14195,N_13589);
nor U17245 (N_17245,N_14076,N_14562);
nand U17246 (N_17246,N_13060,N_13987);
xor U17247 (N_17247,N_13189,N_13605);
or U17248 (N_17248,N_14197,N_14445);
nor U17249 (N_17249,N_13213,N_15398);
nor U17250 (N_17250,N_15318,N_15613);
nor U17251 (N_17251,N_12712,N_13089);
or U17252 (N_17252,N_14069,N_15523);
and U17253 (N_17253,N_15323,N_13653);
nor U17254 (N_17254,N_14316,N_15280);
or U17255 (N_17255,N_13693,N_13527);
nor U17256 (N_17256,N_14443,N_13424);
nand U17257 (N_17257,N_13350,N_15502);
nor U17258 (N_17258,N_14670,N_15387);
or U17259 (N_17259,N_12747,N_13617);
or U17260 (N_17260,N_15095,N_14011);
and U17261 (N_17261,N_14982,N_13814);
and U17262 (N_17262,N_13397,N_13725);
and U17263 (N_17263,N_14050,N_15041);
nand U17264 (N_17264,N_13816,N_13448);
or U17265 (N_17265,N_13003,N_14108);
nor U17266 (N_17266,N_15447,N_14563);
nor U17267 (N_17267,N_13909,N_12605);
nor U17268 (N_17268,N_14116,N_13335);
xor U17269 (N_17269,N_14579,N_14265);
nor U17270 (N_17270,N_14039,N_15574);
nand U17271 (N_17271,N_12917,N_12672);
xor U17272 (N_17272,N_13367,N_14400);
nand U17273 (N_17273,N_14973,N_13959);
nor U17274 (N_17274,N_13516,N_12575);
or U17275 (N_17275,N_14119,N_15386);
and U17276 (N_17276,N_15112,N_15088);
xor U17277 (N_17277,N_14325,N_14500);
nor U17278 (N_17278,N_15182,N_13833);
and U17279 (N_17279,N_13306,N_14868);
or U17280 (N_17280,N_13343,N_14940);
nand U17281 (N_17281,N_13258,N_14915);
nand U17282 (N_17282,N_13097,N_14114);
nand U17283 (N_17283,N_14736,N_13209);
and U17284 (N_17284,N_14829,N_14881);
and U17285 (N_17285,N_13817,N_14735);
nor U17286 (N_17286,N_15074,N_15400);
nand U17287 (N_17287,N_13135,N_14880);
nor U17288 (N_17288,N_13990,N_13299);
xor U17289 (N_17289,N_13298,N_12875);
and U17290 (N_17290,N_14644,N_14823);
or U17291 (N_17291,N_13819,N_13280);
nor U17292 (N_17292,N_12607,N_14925);
nand U17293 (N_17293,N_15270,N_13285);
xnor U17294 (N_17294,N_13997,N_13280);
or U17295 (N_17295,N_13084,N_14564);
nor U17296 (N_17296,N_15591,N_13127);
nor U17297 (N_17297,N_14587,N_12772);
and U17298 (N_17298,N_14420,N_14342);
nand U17299 (N_17299,N_13407,N_13527);
and U17300 (N_17300,N_14925,N_13247);
or U17301 (N_17301,N_14076,N_12921);
or U17302 (N_17302,N_15391,N_13677);
nor U17303 (N_17303,N_13614,N_12669);
or U17304 (N_17304,N_13554,N_13887);
and U17305 (N_17305,N_13884,N_13170);
and U17306 (N_17306,N_15255,N_12657);
and U17307 (N_17307,N_12946,N_12854);
nor U17308 (N_17308,N_14958,N_15047);
and U17309 (N_17309,N_13128,N_13148);
nor U17310 (N_17310,N_14493,N_13778);
nand U17311 (N_17311,N_14344,N_12549);
or U17312 (N_17312,N_14535,N_14708);
nand U17313 (N_17313,N_13833,N_15214);
nor U17314 (N_17314,N_14174,N_13663);
nand U17315 (N_17315,N_12793,N_13735);
xnor U17316 (N_17316,N_13437,N_13222);
or U17317 (N_17317,N_14242,N_13320);
or U17318 (N_17318,N_15119,N_15164);
nor U17319 (N_17319,N_12656,N_15520);
nand U17320 (N_17320,N_15500,N_14145);
and U17321 (N_17321,N_12876,N_15329);
nor U17322 (N_17322,N_13355,N_14600);
nand U17323 (N_17323,N_12977,N_13587);
and U17324 (N_17324,N_13192,N_12987);
and U17325 (N_17325,N_12987,N_13202);
and U17326 (N_17326,N_14651,N_15358);
or U17327 (N_17327,N_13506,N_13078);
xor U17328 (N_17328,N_14883,N_13570);
and U17329 (N_17329,N_13423,N_14180);
nor U17330 (N_17330,N_14537,N_13850);
nor U17331 (N_17331,N_13531,N_14573);
nor U17332 (N_17332,N_13814,N_13372);
xnor U17333 (N_17333,N_14277,N_13347);
nand U17334 (N_17334,N_15117,N_13323);
and U17335 (N_17335,N_13535,N_14473);
and U17336 (N_17336,N_12830,N_13693);
or U17337 (N_17337,N_14290,N_12811);
and U17338 (N_17338,N_14040,N_13032);
xnor U17339 (N_17339,N_14037,N_15197);
or U17340 (N_17340,N_13419,N_13130);
and U17341 (N_17341,N_14099,N_14586);
xor U17342 (N_17342,N_14421,N_15535);
and U17343 (N_17343,N_14849,N_13633);
nand U17344 (N_17344,N_13845,N_13578);
nand U17345 (N_17345,N_15268,N_12755);
and U17346 (N_17346,N_12641,N_15551);
xnor U17347 (N_17347,N_14683,N_15303);
nand U17348 (N_17348,N_14858,N_14515);
and U17349 (N_17349,N_13307,N_13314);
nand U17350 (N_17350,N_13790,N_15030);
xor U17351 (N_17351,N_13621,N_14120);
xnor U17352 (N_17352,N_13316,N_14776);
or U17353 (N_17353,N_14304,N_13113);
and U17354 (N_17354,N_15508,N_12585);
nand U17355 (N_17355,N_14100,N_15620);
or U17356 (N_17356,N_13346,N_12907);
nand U17357 (N_17357,N_14055,N_14316);
nand U17358 (N_17358,N_15326,N_15194);
nand U17359 (N_17359,N_14772,N_13696);
xor U17360 (N_17360,N_12961,N_13134);
or U17361 (N_17361,N_13287,N_14963);
or U17362 (N_17362,N_14849,N_13502);
nand U17363 (N_17363,N_15283,N_15215);
or U17364 (N_17364,N_14635,N_12724);
nor U17365 (N_17365,N_13490,N_12825);
or U17366 (N_17366,N_14009,N_15047);
and U17367 (N_17367,N_13884,N_13685);
nor U17368 (N_17368,N_14708,N_14449);
xnor U17369 (N_17369,N_15017,N_14138);
or U17370 (N_17370,N_13746,N_14831);
nand U17371 (N_17371,N_14881,N_15224);
xnor U17372 (N_17372,N_12895,N_13698);
and U17373 (N_17373,N_12503,N_12772);
xnor U17374 (N_17374,N_14728,N_14917);
nand U17375 (N_17375,N_13876,N_13106);
and U17376 (N_17376,N_12704,N_13612);
and U17377 (N_17377,N_13177,N_13296);
or U17378 (N_17378,N_12663,N_12796);
and U17379 (N_17379,N_13468,N_13976);
xnor U17380 (N_17380,N_12880,N_13003);
nand U17381 (N_17381,N_14957,N_12728);
xor U17382 (N_17382,N_13218,N_14665);
and U17383 (N_17383,N_14943,N_14125);
nand U17384 (N_17384,N_14045,N_14499);
nor U17385 (N_17385,N_14835,N_14389);
or U17386 (N_17386,N_13810,N_12579);
xor U17387 (N_17387,N_12627,N_14819);
and U17388 (N_17388,N_13009,N_12533);
xor U17389 (N_17389,N_14712,N_14173);
and U17390 (N_17390,N_13511,N_13744);
nor U17391 (N_17391,N_13882,N_13235);
nand U17392 (N_17392,N_14077,N_14231);
nand U17393 (N_17393,N_13762,N_13633);
and U17394 (N_17394,N_13283,N_13033);
nor U17395 (N_17395,N_15414,N_15573);
xor U17396 (N_17396,N_14815,N_13234);
nand U17397 (N_17397,N_13525,N_15274);
and U17398 (N_17398,N_13700,N_12673);
or U17399 (N_17399,N_15146,N_14393);
and U17400 (N_17400,N_14465,N_13361);
or U17401 (N_17401,N_14318,N_14959);
nor U17402 (N_17402,N_13221,N_14794);
or U17403 (N_17403,N_13853,N_15408);
and U17404 (N_17404,N_13201,N_13040);
nor U17405 (N_17405,N_13037,N_13157);
or U17406 (N_17406,N_12771,N_15039);
nor U17407 (N_17407,N_15117,N_15088);
xor U17408 (N_17408,N_12940,N_13848);
and U17409 (N_17409,N_14562,N_14313);
nand U17410 (N_17410,N_14161,N_12592);
nand U17411 (N_17411,N_13614,N_13319);
and U17412 (N_17412,N_13580,N_15424);
xor U17413 (N_17413,N_12973,N_14879);
or U17414 (N_17414,N_14163,N_14622);
or U17415 (N_17415,N_15228,N_13732);
nand U17416 (N_17416,N_13763,N_14687);
and U17417 (N_17417,N_13650,N_13980);
nor U17418 (N_17418,N_15553,N_13184);
and U17419 (N_17419,N_14314,N_13919);
and U17420 (N_17420,N_12791,N_13067);
nor U17421 (N_17421,N_15341,N_15061);
or U17422 (N_17422,N_14273,N_14875);
and U17423 (N_17423,N_14068,N_14480);
nor U17424 (N_17424,N_13335,N_13129);
xnor U17425 (N_17425,N_13143,N_14850);
nand U17426 (N_17426,N_14804,N_14285);
or U17427 (N_17427,N_13235,N_12502);
and U17428 (N_17428,N_15614,N_13031);
nand U17429 (N_17429,N_14597,N_14787);
or U17430 (N_17430,N_12868,N_13251);
nand U17431 (N_17431,N_13481,N_13254);
and U17432 (N_17432,N_15523,N_15275);
nand U17433 (N_17433,N_14985,N_14026);
or U17434 (N_17434,N_13986,N_15372);
xor U17435 (N_17435,N_13209,N_14308);
nand U17436 (N_17436,N_14530,N_13787);
or U17437 (N_17437,N_15252,N_15341);
xor U17438 (N_17438,N_13021,N_14733);
and U17439 (N_17439,N_13168,N_13008);
nand U17440 (N_17440,N_15307,N_12677);
or U17441 (N_17441,N_13224,N_12974);
nand U17442 (N_17442,N_14532,N_13217);
nand U17443 (N_17443,N_14486,N_14040);
and U17444 (N_17444,N_14696,N_15453);
xor U17445 (N_17445,N_12881,N_14393);
nand U17446 (N_17446,N_12733,N_14326);
nand U17447 (N_17447,N_13934,N_12960);
and U17448 (N_17448,N_13370,N_15112);
xnor U17449 (N_17449,N_13542,N_14168);
or U17450 (N_17450,N_15258,N_14791);
or U17451 (N_17451,N_12631,N_14055);
nor U17452 (N_17452,N_14966,N_14719);
nor U17453 (N_17453,N_13942,N_13443);
xor U17454 (N_17454,N_14744,N_14657);
xnor U17455 (N_17455,N_13964,N_14429);
xor U17456 (N_17456,N_12661,N_15069);
and U17457 (N_17457,N_12729,N_13662);
or U17458 (N_17458,N_13268,N_15417);
nand U17459 (N_17459,N_14267,N_13091);
and U17460 (N_17460,N_12731,N_14557);
nand U17461 (N_17461,N_13648,N_15017);
or U17462 (N_17462,N_12876,N_15086);
and U17463 (N_17463,N_14565,N_13494);
or U17464 (N_17464,N_13226,N_13121);
nand U17465 (N_17465,N_14255,N_12710);
and U17466 (N_17466,N_13053,N_13101);
nand U17467 (N_17467,N_12661,N_14603);
nand U17468 (N_17468,N_13014,N_12860);
and U17469 (N_17469,N_13334,N_13377);
and U17470 (N_17470,N_13443,N_12569);
and U17471 (N_17471,N_14093,N_13752);
or U17472 (N_17472,N_14030,N_14512);
or U17473 (N_17473,N_13827,N_15116);
nor U17474 (N_17474,N_13172,N_15235);
nor U17475 (N_17475,N_13502,N_13985);
nor U17476 (N_17476,N_14881,N_14360);
or U17477 (N_17477,N_15061,N_13312);
nand U17478 (N_17478,N_13316,N_15095);
and U17479 (N_17479,N_15103,N_14926);
or U17480 (N_17480,N_13424,N_15272);
nor U17481 (N_17481,N_13721,N_15334);
and U17482 (N_17482,N_15309,N_13956);
and U17483 (N_17483,N_13375,N_14912);
nor U17484 (N_17484,N_14886,N_14443);
nor U17485 (N_17485,N_12961,N_15545);
and U17486 (N_17486,N_15117,N_14185);
and U17487 (N_17487,N_15326,N_15203);
nand U17488 (N_17488,N_12572,N_14707);
and U17489 (N_17489,N_15126,N_14910);
nand U17490 (N_17490,N_15119,N_13218);
and U17491 (N_17491,N_13221,N_12808);
nand U17492 (N_17492,N_12784,N_13284);
or U17493 (N_17493,N_13017,N_14999);
and U17494 (N_17494,N_15047,N_14624);
xor U17495 (N_17495,N_12508,N_15077);
xnor U17496 (N_17496,N_12751,N_14053);
or U17497 (N_17497,N_13385,N_14164);
and U17498 (N_17498,N_13328,N_13852);
nor U17499 (N_17499,N_14056,N_13571);
nor U17500 (N_17500,N_15213,N_14097);
or U17501 (N_17501,N_14460,N_13583);
or U17502 (N_17502,N_13169,N_15216);
and U17503 (N_17503,N_14491,N_12977);
or U17504 (N_17504,N_13907,N_15424);
or U17505 (N_17505,N_15102,N_15286);
or U17506 (N_17506,N_13458,N_15073);
xor U17507 (N_17507,N_15183,N_13112);
nor U17508 (N_17508,N_15342,N_13193);
or U17509 (N_17509,N_14852,N_13111);
and U17510 (N_17510,N_15305,N_12647);
and U17511 (N_17511,N_13934,N_15439);
and U17512 (N_17512,N_13080,N_15314);
nor U17513 (N_17513,N_15251,N_14041);
and U17514 (N_17514,N_14299,N_14616);
nand U17515 (N_17515,N_13711,N_12657);
nor U17516 (N_17516,N_12767,N_14115);
nand U17517 (N_17517,N_13743,N_13969);
or U17518 (N_17518,N_12629,N_13356);
nand U17519 (N_17519,N_12646,N_13441);
and U17520 (N_17520,N_14716,N_14589);
and U17521 (N_17521,N_13402,N_13629);
or U17522 (N_17522,N_15028,N_14473);
and U17523 (N_17523,N_14391,N_14740);
or U17524 (N_17524,N_13083,N_13634);
or U17525 (N_17525,N_14912,N_14216);
nand U17526 (N_17526,N_15543,N_12938);
and U17527 (N_17527,N_13838,N_14108);
and U17528 (N_17528,N_14197,N_13815);
nand U17529 (N_17529,N_15409,N_14757);
and U17530 (N_17530,N_14157,N_14637);
or U17531 (N_17531,N_15326,N_13374);
and U17532 (N_17532,N_12875,N_14926);
nand U17533 (N_17533,N_12529,N_14917);
nor U17534 (N_17534,N_13433,N_15258);
nor U17535 (N_17535,N_13804,N_15426);
nand U17536 (N_17536,N_14257,N_14130);
and U17537 (N_17537,N_14509,N_13569);
and U17538 (N_17538,N_12847,N_15129);
xnor U17539 (N_17539,N_13275,N_13448);
nand U17540 (N_17540,N_12565,N_13512);
or U17541 (N_17541,N_15518,N_13899);
nor U17542 (N_17542,N_12921,N_12563);
or U17543 (N_17543,N_13484,N_13091);
nor U17544 (N_17544,N_15004,N_13841);
and U17545 (N_17545,N_14719,N_12517);
or U17546 (N_17546,N_12952,N_13399);
nand U17547 (N_17547,N_13117,N_13062);
nand U17548 (N_17548,N_14199,N_14316);
and U17549 (N_17549,N_14560,N_14092);
and U17550 (N_17550,N_14560,N_13330);
nor U17551 (N_17551,N_12640,N_12909);
and U17552 (N_17552,N_13492,N_13280);
xor U17553 (N_17553,N_12725,N_13526);
nor U17554 (N_17554,N_14114,N_15405);
or U17555 (N_17555,N_12980,N_12597);
and U17556 (N_17556,N_14429,N_13639);
nor U17557 (N_17557,N_14452,N_14227);
nand U17558 (N_17558,N_12585,N_13836);
or U17559 (N_17559,N_14997,N_13092);
and U17560 (N_17560,N_12719,N_13486);
and U17561 (N_17561,N_14895,N_15617);
and U17562 (N_17562,N_13299,N_15050);
nand U17563 (N_17563,N_12651,N_12636);
or U17564 (N_17564,N_14283,N_13801);
nand U17565 (N_17565,N_13902,N_15254);
xor U17566 (N_17566,N_14183,N_13644);
nand U17567 (N_17567,N_14737,N_15620);
nor U17568 (N_17568,N_13194,N_15231);
nor U17569 (N_17569,N_13430,N_15441);
or U17570 (N_17570,N_15176,N_14250);
and U17571 (N_17571,N_13478,N_14871);
nand U17572 (N_17572,N_12778,N_12552);
nand U17573 (N_17573,N_14476,N_13642);
xnor U17574 (N_17574,N_13937,N_13119);
or U17575 (N_17575,N_13800,N_13168);
nand U17576 (N_17576,N_15441,N_14309);
nand U17577 (N_17577,N_14681,N_12966);
or U17578 (N_17578,N_15199,N_13686);
and U17579 (N_17579,N_14080,N_13110);
and U17580 (N_17580,N_14735,N_13964);
nand U17581 (N_17581,N_15140,N_14064);
nand U17582 (N_17582,N_13966,N_15348);
nor U17583 (N_17583,N_12559,N_12585);
and U17584 (N_17584,N_13916,N_14708);
and U17585 (N_17585,N_14937,N_14959);
and U17586 (N_17586,N_15076,N_13658);
or U17587 (N_17587,N_14323,N_14789);
nand U17588 (N_17588,N_14814,N_13038);
or U17589 (N_17589,N_14502,N_14943);
nand U17590 (N_17590,N_15544,N_15532);
nor U17591 (N_17591,N_12759,N_13273);
nand U17592 (N_17592,N_14240,N_12929);
xor U17593 (N_17593,N_13981,N_13480);
and U17594 (N_17594,N_12678,N_14463);
or U17595 (N_17595,N_12831,N_14462);
and U17596 (N_17596,N_15608,N_12873);
nor U17597 (N_17597,N_13681,N_14255);
nor U17598 (N_17598,N_14105,N_12830);
and U17599 (N_17599,N_13607,N_12591);
and U17600 (N_17600,N_13166,N_13009);
nor U17601 (N_17601,N_15039,N_12547);
or U17602 (N_17602,N_13515,N_14443);
xor U17603 (N_17603,N_15191,N_15134);
xor U17604 (N_17604,N_14535,N_13700);
or U17605 (N_17605,N_14627,N_15056);
or U17606 (N_17606,N_12724,N_14337);
and U17607 (N_17607,N_15121,N_13095);
xnor U17608 (N_17608,N_12949,N_13847);
nor U17609 (N_17609,N_15574,N_15151);
or U17610 (N_17610,N_14794,N_15577);
nand U17611 (N_17611,N_15455,N_14040);
nor U17612 (N_17612,N_15510,N_15527);
or U17613 (N_17613,N_15551,N_13830);
and U17614 (N_17614,N_14591,N_14669);
and U17615 (N_17615,N_13640,N_15322);
nor U17616 (N_17616,N_13393,N_13821);
or U17617 (N_17617,N_14667,N_13783);
xnor U17618 (N_17618,N_14223,N_14514);
and U17619 (N_17619,N_14968,N_13760);
and U17620 (N_17620,N_12870,N_13406);
nand U17621 (N_17621,N_14126,N_14909);
and U17622 (N_17622,N_12653,N_12683);
and U17623 (N_17623,N_13085,N_13262);
nand U17624 (N_17624,N_13065,N_12882);
nand U17625 (N_17625,N_14216,N_15473);
and U17626 (N_17626,N_14745,N_13922);
xnor U17627 (N_17627,N_14382,N_13471);
nor U17628 (N_17628,N_13915,N_14927);
and U17629 (N_17629,N_15023,N_12698);
and U17630 (N_17630,N_14898,N_13542);
nor U17631 (N_17631,N_14734,N_15110);
xnor U17632 (N_17632,N_12895,N_13033);
nand U17633 (N_17633,N_13001,N_14016);
or U17634 (N_17634,N_15487,N_13029);
xor U17635 (N_17635,N_13343,N_15509);
or U17636 (N_17636,N_15231,N_14529);
nor U17637 (N_17637,N_13534,N_15432);
nor U17638 (N_17638,N_12971,N_14969);
and U17639 (N_17639,N_13252,N_13050);
nand U17640 (N_17640,N_12791,N_13300);
xnor U17641 (N_17641,N_13342,N_14988);
and U17642 (N_17642,N_13696,N_12784);
and U17643 (N_17643,N_13018,N_13235);
nor U17644 (N_17644,N_15551,N_14916);
nand U17645 (N_17645,N_14383,N_14043);
nand U17646 (N_17646,N_15255,N_14583);
and U17647 (N_17647,N_15297,N_12910);
and U17648 (N_17648,N_13999,N_15022);
and U17649 (N_17649,N_12749,N_13448);
or U17650 (N_17650,N_13763,N_15253);
nor U17651 (N_17651,N_13784,N_14026);
nor U17652 (N_17652,N_15055,N_15316);
or U17653 (N_17653,N_15197,N_13982);
or U17654 (N_17654,N_13565,N_12608);
nor U17655 (N_17655,N_14788,N_14393);
and U17656 (N_17656,N_12647,N_14347);
xnor U17657 (N_17657,N_14781,N_14867);
or U17658 (N_17658,N_14634,N_15523);
or U17659 (N_17659,N_13830,N_13036);
and U17660 (N_17660,N_14804,N_13781);
nand U17661 (N_17661,N_12629,N_15064);
nand U17662 (N_17662,N_12560,N_12887);
nor U17663 (N_17663,N_14341,N_14035);
nand U17664 (N_17664,N_12718,N_13659);
or U17665 (N_17665,N_14361,N_14210);
nand U17666 (N_17666,N_13407,N_15161);
nand U17667 (N_17667,N_13835,N_13126);
and U17668 (N_17668,N_13757,N_13957);
nor U17669 (N_17669,N_13964,N_14002);
nand U17670 (N_17670,N_14919,N_12806);
nor U17671 (N_17671,N_12933,N_13122);
nand U17672 (N_17672,N_12679,N_15292);
or U17673 (N_17673,N_13934,N_15413);
or U17674 (N_17674,N_15044,N_12990);
and U17675 (N_17675,N_14243,N_14466);
nor U17676 (N_17676,N_13555,N_13831);
and U17677 (N_17677,N_13535,N_15413);
nor U17678 (N_17678,N_14834,N_13751);
nor U17679 (N_17679,N_13074,N_14578);
xor U17680 (N_17680,N_15107,N_13419);
and U17681 (N_17681,N_14088,N_15388);
or U17682 (N_17682,N_14008,N_13187);
and U17683 (N_17683,N_14215,N_15312);
or U17684 (N_17684,N_13272,N_12779);
and U17685 (N_17685,N_14116,N_13063);
nand U17686 (N_17686,N_13371,N_13137);
nor U17687 (N_17687,N_14143,N_14773);
nor U17688 (N_17688,N_12668,N_14978);
xnor U17689 (N_17689,N_15542,N_13712);
and U17690 (N_17690,N_13022,N_14312);
xor U17691 (N_17691,N_15017,N_14460);
xnor U17692 (N_17692,N_13866,N_14472);
nand U17693 (N_17693,N_15131,N_13511);
or U17694 (N_17694,N_15300,N_15555);
nand U17695 (N_17695,N_12694,N_13242);
nand U17696 (N_17696,N_15504,N_15230);
and U17697 (N_17697,N_12957,N_12514);
nand U17698 (N_17698,N_13007,N_13551);
nor U17699 (N_17699,N_14205,N_14856);
or U17700 (N_17700,N_13157,N_14433);
and U17701 (N_17701,N_13806,N_14950);
nand U17702 (N_17702,N_14651,N_14799);
nand U17703 (N_17703,N_12753,N_12975);
and U17704 (N_17704,N_15288,N_12875);
nor U17705 (N_17705,N_13768,N_12928);
nand U17706 (N_17706,N_14347,N_14956);
and U17707 (N_17707,N_15520,N_13249);
nand U17708 (N_17708,N_14893,N_13545);
nor U17709 (N_17709,N_15355,N_14560);
nand U17710 (N_17710,N_15508,N_12621);
xor U17711 (N_17711,N_14712,N_15567);
and U17712 (N_17712,N_12947,N_13655);
or U17713 (N_17713,N_12533,N_14127);
nand U17714 (N_17714,N_15305,N_13491);
nand U17715 (N_17715,N_13139,N_14321);
nor U17716 (N_17716,N_14437,N_14260);
and U17717 (N_17717,N_14129,N_14600);
and U17718 (N_17718,N_13995,N_14322);
xor U17719 (N_17719,N_13071,N_14314);
or U17720 (N_17720,N_14283,N_13860);
and U17721 (N_17721,N_14384,N_13690);
xor U17722 (N_17722,N_12768,N_13012);
and U17723 (N_17723,N_13511,N_13049);
nor U17724 (N_17724,N_14352,N_13331);
nor U17725 (N_17725,N_13088,N_12719);
nor U17726 (N_17726,N_13930,N_13874);
nand U17727 (N_17727,N_12968,N_14169);
nor U17728 (N_17728,N_15362,N_14596);
or U17729 (N_17729,N_14638,N_12781);
or U17730 (N_17730,N_14308,N_12690);
nor U17731 (N_17731,N_13823,N_14462);
nor U17732 (N_17732,N_14644,N_13369);
nor U17733 (N_17733,N_14483,N_14556);
and U17734 (N_17734,N_15385,N_14540);
nor U17735 (N_17735,N_13943,N_14202);
nor U17736 (N_17736,N_13232,N_14205);
or U17737 (N_17737,N_14556,N_13045);
or U17738 (N_17738,N_14358,N_13420);
xor U17739 (N_17739,N_14089,N_12684);
and U17740 (N_17740,N_13874,N_13305);
or U17741 (N_17741,N_13952,N_15290);
nor U17742 (N_17742,N_13851,N_15399);
and U17743 (N_17743,N_15263,N_13560);
xor U17744 (N_17744,N_15028,N_14855);
nor U17745 (N_17745,N_14554,N_14340);
and U17746 (N_17746,N_14766,N_14944);
nor U17747 (N_17747,N_12743,N_14804);
and U17748 (N_17748,N_13973,N_13922);
nand U17749 (N_17749,N_13409,N_14498);
and U17750 (N_17750,N_14301,N_14597);
nand U17751 (N_17751,N_13191,N_12928);
nand U17752 (N_17752,N_15491,N_13347);
nor U17753 (N_17753,N_13614,N_12637);
xor U17754 (N_17754,N_14317,N_14102);
and U17755 (N_17755,N_15164,N_13512);
nor U17756 (N_17756,N_14764,N_13338);
or U17757 (N_17757,N_13946,N_13356);
nor U17758 (N_17758,N_14870,N_13760);
xor U17759 (N_17759,N_13445,N_15021);
or U17760 (N_17760,N_12793,N_14211);
nor U17761 (N_17761,N_13827,N_13457);
and U17762 (N_17762,N_15228,N_12903);
and U17763 (N_17763,N_14303,N_15279);
nand U17764 (N_17764,N_12530,N_13673);
and U17765 (N_17765,N_14332,N_13067);
nand U17766 (N_17766,N_13038,N_15451);
nor U17767 (N_17767,N_13121,N_15335);
nor U17768 (N_17768,N_14810,N_15312);
and U17769 (N_17769,N_15422,N_14827);
nand U17770 (N_17770,N_15073,N_12531);
nand U17771 (N_17771,N_14246,N_13985);
nor U17772 (N_17772,N_13033,N_14285);
and U17773 (N_17773,N_13669,N_13401);
nor U17774 (N_17774,N_14627,N_13257);
or U17775 (N_17775,N_14878,N_15157);
or U17776 (N_17776,N_13370,N_13433);
nor U17777 (N_17777,N_15086,N_15056);
xnor U17778 (N_17778,N_13065,N_15126);
or U17779 (N_17779,N_13739,N_13788);
xnor U17780 (N_17780,N_15222,N_12610);
or U17781 (N_17781,N_13815,N_14257);
and U17782 (N_17782,N_13898,N_15137);
and U17783 (N_17783,N_13558,N_12613);
nor U17784 (N_17784,N_14643,N_12768);
nand U17785 (N_17785,N_14723,N_12681);
nand U17786 (N_17786,N_15204,N_14729);
or U17787 (N_17787,N_14558,N_14407);
or U17788 (N_17788,N_14576,N_15157);
or U17789 (N_17789,N_13310,N_14988);
and U17790 (N_17790,N_12843,N_13729);
nand U17791 (N_17791,N_13359,N_14273);
or U17792 (N_17792,N_12964,N_15376);
and U17793 (N_17793,N_14977,N_15487);
and U17794 (N_17794,N_13894,N_15538);
nand U17795 (N_17795,N_15315,N_14829);
or U17796 (N_17796,N_14737,N_15412);
nand U17797 (N_17797,N_12794,N_14479);
nor U17798 (N_17798,N_15115,N_13007);
nor U17799 (N_17799,N_14226,N_14795);
and U17800 (N_17800,N_14428,N_15051);
and U17801 (N_17801,N_15004,N_15609);
or U17802 (N_17802,N_15387,N_15536);
nor U17803 (N_17803,N_15623,N_13953);
nand U17804 (N_17804,N_15596,N_12508);
nor U17805 (N_17805,N_13992,N_14165);
nand U17806 (N_17806,N_14614,N_12827);
nor U17807 (N_17807,N_14564,N_15308);
or U17808 (N_17808,N_13657,N_14002);
or U17809 (N_17809,N_13288,N_13215);
nand U17810 (N_17810,N_14888,N_13629);
and U17811 (N_17811,N_15147,N_14377);
nor U17812 (N_17812,N_12990,N_12595);
or U17813 (N_17813,N_12867,N_14717);
or U17814 (N_17814,N_14715,N_13187);
nand U17815 (N_17815,N_14946,N_14131);
or U17816 (N_17816,N_13133,N_14403);
and U17817 (N_17817,N_15070,N_13530);
nor U17818 (N_17818,N_14386,N_13022);
nor U17819 (N_17819,N_15169,N_15071);
nor U17820 (N_17820,N_14407,N_12501);
xor U17821 (N_17821,N_14691,N_14455);
or U17822 (N_17822,N_14858,N_12535);
nand U17823 (N_17823,N_13417,N_12604);
nand U17824 (N_17824,N_13019,N_15435);
and U17825 (N_17825,N_13672,N_14226);
xor U17826 (N_17826,N_14993,N_15426);
or U17827 (N_17827,N_15307,N_14493);
or U17828 (N_17828,N_13792,N_15003);
and U17829 (N_17829,N_13189,N_12787);
xor U17830 (N_17830,N_14174,N_14832);
nor U17831 (N_17831,N_12649,N_13245);
or U17832 (N_17832,N_13321,N_13536);
and U17833 (N_17833,N_13336,N_14163);
or U17834 (N_17834,N_14224,N_12568);
or U17835 (N_17835,N_13520,N_12530);
xnor U17836 (N_17836,N_14326,N_13362);
and U17837 (N_17837,N_14752,N_12520);
nor U17838 (N_17838,N_13579,N_12791);
xor U17839 (N_17839,N_12711,N_14137);
nor U17840 (N_17840,N_13071,N_13744);
nor U17841 (N_17841,N_14219,N_15450);
xnor U17842 (N_17842,N_12547,N_14710);
nand U17843 (N_17843,N_15350,N_15548);
and U17844 (N_17844,N_12926,N_15350);
or U17845 (N_17845,N_13225,N_15088);
or U17846 (N_17846,N_15251,N_13314);
and U17847 (N_17847,N_13637,N_13977);
nand U17848 (N_17848,N_15551,N_13738);
and U17849 (N_17849,N_14884,N_14827);
and U17850 (N_17850,N_13271,N_13683);
or U17851 (N_17851,N_13808,N_13928);
and U17852 (N_17852,N_14560,N_13476);
xnor U17853 (N_17853,N_13026,N_13295);
xnor U17854 (N_17854,N_14902,N_12710);
xnor U17855 (N_17855,N_14860,N_14672);
nand U17856 (N_17856,N_14579,N_14477);
or U17857 (N_17857,N_13471,N_14135);
xor U17858 (N_17858,N_14541,N_12513);
and U17859 (N_17859,N_14305,N_14079);
nor U17860 (N_17860,N_13797,N_15521);
or U17861 (N_17861,N_15012,N_14316);
and U17862 (N_17862,N_14274,N_14252);
or U17863 (N_17863,N_15323,N_13366);
xor U17864 (N_17864,N_15322,N_13335);
xnor U17865 (N_17865,N_14232,N_14713);
or U17866 (N_17866,N_15520,N_15208);
nor U17867 (N_17867,N_13051,N_15415);
xnor U17868 (N_17868,N_13866,N_15200);
nand U17869 (N_17869,N_14507,N_14272);
or U17870 (N_17870,N_14566,N_13062);
and U17871 (N_17871,N_14448,N_15351);
nand U17872 (N_17872,N_13042,N_13402);
or U17873 (N_17873,N_14690,N_13716);
and U17874 (N_17874,N_13873,N_13251);
or U17875 (N_17875,N_14333,N_14056);
nor U17876 (N_17876,N_13594,N_13337);
or U17877 (N_17877,N_13124,N_12890);
nand U17878 (N_17878,N_12617,N_15106);
and U17879 (N_17879,N_14516,N_14808);
xor U17880 (N_17880,N_15128,N_14392);
nand U17881 (N_17881,N_14984,N_15064);
nand U17882 (N_17882,N_12521,N_15020);
nand U17883 (N_17883,N_12857,N_14548);
nand U17884 (N_17884,N_13903,N_15285);
nor U17885 (N_17885,N_14840,N_14001);
nor U17886 (N_17886,N_14283,N_14416);
xor U17887 (N_17887,N_12808,N_15108);
nand U17888 (N_17888,N_14896,N_13795);
xor U17889 (N_17889,N_15185,N_14858);
nor U17890 (N_17890,N_14718,N_15609);
or U17891 (N_17891,N_13545,N_15455);
xnor U17892 (N_17892,N_14083,N_15256);
xor U17893 (N_17893,N_13326,N_14812);
or U17894 (N_17894,N_14251,N_13860);
nand U17895 (N_17895,N_15556,N_14017);
and U17896 (N_17896,N_12631,N_12853);
or U17897 (N_17897,N_14552,N_12569);
nand U17898 (N_17898,N_13532,N_12905);
and U17899 (N_17899,N_13643,N_12818);
nand U17900 (N_17900,N_14539,N_14858);
nand U17901 (N_17901,N_15429,N_14618);
or U17902 (N_17902,N_12799,N_15262);
nor U17903 (N_17903,N_14862,N_12717);
nor U17904 (N_17904,N_12783,N_15169);
nor U17905 (N_17905,N_14395,N_12982);
nand U17906 (N_17906,N_13995,N_14811);
and U17907 (N_17907,N_15216,N_13519);
xor U17908 (N_17908,N_15367,N_13702);
nand U17909 (N_17909,N_15199,N_14898);
nor U17910 (N_17910,N_13094,N_12857);
or U17911 (N_17911,N_13879,N_13848);
or U17912 (N_17912,N_14918,N_15140);
nor U17913 (N_17913,N_14388,N_14551);
nor U17914 (N_17914,N_14605,N_12930);
or U17915 (N_17915,N_13895,N_13501);
nor U17916 (N_17916,N_14388,N_15514);
and U17917 (N_17917,N_12985,N_15130);
or U17918 (N_17918,N_14315,N_15532);
or U17919 (N_17919,N_13359,N_15542);
nand U17920 (N_17920,N_12987,N_14918);
xnor U17921 (N_17921,N_13614,N_15450);
nand U17922 (N_17922,N_15195,N_13379);
nand U17923 (N_17923,N_14576,N_14209);
nor U17924 (N_17924,N_14420,N_12822);
or U17925 (N_17925,N_13917,N_15285);
nand U17926 (N_17926,N_15196,N_13725);
and U17927 (N_17927,N_14427,N_13214);
and U17928 (N_17928,N_13360,N_14022);
nor U17929 (N_17929,N_15474,N_15242);
nand U17930 (N_17930,N_14567,N_14134);
and U17931 (N_17931,N_12757,N_14251);
or U17932 (N_17932,N_13130,N_14032);
nand U17933 (N_17933,N_14003,N_12763);
or U17934 (N_17934,N_14844,N_14256);
xor U17935 (N_17935,N_13726,N_15217);
or U17936 (N_17936,N_13536,N_13055);
nand U17937 (N_17937,N_13882,N_14904);
nand U17938 (N_17938,N_14405,N_15334);
or U17939 (N_17939,N_14726,N_13973);
nor U17940 (N_17940,N_13139,N_13256);
or U17941 (N_17941,N_14071,N_12609);
nor U17942 (N_17942,N_14072,N_12551);
nor U17943 (N_17943,N_12767,N_14161);
nand U17944 (N_17944,N_14490,N_14814);
nand U17945 (N_17945,N_12871,N_12611);
nor U17946 (N_17946,N_15576,N_14122);
or U17947 (N_17947,N_12634,N_15003);
nand U17948 (N_17948,N_14235,N_14949);
and U17949 (N_17949,N_13394,N_15127);
and U17950 (N_17950,N_13609,N_15014);
and U17951 (N_17951,N_14697,N_14156);
nor U17952 (N_17952,N_15286,N_14403);
nor U17953 (N_17953,N_15318,N_14870);
xnor U17954 (N_17954,N_13575,N_15207);
xnor U17955 (N_17955,N_15299,N_13848);
or U17956 (N_17956,N_15174,N_12559);
nand U17957 (N_17957,N_12757,N_14866);
or U17958 (N_17958,N_12504,N_12929);
and U17959 (N_17959,N_14461,N_13432);
nand U17960 (N_17960,N_13741,N_13241);
or U17961 (N_17961,N_14649,N_13398);
or U17962 (N_17962,N_13210,N_14377);
nand U17963 (N_17963,N_14527,N_13666);
nor U17964 (N_17964,N_12655,N_13000);
and U17965 (N_17965,N_13153,N_14303);
and U17966 (N_17966,N_12627,N_13493);
or U17967 (N_17967,N_15315,N_12548);
nor U17968 (N_17968,N_15175,N_12657);
or U17969 (N_17969,N_15064,N_15262);
nor U17970 (N_17970,N_15528,N_15187);
or U17971 (N_17971,N_13606,N_15166);
nand U17972 (N_17972,N_14020,N_12692);
nor U17973 (N_17973,N_14427,N_14314);
and U17974 (N_17974,N_15003,N_14757);
nand U17975 (N_17975,N_15286,N_13691);
nand U17976 (N_17976,N_12697,N_15401);
and U17977 (N_17977,N_12615,N_12790);
or U17978 (N_17978,N_12817,N_15186);
xor U17979 (N_17979,N_15537,N_14416);
nand U17980 (N_17980,N_13494,N_15013);
and U17981 (N_17981,N_14359,N_14262);
nand U17982 (N_17982,N_14995,N_15373);
or U17983 (N_17983,N_13535,N_12899);
nand U17984 (N_17984,N_15140,N_13433);
and U17985 (N_17985,N_13677,N_15195);
or U17986 (N_17986,N_15258,N_13390);
or U17987 (N_17987,N_15526,N_12747);
xnor U17988 (N_17988,N_13327,N_15481);
or U17989 (N_17989,N_14848,N_14845);
and U17990 (N_17990,N_15115,N_12634);
nand U17991 (N_17991,N_14871,N_14425);
or U17992 (N_17992,N_13181,N_15561);
nand U17993 (N_17993,N_14852,N_13624);
or U17994 (N_17994,N_14059,N_14717);
and U17995 (N_17995,N_13708,N_13333);
or U17996 (N_17996,N_14961,N_14025);
and U17997 (N_17997,N_15298,N_14319);
or U17998 (N_17998,N_13845,N_14264);
and U17999 (N_17999,N_13814,N_15000);
nor U18000 (N_18000,N_12959,N_13590);
and U18001 (N_18001,N_13382,N_14437);
nand U18002 (N_18002,N_14112,N_13459);
nand U18003 (N_18003,N_14047,N_14663);
nand U18004 (N_18004,N_14220,N_12843);
nand U18005 (N_18005,N_15330,N_12512);
nor U18006 (N_18006,N_14375,N_15483);
nand U18007 (N_18007,N_15216,N_12807);
and U18008 (N_18008,N_15115,N_12740);
xor U18009 (N_18009,N_13624,N_12680);
xor U18010 (N_18010,N_14292,N_12818);
or U18011 (N_18011,N_14263,N_13862);
nor U18012 (N_18012,N_12971,N_13214);
nand U18013 (N_18013,N_15458,N_13651);
and U18014 (N_18014,N_13994,N_14334);
nor U18015 (N_18015,N_15233,N_14370);
nor U18016 (N_18016,N_13257,N_14819);
or U18017 (N_18017,N_13447,N_14614);
xor U18018 (N_18018,N_12533,N_14669);
nand U18019 (N_18019,N_15605,N_12670);
xnor U18020 (N_18020,N_15201,N_12693);
or U18021 (N_18021,N_13186,N_13459);
or U18022 (N_18022,N_12565,N_14381);
or U18023 (N_18023,N_15090,N_13096);
or U18024 (N_18024,N_13336,N_14774);
and U18025 (N_18025,N_15027,N_14677);
or U18026 (N_18026,N_14658,N_15138);
nand U18027 (N_18027,N_13996,N_13607);
and U18028 (N_18028,N_14894,N_12906);
xnor U18029 (N_18029,N_14575,N_13442);
and U18030 (N_18030,N_14884,N_12888);
or U18031 (N_18031,N_13014,N_12980);
nor U18032 (N_18032,N_15017,N_15320);
or U18033 (N_18033,N_14248,N_13306);
and U18034 (N_18034,N_15461,N_14162);
xor U18035 (N_18035,N_12996,N_13377);
or U18036 (N_18036,N_14180,N_14183);
nand U18037 (N_18037,N_13929,N_14323);
and U18038 (N_18038,N_12820,N_12902);
and U18039 (N_18039,N_14271,N_14086);
or U18040 (N_18040,N_14156,N_15079);
nor U18041 (N_18041,N_15159,N_15360);
and U18042 (N_18042,N_13111,N_12841);
or U18043 (N_18043,N_15305,N_13904);
nand U18044 (N_18044,N_12909,N_14986);
or U18045 (N_18045,N_13596,N_14827);
nand U18046 (N_18046,N_12907,N_14707);
nand U18047 (N_18047,N_12814,N_14554);
and U18048 (N_18048,N_12687,N_15468);
nor U18049 (N_18049,N_14610,N_13267);
and U18050 (N_18050,N_13075,N_13888);
and U18051 (N_18051,N_14488,N_14569);
nor U18052 (N_18052,N_13486,N_14437);
nor U18053 (N_18053,N_13606,N_13205);
nand U18054 (N_18054,N_13291,N_14431);
xor U18055 (N_18055,N_14347,N_14921);
and U18056 (N_18056,N_13397,N_14749);
nor U18057 (N_18057,N_15495,N_13614);
nand U18058 (N_18058,N_12908,N_15508);
or U18059 (N_18059,N_14159,N_14777);
or U18060 (N_18060,N_14404,N_15218);
and U18061 (N_18061,N_12668,N_14960);
nand U18062 (N_18062,N_13478,N_13341);
and U18063 (N_18063,N_12611,N_12975);
nand U18064 (N_18064,N_14036,N_13371);
or U18065 (N_18065,N_12532,N_14038);
nand U18066 (N_18066,N_13677,N_13694);
nand U18067 (N_18067,N_15300,N_14312);
and U18068 (N_18068,N_13820,N_13842);
and U18069 (N_18069,N_13881,N_14838);
and U18070 (N_18070,N_12571,N_13274);
nor U18071 (N_18071,N_13100,N_15257);
nand U18072 (N_18072,N_13381,N_13282);
nor U18073 (N_18073,N_12703,N_14194);
and U18074 (N_18074,N_12638,N_15009);
nand U18075 (N_18075,N_14950,N_14134);
nand U18076 (N_18076,N_14193,N_13740);
or U18077 (N_18077,N_13649,N_13771);
xnor U18078 (N_18078,N_14736,N_13417);
nand U18079 (N_18079,N_13110,N_12922);
or U18080 (N_18080,N_12616,N_13164);
nor U18081 (N_18081,N_14096,N_15120);
nand U18082 (N_18082,N_14292,N_12980);
and U18083 (N_18083,N_13434,N_13558);
or U18084 (N_18084,N_13308,N_13776);
nand U18085 (N_18085,N_15432,N_14025);
and U18086 (N_18086,N_15322,N_13187);
nor U18087 (N_18087,N_13414,N_12857);
and U18088 (N_18088,N_13832,N_15305);
nand U18089 (N_18089,N_15363,N_13946);
nand U18090 (N_18090,N_14524,N_13174);
nand U18091 (N_18091,N_15041,N_14780);
and U18092 (N_18092,N_14481,N_14664);
xor U18093 (N_18093,N_13401,N_13701);
nand U18094 (N_18094,N_12707,N_13139);
xnor U18095 (N_18095,N_13056,N_15006);
nor U18096 (N_18096,N_13362,N_13318);
or U18097 (N_18097,N_13727,N_13542);
and U18098 (N_18098,N_15176,N_13163);
and U18099 (N_18099,N_15518,N_13707);
xnor U18100 (N_18100,N_14271,N_13501);
and U18101 (N_18101,N_14876,N_12875);
or U18102 (N_18102,N_12826,N_15074);
nor U18103 (N_18103,N_13581,N_15338);
and U18104 (N_18104,N_13624,N_14192);
nor U18105 (N_18105,N_13780,N_15027);
or U18106 (N_18106,N_12970,N_14813);
and U18107 (N_18107,N_12992,N_14701);
nand U18108 (N_18108,N_12737,N_14509);
or U18109 (N_18109,N_13142,N_13512);
or U18110 (N_18110,N_15186,N_15240);
xnor U18111 (N_18111,N_13215,N_15219);
or U18112 (N_18112,N_13433,N_14118);
and U18113 (N_18113,N_14828,N_13785);
nor U18114 (N_18114,N_15296,N_14127);
or U18115 (N_18115,N_15440,N_15170);
or U18116 (N_18116,N_15413,N_14667);
nor U18117 (N_18117,N_14123,N_14455);
xor U18118 (N_18118,N_12548,N_15557);
and U18119 (N_18119,N_13251,N_13953);
or U18120 (N_18120,N_13239,N_15269);
and U18121 (N_18121,N_13910,N_14568);
and U18122 (N_18122,N_13275,N_13918);
nor U18123 (N_18123,N_13096,N_14105);
nor U18124 (N_18124,N_14310,N_12553);
and U18125 (N_18125,N_14656,N_13844);
nor U18126 (N_18126,N_15173,N_14482);
and U18127 (N_18127,N_14237,N_14239);
and U18128 (N_18128,N_14288,N_13959);
xor U18129 (N_18129,N_14017,N_15511);
nor U18130 (N_18130,N_15619,N_13498);
nor U18131 (N_18131,N_14424,N_14873);
nor U18132 (N_18132,N_13004,N_12572);
xnor U18133 (N_18133,N_12830,N_13366);
nor U18134 (N_18134,N_15460,N_14744);
nand U18135 (N_18135,N_15569,N_14293);
and U18136 (N_18136,N_12983,N_15321);
nor U18137 (N_18137,N_13766,N_13555);
or U18138 (N_18138,N_14268,N_12850);
nor U18139 (N_18139,N_13187,N_14173);
and U18140 (N_18140,N_15096,N_12610);
or U18141 (N_18141,N_15077,N_14602);
and U18142 (N_18142,N_13442,N_14868);
and U18143 (N_18143,N_12912,N_13757);
nor U18144 (N_18144,N_15145,N_12591);
or U18145 (N_18145,N_14704,N_12761);
nand U18146 (N_18146,N_15580,N_13261);
xor U18147 (N_18147,N_14060,N_13822);
nor U18148 (N_18148,N_14235,N_13156);
nand U18149 (N_18149,N_14347,N_14085);
and U18150 (N_18150,N_14132,N_12677);
nand U18151 (N_18151,N_15481,N_14071);
and U18152 (N_18152,N_15326,N_14171);
or U18153 (N_18153,N_13421,N_14913);
or U18154 (N_18154,N_14546,N_15377);
or U18155 (N_18155,N_12779,N_14098);
nand U18156 (N_18156,N_14945,N_15268);
nand U18157 (N_18157,N_12794,N_12545);
nor U18158 (N_18158,N_14128,N_13087);
nor U18159 (N_18159,N_14945,N_13953);
or U18160 (N_18160,N_13396,N_13011);
nand U18161 (N_18161,N_12666,N_14035);
or U18162 (N_18162,N_12898,N_14673);
nand U18163 (N_18163,N_15385,N_12833);
or U18164 (N_18164,N_14045,N_14003);
or U18165 (N_18165,N_15043,N_14285);
or U18166 (N_18166,N_15514,N_15118);
nand U18167 (N_18167,N_13969,N_15300);
or U18168 (N_18168,N_14324,N_15340);
xnor U18169 (N_18169,N_13912,N_15199);
nand U18170 (N_18170,N_15144,N_14402);
nor U18171 (N_18171,N_12779,N_14031);
nand U18172 (N_18172,N_15292,N_13568);
xnor U18173 (N_18173,N_14300,N_15497);
and U18174 (N_18174,N_15199,N_14565);
or U18175 (N_18175,N_15225,N_14345);
nor U18176 (N_18176,N_15566,N_12765);
or U18177 (N_18177,N_15123,N_13222);
and U18178 (N_18178,N_13824,N_14500);
nor U18179 (N_18179,N_13555,N_15365);
nand U18180 (N_18180,N_12909,N_13271);
or U18181 (N_18181,N_15072,N_12559);
or U18182 (N_18182,N_12919,N_15426);
nand U18183 (N_18183,N_15193,N_13019);
and U18184 (N_18184,N_12508,N_15571);
or U18185 (N_18185,N_12877,N_14281);
or U18186 (N_18186,N_13359,N_13019);
and U18187 (N_18187,N_13241,N_13561);
xnor U18188 (N_18188,N_14589,N_13588);
xor U18189 (N_18189,N_13133,N_15425);
or U18190 (N_18190,N_13315,N_14994);
and U18191 (N_18191,N_15447,N_13497);
xor U18192 (N_18192,N_13631,N_13496);
nor U18193 (N_18193,N_14761,N_15344);
or U18194 (N_18194,N_13214,N_13502);
nor U18195 (N_18195,N_13825,N_13638);
nor U18196 (N_18196,N_13361,N_13123);
or U18197 (N_18197,N_12732,N_13853);
and U18198 (N_18198,N_12933,N_13270);
or U18199 (N_18199,N_13984,N_13680);
or U18200 (N_18200,N_13958,N_13489);
or U18201 (N_18201,N_13338,N_15437);
nor U18202 (N_18202,N_14545,N_12881);
or U18203 (N_18203,N_12877,N_13227);
nand U18204 (N_18204,N_13899,N_14465);
nor U18205 (N_18205,N_13647,N_13489);
nor U18206 (N_18206,N_14470,N_13585);
nor U18207 (N_18207,N_13148,N_14703);
and U18208 (N_18208,N_14130,N_14344);
nor U18209 (N_18209,N_15397,N_13311);
xor U18210 (N_18210,N_15454,N_15618);
or U18211 (N_18211,N_13818,N_14870);
nand U18212 (N_18212,N_13449,N_15453);
xnor U18213 (N_18213,N_14784,N_14409);
nor U18214 (N_18214,N_13156,N_14107);
xor U18215 (N_18215,N_13337,N_15207);
nand U18216 (N_18216,N_13253,N_14697);
nor U18217 (N_18217,N_15465,N_14615);
or U18218 (N_18218,N_14026,N_13351);
nand U18219 (N_18219,N_12734,N_13914);
nor U18220 (N_18220,N_12563,N_12690);
nand U18221 (N_18221,N_15216,N_14477);
or U18222 (N_18222,N_14491,N_13323);
nand U18223 (N_18223,N_12786,N_14296);
xor U18224 (N_18224,N_14687,N_12844);
xnor U18225 (N_18225,N_14133,N_13735);
and U18226 (N_18226,N_13053,N_13269);
or U18227 (N_18227,N_12523,N_13844);
or U18228 (N_18228,N_15541,N_13334);
or U18229 (N_18229,N_13503,N_14578);
and U18230 (N_18230,N_15112,N_15491);
and U18231 (N_18231,N_12716,N_12874);
or U18232 (N_18232,N_13745,N_13962);
or U18233 (N_18233,N_12703,N_15523);
and U18234 (N_18234,N_14928,N_14458);
and U18235 (N_18235,N_12673,N_13180);
nor U18236 (N_18236,N_13074,N_13733);
nor U18237 (N_18237,N_14268,N_12725);
xnor U18238 (N_18238,N_12619,N_12933);
nand U18239 (N_18239,N_15397,N_14731);
nand U18240 (N_18240,N_14985,N_14642);
and U18241 (N_18241,N_12850,N_13234);
nand U18242 (N_18242,N_15408,N_14396);
nand U18243 (N_18243,N_12936,N_13017);
nand U18244 (N_18244,N_14215,N_13221);
and U18245 (N_18245,N_14065,N_14472);
or U18246 (N_18246,N_14757,N_14664);
nand U18247 (N_18247,N_13315,N_14440);
nand U18248 (N_18248,N_12712,N_12798);
xnor U18249 (N_18249,N_14946,N_13210);
or U18250 (N_18250,N_13294,N_12636);
xor U18251 (N_18251,N_15433,N_13941);
or U18252 (N_18252,N_14345,N_13341);
xnor U18253 (N_18253,N_13416,N_13825);
nand U18254 (N_18254,N_12837,N_13336);
or U18255 (N_18255,N_13892,N_14276);
and U18256 (N_18256,N_12996,N_13933);
and U18257 (N_18257,N_12663,N_13716);
nand U18258 (N_18258,N_14904,N_15010);
nand U18259 (N_18259,N_12619,N_12826);
and U18260 (N_18260,N_13605,N_15104);
and U18261 (N_18261,N_14014,N_14859);
nor U18262 (N_18262,N_13781,N_15281);
nand U18263 (N_18263,N_14390,N_14098);
or U18264 (N_18264,N_12665,N_14388);
nor U18265 (N_18265,N_14413,N_13898);
and U18266 (N_18266,N_15010,N_15425);
and U18267 (N_18267,N_13983,N_13829);
nand U18268 (N_18268,N_13934,N_15271);
nand U18269 (N_18269,N_14191,N_15183);
or U18270 (N_18270,N_12848,N_15420);
nor U18271 (N_18271,N_12827,N_13628);
xnor U18272 (N_18272,N_14855,N_12806);
xor U18273 (N_18273,N_12597,N_13299);
and U18274 (N_18274,N_13345,N_13778);
xnor U18275 (N_18275,N_14408,N_15616);
and U18276 (N_18276,N_15222,N_15552);
nand U18277 (N_18277,N_14183,N_13615);
nand U18278 (N_18278,N_15231,N_15269);
nand U18279 (N_18279,N_15528,N_13677);
nand U18280 (N_18280,N_14195,N_13177);
nand U18281 (N_18281,N_14997,N_14612);
and U18282 (N_18282,N_14621,N_13155);
nand U18283 (N_18283,N_14393,N_12566);
xnor U18284 (N_18284,N_14957,N_15390);
and U18285 (N_18285,N_15517,N_15521);
or U18286 (N_18286,N_13411,N_14437);
or U18287 (N_18287,N_12518,N_15621);
or U18288 (N_18288,N_13243,N_15146);
xor U18289 (N_18289,N_14664,N_13471);
and U18290 (N_18290,N_13756,N_13223);
nor U18291 (N_18291,N_13814,N_13978);
nand U18292 (N_18292,N_13903,N_14315);
nand U18293 (N_18293,N_13154,N_13234);
nand U18294 (N_18294,N_13506,N_13315);
and U18295 (N_18295,N_13711,N_13355);
nor U18296 (N_18296,N_13130,N_15420);
xor U18297 (N_18297,N_12812,N_12705);
xor U18298 (N_18298,N_14766,N_15269);
xnor U18299 (N_18299,N_14460,N_15620);
nor U18300 (N_18300,N_15398,N_13245);
xor U18301 (N_18301,N_15253,N_14847);
or U18302 (N_18302,N_13113,N_13433);
nand U18303 (N_18303,N_15370,N_13610);
and U18304 (N_18304,N_12941,N_13897);
and U18305 (N_18305,N_13217,N_15469);
nand U18306 (N_18306,N_14270,N_12788);
and U18307 (N_18307,N_15588,N_14400);
nand U18308 (N_18308,N_13266,N_13332);
or U18309 (N_18309,N_12895,N_14667);
nor U18310 (N_18310,N_12536,N_12677);
and U18311 (N_18311,N_13288,N_13531);
or U18312 (N_18312,N_13825,N_13839);
and U18313 (N_18313,N_14295,N_14154);
nor U18314 (N_18314,N_14092,N_15473);
or U18315 (N_18315,N_12558,N_14518);
and U18316 (N_18316,N_12627,N_13459);
nand U18317 (N_18317,N_15077,N_14975);
xor U18318 (N_18318,N_14408,N_13538);
nor U18319 (N_18319,N_15383,N_12767);
nand U18320 (N_18320,N_13532,N_14393);
nand U18321 (N_18321,N_15081,N_15284);
nor U18322 (N_18322,N_13366,N_13710);
xnor U18323 (N_18323,N_14250,N_15052);
and U18324 (N_18324,N_13253,N_14780);
and U18325 (N_18325,N_14234,N_12913);
and U18326 (N_18326,N_13709,N_14359);
nand U18327 (N_18327,N_14080,N_14241);
nand U18328 (N_18328,N_12905,N_13188);
nand U18329 (N_18329,N_13492,N_14103);
nand U18330 (N_18330,N_13591,N_12504);
or U18331 (N_18331,N_14318,N_13707);
or U18332 (N_18332,N_15469,N_14065);
nand U18333 (N_18333,N_15536,N_12861);
nand U18334 (N_18334,N_13952,N_13360);
nand U18335 (N_18335,N_12658,N_12675);
xnor U18336 (N_18336,N_13182,N_13271);
xnor U18337 (N_18337,N_15567,N_14380);
or U18338 (N_18338,N_14894,N_13284);
nor U18339 (N_18339,N_13980,N_13546);
xor U18340 (N_18340,N_15261,N_12930);
nor U18341 (N_18341,N_13927,N_15259);
nor U18342 (N_18342,N_15301,N_14858);
xor U18343 (N_18343,N_13362,N_15057);
nand U18344 (N_18344,N_13402,N_15268);
or U18345 (N_18345,N_15580,N_15491);
nand U18346 (N_18346,N_13789,N_13799);
nor U18347 (N_18347,N_15142,N_13069);
nor U18348 (N_18348,N_13104,N_15096);
and U18349 (N_18349,N_14527,N_15517);
nand U18350 (N_18350,N_14194,N_14941);
nor U18351 (N_18351,N_14538,N_12826);
nand U18352 (N_18352,N_15620,N_12678);
or U18353 (N_18353,N_13590,N_13722);
and U18354 (N_18354,N_14581,N_15611);
or U18355 (N_18355,N_15256,N_15485);
or U18356 (N_18356,N_14658,N_13244);
or U18357 (N_18357,N_12580,N_14048);
nor U18358 (N_18358,N_14760,N_13461);
and U18359 (N_18359,N_13038,N_13318);
or U18360 (N_18360,N_14934,N_14727);
and U18361 (N_18361,N_14592,N_13585);
nand U18362 (N_18362,N_14581,N_14355);
or U18363 (N_18363,N_15617,N_12643);
nand U18364 (N_18364,N_13885,N_13513);
nor U18365 (N_18365,N_13270,N_13832);
or U18366 (N_18366,N_15005,N_13295);
or U18367 (N_18367,N_14229,N_14742);
nand U18368 (N_18368,N_14621,N_15084);
nor U18369 (N_18369,N_13451,N_13237);
nor U18370 (N_18370,N_13700,N_13427);
or U18371 (N_18371,N_14267,N_14146);
and U18372 (N_18372,N_13074,N_13281);
nand U18373 (N_18373,N_12520,N_14430);
nand U18374 (N_18374,N_13445,N_13619);
and U18375 (N_18375,N_14675,N_13909);
or U18376 (N_18376,N_15177,N_13999);
nand U18377 (N_18377,N_13764,N_12993);
and U18378 (N_18378,N_13095,N_14467);
or U18379 (N_18379,N_13396,N_15292);
and U18380 (N_18380,N_13810,N_14875);
or U18381 (N_18381,N_15445,N_15006);
or U18382 (N_18382,N_14396,N_13925);
and U18383 (N_18383,N_14608,N_13254);
nand U18384 (N_18384,N_14795,N_15261);
nor U18385 (N_18385,N_13307,N_12719);
and U18386 (N_18386,N_14801,N_13408);
nand U18387 (N_18387,N_13680,N_14947);
or U18388 (N_18388,N_15404,N_12879);
or U18389 (N_18389,N_13649,N_15452);
nand U18390 (N_18390,N_15463,N_13669);
and U18391 (N_18391,N_13123,N_12929);
or U18392 (N_18392,N_12740,N_14242);
nor U18393 (N_18393,N_12712,N_13129);
and U18394 (N_18394,N_13753,N_15523);
xnor U18395 (N_18395,N_15357,N_14830);
nor U18396 (N_18396,N_13279,N_13564);
nand U18397 (N_18397,N_13762,N_14010);
nand U18398 (N_18398,N_15132,N_12825);
nor U18399 (N_18399,N_15540,N_13264);
nor U18400 (N_18400,N_12681,N_13258);
nor U18401 (N_18401,N_13406,N_14443);
or U18402 (N_18402,N_13355,N_13006);
nor U18403 (N_18403,N_14749,N_14526);
and U18404 (N_18404,N_15589,N_13981);
nor U18405 (N_18405,N_13520,N_13971);
nand U18406 (N_18406,N_13368,N_14868);
nor U18407 (N_18407,N_13781,N_13600);
nor U18408 (N_18408,N_15096,N_13001);
nand U18409 (N_18409,N_13263,N_13828);
and U18410 (N_18410,N_13613,N_15092);
nor U18411 (N_18411,N_14521,N_14188);
nand U18412 (N_18412,N_13942,N_14613);
or U18413 (N_18413,N_12752,N_15451);
or U18414 (N_18414,N_14600,N_15423);
or U18415 (N_18415,N_13192,N_14395);
nand U18416 (N_18416,N_15094,N_13526);
nor U18417 (N_18417,N_14093,N_14988);
xnor U18418 (N_18418,N_13135,N_15006);
or U18419 (N_18419,N_14586,N_12832);
nor U18420 (N_18420,N_13665,N_14898);
or U18421 (N_18421,N_15394,N_13588);
and U18422 (N_18422,N_15192,N_15096);
or U18423 (N_18423,N_14781,N_13724);
and U18424 (N_18424,N_14457,N_13002);
xor U18425 (N_18425,N_14887,N_13826);
nor U18426 (N_18426,N_14304,N_14814);
nor U18427 (N_18427,N_14335,N_15323);
or U18428 (N_18428,N_15103,N_15036);
nand U18429 (N_18429,N_13279,N_14400);
nor U18430 (N_18430,N_14465,N_12566);
and U18431 (N_18431,N_14023,N_14201);
nand U18432 (N_18432,N_13700,N_13346);
nor U18433 (N_18433,N_15398,N_14349);
or U18434 (N_18434,N_14775,N_14397);
nor U18435 (N_18435,N_13147,N_14739);
xor U18436 (N_18436,N_14267,N_15103);
nor U18437 (N_18437,N_13759,N_13399);
nor U18438 (N_18438,N_14109,N_12853);
and U18439 (N_18439,N_13598,N_15220);
or U18440 (N_18440,N_13233,N_13213);
and U18441 (N_18441,N_13530,N_14782);
or U18442 (N_18442,N_15399,N_15446);
nand U18443 (N_18443,N_14770,N_15583);
nand U18444 (N_18444,N_14654,N_15299);
and U18445 (N_18445,N_14870,N_15279);
or U18446 (N_18446,N_13221,N_15325);
or U18447 (N_18447,N_13645,N_14198);
nand U18448 (N_18448,N_15097,N_14964);
or U18449 (N_18449,N_14770,N_15387);
nor U18450 (N_18450,N_14980,N_15034);
and U18451 (N_18451,N_12878,N_13971);
nand U18452 (N_18452,N_12632,N_13961);
nor U18453 (N_18453,N_14018,N_15057);
or U18454 (N_18454,N_14483,N_13329);
or U18455 (N_18455,N_15005,N_14500);
and U18456 (N_18456,N_13106,N_12563);
xnor U18457 (N_18457,N_12857,N_14449);
nor U18458 (N_18458,N_12728,N_15496);
nand U18459 (N_18459,N_12512,N_14264);
and U18460 (N_18460,N_13953,N_13484);
and U18461 (N_18461,N_13886,N_13619);
nand U18462 (N_18462,N_13733,N_15259);
or U18463 (N_18463,N_12617,N_15443);
and U18464 (N_18464,N_15036,N_14944);
nor U18465 (N_18465,N_15136,N_13082);
nand U18466 (N_18466,N_14488,N_13028);
xnor U18467 (N_18467,N_12576,N_13688);
and U18468 (N_18468,N_15463,N_15107);
or U18469 (N_18469,N_14107,N_14812);
and U18470 (N_18470,N_12814,N_15102);
and U18471 (N_18471,N_12677,N_14579);
or U18472 (N_18472,N_14057,N_13234);
or U18473 (N_18473,N_13706,N_14746);
or U18474 (N_18474,N_13210,N_15604);
nand U18475 (N_18475,N_15131,N_14957);
and U18476 (N_18476,N_14219,N_13066);
xor U18477 (N_18477,N_15367,N_14392);
and U18478 (N_18478,N_15615,N_13210);
nor U18479 (N_18479,N_13030,N_12660);
nor U18480 (N_18480,N_14317,N_12983);
nor U18481 (N_18481,N_15597,N_14752);
nand U18482 (N_18482,N_13027,N_14279);
nand U18483 (N_18483,N_14872,N_14603);
or U18484 (N_18484,N_12860,N_13799);
and U18485 (N_18485,N_12985,N_13454);
and U18486 (N_18486,N_12860,N_12690);
nor U18487 (N_18487,N_13705,N_13753);
and U18488 (N_18488,N_15178,N_14563);
nor U18489 (N_18489,N_14869,N_12857);
nor U18490 (N_18490,N_13472,N_14909);
nor U18491 (N_18491,N_15141,N_14742);
nor U18492 (N_18492,N_13069,N_13249);
and U18493 (N_18493,N_13792,N_14790);
and U18494 (N_18494,N_13845,N_14813);
xor U18495 (N_18495,N_14235,N_15468);
or U18496 (N_18496,N_13275,N_14112);
xnor U18497 (N_18497,N_12984,N_13205);
and U18498 (N_18498,N_15339,N_13956);
or U18499 (N_18499,N_13051,N_13665);
and U18500 (N_18500,N_12559,N_15327);
nor U18501 (N_18501,N_13240,N_14522);
or U18502 (N_18502,N_15131,N_12662);
or U18503 (N_18503,N_14435,N_13522);
xnor U18504 (N_18504,N_12811,N_14758);
and U18505 (N_18505,N_15320,N_14681);
nand U18506 (N_18506,N_14085,N_13248);
nand U18507 (N_18507,N_13097,N_12891);
or U18508 (N_18508,N_15073,N_14940);
and U18509 (N_18509,N_13345,N_13261);
and U18510 (N_18510,N_14418,N_13484);
and U18511 (N_18511,N_15448,N_14974);
or U18512 (N_18512,N_14018,N_14228);
or U18513 (N_18513,N_14691,N_15470);
and U18514 (N_18514,N_13240,N_13785);
nor U18515 (N_18515,N_12665,N_14193);
xor U18516 (N_18516,N_15555,N_14528);
nand U18517 (N_18517,N_13186,N_14378);
nor U18518 (N_18518,N_13890,N_13977);
and U18519 (N_18519,N_13033,N_13587);
and U18520 (N_18520,N_14537,N_13633);
and U18521 (N_18521,N_13438,N_14293);
or U18522 (N_18522,N_13712,N_15577);
xor U18523 (N_18523,N_14416,N_14897);
or U18524 (N_18524,N_14979,N_14590);
and U18525 (N_18525,N_15154,N_14103);
nor U18526 (N_18526,N_14246,N_15372);
and U18527 (N_18527,N_13429,N_14105);
and U18528 (N_18528,N_14206,N_15562);
and U18529 (N_18529,N_13386,N_13529);
and U18530 (N_18530,N_15101,N_14949);
or U18531 (N_18531,N_14579,N_13758);
nand U18532 (N_18532,N_13539,N_14493);
or U18533 (N_18533,N_12738,N_15541);
nor U18534 (N_18534,N_13410,N_12929);
nand U18535 (N_18535,N_12583,N_13983);
and U18536 (N_18536,N_15453,N_14322);
or U18537 (N_18537,N_12758,N_15100);
and U18538 (N_18538,N_14499,N_15024);
or U18539 (N_18539,N_13310,N_13035);
and U18540 (N_18540,N_15505,N_14695);
or U18541 (N_18541,N_13698,N_13852);
nand U18542 (N_18542,N_14903,N_12980);
and U18543 (N_18543,N_15001,N_14605);
and U18544 (N_18544,N_14590,N_14401);
or U18545 (N_18545,N_13245,N_14108);
nand U18546 (N_18546,N_14137,N_14381);
and U18547 (N_18547,N_14172,N_13832);
and U18548 (N_18548,N_15455,N_15272);
or U18549 (N_18549,N_14404,N_13222);
and U18550 (N_18550,N_14943,N_14872);
or U18551 (N_18551,N_14901,N_14973);
or U18552 (N_18552,N_12934,N_13285);
and U18553 (N_18553,N_12897,N_13310);
nor U18554 (N_18554,N_14059,N_13594);
and U18555 (N_18555,N_12877,N_15043);
nor U18556 (N_18556,N_12806,N_15197);
nor U18557 (N_18557,N_13891,N_14468);
or U18558 (N_18558,N_14948,N_14568);
and U18559 (N_18559,N_15189,N_13336);
or U18560 (N_18560,N_13706,N_13635);
nand U18561 (N_18561,N_12967,N_13642);
and U18562 (N_18562,N_13108,N_15162);
xor U18563 (N_18563,N_13126,N_12526);
or U18564 (N_18564,N_14917,N_14483);
nand U18565 (N_18565,N_13574,N_13201);
nand U18566 (N_18566,N_12668,N_14463);
nand U18567 (N_18567,N_13313,N_12872);
and U18568 (N_18568,N_15227,N_14898);
nor U18569 (N_18569,N_15440,N_13438);
nand U18570 (N_18570,N_12814,N_13842);
or U18571 (N_18571,N_14018,N_13699);
nand U18572 (N_18572,N_12981,N_14904);
nor U18573 (N_18573,N_15207,N_12812);
nand U18574 (N_18574,N_14123,N_15010);
or U18575 (N_18575,N_14604,N_13636);
and U18576 (N_18576,N_13512,N_15378);
nand U18577 (N_18577,N_12660,N_12612);
xor U18578 (N_18578,N_15558,N_13359);
xnor U18579 (N_18579,N_13257,N_13724);
nor U18580 (N_18580,N_14298,N_14214);
or U18581 (N_18581,N_14607,N_14446);
nor U18582 (N_18582,N_13449,N_15086);
or U18583 (N_18583,N_13756,N_14780);
nor U18584 (N_18584,N_13768,N_14615);
and U18585 (N_18585,N_14956,N_13218);
and U18586 (N_18586,N_13760,N_13694);
or U18587 (N_18587,N_14930,N_12525);
xnor U18588 (N_18588,N_12777,N_12913);
nor U18589 (N_18589,N_13049,N_14208);
or U18590 (N_18590,N_13678,N_13710);
and U18591 (N_18591,N_13448,N_13318);
or U18592 (N_18592,N_13324,N_15609);
or U18593 (N_18593,N_13482,N_15563);
or U18594 (N_18594,N_14204,N_13729);
and U18595 (N_18595,N_15212,N_12739);
xor U18596 (N_18596,N_14554,N_14190);
and U18597 (N_18597,N_15125,N_13651);
nor U18598 (N_18598,N_14352,N_13613);
nor U18599 (N_18599,N_14870,N_15352);
or U18600 (N_18600,N_14332,N_12508);
nand U18601 (N_18601,N_13878,N_14385);
nor U18602 (N_18602,N_15363,N_15083);
nand U18603 (N_18603,N_12836,N_14464);
xnor U18604 (N_18604,N_13577,N_13618);
nand U18605 (N_18605,N_13079,N_13578);
or U18606 (N_18606,N_13391,N_12597);
nand U18607 (N_18607,N_15019,N_14866);
or U18608 (N_18608,N_13955,N_13834);
nor U18609 (N_18609,N_13383,N_13742);
nand U18610 (N_18610,N_15018,N_13682);
and U18611 (N_18611,N_14838,N_12548);
nand U18612 (N_18612,N_13010,N_14194);
and U18613 (N_18613,N_14997,N_14210);
nand U18614 (N_18614,N_13604,N_14776);
nor U18615 (N_18615,N_13111,N_13984);
and U18616 (N_18616,N_14860,N_12839);
and U18617 (N_18617,N_15601,N_15380);
and U18618 (N_18618,N_13552,N_12566);
nand U18619 (N_18619,N_13551,N_13606);
nand U18620 (N_18620,N_14982,N_14706);
and U18621 (N_18621,N_12709,N_15083);
or U18622 (N_18622,N_13333,N_15563);
or U18623 (N_18623,N_14107,N_14851);
nand U18624 (N_18624,N_13013,N_14593);
nand U18625 (N_18625,N_13551,N_14232);
nor U18626 (N_18626,N_14900,N_15433);
or U18627 (N_18627,N_13267,N_13500);
nand U18628 (N_18628,N_14585,N_13146);
and U18629 (N_18629,N_14138,N_15120);
nand U18630 (N_18630,N_14218,N_13497);
or U18631 (N_18631,N_13002,N_13406);
xnor U18632 (N_18632,N_12728,N_13290);
and U18633 (N_18633,N_14884,N_14887);
or U18634 (N_18634,N_13345,N_12988);
or U18635 (N_18635,N_13088,N_14971);
and U18636 (N_18636,N_14767,N_12825);
xor U18637 (N_18637,N_14468,N_15156);
nand U18638 (N_18638,N_13373,N_14307);
nand U18639 (N_18639,N_14012,N_14112);
or U18640 (N_18640,N_15617,N_13410);
and U18641 (N_18641,N_12548,N_13254);
and U18642 (N_18642,N_13257,N_15362);
xnor U18643 (N_18643,N_15124,N_13746);
and U18644 (N_18644,N_14628,N_14098);
and U18645 (N_18645,N_14159,N_14950);
or U18646 (N_18646,N_14533,N_14481);
nor U18647 (N_18647,N_13518,N_14863);
nand U18648 (N_18648,N_12906,N_14246);
or U18649 (N_18649,N_13695,N_13772);
nand U18650 (N_18650,N_12649,N_13114);
xor U18651 (N_18651,N_14297,N_14332);
nor U18652 (N_18652,N_15360,N_15146);
nor U18653 (N_18653,N_14926,N_13222);
nor U18654 (N_18654,N_14248,N_14014);
and U18655 (N_18655,N_12692,N_14965);
nand U18656 (N_18656,N_12965,N_15042);
nor U18657 (N_18657,N_13529,N_14575);
and U18658 (N_18658,N_12596,N_14454);
nand U18659 (N_18659,N_13820,N_13029);
nand U18660 (N_18660,N_12834,N_12571);
or U18661 (N_18661,N_14627,N_13711);
nand U18662 (N_18662,N_14247,N_12899);
or U18663 (N_18663,N_14040,N_13879);
nand U18664 (N_18664,N_15066,N_15195);
and U18665 (N_18665,N_12657,N_15333);
nand U18666 (N_18666,N_14438,N_14834);
nor U18667 (N_18667,N_13337,N_13232);
or U18668 (N_18668,N_12841,N_13355);
nand U18669 (N_18669,N_14422,N_12881);
and U18670 (N_18670,N_14953,N_13927);
and U18671 (N_18671,N_12720,N_12919);
and U18672 (N_18672,N_14975,N_15622);
nand U18673 (N_18673,N_13766,N_14198);
or U18674 (N_18674,N_12533,N_14361);
nand U18675 (N_18675,N_14697,N_12618);
or U18676 (N_18676,N_15356,N_14965);
and U18677 (N_18677,N_15308,N_13714);
and U18678 (N_18678,N_13493,N_13543);
nand U18679 (N_18679,N_14538,N_13407);
nand U18680 (N_18680,N_14794,N_15250);
xnor U18681 (N_18681,N_14220,N_13052);
and U18682 (N_18682,N_13316,N_12616);
nor U18683 (N_18683,N_14720,N_14997);
nand U18684 (N_18684,N_13996,N_13375);
and U18685 (N_18685,N_13058,N_13665);
nand U18686 (N_18686,N_14790,N_15180);
nand U18687 (N_18687,N_14287,N_12992);
nand U18688 (N_18688,N_14935,N_13364);
nor U18689 (N_18689,N_14805,N_14975);
and U18690 (N_18690,N_13543,N_13052);
nor U18691 (N_18691,N_12718,N_14981);
nand U18692 (N_18692,N_14951,N_13403);
nor U18693 (N_18693,N_13382,N_13701);
or U18694 (N_18694,N_15033,N_14703);
nand U18695 (N_18695,N_13655,N_15617);
nor U18696 (N_18696,N_13489,N_13669);
xor U18697 (N_18697,N_13818,N_15492);
or U18698 (N_18698,N_13817,N_13348);
and U18699 (N_18699,N_12555,N_14569);
and U18700 (N_18700,N_14985,N_14311);
nand U18701 (N_18701,N_15228,N_15583);
nand U18702 (N_18702,N_12922,N_13695);
nor U18703 (N_18703,N_15426,N_13895);
or U18704 (N_18704,N_13067,N_15427);
or U18705 (N_18705,N_13769,N_14431);
and U18706 (N_18706,N_14365,N_14547);
nor U18707 (N_18707,N_13231,N_12729);
and U18708 (N_18708,N_14623,N_13427);
or U18709 (N_18709,N_12916,N_15571);
nor U18710 (N_18710,N_13201,N_14298);
or U18711 (N_18711,N_13125,N_13171);
nor U18712 (N_18712,N_15241,N_12930);
and U18713 (N_18713,N_15086,N_13296);
or U18714 (N_18714,N_13208,N_13730);
and U18715 (N_18715,N_12713,N_12619);
nand U18716 (N_18716,N_15369,N_14208);
nor U18717 (N_18717,N_14630,N_13408);
xor U18718 (N_18718,N_12592,N_14551);
or U18719 (N_18719,N_15207,N_13748);
nor U18720 (N_18720,N_14603,N_14615);
or U18721 (N_18721,N_13058,N_13185);
nor U18722 (N_18722,N_13574,N_13667);
or U18723 (N_18723,N_15109,N_14260);
nand U18724 (N_18724,N_15419,N_15404);
and U18725 (N_18725,N_12574,N_13455);
xor U18726 (N_18726,N_15016,N_14407);
nand U18727 (N_18727,N_13618,N_14126);
nor U18728 (N_18728,N_15197,N_14713);
and U18729 (N_18729,N_12548,N_13394);
or U18730 (N_18730,N_14433,N_12502);
nor U18731 (N_18731,N_14195,N_14747);
and U18732 (N_18732,N_13301,N_13402);
nand U18733 (N_18733,N_13785,N_14366);
or U18734 (N_18734,N_13824,N_13143);
or U18735 (N_18735,N_15331,N_12972);
or U18736 (N_18736,N_14196,N_15348);
xnor U18737 (N_18737,N_15583,N_15174);
nand U18738 (N_18738,N_15069,N_13825);
or U18739 (N_18739,N_12798,N_13169);
or U18740 (N_18740,N_13004,N_15593);
nand U18741 (N_18741,N_15557,N_12670);
or U18742 (N_18742,N_13806,N_14373);
or U18743 (N_18743,N_15243,N_13633);
nand U18744 (N_18744,N_14060,N_14585);
and U18745 (N_18745,N_14138,N_13426);
nand U18746 (N_18746,N_13943,N_14320);
or U18747 (N_18747,N_14992,N_13651);
nand U18748 (N_18748,N_15378,N_14521);
xnor U18749 (N_18749,N_14118,N_12645);
nor U18750 (N_18750,N_15801,N_18397);
or U18751 (N_18751,N_18527,N_16136);
nand U18752 (N_18752,N_16732,N_15991);
and U18753 (N_18753,N_17244,N_16260);
or U18754 (N_18754,N_15816,N_16350);
nor U18755 (N_18755,N_17833,N_17556);
and U18756 (N_18756,N_18689,N_16676);
or U18757 (N_18757,N_16356,N_15978);
and U18758 (N_18758,N_18291,N_17343);
or U18759 (N_18759,N_18308,N_18332);
and U18760 (N_18760,N_16480,N_16253);
and U18761 (N_18761,N_16493,N_18029);
or U18762 (N_18762,N_16247,N_16347);
or U18763 (N_18763,N_15990,N_15777);
nand U18764 (N_18764,N_16794,N_16543);
or U18765 (N_18765,N_17783,N_16994);
and U18766 (N_18766,N_16161,N_17298);
and U18767 (N_18767,N_18560,N_18662);
and U18768 (N_18768,N_17908,N_18730);
and U18769 (N_18769,N_18558,N_18409);
nor U18770 (N_18770,N_15955,N_18107);
or U18771 (N_18771,N_15819,N_16340);
nor U18772 (N_18772,N_17917,N_16127);
nor U18773 (N_18773,N_18654,N_18040);
and U18774 (N_18774,N_16502,N_15815);
or U18775 (N_18775,N_15793,N_17164);
nand U18776 (N_18776,N_18624,N_17455);
and U18777 (N_18777,N_17224,N_16036);
or U18778 (N_18778,N_16641,N_18283);
nor U18779 (N_18779,N_16984,N_16767);
and U18780 (N_18780,N_18278,N_17717);
or U18781 (N_18781,N_16847,N_18356);
nor U18782 (N_18782,N_16372,N_16640);
and U18783 (N_18783,N_15755,N_15694);
nand U18784 (N_18784,N_16388,N_17179);
or U18785 (N_18785,N_16571,N_16966);
and U18786 (N_18786,N_16780,N_18306);
or U18787 (N_18787,N_18389,N_16913);
and U18788 (N_18788,N_16105,N_17288);
nor U18789 (N_18789,N_16275,N_16169);
nor U18790 (N_18790,N_17046,N_17234);
nor U18791 (N_18791,N_18280,N_15664);
and U18792 (N_18792,N_16692,N_17883);
nor U18793 (N_18793,N_16745,N_17592);
or U18794 (N_18794,N_16657,N_18346);
nand U18795 (N_18795,N_15795,N_15626);
nor U18796 (N_18796,N_18217,N_18083);
and U18797 (N_18797,N_15829,N_17267);
nor U18798 (N_18798,N_16718,N_16018);
nor U18799 (N_18799,N_18252,N_17971);
or U18800 (N_18800,N_18676,N_18454);
nand U18801 (N_18801,N_16370,N_16039);
and U18802 (N_18802,N_15803,N_18208);
or U18803 (N_18803,N_17304,N_18489);
or U18804 (N_18804,N_18472,N_17416);
nand U18805 (N_18805,N_16735,N_15907);
and U18806 (N_18806,N_17182,N_16131);
nor U18807 (N_18807,N_18657,N_15920);
nand U18808 (N_18808,N_15870,N_15960);
nand U18809 (N_18809,N_17894,N_17061);
xnor U18810 (N_18810,N_15715,N_18355);
or U18811 (N_18811,N_16679,N_18392);
nand U18812 (N_18812,N_17710,N_18700);
and U18813 (N_18813,N_15969,N_18432);
nor U18814 (N_18814,N_15862,N_15672);
or U18815 (N_18815,N_17127,N_18644);
nor U18816 (N_18816,N_16695,N_17589);
nand U18817 (N_18817,N_16860,N_18089);
and U18818 (N_18818,N_16301,N_17738);
and U18819 (N_18819,N_16998,N_17200);
nand U18820 (N_18820,N_16896,N_16005);
xor U18821 (N_18821,N_16331,N_17148);
xnor U18822 (N_18822,N_18519,N_18012);
nand U18823 (N_18823,N_18388,N_18206);
xor U18824 (N_18824,N_17866,N_17897);
nor U18825 (N_18825,N_17207,N_15922);
nand U18826 (N_18826,N_16475,N_16077);
nor U18827 (N_18827,N_18600,N_16430);
or U18828 (N_18828,N_17106,N_18627);
nor U18829 (N_18829,N_16868,N_15917);
xnor U18830 (N_18830,N_17612,N_17209);
xnor U18831 (N_18831,N_15660,N_16599);
and U18832 (N_18832,N_18632,N_16007);
and U18833 (N_18833,N_15944,N_15948);
nand U18834 (N_18834,N_18646,N_17568);
or U18835 (N_18835,N_16550,N_15680);
nand U18836 (N_18836,N_16380,N_18652);
nor U18837 (N_18837,N_17566,N_16418);
xor U18838 (N_18838,N_17226,N_16021);
or U18839 (N_18839,N_18157,N_17362);
nor U18840 (N_18840,N_18643,N_15758);
nand U18841 (N_18841,N_15968,N_18670);
nor U18842 (N_18842,N_16216,N_15956);
xor U18843 (N_18843,N_17898,N_17645);
nand U18844 (N_18844,N_17052,N_17481);
or U18845 (N_18845,N_17837,N_17629);
nor U18846 (N_18846,N_17285,N_17730);
nand U18847 (N_18847,N_16920,N_18196);
and U18848 (N_18848,N_15796,N_15988);
or U18849 (N_18849,N_16225,N_18184);
nand U18850 (N_18850,N_15918,N_17047);
or U18851 (N_18851,N_18108,N_17684);
or U18852 (N_18852,N_16773,N_18547);
nand U18853 (N_18853,N_18729,N_17439);
nor U18854 (N_18854,N_17673,N_18578);
xnor U18855 (N_18855,N_17630,N_16511);
or U18856 (N_18856,N_18203,N_17407);
nand U18857 (N_18857,N_17790,N_17396);
or U18858 (N_18858,N_17133,N_15897);
or U18859 (N_18859,N_17900,N_16422);
nand U18860 (N_18860,N_17786,N_16804);
nor U18861 (N_18861,N_16013,N_17767);
or U18862 (N_18862,N_17654,N_15691);
and U18863 (N_18863,N_17518,N_17789);
nor U18864 (N_18864,N_17916,N_16704);
xor U18865 (N_18865,N_17063,N_17505);
nor U18866 (N_18866,N_17554,N_17014);
or U18867 (N_18867,N_16351,N_18200);
nand U18868 (N_18868,N_18188,N_17077);
and U18869 (N_18869,N_16555,N_18185);
nand U18870 (N_18870,N_16165,N_17136);
nand U18871 (N_18871,N_17907,N_16985);
and U18872 (N_18872,N_17252,N_16140);
nand U18873 (N_18873,N_16774,N_17644);
or U18874 (N_18874,N_17201,N_17433);
and U18875 (N_18875,N_18082,N_18164);
and U18876 (N_18876,N_15976,N_16623);
nor U18877 (N_18877,N_15647,N_18622);
xnor U18878 (N_18878,N_18704,N_17575);
nor U18879 (N_18879,N_16393,N_17797);
nand U18880 (N_18880,N_15943,N_17854);
or U18881 (N_18881,N_16783,N_16895);
nor U18882 (N_18882,N_18158,N_16006);
or U18883 (N_18883,N_16273,N_16038);
nor U18884 (N_18884,N_18360,N_16682);
or U18885 (N_18885,N_18366,N_15813);
xnor U18886 (N_18886,N_16609,N_16265);
nand U18887 (N_18887,N_17429,N_16980);
or U18888 (N_18888,N_15797,N_17109);
nand U18889 (N_18889,N_17468,N_17228);
nor U18890 (N_18890,N_16700,N_17183);
or U18891 (N_18891,N_18303,N_16378);
or U18892 (N_18892,N_17636,N_18336);
or U18893 (N_18893,N_15636,N_17778);
or U18894 (N_18894,N_18502,N_15656);
nor U18895 (N_18895,N_15696,N_16115);
or U18896 (N_18896,N_17162,N_18087);
nand U18897 (N_18897,N_17029,N_17752);
xor U18898 (N_18898,N_18016,N_16056);
or U18899 (N_18899,N_18733,N_16806);
and U18900 (N_18900,N_18343,N_16670);
and U18901 (N_18901,N_18615,N_18468);
nor U18902 (N_18902,N_16413,N_15727);
and U18903 (N_18903,N_16689,N_16172);
or U18904 (N_18904,N_18182,N_17159);
and U18905 (N_18905,N_17442,N_18162);
nor U18906 (N_18906,N_15788,N_16330);
and U18907 (N_18907,N_16143,N_18289);
nand U18908 (N_18908,N_16782,N_17422);
xor U18909 (N_18909,N_17300,N_18019);
xnor U18910 (N_18910,N_15842,N_17718);
or U18911 (N_18911,N_16314,N_17983);
or U18912 (N_18912,N_17969,N_18441);
or U18913 (N_18913,N_17191,N_17149);
nand U18914 (N_18914,N_18543,N_15650);
or U18915 (N_18915,N_16989,N_17291);
nand U18916 (N_18916,N_18529,N_17599);
or U18917 (N_18917,N_18501,N_17555);
nor U18918 (N_18918,N_18312,N_16122);
nor U18919 (N_18919,N_17432,N_18344);
nand U18920 (N_18920,N_18491,N_17461);
nand U18921 (N_18921,N_18500,N_15663);
nor U18922 (N_18922,N_17508,N_16589);
nand U18923 (N_18923,N_17277,N_16902);
and U18924 (N_18924,N_16433,N_17841);
or U18925 (N_18925,N_17990,N_17930);
nor U18926 (N_18926,N_16317,N_16646);
xor U18927 (N_18927,N_16389,N_16425);
or U18928 (N_18928,N_16394,N_17744);
nor U18929 (N_18929,N_16524,N_18744);
and U18930 (N_18930,N_16662,N_18212);
or U18931 (N_18931,N_17150,N_15642);
or U18932 (N_18932,N_18126,N_16906);
nor U18933 (N_18933,N_17375,N_16119);
and U18934 (N_18934,N_17009,N_18318);
and U18935 (N_18935,N_16274,N_17751);
or U18936 (N_18936,N_15753,N_16043);
or U18937 (N_18937,N_16016,N_18590);
and U18938 (N_18938,N_16835,N_17156);
and U18939 (N_18939,N_18380,N_17725);
nand U18940 (N_18940,N_17850,N_16278);
and U18941 (N_18941,N_16305,N_18116);
nand U18942 (N_18942,N_16476,N_17492);
and U18943 (N_18943,N_17064,N_18523);
nor U18944 (N_18944,N_15890,N_16941);
or U18945 (N_18945,N_16708,N_17862);
and U18946 (N_18946,N_15834,N_17175);
or U18947 (N_18947,N_15812,N_16492);
nor U18948 (N_18948,N_16009,N_18599);
xor U18949 (N_18949,N_16605,N_17070);
and U18950 (N_18950,N_18740,N_16456);
nor U18951 (N_18951,N_16232,N_16821);
and U18952 (N_18952,N_17485,N_16748);
nor U18953 (N_18953,N_16979,N_15703);
nand U18954 (N_18954,N_17440,N_16282);
and U18955 (N_18955,N_17827,N_16503);
and U18956 (N_18956,N_15669,N_15774);
nand U18957 (N_18957,N_16793,N_17737);
nor U18958 (N_18958,N_16033,N_17932);
xnor U18959 (N_18959,N_18002,N_17548);
or U18960 (N_18960,N_15790,N_16159);
nand U18961 (N_18961,N_15854,N_16720);
nor U18962 (N_18962,N_18139,N_16084);
nor U18963 (N_18963,N_16310,N_17292);
or U18964 (N_18964,N_17859,N_18288);
xnor U18965 (N_18965,N_17391,N_18651);
or U18966 (N_18966,N_15810,N_17262);
and U18967 (N_18967,N_16987,N_16927);
and U18968 (N_18968,N_17863,N_15958);
nand U18969 (N_18969,N_18546,N_18445);
or U18970 (N_18970,N_18358,N_16044);
nand U18971 (N_18971,N_17193,N_16027);
xor U18972 (N_18972,N_18013,N_15912);
nor U18973 (N_18973,N_16992,N_17855);
nand U18974 (N_18974,N_16360,N_17625);
and U18975 (N_18975,N_18717,N_15935);
or U18976 (N_18976,N_18100,N_16103);
nor U18977 (N_18977,N_17160,N_16839);
or U18978 (N_18978,N_17122,N_16775);
and U18979 (N_18979,N_17569,N_18426);
and U18980 (N_18980,N_16706,N_18414);
nand U18981 (N_18981,N_16227,N_15643);
nor U18982 (N_18982,N_16272,N_17289);
or U18983 (N_18983,N_18178,N_17781);
nand U18984 (N_18984,N_16327,N_15895);
and U18985 (N_18985,N_17516,N_17804);
or U18986 (N_18986,N_17558,N_16059);
nand U18987 (N_18987,N_16466,N_16861);
or U18988 (N_18988,N_15817,N_17980);
xnor U18989 (N_18989,N_18368,N_16956);
nand U18990 (N_18990,N_16454,N_16754);
and U18991 (N_18991,N_17506,N_18605);
nor U18992 (N_18992,N_18272,N_18297);
or U18993 (N_18993,N_17669,N_16784);
and U18994 (N_18994,N_15791,N_18150);
or U18995 (N_18995,N_18253,N_15893);
nand U18996 (N_18996,N_17801,N_17089);
or U18997 (N_18997,N_17638,N_17006);
nand U18998 (N_18998,N_15767,N_15689);
nand U18999 (N_18999,N_18498,N_17810);
xor U19000 (N_19000,N_16976,N_18007);
or U19001 (N_19001,N_17927,N_18731);
nor U19002 (N_19002,N_17984,N_16455);
nand U19003 (N_19003,N_17570,N_17614);
nor U19004 (N_19004,N_15732,N_18467);
and U19005 (N_19005,N_17830,N_18540);
or U19006 (N_19006,N_18068,N_18124);
or U19007 (N_19007,N_17661,N_18691);
nand U19008 (N_19008,N_16572,N_15786);
nor U19009 (N_19009,N_17755,N_17536);
and U19010 (N_19010,N_17126,N_15639);
nor U19011 (N_19011,N_17015,N_16551);
and U19012 (N_19012,N_17580,N_16924);
and U19013 (N_19013,N_16545,N_16121);
or U19014 (N_19014,N_18470,N_17988);
nor U19015 (N_19015,N_17271,N_16970);
nor U19016 (N_19016,N_17479,N_17004);
nor U19017 (N_19017,N_17372,N_18128);
and U19018 (N_19018,N_17078,N_15700);
or U19019 (N_19019,N_17315,N_16133);
or U19020 (N_19020,N_18394,N_18403);
or U19021 (N_19021,N_17694,N_18405);
xor U19022 (N_19022,N_16928,N_18055);
nand U19023 (N_19023,N_15825,N_17087);
nand U19024 (N_19024,N_16683,N_17013);
and U19025 (N_19025,N_15923,N_17377);
nand U19026 (N_19026,N_18106,N_17976);
nor U19027 (N_19027,N_16448,N_18473);
and U19028 (N_19028,N_18170,N_15994);
nand U19029 (N_19029,N_18058,N_16423);
or U19030 (N_19030,N_17931,N_16760);
or U19031 (N_19031,N_18550,N_15637);
xnor U19032 (N_19032,N_15823,N_16332);
nand U19033 (N_19033,N_16737,N_15720);
and U19034 (N_19034,N_17828,N_17739);
and U19035 (N_19035,N_16311,N_18216);
and U19036 (N_19036,N_17419,N_16712);
or U19037 (N_19037,N_17543,N_17050);
or U19038 (N_19038,N_17982,N_17280);
and U19039 (N_19039,N_16429,N_17912);
or U19040 (N_19040,N_15878,N_17911);
nand U19041 (N_19041,N_16324,N_16678);
xor U19042 (N_19042,N_16055,N_17116);
or U19043 (N_19043,N_17987,N_18149);
nor U19044 (N_19044,N_18061,N_16579);
and U19045 (N_19045,N_16320,N_17393);
xnor U19046 (N_19046,N_18461,N_18037);
and U19047 (N_19047,N_16163,N_16986);
or U19048 (N_19048,N_18134,N_18373);
or U19049 (N_19049,N_18193,N_16167);
or U19050 (N_19050,N_16101,N_17758);
nor U19051 (N_19051,N_17105,N_17026);
or U19052 (N_19052,N_17297,N_18351);
and U19053 (N_19053,N_17457,N_18245);
or U19054 (N_19054,N_17660,N_16444);
xnor U19055 (N_19055,N_18545,N_16786);
nand U19056 (N_19056,N_17920,N_18034);
xnor U19057 (N_19057,N_17222,N_16065);
nand U19058 (N_19058,N_16063,N_17495);
nand U19059 (N_19059,N_16208,N_15950);
or U19060 (N_19060,N_16538,N_18179);
nor U19061 (N_19061,N_17270,N_17596);
and U19062 (N_19062,N_15759,N_18505);
or U19063 (N_19063,N_17579,N_15760);
nand U19064 (N_19064,N_18737,N_18726);
nand U19065 (N_19065,N_18260,N_17065);
nor U19066 (N_19066,N_18009,N_16075);
nand U19067 (N_19067,N_18001,N_18528);
nand U19068 (N_19068,N_15709,N_18257);
nor U19069 (N_19069,N_16309,N_17449);
or U19070 (N_19070,N_16032,N_18555);
nor U19071 (N_19071,N_16564,N_17074);
nand U19072 (N_19072,N_18091,N_15780);
nor U19073 (N_19073,N_17102,N_17824);
nand U19074 (N_19074,N_18607,N_16749);
and U19075 (N_19075,N_16126,N_17761);
nand U19076 (N_19076,N_18071,N_17296);
or U19077 (N_19077,N_17799,N_16303);
or U19078 (N_19078,N_17978,N_18160);
nor U19079 (N_19079,N_15871,N_18130);
nand U19080 (N_19080,N_16681,N_18228);
xnor U19081 (N_19081,N_17793,N_17177);
nor U19082 (N_19082,N_17329,N_18577);
nor U19083 (N_19083,N_15783,N_16030);
nor U19084 (N_19084,N_15688,N_18492);
nor U19085 (N_19085,N_18172,N_16128);
nor U19086 (N_19086,N_16934,N_18112);
nor U19087 (N_19087,N_17544,N_16299);
xor U19088 (N_19088,N_16222,N_15926);
nand U19089 (N_19089,N_16441,N_18322);
and U19090 (N_19090,N_15718,N_17534);
nand U19091 (N_19091,N_16323,N_16669);
or U19092 (N_19092,N_16613,N_17302);
and U19093 (N_19093,N_16691,N_18140);
or U19094 (N_19094,N_18006,N_17060);
nor U19095 (N_19095,N_18113,N_16498);
nand U19096 (N_19096,N_16880,N_16250);
and U19097 (N_19097,N_18264,N_17722);
or U19098 (N_19098,N_16527,N_17626);
and U19099 (N_19099,N_17748,N_17650);
and U19100 (N_19100,N_16020,N_16089);
nand U19101 (N_19101,N_17732,N_16846);
or U19102 (N_19102,N_18439,N_16965);
and U19103 (N_19103,N_17999,N_18544);
xor U19104 (N_19104,N_16416,N_16522);
or U19105 (N_19105,N_18239,N_15966);
and U19106 (N_19106,N_16473,N_15652);
nor U19107 (N_19107,N_16379,N_18168);
or U19108 (N_19108,N_18635,N_18574);
or U19109 (N_19109,N_16743,N_17158);
nor U19110 (N_19110,N_16533,N_16409);
and U19111 (N_19111,N_16191,N_17510);
or U19112 (N_19112,N_17216,N_17206);
nor U19113 (N_19113,N_17048,N_17099);
nor U19114 (N_19114,N_15739,N_16668);
and U19115 (N_19115,N_15699,N_18310);
and U19116 (N_19116,N_17820,N_17400);
nand U19117 (N_19117,N_16183,N_16787);
and U19118 (N_19118,N_18067,N_16877);
nand U19119 (N_19119,N_18186,N_15939);
nand U19120 (N_19120,N_18442,N_17033);
or U19121 (N_19121,N_16485,N_18003);
nand U19122 (N_19122,N_18420,N_16346);
nand U19123 (N_19123,N_16544,N_17507);
nand U19124 (N_19124,N_16277,N_16813);
nor U19125 (N_19125,N_16325,N_15846);
nor U19126 (N_19126,N_15690,N_17968);
or U19127 (N_19127,N_17782,N_15904);
nor U19128 (N_19128,N_16694,N_18436);
nor U19129 (N_19129,N_15722,N_17151);
nor U19130 (N_19130,N_18549,N_17652);
xnor U19131 (N_19131,N_16242,N_16873);
and U19132 (N_19132,N_15936,N_16603);
and U19133 (N_19133,N_18135,N_18035);
nand U19134 (N_19134,N_18559,N_18483);
or U19135 (N_19135,N_17356,N_16808);
nor U19136 (N_19136,N_17809,N_17111);
nand U19137 (N_19137,N_16050,N_16680);
or U19138 (N_19138,N_17945,N_16628);
nand U19139 (N_19139,N_16845,N_15762);
nor U19140 (N_19140,N_16546,N_16481);
or U19141 (N_19141,N_16888,N_16625);
nor U19142 (N_19142,N_16539,N_17753);
nor U19143 (N_19143,N_17124,N_16637);
nand U19144 (N_19144,N_17016,N_17993);
nand U19145 (N_19145,N_16197,N_16396);
nor U19146 (N_19146,N_15877,N_18099);
or U19147 (N_19147,N_18030,N_16257);
nor U19148 (N_19148,N_15771,N_16442);
xor U19149 (N_19149,N_15998,N_16112);
nor U19150 (N_19150,N_17358,N_18133);
nand U19151 (N_19151,N_17918,N_16893);
nand U19152 (N_19152,N_17573,N_18463);
or U19153 (N_19153,N_17094,N_17379);
or U19154 (N_19154,N_16884,N_16534);
and U19155 (N_19155,N_17635,N_17688);
nand U19156 (N_19156,N_17607,N_16496);
nand U19157 (N_19157,N_16698,N_15894);
xnor U19158 (N_19158,N_17549,N_16184);
or U19159 (N_19159,N_17032,N_17192);
and U19160 (N_19160,N_16096,N_18621);
nor U19161 (N_19161,N_17038,N_18746);
xor U19162 (N_19162,N_18215,N_16536);
or U19163 (N_19163,N_17167,N_17414);
and U19164 (N_19164,N_18518,N_17235);
xnor U19165 (N_19165,N_17276,N_18383);
and U19166 (N_19166,N_17853,N_18451);
nor U19167 (N_19167,N_15919,N_18331);
nor U19168 (N_19168,N_17890,N_18334);
nor U19169 (N_19169,N_17211,N_17282);
or U19170 (N_19170,N_16865,N_16709);
nand U19171 (N_19171,N_18396,N_18353);
xor U19172 (N_19172,N_17500,N_16171);
nand U19173 (N_19173,N_16414,N_17974);
nor U19174 (N_19174,N_17446,N_18235);
nand U19175 (N_19175,N_17483,N_17772);
and U19176 (N_19176,N_18276,N_18121);
and U19177 (N_19177,N_16887,N_16925);
nand U19178 (N_19178,N_16114,N_17585);
or U19179 (N_19179,N_17521,N_18153);
and U19180 (N_19180,N_18000,N_17874);
and U19181 (N_19181,N_16553,N_17686);
or U19182 (N_19182,N_18204,N_16029);
and U19183 (N_19183,N_16195,N_16824);
nor U19184 (N_19184,N_16023,N_17985);
or U19185 (N_19185,N_16621,N_15781);
xor U19186 (N_19186,N_16959,N_16513);
and U19187 (N_19187,N_18370,N_16750);
and U19188 (N_19188,N_16015,N_17602);
and U19189 (N_19189,N_16329,N_17320);
nor U19190 (N_19190,N_17313,N_16932);
nor U19191 (N_19191,N_16437,N_16399);
nor U19192 (N_19192,N_16104,N_16339);
nand U19193 (N_19193,N_16490,N_18084);
nand U19194 (N_19194,N_16082,N_16362);
or U19195 (N_19195,N_17950,N_17595);
nand U19196 (N_19196,N_17463,N_16853);
or U19197 (N_19197,N_17450,N_18189);
nor U19198 (N_19198,N_17250,N_17478);
or U19199 (N_19199,N_18659,N_15980);
nand U19200 (N_19200,N_18633,N_15723);
and U19201 (N_19201,N_16557,N_18649);
or U19202 (N_19202,N_17165,N_16537);
nor U19203 (N_19203,N_17876,N_18410);
nor U19204 (N_19204,N_16060,N_16499);
or U19205 (N_19205,N_18720,N_15951);
nand U19206 (N_19206,N_16058,N_18117);
nand U19207 (N_19207,N_16828,N_16415);
nor U19208 (N_19208,N_16457,N_17293);
and U19209 (N_19209,N_16560,N_17491);
or U19210 (N_19210,N_17232,N_16120);
and U19211 (N_19211,N_15891,N_18125);
nand U19212 (N_19212,N_18137,N_17401);
nor U19213 (N_19213,N_16649,N_18259);
nor U19214 (N_19214,N_16831,N_17245);
or U19215 (N_19215,N_17129,N_15633);
nand U19216 (N_19216,N_18361,N_15908);
xnor U19217 (N_19217,N_17203,N_18275);
and U19218 (N_19218,N_18478,N_15670);
nor U19219 (N_19219,N_16703,N_16482);
nand U19220 (N_19220,N_16449,N_15845);
nor U19221 (N_19221,N_16952,N_17000);
nor U19222 (N_19222,N_16149,N_16259);
and U19223 (N_19223,N_15804,N_18508);
nor U19224 (N_19224,N_17085,N_17873);
or U19225 (N_19225,N_16578,N_18490);
xor U19226 (N_19226,N_17535,N_15822);
nand U19227 (N_19227,N_15757,N_18269);
nand U19228 (N_19228,N_17870,N_18497);
or U19229 (N_19229,N_17954,N_18151);
nand U19230 (N_19230,N_17538,N_17281);
nor U19231 (N_19231,N_15931,N_17671);
nand U19232 (N_19232,N_16474,N_18411);
nor U19233 (N_19233,N_18430,N_15776);
and U19234 (N_19234,N_16252,N_17480);
nor U19235 (N_19235,N_16478,N_18444);
xnor U19236 (N_19236,N_17194,N_17079);
nand U19237 (N_19237,N_16316,N_16001);
nand U19238 (N_19238,N_18052,N_16645);
nand U19239 (N_19239,N_18734,N_17672);
nand U19240 (N_19240,N_16427,N_18715);
nor U19241 (N_19241,N_18266,N_17656);
nor U19242 (N_19242,N_18412,N_16752);
and U19243 (N_19243,N_18023,N_16931);
or U19244 (N_19244,N_16978,N_16954);
nand U19245 (N_19245,N_18422,N_17657);
and U19246 (N_19246,N_16234,N_16917);
nor U19247 (N_19247,N_15867,N_17044);
nor U19248 (N_19248,N_18705,N_18364);
nor U19249 (N_19249,N_18415,N_16147);
and U19250 (N_19250,N_18379,N_17438);
nand U19251 (N_19251,N_16188,N_16298);
or U19252 (N_19252,N_16002,N_18515);
or U19253 (N_19253,N_16520,N_17947);
xor U19254 (N_19254,N_17040,N_15628);
nand U19255 (N_19255,N_15889,N_15833);
and U19256 (N_19256,N_16451,N_17887);
or U19257 (N_19257,N_17019,N_17511);
xnor U19258 (N_19258,N_16465,N_15925);
nand U19259 (N_19259,N_17023,N_17328);
and U19260 (N_19260,N_17723,N_17616);
nand U19261 (N_19261,N_15800,N_17076);
and U19262 (N_19262,N_16666,N_17229);
nand U19263 (N_19263,N_17817,N_17517);
nand U19264 (N_19264,N_17942,N_16019);
and U19265 (N_19265,N_16715,N_18036);
nand U19266 (N_19266,N_17195,N_18057);
nand U19267 (N_19267,N_16686,N_16531);
nand U19268 (N_19268,N_17152,N_15913);
nor U19269 (N_19269,N_16285,N_17103);
nor U19270 (N_19270,N_16193,N_17880);
nor U19271 (N_19271,N_16181,N_16081);
nor U19272 (N_19272,N_17365,N_18026);
and U19273 (N_19273,N_15632,N_16495);
nor U19274 (N_19274,N_18299,N_16607);
and U19275 (N_19275,N_16943,N_17591);
nand U19276 (N_19276,N_16069,N_15701);
and U19277 (N_19277,N_18668,N_16461);
nand U19278 (N_19278,N_18390,N_17803);
nand U19279 (N_19279,N_16816,N_16716);
xnor U19280 (N_19280,N_17404,N_17798);
nor U19281 (N_19281,N_18198,N_16610);
nor U19282 (N_19282,N_18301,N_15738);
or U19283 (N_19283,N_18262,N_16921);
or U19284 (N_19284,N_16955,N_16289);
nand U19285 (N_19285,N_16667,N_16615);
nor U19286 (N_19286,N_18080,N_17423);
and U19287 (N_19287,N_17905,N_17145);
or U19288 (N_19288,N_17588,N_15645);
and U19289 (N_19289,N_16757,N_18488);
nand U19290 (N_19290,N_15992,N_15928);
and U19291 (N_19291,N_17829,N_16135);
nor U19292 (N_19292,N_16664,N_16568);
and U19293 (N_19293,N_17719,N_17331);
and U19294 (N_19294,N_16699,N_18220);
nand U19295 (N_19295,N_18728,N_17254);
or U19296 (N_19296,N_18274,N_18074);
xor U19297 (N_19297,N_17665,N_17696);
or U19298 (N_19298,N_17769,N_17972);
or U19299 (N_19299,N_16850,N_17263);
or U19300 (N_19300,N_16900,N_16674);
or U19301 (N_19301,N_17878,N_18625);
and U19302 (N_19302,N_17119,N_15896);
xnor U19303 (N_19303,N_15770,N_15929);
or U19304 (N_19304,N_18180,N_15785);
xnor U19305 (N_19305,N_16636,N_18608);
and U19306 (N_19306,N_17088,N_18741);
and U19307 (N_19307,N_16858,N_17255);
nand U19308 (N_19308,N_17662,N_17199);
and U19309 (N_19309,N_16653,N_18154);
xnor U19310 (N_19310,N_16525,N_16690);
nor U19311 (N_19311,N_16395,N_15708);
nor U19312 (N_19312,N_16886,N_17699);
or U19313 (N_19313,N_17466,N_16085);
nor U19314 (N_19314,N_18105,N_17024);
nand U19315 (N_19315,N_17622,N_16072);
or U19316 (N_19316,N_17994,N_15856);
and U19317 (N_19317,N_16595,N_16049);
nor U19318 (N_19318,N_16701,N_18697);
nor U19319 (N_19319,N_17791,N_15989);
xor U19320 (N_19320,N_17274,N_16295);
and U19321 (N_19321,N_18342,N_18428);
nor U19322 (N_19322,N_16213,N_18022);
nor U19323 (N_19323,N_17332,N_16095);
nand U19324 (N_19324,N_16230,N_17646);
xor U19325 (N_19325,N_16685,N_16078);
or U19326 (N_19326,N_17754,N_17860);
and U19327 (N_19327,N_18506,N_17906);
or U19328 (N_19328,N_16602,N_16688);
and U19329 (N_19329,N_18330,N_17632);
nor U19330 (N_19330,N_18562,N_16926);
and U19331 (N_19331,N_17843,N_18465);
nor U19332 (N_19332,N_18187,N_16582);
and U19333 (N_19333,N_16064,N_15725);
nand U19334 (N_19334,N_15733,N_18333);
nand U19335 (N_19335,N_18177,N_17210);
or U19336 (N_19336,N_16785,N_16841);
nor U19337 (N_19337,N_16297,N_15784);
nand U19338 (N_19338,N_17173,N_16319);
or U19339 (N_19339,N_16663,N_17904);
and U19340 (N_19340,N_16180,N_18284);
and U19341 (N_19341,N_16964,N_16093);
xor U19342 (N_19342,N_15839,N_18571);
xnor U19343 (N_19343,N_16296,N_18494);
and U19344 (N_19344,N_17899,N_16874);
and U19345 (N_19345,N_18146,N_16730);
xor U19346 (N_19346,N_17387,N_17317);
nand U19347 (N_19347,N_17488,N_17852);
xor U19348 (N_19348,N_16106,N_16957);
nor U19349 (N_19349,N_16796,N_18377);
and U19350 (N_19350,N_16494,N_16182);
nand U19351 (N_19351,N_16432,N_17135);
or U19352 (N_19352,N_17198,N_15901);
nand U19353 (N_19353,N_16644,N_17885);
or U19354 (N_19354,N_17689,N_17034);
nor U19355 (N_19355,N_16530,N_15915);
nor U19356 (N_19356,N_17398,N_17337);
nor U19357 (N_19357,N_18119,N_16509);
nand U19358 (N_19358,N_17227,N_16953);
nor U19359 (N_19359,N_16929,N_18039);
nor U19360 (N_19360,N_16313,N_16629);
xor U19361 (N_19361,N_17677,N_16563);
or U19362 (N_19362,N_17773,N_16562);
or U19363 (N_19363,N_17690,N_18572);
or U19364 (N_19364,N_18211,N_17121);
and U19365 (N_19365,N_18290,N_15729);
and U19366 (N_19366,N_15736,N_16080);
nor U19367 (N_19367,N_17943,N_17886);
and U19368 (N_19368,N_18159,N_15716);
and U19369 (N_19369,N_18433,N_16141);
nand U19370 (N_19370,N_16202,N_17335);
nor U19371 (N_19371,N_18663,N_16764);
and U19372 (N_19372,N_16129,N_15887);
nand U19373 (N_19373,N_16622,N_18381);
or U19374 (N_19374,N_16012,N_16915);
or U19375 (N_19375,N_16408,N_17541);
nand U19376 (N_19376,N_17445,N_16830);
nor U19377 (N_19377,N_17641,N_16073);
or U19378 (N_19378,N_17264,N_17388);
and U19379 (N_19379,N_16446,N_18575);
nand U19380 (N_19380,N_16598,N_17540);
nor U19381 (N_19381,N_17451,N_18101);
or U19382 (N_19382,N_16385,N_18254);
nor U19383 (N_19383,N_18086,N_18045);
or U19384 (N_19384,N_18033,N_17370);
or U19385 (N_19385,N_17168,N_17218);
nand U19386 (N_19386,N_18693,N_15869);
nand U19387 (N_19387,N_18639,N_16744);
and U19388 (N_19388,N_18563,N_17326);
xor U19389 (N_19389,N_16286,N_17357);
nand U19390 (N_19390,N_15705,N_15860);
nand U19391 (N_19391,N_18321,N_18636);
and U19392 (N_19392,N_17134,N_16939);
nand U19393 (N_19393,N_18176,N_17838);
and U19394 (N_19394,N_17587,N_16271);
or U19395 (N_19395,N_17674,N_16588);
xnor U19396 (N_19396,N_17321,N_15909);
nand U19397 (N_19397,N_18238,N_17389);
and U19398 (N_19398,N_17698,N_18350);
nand U19399 (N_19399,N_18323,N_18046);
nand U19400 (N_19400,N_17745,N_17776);
nand U19401 (N_19401,N_17565,N_17237);
nand U19402 (N_19402,N_17241,N_16237);
nor U19403 (N_19403,N_16529,N_16693);
or U19404 (N_19404,N_16899,N_16421);
nand U19405 (N_19405,N_15836,N_16656);
nor U19406 (N_19406,N_16591,N_17604);
nand U19407 (N_19407,N_17430,N_18611);
xnor U19408 (N_19408,N_16584,N_17881);
and U19409 (N_19409,N_18399,N_16288);
nand U19410 (N_19410,N_17301,N_16583);
xnor U19411 (N_19411,N_16742,N_15649);
and U19412 (N_19412,N_17316,N_18213);
nor U19413 (N_19413,N_16769,N_15981);
or U19414 (N_19414,N_18191,N_17995);
and U19415 (N_19415,N_18156,N_18687);
or U19416 (N_19416,N_16223,N_17816);
nor U19417 (N_19417,N_17539,N_17001);
nand U19418 (N_19418,N_17651,N_17946);
xor U19419 (N_19419,N_16175,N_17794);
nand U19420 (N_19420,N_15996,N_16617);
and U19421 (N_19421,N_18684,N_15682);
nor U19422 (N_19422,N_18579,N_18295);
nand U19423 (N_19423,N_17261,N_17025);
or U19424 (N_19424,N_15764,N_16338);
nand U19425 (N_19425,N_17726,N_17266);
nor U19426 (N_19426,N_18169,N_16207);
nand U19427 (N_19427,N_15746,N_18521);
xor U19428 (N_19428,N_15974,N_16788);
and U19429 (N_19429,N_16771,N_17010);
xor U19430 (N_19430,N_16811,N_18049);
nand U19431 (N_19431,N_17057,N_15832);
nand U19432 (N_19432,N_15970,N_18329);
nor U19433 (N_19433,N_15644,N_18460);
xor U19434 (N_19434,N_16261,N_17923);
nand U19435 (N_19435,N_18300,N_17118);
nor U19436 (N_19436,N_16168,N_18354);
nand U19437 (N_19437,N_16062,N_17042);
nand U19438 (N_19438,N_17140,N_18338);
and U19439 (N_19439,N_18267,N_17713);
or U19440 (N_19440,N_18369,N_18664);
nand U19441 (N_19441,N_18735,N_16836);
nand U19442 (N_19442,N_18340,N_16238);
nand U19443 (N_19443,N_17992,N_17533);
nand U19444 (N_19444,N_15900,N_15811);
nand U19445 (N_19445,N_16377,N_18005);
or U19446 (N_19446,N_16046,N_17740);
and U19447 (N_19447,N_17681,N_16194);
nor U19448 (N_19448,N_17498,N_17352);
and U19449 (N_19449,N_17743,N_17800);
xor U19450 (N_19450,N_16540,N_18513);
nor U19451 (N_19451,N_15629,N_16614);
and U19452 (N_19452,N_17527,N_17066);
xor U19453 (N_19453,N_16558,N_16916);
and U19454 (N_19454,N_16728,N_17670);
and U19455 (N_19455,N_16235,N_16411);
nand U19456 (N_19456,N_16940,N_17002);
xnor U19457 (N_19457,N_16053,N_17269);
and U19458 (N_19458,N_17958,N_16326);
and U19459 (N_19459,N_18462,N_17497);
nand U19460 (N_19460,N_15993,N_16717);
and U19461 (N_19461,N_17344,N_16361);
nor U19462 (N_19462,N_17008,N_16108);
nand U19463 (N_19463,N_17640,N_15898);
or U19464 (N_19464,N_18526,N_17188);
nor U19465 (N_19465,N_15984,N_18613);
and U19466 (N_19466,N_15995,N_17312);
or U19467 (N_19467,N_16516,N_18250);
or U19468 (N_19468,N_16995,N_17489);
xor U19469 (N_19469,N_18580,N_17486);
or U19470 (N_19470,N_17997,N_16150);
nand U19471 (N_19471,N_17123,N_16731);
or U19472 (N_19472,N_17678,N_16923);
nor U19473 (N_19473,N_18293,N_18595);
or U19474 (N_19474,N_17272,N_16199);
xor U19475 (N_19475,N_16648,N_17021);
nor U19476 (N_19476,N_16371,N_17373);
nand U19477 (N_19477,N_17336,N_17957);
and U19478 (N_19478,N_17020,N_16497);
nor U19479 (N_19479,N_18714,N_17939);
nor U19480 (N_19480,N_17385,N_15959);
nand U19481 (N_19481,N_15674,N_17139);
and U19482 (N_19482,N_16462,N_17600);
nand U19483 (N_19483,N_16975,N_16170);
nand U19484 (N_19484,N_15971,N_17842);
or U19485 (N_19485,N_18419,N_15772);
nor U19486 (N_19486,N_15731,N_17225);
xor U19487 (N_19487,N_16797,N_18688);
and U19488 (N_19488,N_18395,N_15964);
and U19489 (N_19489,N_18309,N_16827);
or U19490 (N_19490,N_18711,N_17970);
and U19491 (N_19491,N_16130,N_16655);
and U19492 (N_19492,N_18471,N_16947);
nand U19493 (N_19493,N_18173,N_18171);
or U19494 (N_19494,N_16335,N_16762);
nor U19495 (N_19495,N_17406,N_17386);
and U19496 (N_19496,N_17427,N_17073);
xor U19497 (N_19497,N_16407,N_17875);
or U19498 (N_19498,N_15827,N_17458);
nor U19499 (N_19499,N_16526,N_17621);
or U19500 (N_19500,N_18516,N_16179);
or U19501 (N_19501,N_18362,N_18487);
nand U19502 (N_19502,N_15849,N_15735);
nor U19503 (N_19503,N_15792,N_15684);
nor U19504 (N_19504,N_16111,N_18024);
or U19505 (N_19505,N_16635,N_18721);
nor U19506 (N_19506,N_16922,N_15631);
nand U19507 (N_19507,N_15861,N_17253);
nor U19508 (N_19508,N_16647,N_18302);
and U19509 (N_19509,N_17882,N_18292);
nor U19510 (N_19510,N_17903,N_16254);
and U19511 (N_19511,N_17170,N_17308);
and U19512 (N_19512,N_18123,N_18551);
or U19513 (N_19513,N_18271,N_16721);
and U19514 (N_19514,N_18079,N_16025);
and U19515 (N_19515,N_18114,N_16283);
or U19516 (N_19516,N_18421,N_16240);
nor U19517 (N_19517,N_15765,N_16569);
nand U19518 (N_19518,N_16470,N_16146);
nand U19519 (N_19519,N_16435,N_16099);
xnor U19520 (N_19520,N_18534,N_18469);
nor U19521 (N_19521,N_17522,N_16400);
and U19522 (N_19522,N_16003,N_17779);
and U19523 (N_19523,N_18010,N_18685);
and U19524 (N_19524,N_16070,N_16334);
or U19525 (N_19525,N_17775,N_16777);
and U19526 (N_19526,N_17380,N_16083);
xnor U19527 (N_19527,N_17928,N_16097);
nor U19528 (N_19528,N_18387,N_16878);
xor U19529 (N_19529,N_17470,N_18566);
nor U19530 (N_19530,N_16945,N_17340);
nor U19531 (N_19531,N_17155,N_16486);
nand U19532 (N_19532,N_16512,N_15883);
nor U19533 (N_19533,N_18218,N_16107);
nand U19534 (N_19534,N_16566,N_17243);
and U19535 (N_19535,N_18210,N_15805);
and U19536 (N_19536,N_18616,N_17086);
nor U19537 (N_19537,N_18147,N_17703);
and U19538 (N_19538,N_15751,N_15686);
xor U19539 (N_19539,N_16439,N_17056);
xor U19540 (N_19540,N_15737,N_17394);
nand U19541 (N_19541,N_18576,N_18199);
xnor U19542 (N_19542,N_18738,N_16665);
nor U19543 (N_19543,N_17403,N_17821);
and U19544 (N_19544,N_17412,N_16341);
or U19545 (N_19545,N_17323,N_18594);
nand U19546 (N_19546,N_16192,N_15934);
or U19547 (N_19547,N_17892,N_18335);
or U19548 (N_19548,N_18384,N_16766);
nand U19549 (N_19549,N_18230,N_16577);
nand U19550 (N_19550,N_17615,N_18265);
nand U19551 (N_19551,N_16342,N_16304);
nor U19552 (N_19552,N_18708,N_18629);
xnor U19553 (N_19553,N_18614,N_15858);
and U19554 (N_19554,N_17196,N_15728);
or U19555 (N_19555,N_18407,N_16612);
nor U19556 (N_19556,N_15865,N_15627);
nor U19557 (N_19557,N_18104,N_17405);
nor U19558 (N_19558,N_16871,N_16727);
and U19559 (N_19559,N_16398,N_18709);
nor U19560 (N_19560,N_15668,N_16810);
or U19561 (N_19561,N_18314,N_17176);
or U19562 (N_19562,N_16832,N_16972);
xor U19563 (N_19563,N_16559,N_18201);
nor U19564 (N_19564,N_15831,N_18630);
nor U19565 (N_19565,N_17169,N_18286);
and U19566 (N_19566,N_16805,N_17153);
xnor U19567 (N_19567,N_17663,N_18060);
and U19568 (N_19568,N_16477,N_17948);
or U19569 (N_19569,N_17012,N_15673);
xnor U19570 (N_19570,N_16196,N_15714);
nor U19571 (N_19571,N_18435,N_16431);
nand U19572 (N_19572,N_18115,N_16849);
and U19573 (N_19573,N_18589,N_17934);
and U19574 (N_19574,N_16318,N_15659);
nor U19575 (N_19575,N_18591,N_16365);
nor U19576 (N_19576,N_17961,N_16958);
and U19577 (N_19577,N_18557,N_18347);
nand U19578 (N_19578,N_16198,N_15742);
or U19579 (N_19579,N_18618,N_17113);
nor U19580 (N_19580,N_16420,N_16903);
or U19581 (N_19581,N_18246,N_16842);
or U19582 (N_19582,N_17130,N_17597);
and U19583 (N_19583,N_18378,N_18048);
nand U19584 (N_19584,N_15662,N_16642);
nor U19585 (N_19585,N_17007,N_18449);
or U19586 (N_19586,N_15693,N_16825);
and U19587 (N_19587,N_16343,N_18486);
xor U19588 (N_19588,N_16086,N_16306);
or U19589 (N_19589,N_17720,N_15841);
nand U19590 (N_19590,N_18736,N_17760);
nand U19591 (N_19591,N_18581,N_16156);
or U19592 (N_19592,N_17542,N_18698);
nand U19593 (N_19593,N_16650,N_15654);
and U19594 (N_19594,N_16210,N_16624);
or U19595 (N_19595,N_18043,N_18088);
and U19596 (N_19596,N_17764,N_18584);
nand U19597 (N_19597,N_17840,N_18194);
xor U19598 (N_19598,N_16770,N_17826);
nand U19599 (N_19599,N_18694,N_17707);
nor U19600 (N_19600,N_15843,N_17062);
nand U19601 (N_19601,N_18477,N_16643);
xor U19602 (N_19602,N_18437,N_15749);
nand U19603 (N_19603,N_17256,N_16251);
nor U19604 (N_19604,N_17628,N_16778);
nor U19605 (N_19605,N_15651,N_16057);
nand U19606 (N_19606,N_18256,N_16035);
or U19607 (N_19607,N_16710,N_17962);
or U19608 (N_19608,N_18190,N_15724);
and U19609 (N_19609,N_15808,N_17949);
or U19610 (N_19610,N_16322,N_18122);
nand U19611 (N_19611,N_18586,N_16801);
or U19612 (N_19612,N_17759,N_15675);
and U19613 (N_19613,N_17836,N_16949);
nor U19614 (N_19614,N_18539,N_18163);
nand U19615 (N_19615,N_16908,N_16211);
nor U19616 (N_19616,N_16863,N_18226);
xor U19617 (N_19617,N_16593,N_17935);
or U19618 (N_19618,N_17197,N_17441);
or U19619 (N_19619,N_16630,N_18056);
nor U19620 (N_19620,N_17318,N_16228);
nor U19621 (N_19621,N_17879,N_17562);
or U19622 (N_19622,N_16654,N_16834);
and U19623 (N_19623,N_17574,N_16823);
and U19624 (N_19624,N_16523,N_18434);
nand U19625 (N_19625,N_18448,N_15916);
or U19626 (N_19626,N_17161,N_16162);
xor U19627 (N_19627,N_18077,N_18675);
or U19628 (N_19628,N_16279,N_17022);
nor U19629 (N_19629,N_18520,N_15905);
and U19630 (N_19630,N_17822,N_17955);
or U19631 (N_19631,N_17715,N_17531);
nor U19632 (N_19632,N_17731,N_16233);
or U19633 (N_19633,N_18041,N_15766);
xnor U19634 (N_19634,N_17334,N_17682);
nor U19635 (N_19635,N_17347,N_18221);
and U19636 (N_19636,N_17951,N_17584);
nor U19637 (N_19637,N_17576,N_18357);
and U19638 (N_19638,N_16218,N_17784);
or U19639 (N_19639,N_16548,N_17354);
or U19640 (N_19640,N_17763,N_18386);
or U19641 (N_19641,N_16017,N_15666);
nor U19642 (N_19642,N_16606,N_16510);
or U19643 (N_19643,N_18716,N_16392);
xor U19644 (N_19644,N_17659,N_17411);
or U19645 (N_19645,N_17091,N_16528);
or U19646 (N_19646,N_16294,N_17806);
and U19647 (N_19647,N_16776,N_16484);
and U19648 (N_19648,N_17236,N_18175);
nor U19649 (N_19649,N_16844,N_18376);
and U19650 (N_19650,N_16201,N_18452);
xor U19651 (N_19651,N_18669,N_16031);
or U19652 (N_19652,N_15863,N_17452);
or U19653 (N_19653,N_17913,N_16471);
and U19654 (N_19654,N_17647,N_16675);
nand U19655 (N_19655,N_17494,N_16918);
or U19656 (N_19656,N_18143,N_17353);
nor U19657 (N_19657,N_17501,N_17733);
xor U19658 (N_19658,N_17028,N_15704);
xor U19659 (N_19659,N_17037,N_17202);
nor U19660 (N_19660,N_17035,N_15837);
nor U19661 (N_19661,N_18313,N_16852);
nand U19662 (N_19662,N_18440,N_15809);
nand U19663 (N_19663,N_17747,N_18183);
nor U19664 (N_19664,N_16229,N_16542);
or U19665 (N_19665,N_18053,N_16405);
nor U19666 (N_19666,N_17303,N_15717);
or U19667 (N_19667,N_18423,N_17242);
xnor U19668 (N_19668,N_16248,N_15942);
and U19669 (N_19669,N_15824,N_17473);
or U19670 (N_19670,N_18243,N_18455);
and U19671 (N_19671,N_16417,N_18692);
or U19672 (N_19672,N_17884,N_15840);
nand U19673 (N_19673,N_16971,N_17552);
nor U19674 (N_19674,N_18044,N_16364);
nor U19675 (N_19675,N_17503,N_16501);
nand U19676 (N_19676,N_18014,N_17902);
or U19677 (N_19677,N_17110,N_16010);
and U19678 (N_19678,N_17490,N_17178);
or U19679 (N_19679,N_16672,N_18672);
xor U19680 (N_19680,N_17431,N_17163);
nand U19681 (N_19681,N_18723,N_18710);
nor U19682 (N_19682,N_17981,N_18667);
nand U19683 (N_19683,N_17397,N_17096);
nand U19684 (N_19684,N_16580,N_17695);
nor U19685 (N_19685,N_17807,N_16722);
nand U19686 (N_19686,N_16594,N_18311);
nand U19687 (N_19687,N_17676,N_16885);
or U19688 (N_19688,N_17278,N_17359);
or U19689 (N_19689,N_15671,N_16942);
nand U19690 (N_19690,N_18601,N_18385);
nand U19691 (N_19691,N_16946,N_17567);
nor U19692 (N_19692,N_16677,N_18628);
and U19693 (N_19693,N_17205,N_16822);
nor U19694 (N_19694,N_16109,N_15866);
or U19695 (N_19695,N_17059,N_16851);
or U19696 (N_19696,N_18038,N_18416);
nand U19697 (N_19697,N_18680,N_17701);
nor U19698 (N_19698,N_16231,N_18017);
nor U19699 (N_19699,N_18748,N_18219);
or U19700 (N_19700,N_17683,N_17217);
or U19701 (N_19701,N_17941,N_16993);
nand U19702 (N_19702,N_17132,N_17049);
and U19703 (N_19703,N_17290,N_17374);
or U19704 (N_19704,N_17410,N_18138);
nor U19705 (N_19705,N_16697,N_15821);
nand U19706 (N_19706,N_17487,N_15698);
or U19707 (N_19707,N_17618,N_17963);
or U19708 (N_19708,N_17039,N_16164);
or U19709 (N_19709,N_15752,N_16616);
nand U19710 (N_19710,N_15677,N_16791);
nand U19711 (N_19711,N_17526,N_17309);
or U19712 (N_19712,N_16707,N_15798);
and U19713 (N_19713,N_15910,N_16487);
xor U19714 (N_19714,N_16061,N_18382);
or U19715 (N_19715,N_16176,N_18724);
nand U19716 (N_19716,N_18320,N_17189);
and U19717 (N_19717,N_16585,N_16445);
xnor U19718 (N_19718,N_18047,N_18655);
and U19719 (N_19719,N_17901,N_15830);
and U19720 (N_19720,N_17257,N_16246);
nor U19721 (N_19721,N_17351,N_17611);
nor U19722 (N_19722,N_17157,N_17909);
nor U19723 (N_19723,N_18363,N_16576);
nand U19724 (N_19724,N_18681,N_16601);
and U19725 (N_19725,N_18610,N_16187);
nand U19726 (N_19726,N_16659,N_18078);
and U19727 (N_19727,N_16447,N_18294);
xnor U19728 (N_19728,N_16491,N_17742);
nor U19729 (N_19729,N_17219,N_17550);
nand U19730 (N_19730,N_16052,N_17617);
and U19731 (N_19731,N_17092,N_16500);
or U19732 (N_19732,N_15947,N_18051);
nor U19733 (N_19733,N_15794,N_16872);
and U19734 (N_19734,N_18427,N_17606);
nor U19735 (N_19735,N_16733,N_18236);
and U19736 (N_19736,N_18450,N_18141);
or U19737 (N_19737,N_18567,N_17691);
nand U19738 (N_19738,N_15685,N_18371);
nand U19739 (N_19739,N_18367,N_18233);
nor U19740 (N_19740,N_16792,N_16302);
nor U19741 (N_19741,N_17627,N_17117);
nand U19742 (N_19742,N_17054,N_17940);
nor U19743 (N_19743,N_17643,N_17114);
nor U19744 (N_19744,N_16443,N_18612);
nor U19745 (N_19745,N_16587,N_18085);
nor U19746 (N_19746,N_17240,N_18548);
or U19747 (N_19747,N_16219,N_18263);
and U19748 (N_19748,N_15940,N_16434);
and U19749 (N_19749,N_16719,N_17402);
and U19750 (N_19750,N_18227,N_17072);
nand U19751 (N_19751,N_16725,N_16258);
nor U19752 (N_19752,N_17915,N_18732);
nor U19753 (N_19753,N_16206,N_17345);
and U19754 (N_19754,N_16345,N_17273);
and U19755 (N_19755,N_15855,N_15986);
and U19756 (N_19756,N_16894,N_17213);
nand U19757 (N_19757,N_18592,N_16157);
or U19758 (N_19758,N_16397,N_16912);
nor U19759 (N_19759,N_17305,N_16597);
nand U19760 (N_19760,N_17142,N_16561);
xor U19761 (N_19761,N_15884,N_18102);
and U19762 (N_19762,N_18145,N_17083);
or U19763 (N_19763,N_15695,N_17766);
or U19764 (N_19764,N_15692,N_18642);
and U19765 (N_19765,N_17075,N_15938);
or U19766 (N_19766,N_17581,N_18277);
and U19767 (N_19767,N_18665,N_16384);
or U19768 (N_19768,N_16236,N_17067);
nor U19769 (N_19769,N_17469,N_15961);
or U19770 (N_19770,N_17299,N_17053);
nand U19771 (N_19771,N_15962,N_17768);
nor U19772 (N_19772,N_16881,N_16153);
nor U19773 (N_19773,N_16815,N_17551);
nor U19774 (N_19774,N_16308,N_18617);
and U19775 (N_19775,N_17910,N_18097);
nor U19776 (N_19776,N_16284,N_16212);
and U19777 (N_19777,N_15741,N_15814);
xor U19778 (N_19778,N_17482,N_17472);
xor U19779 (N_19779,N_16506,N_16795);
and U19780 (N_19780,N_17504,N_18447);
nor U19781 (N_19781,N_15743,N_17378);
or U19782 (N_19782,N_18096,N_18249);
nor U19783 (N_19783,N_17390,N_17180);
or U19784 (N_19784,N_15880,N_16367);
or U19785 (N_19785,N_16936,N_16739);
nand U19786 (N_19786,N_16068,N_16355);
nor U19787 (N_19787,N_15945,N_16173);
and U19788 (N_19788,N_17027,N_16011);
nor U19789 (N_19789,N_17823,N_17420);
nor U19790 (N_19790,N_17181,N_18021);
nor U19791 (N_19791,N_16469,N_18703);
or U19792 (N_19792,N_18431,N_16054);
nor U19793 (N_19793,N_18285,N_16517);
and U19794 (N_19794,N_18365,N_15853);
xnor U19795 (N_19795,N_16436,N_16209);
xnor U19796 (N_19796,N_16910,N_17399);
and U19797 (N_19797,N_17765,N_16293);
nand U19798 (N_19798,N_16424,N_17251);
or U19799 (N_19799,N_17186,N_17770);
or U19800 (N_19800,N_17642,N_18569);
nor U19801 (N_19801,N_17741,N_16901);
nor U19802 (N_19802,N_18679,N_15906);
or U19803 (N_19803,N_16937,N_17546);
or U19804 (N_19804,N_16554,N_16459);
and U19805 (N_19805,N_17230,N_18604);
nor U19806 (N_19806,N_17426,N_16280);
nand U19807 (N_19807,N_18328,N_18429);
xnor U19808 (N_19808,N_15657,N_18718);
nor U19809 (N_19809,N_17384,N_17421);
or U19810 (N_19810,N_16410,N_16268);
nor U19811 (N_19811,N_17265,N_17966);
nor U19812 (N_19812,N_16866,N_17553);
nor U19813 (N_19813,N_18564,N_18695);
or U19814 (N_19814,N_16359,N_17409);
nand U19815 (N_19815,N_17864,N_18231);
nand U19816 (N_19816,N_17808,N_15973);
nand U19817 (N_19817,N_17960,N_15665);
or U19818 (N_19818,N_16857,N_15987);
nand U19819 (N_19819,N_16983,N_17069);
or U19820 (N_19820,N_17214,N_16962);
and U19821 (N_19821,N_17728,N_16889);
or U19822 (N_19822,N_15702,N_15779);
or U19823 (N_19823,N_18337,N_17756);
and U19824 (N_19824,N_17664,N_17891);
and U19825 (N_19825,N_16067,N_18727);
nor U19826 (N_19826,N_17283,N_17346);
xor U19827 (N_19827,N_17705,N_16034);
xor U19828 (N_19828,N_15787,N_18638);
nor U19829 (N_19829,N_17620,N_17333);
nand U19830 (N_19830,N_15638,N_15879);
or U19831 (N_19831,N_18296,N_17476);
nand U19832 (N_19832,N_17938,N_17557);
or U19833 (N_19833,N_16837,N_16221);
nor U19834 (N_19834,N_17464,N_18503);
xor U19835 (N_19835,N_17249,N_17184);
nand U19836 (N_19836,N_17867,N_16740);
nor U19837 (N_19837,N_18683,N_16891);
nor U19838 (N_19838,N_17959,N_16814);
or U19839 (N_19839,N_17018,N_17146);
nand U19840 (N_19840,N_16729,N_16521);
and U19841 (N_19841,N_16948,N_18372);
nand U19842 (N_19842,N_16217,N_18537);
or U19843 (N_19843,N_16177,N_16552);
and U19844 (N_19844,N_17090,N_16726);
and U19845 (N_19845,N_17471,N_16137);
or U19846 (N_19846,N_17792,N_16768);
nor U19847 (N_19847,N_16604,N_16151);
nand U19848 (N_19848,N_18349,N_16753);
xnor U19849 (N_19849,N_17805,N_18678);
nand U19850 (N_19850,N_17736,N_15721);
and U19851 (N_19851,N_15941,N_18066);
nand U19852 (N_19852,N_16820,N_16967);
nand U19853 (N_19853,N_18725,N_15806);
or U19854 (N_19854,N_17563,N_17721);
nor U19855 (N_19855,N_18623,N_18582);
and U19856 (N_19856,N_17361,N_17093);
nand U19857 (N_19857,N_18524,N_17609);
xnor U19858 (N_19858,N_18650,N_15979);
or U19859 (N_19859,N_15761,N_18304);
or U19860 (N_19860,N_17322,N_15911);
xor U19861 (N_19861,N_17771,N_15953);
or U19862 (N_19862,N_18408,N_17583);
nand U19863 (N_19863,N_16440,N_18237);
and U19864 (N_19864,N_18512,N_16185);
nor U19865 (N_19865,N_16608,N_17525);
and U19866 (N_19866,N_16026,N_17847);
or U19867 (N_19867,N_17871,N_16403);
nand U19868 (N_19868,N_17687,N_17787);
nor U19869 (N_19869,N_18706,N_16464);
xor U19870 (N_19870,N_17750,N_16991);
nand U19871 (N_19871,N_18481,N_17260);
nor U19872 (N_19872,N_16174,N_17872);
nor U19873 (N_19873,N_16626,N_16658);
nor U19874 (N_19874,N_18531,N_17832);
or U19875 (N_19875,N_15886,N_16864);
nand U19876 (N_19876,N_17376,N_17865);
or U19877 (N_19877,N_15820,N_17603);
or U19878 (N_19878,N_18244,N_16736);
xor U19879 (N_19879,N_15683,N_15965);
nor U19880 (N_19880,N_15930,N_17314);
and U19881 (N_19881,N_16452,N_17577);
nor U19882 (N_19882,N_15937,N_16189);
or U19883 (N_19883,N_15921,N_17868);
nand U19884 (N_19884,N_17693,N_16292);
and U19885 (N_19885,N_17107,N_17137);
and U19886 (N_19886,N_17711,N_18004);
nor U19887 (N_19887,N_15678,N_15885);
nor U19888 (N_19888,N_17848,N_16241);
nand U19889 (N_19889,N_17895,N_17392);
and U19890 (N_19890,N_18696,N_16402);
nor U19891 (N_19891,N_16215,N_16826);
or U19892 (N_19892,N_17729,N_18641);
nor U19893 (N_19893,N_16139,N_17530);
nand U19894 (N_19894,N_16812,N_15711);
or U19895 (N_19895,N_15949,N_18701);
nor U19896 (N_19896,N_17633,N_16883);
and U19897 (N_19897,N_18316,N_16134);
nor U19898 (N_19898,N_16467,N_16673);
nand U19899 (N_19899,N_18095,N_15745);
nand U19900 (N_19900,N_16633,N_15726);
and U19901 (N_19901,N_18593,N_17857);
and U19902 (N_19902,N_16203,N_17929);
nand U19903 (N_19903,N_16907,N_16245);
and U19904 (N_19904,N_17979,N_15859);
and U19905 (N_19905,N_16800,N_17467);
nor U19906 (N_19906,N_17338,N_15676);
nor U19907 (N_19907,N_16968,N_17381);
and U19908 (N_19908,N_16307,N_18192);
nand U19909 (N_19909,N_16428,N_18682);
and U19910 (N_19910,N_17475,N_15634);
or U19911 (N_19911,N_17582,N_17749);
nor U19912 (N_19912,N_17417,N_17259);
nor U19913 (N_19913,N_16333,N_16573);
and U19914 (N_19914,N_16930,N_17408);
or U19915 (N_19915,N_15874,N_16586);
xor U19916 (N_19916,N_17519,N_17936);
and U19917 (N_19917,N_17474,N_18417);
nand U19918 (N_19918,N_18597,N_15740);
and U19919 (N_19919,N_18443,N_16898);
nand U19920 (N_19920,N_16066,N_17097);
or U19921 (N_19921,N_16746,N_15681);
nand U19922 (N_19922,N_18476,N_17712);
nor U19923 (N_19923,N_17051,N_18406);
or U19924 (N_19924,N_17914,N_16803);
or U19925 (N_19925,N_15851,N_15754);
and U19926 (N_19926,N_17965,N_17413);
nor U19927 (N_19927,N_17818,N_15707);
or U19928 (N_19928,N_15826,N_18425);
nor U19929 (N_19929,N_16876,N_17141);
nand U19930 (N_19930,N_17058,N_17655);
or U19931 (N_19931,N_15997,N_16269);
and U19932 (N_19932,N_16426,N_16859);
nor U19933 (N_19933,N_17564,N_17839);
nor U19934 (N_19934,N_16178,N_16024);
or U19935 (N_19935,N_16519,N_17952);
nand U19936 (N_19936,N_16840,N_17819);
nor U19937 (N_19937,N_18482,N_18094);
and U19938 (N_19938,N_16040,N_16091);
or U19939 (N_19939,N_18136,N_18375);
or U19940 (N_19940,N_17350,N_18127);
nor U19941 (N_19941,N_15625,N_17815);
or U19942 (N_19942,N_16387,N_18553);
and U19943 (N_19943,N_16590,N_17327);
or U19944 (N_19944,N_18656,N_18686);
or U19945 (N_19945,N_18446,N_15899);
nand U19946 (N_19946,N_17708,N_16369);
nand U19947 (N_19947,N_18050,N_18637);
nor U19948 (N_19948,N_16145,N_15655);
and U19949 (N_19949,N_18484,N_16450);
nand U19950 (N_19950,N_16856,N_16504);
nand U19951 (N_19951,N_16041,N_18307);
nor U19952 (N_19952,N_15873,N_18339);
or U19953 (N_19953,N_18287,N_16138);
or U19954 (N_19954,N_16981,N_17623);
or U19955 (N_19955,N_17115,N_16160);
or U19956 (N_19956,N_18359,N_18120);
nor U19957 (N_19957,N_16037,N_17082);
or U19958 (N_19958,N_16911,N_15954);
nand U19959 (N_19959,N_17003,N_18223);
nand U19960 (N_19960,N_16779,N_16074);
xor U19961 (N_19961,N_18073,N_17125);
or U19962 (N_19962,N_18587,N_16008);
and U19963 (N_19963,N_16244,N_18240);
nand U19964 (N_19964,N_17425,N_16000);
nor U19965 (N_19965,N_18674,N_16819);
nand U19966 (N_19966,N_18404,N_17284);
and U19967 (N_19967,N_18258,N_17998);
or U19968 (N_19968,N_18018,N_17279);
nand U19969 (N_19969,N_17762,N_18493);
nor U19970 (N_19970,N_17383,N_17925);
nand U19971 (N_19971,N_18166,N_16532);
nand U19972 (N_19972,N_16696,N_18197);
or U19973 (N_19973,N_17220,N_18424);
and U19974 (N_19974,N_17788,N_18401);
nor U19975 (N_19975,N_17637,N_15807);
xor U19976 (N_19976,N_17706,N_17045);
xor U19977 (N_19977,N_18319,N_16468);
and U19978 (N_19978,N_18391,N_15748);
nand U19979 (N_19979,N_16862,N_18713);
and U19980 (N_19980,N_17311,N_17973);
nor U19981 (N_19981,N_17700,N_17349);
and U19982 (N_19982,N_17590,N_18015);
and U19983 (N_19983,N_17537,N_17889);
and U19984 (N_19984,N_17921,N_18270);
nor U19985 (N_19985,N_16357,N_16652);
nand U19986 (N_19986,N_18722,N_18648);
or U19987 (N_19987,N_16092,N_17496);
nand U19988 (N_19988,N_17825,N_18129);
and U19989 (N_19989,N_16483,N_17716);
and U19990 (N_19990,N_16661,N_16974);
or U19991 (N_19991,N_18496,N_16950);
nand U19992 (N_19992,N_18561,N_18702);
nor U19993 (N_19993,N_18118,N_18699);
and U19994 (N_19994,N_18480,N_17679);
nor U19995 (N_19995,N_16102,N_17780);
xnor U19996 (N_19996,N_15914,N_18749);
and U19997 (N_19997,N_15927,N_18224);
and U19998 (N_19998,N_16963,N_18069);
or U19999 (N_19999,N_15775,N_16042);
nor U20000 (N_20000,N_16110,N_17084);
or U20001 (N_20001,N_17437,N_16118);
nand U20002 (N_20002,N_16123,N_18225);
nand U20003 (N_20003,N_18413,N_18743);
nand U20004 (N_20004,N_16807,N_16249);
nor U20005 (N_20005,N_16022,N_15844);
and U20006 (N_20006,N_17295,N_18485);
xor U20007 (N_20007,N_18542,N_18054);
nor U20008 (N_20008,N_18514,N_18081);
nor U20009 (N_20009,N_16882,N_16205);
or U20010 (N_20010,N_17248,N_17796);
xnor U20011 (N_20011,N_17360,N_17212);
xor U20012 (N_20012,N_16982,N_16734);
or U20013 (N_20013,N_17601,N_16344);
nor U20014 (N_20014,N_16144,N_18573);
nor U20015 (N_20015,N_17324,N_17247);
and U20016 (N_20016,N_15640,N_15882);
nor U20017 (N_20017,N_16567,N_16627);
or U20018 (N_20018,N_17275,N_17835);
or U20019 (N_20019,N_17680,N_17231);
nand U20020 (N_20020,N_16515,N_17144);
or U20021 (N_20021,N_16158,N_17944);
or U20022 (N_20022,N_16472,N_15933);
nand U20023 (N_20023,N_15687,N_17896);
nand U20024 (N_20024,N_16098,N_16671);
and U20025 (N_20025,N_18232,N_17477);
nor U20026 (N_20026,N_17991,N_16375);
or U20027 (N_20027,N_18144,N_15734);
nand U20028 (N_20028,N_16116,N_17095);
xnor U20029 (N_20029,N_15852,N_18251);
nand U20030 (N_20030,N_15653,N_17702);
and U20031 (N_20031,N_16904,N_18418);
nand U20032 (N_20032,N_17844,N_18626);
xnor U20033 (N_20033,N_17355,N_16489);
nor U20034 (N_20034,N_17735,N_16618);
nor U20035 (N_20035,N_16761,N_16723);
or U20036 (N_20036,N_16518,N_16631);
or U20037 (N_20037,N_16756,N_16781);
nand U20038 (N_20038,N_16488,N_16818);
or U20039 (N_20039,N_17204,N_17560);
nand U20040 (N_20040,N_15946,N_17869);
or U20041 (N_20041,N_15828,N_17509);
nor U20042 (N_20042,N_18398,N_17424);
and U20043 (N_20043,N_17112,N_17462);
and U20044 (N_20044,N_17774,N_17532);
xor U20045 (N_20045,N_17185,N_18281);
and U20046 (N_20046,N_16724,N_16028);
nor U20047 (N_20047,N_18161,N_15932);
nand U20048 (N_20048,N_18324,N_16366);
nand U20049 (N_20049,N_16048,N_18565);
or U20050 (N_20050,N_18032,N_18222);
nor U20051 (N_20051,N_16620,N_17734);
xor U20052 (N_20052,N_18317,N_15847);
nor U20053 (N_20053,N_18207,N_17147);
nor U20054 (N_20054,N_15744,N_16592);
nand U20055 (N_20055,N_18174,N_16220);
and U20056 (N_20056,N_16166,N_16373);
xor U20057 (N_20057,N_18165,N_15747);
xor U20058 (N_20058,N_16076,N_16684);
and U20059 (N_20059,N_16619,N_16090);
nand U20060 (N_20060,N_16353,N_16763);
nor U20061 (N_20061,N_16507,N_16152);
nor U20062 (N_20062,N_18598,N_16632);
and U20063 (N_20063,N_18202,N_18530);
nor U20064 (N_20064,N_17465,N_17996);
or U20065 (N_20065,N_16508,N_17238);
nand U20066 (N_20066,N_16186,N_17845);
nand U20067 (N_20067,N_17081,N_16276);
or U20068 (N_20068,N_18556,N_15648);
or U20069 (N_20069,N_18028,N_15872);
and U20070 (N_20070,N_17005,N_17594);
nand U20071 (N_20071,N_17528,N_18152);
nand U20072 (N_20072,N_17363,N_17724);
and U20073 (N_20073,N_17138,N_17529);
or U20074 (N_20074,N_17011,N_16154);
nor U20075 (N_20075,N_17524,N_16281);
nor U20076 (N_20076,N_17418,N_18241);
nand U20077 (N_20077,N_15848,N_17172);
or U20078 (N_20078,N_17619,N_18660);
nor U20079 (N_20079,N_17667,N_17515);
nor U20080 (N_20080,N_16639,N_17608);
or U20081 (N_20081,N_16611,N_18583);
nor U20082 (N_20082,N_16570,N_18402);
nand U20083 (N_20083,N_16363,N_16419);
or U20084 (N_20084,N_17348,N_16406);
nand U20085 (N_20085,N_15875,N_17325);
and U20086 (N_20086,N_15835,N_16869);
nor U20087 (N_20087,N_17435,N_18438);
nand U20088 (N_20088,N_18092,N_15972);
nand U20089 (N_20089,N_17858,N_18541);
and U20090 (N_20090,N_17460,N_17367);
nor U20091 (N_20091,N_17068,N_15838);
or U20092 (N_20092,N_16155,N_15881);
nand U20093 (N_20093,N_16321,N_18507);
and U20094 (N_20094,N_17443,N_17685);
or U20095 (N_20095,N_17310,N_18739);
or U20096 (N_20096,N_17187,N_18645);
nand U20097 (N_20097,N_16124,N_17513);
nand U20098 (N_20098,N_15975,N_18712);
xnor U20099 (N_20099,N_17922,N_17709);
and U20100 (N_20100,N_17610,N_17956);
nor U20101 (N_20101,N_17190,N_17834);
or U20102 (N_20102,N_16867,N_16575);
xnor U20103 (N_20103,N_16596,N_15868);
nor U20104 (N_20104,N_17937,N_17547);
nand U20105 (N_20105,N_15667,N_17666);
and U20106 (N_20106,N_18596,N_18315);
nor U20107 (N_20107,N_18690,N_16463);
nand U20108 (N_20108,N_16565,N_17108);
and U20109 (N_20109,N_17653,N_16574);
nand U20110 (N_20110,N_16809,N_16505);
nand U20111 (N_20111,N_18588,N_15818);
xor U20112 (N_20112,N_18103,N_15730);
xnor U20113 (N_20113,N_16765,N_18062);
and U20114 (N_20114,N_18042,N_15983);
nand U20115 (N_20115,N_15957,N_18305);
nand U20116 (N_20116,N_17131,N_16266);
or U20117 (N_20117,N_16535,N_15763);
and U20118 (N_20118,N_15661,N_15864);
and U20119 (N_20119,N_16312,N_18229);
or U20120 (N_20120,N_16190,N_17888);
nand U20121 (N_20121,N_16125,N_18142);
or U20122 (N_20122,N_18538,N_18341);
xor U20123 (N_20123,N_18509,N_16634);
and U20124 (N_20124,N_16713,N_17055);
nand U20125 (N_20125,N_17342,N_18025);
nand U20126 (N_20126,N_17924,N_17975);
or U20127 (N_20127,N_16264,N_17434);
and U20128 (N_20128,N_16239,N_17287);
and U20129 (N_20129,N_17030,N_18458);
nand U20130 (N_20130,N_16386,N_16789);
nor U20131 (N_20131,N_17456,N_16833);
nand U20132 (N_20132,N_18532,N_15635);
or U20133 (N_20133,N_17926,N_16438);
nand U20134 (N_20134,N_18745,N_16838);
and U20135 (N_20135,N_17294,N_17813);
nor U20136 (N_20136,N_17459,N_16638);
or U20137 (N_20137,N_18609,N_17561);
and U20138 (N_20138,N_16142,N_18647);
nand U20139 (N_20139,N_16255,N_18552);
or U20140 (N_20140,N_17846,N_16798);
and U20141 (N_20141,N_16349,N_16897);
or U20142 (N_20142,N_15789,N_15982);
nand U20143 (N_20143,N_18533,N_18234);
xor U20144 (N_20144,N_17395,N_17371);
nor U20145 (N_20145,N_16988,N_16711);
nor U20146 (N_20146,N_18619,N_16263);
nand U20147 (N_20147,N_18090,N_17697);
nand U20148 (N_20148,N_18719,N_18070);
or U20149 (N_20149,N_16997,N_17415);
and U20150 (N_20150,N_15756,N_16224);
nand U20151 (N_20151,N_16875,N_16758);
and U20152 (N_20152,N_15802,N_16996);
nor U20153 (N_20153,N_17593,N_16687);
nor U20154 (N_20154,N_15888,N_16990);
and U20155 (N_20155,N_18268,N_16226);
or U20156 (N_20156,N_17795,N_18075);
nor U20157 (N_20157,N_17523,N_17239);
or U20158 (N_20158,N_17366,N_17631);
nand U20159 (N_20159,N_17436,N_17977);
or U20160 (N_20160,N_16256,N_16004);
and U20161 (N_20161,N_16905,N_18457);
or U20162 (N_20162,N_16287,N_17080);
nand U20163 (N_20163,N_17814,N_18666);
or U20164 (N_20164,N_17964,N_16374);
xnor U20165 (N_20165,N_18466,N_17031);
or U20166 (N_20166,N_17877,N_17727);
nor U20167 (N_20167,N_17953,N_15903);
xor U20168 (N_20168,N_17499,N_16951);
nand U20169 (N_20169,N_17444,N_15630);
or U20170 (N_20170,N_18167,N_15719);
xnor U20171 (N_20171,N_17382,N_16772);
nand U20172 (N_20172,N_17520,N_18155);
or U20173 (N_20173,N_17246,N_16547);
nand U20174 (N_20174,N_18535,N_18658);
nand U20175 (N_20175,N_16817,N_16404);
nor U20176 (N_20176,N_16747,N_18065);
or U20177 (N_20177,N_17319,N_18109);
xnor U20178 (N_20178,N_16382,N_18568);
nand U20179 (N_20179,N_16336,N_17856);
and U20180 (N_20180,N_16977,N_16909);
xnor U20181 (N_20181,N_16660,N_15892);
xor U20182 (N_20182,N_16100,N_16879);
nand U20183 (N_20183,N_18453,N_16848);
nand U20184 (N_20184,N_17512,N_18209);
nand U20185 (N_20185,N_16148,N_17369);
and U20186 (N_20186,N_17493,N_18707);
xor U20187 (N_20187,N_18063,N_18027);
xnor U20188 (N_20188,N_15977,N_17634);
and U20189 (N_20189,N_18585,N_15902);
nor U20190 (N_20190,N_18374,N_15679);
nor U20191 (N_20191,N_16854,N_17649);
or U20192 (N_20192,N_18247,N_17605);
xor U20193 (N_20193,N_15769,N_18110);
nor U20194 (N_20194,N_16383,N_15999);
and U20195 (N_20195,N_16973,N_16458);
and U20196 (N_20196,N_17143,N_18459);
or U20197 (N_20197,N_17849,N_16391);
nand U20198 (N_20198,N_16802,N_16094);
or U20199 (N_20199,N_15768,N_17986);
nor U20200 (N_20200,N_17448,N_17648);
and U20201 (N_20201,N_16702,N_15924);
and U20202 (N_20202,N_18603,N_18570);
and U20203 (N_20203,N_17861,N_15850);
nand U20204 (N_20204,N_16381,N_17258);
and U20205 (N_20205,N_15799,N_16214);
and U20206 (N_20206,N_16390,N_16960);
and U20207 (N_20207,N_17098,N_18606);
xnor U20208 (N_20208,N_17215,N_17484);
or U20209 (N_20209,N_16368,N_17831);
nand U20210 (N_20210,N_16358,N_17208);
nand U20211 (N_20211,N_16051,N_16890);
and U20212 (N_20212,N_16045,N_16935);
and U20213 (N_20213,N_16714,N_16870);
or U20214 (N_20214,N_16079,N_16352);
or U20215 (N_20215,N_17668,N_17428);
nand U20216 (N_20216,N_16479,N_17851);
and U20217 (N_20217,N_18348,N_18011);
or U20218 (N_20218,N_18475,N_17613);
and U20219 (N_20219,N_16914,N_16376);
and U20220 (N_20220,N_16751,N_18456);
nand U20221 (N_20221,N_16014,N_18474);
or U20222 (N_20222,N_18131,N_17368);
nand U20223 (N_20223,N_16290,N_18181);
nor U20224 (N_20224,N_16705,N_16117);
xor U20225 (N_20225,N_17559,N_18072);
xnor U20226 (N_20226,N_18479,N_18205);
or U20227 (N_20227,N_17041,N_17893);
nand U20228 (N_20228,N_18111,N_16855);
nand U20229 (N_20229,N_18525,N_16738);
and U20230 (N_20230,N_18554,N_16354);
or U20231 (N_20231,N_17104,N_15697);
or U20232 (N_20232,N_16969,N_18634);
nor U20233 (N_20233,N_16071,N_15985);
xor U20234 (N_20234,N_17598,N_16132);
nand U20235 (N_20235,N_17502,N_17919);
nor U20236 (N_20236,N_18499,N_15713);
or U20237 (N_20237,N_17545,N_17128);
nand U20238 (N_20238,N_17306,N_17514);
or U20239 (N_20239,N_15963,N_15967);
xor U20240 (N_20240,N_18536,N_17802);
and U20241 (N_20241,N_18352,N_16262);
or U20242 (N_20242,N_18076,N_16541);
or U20243 (N_20243,N_17017,N_17624);
and U20244 (N_20244,N_18661,N_17286);
nand U20245 (N_20245,N_17154,N_17675);
and U20246 (N_20246,N_15712,N_16790);
nor U20247 (N_20247,N_17071,N_17120);
nand U20248 (N_20248,N_16651,N_18214);
or U20249 (N_20249,N_15773,N_18640);
nor U20250 (N_20250,N_18242,N_17233);
nor U20251 (N_20251,N_17221,N_16270);
xor U20252 (N_20252,N_18273,N_18248);
or U20253 (N_20253,N_17967,N_17777);
and U20254 (N_20254,N_18282,N_16549);
xor U20255 (N_20255,N_17453,N_17454);
and U20256 (N_20256,N_17989,N_16999);
nor U20257 (N_20257,N_17100,N_17704);
nor U20258 (N_20258,N_16961,N_17341);
and U20259 (N_20259,N_17036,N_18326);
nand U20260 (N_20260,N_16741,N_17692);
or U20261 (N_20261,N_18400,N_16300);
nor U20262 (N_20262,N_16113,N_17043);
nand U20263 (N_20263,N_18464,N_17811);
and U20264 (N_20264,N_17933,N_18298);
and U20265 (N_20265,N_18602,N_16938);
nor U20266 (N_20266,N_15782,N_18677);
and U20267 (N_20267,N_17268,N_15646);
xor U20268 (N_20268,N_18345,N_16401);
and U20269 (N_20269,N_15658,N_18517);
and U20270 (N_20270,N_16348,N_17223);
or U20271 (N_20271,N_17572,N_17714);
xnor U20272 (N_20272,N_16460,N_17586);
nand U20273 (N_20273,N_17658,N_16047);
xor U20274 (N_20274,N_15778,N_16581);
xnor U20275 (N_20275,N_18064,N_16892);
nand U20276 (N_20276,N_18511,N_16514);
nand U20277 (N_20277,N_18325,N_16829);
or U20278 (N_20278,N_17447,N_18327);
and U20279 (N_20279,N_17571,N_16337);
and U20280 (N_20280,N_15641,N_18059);
or U20281 (N_20281,N_15710,N_18098);
or U20282 (N_20282,N_15750,N_18504);
and U20283 (N_20283,N_16315,N_17578);
and U20284 (N_20284,N_18631,N_18255);
nand U20285 (N_20285,N_16328,N_17812);
and U20286 (N_20286,N_17757,N_17166);
and U20287 (N_20287,N_16944,N_18620);
and U20288 (N_20288,N_17101,N_15952);
nand U20289 (N_20289,N_16600,N_18008);
xor U20290 (N_20290,N_16843,N_15857);
or U20291 (N_20291,N_18195,N_18093);
nand U20292 (N_20292,N_18020,N_16755);
nand U20293 (N_20293,N_16412,N_16556);
nor U20294 (N_20294,N_18742,N_18261);
nand U20295 (N_20295,N_17330,N_18671);
nand U20296 (N_20296,N_16453,N_17171);
xnor U20297 (N_20297,N_16200,N_16919);
nor U20298 (N_20298,N_18747,N_16267);
and U20299 (N_20299,N_18653,N_17339);
or U20300 (N_20300,N_15706,N_18148);
or U20301 (N_20301,N_18279,N_16204);
nand U20302 (N_20302,N_16291,N_18522);
and U20303 (N_20303,N_17639,N_16933);
and U20304 (N_20304,N_17307,N_17364);
nor U20305 (N_20305,N_18132,N_16243);
xor U20306 (N_20306,N_18510,N_18031);
nand U20307 (N_20307,N_15876,N_17746);
and U20308 (N_20308,N_16799,N_17174);
or U20309 (N_20309,N_16759,N_18495);
or U20310 (N_20310,N_18673,N_16087);
or U20311 (N_20311,N_18393,N_16088);
or U20312 (N_20312,N_17785,N_18361);
or U20313 (N_20313,N_16749,N_18252);
xor U20314 (N_20314,N_17134,N_15685);
nor U20315 (N_20315,N_18654,N_16835);
or U20316 (N_20316,N_15848,N_17264);
nor U20317 (N_20317,N_17655,N_17882);
nor U20318 (N_20318,N_18024,N_17317);
and U20319 (N_20319,N_18138,N_16961);
and U20320 (N_20320,N_17825,N_17908);
nand U20321 (N_20321,N_17154,N_18379);
or U20322 (N_20322,N_16784,N_16759);
nand U20323 (N_20323,N_17376,N_16818);
or U20324 (N_20324,N_18490,N_16850);
and U20325 (N_20325,N_16850,N_17733);
or U20326 (N_20326,N_17874,N_15928);
nand U20327 (N_20327,N_18578,N_15763);
or U20328 (N_20328,N_18539,N_17379);
and U20329 (N_20329,N_17996,N_17426);
nor U20330 (N_20330,N_17662,N_17457);
and U20331 (N_20331,N_15701,N_17390);
xnor U20332 (N_20332,N_16315,N_18316);
nor U20333 (N_20333,N_16784,N_17435);
and U20334 (N_20334,N_17253,N_17459);
xnor U20335 (N_20335,N_15835,N_17044);
or U20336 (N_20336,N_17029,N_16401);
nand U20337 (N_20337,N_17972,N_17037);
and U20338 (N_20338,N_18370,N_16976);
or U20339 (N_20339,N_16202,N_15690);
nor U20340 (N_20340,N_15865,N_18402);
nor U20341 (N_20341,N_15923,N_16363);
nand U20342 (N_20342,N_17906,N_16052);
nor U20343 (N_20343,N_16199,N_16571);
nand U20344 (N_20344,N_16163,N_15985);
xnor U20345 (N_20345,N_17598,N_16068);
or U20346 (N_20346,N_16262,N_16366);
and U20347 (N_20347,N_17080,N_18195);
and U20348 (N_20348,N_15950,N_15732);
nand U20349 (N_20349,N_18232,N_16130);
and U20350 (N_20350,N_16118,N_16669);
or U20351 (N_20351,N_15929,N_16456);
or U20352 (N_20352,N_16667,N_17025);
and U20353 (N_20353,N_18333,N_15750);
nor U20354 (N_20354,N_15812,N_16738);
and U20355 (N_20355,N_18649,N_18237);
nor U20356 (N_20356,N_16213,N_16871);
or U20357 (N_20357,N_16361,N_18121);
nand U20358 (N_20358,N_15656,N_16973);
nand U20359 (N_20359,N_17522,N_17644);
or U20360 (N_20360,N_17749,N_16312);
and U20361 (N_20361,N_17410,N_16601);
or U20362 (N_20362,N_16243,N_15924);
and U20363 (N_20363,N_18674,N_17756);
nand U20364 (N_20364,N_18226,N_18706);
nor U20365 (N_20365,N_17015,N_18327);
nor U20366 (N_20366,N_16555,N_18649);
or U20367 (N_20367,N_17562,N_15656);
nand U20368 (N_20368,N_17346,N_15867);
or U20369 (N_20369,N_18143,N_18572);
and U20370 (N_20370,N_18591,N_17741);
nand U20371 (N_20371,N_16640,N_17701);
or U20372 (N_20372,N_18530,N_15904);
xor U20373 (N_20373,N_17655,N_16047);
and U20374 (N_20374,N_15981,N_18447);
nor U20375 (N_20375,N_17555,N_16492);
nor U20376 (N_20376,N_17215,N_17703);
nor U20377 (N_20377,N_18137,N_16615);
nor U20378 (N_20378,N_16954,N_16524);
nand U20379 (N_20379,N_18263,N_17824);
or U20380 (N_20380,N_16366,N_15780);
and U20381 (N_20381,N_18275,N_17683);
nor U20382 (N_20382,N_17582,N_16094);
nand U20383 (N_20383,N_18110,N_16149);
and U20384 (N_20384,N_17258,N_17567);
or U20385 (N_20385,N_17219,N_15772);
and U20386 (N_20386,N_16503,N_17790);
nand U20387 (N_20387,N_16886,N_17217);
nand U20388 (N_20388,N_17643,N_15666);
and U20389 (N_20389,N_18634,N_15898);
nand U20390 (N_20390,N_15679,N_18597);
nand U20391 (N_20391,N_18184,N_16572);
nand U20392 (N_20392,N_17558,N_18528);
nand U20393 (N_20393,N_16777,N_16288);
and U20394 (N_20394,N_16300,N_15842);
or U20395 (N_20395,N_16597,N_18263);
nor U20396 (N_20396,N_15818,N_17714);
and U20397 (N_20397,N_18466,N_15967);
or U20398 (N_20398,N_18409,N_18530);
or U20399 (N_20399,N_16958,N_18204);
or U20400 (N_20400,N_18096,N_15671);
xor U20401 (N_20401,N_18229,N_16779);
or U20402 (N_20402,N_16907,N_17063);
or U20403 (N_20403,N_17284,N_17987);
and U20404 (N_20404,N_15897,N_18307);
or U20405 (N_20405,N_16364,N_17784);
or U20406 (N_20406,N_17563,N_16774);
xnor U20407 (N_20407,N_17693,N_17026);
or U20408 (N_20408,N_17014,N_15881);
nor U20409 (N_20409,N_16264,N_16799);
nor U20410 (N_20410,N_16230,N_18519);
nor U20411 (N_20411,N_17953,N_17072);
nand U20412 (N_20412,N_16323,N_15755);
nand U20413 (N_20413,N_15626,N_16816);
or U20414 (N_20414,N_18085,N_17051);
or U20415 (N_20415,N_16156,N_17425);
nor U20416 (N_20416,N_16377,N_18144);
or U20417 (N_20417,N_17178,N_16820);
or U20418 (N_20418,N_15792,N_16913);
nand U20419 (N_20419,N_16517,N_16699);
nand U20420 (N_20420,N_18461,N_17301);
and U20421 (N_20421,N_18563,N_18180);
or U20422 (N_20422,N_16335,N_16608);
or U20423 (N_20423,N_18673,N_18042);
xor U20424 (N_20424,N_18725,N_15782);
and U20425 (N_20425,N_17703,N_18316);
nor U20426 (N_20426,N_16415,N_18681);
or U20427 (N_20427,N_16476,N_18561);
and U20428 (N_20428,N_17258,N_18589);
xnor U20429 (N_20429,N_16925,N_16277);
or U20430 (N_20430,N_18351,N_17023);
xor U20431 (N_20431,N_15926,N_16995);
nor U20432 (N_20432,N_16379,N_17278);
xnor U20433 (N_20433,N_16655,N_15778);
or U20434 (N_20434,N_17425,N_17230);
or U20435 (N_20435,N_18649,N_17365);
or U20436 (N_20436,N_16796,N_17663);
nor U20437 (N_20437,N_16375,N_18089);
nand U20438 (N_20438,N_16699,N_16414);
nor U20439 (N_20439,N_15873,N_16027);
nor U20440 (N_20440,N_16414,N_16657);
xnor U20441 (N_20441,N_16382,N_18087);
or U20442 (N_20442,N_16884,N_18507);
or U20443 (N_20443,N_16586,N_18170);
or U20444 (N_20444,N_17654,N_15696);
xnor U20445 (N_20445,N_17385,N_18263);
nand U20446 (N_20446,N_15878,N_18482);
and U20447 (N_20447,N_16119,N_16963);
and U20448 (N_20448,N_15742,N_15993);
and U20449 (N_20449,N_18126,N_18237);
xor U20450 (N_20450,N_17664,N_18622);
or U20451 (N_20451,N_17004,N_16419);
nand U20452 (N_20452,N_17317,N_17900);
and U20453 (N_20453,N_17524,N_18519);
and U20454 (N_20454,N_15975,N_17734);
or U20455 (N_20455,N_18336,N_17448);
xor U20456 (N_20456,N_17214,N_16129);
nor U20457 (N_20457,N_16164,N_16844);
nor U20458 (N_20458,N_16025,N_17074);
xor U20459 (N_20459,N_17511,N_17912);
nor U20460 (N_20460,N_16729,N_17593);
or U20461 (N_20461,N_16001,N_16924);
and U20462 (N_20462,N_17747,N_15682);
xor U20463 (N_20463,N_16277,N_17897);
nand U20464 (N_20464,N_17614,N_16027);
or U20465 (N_20465,N_17976,N_16285);
nor U20466 (N_20466,N_16160,N_17660);
or U20467 (N_20467,N_15771,N_17180);
nand U20468 (N_20468,N_18607,N_15773);
nor U20469 (N_20469,N_17228,N_17131);
nor U20470 (N_20470,N_17126,N_17501);
or U20471 (N_20471,N_16412,N_16011);
nor U20472 (N_20472,N_16003,N_16505);
xnor U20473 (N_20473,N_16227,N_17218);
or U20474 (N_20474,N_16590,N_16301);
nand U20475 (N_20475,N_15744,N_17193);
and U20476 (N_20476,N_18692,N_15908);
nand U20477 (N_20477,N_17332,N_18113);
and U20478 (N_20478,N_15928,N_18741);
or U20479 (N_20479,N_15689,N_18524);
or U20480 (N_20480,N_16129,N_15770);
nor U20481 (N_20481,N_18448,N_15890);
or U20482 (N_20482,N_18721,N_17782);
and U20483 (N_20483,N_17511,N_18438);
xor U20484 (N_20484,N_16271,N_18171);
or U20485 (N_20485,N_17641,N_18479);
nor U20486 (N_20486,N_17385,N_17050);
nor U20487 (N_20487,N_17047,N_15899);
nand U20488 (N_20488,N_16782,N_15666);
or U20489 (N_20489,N_16463,N_18073);
or U20490 (N_20490,N_18504,N_18309);
or U20491 (N_20491,N_16993,N_17417);
xnor U20492 (N_20492,N_16658,N_15887);
or U20493 (N_20493,N_16622,N_16709);
or U20494 (N_20494,N_18133,N_17250);
nand U20495 (N_20495,N_16406,N_16124);
nor U20496 (N_20496,N_16214,N_18169);
or U20497 (N_20497,N_17514,N_16638);
nand U20498 (N_20498,N_15957,N_15910);
and U20499 (N_20499,N_18317,N_17475);
or U20500 (N_20500,N_16479,N_15824);
or U20501 (N_20501,N_17124,N_15801);
or U20502 (N_20502,N_18161,N_17240);
nand U20503 (N_20503,N_17600,N_16910);
nor U20504 (N_20504,N_18058,N_17237);
or U20505 (N_20505,N_18492,N_17101);
and U20506 (N_20506,N_17696,N_18596);
nor U20507 (N_20507,N_16562,N_15693);
xor U20508 (N_20508,N_18041,N_16299);
or U20509 (N_20509,N_17246,N_17535);
nand U20510 (N_20510,N_16242,N_15667);
nor U20511 (N_20511,N_18599,N_16979);
or U20512 (N_20512,N_16854,N_16666);
nor U20513 (N_20513,N_17775,N_15842);
nand U20514 (N_20514,N_15920,N_15851);
and U20515 (N_20515,N_16113,N_16021);
or U20516 (N_20516,N_17294,N_16036);
nand U20517 (N_20517,N_17756,N_17161);
nor U20518 (N_20518,N_17216,N_16983);
or U20519 (N_20519,N_18070,N_18738);
and U20520 (N_20520,N_17313,N_17661);
and U20521 (N_20521,N_17691,N_16573);
and U20522 (N_20522,N_18182,N_16335);
nand U20523 (N_20523,N_15725,N_16412);
nand U20524 (N_20524,N_17774,N_17951);
xor U20525 (N_20525,N_16290,N_16503);
nor U20526 (N_20526,N_17267,N_16279);
nand U20527 (N_20527,N_18320,N_17990);
or U20528 (N_20528,N_18217,N_15791);
nand U20529 (N_20529,N_18621,N_17956);
nand U20530 (N_20530,N_16446,N_18056);
nor U20531 (N_20531,N_18732,N_16199);
or U20532 (N_20532,N_17476,N_18203);
xor U20533 (N_20533,N_18493,N_18104);
and U20534 (N_20534,N_17472,N_18520);
and U20535 (N_20535,N_17070,N_15950);
xnor U20536 (N_20536,N_17296,N_18314);
nor U20537 (N_20537,N_15729,N_16237);
nand U20538 (N_20538,N_18572,N_17498);
or U20539 (N_20539,N_16040,N_16798);
or U20540 (N_20540,N_16106,N_18110);
xor U20541 (N_20541,N_17497,N_18309);
nand U20542 (N_20542,N_17103,N_17071);
and U20543 (N_20543,N_16157,N_15808);
and U20544 (N_20544,N_17628,N_15949);
or U20545 (N_20545,N_17917,N_18147);
or U20546 (N_20546,N_17717,N_16625);
nor U20547 (N_20547,N_15722,N_18610);
and U20548 (N_20548,N_17589,N_18159);
nor U20549 (N_20549,N_17258,N_15957);
nand U20550 (N_20550,N_17086,N_17296);
or U20551 (N_20551,N_18604,N_18580);
nand U20552 (N_20552,N_17288,N_18236);
xor U20553 (N_20553,N_18016,N_16180);
nor U20554 (N_20554,N_17962,N_18707);
and U20555 (N_20555,N_16379,N_16275);
nand U20556 (N_20556,N_17790,N_16714);
nor U20557 (N_20557,N_16017,N_16642);
or U20558 (N_20558,N_16759,N_17016);
and U20559 (N_20559,N_15950,N_17151);
nor U20560 (N_20560,N_17523,N_17238);
or U20561 (N_20561,N_16068,N_16251);
nand U20562 (N_20562,N_18350,N_15845);
nand U20563 (N_20563,N_16640,N_18522);
nand U20564 (N_20564,N_17709,N_18394);
nor U20565 (N_20565,N_16915,N_16322);
and U20566 (N_20566,N_17581,N_16244);
and U20567 (N_20567,N_18684,N_16001);
nand U20568 (N_20568,N_17153,N_15887);
xor U20569 (N_20569,N_16121,N_18369);
or U20570 (N_20570,N_17454,N_18065);
nand U20571 (N_20571,N_18440,N_16977);
xnor U20572 (N_20572,N_17846,N_16638);
or U20573 (N_20573,N_15835,N_17901);
and U20574 (N_20574,N_16296,N_17475);
nor U20575 (N_20575,N_16875,N_17634);
nor U20576 (N_20576,N_16537,N_17374);
or U20577 (N_20577,N_16120,N_17956);
nor U20578 (N_20578,N_16402,N_16613);
nand U20579 (N_20579,N_17129,N_16376);
or U20580 (N_20580,N_16723,N_16383);
or U20581 (N_20581,N_17997,N_18165);
nand U20582 (N_20582,N_16052,N_18308);
xnor U20583 (N_20583,N_16636,N_18568);
nand U20584 (N_20584,N_16004,N_16485);
and U20585 (N_20585,N_15881,N_18070);
and U20586 (N_20586,N_17695,N_18573);
or U20587 (N_20587,N_17544,N_17645);
or U20588 (N_20588,N_16595,N_17806);
and U20589 (N_20589,N_16920,N_15812);
nor U20590 (N_20590,N_16408,N_17122);
nor U20591 (N_20591,N_15639,N_15861);
or U20592 (N_20592,N_17422,N_17053);
and U20593 (N_20593,N_16655,N_18008);
or U20594 (N_20594,N_15908,N_18695);
nand U20595 (N_20595,N_16912,N_17934);
nand U20596 (N_20596,N_16231,N_18220);
nand U20597 (N_20597,N_17307,N_17623);
or U20598 (N_20598,N_18246,N_17295);
nand U20599 (N_20599,N_16635,N_17203);
or U20600 (N_20600,N_17211,N_15940);
nand U20601 (N_20601,N_17742,N_18467);
or U20602 (N_20602,N_18678,N_16263);
nor U20603 (N_20603,N_17179,N_16150);
nor U20604 (N_20604,N_17140,N_17719);
nor U20605 (N_20605,N_15651,N_16461);
or U20606 (N_20606,N_15756,N_17609);
and U20607 (N_20607,N_16231,N_17261);
nand U20608 (N_20608,N_17439,N_17688);
nor U20609 (N_20609,N_18259,N_16109);
nor U20610 (N_20610,N_15908,N_16438);
nand U20611 (N_20611,N_16818,N_16123);
or U20612 (N_20612,N_16353,N_16856);
nand U20613 (N_20613,N_18481,N_16421);
nand U20614 (N_20614,N_15953,N_16064);
or U20615 (N_20615,N_15655,N_18460);
xor U20616 (N_20616,N_18256,N_18255);
and U20617 (N_20617,N_16940,N_17501);
or U20618 (N_20618,N_16937,N_17563);
nand U20619 (N_20619,N_15761,N_17027);
nor U20620 (N_20620,N_18191,N_18646);
or U20621 (N_20621,N_17726,N_18430);
xor U20622 (N_20622,N_16756,N_18354);
xor U20623 (N_20623,N_16201,N_17986);
nand U20624 (N_20624,N_15847,N_18683);
or U20625 (N_20625,N_18387,N_17517);
or U20626 (N_20626,N_16555,N_18407);
and U20627 (N_20627,N_16656,N_17432);
and U20628 (N_20628,N_17013,N_17369);
nor U20629 (N_20629,N_18597,N_18071);
and U20630 (N_20630,N_17854,N_16421);
or U20631 (N_20631,N_18107,N_18216);
nand U20632 (N_20632,N_17161,N_16773);
nor U20633 (N_20633,N_15808,N_18333);
and U20634 (N_20634,N_17710,N_16382);
or U20635 (N_20635,N_17517,N_17657);
or U20636 (N_20636,N_17723,N_15779);
nor U20637 (N_20637,N_15675,N_16226);
nand U20638 (N_20638,N_16284,N_18256);
xor U20639 (N_20639,N_16759,N_17619);
nand U20640 (N_20640,N_17242,N_17373);
nand U20641 (N_20641,N_17819,N_16261);
and U20642 (N_20642,N_18230,N_18065);
and U20643 (N_20643,N_16558,N_16657);
or U20644 (N_20644,N_18588,N_16997);
nand U20645 (N_20645,N_18547,N_17885);
or U20646 (N_20646,N_18142,N_17892);
and U20647 (N_20647,N_17908,N_16782);
nand U20648 (N_20648,N_16285,N_17056);
xnor U20649 (N_20649,N_17430,N_18199);
nand U20650 (N_20650,N_16618,N_17704);
nand U20651 (N_20651,N_15664,N_17546);
or U20652 (N_20652,N_17544,N_18025);
xnor U20653 (N_20653,N_18465,N_17204);
or U20654 (N_20654,N_16634,N_16166);
nand U20655 (N_20655,N_16707,N_18147);
and U20656 (N_20656,N_16953,N_16751);
or U20657 (N_20657,N_17782,N_17898);
or U20658 (N_20658,N_17190,N_18107);
or U20659 (N_20659,N_16693,N_15710);
xor U20660 (N_20660,N_18559,N_17260);
nor U20661 (N_20661,N_16554,N_15905);
nand U20662 (N_20662,N_18703,N_16256);
and U20663 (N_20663,N_17741,N_16624);
and U20664 (N_20664,N_18543,N_18703);
and U20665 (N_20665,N_16489,N_18715);
and U20666 (N_20666,N_16392,N_16860);
or U20667 (N_20667,N_15863,N_16359);
nand U20668 (N_20668,N_16915,N_18366);
or U20669 (N_20669,N_18737,N_17112);
and U20670 (N_20670,N_16056,N_17277);
and U20671 (N_20671,N_16374,N_16556);
nand U20672 (N_20672,N_15903,N_16544);
and U20673 (N_20673,N_17947,N_16135);
nor U20674 (N_20674,N_17896,N_16907);
nor U20675 (N_20675,N_17798,N_16904);
nor U20676 (N_20676,N_17733,N_17901);
or U20677 (N_20677,N_17301,N_17431);
nand U20678 (N_20678,N_18051,N_15770);
and U20679 (N_20679,N_16916,N_17549);
nand U20680 (N_20680,N_15863,N_16470);
nand U20681 (N_20681,N_17004,N_18224);
nand U20682 (N_20682,N_16550,N_18022);
xnor U20683 (N_20683,N_17626,N_17847);
and U20684 (N_20684,N_17389,N_18377);
nor U20685 (N_20685,N_16449,N_16780);
or U20686 (N_20686,N_16127,N_17511);
and U20687 (N_20687,N_18020,N_15965);
nand U20688 (N_20688,N_18136,N_16643);
or U20689 (N_20689,N_16881,N_15635);
and U20690 (N_20690,N_16583,N_18416);
nor U20691 (N_20691,N_17017,N_17645);
and U20692 (N_20692,N_17408,N_17312);
or U20693 (N_20693,N_18428,N_16537);
xnor U20694 (N_20694,N_17033,N_17472);
nor U20695 (N_20695,N_16154,N_17595);
and U20696 (N_20696,N_18437,N_18206);
nand U20697 (N_20697,N_17700,N_17765);
nand U20698 (N_20698,N_18230,N_17287);
nor U20699 (N_20699,N_16080,N_16850);
and U20700 (N_20700,N_18582,N_16280);
nor U20701 (N_20701,N_16539,N_16882);
and U20702 (N_20702,N_18213,N_16367);
nand U20703 (N_20703,N_16028,N_18263);
and U20704 (N_20704,N_18638,N_17502);
nor U20705 (N_20705,N_18225,N_18123);
nor U20706 (N_20706,N_16271,N_15966);
and U20707 (N_20707,N_15835,N_16711);
nand U20708 (N_20708,N_15952,N_16868);
nand U20709 (N_20709,N_18511,N_15707);
nor U20710 (N_20710,N_18583,N_17934);
and U20711 (N_20711,N_16401,N_16307);
or U20712 (N_20712,N_18549,N_17136);
nor U20713 (N_20713,N_15711,N_18367);
or U20714 (N_20714,N_16766,N_17538);
xnor U20715 (N_20715,N_17065,N_17850);
or U20716 (N_20716,N_17270,N_18469);
nor U20717 (N_20717,N_17839,N_18160);
or U20718 (N_20718,N_15847,N_16027);
nor U20719 (N_20719,N_18722,N_17828);
and U20720 (N_20720,N_16179,N_17907);
nor U20721 (N_20721,N_17124,N_16003);
and U20722 (N_20722,N_17592,N_16246);
and U20723 (N_20723,N_16652,N_16969);
nand U20724 (N_20724,N_16473,N_17465);
nand U20725 (N_20725,N_17185,N_16924);
and U20726 (N_20726,N_17156,N_18577);
or U20727 (N_20727,N_17418,N_15668);
nor U20728 (N_20728,N_17329,N_17255);
nand U20729 (N_20729,N_16905,N_17581);
or U20730 (N_20730,N_16681,N_17538);
xnor U20731 (N_20731,N_16182,N_16872);
or U20732 (N_20732,N_18448,N_17972);
and U20733 (N_20733,N_16414,N_17748);
nand U20734 (N_20734,N_17701,N_15663);
nand U20735 (N_20735,N_15824,N_16439);
nand U20736 (N_20736,N_15842,N_15878);
or U20737 (N_20737,N_17023,N_16662);
xor U20738 (N_20738,N_16621,N_18085);
nor U20739 (N_20739,N_16344,N_17228);
xnor U20740 (N_20740,N_16580,N_18615);
and U20741 (N_20741,N_17119,N_17141);
nor U20742 (N_20742,N_18581,N_18106);
nor U20743 (N_20743,N_17645,N_16382);
nor U20744 (N_20744,N_17793,N_16773);
nor U20745 (N_20745,N_17463,N_17065);
or U20746 (N_20746,N_17552,N_17021);
xnor U20747 (N_20747,N_18689,N_16383);
nand U20748 (N_20748,N_15904,N_16852);
xnor U20749 (N_20749,N_18563,N_17346);
nand U20750 (N_20750,N_15674,N_18358);
or U20751 (N_20751,N_15680,N_17807);
nor U20752 (N_20752,N_16177,N_17332);
nand U20753 (N_20753,N_17028,N_17342);
or U20754 (N_20754,N_15899,N_17471);
or U20755 (N_20755,N_17450,N_16611);
nor U20756 (N_20756,N_15894,N_17907);
nand U20757 (N_20757,N_18162,N_16857);
and U20758 (N_20758,N_17573,N_16399);
nand U20759 (N_20759,N_18418,N_15822);
and U20760 (N_20760,N_17501,N_15927);
and U20761 (N_20761,N_18023,N_17641);
and U20762 (N_20762,N_18587,N_16092);
or U20763 (N_20763,N_18011,N_17874);
and U20764 (N_20764,N_18132,N_17162);
nor U20765 (N_20765,N_17590,N_17457);
or U20766 (N_20766,N_16555,N_17487);
nand U20767 (N_20767,N_17271,N_17841);
nand U20768 (N_20768,N_16442,N_17724);
xnor U20769 (N_20769,N_18062,N_16657);
nand U20770 (N_20770,N_16217,N_18706);
nor U20771 (N_20771,N_15787,N_16259);
or U20772 (N_20772,N_16817,N_15724);
nor U20773 (N_20773,N_15764,N_16904);
nand U20774 (N_20774,N_16491,N_15721);
nand U20775 (N_20775,N_17525,N_16868);
and U20776 (N_20776,N_16017,N_18312);
or U20777 (N_20777,N_17931,N_15992);
or U20778 (N_20778,N_17215,N_17452);
xor U20779 (N_20779,N_16218,N_16932);
and U20780 (N_20780,N_17074,N_15942);
nor U20781 (N_20781,N_15680,N_15809);
nand U20782 (N_20782,N_16064,N_16871);
nand U20783 (N_20783,N_17476,N_17929);
nor U20784 (N_20784,N_16092,N_18671);
or U20785 (N_20785,N_16266,N_17545);
and U20786 (N_20786,N_15626,N_16852);
xnor U20787 (N_20787,N_18391,N_15756);
nand U20788 (N_20788,N_18160,N_16289);
nor U20789 (N_20789,N_18617,N_17710);
nor U20790 (N_20790,N_17668,N_17141);
and U20791 (N_20791,N_18484,N_17982);
nand U20792 (N_20792,N_18241,N_16514);
nand U20793 (N_20793,N_15946,N_18082);
nor U20794 (N_20794,N_16045,N_15741);
nor U20795 (N_20795,N_16129,N_17434);
nor U20796 (N_20796,N_16475,N_17000);
xor U20797 (N_20797,N_18181,N_18080);
nor U20798 (N_20798,N_15982,N_17071);
xnor U20799 (N_20799,N_18391,N_18323);
nor U20800 (N_20800,N_16481,N_17962);
nand U20801 (N_20801,N_16724,N_16530);
or U20802 (N_20802,N_17995,N_16361);
nor U20803 (N_20803,N_17263,N_15725);
nand U20804 (N_20804,N_16928,N_17269);
nand U20805 (N_20805,N_15950,N_18545);
xor U20806 (N_20806,N_17047,N_16641);
and U20807 (N_20807,N_16998,N_16575);
and U20808 (N_20808,N_15877,N_16809);
and U20809 (N_20809,N_16040,N_17810);
and U20810 (N_20810,N_16674,N_17963);
nor U20811 (N_20811,N_18276,N_18267);
or U20812 (N_20812,N_17481,N_16288);
nor U20813 (N_20813,N_16533,N_16277);
or U20814 (N_20814,N_16450,N_16457);
or U20815 (N_20815,N_16908,N_18020);
nand U20816 (N_20816,N_17116,N_18682);
nand U20817 (N_20817,N_17976,N_16407);
nor U20818 (N_20818,N_17151,N_18600);
xor U20819 (N_20819,N_18475,N_18240);
or U20820 (N_20820,N_15644,N_17303);
nor U20821 (N_20821,N_16497,N_18278);
xor U20822 (N_20822,N_17986,N_17718);
or U20823 (N_20823,N_17950,N_18359);
nor U20824 (N_20824,N_18577,N_18214);
or U20825 (N_20825,N_17102,N_17474);
or U20826 (N_20826,N_17521,N_16303);
nand U20827 (N_20827,N_16937,N_17488);
xnor U20828 (N_20828,N_18607,N_18394);
and U20829 (N_20829,N_16832,N_16335);
nor U20830 (N_20830,N_16005,N_18693);
nand U20831 (N_20831,N_17146,N_18460);
or U20832 (N_20832,N_17257,N_16010);
nor U20833 (N_20833,N_18087,N_15673);
nand U20834 (N_20834,N_17575,N_16646);
nand U20835 (N_20835,N_18686,N_18443);
and U20836 (N_20836,N_16107,N_18175);
and U20837 (N_20837,N_17698,N_17759);
nand U20838 (N_20838,N_17859,N_17134);
or U20839 (N_20839,N_17603,N_17679);
or U20840 (N_20840,N_16576,N_16747);
and U20841 (N_20841,N_15863,N_17207);
xnor U20842 (N_20842,N_16623,N_16962);
and U20843 (N_20843,N_17045,N_15980);
and U20844 (N_20844,N_16180,N_17929);
nand U20845 (N_20845,N_16208,N_16003);
xnor U20846 (N_20846,N_18590,N_17653);
nor U20847 (N_20847,N_16523,N_18104);
nor U20848 (N_20848,N_15726,N_16910);
or U20849 (N_20849,N_18526,N_17205);
and U20850 (N_20850,N_17671,N_17163);
nor U20851 (N_20851,N_18662,N_17379);
or U20852 (N_20852,N_15748,N_15888);
or U20853 (N_20853,N_17922,N_15701);
and U20854 (N_20854,N_16025,N_16531);
or U20855 (N_20855,N_16768,N_18002);
or U20856 (N_20856,N_18249,N_16769);
and U20857 (N_20857,N_18190,N_17541);
nand U20858 (N_20858,N_17068,N_15782);
or U20859 (N_20859,N_15733,N_16129);
and U20860 (N_20860,N_15938,N_16617);
nor U20861 (N_20861,N_17978,N_16565);
or U20862 (N_20862,N_16496,N_16217);
and U20863 (N_20863,N_15695,N_17205);
nor U20864 (N_20864,N_16618,N_17027);
xnor U20865 (N_20865,N_15948,N_18484);
or U20866 (N_20866,N_16736,N_17408);
or U20867 (N_20867,N_18166,N_18489);
nand U20868 (N_20868,N_15943,N_17826);
nor U20869 (N_20869,N_17940,N_18233);
nand U20870 (N_20870,N_17946,N_15996);
or U20871 (N_20871,N_17287,N_16336);
and U20872 (N_20872,N_18520,N_18509);
nor U20873 (N_20873,N_16768,N_18582);
nand U20874 (N_20874,N_16350,N_16644);
xnor U20875 (N_20875,N_16050,N_17032);
nand U20876 (N_20876,N_15897,N_16855);
nand U20877 (N_20877,N_18388,N_16189);
or U20878 (N_20878,N_18310,N_15848);
and U20879 (N_20879,N_17007,N_17065);
xnor U20880 (N_20880,N_17722,N_18641);
xor U20881 (N_20881,N_17334,N_17034);
nor U20882 (N_20882,N_17942,N_17661);
xor U20883 (N_20883,N_18124,N_17082);
or U20884 (N_20884,N_16815,N_16993);
nor U20885 (N_20885,N_16203,N_16204);
nor U20886 (N_20886,N_16144,N_17689);
and U20887 (N_20887,N_16236,N_16213);
and U20888 (N_20888,N_18046,N_16737);
nand U20889 (N_20889,N_17648,N_16937);
and U20890 (N_20890,N_16389,N_17471);
nand U20891 (N_20891,N_17657,N_15788);
and U20892 (N_20892,N_16598,N_17067);
or U20893 (N_20893,N_18004,N_16196);
or U20894 (N_20894,N_18067,N_17829);
nand U20895 (N_20895,N_17395,N_17653);
nor U20896 (N_20896,N_15966,N_17981);
nor U20897 (N_20897,N_16434,N_18237);
nand U20898 (N_20898,N_16454,N_17596);
or U20899 (N_20899,N_17379,N_18735);
or U20900 (N_20900,N_16315,N_17079);
and U20901 (N_20901,N_17529,N_16420);
nand U20902 (N_20902,N_18449,N_18415);
and U20903 (N_20903,N_18732,N_16117);
nor U20904 (N_20904,N_18553,N_17993);
and U20905 (N_20905,N_18012,N_16522);
nor U20906 (N_20906,N_17801,N_16386);
and U20907 (N_20907,N_16075,N_15951);
xnor U20908 (N_20908,N_17219,N_17495);
or U20909 (N_20909,N_18514,N_18538);
nor U20910 (N_20910,N_16678,N_15765);
nand U20911 (N_20911,N_16990,N_18219);
and U20912 (N_20912,N_18146,N_16493);
nor U20913 (N_20913,N_16239,N_16005);
and U20914 (N_20914,N_18030,N_16605);
or U20915 (N_20915,N_18482,N_17907);
and U20916 (N_20916,N_16388,N_16534);
nor U20917 (N_20917,N_17239,N_16207);
nand U20918 (N_20918,N_16525,N_18732);
nor U20919 (N_20919,N_18155,N_17631);
and U20920 (N_20920,N_18521,N_16024);
nor U20921 (N_20921,N_18088,N_17025);
xnor U20922 (N_20922,N_16544,N_16421);
and U20923 (N_20923,N_15865,N_15723);
nand U20924 (N_20924,N_16529,N_16057);
xnor U20925 (N_20925,N_16781,N_18073);
or U20926 (N_20926,N_17169,N_16932);
or U20927 (N_20927,N_17220,N_15832);
nand U20928 (N_20928,N_17270,N_16455);
or U20929 (N_20929,N_17037,N_16768);
and U20930 (N_20930,N_17963,N_17909);
nand U20931 (N_20931,N_16257,N_18249);
nor U20932 (N_20932,N_16864,N_16537);
or U20933 (N_20933,N_18075,N_16551);
xnor U20934 (N_20934,N_16113,N_18267);
nand U20935 (N_20935,N_17229,N_16739);
and U20936 (N_20936,N_16530,N_17600);
and U20937 (N_20937,N_17219,N_18430);
and U20938 (N_20938,N_16545,N_17312);
nor U20939 (N_20939,N_17755,N_16784);
and U20940 (N_20940,N_15751,N_17937);
nand U20941 (N_20941,N_15693,N_18425);
xnor U20942 (N_20942,N_17620,N_18040);
nand U20943 (N_20943,N_17012,N_17828);
xor U20944 (N_20944,N_15965,N_16509);
or U20945 (N_20945,N_18612,N_17169);
and U20946 (N_20946,N_16619,N_17325);
nor U20947 (N_20947,N_15871,N_16045);
nor U20948 (N_20948,N_18611,N_16791);
or U20949 (N_20949,N_15760,N_18483);
and U20950 (N_20950,N_18154,N_16826);
and U20951 (N_20951,N_15667,N_16602);
nor U20952 (N_20952,N_15852,N_18600);
and U20953 (N_20953,N_16592,N_17261);
nand U20954 (N_20954,N_18042,N_18288);
or U20955 (N_20955,N_18343,N_18000);
nor U20956 (N_20956,N_18162,N_15942);
xnor U20957 (N_20957,N_16726,N_17703);
and U20958 (N_20958,N_18330,N_16593);
or U20959 (N_20959,N_17929,N_18480);
and U20960 (N_20960,N_18348,N_15662);
xnor U20961 (N_20961,N_17271,N_18664);
nor U20962 (N_20962,N_18088,N_16128);
and U20963 (N_20963,N_17611,N_17206);
or U20964 (N_20964,N_16069,N_16923);
xnor U20965 (N_20965,N_15944,N_17846);
nand U20966 (N_20966,N_17193,N_16249);
or U20967 (N_20967,N_17821,N_16958);
and U20968 (N_20968,N_18448,N_17524);
and U20969 (N_20969,N_16106,N_18010);
and U20970 (N_20970,N_18735,N_16619);
nor U20971 (N_20971,N_16761,N_18662);
xnor U20972 (N_20972,N_17016,N_16316);
nand U20973 (N_20973,N_16547,N_18355);
or U20974 (N_20974,N_18734,N_15633);
nor U20975 (N_20975,N_16925,N_17526);
and U20976 (N_20976,N_16295,N_16174);
nand U20977 (N_20977,N_17969,N_17977);
nor U20978 (N_20978,N_18666,N_17849);
xor U20979 (N_20979,N_18217,N_17890);
nor U20980 (N_20980,N_16589,N_18198);
or U20981 (N_20981,N_17700,N_17242);
or U20982 (N_20982,N_16062,N_17470);
or U20983 (N_20983,N_18064,N_16226);
nor U20984 (N_20984,N_15837,N_15673);
nor U20985 (N_20985,N_16161,N_18180);
or U20986 (N_20986,N_18645,N_16958);
nand U20987 (N_20987,N_16498,N_16648);
nand U20988 (N_20988,N_18235,N_16580);
or U20989 (N_20989,N_17546,N_16009);
and U20990 (N_20990,N_18009,N_15712);
nor U20991 (N_20991,N_17501,N_17800);
or U20992 (N_20992,N_17375,N_16994);
nor U20993 (N_20993,N_17996,N_17286);
and U20994 (N_20994,N_15932,N_16941);
and U20995 (N_20995,N_18054,N_16970);
nor U20996 (N_20996,N_15889,N_17236);
and U20997 (N_20997,N_16388,N_18499);
nor U20998 (N_20998,N_16397,N_17499);
nand U20999 (N_20999,N_16079,N_16978);
or U21000 (N_21000,N_18259,N_16031);
or U21001 (N_21001,N_17148,N_16713);
nand U21002 (N_21002,N_15991,N_18220);
nand U21003 (N_21003,N_18659,N_16624);
nor U21004 (N_21004,N_16204,N_18380);
and U21005 (N_21005,N_15671,N_16097);
and U21006 (N_21006,N_18402,N_16835);
nor U21007 (N_21007,N_18427,N_17788);
or U21008 (N_21008,N_15929,N_16307);
xor U21009 (N_21009,N_15951,N_17018);
and U21010 (N_21010,N_15670,N_15825);
nor U21011 (N_21011,N_18354,N_17590);
and U21012 (N_21012,N_17648,N_18265);
or U21013 (N_21013,N_17919,N_16137);
and U21014 (N_21014,N_16808,N_18273);
nand U21015 (N_21015,N_16254,N_16518);
and U21016 (N_21016,N_18627,N_16875);
or U21017 (N_21017,N_15837,N_16533);
and U21018 (N_21018,N_16172,N_17422);
nor U21019 (N_21019,N_18178,N_15883);
or U21020 (N_21020,N_15681,N_17108);
nand U21021 (N_21021,N_16119,N_15846);
xor U21022 (N_21022,N_15938,N_17749);
nor U21023 (N_21023,N_16181,N_17464);
nor U21024 (N_21024,N_17397,N_15739);
nand U21025 (N_21025,N_16707,N_15954);
and U21026 (N_21026,N_17396,N_17173);
or U21027 (N_21027,N_17957,N_18382);
and U21028 (N_21028,N_18571,N_16679);
or U21029 (N_21029,N_15819,N_17689);
xnor U21030 (N_21030,N_17064,N_16310);
or U21031 (N_21031,N_17465,N_16214);
nor U21032 (N_21032,N_16225,N_17624);
or U21033 (N_21033,N_18338,N_18347);
nor U21034 (N_21034,N_16711,N_17394);
nand U21035 (N_21035,N_16210,N_16681);
or U21036 (N_21036,N_16360,N_16592);
and U21037 (N_21037,N_18186,N_18275);
or U21038 (N_21038,N_17309,N_18225);
or U21039 (N_21039,N_17082,N_17713);
nor U21040 (N_21040,N_16725,N_17318);
and U21041 (N_21041,N_16081,N_16288);
or U21042 (N_21042,N_16750,N_15783);
nor U21043 (N_21043,N_16847,N_16594);
or U21044 (N_21044,N_16884,N_16970);
or U21045 (N_21045,N_17473,N_17783);
nand U21046 (N_21046,N_15948,N_16522);
nand U21047 (N_21047,N_17213,N_16300);
xnor U21048 (N_21048,N_16064,N_18548);
nor U21049 (N_21049,N_16251,N_16893);
nor U21050 (N_21050,N_15762,N_18701);
or U21051 (N_21051,N_17208,N_15760);
or U21052 (N_21052,N_15774,N_16275);
and U21053 (N_21053,N_18583,N_17508);
or U21054 (N_21054,N_16509,N_16161);
nand U21055 (N_21055,N_15796,N_18077);
or U21056 (N_21056,N_17779,N_18708);
nor U21057 (N_21057,N_18204,N_18483);
xnor U21058 (N_21058,N_16560,N_17414);
nor U21059 (N_21059,N_16225,N_17444);
nand U21060 (N_21060,N_16880,N_18675);
or U21061 (N_21061,N_15941,N_18565);
and U21062 (N_21062,N_18641,N_16806);
and U21063 (N_21063,N_16378,N_17291);
and U21064 (N_21064,N_18527,N_17182);
xor U21065 (N_21065,N_16960,N_17506);
and U21066 (N_21066,N_16796,N_15912);
and U21067 (N_21067,N_16910,N_15809);
nand U21068 (N_21068,N_16356,N_16798);
nand U21069 (N_21069,N_18482,N_15727);
xor U21070 (N_21070,N_15957,N_17069);
and U21071 (N_21071,N_15833,N_18683);
and U21072 (N_21072,N_17734,N_16262);
and U21073 (N_21073,N_17191,N_16589);
or U21074 (N_21074,N_16878,N_17915);
or U21075 (N_21075,N_16427,N_15637);
xnor U21076 (N_21076,N_15956,N_17484);
or U21077 (N_21077,N_18610,N_18639);
nand U21078 (N_21078,N_17691,N_17743);
nor U21079 (N_21079,N_18690,N_16151);
nor U21080 (N_21080,N_17081,N_18705);
xnor U21081 (N_21081,N_16315,N_16745);
or U21082 (N_21082,N_18489,N_16987);
xor U21083 (N_21083,N_15787,N_17313);
xnor U21084 (N_21084,N_16624,N_16637);
or U21085 (N_21085,N_17895,N_17683);
and U21086 (N_21086,N_18195,N_18451);
or U21087 (N_21087,N_16417,N_16004);
and U21088 (N_21088,N_16378,N_16118);
nor U21089 (N_21089,N_16525,N_16306);
nor U21090 (N_21090,N_16340,N_16589);
nor U21091 (N_21091,N_16668,N_17196);
xnor U21092 (N_21092,N_16322,N_18309);
and U21093 (N_21093,N_17518,N_17345);
or U21094 (N_21094,N_16848,N_16405);
or U21095 (N_21095,N_17066,N_16112);
xnor U21096 (N_21096,N_15917,N_16368);
or U21097 (N_21097,N_16898,N_15917);
or U21098 (N_21098,N_17696,N_18720);
nor U21099 (N_21099,N_17871,N_16744);
nor U21100 (N_21100,N_17429,N_18184);
xnor U21101 (N_21101,N_17865,N_17380);
or U21102 (N_21102,N_17533,N_16933);
and U21103 (N_21103,N_17570,N_16216);
nand U21104 (N_21104,N_17469,N_16201);
or U21105 (N_21105,N_18725,N_15928);
nand U21106 (N_21106,N_18279,N_18424);
nor U21107 (N_21107,N_15813,N_18644);
or U21108 (N_21108,N_18395,N_17384);
nand U21109 (N_21109,N_16331,N_17729);
nand U21110 (N_21110,N_16251,N_16220);
or U21111 (N_21111,N_17836,N_15660);
or U21112 (N_21112,N_16107,N_16879);
nand U21113 (N_21113,N_18577,N_17240);
or U21114 (N_21114,N_16474,N_16550);
and U21115 (N_21115,N_18117,N_18150);
or U21116 (N_21116,N_17418,N_16682);
nand U21117 (N_21117,N_17857,N_15992);
xnor U21118 (N_21118,N_16655,N_17300);
nor U21119 (N_21119,N_18704,N_17509);
and U21120 (N_21120,N_16588,N_17965);
or U21121 (N_21121,N_16691,N_15771);
nor U21122 (N_21122,N_17077,N_16643);
nand U21123 (N_21123,N_16065,N_16944);
nor U21124 (N_21124,N_17051,N_16917);
or U21125 (N_21125,N_18062,N_16759);
nor U21126 (N_21126,N_16784,N_16934);
nor U21127 (N_21127,N_18344,N_18072);
and U21128 (N_21128,N_16666,N_17322);
nor U21129 (N_21129,N_17361,N_17372);
nor U21130 (N_21130,N_17369,N_17081);
nor U21131 (N_21131,N_15655,N_17161);
nor U21132 (N_21132,N_18586,N_15867);
xor U21133 (N_21133,N_16902,N_16773);
or U21134 (N_21134,N_16132,N_16585);
and U21135 (N_21135,N_18017,N_17825);
or U21136 (N_21136,N_16493,N_15868);
xnor U21137 (N_21137,N_15908,N_16230);
nand U21138 (N_21138,N_17595,N_18431);
nor U21139 (N_21139,N_16094,N_15632);
nand U21140 (N_21140,N_15692,N_17323);
xnor U21141 (N_21141,N_15764,N_17053);
nand U21142 (N_21142,N_15689,N_17627);
or U21143 (N_21143,N_16396,N_18370);
nor U21144 (N_21144,N_17172,N_16966);
nand U21145 (N_21145,N_18678,N_17264);
nor U21146 (N_21146,N_17074,N_17519);
nand U21147 (N_21147,N_17499,N_16969);
or U21148 (N_21148,N_17637,N_18603);
nor U21149 (N_21149,N_18418,N_16582);
nand U21150 (N_21150,N_15954,N_16691);
and U21151 (N_21151,N_15695,N_17541);
nor U21152 (N_21152,N_16601,N_18110);
or U21153 (N_21153,N_16764,N_17627);
xnor U21154 (N_21154,N_18126,N_16031);
nand U21155 (N_21155,N_18515,N_16117);
or U21156 (N_21156,N_18700,N_16654);
nor U21157 (N_21157,N_15951,N_15759);
nor U21158 (N_21158,N_15955,N_15695);
nor U21159 (N_21159,N_17885,N_17464);
nor U21160 (N_21160,N_17003,N_18199);
or U21161 (N_21161,N_16566,N_17508);
nor U21162 (N_21162,N_17202,N_16770);
and U21163 (N_21163,N_18290,N_18317);
and U21164 (N_21164,N_15819,N_18109);
nand U21165 (N_21165,N_17047,N_16897);
nor U21166 (N_21166,N_15764,N_15715);
or U21167 (N_21167,N_15642,N_16818);
and U21168 (N_21168,N_15626,N_15896);
or U21169 (N_21169,N_18265,N_16872);
or U21170 (N_21170,N_17641,N_18302);
nor U21171 (N_21171,N_17956,N_16918);
and U21172 (N_21172,N_17609,N_18013);
and U21173 (N_21173,N_17307,N_17850);
or U21174 (N_21174,N_17645,N_17875);
and U21175 (N_21175,N_16576,N_16700);
nor U21176 (N_21176,N_15997,N_18270);
nor U21177 (N_21177,N_18711,N_17268);
xnor U21178 (N_21178,N_17971,N_18529);
and U21179 (N_21179,N_18640,N_18562);
nor U21180 (N_21180,N_18332,N_17675);
nor U21181 (N_21181,N_18243,N_15910);
or U21182 (N_21182,N_18163,N_16573);
nor U21183 (N_21183,N_16611,N_17953);
and U21184 (N_21184,N_17025,N_17677);
nand U21185 (N_21185,N_18599,N_18324);
and U21186 (N_21186,N_18202,N_17962);
and U21187 (N_21187,N_16428,N_17941);
nand U21188 (N_21188,N_18324,N_18517);
nand U21189 (N_21189,N_15680,N_18245);
xor U21190 (N_21190,N_16566,N_18250);
nor U21191 (N_21191,N_17937,N_15669);
and U21192 (N_21192,N_17816,N_18621);
and U21193 (N_21193,N_16368,N_16275);
or U21194 (N_21194,N_18328,N_16039);
and U21195 (N_21195,N_17205,N_16074);
nor U21196 (N_21196,N_17201,N_17801);
xnor U21197 (N_21197,N_16242,N_17696);
and U21198 (N_21198,N_17249,N_16820);
nor U21199 (N_21199,N_17339,N_17643);
and U21200 (N_21200,N_17118,N_17160);
xor U21201 (N_21201,N_15840,N_17145);
and U21202 (N_21202,N_17226,N_17236);
or U21203 (N_21203,N_16416,N_16155);
xor U21204 (N_21204,N_18489,N_18628);
xnor U21205 (N_21205,N_17336,N_17751);
and U21206 (N_21206,N_17026,N_16688);
and U21207 (N_21207,N_17204,N_15947);
nor U21208 (N_21208,N_18068,N_16058);
and U21209 (N_21209,N_16403,N_18167);
nor U21210 (N_21210,N_17741,N_17218);
nand U21211 (N_21211,N_17365,N_18687);
nand U21212 (N_21212,N_18298,N_17246);
nand U21213 (N_21213,N_17623,N_17471);
and U21214 (N_21214,N_18367,N_17485);
or U21215 (N_21215,N_17775,N_16296);
nand U21216 (N_21216,N_18683,N_16040);
xnor U21217 (N_21217,N_18638,N_15628);
nor U21218 (N_21218,N_17028,N_16114);
or U21219 (N_21219,N_17836,N_16632);
nand U21220 (N_21220,N_16364,N_18455);
nor U21221 (N_21221,N_18038,N_17061);
nand U21222 (N_21222,N_18665,N_17325);
nor U21223 (N_21223,N_18399,N_18625);
nand U21224 (N_21224,N_18635,N_16858);
and U21225 (N_21225,N_18378,N_15890);
and U21226 (N_21226,N_18573,N_17325);
or U21227 (N_21227,N_17062,N_18174);
and U21228 (N_21228,N_18280,N_16508);
nand U21229 (N_21229,N_15706,N_17084);
and U21230 (N_21230,N_16900,N_16586);
and U21231 (N_21231,N_18059,N_16357);
and U21232 (N_21232,N_16827,N_17511);
and U21233 (N_21233,N_16558,N_16631);
or U21234 (N_21234,N_15828,N_17056);
or U21235 (N_21235,N_17874,N_18523);
nor U21236 (N_21236,N_15834,N_15820);
or U21237 (N_21237,N_15840,N_16207);
or U21238 (N_21238,N_16133,N_18249);
nand U21239 (N_21239,N_18561,N_18443);
and U21240 (N_21240,N_18077,N_16368);
and U21241 (N_21241,N_16266,N_16669);
nor U21242 (N_21242,N_18541,N_17990);
nor U21243 (N_21243,N_17862,N_18018);
nor U21244 (N_21244,N_15816,N_17920);
nor U21245 (N_21245,N_18018,N_16556);
nand U21246 (N_21246,N_18527,N_15826);
xnor U21247 (N_21247,N_18105,N_18247);
xnor U21248 (N_21248,N_17310,N_17987);
nand U21249 (N_21249,N_16156,N_17759);
or U21250 (N_21250,N_16610,N_18471);
nor U21251 (N_21251,N_18212,N_17070);
nand U21252 (N_21252,N_16549,N_17326);
or U21253 (N_21253,N_18289,N_16728);
nand U21254 (N_21254,N_18339,N_17891);
and U21255 (N_21255,N_15947,N_18590);
nor U21256 (N_21256,N_17925,N_17894);
nor U21257 (N_21257,N_15968,N_16745);
xor U21258 (N_21258,N_17308,N_17603);
and U21259 (N_21259,N_15933,N_17543);
nor U21260 (N_21260,N_18467,N_15819);
nor U21261 (N_21261,N_16242,N_17459);
and U21262 (N_21262,N_17464,N_18130);
nand U21263 (N_21263,N_17804,N_16737);
nor U21264 (N_21264,N_18551,N_18594);
nor U21265 (N_21265,N_15942,N_16187);
nor U21266 (N_21266,N_17003,N_16997);
xor U21267 (N_21267,N_18391,N_15880);
xnor U21268 (N_21268,N_17534,N_15791);
nor U21269 (N_21269,N_18190,N_18084);
nand U21270 (N_21270,N_17922,N_17867);
nor U21271 (N_21271,N_16384,N_18405);
or U21272 (N_21272,N_16612,N_15899);
nor U21273 (N_21273,N_17687,N_17819);
or U21274 (N_21274,N_17161,N_18204);
or U21275 (N_21275,N_18651,N_17687);
and U21276 (N_21276,N_17222,N_15817);
nand U21277 (N_21277,N_17969,N_17232);
nand U21278 (N_21278,N_18432,N_16923);
or U21279 (N_21279,N_16157,N_18182);
and U21280 (N_21280,N_18179,N_17465);
xnor U21281 (N_21281,N_15737,N_18097);
nand U21282 (N_21282,N_18138,N_15804);
and U21283 (N_21283,N_17413,N_16082);
nor U21284 (N_21284,N_17903,N_17525);
and U21285 (N_21285,N_17952,N_18347);
nand U21286 (N_21286,N_17854,N_17893);
nand U21287 (N_21287,N_17703,N_17123);
and U21288 (N_21288,N_17518,N_18028);
nand U21289 (N_21289,N_16426,N_18254);
nor U21290 (N_21290,N_18609,N_17810);
nor U21291 (N_21291,N_18385,N_18681);
nand U21292 (N_21292,N_18565,N_17999);
or U21293 (N_21293,N_16345,N_15812);
nor U21294 (N_21294,N_17644,N_17759);
xor U21295 (N_21295,N_18280,N_17954);
or U21296 (N_21296,N_18582,N_16780);
nand U21297 (N_21297,N_17468,N_15827);
or U21298 (N_21298,N_16112,N_16963);
nor U21299 (N_21299,N_16592,N_16530);
and U21300 (N_21300,N_16454,N_18054);
or U21301 (N_21301,N_18577,N_16980);
xnor U21302 (N_21302,N_15720,N_17634);
nor U21303 (N_21303,N_17750,N_17954);
nand U21304 (N_21304,N_16585,N_17594);
and U21305 (N_21305,N_16329,N_18334);
nor U21306 (N_21306,N_17281,N_16442);
xnor U21307 (N_21307,N_17746,N_18693);
or U21308 (N_21308,N_16416,N_16694);
nand U21309 (N_21309,N_18513,N_17500);
xnor U21310 (N_21310,N_18526,N_17745);
nand U21311 (N_21311,N_15924,N_16313);
xnor U21312 (N_21312,N_15771,N_17985);
or U21313 (N_21313,N_18476,N_15697);
nor U21314 (N_21314,N_16448,N_17970);
or U21315 (N_21315,N_18246,N_16669);
or U21316 (N_21316,N_16789,N_16160);
or U21317 (N_21317,N_15844,N_18398);
nand U21318 (N_21318,N_17686,N_16475);
nand U21319 (N_21319,N_18351,N_15721);
nor U21320 (N_21320,N_17992,N_16720);
nor U21321 (N_21321,N_16542,N_15727);
xor U21322 (N_21322,N_17850,N_17554);
and U21323 (N_21323,N_16410,N_15919);
and U21324 (N_21324,N_15899,N_18371);
or U21325 (N_21325,N_18267,N_18673);
or U21326 (N_21326,N_16067,N_17002);
and U21327 (N_21327,N_16821,N_16898);
and U21328 (N_21328,N_17167,N_18553);
nor U21329 (N_21329,N_15796,N_16328);
xor U21330 (N_21330,N_16164,N_16116);
nor U21331 (N_21331,N_16227,N_16279);
or U21332 (N_21332,N_17364,N_17084);
nor U21333 (N_21333,N_17575,N_15659);
nor U21334 (N_21334,N_17876,N_18034);
xnor U21335 (N_21335,N_17620,N_16184);
nand U21336 (N_21336,N_16802,N_17531);
xnor U21337 (N_21337,N_16610,N_17701);
and U21338 (N_21338,N_16846,N_16224);
xor U21339 (N_21339,N_18433,N_15973);
nor U21340 (N_21340,N_16656,N_17195);
nor U21341 (N_21341,N_16412,N_16907);
xnor U21342 (N_21342,N_17171,N_16019);
and U21343 (N_21343,N_16784,N_16921);
and U21344 (N_21344,N_15794,N_18396);
and U21345 (N_21345,N_18704,N_17108);
nand U21346 (N_21346,N_16248,N_18211);
nor U21347 (N_21347,N_17751,N_17508);
nand U21348 (N_21348,N_17165,N_16219);
and U21349 (N_21349,N_15827,N_17071);
and U21350 (N_21350,N_16353,N_15626);
nand U21351 (N_21351,N_17116,N_15912);
or U21352 (N_21352,N_18059,N_16228);
and U21353 (N_21353,N_16964,N_18652);
nand U21354 (N_21354,N_16299,N_17434);
nor U21355 (N_21355,N_18302,N_17336);
and U21356 (N_21356,N_15841,N_17773);
or U21357 (N_21357,N_16053,N_16777);
nand U21358 (N_21358,N_15807,N_16561);
and U21359 (N_21359,N_17923,N_16687);
or U21360 (N_21360,N_18695,N_17594);
and U21361 (N_21361,N_17293,N_17213);
nor U21362 (N_21362,N_17503,N_16960);
nand U21363 (N_21363,N_16716,N_17245);
or U21364 (N_21364,N_16939,N_17965);
or U21365 (N_21365,N_16829,N_16465);
nand U21366 (N_21366,N_17389,N_18436);
and U21367 (N_21367,N_16424,N_17434);
nand U21368 (N_21368,N_16401,N_18604);
nor U21369 (N_21369,N_16424,N_16704);
and U21370 (N_21370,N_17654,N_15746);
nor U21371 (N_21371,N_15831,N_16001);
nor U21372 (N_21372,N_16019,N_17128);
and U21373 (N_21373,N_16332,N_17589);
or U21374 (N_21374,N_16667,N_17973);
and U21375 (N_21375,N_17144,N_15726);
nor U21376 (N_21376,N_18705,N_17765);
and U21377 (N_21377,N_17513,N_16374);
nand U21378 (N_21378,N_17486,N_18452);
or U21379 (N_21379,N_15625,N_18278);
nand U21380 (N_21380,N_16912,N_18194);
nand U21381 (N_21381,N_16068,N_17015);
nand U21382 (N_21382,N_17499,N_15907);
nand U21383 (N_21383,N_17480,N_17874);
or U21384 (N_21384,N_15840,N_15843);
nor U21385 (N_21385,N_17885,N_16527);
nor U21386 (N_21386,N_16759,N_16701);
and U21387 (N_21387,N_15904,N_17833);
nand U21388 (N_21388,N_16941,N_18331);
nor U21389 (N_21389,N_18450,N_17304);
and U21390 (N_21390,N_16125,N_18652);
nand U21391 (N_21391,N_16010,N_17761);
and U21392 (N_21392,N_15933,N_15801);
nand U21393 (N_21393,N_17471,N_18358);
xnor U21394 (N_21394,N_18510,N_18062);
and U21395 (N_21395,N_17150,N_18680);
xor U21396 (N_21396,N_16109,N_18428);
nand U21397 (N_21397,N_16708,N_17542);
and U21398 (N_21398,N_16144,N_16057);
nor U21399 (N_21399,N_18316,N_15850);
or U21400 (N_21400,N_17077,N_17582);
or U21401 (N_21401,N_17387,N_17134);
or U21402 (N_21402,N_16244,N_18650);
and U21403 (N_21403,N_17657,N_18665);
xor U21404 (N_21404,N_18257,N_16277);
or U21405 (N_21405,N_16395,N_17599);
or U21406 (N_21406,N_16750,N_15893);
nor U21407 (N_21407,N_15801,N_17808);
or U21408 (N_21408,N_16892,N_17805);
xor U21409 (N_21409,N_17486,N_16219);
nor U21410 (N_21410,N_18568,N_16448);
and U21411 (N_21411,N_15857,N_17835);
and U21412 (N_21412,N_15875,N_15934);
or U21413 (N_21413,N_18377,N_17173);
nand U21414 (N_21414,N_17661,N_18591);
and U21415 (N_21415,N_18541,N_17943);
or U21416 (N_21416,N_18494,N_16403);
or U21417 (N_21417,N_17492,N_17600);
nor U21418 (N_21418,N_16835,N_15749);
and U21419 (N_21419,N_18689,N_16977);
and U21420 (N_21420,N_15714,N_17437);
and U21421 (N_21421,N_17085,N_16105);
xnor U21422 (N_21422,N_17421,N_16854);
or U21423 (N_21423,N_15936,N_18135);
nor U21424 (N_21424,N_15766,N_17802);
nand U21425 (N_21425,N_15966,N_18746);
nor U21426 (N_21426,N_17677,N_15765);
nand U21427 (N_21427,N_16793,N_15633);
nor U21428 (N_21428,N_16058,N_18470);
nand U21429 (N_21429,N_17369,N_18540);
nand U21430 (N_21430,N_18187,N_17907);
nand U21431 (N_21431,N_17086,N_17590);
nand U21432 (N_21432,N_17968,N_18311);
and U21433 (N_21433,N_18061,N_18704);
nand U21434 (N_21434,N_18568,N_16214);
nor U21435 (N_21435,N_17225,N_15714);
nor U21436 (N_21436,N_17858,N_17535);
nor U21437 (N_21437,N_16115,N_17616);
nand U21438 (N_21438,N_17942,N_18655);
and U21439 (N_21439,N_17239,N_17947);
nor U21440 (N_21440,N_18123,N_15663);
or U21441 (N_21441,N_18081,N_16046);
and U21442 (N_21442,N_16332,N_17225);
nor U21443 (N_21443,N_17679,N_16568);
xnor U21444 (N_21444,N_17370,N_16422);
and U21445 (N_21445,N_15839,N_17664);
xor U21446 (N_21446,N_16636,N_16817);
nand U21447 (N_21447,N_16284,N_18267);
nand U21448 (N_21448,N_16723,N_15714);
or U21449 (N_21449,N_16249,N_16339);
nand U21450 (N_21450,N_17815,N_15903);
nand U21451 (N_21451,N_18003,N_18627);
xor U21452 (N_21452,N_18230,N_17493);
or U21453 (N_21453,N_18326,N_18223);
or U21454 (N_21454,N_16171,N_18250);
or U21455 (N_21455,N_15889,N_16245);
nor U21456 (N_21456,N_16368,N_16458);
nor U21457 (N_21457,N_16660,N_17700);
or U21458 (N_21458,N_17583,N_17166);
nand U21459 (N_21459,N_18452,N_17763);
and U21460 (N_21460,N_17972,N_17319);
or U21461 (N_21461,N_18148,N_17762);
xor U21462 (N_21462,N_18415,N_16811);
or U21463 (N_21463,N_17176,N_17627);
and U21464 (N_21464,N_17332,N_16733);
nor U21465 (N_21465,N_15952,N_18677);
nor U21466 (N_21466,N_15791,N_15999);
nand U21467 (N_21467,N_18358,N_16516);
xor U21468 (N_21468,N_18020,N_18387);
nor U21469 (N_21469,N_16955,N_17518);
and U21470 (N_21470,N_18253,N_18297);
xnor U21471 (N_21471,N_18538,N_16122);
and U21472 (N_21472,N_17201,N_16274);
or U21473 (N_21473,N_17006,N_16676);
and U21474 (N_21474,N_16972,N_15873);
nor U21475 (N_21475,N_18367,N_15868);
nor U21476 (N_21476,N_17922,N_18340);
nand U21477 (N_21477,N_16101,N_18589);
nor U21478 (N_21478,N_18452,N_16196);
or U21479 (N_21479,N_16855,N_16155);
and U21480 (N_21480,N_18488,N_16237);
nand U21481 (N_21481,N_16365,N_16819);
and U21482 (N_21482,N_17432,N_16647);
nor U21483 (N_21483,N_18013,N_17773);
nor U21484 (N_21484,N_17632,N_16837);
nor U21485 (N_21485,N_17643,N_17192);
nand U21486 (N_21486,N_16025,N_16072);
or U21487 (N_21487,N_18275,N_17389);
and U21488 (N_21488,N_17474,N_17332);
and U21489 (N_21489,N_17745,N_17307);
or U21490 (N_21490,N_18010,N_17990);
or U21491 (N_21491,N_16329,N_17327);
nor U21492 (N_21492,N_17015,N_17309);
nand U21493 (N_21493,N_18593,N_17756);
nor U21494 (N_21494,N_18474,N_18242);
or U21495 (N_21495,N_15776,N_16344);
or U21496 (N_21496,N_16660,N_17798);
or U21497 (N_21497,N_18579,N_17672);
xnor U21498 (N_21498,N_16046,N_17029);
nor U21499 (N_21499,N_16178,N_17250);
and U21500 (N_21500,N_17213,N_17477);
and U21501 (N_21501,N_16321,N_17841);
and U21502 (N_21502,N_15818,N_17710);
xor U21503 (N_21503,N_16453,N_17073);
xnor U21504 (N_21504,N_17450,N_15844);
or U21505 (N_21505,N_15915,N_16586);
or U21506 (N_21506,N_18494,N_18571);
xor U21507 (N_21507,N_17209,N_15786);
nand U21508 (N_21508,N_17474,N_18624);
nor U21509 (N_21509,N_17978,N_15684);
nor U21510 (N_21510,N_18145,N_17767);
or U21511 (N_21511,N_17524,N_18138);
nand U21512 (N_21512,N_18221,N_18226);
and U21513 (N_21513,N_18096,N_17569);
or U21514 (N_21514,N_18402,N_17233);
nor U21515 (N_21515,N_15629,N_15739);
or U21516 (N_21516,N_17501,N_18411);
xor U21517 (N_21517,N_17105,N_16090);
nand U21518 (N_21518,N_18673,N_18579);
nand U21519 (N_21519,N_18440,N_17839);
and U21520 (N_21520,N_18042,N_15991);
nor U21521 (N_21521,N_17829,N_17925);
nor U21522 (N_21522,N_17447,N_16778);
and U21523 (N_21523,N_16189,N_17970);
or U21524 (N_21524,N_16148,N_15912);
or U21525 (N_21525,N_16747,N_15679);
nor U21526 (N_21526,N_15698,N_16079);
and U21527 (N_21527,N_18166,N_15975);
xor U21528 (N_21528,N_16267,N_17836);
and U21529 (N_21529,N_17463,N_15694);
xnor U21530 (N_21530,N_17854,N_16801);
nand U21531 (N_21531,N_18410,N_16825);
or U21532 (N_21532,N_17683,N_17867);
nor U21533 (N_21533,N_16898,N_16340);
and U21534 (N_21534,N_16929,N_16485);
nand U21535 (N_21535,N_16319,N_16697);
or U21536 (N_21536,N_16942,N_17112);
xnor U21537 (N_21537,N_17167,N_17887);
and U21538 (N_21538,N_17270,N_16884);
xor U21539 (N_21539,N_16109,N_16887);
or U21540 (N_21540,N_17747,N_17015);
and U21541 (N_21541,N_15878,N_18529);
xnor U21542 (N_21542,N_17300,N_17057);
nand U21543 (N_21543,N_16269,N_16104);
nand U21544 (N_21544,N_16563,N_17313);
and U21545 (N_21545,N_16440,N_15774);
nor U21546 (N_21546,N_16014,N_17411);
nor U21547 (N_21547,N_17661,N_17915);
nand U21548 (N_21548,N_15854,N_15772);
or U21549 (N_21549,N_15874,N_16183);
nor U21550 (N_21550,N_17490,N_16882);
or U21551 (N_21551,N_16898,N_16595);
nand U21552 (N_21552,N_16896,N_17436);
nor U21553 (N_21553,N_15714,N_17451);
and U21554 (N_21554,N_16267,N_17803);
nand U21555 (N_21555,N_16641,N_18613);
nand U21556 (N_21556,N_15847,N_18616);
and U21557 (N_21557,N_16763,N_16875);
nand U21558 (N_21558,N_16448,N_17287);
and U21559 (N_21559,N_16151,N_15916);
and U21560 (N_21560,N_18581,N_16016);
and U21561 (N_21561,N_16901,N_15711);
nand U21562 (N_21562,N_16234,N_16775);
or U21563 (N_21563,N_17313,N_18569);
xor U21564 (N_21564,N_16231,N_18222);
and U21565 (N_21565,N_16581,N_16266);
nor U21566 (N_21566,N_18476,N_15929);
and U21567 (N_21567,N_17549,N_16323);
and U21568 (N_21568,N_15903,N_17394);
nand U21569 (N_21569,N_16128,N_18486);
nand U21570 (N_21570,N_16570,N_18365);
nor U21571 (N_21571,N_18265,N_18539);
nand U21572 (N_21572,N_15745,N_17777);
nor U21573 (N_21573,N_16458,N_18427);
and U21574 (N_21574,N_18215,N_16205);
nand U21575 (N_21575,N_16481,N_18416);
nor U21576 (N_21576,N_16633,N_16084);
nor U21577 (N_21577,N_16283,N_15943);
nand U21578 (N_21578,N_17702,N_15794);
and U21579 (N_21579,N_16321,N_18338);
xnor U21580 (N_21580,N_17550,N_17239);
nand U21581 (N_21581,N_17353,N_18694);
nand U21582 (N_21582,N_18374,N_16370);
or U21583 (N_21583,N_18147,N_17759);
or U21584 (N_21584,N_17647,N_16680);
nor U21585 (N_21585,N_17451,N_18437);
or U21586 (N_21586,N_18435,N_17823);
xnor U21587 (N_21587,N_17425,N_17506);
or U21588 (N_21588,N_17128,N_18499);
or U21589 (N_21589,N_18608,N_17952);
and U21590 (N_21590,N_18379,N_16288);
and U21591 (N_21591,N_17586,N_17173);
nand U21592 (N_21592,N_15919,N_15897);
or U21593 (N_21593,N_15647,N_18492);
or U21594 (N_21594,N_18141,N_18744);
nand U21595 (N_21595,N_16037,N_17283);
xnor U21596 (N_21596,N_16972,N_17737);
nand U21597 (N_21597,N_15868,N_18519);
nor U21598 (N_21598,N_16797,N_16947);
nor U21599 (N_21599,N_18519,N_16080);
nor U21600 (N_21600,N_18305,N_18723);
nand U21601 (N_21601,N_16863,N_15740);
nor U21602 (N_21602,N_16976,N_17418);
and U21603 (N_21603,N_17435,N_17397);
nand U21604 (N_21604,N_18246,N_17081);
and U21605 (N_21605,N_17882,N_17074);
xnor U21606 (N_21606,N_16460,N_17485);
nor U21607 (N_21607,N_18388,N_18126);
and U21608 (N_21608,N_16113,N_16798);
and U21609 (N_21609,N_17657,N_17649);
nand U21610 (N_21610,N_18512,N_16146);
nor U21611 (N_21611,N_17348,N_18266);
nor U21612 (N_21612,N_17996,N_15950);
or U21613 (N_21613,N_15813,N_18159);
nor U21614 (N_21614,N_18083,N_16358);
or U21615 (N_21615,N_16839,N_15727);
or U21616 (N_21616,N_18510,N_15805);
nor U21617 (N_21617,N_18514,N_17771);
and U21618 (N_21618,N_16459,N_16943);
xnor U21619 (N_21619,N_16673,N_17606);
or U21620 (N_21620,N_16601,N_16122);
or U21621 (N_21621,N_17871,N_15731);
nand U21622 (N_21622,N_16904,N_16508);
or U21623 (N_21623,N_16178,N_16260);
nand U21624 (N_21624,N_18159,N_16096);
or U21625 (N_21625,N_16136,N_18606);
nor U21626 (N_21626,N_18466,N_18461);
xnor U21627 (N_21627,N_18409,N_17218);
nand U21628 (N_21628,N_17280,N_16936);
xor U21629 (N_21629,N_15681,N_18661);
xor U21630 (N_21630,N_16318,N_17961);
nand U21631 (N_21631,N_18175,N_18675);
xor U21632 (N_21632,N_17839,N_16882);
and U21633 (N_21633,N_16152,N_17457);
or U21634 (N_21634,N_18066,N_16156);
xor U21635 (N_21635,N_18612,N_16074);
or U21636 (N_21636,N_17829,N_16225);
or U21637 (N_21637,N_17563,N_18419);
xor U21638 (N_21638,N_16088,N_18381);
and U21639 (N_21639,N_18339,N_18607);
and U21640 (N_21640,N_18293,N_18372);
and U21641 (N_21641,N_17962,N_18457);
xor U21642 (N_21642,N_18737,N_16273);
xor U21643 (N_21643,N_18487,N_17195);
and U21644 (N_21644,N_15802,N_17916);
nor U21645 (N_21645,N_16922,N_18057);
or U21646 (N_21646,N_17216,N_17697);
or U21647 (N_21647,N_17865,N_16651);
and U21648 (N_21648,N_16196,N_15956);
nor U21649 (N_21649,N_16025,N_17048);
nand U21650 (N_21650,N_16261,N_18620);
and U21651 (N_21651,N_16426,N_15806);
xnor U21652 (N_21652,N_16338,N_16965);
nor U21653 (N_21653,N_16664,N_17875);
nand U21654 (N_21654,N_18657,N_18185);
and U21655 (N_21655,N_17393,N_18139);
or U21656 (N_21656,N_16007,N_17196);
nand U21657 (N_21657,N_17733,N_17257);
or U21658 (N_21658,N_16170,N_18337);
nor U21659 (N_21659,N_16175,N_17942);
and U21660 (N_21660,N_15743,N_18282);
nor U21661 (N_21661,N_16844,N_17602);
or U21662 (N_21662,N_16734,N_17105);
and U21663 (N_21663,N_17284,N_18191);
nand U21664 (N_21664,N_17449,N_16719);
and U21665 (N_21665,N_16014,N_17442);
or U21666 (N_21666,N_17821,N_16348);
nor U21667 (N_21667,N_16462,N_16904);
nand U21668 (N_21668,N_15849,N_17325);
or U21669 (N_21669,N_18694,N_17662);
or U21670 (N_21670,N_16743,N_16694);
nand U21671 (N_21671,N_18525,N_17682);
nand U21672 (N_21672,N_17553,N_18314);
and U21673 (N_21673,N_17877,N_16025);
nor U21674 (N_21674,N_17516,N_15671);
nand U21675 (N_21675,N_15879,N_16552);
xor U21676 (N_21676,N_17713,N_16611);
xnor U21677 (N_21677,N_17308,N_18660);
nand U21678 (N_21678,N_17764,N_16948);
nor U21679 (N_21679,N_16949,N_17156);
or U21680 (N_21680,N_16938,N_17989);
and U21681 (N_21681,N_18154,N_15935);
nor U21682 (N_21682,N_17532,N_17417);
nor U21683 (N_21683,N_17777,N_16993);
xor U21684 (N_21684,N_16637,N_17517);
nand U21685 (N_21685,N_17287,N_16469);
or U21686 (N_21686,N_17385,N_16121);
or U21687 (N_21687,N_17311,N_16909);
and U21688 (N_21688,N_18585,N_16634);
nor U21689 (N_21689,N_18118,N_17112);
and U21690 (N_21690,N_16297,N_16444);
and U21691 (N_21691,N_17763,N_16938);
nor U21692 (N_21692,N_16012,N_16947);
or U21693 (N_21693,N_18617,N_16313);
or U21694 (N_21694,N_15956,N_16021);
and U21695 (N_21695,N_17159,N_18417);
and U21696 (N_21696,N_16344,N_17545);
nor U21697 (N_21697,N_16342,N_16034);
nand U21698 (N_21698,N_16192,N_15998);
or U21699 (N_21699,N_16031,N_16546);
or U21700 (N_21700,N_17615,N_18111);
and U21701 (N_21701,N_16203,N_17073);
nand U21702 (N_21702,N_15827,N_16353);
and U21703 (N_21703,N_18155,N_17111);
nand U21704 (N_21704,N_17169,N_17708);
nand U21705 (N_21705,N_16673,N_18729);
or U21706 (N_21706,N_16318,N_15667);
and U21707 (N_21707,N_17110,N_16967);
and U21708 (N_21708,N_15884,N_16192);
or U21709 (N_21709,N_15650,N_16754);
nand U21710 (N_21710,N_15683,N_18011);
nor U21711 (N_21711,N_16288,N_18390);
nor U21712 (N_21712,N_18253,N_16659);
or U21713 (N_21713,N_16026,N_17284);
nand U21714 (N_21714,N_17822,N_16321);
and U21715 (N_21715,N_18459,N_16272);
nand U21716 (N_21716,N_17803,N_17654);
nand U21717 (N_21717,N_17046,N_16520);
or U21718 (N_21718,N_17423,N_15798);
nand U21719 (N_21719,N_17524,N_15740);
or U21720 (N_21720,N_17950,N_15640);
nor U21721 (N_21721,N_16150,N_18361);
nand U21722 (N_21722,N_18263,N_16100);
nor U21723 (N_21723,N_17277,N_16550);
nand U21724 (N_21724,N_17119,N_17915);
nand U21725 (N_21725,N_16088,N_18565);
xnor U21726 (N_21726,N_17335,N_15662);
and U21727 (N_21727,N_16941,N_17856);
nand U21728 (N_21728,N_16916,N_17257);
nor U21729 (N_21729,N_16050,N_18335);
and U21730 (N_21730,N_16736,N_16671);
xor U21731 (N_21731,N_18204,N_16396);
nand U21732 (N_21732,N_16089,N_16285);
or U21733 (N_21733,N_17263,N_16406);
nand U21734 (N_21734,N_17396,N_15990);
or U21735 (N_21735,N_17741,N_17193);
nor U21736 (N_21736,N_17363,N_18072);
nor U21737 (N_21737,N_17139,N_17755);
xor U21738 (N_21738,N_18492,N_16733);
nor U21739 (N_21739,N_17761,N_17660);
or U21740 (N_21740,N_15962,N_15832);
nand U21741 (N_21741,N_18552,N_15852);
or U21742 (N_21742,N_17792,N_15779);
nor U21743 (N_21743,N_17845,N_16935);
nand U21744 (N_21744,N_16421,N_16016);
nor U21745 (N_21745,N_17063,N_17054);
and U21746 (N_21746,N_16642,N_18437);
and U21747 (N_21747,N_18616,N_18534);
or U21748 (N_21748,N_18739,N_18524);
nand U21749 (N_21749,N_16233,N_17582);
xor U21750 (N_21750,N_16200,N_16907);
nor U21751 (N_21751,N_17140,N_18400);
nor U21752 (N_21752,N_17990,N_17790);
or U21753 (N_21753,N_15857,N_16327);
and U21754 (N_21754,N_17871,N_17901);
or U21755 (N_21755,N_15979,N_18112);
and U21756 (N_21756,N_18111,N_17276);
nor U21757 (N_21757,N_17674,N_17319);
nor U21758 (N_21758,N_17809,N_15764);
or U21759 (N_21759,N_18026,N_16439);
and U21760 (N_21760,N_17688,N_18008);
and U21761 (N_21761,N_16373,N_16072);
nand U21762 (N_21762,N_18278,N_15821);
nor U21763 (N_21763,N_16987,N_16310);
nand U21764 (N_21764,N_18176,N_18395);
nand U21765 (N_21765,N_16833,N_17749);
nand U21766 (N_21766,N_17423,N_18031);
or U21767 (N_21767,N_17358,N_17910);
or U21768 (N_21768,N_15955,N_16210);
nor U21769 (N_21769,N_18423,N_15722);
nor U21770 (N_21770,N_16098,N_18240);
nand U21771 (N_21771,N_16784,N_17683);
xnor U21772 (N_21772,N_17350,N_16687);
or U21773 (N_21773,N_18608,N_16308);
or U21774 (N_21774,N_18408,N_16308);
or U21775 (N_21775,N_17659,N_17902);
or U21776 (N_21776,N_17685,N_18280);
or U21777 (N_21777,N_16735,N_16185);
and U21778 (N_21778,N_18162,N_16833);
or U21779 (N_21779,N_17104,N_17182);
or U21780 (N_21780,N_15863,N_17631);
xor U21781 (N_21781,N_17825,N_17331);
or U21782 (N_21782,N_17131,N_15842);
nand U21783 (N_21783,N_18224,N_18091);
nand U21784 (N_21784,N_16637,N_16792);
or U21785 (N_21785,N_18356,N_15938);
nor U21786 (N_21786,N_16584,N_18662);
nand U21787 (N_21787,N_16899,N_18057);
nor U21788 (N_21788,N_18259,N_18502);
nor U21789 (N_21789,N_17130,N_17295);
nor U21790 (N_21790,N_17175,N_15671);
or U21791 (N_21791,N_16298,N_16932);
or U21792 (N_21792,N_16821,N_16345);
or U21793 (N_21793,N_17507,N_17140);
nand U21794 (N_21794,N_16711,N_16918);
and U21795 (N_21795,N_18703,N_17490);
and U21796 (N_21796,N_18222,N_18485);
xor U21797 (N_21797,N_15688,N_18104);
and U21798 (N_21798,N_18402,N_16623);
nand U21799 (N_21799,N_18742,N_17206);
or U21800 (N_21800,N_17653,N_16385);
nor U21801 (N_21801,N_15977,N_18017);
and U21802 (N_21802,N_17881,N_17643);
and U21803 (N_21803,N_17752,N_17787);
nor U21804 (N_21804,N_15884,N_17856);
nand U21805 (N_21805,N_18614,N_16488);
and U21806 (N_21806,N_18448,N_16131);
or U21807 (N_21807,N_18454,N_16991);
and U21808 (N_21808,N_17114,N_17931);
xnor U21809 (N_21809,N_18647,N_15737);
nand U21810 (N_21810,N_15806,N_17120);
nor U21811 (N_21811,N_18352,N_17286);
nor U21812 (N_21812,N_18684,N_16795);
and U21813 (N_21813,N_15967,N_17084);
nand U21814 (N_21814,N_17114,N_16685);
or U21815 (N_21815,N_16866,N_17293);
or U21816 (N_21816,N_17625,N_18580);
nand U21817 (N_21817,N_16072,N_16202);
xnor U21818 (N_21818,N_15731,N_16392);
or U21819 (N_21819,N_17731,N_16906);
and U21820 (N_21820,N_16325,N_16160);
nand U21821 (N_21821,N_17289,N_15881);
nand U21822 (N_21822,N_15927,N_16349);
and U21823 (N_21823,N_17217,N_17456);
nand U21824 (N_21824,N_18546,N_18713);
and U21825 (N_21825,N_18552,N_17757);
nand U21826 (N_21826,N_17007,N_16040);
nand U21827 (N_21827,N_17732,N_15876);
or U21828 (N_21828,N_15654,N_18430);
or U21829 (N_21829,N_17652,N_18300);
and U21830 (N_21830,N_17161,N_16778);
and U21831 (N_21831,N_15847,N_16165);
nor U21832 (N_21832,N_18009,N_17438);
or U21833 (N_21833,N_16149,N_18379);
or U21834 (N_21834,N_16882,N_17009);
nor U21835 (N_21835,N_18370,N_17323);
nor U21836 (N_21836,N_16920,N_18016);
nor U21837 (N_21837,N_17329,N_18740);
nor U21838 (N_21838,N_16022,N_17839);
or U21839 (N_21839,N_16280,N_16574);
nand U21840 (N_21840,N_17905,N_16099);
nor U21841 (N_21841,N_16955,N_16297);
nand U21842 (N_21842,N_16016,N_18717);
or U21843 (N_21843,N_16641,N_15736);
nor U21844 (N_21844,N_16321,N_15639);
nor U21845 (N_21845,N_18402,N_18232);
nand U21846 (N_21846,N_17937,N_16046);
and U21847 (N_21847,N_15706,N_17574);
and U21848 (N_21848,N_17872,N_18739);
and U21849 (N_21849,N_16604,N_16943);
or U21850 (N_21850,N_17881,N_18003);
xnor U21851 (N_21851,N_16080,N_16041);
nor U21852 (N_21852,N_16535,N_17200);
nor U21853 (N_21853,N_16810,N_16181);
or U21854 (N_21854,N_16904,N_17758);
and U21855 (N_21855,N_17937,N_16307);
nand U21856 (N_21856,N_15688,N_16965);
nor U21857 (N_21857,N_16043,N_18595);
nor U21858 (N_21858,N_18431,N_16640);
nand U21859 (N_21859,N_16632,N_16726);
and U21860 (N_21860,N_16828,N_17281);
nor U21861 (N_21861,N_17635,N_17472);
nor U21862 (N_21862,N_16346,N_16290);
and U21863 (N_21863,N_15856,N_17996);
and U21864 (N_21864,N_16663,N_15853);
nand U21865 (N_21865,N_16597,N_16364);
and U21866 (N_21866,N_17692,N_16316);
nor U21867 (N_21867,N_18283,N_18489);
xor U21868 (N_21868,N_16597,N_18590);
nand U21869 (N_21869,N_17140,N_17214);
or U21870 (N_21870,N_16265,N_17862);
nor U21871 (N_21871,N_17435,N_18675);
and U21872 (N_21872,N_17682,N_15730);
and U21873 (N_21873,N_17443,N_17233);
and U21874 (N_21874,N_15935,N_18673);
nand U21875 (N_21875,N_20218,N_19430);
nand U21876 (N_21876,N_19780,N_21055);
nor U21877 (N_21877,N_21485,N_21279);
and U21878 (N_21878,N_19192,N_19653);
nor U21879 (N_21879,N_19909,N_20100);
nor U21880 (N_21880,N_20280,N_20820);
nor U21881 (N_21881,N_21084,N_18882);
nor U21882 (N_21882,N_21200,N_20053);
xor U21883 (N_21883,N_20604,N_19468);
nand U21884 (N_21884,N_21840,N_19530);
and U21885 (N_21885,N_20360,N_20346);
and U21886 (N_21886,N_20096,N_20467);
or U21887 (N_21887,N_20716,N_20476);
or U21888 (N_21888,N_21805,N_20259);
and U21889 (N_21889,N_20037,N_19835);
or U21890 (N_21890,N_21305,N_19828);
and U21891 (N_21891,N_19873,N_19386);
nand U21892 (N_21892,N_19338,N_19638);
nand U21893 (N_21893,N_18814,N_20244);
xnor U21894 (N_21894,N_19552,N_18995);
xor U21895 (N_21895,N_20021,N_18853);
and U21896 (N_21896,N_20181,N_21429);
nor U21897 (N_21897,N_19993,N_21071);
nand U21898 (N_21898,N_21235,N_20433);
and U21899 (N_21899,N_19082,N_21268);
and U21900 (N_21900,N_21580,N_20395);
and U21901 (N_21901,N_19499,N_18850);
and U21902 (N_21902,N_19469,N_21536);
nand U21903 (N_21903,N_19436,N_19704);
or U21904 (N_21904,N_21064,N_18799);
and U21905 (N_21905,N_20928,N_18880);
or U21906 (N_21906,N_20863,N_19396);
and U21907 (N_21907,N_20664,N_20800);
xnor U21908 (N_21908,N_19830,N_21099);
and U21909 (N_21909,N_21865,N_20355);
or U21910 (N_21910,N_20042,N_21868);
nor U21911 (N_21911,N_18779,N_19786);
nand U21912 (N_21912,N_19603,N_20164);
nor U21913 (N_21913,N_20076,N_19076);
xor U21914 (N_21914,N_21339,N_19551);
xnor U21915 (N_21915,N_19990,N_20421);
and U21916 (N_21916,N_20298,N_20271);
nand U21917 (N_21917,N_19750,N_19762);
or U21918 (N_21918,N_20990,N_21301);
nor U21919 (N_21919,N_18849,N_19269);
nor U21920 (N_21920,N_19311,N_20032);
and U21921 (N_21921,N_19688,N_20058);
nor U21922 (N_21922,N_20529,N_21665);
or U21923 (N_21923,N_21440,N_19196);
nor U21924 (N_21924,N_20815,N_21802);
nor U21925 (N_21925,N_20892,N_18948);
nor U21926 (N_21926,N_21004,N_20835);
and U21927 (N_21927,N_20370,N_20029);
and U21928 (N_21928,N_18824,N_19191);
and U21929 (N_21929,N_20180,N_20153);
nand U21930 (N_21930,N_18816,N_20419);
nand U21931 (N_21931,N_19014,N_19033);
and U21932 (N_21932,N_20002,N_19091);
nand U21933 (N_21933,N_20673,N_21834);
nor U21934 (N_21934,N_21025,N_19781);
and U21935 (N_21935,N_21843,N_20507);
and U21936 (N_21936,N_20920,N_21214);
and U21937 (N_21937,N_18841,N_19732);
nand U21938 (N_21938,N_21428,N_19952);
or U21939 (N_21939,N_20817,N_21558);
xor U21940 (N_21940,N_21596,N_21330);
or U21941 (N_21941,N_20812,N_21056);
and U21942 (N_21942,N_18900,N_21647);
nor U21943 (N_21943,N_20225,N_21143);
nand U21944 (N_21944,N_21780,N_18913);
or U21945 (N_21945,N_20022,N_20099);
and U21946 (N_21946,N_19544,N_21572);
or U21947 (N_21947,N_18840,N_21737);
or U21948 (N_21948,N_20547,N_21541);
or U21949 (N_21949,N_21273,N_20450);
nor U21950 (N_21950,N_21545,N_19339);
nand U21951 (N_21951,N_19838,N_19372);
nor U21952 (N_21952,N_19517,N_21808);
or U21953 (N_21953,N_21848,N_20951);
xor U21954 (N_21954,N_21569,N_19641);
or U21955 (N_21955,N_21197,N_19047);
nand U21956 (N_21956,N_19111,N_20803);
and U21957 (N_21957,N_19337,N_19153);
or U21958 (N_21958,N_20160,N_19418);
nand U21959 (N_21959,N_19102,N_20456);
nor U21960 (N_21960,N_18886,N_21019);
xnor U21961 (N_21961,N_21123,N_19371);
nor U21962 (N_21962,N_21542,N_20434);
nand U21963 (N_21963,N_20030,N_20762);
nor U21964 (N_21964,N_21576,N_19237);
or U21965 (N_21965,N_20212,N_19158);
and U21966 (N_21966,N_21109,N_19996);
nor U21967 (N_21967,N_20177,N_21151);
or U21968 (N_21968,N_19836,N_20430);
nand U21969 (N_21969,N_19813,N_21613);
nand U21970 (N_21970,N_20861,N_21491);
or U21971 (N_21971,N_19722,N_19821);
or U21972 (N_21972,N_18844,N_21163);
or U21973 (N_21973,N_19204,N_20124);
or U21974 (N_21974,N_19861,N_20324);
nor U21975 (N_21975,N_21207,N_20125);
xor U21976 (N_21976,N_19009,N_19325);
and U21977 (N_21977,N_19506,N_21815);
or U21978 (N_21978,N_19380,N_20031);
and U21979 (N_21979,N_20926,N_20921);
nor U21980 (N_21980,N_19934,N_19353);
nor U21981 (N_21981,N_20953,N_20734);
and U21982 (N_21982,N_19531,N_19706);
nor U21983 (N_21983,N_21680,N_21872);
or U21984 (N_21984,N_19957,N_21586);
and U21985 (N_21985,N_21540,N_20832);
nand U21986 (N_21986,N_21487,N_20714);
and U21987 (N_21987,N_19774,N_21756);
or U21988 (N_21988,N_20742,N_19299);
or U21989 (N_21989,N_19730,N_20767);
nor U21990 (N_21990,N_20189,N_20655);
nand U21991 (N_21991,N_18883,N_21316);
nand U21992 (N_21992,N_20389,N_19363);
or U21993 (N_21993,N_21749,N_21068);
and U21994 (N_21994,N_19583,N_20797);
nor U21995 (N_21995,N_20003,N_19385);
nand U21996 (N_21996,N_20750,N_19019);
nand U21997 (N_21997,N_19526,N_21841);
or U21998 (N_21998,N_19570,N_19634);
nor U21999 (N_21999,N_18968,N_21451);
nand U22000 (N_22000,N_19218,N_20846);
nand U22001 (N_22001,N_20935,N_19301);
nand U22002 (N_22002,N_20975,N_20545);
and U22003 (N_22003,N_21827,N_21721);
nor U22004 (N_22004,N_18997,N_19733);
nand U22005 (N_22005,N_20348,N_20005);
nand U22006 (N_22006,N_20410,N_18927);
nand U22007 (N_22007,N_21061,N_20985);
nand U22008 (N_22008,N_21522,N_19001);
or U22009 (N_22009,N_19248,N_18996);
and U22010 (N_22010,N_19516,N_20241);
and U22011 (N_22011,N_20878,N_20642);
or U22012 (N_22012,N_19484,N_20060);
nor U22013 (N_22013,N_20741,N_19403);
nor U22014 (N_22014,N_19746,N_19520);
or U22015 (N_22015,N_20633,N_19441);
or U22016 (N_22016,N_21725,N_19253);
or U22017 (N_22017,N_20701,N_19765);
or U22018 (N_22018,N_21332,N_19627);
and U22019 (N_22019,N_21103,N_19394);
nor U22020 (N_22020,N_19171,N_21619);
nor U22021 (N_22021,N_18767,N_19295);
nor U22022 (N_22022,N_20033,N_21139);
nor U22023 (N_22023,N_21436,N_21464);
or U22024 (N_22024,N_20302,N_21626);
nand U22025 (N_22025,N_19362,N_21248);
or U22026 (N_22026,N_20868,N_21810);
and U22027 (N_22027,N_20710,N_21473);
and U22028 (N_22028,N_21229,N_19005);
and U22029 (N_22029,N_20167,N_21191);
and U22030 (N_22030,N_19984,N_21469);
nor U22031 (N_22031,N_19265,N_18879);
xor U22032 (N_22032,N_20810,N_20535);
nand U22033 (N_22033,N_20713,N_19720);
xor U22034 (N_22034,N_20080,N_21657);
xor U22035 (N_22035,N_20974,N_20605);
nand U22036 (N_22036,N_19814,N_21635);
or U22037 (N_22037,N_18932,N_19951);
or U22038 (N_22038,N_20704,N_20027);
nor U22039 (N_22039,N_20161,N_19271);
and U22040 (N_22040,N_19025,N_21551);
nand U22041 (N_22041,N_19919,N_20579);
or U22042 (N_22042,N_21298,N_20196);
nor U22043 (N_22043,N_19837,N_20310);
or U22044 (N_22044,N_21049,N_20245);
or U22045 (N_22045,N_18805,N_19854);
nor U22046 (N_22046,N_21477,N_20035);
and U22047 (N_22047,N_20598,N_19041);
and U22048 (N_22048,N_19642,N_21465);
nor U22049 (N_22049,N_19756,N_21766);
or U22050 (N_22050,N_19564,N_19938);
and U22051 (N_22051,N_20268,N_20536);
nor U22052 (N_22052,N_21475,N_20538);
or U22053 (N_22053,N_21864,N_19616);
nor U22054 (N_22054,N_20504,N_20544);
and U22055 (N_22055,N_20007,N_19841);
or U22056 (N_22056,N_20093,N_20277);
nand U22057 (N_22057,N_20864,N_20250);
nand U22058 (N_22058,N_20045,N_20192);
xnor U22059 (N_22059,N_19929,N_21026);
nand U22060 (N_22060,N_20632,N_21342);
and U22061 (N_22061,N_18830,N_21304);
nor U22062 (N_22062,N_21589,N_20749);
and U22063 (N_22063,N_21320,N_18867);
nand U22064 (N_22064,N_18977,N_20776);
xor U22065 (N_22065,N_19416,N_19630);
nor U22066 (N_22066,N_18862,N_20191);
and U22067 (N_22067,N_20667,N_18833);
nor U22068 (N_22068,N_19581,N_20429);
nand U22069 (N_22069,N_21459,N_21696);
nand U22070 (N_22070,N_21242,N_18916);
nor U22071 (N_22071,N_19450,N_19163);
or U22072 (N_22072,N_21801,N_19715);
nor U22073 (N_22073,N_21387,N_20765);
nor U22074 (N_22074,N_18922,N_20374);
nand U22075 (N_22075,N_19661,N_19840);
nand U22076 (N_22076,N_21524,N_21760);
and U22077 (N_22077,N_18838,N_20373);
nand U22078 (N_22078,N_21390,N_18768);
nand U22079 (N_22079,N_20318,N_19423);
nor U22080 (N_22080,N_20929,N_18896);
nand U22081 (N_22081,N_19930,N_21411);
nor U22082 (N_22082,N_18852,N_20681);
or U22083 (N_22083,N_21720,N_18764);
and U22084 (N_22084,N_21328,N_19702);
and U22085 (N_22085,N_21627,N_19698);
nor U22086 (N_22086,N_19580,N_21643);
xor U22087 (N_22087,N_20722,N_21188);
nand U22088 (N_22088,N_21137,N_21272);
and U22089 (N_22089,N_20871,N_19947);
and U22090 (N_22090,N_21554,N_19536);
nand U22091 (N_22091,N_20262,N_21670);
or U22092 (N_22092,N_19096,N_19390);
nor U22093 (N_22093,N_21098,N_18935);
nand U22094 (N_22094,N_19816,N_19547);
xor U22095 (N_22095,N_20018,N_20548);
and U22096 (N_22096,N_19176,N_21434);
or U22097 (N_22097,N_19135,N_18750);
nand U22098 (N_22098,N_20630,N_20121);
xor U22099 (N_22099,N_21507,N_18857);
or U22100 (N_22100,N_21419,N_21870);
or U22101 (N_22101,N_19791,N_20565);
nor U22102 (N_22102,N_21127,N_20013);
and U22103 (N_22103,N_21383,N_21422);
and U22104 (N_22104,N_18837,N_19618);
and U22105 (N_22105,N_19454,N_21605);
and U22106 (N_22106,N_19666,N_21562);
nor U22107 (N_22107,N_19721,N_19637);
or U22108 (N_22108,N_19562,N_20702);
nor U22109 (N_22109,N_20391,N_19682);
and U22110 (N_22110,N_19649,N_19480);
nand U22111 (N_22111,N_21511,N_20933);
and U22112 (N_22112,N_20014,N_21822);
nor U22113 (N_22113,N_20672,N_20345);
and U22114 (N_22114,N_20983,N_21578);
nor U22115 (N_22115,N_18917,N_20133);
nor U22116 (N_22116,N_21832,N_20226);
or U22117 (N_22117,N_19458,N_20534);
nor U22118 (N_22118,N_20119,N_21282);
nor U22119 (N_22119,N_21276,N_18826);
and U22120 (N_22120,N_21639,N_20743);
xor U22121 (N_22121,N_19757,N_19407);
and U22122 (N_22122,N_20554,N_21168);
xor U22123 (N_22123,N_20221,N_19056);
nand U22124 (N_22124,N_21468,N_20500);
nor U22125 (N_22125,N_19261,N_19515);
or U22126 (N_22126,N_21615,N_19665);
nand U22127 (N_22127,N_20201,N_20441);
or U22128 (N_22128,N_20889,N_19745);
or U22129 (N_22129,N_19400,N_19148);
and U22130 (N_22130,N_21510,N_21287);
or U22131 (N_22131,N_19933,N_18806);
or U22132 (N_22132,N_20350,N_20256);
xnor U22133 (N_22133,N_20165,N_19632);
nor U22134 (N_22134,N_19592,N_19556);
or U22135 (N_22135,N_19635,N_20130);
nor U22136 (N_22136,N_20830,N_20838);
nor U22137 (N_22137,N_21764,N_19509);
or U22138 (N_22138,N_21245,N_19811);
and U22139 (N_22139,N_18789,N_19227);
or U22140 (N_22140,N_20780,N_18982);
and U22141 (N_22141,N_19471,N_21755);
or U22142 (N_22142,N_18998,N_21817);
or U22143 (N_22143,N_20621,N_21021);
and U22144 (N_22144,N_19655,N_19086);
xor U22145 (N_22145,N_18920,N_20590);
nor U22146 (N_22146,N_20764,N_20782);
nor U22147 (N_22147,N_19845,N_21426);
nor U22148 (N_22148,N_20291,N_21231);
nand U22149 (N_22149,N_20850,N_19029);
nand U22150 (N_22150,N_21753,N_21223);
and U22151 (N_22151,N_21553,N_20103);
and U22152 (N_22152,N_18868,N_19879);
xor U22153 (N_22153,N_20073,N_20980);
and U22154 (N_22154,N_20730,N_21311);
nor U22155 (N_22155,N_19870,N_19998);
nor U22156 (N_22156,N_19586,N_20752);
or U22157 (N_22157,N_21280,N_20139);
xnor U22158 (N_22158,N_20786,N_19350);
or U22159 (N_22159,N_18786,N_19659);
nand U22160 (N_22160,N_21326,N_20445);
nor U22161 (N_22161,N_20969,N_20608);
and U22162 (N_22162,N_18780,N_19856);
or U22163 (N_22163,N_21660,N_20383);
nand U22164 (N_22164,N_19654,N_21263);
or U22165 (N_22165,N_20745,N_20267);
nor U22166 (N_22166,N_20332,N_20942);
or U22167 (N_22167,N_18999,N_19678);
and U22168 (N_22168,N_19032,N_21396);
nand U22169 (N_22169,N_21042,N_21687);
nor U22170 (N_22170,N_19815,N_21839);
or U22171 (N_22171,N_20772,N_20727);
and U22172 (N_22172,N_21382,N_19123);
or U22173 (N_22173,N_21686,N_21862);
or U22174 (N_22174,N_20187,N_20106);
nand U22175 (N_22175,N_21782,N_21495);
or U22176 (N_22176,N_21120,N_20530);
and U22177 (N_22177,N_19226,N_19905);
or U22178 (N_22178,N_21166,N_20769);
nand U22179 (N_22179,N_20138,N_20305);
or U22180 (N_22180,N_18847,N_20062);
and U22181 (N_22181,N_19554,N_20089);
nand U22182 (N_22182,N_20307,N_19315);
nand U22183 (N_22183,N_21857,N_21077);
nor U22184 (N_22184,N_21117,N_19972);
or U22185 (N_22185,N_21238,N_18865);
or U22186 (N_22186,N_19072,N_18760);
or U22187 (N_22187,N_20426,N_20930);
and U22188 (N_22188,N_21852,N_19297);
nor U22189 (N_22189,N_19366,N_19281);
nor U22190 (N_22190,N_19831,N_20174);
nor U22191 (N_22191,N_19557,N_20872);
or U22192 (N_22192,N_20614,N_20394);
nor U22193 (N_22193,N_19048,N_21296);
nand U22194 (N_22194,N_20276,N_18877);
nor U22195 (N_22195,N_21446,N_20993);
nor U22196 (N_22196,N_19863,N_18926);
nand U22197 (N_22197,N_20179,N_21778);
and U22198 (N_22198,N_19069,N_21048);
or U22199 (N_22199,N_20477,N_19968);
nand U22200 (N_22200,N_21013,N_20966);
and U22201 (N_22201,N_21492,N_21552);
and U22202 (N_22202,N_20626,N_18859);
nor U22203 (N_22203,N_21407,N_20490);
nor U22204 (N_22204,N_21823,N_19270);
nand U22205 (N_22205,N_20322,N_19925);
and U22206 (N_22206,N_21192,N_18866);
nand U22207 (N_22207,N_19073,N_21813);
or U22208 (N_22208,N_20399,N_20246);
or U22209 (N_22209,N_21338,N_21178);
and U22210 (N_22210,N_21763,N_19883);
xnor U22211 (N_22211,N_20881,N_20746);
nor U22212 (N_22212,N_19614,N_19387);
nor U22213 (N_22213,N_20676,N_21362);
or U22214 (N_22214,N_20593,N_19264);
and U22215 (N_22215,N_19244,N_20697);
or U22216 (N_22216,N_18793,N_19277);
nor U22217 (N_22217,N_21222,N_18762);
xor U22218 (N_22218,N_21692,N_19116);
xnor U22219 (N_22219,N_20844,N_19426);
or U22220 (N_22220,N_20065,N_19617);
nor U22221 (N_22221,N_20773,N_19074);
and U22222 (N_22222,N_19956,N_20813);
xor U22223 (N_22223,N_19798,N_20634);
xor U22224 (N_22224,N_19120,N_19274);
and U22225 (N_22225,N_21591,N_20996);
nor U22226 (N_22226,N_19608,N_21063);
and U22227 (N_22227,N_21757,N_21788);
nor U22228 (N_22228,N_21190,N_19293);
nor U22229 (N_22229,N_20855,N_20357);
and U22230 (N_22230,N_20026,N_19252);
nand U22231 (N_22231,N_21136,N_21636);
or U22232 (N_22232,N_19448,N_18911);
or U22233 (N_22233,N_20973,N_19707);
or U22234 (N_22234,N_19010,N_21145);
or U22235 (N_22235,N_20950,N_18751);
nor U22236 (N_22236,N_19548,N_19037);
and U22237 (N_22237,N_21818,N_21275);
nand U22238 (N_22238,N_19291,N_19729);
or U22239 (N_22239,N_19119,N_19006);
xnor U22240 (N_22240,N_20690,N_20568);
nand U22241 (N_22241,N_19943,N_19523);
and U22242 (N_22242,N_18777,N_19725);
nor U22243 (N_22243,N_20049,N_20757);
nand U22244 (N_22244,N_21471,N_19190);
nand U22245 (N_22245,N_20827,N_21331);
and U22246 (N_22246,N_19173,N_20118);
nand U22247 (N_22247,N_19687,N_19950);
or U22248 (N_22248,N_19761,N_18803);
and U22249 (N_22249,N_19328,N_20193);
and U22250 (N_22250,N_19810,N_21097);
or U22251 (N_22251,N_20686,N_19693);
and U22252 (N_22252,N_20687,N_18819);
nor U22253 (N_22253,N_20852,N_19439);
nor U22254 (N_22254,N_21571,N_20890);
or U22255 (N_22255,N_18757,N_21566);
and U22256 (N_22256,N_19827,N_20249);
or U22257 (N_22257,N_19130,N_21079);
nor U22258 (N_22258,N_20081,N_18836);
xor U22259 (N_22259,N_20253,N_19125);
nand U22260 (N_22260,N_20078,N_20116);
nand U22261 (N_22261,N_20848,N_21360);
xnor U22262 (N_22262,N_21167,N_21230);
nor U22263 (N_22263,N_21257,N_20142);
and U22264 (N_22264,N_19206,N_19164);
or U22265 (N_22265,N_19594,N_21470);
nor U22266 (N_22266,N_19329,N_20279);
nand U22267 (N_22267,N_20329,N_20292);
nor U22268 (N_22268,N_19283,N_20822);
xnor U22269 (N_22269,N_20662,N_20651);
nand U22270 (N_22270,N_21286,N_21652);
or U22271 (N_22271,N_21095,N_20705);
or U22272 (N_22272,N_21825,N_21046);
or U22273 (N_22273,N_19059,N_21244);
nand U22274 (N_22274,N_19874,N_19429);
xnor U22275 (N_22275,N_21406,N_21836);
nor U22276 (N_22276,N_21258,N_19310);
nor U22277 (N_22277,N_19964,N_21460);
and U22278 (N_22278,N_20785,N_19485);
nand U22279 (N_22279,N_20923,N_21088);
nand U22280 (N_22280,N_20971,N_20495);
nand U22281 (N_22281,N_21154,N_21144);
nor U22282 (N_22282,N_21641,N_20023);
and U22283 (N_22283,N_20135,N_21124);
nor U22284 (N_22284,N_19267,N_19170);
and U22285 (N_22285,N_21774,N_20668);
xnor U22286 (N_22286,N_19289,N_20126);
xnor U22287 (N_22287,N_19042,N_21252);
nand U22288 (N_22288,N_18842,N_19185);
nand U22289 (N_22289,N_19657,N_20541);
and U22290 (N_22290,N_19121,N_19323);
nand U22291 (N_22291,N_19279,N_21685);
nand U22292 (N_22292,N_20558,N_20557);
xnor U22293 (N_22293,N_19210,N_20480);
or U22294 (N_22294,N_21441,N_21821);
nand U22295 (N_22295,N_20689,N_21353);
or U22296 (N_22296,N_21784,N_18787);
and U22297 (N_22297,N_20919,N_21447);
nand U22298 (N_22298,N_21072,N_20435);
and U22299 (N_22299,N_21726,N_18931);
or U22300 (N_22300,N_20208,N_19445);
xnor U22301 (N_22301,N_20281,N_20228);
nor U22302 (N_22302,N_19200,N_20523);
and U22303 (N_22303,N_19926,N_20371);
or U22304 (N_22304,N_19582,N_21773);
or U22305 (N_22305,N_20927,N_19446);
and U22306 (N_22306,N_19107,N_21804);
nand U22307 (N_22307,N_21744,N_21642);
and U22308 (N_22308,N_19705,N_19710);
nand U22309 (N_22309,N_18912,N_19359);
nand U22310 (N_22310,N_19075,N_20914);
nand U22311 (N_22311,N_20650,N_19979);
or U22312 (N_22312,N_18798,N_20674);
and U22313 (N_22313,N_19078,N_20064);
nand U22314 (N_22314,N_20723,N_19794);
nor U22315 (N_22315,N_20255,N_20638);
nand U22316 (N_22316,N_19629,N_19684);
xnor U22317 (N_22317,N_18923,N_19198);
or U22318 (N_22318,N_21211,N_21432);
or U22319 (N_22319,N_20619,N_20295);
nand U22320 (N_22320,N_18832,N_21873);
and U22321 (N_22321,N_19595,N_20533);
and U22322 (N_22322,N_20328,N_21729);
nand U22323 (N_22323,N_19054,N_20599);
or U22324 (N_22324,N_21518,N_19709);
nand U22325 (N_22325,N_20870,N_20008);
and U22326 (N_22326,N_20217,N_19824);
nor U22327 (N_22327,N_18858,N_21195);
nor U22328 (N_22328,N_20427,N_19826);
or U22329 (N_22329,N_21577,N_19476);
nand U22330 (N_22330,N_20289,N_21085);
xnor U22331 (N_22331,N_19532,N_19829);
xnor U22332 (N_22332,N_20866,N_21567);
and U22333 (N_22333,N_18966,N_21502);
nor U22334 (N_22334,N_19098,N_21062);
or U22335 (N_22335,N_19755,N_19208);
or U22336 (N_22336,N_20323,N_20594);
or U22337 (N_22337,N_20284,N_18827);
xnor U22338 (N_22338,N_21381,N_21300);
and U22339 (N_22339,N_21074,N_21113);
and U22340 (N_22340,N_18934,N_20586);
nand U22341 (N_22341,N_21176,N_20054);
or U22342 (N_22342,N_21564,N_19280);
or U22343 (N_22343,N_20944,N_20610);
nand U22344 (N_22344,N_20511,N_21116);
nand U22345 (N_22345,N_19999,N_19194);
nor U22346 (N_22346,N_20147,N_19129);
nand U22347 (N_22347,N_21140,N_19803);
nor U22348 (N_22348,N_19410,N_20875);
nor U22349 (N_22349,N_19872,N_21052);
and U22350 (N_22350,N_19146,N_21565);
nand U22351 (N_22351,N_20205,N_19994);
and U22352 (N_22352,N_21308,N_20620);
nand U22353 (N_22353,N_20688,N_20898);
xor U22354 (N_22354,N_20252,N_21746);
and U22355 (N_22355,N_21479,N_21561);
nand U22356 (N_22356,N_20945,N_20265);
or U22357 (N_22357,N_19626,N_19420);
nor U22358 (N_22358,N_19859,N_19540);
and U22359 (N_22359,N_20521,N_21799);
and U22360 (N_22360,N_19850,N_20987);
and U22361 (N_22361,N_21820,N_21498);
xnor U22362 (N_22362,N_19016,N_20431);
or U22363 (N_22363,N_19401,N_21196);
nor U22364 (N_22364,N_20260,N_19195);
and U22365 (N_22365,N_19483,N_19559);
nand U22366 (N_22366,N_21829,N_19199);
nor U22367 (N_22367,N_20814,N_19670);
nor U22368 (N_22368,N_21844,N_20117);
or U22369 (N_22369,N_20787,N_19159);
nand U22370 (N_22370,N_21538,N_19970);
and U22371 (N_22371,N_20137,N_19038);
nand U22372 (N_22372,N_20644,N_21584);
nor U22373 (N_22373,N_21633,N_19172);
nor U22374 (N_22374,N_19853,N_21676);
nor U22375 (N_22375,N_21334,N_19321);
nand U22376 (N_22376,N_18851,N_19275);
xor U22377 (N_22377,N_21126,N_18876);
and U22378 (N_22378,N_20290,N_20853);
nand U22379 (N_22379,N_19395,N_19260);
nand U22380 (N_22380,N_19051,N_19525);
and U22381 (N_22381,N_21015,N_19593);
and U22382 (N_22382,N_20308,N_19273);
nor U22383 (N_22383,N_21271,N_20266);
or U22384 (N_22384,N_18772,N_20551);
nor U22385 (N_22385,N_19691,N_21213);
nor U22386 (N_22386,N_19946,N_19513);
nor U22387 (N_22387,N_21745,N_21467);
or U22388 (N_22388,N_18754,N_20525);
and U22389 (N_22389,N_21110,N_19681);
nand U22390 (N_22390,N_20999,N_21012);
or U22391 (N_22391,N_19640,N_20238);
and U22392 (N_22392,N_20185,N_19864);
nor U22393 (N_22393,N_21672,N_19364);
nand U22394 (N_22394,N_21153,N_20090);
xnor U22395 (N_22395,N_20352,N_19696);
nor U22396 (N_22396,N_19202,N_18949);
nand U22397 (N_22397,N_19599,N_20622);
and U22398 (N_22398,N_20589,N_20961);
nand U22399 (N_22399,N_21712,N_21184);
and U22400 (N_22400,N_21587,N_19676);
or U22401 (N_22401,N_19522,N_21658);
nand U22402 (N_22402,N_19882,N_20732);
or U22403 (N_22403,N_20059,N_21105);
nor U22404 (N_22404,N_19607,N_18785);
nand U22405 (N_22405,N_19478,N_20409);
and U22406 (N_22406,N_19486,N_20274);
or U22407 (N_22407,N_18958,N_20733);
or U22408 (N_22408,N_20460,N_21456);
nor U22409 (N_22409,N_19419,N_21546);
xor U22410 (N_22410,N_20724,N_19399);
and U22411 (N_22411,N_19050,N_19017);
or U22412 (N_22412,N_20901,N_20316);
and U22413 (N_22413,N_21047,N_20997);
and U22414 (N_22414,N_21529,N_21373);
nand U22415 (N_22415,N_21499,N_21442);
or U22416 (N_22416,N_19367,N_19865);
nor U22417 (N_22417,N_21673,N_21029);
or U22418 (N_22418,N_19049,N_18753);
nand U22419 (N_22419,N_20869,N_20570);
nand U22420 (N_22420,N_21000,N_19092);
and U22421 (N_22421,N_21115,N_21637);
or U22422 (N_22422,N_21752,N_20188);
and U22423 (N_22423,N_19903,N_19262);
or U22424 (N_22424,N_20407,N_21107);
nand U22425 (N_22425,N_18946,N_19656);
nand U22426 (N_22426,N_19045,N_21194);
and U22427 (N_22427,N_21679,N_19492);
and U22428 (N_22428,N_20009,N_19223);
xor U22429 (N_22429,N_19365,N_21329);
nor U22430 (N_22430,N_20239,N_18955);
or U22431 (N_22431,N_20105,N_19108);
nor U22432 (N_22432,N_20004,N_18954);
and U22433 (N_22433,N_20527,N_20783);
nand U22434 (N_22434,N_20327,N_19651);
nor U22435 (N_22435,N_21321,N_21108);
xor U22436 (N_22436,N_21152,N_20084);
nor U22437 (N_22437,N_19213,N_21609);
nor U22438 (N_22438,N_19391,N_20028);
and U22439 (N_22439,N_18808,N_19249);
or U22440 (N_22440,N_20285,N_20498);
or U22441 (N_22441,N_18812,N_19241);
or U22442 (N_22442,N_21850,N_19631);
nor U22443 (N_22443,N_20580,N_20091);
and U22444 (N_22444,N_19563,N_20731);
nand U22445 (N_22445,N_20949,N_20675);
nand U22446 (N_22446,N_19370,N_20462);
xnor U22447 (N_22447,N_21418,N_21288);
xor U22448 (N_22448,N_20834,N_19490);
nor U22449 (N_22449,N_19974,N_21693);
nand U22450 (N_22450,N_20899,N_20660);
nor U22451 (N_22451,N_18863,N_20144);
xor U22452 (N_22452,N_19675,N_19118);
and U22453 (N_22453,N_20254,N_21772);
or U22454 (N_22454,N_19579,N_21023);
or U22455 (N_22455,N_21550,N_20851);
nor U22456 (N_22456,N_20077,N_19472);
and U22457 (N_22457,N_20403,N_20678);
nor U22458 (N_22458,N_19962,N_18974);
nand U22459 (N_22459,N_18964,N_20631);
nor U22460 (N_22460,N_21681,N_19685);
nor U22461 (N_22461,N_20455,N_20503);
and U22462 (N_22462,N_21616,N_19489);
and U22463 (N_22463,N_19136,N_19533);
and U22464 (N_22464,N_20356,N_21169);
nand U22465 (N_22465,N_19584,N_21714);
nand U22466 (N_22466,N_19801,N_19959);
or U22467 (N_22467,N_20671,N_21059);
nor U22468 (N_22468,N_19932,N_19080);
or U22469 (N_22469,N_20659,N_21724);
or U22470 (N_22470,N_21067,N_21433);
or U22471 (N_22471,N_19708,N_20518);
nand U22472 (N_22472,N_20794,N_21227);
or U22473 (N_22473,N_20501,N_19812);
nor U22474 (N_22474,N_20640,N_20294);
and U22475 (N_22475,N_20197,N_21659);
and U22476 (N_22476,N_21002,N_20952);
and U22477 (N_22477,N_19565,N_20563);
nand U22478 (N_22478,N_20234,N_20485);
nor U22479 (N_22479,N_19683,N_20206);
or U22480 (N_22480,N_21603,N_18802);
nor U22481 (N_22481,N_20296,N_20712);
nor U22482 (N_22482,N_19784,N_18810);
or U22483 (N_22483,N_20790,N_21845);
and U22484 (N_22484,N_20447,N_20364);
nor U22485 (N_22485,N_19914,N_20288);
or U22486 (N_22486,N_21824,N_21044);
or U22487 (N_22487,N_19272,N_20071);
or U22488 (N_22488,N_19369,N_20826);
nor U22489 (N_22489,N_19887,N_19988);
and U22490 (N_22490,N_21147,N_20494);
nand U22491 (N_22491,N_20016,N_21650);
xnor U22492 (N_22492,N_18990,N_21806);
nand U22493 (N_22493,N_21078,N_21142);
and U22494 (N_22494,N_20613,N_20492);
and U22495 (N_22495,N_20968,N_19508);
or U22496 (N_22496,N_20947,N_20287);
and U22497 (N_22497,N_21394,N_21045);
or U22498 (N_22498,N_20611,N_21854);
nor U22499 (N_22499,N_19966,N_19892);
nor U22500 (N_22500,N_20104,N_20726);
nand U22501 (N_22501,N_19935,N_19243);
or U22502 (N_22502,N_21556,N_20362);
nor U22503 (N_22503,N_20411,N_19233);
and U22504 (N_22504,N_19375,N_20934);
and U22505 (N_22505,N_20791,N_20884);
and U22506 (N_22506,N_21290,N_20958);
nor U22507 (N_22507,N_20481,N_21769);
nor U22508 (N_22508,N_21016,N_20542);
or U22509 (N_22509,N_21384,N_20842);
or U22510 (N_22510,N_21253,N_21594);
nand U22511 (N_22511,N_20396,N_18957);
xor U22512 (N_22512,N_18791,N_19646);
and U22513 (N_22513,N_19333,N_19447);
xnor U22514 (N_22514,N_20577,N_19404);
xor U22515 (N_22515,N_19142,N_20954);
nand U22516 (N_22516,N_20386,N_21114);
and U22517 (N_22517,N_19345,N_20978);
and U22518 (N_22518,N_21208,N_19542);
nor U22519 (N_22519,N_20768,N_19292);
and U22520 (N_22520,N_20931,N_19298);
nand U22521 (N_22521,N_18902,N_20806);
or U22522 (N_22522,N_19155,N_20219);
nand U22523 (N_22523,N_18854,N_20349);
nand U22524 (N_22524,N_21666,N_20685);
nand U22525 (N_22525,N_18820,N_21156);
or U22526 (N_22526,N_20699,N_20957);
and U22527 (N_22527,N_20559,N_20849);
or U22528 (N_22528,N_20401,N_21794);
nand U22529 (N_22529,N_21314,N_21415);
xnor U22530 (N_22530,N_19197,N_21600);
and U22531 (N_22531,N_20932,N_21204);
nor U22532 (N_22532,N_19759,N_20867);
nand U22533 (N_22533,N_21217,N_20761);
and U22534 (N_22534,N_19820,N_19622);
and U22535 (N_22535,N_21171,N_20771);
nand U22536 (N_22536,N_20663,N_19658);
and U22537 (N_22537,N_21361,N_20588);
nand U22538 (N_22538,N_19113,N_19911);
or U22539 (N_22539,N_21001,N_21489);
nor U22540 (N_22540,N_19465,N_20321);
xnor U22541 (N_22541,N_20140,N_19140);
xor U22542 (N_22542,N_19063,N_18846);
nor U22543 (N_22543,N_19799,N_19493);
xor U22544 (N_22544,N_21285,N_19230);
or U22545 (N_22545,N_20207,N_21277);
xnor U22546 (N_22546,N_20453,N_20574);
nand U22547 (N_22547,N_20564,N_21243);
or U22548 (N_22548,N_21219,N_19036);
or U22549 (N_22549,N_19433,N_18915);
nand U22550 (N_22550,N_20039,N_19068);
and U22551 (N_22551,N_19939,N_18794);
nand U22552 (N_22552,N_19497,N_19904);
nor U22553 (N_22553,N_19529,N_21573);
nand U22554 (N_22554,N_19217,N_21508);
nor U22555 (N_22555,N_21695,N_19250);
nand U22556 (N_22556,N_19101,N_20341);
and U22557 (N_22557,N_20939,N_21509);
nand U22558 (N_22558,N_19398,N_19077);
nor U22559 (N_22559,N_20102,N_20108);
or U22560 (N_22560,N_21651,N_20804);
and U22561 (N_22561,N_18980,N_21606);
nor U22562 (N_22562,N_19767,N_20720);
nor U22563 (N_22563,N_18991,N_19699);
nand U22564 (N_22564,N_20344,N_19783);
nor U22565 (N_22565,N_20278,N_19306);
and U22566 (N_22566,N_19923,N_19201);
and U22567 (N_22567,N_21111,N_20831);
or U22568 (N_22568,N_20368,N_21040);
or U22569 (N_22569,N_21560,N_19920);
and U22570 (N_22570,N_20882,N_18804);
xor U22571 (N_22571,N_20497,N_20753);
nand U22572 (N_22572,N_19214,N_19457);
or U22573 (N_22573,N_20656,N_19965);
xnor U22574 (N_22574,N_21648,N_21795);
nand U22575 (N_22575,N_18811,N_21601);
nand U22576 (N_22576,N_19421,N_18829);
and U22577 (N_22577,N_19341,N_21122);
nor U22578 (N_22578,N_20380,N_21425);
and U22579 (N_22579,N_18885,N_19539);
or U22580 (N_22580,N_20981,N_19507);
or U22581 (N_22581,N_19921,N_21033);
and U22582 (N_22582,N_19944,N_20522);
or U22583 (N_22583,N_20648,N_21354);
xor U22584 (N_22584,N_19949,N_19152);
nand U22585 (N_22585,N_21141,N_20182);
and U22586 (N_22586,N_20711,N_19995);
and U22587 (N_22587,N_20778,N_21031);
and U22588 (N_22588,N_19026,N_20043);
or U22589 (N_22589,N_19384,N_20754);
nor U22590 (N_22590,N_19808,N_20502);
and U22591 (N_22591,N_20744,N_20641);
or U22592 (N_22592,N_21743,N_19878);
xor U22593 (N_22593,N_19566,N_21582);
or U22594 (N_22594,N_19671,N_19143);
and U22595 (N_22595,N_21691,N_20624);
nand U22596 (N_22596,N_20075,N_19083);
or U22597 (N_22597,N_19677,N_20576);
or U22598 (N_22598,N_20097,N_19373);
and U22599 (N_22599,N_20151,N_21364);
nand U22600 (N_22600,N_20661,N_21667);
nand U22601 (N_22601,N_20860,N_21662);
xnor U22602 (N_22602,N_20992,N_19734);
xor U22603 (N_22603,N_21351,N_19717);
nand U22604 (N_22604,N_20904,N_19276);
nand U22605 (N_22605,N_20818,N_21039);
nand U22606 (N_22606,N_21054,N_21575);
nor U22607 (N_22607,N_20367,N_20680);
nand U22608 (N_22608,N_21678,N_21740);
nor U22609 (N_22609,N_18782,N_19724);
or U22610 (N_22610,N_20240,N_18988);
nand U22611 (N_22611,N_21215,N_20566);
nand U22612 (N_22612,N_19313,N_19327);
or U22613 (N_22613,N_19079,N_19936);
nand U22614 (N_22614,N_19852,N_19895);
nor U22615 (N_22615,N_19839,N_20520);
nor U22616 (N_22616,N_21408,N_21770);
nand U22617 (N_22617,N_21134,N_21283);
or U22618 (N_22618,N_20775,N_21621);
or U22619 (N_22619,N_20528,N_20275);
nor U22620 (N_22620,N_21372,N_19470);
xor U22621 (N_22621,N_19251,N_21086);
nor U22622 (N_22622,N_18899,N_21292);
xnor U22623 (N_22623,N_21352,N_19466);
nand U22624 (N_22624,N_20519,N_20777);
nand U22625 (N_22625,N_19288,N_21028);
nand U22626 (N_22626,N_21090,N_21203);
and U22627 (N_22627,N_19424,N_21768);
nand U22628 (N_22628,N_21341,N_21480);
nor U22629 (N_22629,N_18801,N_21607);
and U22630 (N_22630,N_21395,N_20006);
nand U22631 (N_22631,N_21694,N_20314);
and U22632 (N_22632,N_19461,N_18843);
nor U22633 (N_22633,N_19156,N_20496);
xor U22634 (N_22634,N_19621,N_21201);
and U22635 (N_22635,N_20198,N_20618);
or U22636 (N_22636,N_19431,N_20883);
and U22637 (N_22637,N_20222,N_18869);
and U22638 (N_22638,N_21735,N_20479);
nand U22639 (N_22639,N_21501,N_19103);
nand U22640 (N_22640,N_19084,N_20051);
nor U22641 (N_22641,N_19408,N_19031);
nor U22642 (N_22642,N_19035,N_21010);
nand U22643 (N_22643,N_19869,N_18894);
nor U22644 (N_22644,N_21513,N_20756);
xor U22645 (N_22645,N_21075,N_18781);
nand U22646 (N_22646,N_21494,N_19669);
and U22647 (N_22647,N_20692,N_21608);
nand U22648 (N_22648,N_19334,N_21069);
xnor U22649 (N_22649,N_19360,N_21284);
nand U22650 (N_22650,N_21532,N_21846);
nor U22651 (N_22651,N_21377,N_18936);
or U22652 (N_22652,N_19981,N_19910);
nand U22653 (N_22653,N_21671,N_20158);
nor U22654 (N_22654,N_19349,N_21212);
xor U22655 (N_22655,N_19114,N_19043);
nand U22656 (N_22656,N_19188,N_20994);
nor U22657 (N_22657,N_19703,N_20417);
or U22658 (N_22658,N_20034,N_18834);
and U22659 (N_22659,N_21614,N_20046);
nor U22660 (N_22660,N_19753,N_21409);
and U22661 (N_22661,N_19598,N_19039);
nor U22662 (N_22662,N_19207,N_21544);
nor U22663 (N_22663,N_19456,N_19347);
nor U22664 (N_22664,N_21506,N_20924);
and U22665 (N_22665,N_20821,N_21365);
and U22666 (N_22666,N_21863,N_19834);
xnor U22667 (N_22667,N_18861,N_20070);
nand U22668 (N_22668,N_21443,N_19560);
or U22669 (N_22669,N_21861,N_20895);
nor U22670 (N_22670,N_20388,N_20025);
nor U22671 (N_22671,N_21574,N_19960);
and U22672 (N_22672,N_19263,N_21697);
and U22673 (N_22673,N_19320,N_21187);
or U22674 (N_22674,N_20334,N_21017);
or U22675 (N_22675,N_21654,N_21624);
nand U22676 (N_22676,N_19134,N_19941);
and U22677 (N_22677,N_21155,N_20896);
or U22678 (N_22678,N_20666,N_19307);
nor U22679 (N_22679,N_19719,N_21036);
or U22680 (N_22680,N_20300,N_19167);
nor U22681 (N_22681,N_20333,N_19071);
or U22682 (N_22682,N_21081,N_19898);
xor U22683 (N_22683,N_19510,N_19512);
xor U22684 (N_22684,N_20313,N_20478);
nand U22685 (N_22685,N_21024,N_21668);
or U22686 (N_22686,N_21101,N_19585);
xor U22687 (N_22687,N_20569,N_19601);
nor U22688 (N_22688,N_19690,N_20406);
nor U22689 (N_22689,N_21630,N_19543);
and U22690 (N_22690,N_20693,N_21438);
nor U22691 (N_22691,N_19519,N_21708);
nor U22692 (N_22692,N_20361,N_18792);
and U22693 (N_22693,N_18823,N_21399);
and U22694 (N_22694,N_20967,N_19090);
nor U22695 (N_22695,N_21233,N_19958);
nor U22696 (N_22696,N_21484,N_19500);
and U22697 (N_22697,N_20247,N_20858);
or U22698 (N_22698,N_21043,N_20484);
and U22699 (N_22699,N_21249,N_20540);
nor U22700 (N_22700,N_20788,N_18797);
or U22701 (N_22701,N_20402,N_20859);
or U22702 (N_22702,N_21791,N_20658);
nand U22703 (N_22703,N_21291,N_19314);
nand U22704 (N_22704,N_18825,N_19442);
xor U22705 (N_22705,N_20141,N_20458);
xnor U22706 (N_22706,N_21093,N_19823);
or U22707 (N_22707,N_19023,N_21177);
nor U22708 (N_22708,N_20874,N_18855);
and U22709 (N_22709,N_20444,N_19728);
or U22710 (N_22710,N_20398,N_21259);
nor U22711 (N_22711,N_21711,N_19239);
or U22712 (N_22712,N_20114,N_20040);
or U22713 (N_22713,N_20113,N_21018);
or U22714 (N_22714,N_18788,N_20602);
or U22715 (N_22715,N_21132,N_20488);
or U22716 (N_22716,N_19425,N_18835);
nand U22717 (N_22717,N_21786,N_20888);
nor U22718 (N_22718,N_21037,N_21336);
or U22719 (N_22719,N_20111,N_20816);
nand U22720 (N_22720,N_20264,N_21455);
nand U22721 (N_22721,N_20700,N_19491);
xor U22722 (N_22722,N_21583,N_20795);
or U22723 (N_22723,N_21526,N_20543);
nor U22724 (N_22724,N_19064,N_21701);
and U22725 (N_22725,N_20050,N_20751);
and U22726 (N_22726,N_18984,N_19992);
nand U22727 (N_22727,N_19505,N_20454);
and U22728 (N_22728,N_21732,N_21367);
xor U22729 (N_22729,N_20893,N_21112);
xnor U22730 (N_22730,N_20312,N_21413);
nand U22731 (N_22731,N_19615,N_19817);
nor U22732 (N_22732,N_19258,N_20412);
and U22733 (N_22733,N_19567,N_21838);
and U22734 (N_22734,N_19257,N_21461);
nor U22735 (N_22735,N_19319,N_18815);
or U22736 (N_22736,N_20956,N_20257);
nor U22737 (N_22737,N_20796,N_20735);
nand U22738 (N_22738,N_20461,N_19743);
xnor U22739 (N_22739,N_21414,N_20824);
and U22740 (N_22740,N_21182,N_21034);
and U22741 (N_22741,N_20390,N_19997);
or U22742 (N_22742,N_19550,N_19538);
or U22743 (N_22743,N_21080,N_20915);
and U22744 (N_22744,N_20220,N_19141);
nor U22745 (N_22745,N_21530,N_21427);
nor U22746 (N_22746,N_20336,N_19247);
nand U22747 (N_22747,N_20903,N_19866);
or U22748 (N_22748,N_20508,N_18875);
nand U22749 (N_22749,N_20940,N_20178);
nand U22750 (N_22750,N_19569,N_19012);
nor U22751 (N_22751,N_21295,N_18870);
nor U22752 (N_22752,N_18981,N_19982);
nor U22753 (N_22753,N_21106,N_19175);
and U22754 (N_22754,N_19348,N_21220);
nand U22755 (N_22755,N_19800,N_20236);
xnor U22756 (N_22756,N_21423,N_20583);
and U22757 (N_22757,N_20233,N_21858);
nor U22758 (N_22758,N_19287,N_20363);
and U22759 (N_22759,N_19406,N_20906);
nor U22760 (N_22760,N_19546,N_20282);
or U22761 (N_22761,N_19679,N_21761);
and U22762 (N_22762,N_21706,N_20717);
or U22763 (N_22763,N_19590,N_20789);
or U22764 (N_22764,N_19177,N_21149);
nor U22765 (N_22765,N_20393,N_21520);
or U22766 (N_22766,N_21032,N_19104);
nand U22767 (N_22767,N_19738,N_20581);
and U22768 (N_22768,N_19534,N_19877);
or U22769 (N_22769,N_20152,N_20989);
nand U22770 (N_22770,N_19309,N_21779);
and U22771 (N_22771,N_19236,N_20770);
and U22772 (N_22772,N_20415,N_20055);
and U22773 (N_22773,N_21092,N_20376);
nand U22774 (N_22774,N_19215,N_21404);
nand U22775 (N_22775,N_19792,N_21512);
nand U22776 (N_22776,N_21748,N_20337);
nor U22777 (N_22777,N_20150,N_18947);
nand U22778 (N_22778,N_20808,N_20670);
and U22779 (N_22779,N_19764,N_18963);
nand U22780 (N_22780,N_21623,N_21527);
or U22781 (N_22781,N_20499,N_21462);
or U22782 (N_22782,N_18784,N_19417);
nand U22783 (N_22783,N_19067,N_20617);
and U22784 (N_22784,N_21239,N_18765);
xnor U22785 (N_22785,N_20913,N_19030);
and U22786 (N_22786,N_21391,N_20420);
and U22787 (N_22787,N_21100,N_19128);
or U22788 (N_22788,N_20112,N_18774);
nand U22789 (N_22789,N_20755,N_20972);
nand U22790 (N_22790,N_21750,N_20799);
xor U22791 (N_22791,N_21751,N_19612);
nand U22792 (N_22792,N_18983,N_21622);
and U22793 (N_22793,N_20682,N_20183);
nand U22794 (N_22794,N_20184,N_19305);
nor U22795 (N_22795,N_21159,N_21759);
nor U22796 (N_22796,N_19284,N_21348);
nor U22797 (N_22797,N_21198,N_19168);
and U22798 (N_22798,N_21421,N_19680);
xnor U22799 (N_22799,N_18752,N_21856);
or U22800 (N_22800,N_21629,N_19511);
or U22801 (N_22801,N_20486,N_20330);
and U22802 (N_22802,N_20397,N_20331);
or U22803 (N_22803,N_21645,N_21653);
xnor U22804 (N_22804,N_20405,N_20532);
or U22805 (N_22805,N_18761,N_21179);
or U22806 (N_22806,N_21517,N_19097);
nor U22807 (N_22807,N_19846,N_19976);
and U22808 (N_22808,N_19605,N_18845);
nor U22809 (N_22809,N_20691,N_20524);
xor U22810 (N_22810,N_19636,N_19256);
nor U22811 (N_22811,N_21682,N_20442);
and U22812 (N_22812,N_18878,N_20335);
nand U22813 (N_22813,N_19524,N_19150);
nand U22814 (N_22814,N_19891,N_18828);
or U22815 (N_22815,N_20811,N_18952);
and U22816 (N_22816,N_20297,N_20092);
and U22817 (N_22817,N_20339,N_20326);
and U22818 (N_22818,N_20057,N_19331);
xnor U22819 (N_22819,N_20448,N_21294);
or U22820 (N_22820,N_18943,N_21661);
nor U22821 (N_22821,N_21346,N_19203);
and U22822 (N_22822,N_20470,N_18951);
nand U22823 (N_22823,N_20925,N_20168);
or U22824 (N_22824,N_21859,N_19624);
and U22825 (N_22825,N_19183,N_19890);
xor U22826 (N_22826,N_20468,N_21602);
and U22827 (N_22827,N_21797,N_21265);
or U22828 (N_22828,N_19625,N_21087);
or U22829 (N_22829,N_21723,N_19504);
or U22830 (N_22830,N_20304,N_18889);
and U22831 (N_22831,N_20283,N_19889);
xor U22832 (N_22832,N_21205,N_18871);
or U22833 (N_22833,N_19434,N_20446);
xor U22834 (N_22834,N_20472,N_21476);
or U22835 (N_22835,N_18907,N_18817);
nor U22836 (N_22836,N_19462,N_19028);
nor U22837 (N_22837,N_20375,N_19322);
and U22838 (N_22838,N_20553,N_20873);
xnor U22839 (N_22839,N_19147,N_19793);
and U22840 (N_22840,N_21380,N_21568);
xor U22841 (N_22841,N_19444,N_19805);
or U22842 (N_22842,N_20902,N_21303);
nor U22843 (N_22843,N_19983,N_21181);
nor U22844 (N_22844,N_20082,N_20044);
nand U22845 (N_22845,N_20515,N_21481);
nand U22846 (N_22846,N_20698,N_19848);
nor U22847 (N_22847,N_20083,N_20781);
nand U22848 (N_22848,N_19521,N_21814);
nor U22849 (N_22849,N_19574,N_19455);
and U22850 (N_22850,N_21787,N_19008);
or U22851 (N_22851,N_19961,N_19240);
and U22852 (N_22852,N_20845,N_20916);
and U22853 (N_22853,N_19804,N_18976);
and U22854 (N_22854,N_21343,N_19771);
or U22855 (N_22855,N_20408,N_20729);
and U22856 (N_22856,N_18881,N_19700);
nand U22857 (N_22857,N_20986,N_19843);
nor U22858 (N_22858,N_19022,N_19304);
and U22859 (N_22859,N_21739,N_18790);
nor U22860 (N_22860,N_21312,N_19034);
nand U22861 (N_22861,N_20784,N_20052);
nand U22862 (N_22862,N_19752,N_19343);
nor U22863 (N_22863,N_20107,N_20549);
and U22864 (N_22864,N_21765,N_18959);
nor U22865 (N_22865,N_20837,N_19053);
nor U22866 (N_22866,N_20143,N_19340);
nand U22867 (N_22867,N_20552,N_19596);
or U22868 (N_22868,N_19060,N_19238);
nand U22869 (N_22869,N_20162,N_21131);
xnor U22870 (N_22870,N_18874,N_19357);
nor U22871 (N_22871,N_21598,N_21617);
nand U22872 (N_22872,N_20654,N_20358);
nand U22873 (N_22873,N_20955,N_21089);
and U22874 (N_22874,N_21831,N_20428);
nand U22875 (N_22875,N_21709,N_19402);
or U22876 (N_22876,N_19674,N_19940);
and U22877 (N_22877,N_21096,N_20132);
or U22878 (N_22878,N_20679,N_21698);
nor U22879 (N_22879,N_20636,N_19002);
nor U22880 (N_22880,N_21009,N_21528);
xor U22881 (N_22881,N_21315,N_20988);
nor U22882 (N_22882,N_19379,N_18928);
or U22883 (N_22883,N_19356,N_21264);
nor U22884 (N_22884,N_18809,N_19875);
nor U22885 (N_22885,N_19412,N_20056);
nor U22886 (N_22886,N_21777,N_20325);
nand U22887 (N_22887,N_21559,N_20157);
or U22888 (N_22888,N_20965,N_19007);
and U22889 (N_22889,N_20669,N_20387);
and U22890 (N_22890,N_21807,N_21547);
nand U22891 (N_22891,N_19885,N_20136);
or U22892 (N_22892,N_21146,N_20900);
nor U22893 (N_22893,N_18892,N_19165);
xor U22894 (N_22894,N_20561,N_21516);
or U22895 (N_22895,N_20962,N_19673);
nand U22896 (N_22896,N_20109,N_21389);
nor U22897 (N_22897,N_19011,N_19748);
or U22898 (N_22898,N_21082,N_19482);
nand U22899 (N_22899,N_21466,N_20230);
nor U22900 (N_22900,N_18770,N_19768);
and U22901 (N_22901,N_18769,N_20585);
nand U22902 (N_22902,N_20854,N_18773);
xnor U22903 (N_22903,N_19953,N_19110);
and U22904 (N_22904,N_20647,N_21715);
nor U22905 (N_22905,N_20959,N_21548);
or U22906 (N_22906,N_21226,N_19969);
nand U22907 (N_22907,N_20041,N_21254);
or U22908 (N_22908,N_20471,N_20607);
nand U22909 (N_22909,N_18986,N_21157);
xnor U22910 (N_22910,N_20303,N_19857);
or U22911 (N_22911,N_19105,N_19736);
nor U22912 (N_22912,N_20809,N_20627);
and U22913 (N_22913,N_19643,N_20418);
or U22914 (N_22914,N_18796,N_20366);
and U22915 (N_22915,N_21255,N_20459);
nand U22916 (N_22916,N_20474,N_19855);
or U22917 (N_22917,N_20891,N_20643);
and U22918 (N_22918,N_19561,N_20203);
nand U22919 (N_22919,N_19162,N_19514);
xor U22920 (N_22920,N_20359,N_19169);
nand U22921 (N_22921,N_20894,N_19242);
nand U22922 (N_22922,N_20439,N_21819);
or U22923 (N_22923,N_21118,N_20759);
nand U22924 (N_22924,N_19751,N_19020);
or U22925 (N_22925,N_19578,N_19739);
or U22926 (N_22926,N_21210,N_21792);
nor U22927 (N_22927,N_20319,N_19464);
nand U22928 (N_22928,N_21472,N_21719);
xnor U22929 (N_22929,N_20908,N_20372);
and U22930 (N_22930,N_19763,N_21738);
nand U22931 (N_22931,N_21519,N_21060);
nand U22932 (N_22932,N_21449,N_20829);
and U22933 (N_22933,N_19902,N_20943);
nand U22934 (N_22934,N_21073,N_21317);
and U22935 (N_22935,N_19571,N_21702);
nand U22936 (N_22936,N_20120,N_21847);
nand U22937 (N_22937,N_19588,N_19109);
xor U22938 (N_22938,N_19986,N_21228);
and U22939 (N_22939,N_19623,N_21393);
nor U22940 (N_22940,N_19467,N_19908);
nor U22941 (N_22941,N_20465,N_20094);
and U22942 (N_22942,N_19057,N_19609);
and U22943 (N_22943,N_20877,N_19160);
and U22944 (N_22944,N_19040,N_20175);
or U22945 (N_22945,N_20912,N_20489);
or U22946 (N_22946,N_19414,N_19184);
or U22947 (N_22947,N_21310,N_18942);
nor U22948 (N_22948,N_21445,N_19443);
nor U22949 (N_22949,N_19449,N_21065);
or U22950 (N_22950,N_19723,N_18901);
nand U22951 (N_22951,N_21742,N_20615);
nand U22952 (N_22952,N_19027,N_20623);
and U22953 (N_22953,N_19225,N_18822);
and U22954 (N_22954,N_20719,N_21251);
nor U22955 (N_22955,N_19115,N_20422);
nand U22956 (N_22956,N_19126,N_21689);
nor U22957 (N_22957,N_20086,N_20449);
and U22958 (N_22958,N_19899,N_21150);
or U22959 (N_22959,N_19409,N_21038);
or U22960 (N_22960,N_20625,N_20706);
and U22961 (N_22961,N_19290,N_21297);
or U22962 (N_22962,N_19388,N_20819);
nor U22963 (N_22963,N_18763,N_19779);
nor U22964 (N_22964,N_21669,N_18895);
nand U22965 (N_22965,N_21162,N_21453);
nor U22966 (N_22966,N_20229,N_18994);
or U22967 (N_22967,N_20708,N_21490);
or U22968 (N_22968,N_21405,N_20400);
nand U22969 (N_22969,N_21431,N_19718);
and U22970 (N_22970,N_20823,N_19004);
or U22971 (N_22971,N_18919,N_19496);
or U22972 (N_22972,N_19576,N_18766);
or U22973 (N_22973,N_19573,N_19463);
nor U22974 (N_22974,N_18972,N_20011);
and U22975 (N_22975,N_21731,N_20404);
and U22976 (N_22976,N_19663,N_20582);
nor U22977 (N_22977,N_19644,N_20862);
nor U22978 (N_22978,N_21478,N_20263);
xor U22979 (N_22979,N_21158,N_20123);
nor U22980 (N_22980,N_21579,N_18930);
nand U22981 (N_22981,N_21713,N_20917);
and U22982 (N_22982,N_19133,N_21733);
nor U22983 (N_22983,N_19769,N_20392);
and U22984 (N_22984,N_19647,N_21595);
xnor U22985 (N_22985,N_19021,N_19527);
nand U22986 (N_22986,N_20437,N_20918);
and U22987 (N_22987,N_20505,N_20737);
nor U22988 (N_22988,N_18888,N_19494);
or U22989 (N_22989,N_21783,N_20509);
xnor U22990 (N_22990,N_19537,N_20843);
xor U22991 (N_22991,N_19234,N_20725);
nor U22992 (N_22992,N_18758,N_21323);
or U22993 (N_22993,N_20825,N_20195);
nand U22994 (N_22994,N_19577,N_20984);
nand U22995 (N_22995,N_21855,N_21164);
nor U22996 (N_22996,N_19937,N_21664);
and U22997 (N_22997,N_21457,N_20063);
or U22998 (N_22998,N_20145,N_19174);
and U22999 (N_22999,N_21736,N_20516);
nand U23000 (N_23000,N_21707,N_21376);
and U23001 (N_23001,N_21762,N_19228);
nor U23002 (N_23002,N_19694,N_19335);
and U23003 (N_23003,N_20237,N_20299);
and U23004 (N_23004,N_19597,N_20491);
and U23005 (N_23005,N_20885,N_18975);
or U23006 (N_23006,N_21209,N_21771);
nor U23007 (N_23007,N_21767,N_20718);
and U23008 (N_23008,N_21267,N_18960);
or U23009 (N_23009,N_19316,N_19144);
nand U23010 (N_23010,N_20340,N_20739);
or U23011 (N_23011,N_21646,N_19849);
and U23012 (N_23012,N_20506,N_21866);
nor U23013 (N_23013,N_20475,N_20979);
nor U23014 (N_23014,N_19460,N_21448);
nand U23015 (N_23015,N_20354,N_19358);
or U23016 (N_23016,N_21776,N_20616);
and U23017 (N_23017,N_20469,N_20560);
or U23018 (N_23018,N_18937,N_19209);
and U23019 (N_23019,N_20936,N_21130);
nand U23020 (N_23020,N_21322,N_21871);
nand U23021 (N_23021,N_21585,N_18898);
or U23022 (N_23022,N_21375,N_20513);
xnor U23023 (N_23023,N_19070,N_21347);
or U23024 (N_23024,N_20110,N_21324);
nor U23025 (N_23025,N_19528,N_20938);
and U23026 (N_23026,N_20828,N_19871);
xor U23027 (N_23027,N_18950,N_19393);
or U23028 (N_23028,N_20510,N_21741);
nand U23029 (N_23029,N_20223,N_21403);
or U23030 (N_23030,N_21260,N_19664);
nand U23031 (N_23031,N_19336,N_19772);
nand U23032 (N_23032,N_19303,N_19787);
or U23033 (N_23033,N_20941,N_20792);
and U23034 (N_23034,N_21611,N_19518);
xnor U23035 (N_23035,N_19124,N_21325);
and U23036 (N_23036,N_20721,N_20597);
nor U23037 (N_23037,N_21221,N_21704);
nand U23038 (N_23038,N_21699,N_20369);
or U23039 (N_23039,N_20273,N_21496);
and U23040 (N_23040,N_20074,N_19712);
nor U23041 (N_23041,N_21358,N_20451);
xnor U23042 (N_23042,N_19065,N_21189);
and U23043 (N_23043,N_20514,N_20998);
and U23044 (N_23044,N_19591,N_21269);
nor U23045 (N_23045,N_21703,N_19697);
or U23046 (N_23046,N_19085,N_20235);
nor U23047 (N_23047,N_21812,N_21705);
and U23048 (N_23048,N_19971,N_20146);
and U23049 (N_23049,N_21337,N_20740);
nor U23050 (N_23050,N_20258,N_21193);
nand U23051 (N_23051,N_20694,N_19945);
nand U23052 (N_23052,N_21366,N_19161);
nor U23053 (N_23053,N_20270,N_20061);
and U23054 (N_23054,N_20905,N_21289);
and U23055 (N_23055,N_20463,N_18860);
nand U23056 (N_23056,N_21051,N_21592);
or U23057 (N_23057,N_19604,N_20204);
and U23058 (N_23058,N_19985,N_19928);
nand U23059 (N_23059,N_19894,N_18992);
xnor U23060 (N_23060,N_19744,N_19980);
nor U23061 (N_23061,N_21497,N_20982);
or U23062 (N_23062,N_19392,N_20839);
nor U23063 (N_23063,N_21370,N_19660);
nand U23064 (N_23064,N_21758,N_20381);
or U23065 (N_23065,N_18956,N_21677);
or U23066 (N_23066,N_20537,N_18914);
nor U23067 (N_23067,N_20343,N_20186);
nand U23068 (N_23068,N_19346,N_21218);
nor U23069 (N_23069,N_20127,N_19149);
nand U23070 (N_23070,N_21281,N_19611);
nor U23071 (N_23071,N_19317,N_21104);
and U23072 (N_23072,N_20703,N_19018);
nor U23073 (N_23073,N_21690,N_19166);
nor U23074 (N_23074,N_19459,N_19312);
nor U23075 (N_23075,N_21066,N_20857);
nor U23076 (N_23076,N_19868,N_18906);
or U23077 (N_23077,N_21121,N_20068);
or U23078 (N_23078,N_19355,N_20315);
and U23079 (N_23079,N_18771,N_20601);
xnor U23080 (N_23080,N_21385,N_19782);
nor U23081 (N_23081,N_21634,N_20964);
nand U23082 (N_23082,N_19716,N_20272);
nor U23083 (N_23083,N_21454,N_18908);
and U23084 (N_23084,N_21515,N_21488);
nand U23085 (N_23085,N_18864,N_19122);
nand U23086 (N_23086,N_19555,N_20748);
or U23087 (N_23087,N_19807,N_19806);
nand U23088 (N_23088,N_21826,N_19058);
and U23089 (N_23089,N_19987,N_21700);
and U23090 (N_23090,N_19610,N_19991);
or U23091 (N_23091,N_19205,N_21247);
and U23092 (N_23092,N_19193,N_21307);
and U23093 (N_23093,N_21299,N_21216);
or U23094 (N_23094,N_19773,N_19770);
or U23095 (N_23095,N_18953,N_21444);
and U23096 (N_23096,N_19106,N_21599);
nor U23097 (N_23097,N_21610,N_18925);
and U23098 (N_23098,N_20707,N_19620);
nor U23099 (N_23099,N_21057,N_21828);
xnor U23100 (N_23100,N_21800,N_20573);
or U23101 (N_23101,N_19099,N_19668);
or U23102 (N_23102,N_21125,N_18890);
nand U23103 (N_23103,N_20683,N_19046);
and U23104 (N_23104,N_21027,N_21070);
or U23105 (N_23105,N_21133,N_20977);
and U23106 (N_23106,N_21417,N_19880);
xnor U23107 (N_23107,N_20684,N_19296);
nor U23108 (N_23108,N_20424,N_19332);
nor U23109 (N_23109,N_21135,N_21183);
nand U23110 (N_23110,N_18967,N_19220);
nor U23111 (N_23111,N_19754,N_21148);
nor U23112 (N_23112,N_20020,N_21278);
and U23113 (N_23113,N_20209,N_19893);
xor U23114 (N_23114,N_18918,N_20069);
and U23115 (N_23115,N_20036,N_20946);
nand U23116 (N_23116,N_19216,N_19652);
nor U23117 (N_23117,N_20922,N_19415);
or U23118 (N_23118,N_18872,N_20709);
nand U23119 (N_23119,N_19978,N_20438);
xor U23120 (N_23120,N_20365,N_18891);
nand U23121 (N_23121,N_19354,N_19686);
nand U23122 (N_23122,N_21811,N_19112);
and U23123 (N_23123,N_21388,N_18884);
nor U23124 (N_23124,N_21363,N_20487);
and U23125 (N_23125,N_21302,N_21234);
or U23126 (N_23126,N_19711,N_21241);
xor U23127 (N_23127,N_21523,N_19473);
nor U23128 (N_23128,N_21505,N_19778);
xnor U23129 (N_23129,N_19015,N_20645);
nor U23130 (N_23130,N_21020,N_19795);
xnor U23131 (N_23131,N_18987,N_20038);
nand U23132 (N_23132,N_19254,N_19842);
nor U23133 (N_23133,N_21206,N_20779);
nor U23134 (N_23134,N_20019,N_21357);
or U23135 (N_23135,N_19572,N_19117);
nor U23136 (N_23136,N_20578,N_20293);
nor U23137 (N_23137,N_18821,N_20738);
nor U23138 (N_23138,N_20017,N_19182);
nor U23139 (N_23139,N_19266,N_20758);
or U23140 (N_23140,N_18783,N_21803);
nor U23141 (N_23141,N_20728,N_19589);
nand U23142 (N_23142,N_21345,N_19775);
and U23143 (N_23143,N_20101,N_21833);
nand U23144 (N_23144,N_19326,N_21649);
xor U23145 (N_23145,N_18961,N_21246);
and U23146 (N_23146,N_19352,N_21386);
nand U23147 (N_23147,N_19672,N_21172);
or U23148 (N_23148,N_20213,N_20801);
nand U23149 (N_23149,N_20457,N_20606);
nor U23150 (N_23150,N_21620,N_21102);
nand U23151 (N_23151,N_20215,N_19137);
and U23152 (N_23152,N_21340,N_19825);
or U23153 (N_23153,N_19259,N_19973);
and U23154 (N_23154,N_19790,N_21534);
nor U23155 (N_23155,N_21091,N_21486);
nand U23156 (N_23156,N_19809,N_20155);
and U23157 (N_23157,N_20000,N_21474);
nor U23158 (N_23158,N_21261,N_18807);
or U23159 (N_23159,N_19089,N_19701);
xnor U23160 (N_23160,N_19907,N_21539);
xor U23161 (N_23161,N_18818,N_19975);
or U23162 (N_23162,N_20696,N_18924);
and U23163 (N_23163,N_21378,N_19440);
nor U23164 (N_23164,N_19888,N_21830);
nand U23165 (N_23165,N_21775,N_20512);
nor U23166 (N_23166,N_18938,N_19915);
nor U23167 (N_23167,N_20591,N_20087);
nand U23168 (N_23168,N_21644,N_18909);
nand U23169 (N_23169,N_21500,N_21225);
or U23170 (N_23170,N_20012,N_18759);
nor U23171 (N_23171,N_20609,N_21368);
nand U23172 (N_23172,N_20856,N_18973);
nor U23173 (N_23173,N_19211,N_20443);
nor U23174 (N_23174,N_20214,N_20911);
xnor U23175 (N_23175,N_20910,N_20149);
and U23176 (N_23176,N_21165,N_21003);
and U23177 (N_23177,N_20134,N_19760);
and U23178 (N_23178,N_20805,N_21604);
xnor U23179 (N_23179,N_21306,N_19066);
xor U23180 (N_23180,N_21007,N_20286);
xnor U23181 (N_23181,N_19061,N_19294);
or U23182 (N_23182,N_18755,N_20948);
nor U23183 (N_23183,N_19789,N_20493);
and U23184 (N_23184,N_19881,N_21014);
or U23185 (N_23185,N_21793,N_20425);
nand U23186 (N_23186,N_21175,N_19246);
or U23187 (N_23187,N_18939,N_19330);
nor U23188 (N_23188,N_18989,N_19368);
or U23189 (N_23189,N_21379,N_20483);
and U23190 (N_23190,N_21138,N_21718);
nor U23191 (N_23191,N_20807,N_19633);
xnor U23192 (N_23192,N_19324,N_19378);
nand U23193 (N_23193,N_19600,N_20338);
nand U23194 (N_23194,N_19727,N_18839);
and U23195 (N_23195,N_20567,N_19737);
nand U23196 (N_23196,N_19886,N_19435);
nand U23197 (N_23197,N_19231,N_21318);
nand U23198 (N_23198,N_20416,N_19847);
nand U23199 (N_23199,N_19862,N_21688);
nand U23200 (N_23200,N_19302,N_19788);
or U23201 (N_23201,N_21463,N_18775);
nor U23202 (N_23202,N_21504,N_21250);
and U23203 (N_23203,N_20190,N_18778);
nand U23204 (N_23204,N_19740,N_19549);
or U23205 (N_23205,N_18776,N_21734);
nor U23206 (N_23206,N_19602,N_19062);
and U23207 (N_23207,N_19224,N_21663);
nor U23208 (N_23208,N_19451,N_20836);
xor U23209 (N_23209,N_19180,N_19553);
and U23210 (N_23210,N_20377,N_20637);
or U23211 (N_23211,N_19501,N_20575);
nand U23212 (N_23212,N_20970,N_21392);
nand U23213 (N_23213,N_20163,N_21483);
nor U23214 (N_23214,N_19487,N_21350);
nor U23215 (N_23215,N_19100,N_21722);
or U23216 (N_23216,N_21128,N_20261);
and U23217 (N_23217,N_20232,N_20242);
nor U23218 (N_23218,N_19977,N_21842);
nor U23219 (N_23219,N_21450,N_20907);
nand U23220 (N_23220,N_18940,N_19235);
or U23221 (N_23221,N_18941,N_21728);
or U23222 (N_23222,N_19796,N_18945);
or U23223 (N_23223,N_20793,N_20088);
or U23224 (N_23224,N_20156,N_18970);
or U23225 (N_23225,N_19187,N_18921);
xnor U23226 (N_23226,N_21683,N_20847);
nand U23227 (N_23227,N_20865,N_19785);
nor U23228 (N_23228,N_20526,N_20995);
nand U23229 (N_23229,N_20584,N_19132);
nand U23230 (N_23230,N_19662,N_18979);
and U23231 (N_23231,N_20628,N_19503);
nand U23232 (N_23232,N_19437,N_21173);
and U23233 (N_23233,N_21796,N_19285);
and U23234 (N_23234,N_20937,N_21581);
and U23235 (N_23235,N_18800,N_19906);
and U23236 (N_23236,N_20015,N_21416);
xnor U23237 (N_23237,N_21543,N_19413);
nor U23238 (N_23238,N_19558,N_21458);
nor U23239 (N_23239,N_21790,N_21570);
nor U23240 (N_23240,N_19989,N_19361);
nor U23241 (N_23241,N_21035,N_20649);
or U23242 (N_23242,N_21638,N_21185);
nor U23243 (N_23243,N_21710,N_19000);
and U23244 (N_23244,N_21628,N_19639);
and U23245 (N_23245,N_19411,N_19650);
nand U23246 (N_23246,N_18969,N_21533);
or U23247 (N_23247,N_20131,N_20269);
nor U23248 (N_23248,N_21555,N_20976);
nand U23249 (N_23249,N_20715,N_19422);
and U23250 (N_23250,N_20384,N_20562);
and U23251 (N_23251,N_20353,N_19955);
or U23252 (N_23252,N_21521,N_21860);
xor U23253 (N_23253,N_20571,N_21420);
nand U23254 (N_23254,N_21180,N_20243);
nor U23255 (N_23255,N_20320,N_20665);
nand U23256 (N_23256,N_21640,N_20176);
nor U23257 (N_23257,N_20798,N_18903);
or U23258 (N_23258,N_19452,N_19912);
xnor U23259 (N_23259,N_21083,N_19475);
nor U23260 (N_23260,N_21837,N_21371);
and U23261 (N_23261,N_19278,N_20170);
nand U23262 (N_23262,N_18944,N_21747);
nor U23263 (N_23263,N_19481,N_21266);
nor U23264 (N_23264,N_19714,N_21537);
and U23265 (N_23265,N_20128,N_19867);
and U23266 (N_23266,N_21356,N_19376);
nor U23267 (N_23267,N_19488,N_19822);
and U23268 (N_23268,N_19178,N_21798);
and U23269 (N_23269,N_20414,N_20301);
nor U23270 (N_23270,N_19342,N_21053);
nand U23271 (N_23271,N_20432,N_21174);
and U23272 (N_23272,N_21344,N_21319);
nor U23273 (N_23273,N_20048,N_19917);
nand U23274 (N_23274,N_20657,N_19052);
or U23275 (N_23275,N_19245,N_21730);
and U23276 (N_23276,N_20024,N_21849);
or U23277 (N_23277,N_18985,N_19268);
nand U23278 (N_23278,N_21161,N_21514);
xnor U23279 (N_23279,N_21631,N_19922);
and U23280 (N_23280,N_19344,N_19777);
and U23281 (N_23281,N_20317,N_20887);
nand U23282 (N_23282,N_20909,N_21590);
and U23283 (N_23283,N_20886,N_18813);
nor U23284 (N_23284,N_19318,N_19432);
nand U23285 (N_23285,N_19758,N_19308);
xnor U23286 (N_23286,N_19154,N_20095);
and U23287 (N_23287,N_19186,N_19232);
nor U23288 (N_23288,N_20413,N_21656);
xnor U23289 (N_23289,N_19013,N_19884);
or U23290 (N_23290,N_20774,N_21435);
nor U23291 (N_23291,N_19628,N_20880);
nor U23292 (N_23292,N_20482,N_19695);
and U23293 (N_23293,N_19377,N_18905);
nor U23294 (N_23294,N_21588,N_18848);
nand U23295 (N_23295,N_20841,N_21809);
and U23296 (N_23296,N_21335,N_19689);
nor U23297 (N_23297,N_19189,N_20166);
and U23298 (N_23298,N_21867,N_18978);
and U23299 (N_23299,N_20555,N_19876);
or U23300 (N_23300,N_19575,N_20436);
or U23301 (N_23301,N_19819,N_19212);
nand U23302 (N_23302,N_19131,N_21262);
nand U23303 (N_23303,N_21452,N_19179);
nand U23304 (N_23304,N_19474,N_21058);
xor U23305 (N_23305,N_21785,N_21727);
nor U23306 (N_23306,N_21684,N_21612);
nor U23307 (N_23307,N_21781,N_21313);
nor U23308 (N_23308,N_19918,N_21439);
or U23309 (N_23309,N_21655,N_20216);
nor U23310 (N_23310,N_19535,N_19541);
or U23311 (N_23311,N_20382,N_20347);
or U23312 (N_23312,N_19735,N_20473);
and U23313 (N_23313,N_21625,N_19094);
and U23314 (N_23314,N_20646,N_19427);
xnor U23315 (N_23315,N_19713,N_19397);
or U23316 (N_23316,N_20115,N_19613);
nor U23317 (N_23317,N_19221,N_18795);
and U23318 (N_23318,N_21349,N_21410);
nand U23319 (N_23319,N_18929,N_20231);
xor U23320 (N_23320,N_20342,N_19741);
or U23321 (N_23321,N_18971,N_21119);
nand U23322 (N_23322,N_20122,N_20224);
or U23323 (N_23323,N_19963,N_19300);
and U23324 (N_23324,N_19942,N_20677);
and U23325 (N_23325,N_20159,N_19896);
nand U23326 (N_23326,N_20763,N_21503);
or U23327 (N_23327,N_19776,N_20596);
nor U23328 (N_23328,N_19948,N_19024);
nor U23329 (N_23329,N_19151,N_19860);
and U23330 (N_23330,N_21851,N_19900);
nor U23331 (N_23331,N_20169,N_19081);
nand U23332 (N_23332,N_19453,N_19833);
nor U23333 (N_23333,N_21309,N_21874);
or U23334 (N_23334,N_20210,N_21186);
or U23335 (N_23335,N_21129,N_21482);
nor U23336 (N_23336,N_20378,N_19924);
or U23337 (N_23337,N_20603,N_20148);
nor U23338 (N_23338,N_19498,N_20833);
and U23339 (N_23339,N_19286,N_20600);
xnor U23340 (N_23340,N_18910,N_21006);
and U23341 (N_23341,N_20129,N_20550);
nand U23342 (N_23342,N_21170,N_21531);
nand U23343 (N_23343,N_21412,N_19692);
or U23344 (N_23344,N_21274,N_20592);
xnor U23345 (N_23345,N_21424,N_19222);
nand U23346 (N_23346,N_20066,N_19095);
or U23347 (N_23347,N_19139,N_19055);
or U23348 (N_23348,N_19818,N_21202);
nor U23349 (N_23349,N_19913,N_19645);
nand U23350 (N_23350,N_20840,N_19731);
xor U23351 (N_23351,N_20001,N_19851);
or U23352 (N_23352,N_21397,N_19477);
or U23353 (N_23353,N_20960,N_21401);
or U23354 (N_23354,N_20154,N_18873);
xnor U23355 (N_23355,N_19127,N_19219);
nor U23356 (N_23356,N_20440,N_19157);
and U23357 (N_23357,N_20085,N_21041);
or U23358 (N_23358,N_20736,N_21493);
and U23359 (N_23359,N_21333,N_21355);
nor U23360 (N_23360,N_21557,N_19832);
nor U23361 (N_23361,N_21240,N_19229);
or U23362 (N_23362,N_19967,N_20172);
or U23363 (N_23363,N_19901,N_21430);
or U23364 (N_23364,N_20595,N_19382);
or U23365 (N_23365,N_20653,N_20047);
or U23366 (N_23366,N_21224,N_20173);
or U23367 (N_23367,N_20639,N_21597);
nor U23368 (N_23368,N_20309,N_19381);
or U23369 (N_23369,N_21563,N_20379);
nor U23370 (N_23370,N_19138,N_21022);
nand U23371 (N_23371,N_20202,N_20351);
or U23372 (N_23372,N_21076,N_21593);
and U23373 (N_23373,N_19374,N_20072);
nand U23374 (N_23374,N_20766,N_21369);
or U23375 (N_23375,N_20248,N_20879);
nor U23376 (N_23376,N_19568,N_20200);
or U23377 (N_23377,N_21869,N_20079);
xnor U23378 (N_23378,N_21618,N_21632);
nand U23379 (N_23379,N_21402,N_21374);
nor U23380 (N_23380,N_18962,N_19749);
xor U23381 (N_23381,N_20423,N_21327);
nand U23382 (N_23382,N_21359,N_19766);
or U23383 (N_23383,N_18893,N_21535);
or U23384 (N_23384,N_20311,N_21717);
nand U23385 (N_23385,N_20199,N_19087);
and U23386 (N_23386,N_18965,N_20897);
nor U23387 (N_23387,N_19587,N_20587);
and U23388 (N_23388,N_19858,N_21674);
nand U23389 (N_23389,N_21675,N_20629);
nand U23390 (N_23390,N_21270,N_20556);
xor U23391 (N_23391,N_20652,N_19797);
and U23392 (N_23392,N_20695,N_21050);
nand U23393 (N_23393,N_21293,N_19667);
nor U23394 (N_23394,N_21437,N_20963);
nor U23395 (N_23395,N_19428,N_18887);
xor U23396 (N_23396,N_21853,N_19742);
and U23397 (N_23397,N_18897,N_19383);
nor U23398 (N_23398,N_19931,N_20539);
xor U23399 (N_23399,N_19606,N_21398);
nand U23400 (N_23400,N_20760,N_19619);
nand U23401 (N_23401,N_19916,N_20802);
nor U23402 (N_23402,N_19927,N_21232);
nor U23403 (N_23403,N_18993,N_20572);
nor U23404 (N_23404,N_21525,N_19502);
and U23405 (N_23405,N_20385,N_18904);
nand U23406 (N_23406,N_19088,N_20306);
or U23407 (N_23407,N_20227,N_21008);
xor U23408 (N_23408,N_20452,N_19545);
and U23409 (N_23409,N_19438,N_21754);
nand U23410 (N_23410,N_18933,N_19145);
nor U23411 (N_23411,N_21236,N_19003);
and U23412 (N_23412,N_19495,N_21094);
xnor U23413 (N_23413,N_19479,N_21199);
or U23414 (N_23414,N_21256,N_20747);
xor U23415 (N_23415,N_19897,N_20876);
and U23416 (N_23416,N_20635,N_19405);
nor U23417 (N_23417,N_21237,N_20466);
nor U23418 (N_23418,N_20010,N_19351);
nor U23419 (N_23419,N_19044,N_19389);
nor U23420 (N_23420,N_19648,N_20531);
nand U23421 (N_23421,N_20171,N_21549);
nand U23422 (N_23422,N_19747,N_20194);
or U23423 (N_23423,N_19093,N_20211);
nand U23424 (N_23424,N_19255,N_20464);
or U23425 (N_23425,N_21030,N_18831);
nand U23426 (N_23426,N_21160,N_19282);
nand U23427 (N_23427,N_18756,N_20251);
or U23428 (N_23428,N_21835,N_20067);
nand U23429 (N_23429,N_18856,N_19802);
and U23430 (N_23430,N_21789,N_20991);
or U23431 (N_23431,N_21011,N_21716);
nor U23432 (N_23432,N_20517,N_19954);
nor U23433 (N_23433,N_20098,N_20612);
nand U23434 (N_23434,N_20546,N_19844);
nor U23435 (N_23435,N_21400,N_19726);
nor U23436 (N_23436,N_19181,N_21816);
and U23437 (N_23437,N_21005,N_20359);
or U23438 (N_23438,N_21539,N_19682);
nor U23439 (N_23439,N_19732,N_20396);
and U23440 (N_23440,N_20160,N_20989);
xor U23441 (N_23441,N_19034,N_20114);
nand U23442 (N_23442,N_19309,N_19178);
and U23443 (N_23443,N_20738,N_21003);
nand U23444 (N_23444,N_21171,N_21455);
or U23445 (N_23445,N_21497,N_21502);
or U23446 (N_23446,N_20467,N_18825);
or U23447 (N_23447,N_20207,N_19980);
or U23448 (N_23448,N_19571,N_20711);
or U23449 (N_23449,N_19114,N_19059);
or U23450 (N_23450,N_19886,N_21710);
nor U23451 (N_23451,N_20572,N_19187);
and U23452 (N_23452,N_19961,N_19552);
nor U23453 (N_23453,N_21207,N_21438);
nor U23454 (N_23454,N_21243,N_18992);
nand U23455 (N_23455,N_21626,N_19697);
and U23456 (N_23456,N_21392,N_21668);
nand U23457 (N_23457,N_20862,N_21490);
or U23458 (N_23458,N_18774,N_19466);
nand U23459 (N_23459,N_20922,N_21660);
nor U23460 (N_23460,N_21768,N_21323);
or U23461 (N_23461,N_18944,N_19490);
and U23462 (N_23462,N_20481,N_21037);
or U23463 (N_23463,N_21703,N_18988);
and U23464 (N_23464,N_19588,N_19124);
nor U23465 (N_23465,N_19089,N_21114);
and U23466 (N_23466,N_21697,N_20105);
or U23467 (N_23467,N_19093,N_21792);
nand U23468 (N_23468,N_20807,N_20901);
or U23469 (N_23469,N_19937,N_19159);
and U23470 (N_23470,N_20599,N_19991);
or U23471 (N_23471,N_19901,N_19309);
or U23472 (N_23472,N_20069,N_20757);
and U23473 (N_23473,N_21555,N_20619);
or U23474 (N_23474,N_19113,N_21189);
and U23475 (N_23475,N_19572,N_19157);
or U23476 (N_23476,N_19889,N_20033);
nor U23477 (N_23477,N_19628,N_19094);
nand U23478 (N_23478,N_19171,N_19705);
nor U23479 (N_23479,N_20327,N_20864);
nand U23480 (N_23480,N_20086,N_19197);
xnor U23481 (N_23481,N_21767,N_19642);
and U23482 (N_23482,N_19606,N_20416);
or U23483 (N_23483,N_21783,N_19343);
nand U23484 (N_23484,N_21508,N_19446);
and U23485 (N_23485,N_20730,N_18770);
nor U23486 (N_23486,N_20076,N_19925);
nor U23487 (N_23487,N_20861,N_21721);
xnor U23488 (N_23488,N_19159,N_18845);
nand U23489 (N_23489,N_20683,N_20092);
nand U23490 (N_23490,N_20367,N_20780);
nand U23491 (N_23491,N_19634,N_19898);
nor U23492 (N_23492,N_21650,N_20629);
or U23493 (N_23493,N_20513,N_19724);
or U23494 (N_23494,N_20636,N_19344);
or U23495 (N_23495,N_21535,N_18934);
or U23496 (N_23496,N_19050,N_21358);
nor U23497 (N_23497,N_19028,N_19099);
nor U23498 (N_23498,N_18862,N_21386);
nor U23499 (N_23499,N_20908,N_20022);
nand U23500 (N_23500,N_19012,N_18865);
nor U23501 (N_23501,N_21352,N_20356);
nor U23502 (N_23502,N_19247,N_19915);
nand U23503 (N_23503,N_20321,N_19169);
or U23504 (N_23504,N_20748,N_19169);
and U23505 (N_23505,N_20210,N_19131);
nand U23506 (N_23506,N_19714,N_20849);
and U23507 (N_23507,N_20032,N_20307);
xnor U23508 (N_23508,N_20205,N_18770);
or U23509 (N_23509,N_19549,N_18809);
nand U23510 (N_23510,N_19093,N_20333);
and U23511 (N_23511,N_21704,N_21089);
xnor U23512 (N_23512,N_20486,N_20229);
nand U23513 (N_23513,N_20283,N_20590);
nand U23514 (N_23514,N_20538,N_20432);
nand U23515 (N_23515,N_18859,N_19094);
xnor U23516 (N_23516,N_20224,N_19791);
or U23517 (N_23517,N_20198,N_21241);
nor U23518 (N_23518,N_21316,N_20300);
and U23519 (N_23519,N_21169,N_19801);
and U23520 (N_23520,N_19705,N_21801);
xor U23521 (N_23521,N_20740,N_21761);
or U23522 (N_23522,N_20237,N_20253);
and U23523 (N_23523,N_19053,N_21810);
xor U23524 (N_23524,N_19187,N_19042);
nor U23525 (N_23525,N_19124,N_18861);
and U23526 (N_23526,N_18944,N_20791);
and U23527 (N_23527,N_19643,N_19855);
or U23528 (N_23528,N_19046,N_20270);
nor U23529 (N_23529,N_20654,N_20171);
nor U23530 (N_23530,N_20030,N_20197);
xnor U23531 (N_23531,N_19973,N_20195);
nand U23532 (N_23532,N_20485,N_19393);
or U23533 (N_23533,N_19343,N_20466);
and U23534 (N_23534,N_20238,N_18899);
nand U23535 (N_23535,N_19545,N_20221);
or U23536 (N_23536,N_19452,N_20968);
and U23537 (N_23537,N_19754,N_20491);
nand U23538 (N_23538,N_18891,N_20796);
nor U23539 (N_23539,N_19294,N_20853);
xor U23540 (N_23540,N_20498,N_20361);
xor U23541 (N_23541,N_20043,N_20544);
nor U23542 (N_23542,N_19632,N_19065);
nand U23543 (N_23543,N_19362,N_21483);
or U23544 (N_23544,N_20239,N_21119);
nand U23545 (N_23545,N_19513,N_19225);
and U23546 (N_23546,N_19355,N_19644);
nor U23547 (N_23547,N_18844,N_20586);
nand U23548 (N_23548,N_18782,N_19984);
nand U23549 (N_23549,N_20945,N_21024);
nand U23550 (N_23550,N_20717,N_19789);
or U23551 (N_23551,N_19389,N_20732);
nor U23552 (N_23552,N_19880,N_20073);
nor U23553 (N_23553,N_19555,N_19706);
or U23554 (N_23554,N_18797,N_20991);
nand U23555 (N_23555,N_19949,N_19694);
nand U23556 (N_23556,N_21865,N_20060);
or U23557 (N_23557,N_19749,N_20338);
and U23558 (N_23558,N_19991,N_19044);
and U23559 (N_23559,N_19258,N_19907);
nor U23560 (N_23560,N_19499,N_20338);
or U23561 (N_23561,N_20932,N_20594);
nor U23562 (N_23562,N_19572,N_19837);
nor U23563 (N_23563,N_21020,N_21151);
and U23564 (N_23564,N_20969,N_20533);
or U23565 (N_23565,N_18916,N_20565);
xor U23566 (N_23566,N_21455,N_19267);
or U23567 (N_23567,N_18997,N_20559);
xnor U23568 (N_23568,N_21263,N_20465);
nor U23569 (N_23569,N_19867,N_18764);
nor U23570 (N_23570,N_20553,N_19099);
nand U23571 (N_23571,N_19590,N_19906);
nor U23572 (N_23572,N_19025,N_18751);
nand U23573 (N_23573,N_21644,N_21508);
nor U23574 (N_23574,N_20659,N_20453);
xor U23575 (N_23575,N_20497,N_19210);
or U23576 (N_23576,N_20401,N_19170);
nor U23577 (N_23577,N_19176,N_19054);
and U23578 (N_23578,N_19118,N_20031);
nand U23579 (N_23579,N_20256,N_18970);
and U23580 (N_23580,N_20362,N_19811);
nor U23581 (N_23581,N_18995,N_19641);
nor U23582 (N_23582,N_21599,N_20362);
and U23583 (N_23583,N_19573,N_21523);
nor U23584 (N_23584,N_20706,N_21042);
nand U23585 (N_23585,N_18857,N_19759);
or U23586 (N_23586,N_19083,N_20112);
nor U23587 (N_23587,N_20508,N_19283);
or U23588 (N_23588,N_19720,N_21275);
or U23589 (N_23589,N_18861,N_18808);
nand U23590 (N_23590,N_20406,N_20521);
nor U23591 (N_23591,N_21064,N_20977);
or U23592 (N_23592,N_21750,N_19101);
nand U23593 (N_23593,N_18825,N_20945);
nand U23594 (N_23594,N_20412,N_18792);
nor U23595 (N_23595,N_19733,N_20490);
nor U23596 (N_23596,N_21790,N_20077);
xnor U23597 (N_23597,N_21409,N_20709);
nor U23598 (N_23598,N_18776,N_20447);
and U23599 (N_23599,N_20254,N_21624);
and U23600 (N_23600,N_20150,N_20886);
and U23601 (N_23601,N_20680,N_20803);
nor U23602 (N_23602,N_19489,N_21075);
nor U23603 (N_23603,N_19922,N_21512);
xor U23604 (N_23604,N_19698,N_21519);
xor U23605 (N_23605,N_18919,N_19839);
and U23606 (N_23606,N_20263,N_20294);
and U23607 (N_23607,N_21431,N_20129);
and U23608 (N_23608,N_20702,N_20612);
or U23609 (N_23609,N_20035,N_19431);
nor U23610 (N_23610,N_21673,N_21642);
or U23611 (N_23611,N_21704,N_21098);
or U23612 (N_23612,N_20406,N_20335);
nand U23613 (N_23613,N_20059,N_19586);
nand U23614 (N_23614,N_19454,N_20002);
nand U23615 (N_23615,N_19837,N_19110);
nor U23616 (N_23616,N_21347,N_20498);
nand U23617 (N_23617,N_19932,N_21618);
nor U23618 (N_23618,N_19037,N_21676);
or U23619 (N_23619,N_19850,N_20473);
xor U23620 (N_23620,N_20625,N_21576);
nand U23621 (N_23621,N_21420,N_20080);
or U23622 (N_23622,N_20947,N_20270);
xnor U23623 (N_23623,N_19135,N_19399);
or U23624 (N_23624,N_18754,N_20062);
and U23625 (N_23625,N_21265,N_21424);
nand U23626 (N_23626,N_20443,N_19992);
nor U23627 (N_23627,N_19431,N_19942);
nand U23628 (N_23628,N_21330,N_21413);
nor U23629 (N_23629,N_20312,N_19654);
and U23630 (N_23630,N_20380,N_19227);
nand U23631 (N_23631,N_19400,N_18933);
and U23632 (N_23632,N_21718,N_19937);
nor U23633 (N_23633,N_21693,N_20623);
or U23634 (N_23634,N_20231,N_20596);
and U23635 (N_23635,N_21469,N_20329);
and U23636 (N_23636,N_19673,N_19389);
xor U23637 (N_23637,N_19119,N_20080);
and U23638 (N_23638,N_20524,N_18820);
and U23639 (N_23639,N_19498,N_18933);
xor U23640 (N_23640,N_19407,N_21105);
or U23641 (N_23641,N_20005,N_19434);
xor U23642 (N_23642,N_19168,N_21021);
nand U23643 (N_23643,N_21701,N_18865);
nor U23644 (N_23644,N_19701,N_20642);
nand U23645 (N_23645,N_21686,N_20357);
nor U23646 (N_23646,N_19886,N_21634);
xor U23647 (N_23647,N_21836,N_20153);
and U23648 (N_23648,N_21644,N_19630);
nand U23649 (N_23649,N_18765,N_21028);
nand U23650 (N_23650,N_19500,N_20076);
or U23651 (N_23651,N_20891,N_21821);
and U23652 (N_23652,N_21710,N_18985);
xnor U23653 (N_23653,N_19473,N_21763);
nor U23654 (N_23654,N_21602,N_19378);
nand U23655 (N_23655,N_19067,N_20423);
nand U23656 (N_23656,N_19823,N_19793);
nor U23657 (N_23657,N_19971,N_21726);
or U23658 (N_23658,N_19655,N_19580);
nand U23659 (N_23659,N_20320,N_18886);
nor U23660 (N_23660,N_19387,N_19102);
xnor U23661 (N_23661,N_21163,N_20090);
or U23662 (N_23662,N_20577,N_18775);
or U23663 (N_23663,N_19580,N_21182);
nand U23664 (N_23664,N_19193,N_20700);
nand U23665 (N_23665,N_18944,N_19793);
and U23666 (N_23666,N_20324,N_19229);
or U23667 (N_23667,N_19256,N_21307);
or U23668 (N_23668,N_20742,N_21124);
nand U23669 (N_23669,N_20087,N_20697);
and U23670 (N_23670,N_20840,N_21111);
or U23671 (N_23671,N_20878,N_20234);
nor U23672 (N_23672,N_19553,N_21505);
or U23673 (N_23673,N_19328,N_18751);
nand U23674 (N_23674,N_21791,N_19547);
and U23675 (N_23675,N_20280,N_19329);
nand U23676 (N_23676,N_20539,N_19393);
nand U23677 (N_23677,N_21014,N_18811);
nand U23678 (N_23678,N_20718,N_21063);
and U23679 (N_23679,N_20395,N_21366);
nor U23680 (N_23680,N_19656,N_21466);
or U23681 (N_23681,N_20606,N_21184);
or U23682 (N_23682,N_19636,N_19456);
nor U23683 (N_23683,N_18819,N_19743);
and U23684 (N_23684,N_20008,N_20348);
or U23685 (N_23685,N_18923,N_19885);
and U23686 (N_23686,N_18795,N_20757);
and U23687 (N_23687,N_20495,N_21269);
xor U23688 (N_23688,N_21066,N_21136);
xor U23689 (N_23689,N_18829,N_19208);
or U23690 (N_23690,N_19872,N_20289);
nand U23691 (N_23691,N_20157,N_18900);
nand U23692 (N_23692,N_19444,N_21113);
or U23693 (N_23693,N_19235,N_20424);
nand U23694 (N_23694,N_19434,N_19863);
nand U23695 (N_23695,N_20288,N_19411);
nor U23696 (N_23696,N_20251,N_19736);
nand U23697 (N_23697,N_20068,N_21538);
nand U23698 (N_23698,N_21794,N_20731);
nand U23699 (N_23699,N_21072,N_19676);
and U23700 (N_23700,N_19670,N_19279);
or U23701 (N_23701,N_21312,N_19737);
or U23702 (N_23702,N_20858,N_18963);
nor U23703 (N_23703,N_20828,N_20183);
and U23704 (N_23704,N_21267,N_21793);
nor U23705 (N_23705,N_20936,N_21388);
nand U23706 (N_23706,N_20769,N_19352);
nor U23707 (N_23707,N_20107,N_19879);
nor U23708 (N_23708,N_19293,N_19197);
nand U23709 (N_23709,N_20184,N_19638);
nor U23710 (N_23710,N_20840,N_20874);
or U23711 (N_23711,N_19066,N_20177);
nor U23712 (N_23712,N_21732,N_21425);
xor U23713 (N_23713,N_20024,N_19383);
or U23714 (N_23714,N_21421,N_20222);
xor U23715 (N_23715,N_20727,N_20579);
and U23716 (N_23716,N_19049,N_19981);
nor U23717 (N_23717,N_19980,N_21062);
and U23718 (N_23718,N_20523,N_20804);
or U23719 (N_23719,N_19314,N_21355);
and U23720 (N_23720,N_18975,N_19500);
nand U23721 (N_23721,N_21423,N_18886);
and U23722 (N_23722,N_20234,N_19095);
nor U23723 (N_23723,N_20453,N_20132);
or U23724 (N_23724,N_21581,N_19209);
nor U23725 (N_23725,N_18822,N_21243);
nand U23726 (N_23726,N_21221,N_21763);
nor U23727 (N_23727,N_21784,N_21291);
xnor U23728 (N_23728,N_21239,N_19500);
and U23729 (N_23729,N_21467,N_20358);
and U23730 (N_23730,N_21724,N_19540);
nor U23731 (N_23731,N_21374,N_21227);
and U23732 (N_23732,N_21871,N_21596);
nor U23733 (N_23733,N_20781,N_20280);
or U23734 (N_23734,N_21447,N_20745);
nand U23735 (N_23735,N_18827,N_20873);
nor U23736 (N_23736,N_19144,N_19612);
nand U23737 (N_23737,N_21058,N_19230);
or U23738 (N_23738,N_19537,N_19605);
nand U23739 (N_23739,N_19406,N_18835);
nor U23740 (N_23740,N_21416,N_21003);
xnor U23741 (N_23741,N_20365,N_20022);
nand U23742 (N_23742,N_21379,N_19477);
nor U23743 (N_23743,N_21396,N_21840);
xor U23744 (N_23744,N_19882,N_21298);
nor U23745 (N_23745,N_19767,N_19148);
nor U23746 (N_23746,N_21075,N_20031);
and U23747 (N_23747,N_21065,N_19836);
xnor U23748 (N_23748,N_20299,N_20017);
nand U23749 (N_23749,N_21538,N_19928);
nor U23750 (N_23750,N_20753,N_20274);
nor U23751 (N_23751,N_19913,N_20345);
and U23752 (N_23752,N_19254,N_20706);
and U23753 (N_23753,N_18920,N_20172);
xnor U23754 (N_23754,N_20882,N_20890);
nor U23755 (N_23755,N_19636,N_19068);
or U23756 (N_23756,N_18816,N_21412);
and U23757 (N_23757,N_20720,N_19830);
nor U23758 (N_23758,N_21554,N_20374);
and U23759 (N_23759,N_19510,N_20841);
or U23760 (N_23760,N_19750,N_19051);
or U23761 (N_23761,N_20458,N_20718);
nand U23762 (N_23762,N_19750,N_19067);
nor U23763 (N_23763,N_19691,N_20980);
nor U23764 (N_23764,N_21871,N_21418);
xor U23765 (N_23765,N_20821,N_19260);
and U23766 (N_23766,N_21313,N_21484);
nor U23767 (N_23767,N_18879,N_20487);
nor U23768 (N_23768,N_21674,N_19896);
or U23769 (N_23769,N_19280,N_21871);
and U23770 (N_23770,N_19773,N_19935);
or U23771 (N_23771,N_21236,N_21862);
nand U23772 (N_23772,N_18981,N_18908);
nand U23773 (N_23773,N_21857,N_21844);
nor U23774 (N_23774,N_19558,N_19030);
nor U23775 (N_23775,N_19025,N_19277);
nand U23776 (N_23776,N_20644,N_20432);
and U23777 (N_23777,N_20427,N_18890);
xor U23778 (N_23778,N_21815,N_20977);
or U23779 (N_23779,N_19596,N_21377);
and U23780 (N_23780,N_21846,N_20877);
and U23781 (N_23781,N_18782,N_19171);
xor U23782 (N_23782,N_21854,N_21161);
nand U23783 (N_23783,N_21056,N_20429);
nor U23784 (N_23784,N_20399,N_19730);
xnor U23785 (N_23785,N_18959,N_21453);
nor U23786 (N_23786,N_19644,N_19288);
nor U23787 (N_23787,N_18914,N_19468);
and U23788 (N_23788,N_20804,N_19642);
nand U23789 (N_23789,N_19384,N_20218);
or U23790 (N_23790,N_20155,N_19657);
nor U23791 (N_23791,N_20505,N_18849);
or U23792 (N_23792,N_19624,N_20290);
xnor U23793 (N_23793,N_18895,N_19922);
or U23794 (N_23794,N_18804,N_20626);
nand U23795 (N_23795,N_21622,N_20302);
nor U23796 (N_23796,N_21093,N_18810);
nor U23797 (N_23797,N_20466,N_19887);
and U23798 (N_23798,N_20675,N_20231);
nor U23799 (N_23799,N_19547,N_20543);
and U23800 (N_23800,N_19731,N_20852);
nor U23801 (N_23801,N_18831,N_20728);
nand U23802 (N_23802,N_20370,N_21071);
nand U23803 (N_23803,N_20467,N_20360);
or U23804 (N_23804,N_21597,N_19012);
xor U23805 (N_23805,N_19257,N_20765);
nor U23806 (N_23806,N_19364,N_20793);
and U23807 (N_23807,N_18913,N_20830);
nand U23808 (N_23808,N_21828,N_18774);
xnor U23809 (N_23809,N_20624,N_19683);
nand U23810 (N_23810,N_18869,N_20480);
nand U23811 (N_23811,N_20485,N_21328);
xor U23812 (N_23812,N_20301,N_20340);
nor U23813 (N_23813,N_20639,N_19704);
nand U23814 (N_23814,N_18831,N_20974);
nand U23815 (N_23815,N_19467,N_19259);
and U23816 (N_23816,N_19502,N_20464);
nor U23817 (N_23817,N_21569,N_20100);
nand U23818 (N_23818,N_19176,N_20327);
or U23819 (N_23819,N_19436,N_19136);
and U23820 (N_23820,N_19472,N_19224);
nor U23821 (N_23821,N_21280,N_20482);
and U23822 (N_23822,N_19250,N_18764);
nor U23823 (N_23823,N_20765,N_21453);
nand U23824 (N_23824,N_21391,N_19845);
nand U23825 (N_23825,N_18797,N_21189);
nand U23826 (N_23826,N_20157,N_19708);
nor U23827 (N_23827,N_19652,N_18925);
nand U23828 (N_23828,N_21055,N_20075);
xnor U23829 (N_23829,N_19141,N_19061);
nor U23830 (N_23830,N_21621,N_21212);
nand U23831 (N_23831,N_19859,N_19342);
nor U23832 (N_23832,N_20681,N_20602);
nor U23833 (N_23833,N_20122,N_21626);
or U23834 (N_23834,N_21027,N_20244);
nand U23835 (N_23835,N_20114,N_21520);
nor U23836 (N_23836,N_18997,N_19711);
and U23837 (N_23837,N_18832,N_20228);
or U23838 (N_23838,N_19267,N_20184);
and U23839 (N_23839,N_20673,N_18788);
or U23840 (N_23840,N_20140,N_19236);
or U23841 (N_23841,N_20041,N_19320);
or U23842 (N_23842,N_21820,N_19503);
nand U23843 (N_23843,N_21634,N_21778);
and U23844 (N_23844,N_20844,N_18824);
or U23845 (N_23845,N_19780,N_18991);
nor U23846 (N_23846,N_19155,N_20460);
nor U23847 (N_23847,N_20522,N_20620);
or U23848 (N_23848,N_21171,N_19150);
or U23849 (N_23849,N_19361,N_19165);
xnor U23850 (N_23850,N_19584,N_21647);
or U23851 (N_23851,N_18958,N_18900);
or U23852 (N_23852,N_19470,N_18801);
and U23853 (N_23853,N_21749,N_19142);
or U23854 (N_23854,N_20031,N_19723);
nor U23855 (N_23855,N_20850,N_21016);
nor U23856 (N_23856,N_21175,N_19411);
and U23857 (N_23857,N_21380,N_19973);
and U23858 (N_23858,N_19682,N_21842);
nand U23859 (N_23859,N_19822,N_19119);
and U23860 (N_23860,N_20638,N_20291);
or U23861 (N_23861,N_21444,N_21120);
nand U23862 (N_23862,N_20684,N_20192);
nand U23863 (N_23863,N_21226,N_19303);
or U23864 (N_23864,N_20139,N_20130);
nand U23865 (N_23865,N_21284,N_19953);
or U23866 (N_23866,N_19557,N_20877);
and U23867 (N_23867,N_21697,N_21489);
and U23868 (N_23868,N_20726,N_20680);
or U23869 (N_23869,N_19316,N_20060);
or U23870 (N_23870,N_21778,N_21297);
and U23871 (N_23871,N_21563,N_20078);
nor U23872 (N_23872,N_21205,N_20196);
and U23873 (N_23873,N_20758,N_19886);
and U23874 (N_23874,N_21075,N_20231);
nor U23875 (N_23875,N_19534,N_19646);
nand U23876 (N_23876,N_20763,N_21740);
and U23877 (N_23877,N_21338,N_20817);
nor U23878 (N_23878,N_21343,N_20470);
nand U23879 (N_23879,N_19983,N_19804);
or U23880 (N_23880,N_20048,N_20569);
and U23881 (N_23881,N_21725,N_20753);
or U23882 (N_23882,N_19696,N_21570);
nor U23883 (N_23883,N_20766,N_19176);
nand U23884 (N_23884,N_20772,N_19307);
nor U23885 (N_23885,N_20276,N_19773);
and U23886 (N_23886,N_21254,N_20009);
and U23887 (N_23887,N_20286,N_19469);
nor U23888 (N_23888,N_20627,N_19018);
or U23889 (N_23889,N_21601,N_21321);
nor U23890 (N_23890,N_20997,N_20390);
nand U23891 (N_23891,N_21096,N_19606);
or U23892 (N_23892,N_20020,N_20154);
and U23893 (N_23893,N_19229,N_20577);
and U23894 (N_23894,N_19636,N_21868);
nand U23895 (N_23895,N_18987,N_20793);
nand U23896 (N_23896,N_21639,N_20890);
or U23897 (N_23897,N_18934,N_19238);
nor U23898 (N_23898,N_19321,N_20392);
or U23899 (N_23899,N_19113,N_19029);
or U23900 (N_23900,N_18876,N_20171);
or U23901 (N_23901,N_18817,N_21184);
or U23902 (N_23902,N_20303,N_21398);
or U23903 (N_23903,N_20303,N_21103);
nand U23904 (N_23904,N_19576,N_20838);
or U23905 (N_23905,N_18870,N_20034);
nand U23906 (N_23906,N_20196,N_19385);
nand U23907 (N_23907,N_19884,N_21133);
nand U23908 (N_23908,N_21121,N_21741);
nand U23909 (N_23909,N_21681,N_20536);
nand U23910 (N_23910,N_21300,N_20694);
nor U23911 (N_23911,N_20423,N_18751);
nand U23912 (N_23912,N_21273,N_20170);
xor U23913 (N_23913,N_20895,N_19680);
and U23914 (N_23914,N_21357,N_19620);
and U23915 (N_23915,N_19247,N_19425);
or U23916 (N_23916,N_21611,N_21063);
nor U23917 (N_23917,N_19614,N_19939);
and U23918 (N_23918,N_21343,N_21184);
xor U23919 (N_23919,N_19429,N_20018);
or U23920 (N_23920,N_20384,N_21236);
and U23921 (N_23921,N_19294,N_21767);
and U23922 (N_23922,N_20442,N_20446);
and U23923 (N_23923,N_18895,N_21298);
nand U23924 (N_23924,N_19628,N_20470);
and U23925 (N_23925,N_20895,N_19556);
nand U23926 (N_23926,N_20196,N_19877);
or U23927 (N_23927,N_21129,N_21303);
and U23928 (N_23928,N_19249,N_20240);
nand U23929 (N_23929,N_20740,N_20873);
nand U23930 (N_23930,N_19394,N_19112);
and U23931 (N_23931,N_20815,N_19389);
nor U23932 (N_23932,N_20788,N_20234);
nor U23933 (N_23933,N_19079,N_20653);
and U23934 (N_23934,N_19666,N_20578);
nand U23935 (N_23935,N_20121,N_19635);
nand U23936 (N_23936,N_19495,N_18779);
nor U23937 (N_23937,N_21654,N_18768);
and U23938 (N_23938,N_19830,N_19211);
xnor U23939 (N_23939,N_21004,N_19639);
and U23940 (N_23940,N_20300,N_18838);
and U23941 (N_23941,N_21651,N_19356);
and U23942 (N_23942,N_20551,N_19410);
and U23943 (N_23943,N_20984,N_21250);
nor U23944 (N_23944,N_20100,N_18986);
and U23945 (N_23945,N_20005,N_20890);
nand U23946 (N_23946,N_19916,N_20788);
and U23947 (N_23947,N_19275,N_21070);
or U23948 (N_23948,N_21288,N_21729);
nand U23949 (N_23949,N_19225,N_19171);
nand U23950 (N_23950,N_21325,N_21768);
nor U23951 (N_23951,N_21460,N_19811);
nor U23952 (N_23952,N_19999,N_19417);
or U23953 (N_23953,N_19181,N_21422);
nor U23954 (N_23954,N_21447,N_20164);
nor U23955 (N_23955,N_20745,N_20707);
nand U23956 (N_23956,N_21036,N_19957);
nor U23957 (N_23957,N_19594,N_21083);
or U23958 (N_23958,N_19380,N_20096);
xor U23959 (N_23959,N_21776,N_19638);
nand U23960 (N_23960,N_19834,N_19392);
nand U23961 (N_23961,N_20589,N_21173);
and U23962 (N_23962,N_21751,N_20815);
and U23963 (N_23963,N_20876,N_20774);
nor U23964 (N_23964,N_19933,N_20126);
nand U23965 (N_23965,N_21719,N_19647);
xnor U23966 (N_23966,N_20973,N_21357);
or U23967 (N_23967,N_19957,N_19435);
nor U23968 (N_23968,N_19799,N_19165);
nand U23969 (N_23969,N_20666,N_20165);
nor U23970 (N_23970,N_20784,N_21188);
nand U23971 (N_23971,N_21866,N_21635);
nor U23972 (N_23972,N_20675,N_18813);
nand U23973 (N_23973,N_20346,N_21874);
nor U23974 (N_23974,N_19115,N_21494);
and U23975 (N_23975,N_19187,N_19517);
and U23976 (N_23976,N_19262,N_19335);
nand U23977 (N_23977,N_20421,N_20863);
xnor U23978 (N_23978,N_20011,N_19530);
or U23979 (N_23979,N_20539,N_20054);
xnor U23980 (N_23980,N_19680,N_19191);
xnor U23981 (N_23981,N_21123,N_18769);
nor U23982 (N_23982,N_20609,N_18873);
nand U23983 (N_23983,N_19867,N_19213);
nand U23984 (N_23984,N_20268,N_21394);
nand U23985 (N_23985,N_19831,N_18789);
xor U23986 (N_23986,N_21461,N_19357);
nand U23987 (N_23987,N_21052,N_20684);
nand U23988 (N_23988,N_19105,N_21713);
or U23989 (N_23989,N_20755,N_19281);
xor U23990 (N_23990,N_20421,N_20518);
nor U23991 (N_23991,N_20090,N_21208);
nand U23992 (N_23992,N_21407,N_19177);
or U23993 (N_23993,N_21462,N_20362);
and U23994 (N_23994,N_18928,N_21026);
nand U23995 (N_23995,N_20412,N_19146);
nor U23996 (N_23996,N_19601,N_21111);
nand U23997 (N_23997,N_21538,N_20686);
nor U23998 (N_23998,N_21459,N_19662);
xnor U23999 (N_23999,N_19978,N_20489);
and U24000 (N_24000,N_20511,N_20590);
and U24001 (N_24001,N_19995,N_20020);
xor U24002 (N_24002,N_21104,N_19098);
nand U24003 (N_24003,N_21600,N_20596);
and U24004 (N_24004,N_19073,N_19200);
and U24005 (N_24005,N_21867,N_19926);
nor U24006 (N_24006,N_21127,N_19630);
or U24007 (N_24007,N_19870,N_19230);
xor U24008 (N_24008,N_20128,N_20635);
nand U24009 (N_24009,N_19820,N_20797);
nor U24010 (N_24010,N_20467,N_19770);
nand U24011 (N_24011,N_20805,N_21029);
and U24012 (N_24012,N_21793,N_19868);
or U24013 (N_24013,N_19482,N_19910);
nor U24014 (N_24014,N_21572,N_20917);
and U24015 (N_24015,N_20191,N_21515);
nor U24016 (N_24016,N_21656,N_21548);
and U24017 (N_24017,N_20882,N_21270);
nand U24018 (N_24018,N_20017,N_19963);
nand U24019 (N_24019,N_21203,N_19239);
nand U24020 (N_24020,N_21222,N_19703);
or U24021 (N_24021,N_18779,N_20585);
xnor U24022 (N_24022,N_18765,N_21128);
nand U24023 (N_24023,N_21712,N_18836);
and U24024 (N_24024,N_21690,N_20286);
or U24025 (N_24025,N_19785,N_20531);
nor U24026 (N_24026,N_20762,N_18830);
nand U24027 (N_24027,N_18756,N_20037);
nor U24028 (N_24028,N_21616,N_21871);
and U24029 (N_24029,N_19271,N_21612);
or U24030 (N_24030,N_19834,N_19218);
nor U24031 (N_24031,N_19856,N_21315);
or U24032 (N_24032,N_19014,N_19358);
nor U24033 (N_24033,N_19089,N_20802);
nor U24034 (N_24034,N_21735,N_19722);
and U24035 (N_24035,N_20812,N_21675);
or U24036 (N_24036,N_19292,N_21419);
nor U24037 (N_24037,N_19522,N_21522);
nor U24038 (N_24038,N_21409,N_18857);
nor U24039 (N_24039,N_20132,N_18815);
and U24040 (N_24040,N_20209,N_20773);
and U24041 (N_24041,N_21296,N_21860);
nand U24042 (N_24042,N_20214,N_19702);
nand U24043 (N_24043,N_20011,N_20686);
nand U24044 (N_24044,N_20327,N_20754);
nor U24045 (N_24045,N_19873,N_20288);
and U24046 (N_24046,N_21431,N_21293);
xor U24047 (N_24047,N_18871,N_19877);
and U24048 (N_24048,N_20906,N_19095);
or U24049 (N_24049,N_18895,N_21061);
or U24050 (N_24050,N_20098,N_19646);
nand U24051 (N_24051,N_21315,N_21564);
nand U24052 (N_24052,N_19171,N_21488);
nor U24053 (N_24053,N_19662,N_19219);
or U24054 (N_24054,N_19491,N_19960);
nor U24055 (N_24055,N_19560,N_19172);
and U24056 (N_24056,N_20376,N_21354);
nor U24057 (N_24057,N_19850,N_20884);
nand U24058 (N_24058,N_20349,N_21220);
and U24059 (N_24059,N_19721,N_20845);
and U24060 (N_24060,N_20723,N_19249);
xnor U24061 (N_24061,N_18846,N_21780);
nor U24062 (N_24062,N_19577,N_21667);
or U24063 (N_24063,N_18962,N_20209);
or U24064 (N_24064,N_20173,N_20133);
and U24065 (N_24065,N_19239,N_21273);
nor U24066 (N_24066,N_19070,N_21593);
and U24067 (N_24067,N_20719,N_19544);
and U24068 (N_24068,N_18796,N_20879);
nand U24069 (N_24069,N_20714,N_21581);
nor U24070 (N_24070,N_20317,N_21730);
or U24071 (N_24071,N_19431,N_19820);
or U24072 (N_24072,N_21684,N_21011);
and U24073 (N_24073,N_18970,N_19853);
and U24074 (N_24074,N_20358,N_21623);
nand U24075 (N_24075,N_19009,N_19542);
or U24076 (N_24076,N_21802,N_21832);
or U24077 (N_24077,N_20535,N_20710);
or U24078 (N_24078,N_21751,N_20260);
nor U24079 (N_24079,N_20239,N_18837);
nor U24080 (N_24080,N_20340,N_19635);
xor U24081 (N_24081,N_20658,N_21670);
and U24082 (N_24082,N_19979,N_21000);
nor U24083 (N_24083,N_21783,N_21102);
nor U24084 (N_24084,N_18937,N_21470);
and U24085 (N_24085,N_20575,N_21232);
nand U24086 (N_24086,N_19020,N_21420);
xnor U24087 (N_24087,N_21591,N_20580);
xor U24088 (N_24088,N_20489,N_19986);
or U24089 (N_24089,N_20705,N_20288);
or U24090 (N_24090,N_18900,N_19560);
or U24091 (N_24091,N_21632,N_20195);
or U24092 (N_24092,N_20638,N_20931);
and U24093 (N_24093,N_18931,N_20925);
or U24094 (N_24094,N_21556,N_20821);
or U24095 (N_24095,N_20651,N_21707);
or U24096 (N_24096,N_21188,N_19086);
and U24097 (N_24097,N_20825,N_19949);
and U24098 (N_24098,N_19121,N_20104);
nor U24099 (N_24099,N_18936,N_21756);
or U24100 (N_24100,N_20217,N_20980);
nand U24101 (N_24101,N_19680,N_20596);
xor U24102 (N_24102,N_20421,N_21812);
and U24103 (N_24103,N_21466,N_19466);
nor U24104 (N_24104,N_19539,N_18818);
nor U24105 (N_24105,N_21186,N_19218);
nand U24106 (N_24106,N_20381,N_20241);
nand U24107 (N_24107,N_21394,N_20778);
or U24108 (N_24108,N_19084,N_21318);
and U24109 (N_24109,N_20321,N_19704);
and U24110 (N_24110,N_19751,N_19107);
and U24111 (N_24111,N_19054,N_19788);
nand U24112 (N_24112,N_21790,N_19705);
and U24113 (N_24113,N_21031,N_19632);
nand U24114 (N_24114,N_21539,N_20384);
nand U24115 (N_24115,N_21480,N_19951);
and U24116 (N_24116,N_20133,N_20513);
or U24117 (N_24117,N_19689,N_20894);
and U24118 (N_24118,N_19699,N_20771);
nand U24119 (N_24119,N_21350,N_21591);
nand U24120 (N_24120,N_21224,N_19104);
nor U24121 (N_24121,N_20819,N_20017);
and U24122 (N_24122,N_20808,N_19472);
xnor U24123 (N_24123,N_21187,N_19302);
and U24124 (N_24124,N_20059,N_20570);
and U24125 (N_24125,N_20086,N_19607);
nand U24126 (N_24126,N_21669,N_21210);
xnor U24127 (N_24127,N_19418,N_20549);
and U24128 (N_24128,N_20805,N_20344);
and U24129 (N_24129,N_18824,N_20202);
nand U24130 (N_24130,N_19700,N_20144);
nor U24131 (N_24131,N_21181,N_18813);
and U24132 (N_24132,N_20956,N_19447);
nor U24133 (N_24133,N_18934,N_20813);
nand U24134 (N_24134,N_19063,N_20371);
xor U24135 (N_24135,N_19626,N_18940);
nand U24136 (N_24136,N_20726,N_20019);
nand U24137 (N_24137,N_21066,N_21323);
or U24138 (N_24138,N_19016,N_20117);
nor U24139 (N_24139,N_20303,N_19225);
nor U24140 (N_24140,N_18770,N_21718);
or U24141 (N_24141,N_18756,N_20135);
nor U24142 (N_24142,N_20220,N_21158);
or U24143 (N_24143,N_19468,N_21628);
or U24144 (N_24144,N_21154,N_21127);
and U24145 (N_24145,N_20749,N_18888);
and U24146 (N_24146,N_19646,N_20885);
nor U24147 (N_24147,N_20879,N_21040);
nor U24148 (N_24148,N_20796,N_20670);
or U24149 (N_24149,N_19298,N_19562);
and U24150 (N_24150,N_21199,N_21214);
and U24151 (N_24151,N_20134,N_20868);
and U24152 (N_24152,N_21501,N_18935);
and U24153 (N_24153,N_18986,N_19322);
nor U24154 (N_24154,N_21796,N_20955);
and U24155 (N_24155,N_20903,N_19332);
xor U24156 (N_24156,N_19169,N_21508);
and U24157 (N_24157,N_19519,N_21494);
nand U24158 (N_24158,N_21501,N_21656);
or U24159 (N_24159,N_21859,N_21558);
xnor U24160 (N_24160,N_19980,N_21095);
xor U24161 (N_24161,N_19563,N_20322);
or U24162 (N_24162,N_19489,N_19463);
or U24163 (N_24163,N_18968,N_21315);
nand U24164 (N_24164,N_20325,N_19078);
nand U24165 (N_24165,N_21025,N_20247);
or U24166 (N_24166,N_21689,N_19303);
nand U24167 (N_24167,N_19250,N_19439);
or U24168 (N_24168,N_19999,N_19983);
nand U24169 (N_24169,N_19423,N_18763);
and U24170 (N_24170,N_18750,N_20502);
nand U24171 (N_24171,N_19335,N_20897);
nor U24172 (N_24172,N_20909,N_19118);
nor U24173 (N_24173,N_19024,N_21547);
nand U24174 (N_24174,N_21584,N_21373);
and U24175 (N_24175,N_20873,N_19867);
nand U24176 (N_24176,N_20015,N_21674);
nand U24177 (N_24177,N_20556,N_21172);
or U24178 (N_24178,N_21373,N_20358);
and U24179 (N_24179,N_19632,N_20987);
and U24180 (N_24180,N_20865,N_19389);
and U24181 (N_24181,N_18840,N_21852);
nand U24182 (N_24182,N_20598,N_19869);
and U24183 (N_24183,N_20858,N_21445);
and U24184 (N_24184,N_18936,N_19826);
nor U24185 (N_24185,N_19915,N_20601);
or U24186 (N_24186,N_20070,N_20346);
nand U24187 (N_24187,N_20226,N_21704);
nor U24188 (N_24188,N_20370,N_19146);
nor U24189 (N_24189,N_20337,N_19494);
xnor U24190 (N_24190,N_19372,N_18767);
nand U24191 (N_24191,N_20485,N_21547);
xor U24192 (N_24192,N_19116,N_21492);
nand U24193 (N_24193,N_18828,N_21163);
or U24194 (N_24194,N_21862,N_19938);
or U24195 (N_24195,N_18814,N_21398);
and U24196 (N_24196,N_19786,N_21464);
nand U24197 (N_24197,N_19531,N_20578);
or U24198 (N_24198,N_19917,N_20902);
or U24199 (N_24199,N_21437,N_20489);
nor U24200 (N_24200,N_20609,N_18811);
and U24201 (N_24201,N_20953,N_20932);
nand U24202 (N_24202,N_20837,N_21225);
nor U24203 (N_24203,N_20739,N_18929);
nand U24204 (N_24204,N_19890,N_19369);
nand U24205 (N_24205,N_20524,N_21748);
or U24206 (N_24206,N_21562,N_19580);
nand U24207 (N_24207,N_20672,N_20391);
and U24208 (N_24208,N_19078,N_19411);
and U24209 (N_24209,N_20938,N_21726);
nand U24210 (N_24210,N_19028,N_21715);
and U24211 (N_24211,N_20277,N_20125);
nand U24212 (N_24212,N_20438,N_21763);
and U24213 (N_24213,N_20975,N_18836);
xnor U24214 (N_24214,N_20421,N_20894);
nor U24215 (N_24215,N_18955,N_18987);
or U24216 (N_24216,N_19327,N_21837);
xor U24217 (N_24217,N_21667,N_19455);
nand U24218 (N_24218,N_20868,N_20157);
nand U24219 (N_24219,N_20867,N_20742);
nand U24220 (N_24220,N_19298,N_20255);
and U24221 (N_24221,N_19313,N_18828);
and U24222 (N_24222,N_20429,N_19774);
or U24223 (N_24223,N_21310,N_21712);
and U24224 (N_24224,N_20918,N_20214);
and U24225 (N_24225,N_19558,N_20844);
and U24226 (N_24226,N_20640,N_21590);
or U24227 (N_24227,N_21554,N_19595);
and U24228 (N_24228,N_18892,N_19092);
or U24229 (N_24229,N_20102,N_20809);
or U24230 (N_24230,N_20978,N_21311);
or U24231 (N_24231,N_18788,N_20511);
and U24232 (N_24232,N_21699,N_19422);
nand U24233 (N_24233,N_20126,N_19128);
and U24234 (N_24234,N_20605,N_19875);
and U24235 (N_24235,N_19552,N_20436);
and U24236 (N_24236,N_19666,N_21590);
or U24237 (N_24237,N_19735,N_21472);
nand U24238 (N_24238,N_21393,N_19583);
and U24239 (N_24239,N_21014,N_21231);
nor U24240 (N_24240,N_18967,N_19537);
nor U24241 (N_24241,N_21097,N_20953);
nand U24242 (N_24242,N_19778,N_19747);
and U24243 (N_24243,N_20563,N_20253);
nand U24244 (N_24244,N_20619,N_20289);
nor U24245 (N_24245,N_20857,N_20543);
or U24246 (N_24246,N_19352,N_21352);
and U24247 (N_24247,N_20834,N_19229);
xnor U24248 (N_24248,N_18778,N_19007);
or U24249 (N_24249,N_20183,N_20097);
xnor U24250 (N_24250,N_19697,N_20997);
or U24251 (N_24251,N_19988,N_18827);
or U24252 (N_24252,N_21328,N_20381);
and U24253 (N_24253,N_21411,N_20371);
or U24254 (N_24254,N_21625,N_19627);
nand U24255 (N_24255,N_19197,N_19616);
nand U24256 (N_24256,N_21011,N_20260);
nor U24257 (N_24257,N_19663,N_20252);
and U24258 (N_24258,N_21657,N_18843);
nor U24259 (N_24259,N_20839,N_20947);
xor U24260 (N_24260,N_21267,N_19046);
or U24261 (N_24261,N_20784,N_19767);
or U24262 (N_24262,N_21026,N_21040);
or U24263 (N_24263,N_19251,N_20660);
nand U24264 (N_24264,N_19497,N_20118);
nor U24265 (N_24265,N_19467,N_21851);
xnor U24266 (N_24266,N_19390,N_18804);
or U24267 (N_24267,N_21538,N_21574);
nand U24268 (N_24268,N_20005,N_20881);
nor U24269 (N_24269,N_21366,N_20618);
nor U24270 (N_24270,N_21101,N_20037);
nand U24271 (N_24271,N_20960,N_19674);
nand U24272 (N_24272,N_21135,N_21686);
and U24273 (N_24273,N_18815,N_20281);
or U24274 (N_24274,N_20318,N_21187);
and U24275 (N_24275,N_20954,N_19146);
nor U24276 (N_24276,N_20678,N_21541);
nand U24277 (N_24277,N_21266,N_21392);
and U24278 (N_24278,N_21689,N_21746);
and U24279 (N_24279,N_19312,N_19635);
or U24280 (N_24280,N_20925,N_21829);
xnor U24281 (N_24281,N_20042,N_19006);
nor U24282 (N_24282,N_19923,N_19630);
nand U24283 (N_24283,N_20232,N_19596);
and U24284 (N_24284,N_19351,N_18777);
and U24285 (N_24285,N_19830,N_21815);
and U24286 (N_24286,N_20441,N_20140);
or U24287 (N_24287,N_20073,N_20218);
or U24288 (N_24288,N_21804,N_21056);
xor U24289 (N_24289,N_20119,N_21127);
nand U24290 (N_24290,N_21402,N_20046);
nand U24291 (N_24291,N_18943,N_21030);
or U24292 (N_24292,N_20297,N_20562);
nor U24293 (N_24293,N_19734,N_20062);
xor U24294 (N_24294,N_20893,N_20325);
or U24295 (N_24295,N_20304,N_20144);
xor U24296 (N_24296,N_21301,N_20592);
nor U24297 (N_24297,N_20291,N_20233);
nor U24298 (N_24298,N_20422,N_21172);
or U24299 (N_24299,N_20552,N_19273);
nand U24300 (N_24300,N_19802,N_20337);
or U24301 (N_24301,N_21173,N_20958);
nor U24302 (N_24302,N_20055,N_20443);
nand U24303 (N_24303,N_18786,N_20145);
or U24304 (N_24304,N_20080,N_19042);
nand U24305 (N_24305,N_20401,N_18865);
and U24306 (N_24306,N_20391,N_19384);
or U24307 (N_24307,N_20715,N_21496);
nand U24308 (N_24308,N_19275,N_20114);
and U24309 (N_24309,N_19495,N_21437);
nor U24310 (N_24310,N_19527,N_20968);
or U24311 (N_24311,N_21836,N_19897);
or U24312 (N_24312,N_20974,N_20172);
nand U24313 (N_24313,N_20964,N_20777);
and U24314 (N_24314,N_20786,N_20709);
xnor U24315 (N_24315,N_18864,N_19555);
or U24316 (N_24316,N_19898,N_20032);
nor U24317 (N_24317,N_21419,N_19056);
or U24318 (N_24318,N_20359,N_20108);
or U24319 (N_24319,N_20889,N_21833);
nor U24320 (N_24320,N_21223,N_20027);
nor U24321 (N_24321,N_19382,N_20098);
and U24322 (N_24322,N_21308,N_21433);
and U24323 (N_24323,N_19086,N_20275);
nor U24324 (N_24324,N_21132,N_20776);
and U24325 (N_24325,N_20264,N_21228);
or U24326 (N_24326,N_20651,N_18868);
and U24327 (N_24327,N_21245,N_18855);
and U24328 (N_24328,N_19880,N_20268);
and U24329 (N_24329,N_20165,N_21260);
nand U24330 (N_24330,N_20363,N_21104);
nand U24331 (N_24331,N_20080,N_19970);
nor U24332 (N_24332,N_19881,N_18794);
nand U24333 (N_24333,N_20732,N_19191);
and U24334 (N_24334,N_21156,N_21761);
and U24335 (N_24335,N_19076,N_21659);
nor U24336 (N_24336,N_19508,N_21420);
or U24337 (N_24337,N_20223,N_20311);
or U24338 (N_24338,N_19413,N_20782);
or U24339 (N_24339,N_21076,N_21062);
nor U24340 (N_24340,N_19738,N_18865);
nand U24341 (N_24341,N_19625,N_20978);
or U24342 (N_24342,N_21121,N_19814);
nor U24343 (N_24343,N_20183,N_20160);
nor U24344 (N_24344,N_18791,N_21671);
and U24345 (N_24345,N_20924,N_21427);
nor U24346 (N_24346,N_19301,N_18889);
or U24347 (N_24347,N_19050,N_20437);
or U24348 (N_24348,N_18975,N_21661);
nand U24349 (N_24349,N_20813,N_19986);
nand U24350 (N_24350,N_21586,N_20496);
or U24351 (N_24351,N_18762,N_21780);
and U24352 (N_24352,N_19441,N_19363);
or U24353 (N_24353,N_19524,N_19276);
nand U24354 (N_24354,N_20711,N_19778);
nand U24355 (N_24355,N_19243,N_21205);
or U24356 (N_24356,N_19395,N_18846);
nor U24357 (N_24357,N_19876,N_20994);
or U24358 (N_24358,N_19430,N_21555);
or U24359 (N_24359,N_21002,N_21599);
nor U24360 (N_24360,N_20010,N_19492);
nor U24361 (N_24361,N_19549,N_19772);
nand U24362 (N_24362,N_19446,N_21745);
and U24363 (N_24363,N_21171,N_21342);
nand U24364 (N_24364,N_19325,N_21161);
xnor U24365 (N_24365,N_21616,N_19025);
or U24366 (N_24366,N_18869,N_20975);
nand U24367 (N_24367,N_21285,N_20946);
nand U24368 (N_24368,N_19589,N_20187);
and U24369 (N_24369,N_20128,N_21598);
nand U24370 (N_24370,N_21370,N_19815);
nor U24371 (N_24371,N_21471,N_20718);
nor U24372 (N_24372,N_19195,N_21855);
or U24373 (N_24373,N_20628,N_21727);
xor U24374 (N_24374,N_21059,N_19774);
nor U24375 (N_24375,N_20907,N_19381);
nand U24376 (N_24376,N_18752,N_20386);
nand U24377 (N_24377,N_21565,N_19515);
or U24378 (N_24378,N_20145,N_18917);
xor U24379 (N_24379,N_20708,N_18986);
nor U24380 (N_24380,N_21162,N_19291);
and U24381 (N_24381,N_21656,N_21130);
nor U24382 (N_24382,N_18793,N_19426);
nor U24383 (N_24383,N_19583,N_20478);
or U24384 (N_24384,N_21180,N_21142);
or U24385 (N_24385,N_21743,N_20627);
nor U24386 (N_24386,N_21157,N_19530);
nor U24387 (N_24387,N_19095,N_19752);
or U24388 (N_24388,N_18753,N_21105);
nor U24389 (N_24389,N_18971,N_20250);
nor U24390 (N_24390,N_20817,N_21150);
or U24391 (N_24391,N_19805,N_21280);
nand U24392 (N_24392,N_20764,N_21324);
xnor U24393 (N_24393,N_20134,N_20916);
nor U24394 (N_24394,N_21677,N_19753);
nand U24395 (N_24395,N_19930,N_21145);
and U24396 (N_24396,N_19616,N_20317);
nor U24397 (N_24397,N_20784,N_21861);
and U24398 (N_24398,N_20409,N_20936);
xnor U24399 (N_24399,N_20893,N_21001);
nand U24400 (N_24400,N_20989,N_20291);
or U24401 (N_24401,N_20520,N_20025);
or U24402 (N_24402,N_20748,N_21485);
nor U24403 (N_24403,N_20117,N_19717);
nor U24404 (N_24404,N_21246,N_21824);
or U24405 (N_24405,N_20311,N_21664);
nor U24406 (N_24406,N_20381,N_21230);
xor U24407 (N_24407,N_20985,N_20237);
nor U24408 (N_24408,N_21279,N_19366);
and U24409 (N_24409,N_20446,N_20240);
nor U24410 (N_24410,N_18795,N_21748);
or U24411 (N_24411,N_19854,N_19683);
or U24412 (N_24412,N_20167,N_21038);
nor U24413 (N_24413,N_20388,N_20865);
and U24414 (N_24414,N_20747,N_19108);
nand U24415 (N_24415,N_19546,N_19573);
nor U24416 (N_24416,N_20126,N_19323);
nor U24417 (N_24417,N_20552,N_21195);
nor U24418 (N_24418,N_19379,N_21745);
and U24419 (N_24419,N_20022,N_19939);
nand U24420 (N_24420,N_19820,N_19718);
nand U24421 (N_24421,N_21700,N_20050);
nand U24422 (N_24422,N_19387,N_19314);
or U24423 (N_24423,N_19603,N_21422);
and U24424 (N_24424,N_19619,N_20929);
or U24425 (N_24425,N_21357,N_20492);
nand U24426 (N_24426,N_20683,N_19998);
nand U24427 (N_24427,N_19618,N_20827);
nand U24428 (N_24428,N_19620,N_18802);
nand U24429 (N_24429,N_19405,N_19778);
nand U24430 (N_24430,N_19370,N_19064);
nor U24431 (N_24431,N_18863,N_19564);
and U24432 (N_24432,N_20650,N_19776);
nor U24433 (N_24433,N_21027,N_20696);
nand U24434 (N_24434,N_20963,N_20337);
and U24435 (N_24435,N_20296,N_21039);
nor U24436 (N_24436,N_19616,N_21549);
and U24437 (N_24437,N_19775,N_21051);
nand U24438 (N_24438,N_21421,N_21822);
nor U24439 (N_24439,N_21076,N_19615);
nor U24440 (N_24440,N_19108,N_19967);
nand U24441 (N_24441,N_20504,N_18976);
and U24442 (N_24442,N_19922,N_19433);
nor U24443 (N_24443,N_19929,N_21694);
nand U24444 (N_24444,N_19960,N_19844);
and U24445 (N_24445,N_19515,N_21591);
nand U24446 (N_24446,N_20537,N_21091);
nor U24447 (N_24447,N_21090,N_19130);
nor U24448 (N_24448,N_20277,N_19299);
nand U24449 (N_24449,N_19865,N_21551);
or U24450 (N_24450,N_19879,N_21313);
nor U24451 (N_24451,N_19404,N_21058);
or U24452 (N_24452,N_21368,N_20097);
and U24453 (N_24453,N_21782,N_18825);
or U24454 (N_24454,N_19859,N_19242);
or U24455 (N_24455,N_20517,N_21487);
nor U24456 (N_24456,N_19155,N_19570);
nor U24457 (N_24457,N_18964,N_19232);
or U24458 (N_24458,N_19599,N_21605);
nor U24459 (N_24459,N_20345,N_21556);
and U24460 (N_24460,N_19575,N_19558);
nor U24461 (N_24461,N_19280,N_21648);
or U24462 (N_24462,N_20473,N_19747);
or U24463 (N_24463,N_21687,N_19046);
or U24464 (N_24464,N_21317,N_21435);
nor U24465 (N_24465,N_20520,N_20803);
nor U24466 (N_24466,N_18991,N_19185);
nor U24467 (N_24467,N_20922,N_19870);
and U24468 (N_24468,N_21372,N_21677);
or U24469 (N_24469,N_21335,N_18818);
nor U24470 (N_24470,N_21194,N_21105);
nand U24471 (N_24471,N_19747,N_20689);
or U24472 (N_24472,N_21320,N_21873);
or U24473 (N_24473,N_21029,N_19913);
nor U24474 (N_24474,N_19102,N_18779);
xor U24475 (N_24475,N_20020,N_21196);
or U24476 (N_24476,N_19524,N_20676);
nor U24477 (N_24477,N_19417,N_18780);
nand U24478 (N_24478,N_20057,N_20852);
or U24479 (N_24479,N_18824,N_20288);
nor U24480 (N_24480,N_19423,N_21061);
and U24481 (N_24481,N_20110,N_19439);
nand U24482 (N_24482,N_20181,N_21352);
nor U24483 (N_24483,N_20449,N_21693);
nor U24484 (N_24484,N_21053,N_19189);
and U24485 (N_24485,N_19804,N_20513);
or U24486 (N_24486,N_19448,N_20188);
nand U24487 (N_24487,N_20770,N_19673);
nand U24488 (N_24488,N_19767,N_21394);
xnor U24489 (N_24489,N_20703,N_19481);
and U24490 (N_24490,N_19000,N_19540);
xnor U24491 (N_24491,N_21797,N_19240);
nor U24492 (N_24492,N_19832,N_20103);
nand U24493 (N_24493,N_20144,N_19148);
nand U24494 (N_24494,N_18895,N_19832);
and U24495 (N_24495,N_19961,N_21618);
xnor U24496 (N_24496,N_21321,N_19951);
or U24497 (N_24497,N_19474,N_21092);
nand U24498 (N_24498,N_21571,N_20906);
nand U24499 (N_24499,N_19787,N_20377);
xor U24500 (N_24500,N_21763,N_18875);
or U24501 (N_24501,N_20188,N_20197);
or U24502 (N_24502,N_20562,N_19095);
or U24503 (N_24503,N_19931,N_20101);
nand U24504 (N_24504,N_20757,N_21220);
and U24505 (N_24505,N_21872,N_20786);
nand U24506 (N_24506,N_18975,N_21684);
nand U24507 (N_24507,N_21549,N_19469);
nand U24508 (N_24508,N_19774,N_21333);
nor U24509 (N_24509,N_21235,N_19431);
nand U24510 (N_24510,N_19704,N_20134);
and U24511 (N_24511,N_18752,N_19901);
and U24512 (N_24512,N_20984,N_20231);
nand U24513 (N_24513,N_21714,N_19239);
and U24514 (N_24514,N_19980,N_21108);
or U24515 (N_24515,N_20464,N_20628);
or U24516 (N_24516,N_18801,N_20440);
or U24517 (N_24517,N_19630,N_19786);
xor U24518 (N_24518,N_21558,N_19708);
xor U24519 (N_24519,N_20887,N_20499);
nor U24520 (N_24520,N_21542,N_19545);
nand U24521 (N_24521,N_21048,N_21130);
or U24522 (N_24522,N_20190,N_20900);
nor U24523 (N_24523,N_20338,N_20649);
nor U24524 (N_24524,N_20461,N_19207);
or U24525 (N_24525,N_18936,N_18979);
or U24526 (N_24526,N_20270,N_20526);
xnor U24527 (N_24527,N_19331,N_19691);
or U24528 (N_24528,N_20133,N_19058);
nor U24529 (N_24529,N_18825,N_19415);
nor U24530 (N_24530,N_20782,N_21611);
nor U24531 (N_24531,N_21251,N_20836);
nand U24532 (N_24532,N_20205,N_20865);
nor U24533 (N_24533,N_20497,N_21036);
xor U24534 (N_24534,N_19359,N_20572);
and U24535 (N_24535,N_20177,N_18867);
nor U24536 (N_24536,N_20619,N_21171);
or U24537 (N_24537,N_21197,N_20853);
and U24538 (N_24538,N_18999,N_21761);
nand U24539 (N_24539,N_21340,N_20649);
nand U24540 (N_24540,N_20325,N_19874);
nor U24541 (N_24541,N_19553,N_21398);
nand U24542 (N_24542,N_19527,N_21139);
nor U24543 (N_24543,N_20394,N_20371);
nand U24544 (N_24544,N_20549,N_21141);
nand U24545 (N_24545,N_20906,N_20644);
and U24546 (N_24546,N_18941,N_20743);
and U24547 (N_24547,N_19813,N_18788);
and U24548 (N_24548,N_20527,N_21490);
nand U24549 (N_24549,N_20294,N_20884);
nor U24550 (N_24550,N_19242,N_18936);
xnor U24551 (N_24551,N_21542,N_20307);
or U24552 (N_24552,N_21192,N_20356);
and U24553 (N_24553,N_20194,N_20357);
or U24554 (N_24554,N_20076,N_21790);
or U24555 (N_24555,N_20457,N_20061);
nand U24556 (N_24556,N_20043,N_19916);
nand U24557 (N_24557,N_20261,N_19498);
nand U24558 (N_24558,N_18964,N_19894);
and U24559 (N_24559,N_20512,N_19083);
and U24560 (N_24560,N_20632,N_19281);
or U24561 (N_24561,N_20698,N_19118);
nand U24562 (N_24562,N_19490,N_18867);
nor U24563 (N_24563,N_19413,N_19517);
nand U24564 (N_24564,N_21722,N_19012);
and U24565 (N_24565,N_21563,N_19102);
or U24566 (N_24566,N_20196,N_20384);
xor U24567 (N_24567,N_19530,N_19808);
and U24568 (N_24568,N_20962,N_19927);
nand U24569 (N_24569,N_18842,N_19650);
nor U24570 (N_24570,N_19407,N_21587);
and U24571 (N_24571,N_19647,N_20542);
and U24572 (N_24572,N_18967,N_21765);
nor U24573 (N_24573,N_19957,N_21116);
or U24574 (N_24574,N_21069,N_19093);
nor U24575 (N_24575,N_21519,N_21155);
or U24576 (N_24576,N_20942,N_19538);
xnor U24577 (N_24577,N_21506,N_19070);
and U24578 (N_24578,N_21243,N_21042);
or U24579 (N_24579,N_21554,N_19653);
and U24580 (N_24580,N_19733,N_19910);
nand U24581 (N_24581,N_19289,N_20311);
and U24582 (N_24582,N_19974,N_20265);
nor U24583 (N_24583,N_20320,N_19338);
nand U24584 (N_24584,N_19504,N_20440);
and U24585 (N_24585,N_19939,N_19222);
and U24586 (N_24586,N_20842,N_19495);
or U24587 (N_24587,N_20725,N_20443);
nor U24588 (N_24588,N_20465,N_20632);
nand U24589 (N_24589,N_18764,N_19528);
nand U24590 (N_24590,N_21277,N_19163);
nand U24591 (N_24591,N_18808,N_21167);
xor U24592 (N_24592,N_20735,N_20563);
xnor U24593 (N_24593,N_21461,N_19787);
nor U24594 (N_24594,N_20998,N_19331);
or U24595 (N_24595,N_19486,N_21563);
xnor U24596 (N_24596,N_20710,N_20059);
xnor U24597 (N_24597,N_20360,N_21837);
and U24598 (N_24598,N_19771,N_21203);
or U24599 (N_24599,N_18950,N_21266);
nor U24600 (N_24600,N_21011,N_20421);
nor U24601 (N_24601,N_20835,N_20885);
and U24602 (N_24602,N_20951,N_18869);
or U24603 (N_24603,N_20010,N_21794);
nor U24604 (N_24604,N_19074,N_21848);
nor U24605 (N_24605,N_21063,N_19594);
nor U24606 (N_24606,N_19793,N_20957);
and U24607 (N_24607,N_20683,N_20680);
nand U24608 (N_24608,N_21802,N_20535);
and U24609 (N_24609,N_21692,N_20424);
nand U24610 (N_24610,N_21215,N_20055);
nand U24611 (N_24611,N_21404,N_19842);
nand U24612 (N_24612,N_18979,N_20733);
and U24613 (N_24613,N_20703,N_19496);
or U24614 (N_24614,N_20629,N_19349);
nor U24615 (N_24615,N_20046,N_20058);
nor U24616 (N_24616,N_19089,N_20562);
and U24617 (N_24617,N_18976,N_20477);
nor U24618 (N_24618,N_21172,N_18856);
or U24619 (N_24619,N_19007,N_19303);
nand U24620 (N_24620,N_20034,N_19080);
nor U24621 (N_24621,N_20338,N_21745);
nand U24622 (N_24622,N_20012,N_19290);
and U24623 (N_24623,N_20819,N_21494);
nand U24624 (N_24624,N_19072,N_18953);
or U24625 (N_24625,N_19117,N_19916);
or U24626 (N_24626,N_18953,N_19037);
nand U24627 (N_24627,N_21110,N_19792);
or U24628 (N_24628,N_19068,N_21598);
xor U24629 (N_24629,N_20838,N_21757);
nor U24630 (N_24630,N_20050,N_19832);
nor U24631 (N_24631,N_21203,N_21833);
nand U24632 (N_24632,N_19462,N_21474);
nand U24633 (N_24633,N_19387,N_21737);
and U24634 (N_24634,N_20346,N_21428);
and U24635 (N_24635,N_19842,N_21545);
or U24636 (N_24636,N_20406,N_20879);
nor U24637 (N_24637,N_19223,N_21611);
nor U24638 (N_24638,N_21836,N_19055);
nand U24639 (N_24639,N_19697,N_20152);
and U24640 (N_24640,N_20570,N_20523);
and U24641 (N_24641,N_19541,N_21813);
nor U24642 (N_24642,N_21519,N_20754);
nor U24643 (N_24643,N_21458,N_21257);
xnor U24644 (N_24644,N_20032,N_20738);
nor U24645 (N_24645,N_21285,N_21092);
nor U24646 (N_24646,N_21079,N_19162);
and U24647 (N_24647,N_20323,N_20446);
nor U24648 (N_24648,N_19551,N_21720);
nand U24649 (N_24649,N_19636,N_19494);
nor U24650 (N_24650,N_18789,N_19724);
and U24651 (N_24651,N_19883,N_19094);
and U24652 (N_24652,N_21842,N_19065);
nor U24653 (N_24653,N_19779,N_20833);
nand U24654 (N_24654,N_21054,N_21416);
or U24655 (N_24655,N_21351,N_21707);
nand U24656 (N_24656,N_20897,N_20706);
and U24657 (N_24657,N_21409,N_19584);
nand U24658 (N_24658,N_18785,N_20035);
and U24659 (N_24659,N_19726,N_19021);
or U24660 (N_24660,N_21835,N_19268);
or U24661 (N_24661,N_19700,N_20172);
or U24662 (N_24662,N_19328,N_18759);
nand U24663 (N_24663,N_19366,N_21431);
or U24664 (N_24664,N_19080,N_21855);
or U24665 (N_24665,N_21086,N_21381);
xnor U24666 (N_24666,N_19919,N_19096);
nand U24667 (N_24667,N_20074,N_21595);
and U24668 (N_24668,N_21550,N_20359);
and U24669 (N_24669,N_21805,N_20168);
and U24670 (N_24670,N_19279,N_19233);
nand U24671 (N_24671,N_21721,N_21479);
xnor U24672 (N_24672,N_18957,N_20180);
or U24673 (N_24673,N_21693,N_21755);
and U24674 (N_24674,N_19521,N_21364);
nand U24675 (N_24675,N_20531,N_21217);
xnor U24676 (N_24676,N_21397,N_19182);
nand U24677 (N_24677,N_21068,N_19944);
and U24678 (N_24678,N_19911,N_21424);
nor U24679 (N_24679,N_20802,N_20132);
and U24680 (N_24680,N_19865,N_20599);
and U24681 (N_24681,N_21436,N_19366);
or U24682 (N_24682,N_21197,N_21735);
nand U24683 (N_24683,N_20445,N_21206);
nand U24684 (N_24684,N_21384,N_21189);
nor U24685 (N_24685,N_19303,N_20802);
nor U24686 (N_24686,N_19289,N_20068);
or U24687 (N_24687,N_21519,N_21689);
or U24688 (N_24688,N_19926,N_19517);
nor U24689 (N_24689,N_18957,N_20233);
nor U24690 (N_24690,N_20742,N_20786);
and U24691 (N_24691,N_21288,N_19651);
nand U24692 (N_24692,N_21330,N_21819);
or U24693 (N_24693,N_19974,N_20370);
nor U24694 (N_24694,N_21389,N_20034);
or U24695 (N_24695,N_19755,N_20569);
xor U24696 (N_24696,N_19084,N_19066);
nor U24697 (N_24697,N_19970,N_19448);
nor U24698 (N_24698,N_18982,N_19446);
and U24699 (N_24699,N_21790,N_19063);
and U24700 (N_24700,N_19519,N_20348);
nand U24701 (N_24701,N_19139,N_20422);
and U24702 (N_24702,N_19751,N_19659);
and U24703 (N_24703,N_21191,N_19051);
nor U24704 (N_24704,N_19774,N_19568);
and U24705 (N_24705,N_19191,N_18906);
or U24706 (N_24706,N_20318,N_20955);
or U24707 (N_24707,N_21183,N_19197);
or U24708 (N_24708,N_21205,N_21242);
nor U24709 (N_24709,N_20321,N_21847);
nor U24710 (N_24710,N_18776,N_19320);
nand U24711 (N_24711,N_20580,N_19265);
nor U24712 (N_24712,N_21017,N_18894);
nand U24713 (N_24713,N_20543,N_21170);
nor U24714 (N_24714,N_20607,N_19986);
nand U24715 (N_24715,N_18763,N_21745);
nor U24716 (N_24716,N_20074,N_19370);
nand U24717 (N_24717,N_20137,N_19613);
and U24718 (N_24718,N_20241,N_20742);
or U24719 (N_24719,N_20006,N_21136);
and U24720 (N_24720,N_21265,N_20746);
nor U24721 (N_24721,N_18922,N_20833);
xnor U24722 (N_24722,N_19308,N_20381);
and U24723 (N_24723,N_19848,N_20277);
nor U24724 (N_24724,N_20438,N_19994);
or U24725 (N_24725,N_21864,N_21367);
nand U24726 (N_24726,N_21458,N_20786);
nor U24727 (N_24727,N_21523,N_21283);
nand U24728 (N_24728,N_20105,N_19147);
and U24729 (N_24729,N_21025,N_19598);
nand U24730 (N_24730,N_19785,N_21675);
and U24731 (N_24731,N_19652,N_20826);
nor U24732 (N_24732,N_20587,N_21452);
or U24733 (N_24733,N_20480,N_21484);
or U24734 (N_24734,N_21039,N_20542);
and U24735 (N_24735,N_18789,N_20352);
and U24736 (N_24736,N_21336,N_19471);
and U24737 (N_24737,N_20378,N_20775);
nand U24738 (N_24738,N_19629,N_20092);
or U24739 (N_24739,N_20844,N_20309);
or U24740 (N_24740,N_19841,N_19608);
nor U24741 (N_24741,N_21556,N_19022);
nor U24742 (N_24742,N_19678,N_20921);
or U24743 (N_24743,N_21316,N_21697);
or U24744 (N_24744,N_18981,N_20527);
or U24745 (N_24745,N_21807,N_20148);
and U24746 (N_24746,N_20191,N_20769);
nor U24747 (N_24747,N_19706,N_18936);
nor U24748 (N_24748,N_19387,N_18963);
nor U24749 (N_24749,N_19441,N_18976);
or U24750 (N_24750,N_21080,N_19454);
or U24751 (N_24751,N_19358,N_20115);
and U24752 (N_24752,N_19895,N_19507);
nand U24753 (N_24753,N_19923,N_20497);
and U24754 (N_24754,N_19677,N_19163);
and U24755 (N_24755,N_21480,N_19581);
nand U24756 (N_24756,N_20894,N_19926);
xor U24757 (N_24757,N_18941,N_19844);
and U24758 (N_24758,N_21214,N_20358);
nand U24759 (N_24759,N_21338,N_20925);
or U24760 (N_24760,N_19465,N_18897);
nor U24761 (N_24761,N_19904,N_20935);
xor U24762 (N_24762,N_19261,N_19089);
nor U24763 (N_24763,N_20292,N_19161);
nand U24764 (N_24764,N_21344,N_19719);
nand U24765 (N_24765,N_19872,N_21776);
nand U24766 (N_24766,N_19807,N_20740);
or U24767 (N_24767,N_18789,N_20106);
nor U24768 (N_24768,N_19915,N_21805);
nand U24769 (N_24769,N_20077,N_21096);
and U24770 (N_24770,N_19400,N_21595);
and U24771 (N_24771,N_21106,N_21000);
or U24772 (N_24772,N_21178,N_19526);
nor U24773 (N_24773,N_19725,N_19175);
and U24774 (N_24774,N_19711,N_19382);
or U24775 (N_24775,N_21739,N_19597);
nor U24776 (N_24776,N_21328,N_21115);
or U24777 (N_24777,N_20732,N_21054);
or U24778 (N_24778,N_21241,N_20734);
and U24779 (N_24779,N_19499,N_19120);
and U24780 (N_24780,N_20414,N_19594);
or U24781 (N_24781,N_18796,N_18793);
nand U24782 (N_24782,N_20777,N_19782);
nand U24783 (N_24783,N_20745,N_21257);
or U24784 (N_24784,N_19501,N_19417);
nand U24785 (N_24785,N_19942,N_20052);
and U24786 (N_24786,N_20963,N_21628);
or U24787 (N_24787,N_21130,N_21114);
nor U24788 (N_24788,N_19948,N_19011);
nand U24789 (N_24789,N_19493,N_19070);
nand U24790 (N_24790,N_20250,N_20851);
and U24791 (N_24791,N_21384,N_19986);
nor U24792 (N_24792,N_19223,N_19569);
nor U24793 (N_24793,N_21630,N_19388);
and U24794 (N_24794,N_19669,N_19466);
or U24795 (N_24795,N_20380,N_21129);
nor U24796 (N_24796,N_21212,N_21525);
or U24797 (N_24797,N_19728,N_19898);
nor U24798 (N_24798,N_18956,N_20545);
or U24799 (N_24799,N_20850,N_21805);
or U24800 (N_24800,N_20925,N_21518);
or U24801 (N_24801,N_20667,N_19211);
nand U24802 (N_24802,N_20028,N_21638);
nand U24803 (N_24803,N_19916,N_20942);
nand U24804 (N_24804,N_20511,N_19189);
or U24805 (N_24805,N_19053,N_19975);
or U24806 (N_24806,N_20411,N_20677);
and U24807 (N_24807,N_21321,N_21723);
and U24808 (N_24808,N_19381,N_21535);
and U24809 (N_24809,N_20325,N_20287);
and U24810 (N_24810,N_21601,N_19627);
and U24811 (N_24811,N_21403,N_21371);
and U24812 (N_24812,N_21778,N_19260);
nor U24813 (N_24813,N_20449,N_20404);
nor U24814 (N_24814,N_19891,N_21407);
nor U24815 (N_24815,N_21807,N_20592);
and U24816 (N_24816,N_21791,N_19918);
and U24817 (N_24817,N_20294,N_20759);
or U24818 (N_24818,N_19724,N_19589);
nand U24819 (N_24819,N_18919,N_20317);
nor U24820 (N_24820,N_20223,N_20568);
nand U24821 (N_24821,N_19276,N_20709);
nor U24822 (N_24822,N_19068,N_20803);
xnor U24823 (N_24823,N_21170,N_19729);
nand U24824 (N_24824,N_19639,N_21437);
or U24825 (N_24825,N_21508,N_21051);
or U24826 (N_24826,N_19913,N_21632);
nand U24827 (N_24827,N_21250,N_19497);
nor U24828 (N_24828,N_20331,N_19620);
nor U24829 (N_24829,N_19895,N_20396);
and U24830 (N_24830,N_21490,N_20830);
or U24831 (N_24831,N_20168,N_19202);
nand U24832 (N_24832,N_20857,N_20922);
and U24833 (N_24833,N_21711,N_21302);
nor U24834 (N_24834,N_20449,N_18841);
nand U24835 (N_24835,N_19706,N_20153);
xor U24836 (N_24836,N_18906,N_20729);
or U24837 (N_24837,N_19413,N_19291);
and U24838 (N_24838,N_20669,N_19709);
or U24839 (N_24839,N_18841,N_21717);
nand U24840 (N_24840,N_20905,N_20692);
xor U24841 (N_24841,N_19629,N_20444);
nor U24842 (N_24842,N_21406,N_18795);
nand U24843 (N_24843,N_19368,N_20160);
nand U24844 (N_24844,N_21780,N_18868);
xor U24845 (N_24845,N_21399,N_20029);
nor U24846 (N_24846,N_20199,N_20640);
nand U24847 (N_24847,N_19948,N_20437);
nand U24848 (N_24848,N_20550,N_19833);
nand U24849 (N_24849,N_19318,N_19966);
nand U24850 (N_24850,N_20369,N_19998);
nor U24851 (N_24851,N_20385,N_19808);
nor U24852 (N_24852,N_19058,N_21612);
and U24853 (N_24853,N_20508,N_21287);
nand U24854 (N_24854,N_18793,N_19692);
and U24855 (N_24855,N_20633,N_21713);
and U24856 (N_24856,N_20065,N_21320);
nand U24857 (N_24857,N_20184,N_20285);
nor U24858 (N_24858,N_19562,N_20018);
nand U24859 (N_24859,N_21234,N_21151);
or U24860 (N_24860,N_20408,N_21770);
or U24861 (N_24861,N_20304,N_19894);
and U24862 (N_24862,N_20762,N_21633);
nand U24863 (N_24863,N_19481,N_20417);
or U24864 (N_24864,N_21721,N_18766);
and U24865 (N_24865,N_21063,N_21257);
and U24866 (N_24866,N_20936,N_20163);
xnor U24867 (N_24867,N_19469,N_21441);
nor U24868 (N_24868,N_20167,N_20569);
and U24869 (N_24869,N_19265,N_20138);
or U24870 (N_24870,N_21627,N_19181);
or U24871 (N_24871,N_21514,N_18842);
or U24872 (N_24872,N_20512,N_19244);
nor U24873 (N_24873,N_20248,N_18757);
or U24874 (N_24874,N_19803,N_21466);
or U24875 (N_24875,N_19187,N_21479);
and U24876 (N_24876,N_21439,N_21831);
and U24877 (N_24877,N_21848,N_18836);
and U24878 (N_24878,N_19699,N_20495);
nor U24879 (N_24879,N_19641,N_21788);
or U24880 (N_24880,N_18805,N_21196);
and U24881 (N_24881,N_19269,N_21684);
nand U24882 (N_24882,N_20459,N_21501);
nand U24883 (N_24883,N_20986,N_20706);
nor U24884 (N_24884,N_19753,N_20173);
and U24885 (N_24885,N_19569,N_20385);
nand U24886 (N_24886,N_19859,N_21535);
and U24887 (N_24887,N_21588,N_19358);
nand U24888 (N_24888,N_19762,N_21032);
xor U24889 (N_24889,N_20972,N_21501);
nand U24890 (N_24890,N_21592,N_21376);
nand U24891 (N_24891,N_21865,N_20698);
nor U24892 (N_24892,N_19027,N_18976);
xor U24893 (N_24893,N_19619,N_20875);
or U24894 (N_24894,N_20162,N_20001);
nand U24895 (N_24895,N_20277,N_18945);
and U24896 (N_24896,N_19732,N_19643);
or U24897 (N_24897,N_19756,N_20918);
and U24898 (N_24898,N_21536,N_21686);
and U24899 (N_24899,N_20356,N_21367);
nor U24900 (N_24900,N_19376,N_18910);
and U24901 (N_24901,N_18759,N_20165);
nor U24902 (N_24902,N_21856,N_20047);
and U24903 (N_24903,N_19790,N_20001);
nor U24904 (N_24904,N_19441,N_20555);
or U24905 (N_24905,N_19156,N_21209);
nand U24906 (N_24906,N_19566,N_19462);
and U24907 (N_24907,N_20485,N_18948);
or U24908 (N_24908,N_20713,N_19986);
nand U24909 (N_24909,N_19881,N_21370);
nor U24910 (N_24910,N_19814,N_19837);
nand U24911 (N_24911,N_20584,N_19297);
nor U24912 (N_24912,N_19119,N_20306);
nand U24913 (N_24913,N_20044,N_18924);
or U24914 (N_24914,N_20896,N_20547);
xor U24915 (N_24915,N_19503,N_21750);
and U24916 (N_24916,N_20293,N_21551);
nand U24917 (N_24917,N_18870,N_18966);
xnor U24918 (N_24918,N_18974,N_21183);
or U24919 (N_24919,N_18957,N_21803);
nor U24920 (N_24920,N_21628,N_20444);
xor U24921 (N_24921,N_21253,N_21657);
nor U24922 (N_24922,N_19152,N_19286);
or U24923 (N_24923,N_19381,N_19650);
nand U24924 (N_24924,N_21073,N_19340);
nor U24925 (N_24925,N_21234,N_20702);
or U24926 (N_24926,N_20143,N_20527);
and U24927 (N_24927,N_20839,N_19674);
nand U24928 (N_24928,N_18858,N_19798);
nand U24929 (N_24929,N_20456,N_21505);
or U24930 (N_24930,N_20386,N_21722);
or U24931 (N_24931,N_21339,N_19741);
nand U24932 (N_24932,N_19413,N_21397);
nor U24933 (N_24933,N_19904,N_19840);
nand U24934 (N_24934,N_19070,N_20676);
nor U24935 (N_24935,N_20063,N_19688);
or U24936 (N_24936,N_20161,N_19855);
and U24937 (N_24937,N_21732,N_19111);
nand U24938 (N_24938,N_21008,N_21376);
and U24939 (N_24939,N_21220,N_19926);
and U24940 (N_24940,N_19490,N_19796);
nand U24941 (N_24941,N_21011,N_19363);
xor U24942 (N_24942,N_21698,N_21275);
nor U24943 (N_24943,N_19832,N_21821);
and U24944 (N_24944,N_19702,N_19482);
nor U24945 (N_24945,N_20036,N_21394);
and U24946 (N_24946,N_20158,N_18805);
or U24947 (N_24947,N_20768,N_20778);
or U24948 (N_24948,N_20065,N_19912);
or U24949 (N_24949,N_21576,N_20860);
nand U24950 (N_24950,N_20060,N_21043);
xor U24951 (N_24951,N_21239,N_19493);
and U24952 (N_24952,N_21122,N_20167);
or U24953 (N_24953,N_20781,N_19936);
nand U24954 (N_24954,N_19156,N_21257);
or U24955 (N_24955,N_19901,N_21217);
or U24956 (N_24956,N_21774,N_21024);
nand U24957 (N_24957,N_21426,N_20848);
nor U24958 (N_24958,N_19948,N_18880);
or U24959 (N_24959,N_19717,N_19629);
xor U24960 (N_24960,N_21437,N_19028);
or U24961 (N_24961,N_21566,N_20513);
nor U24962 (N_24962,N_20831,N_19690);
or U24963 (N_24963,N_19934,N_21225);
or U24964 (N_24964,N_20193,N_18867);
xnor U24965 (N_24965,N_20988,N_19817);
nand U24966 (N_24966,N_20852,N_21248);
or U24967 (N_24967,N_20390,N_20637);
nand U24968 (N_24968,N_20997,N_18755);
nand U24969 (N_24969,N_19946,N_20339);
or U24970 (N_24970,N_21309,N_19891);
nand U24971 (N_24971,N_20944,N_21320);
nor U24972 (N_24972,N_18857,N_19770);
nor U24973 (N_24973,N_21282,N_21344);
and U24974 (N_24974,N_20457,N_20205);
nand U24975 (N_24975,N_19360,N_19629);
nand U24976 (N_24976,N_21539,N_20972);
and U24977 (N_24977,N_18847,N_19719);
xnor U24978 (N_24978,N_21507,N_19646);
nor U24979 (N_24979,N_20196,N_19571);
nor U24980 (N_24980,N_20440,N_20029);
nand U24981 (N_24981,N_20653,N_21811);
nand U24982 (N_24982,N_19882,N_19976);
and U24983 (N_24983,N_20427,N_21103);
nand U24984 (N_24984,N_20685,N_21216);
nand U24985 (N_24985,N_19806,N_21058);
or U24986 (N_24986,N_21475,N_20632);
nand U24987 (N_24987,N_19693,N_20586);
or U24988 (N_24988,N_20656,N_20813);
nand U24989 (N_24989,N_21420,N_19003);
nand U24990 (N_24990,N_21192,N_21052);
nor U24991 (N_24991,N_19400,N_21772);
and U24992 (N_24992,N_19379,N_20967);
and U24993 (N_24993,N_20739,N_21167);
or U24994 (N_24994,N_21209,N_19791);
nor U24995 (N_24995,N_21167,N_20936);
nand U24996 (N_24996,N_18993,N_21293);
xnor U24997 (N_24997,N_19519,N_18861);
nor U24998 (N_24998,N_20831,N_19970);
nand U24999 (N_24999,N_19091,N_19561);
nor UO_0 (O_0,N_23719,N_23810);
and UO_1 (O_1,N_23300,N_22914);
nor UO_2 (O_2,N_23524,N_24716);
xor UO_3 (O_3,N_24628,N_24599);
nor UO_4 (O_4,N_24002,N_23016);
and UO_5 (O_5,N_22208,N_22248);
nand UO_6 (O_6,N_23648,N_23462);
and UO_7 (O_7,N_22708,N_22245);
xor UO_8 (O_8,N_23223,N_23705);
xor UO_9 (O_9,N_22060,N_23944);
nor UO_10 (O_10,N_24784,N_24634);
xor UO_11 (O_11,N_21964,N_23180);
or UO_12 (O_12,N_24683,N_24024);
nor UO_13 (O_13,N_24162,N_23573);
nand UO_14 (O_14,N_22606,N_23495);
xor UO_15 (O_15,N_23616,N_23100);
and UO_16 (O_16,N_22927,N_23094);
and UO_17 (O_17,N_24943,N_22589);
and UO_18 (O_18,N_22316,N_22607);
or UO_19 (O_19,N_24397,N_24865);
or UO_20 (O_20,N_22683,N_23506);
or UO_21 (O_21,N_24228,N_24772);
nor UO_22 (O_22,N_22077,N_24998);
and UO_23 (O_23,N_24500,N_24991);
nand UO_24 (O_24,N_23844,N_22337);
nor UO_25 (O_25,N_24733,N_23988);
or UO_26 (O_26,N_22534,N_23665);
and UO_27 (O_27,N_22151,N_23168);
xor UO_28 (O_28,N_24742,N_21967);
and UO_29 (O_29,N_24803,N_23240);
and UO_30 (O_30,N_22089,N_22689);
or UO_31 (O_31,N_24701,N_24040);
nand UO_32 (O_32,N_22545,N_22419);
or UO_33 (O_33,N_24199,N_23942);
and UO_34 (O_34,N_22229,N_24068);
nand UO_35 (O_35,N_24677,N_24556);
and UO_36 (O_36,N_24714,N_22520);
nor UO_37 (O_37,N_24394,N_23801);
and UO_38 (O_38,N_22065,N_22351);
and UO_39 (O_39,N_24353,N_22891);
nand UO_40 (O_40,N_23649,N_22672);
nor UO_41 (O_41,N_23184,N_24313);
and UO_42 (O_42,N_22384,N_21917);
and UO_43 (O_43,N_24250,N_24477);
nor UO_44 (O_44,N_23429,N_23785);
or UO_45 (O_45,N_24052,N_23015);
or UO_46 (O_46,N_22124,N_23087);
or UO_47 (O_47,N_22734,N_22451);
nor UO_48 (O_48,N_24632,N_22243);
and UO_49 (O_49,N_23084,N_24091);
nand UO_50 (O_50,N_21999,N_24098);
or UO_51 (O_51,N_22438,N_24764);
xnor UO_52 (O_52,N_23272,N_24910);
nand UO_53 (O_53,N_24799,N_24782);
xnor UO_54 (O_54,N_23046,N_24125);
nand UO_55 (O_55,N_24017,N_22619);
nand UO_56 (O_56,N_23940,N_22241);
or UO_57 (O_57,N_22043,N_22705);
or UO_58 (O_58,N_23805,N_24331);
and UO_59 (O_59,N_24303,N_24592);
nand UO_60 (O_60,N_24456,N_24623);
nand UO_61 (O_61,N_22885,N_24438);
or UO_62 (O_62,N_24375,N_22174);
and UO_63 (O_63,N_22614,N_22573);
nor UO_64 (O_64,N_22758,N_22709);
nand UO_65 (O_65,N_23893,N_23259);
nand UO_66 (O_66,N_23872,N_22706);
and UO_67 (O_67,N_24395,N_24618);
or UO_68 (O_68,N_22293,N_22697);
and UO_69 (O_69,N_22536,N_22602);
and UO_70 (O_70,N_24740,N_22583);
and UO_71 (O_71,N_24968,N_22290);
xnor UO_72 (O_72,N_23209,N_24439);
xor UO_73 (O_73,N_23400,N_22329);
nor UO_74 (O_74,N_23271,N_24458);
or UO_75 (O_75,N_23324,N_23936);
or UO_76 (O_76,N_24342,N_22559);
and UO_77 (O_77,N_21927,N_22235);
nor UO_78 (O_78,N_24014,N_22232);
nand UO_79 (O_79,N_23512,N_24702);
and UO_80 (O_80,N_24806,N_23191);
and UO_81 (O_81,N_23814,N_23569);
nand UO_82 (O_82,N_23956,N_22464);
nand UO_83 (O_83,N_23832,N_21928);
or UO_84 (O_84,N_23855,N_24792);
nand UO_85 (O_85,N_22433,N_22122);
or UO_86 (O_86,N_22853,N_21909);
nor UO_87 (O_87,N_22244,N_22187);
nand UO_88 (O_88,N_21933,N_22524);
nand UO_89 (O_89,N_23018,N_24452);
nand UO_90 (O_90,N_22681,N_23663);
and UO_91 (O_91,N_23234,N_23221);
nand UO_92 (O_92,N_24744,N_23886);
and UO_93 (O_93,N_22726,N_24533);
or UO_94 (O_94,N_22106,N_22677);
and UO_95 (O_95,N_24494,N_22572);
nor UO_96 (O_96,N_22056,N_23771);
nor UO_97 (O_97,N_23291,N_22225);
and UO_98 (O_98,N_24150,N_23391);
or UO_99 (O_99,N_24185,N_23717);
or UO_100 (O_100,N_24406,N_23837);
nor UO_101 (O_101,N_24271,N_22813);
nand UO_102 (O_102,N_22470,N_23135);
nand UO_103 (O_103,N_24774,N_23390);
nand UO_104 (O_104,N_24606,N_22586);
nor UO_105 (O_105,N_24905,N_23615);
or UO_106 (O_106,N_23434,N_23368);
and UO_107 (O_107,N_23147,N_24027);
nor UO_108 (O_108,N_22529,N_22805);
or UO_109 (O_109,N_22367,N_23661);
nand UO_110 (O_110,N_23525,N_23971);
nand UO_111 (O_111,N_22019,N_22539);
xor UO_112 (O_112,N_23351,N_24647);
nand UO_113 (O_113,N_23668,N_23593);
nand UO_114 (O_114,N_22675,N_24976);
nand UO_115 (O_115,N_22195,N_23114);
nand UO_116 (O_116,N_23773,N_24444);
or UO_117 (O_117,N_22863,N_22100);
or UO_118 (O_118,N_24895,N_22003);
or UO_119 (O_119,N_24107,N_24723);
nand UO_120 (O_120,N_23210,N_23739);
nand UO_121 (O_121,N_23786,N_23652);
nor UO_122 (O_122,N_23000,N_24241);
xnor UO_123 (O_123,N_23533,N_23582);
and UO_124 (O_124,N_23458,N_24621);
or UO_125 (O_125,N_24385,N_24255);
or UO_126 (O_126,N_23357,N_24745);
or UO_127 (O_127,N_23348,N_24420);
nor UO_128 (O_128,N_23857,N_22047);
nand UO_129 (O_129,N_23938,N_24022);
and UO_130 (O_130,N_22652,N_24167);
nor UO_131 (O_131,N_24209,N_22514);
xnor UO_132 (O_132,N_23023,N_23897);
nand UO_133 (O_133,N_22009,N_22458);
xnor UO_134 (O_134,N_24163,N_24585);
and UO_135 (O_135,N_22303,N_23726);
nand UO_136 (O_136,N_22411,N_23662);
and UO_137 (O_137,N_24748,N_23101);
and UO_138 (O_138,N_23774,N_22829);
or UO_139 (O_139,N_22560,N_24448);
or UO_140 (O_140,N_24773,N_24622);
or UO_141 (O_141,N_23748,N_23123);
xnor UO_142 (O_142,N_23288,N_23407);
nand UO_143 (O_143,N_24627,N_23039);
or UO_144 (O_144,N_24902,N_23061);
nor UO_145 (O_145,N_22111,N_23102);
and UO_146 (O_146,N_22157,N_23231);
nand UO_147 (O_147,N_23678,N_23409);
nor UO_148 (O_148,N_24405,N_22716);
nand UO_149 (O_149,N_24089,N_21876);
xnor UO_150 (O_150,N_23451,N_23833);
nand UO_151 (O_151,N_24478,N_24364);
nor UO_152 (O_152,N_23667,N_22873);
xnor UO_153 (O_153,N_24609,N_24785);
and UO_154 (O_154,N_24328,N_21958);
nor UO_155 (O_155,N_24301,N_23729);
nand UO_156 (O_156,N_23762,N_22158);
nor UO_157 (O_157,N_22605,N_22335);
nand UO_158 (O_158,N_24314,N_22966);
nor UO_159 (O_159,N_24189,N_23268);
nand UO_160 (O_160,N_24577,N_23213);
and UO_161 (O_161,N_23378,N_22204);
and UO_162 (O_162,N_22727,N_22240);
xnor UO_163 (O_163,N_24260,N_23284);
nor UO_164 (O_164,N_23881,N_23037);
and UO_165 (O_165,N_24276,N_23267);
nand UO_166 (O_166,N_24690,N_24719);
nor UO_167 (O_167,N_23585,N_23352);
or UO_168 (O_168,N_24750,N_22164);
or UO_169 (O_169,N_23469,N_23232);
and UO_170 (O_170,N_23260,N_22661);
nor UO_171 (O_171,N_22183,N_22112);
nor UO_172 (O_172,N_24761,N_24265);
xnor UO_173 (O_173,N_23273,N_22944);
or UO_174 (O_174,N_22078,N_23962);
nand UO_175 (O_175,N_23594,N_22830);
xnor UO_176 (O_176,N_23555,N_24198);
nand UO_177 (O_177,N_24629,N_22742);
nand UO_178 (O_178,N_24411,N_21994);
nand UO_179 (O_179,N_22025,N_24009);
xor UO_180 (O_180,N_23425,N_23176);
or UO_181 (O_181,N_21990,N_24807);
nand UO_182 (O_182,N_22334,N_22063);
and UO_183 (O_183,N_21893,N_24156);
xor UO_184 (O_184,N_22656,N_22013);
nor UO_185 (O_185,N_23941,N_21978);
nor UO_186 (O_186,N_22379,N_22205);
and UO_187 (O_187,N_24416,N_24994);
and UO_188 (O_188,N_22259,N_22173);
and UO_189 (O_189,N_22937,N_23250);
or UO_190 (O_190,N_24642,N_22511);
or UO_191 (O_191,N_23170,N_22506);
or UO_192 (O_192,N_24065,N_24694);
or UO_193 (O_193,N_23518,N_24915);
or UO_194 (O_194,N_22882,N_23758);
nand UO_195 (O_195,N_22048,N_23295);
nor UO_196 (O_196,N_23611,N_23638);
and UO_197 (O_197,N_22980,N_23013);
nor UO_198 (O_198,N_22234,N_24933);
and UO_199 (O_199,N_22219,N_22986);
nand UO_200 (O_200,N_22880,N_24412);
or UO_201 (O_201,N_24111,N_23924);
nand UO_202 (O_202,N_22509,N_22531);
or UO_203 (O_203,N_22185,N_22081);
and UO_204 (O_204,N_23241,N_22167);
or UO_205 (O_205,N_24979,N_22866);
or UO_206 (O_206,N_22749,N_24114);
or UO_207 (O_207,N_22938,N_22249);
xnor UO_208 (O_208,N_24851,N_24259);
xor UO_209 (O_209,N_23394,N_22220);
nand UO_210 (O_210,N_22069,N_23831);
or UO_211 (O_211,N_24455,N_24842);
and UO_212 (O_212,N_23970,N_24832);
nand UO_213 (O_213,N_22859,N_24866);
and UO_214 (O_214,N_23601,N_22038);
and UO_215 (O_215,N_23050,N_24435);
nand UO_216 (O_216,N_24984,N_24318);
nand UO_217 (O_217,N_22997,N_24018);
xor UO_218 (O_218,N_24214,N_22800);
nor UO_219 (O_219,N_24769,N_24777);
or UO_220 (O_220,N_22094,N_24044);
nand UO_221 (O_221,N_23850,N_22169);
or UO_222 (O_222,N_22551,N_23497);
or UO_223 (O_223,N_24124,N_23787);
or UO_224 (O_224,N_23825,N_23858);
nor UO_225 (O_225,N_24703,N_23381);
nand UO_226 (O_226,N_24952,N_22504);
and UO_227 (O_227,N_23575,N_24559);
or UO_228 (O_228,N_22600,N_22999);
or UO_229 (O_229,N_23520,N_24864);
nor UO_230 (O_230,N_22816,N_22155);
nand UO_231 (O_231,N_24457,N_23728);
or UO_232 (O_232,N_24853,N_23182);
or UO_233 (O_233,N_21985,N_22945);
or UO_234 (O_234,N_23522,N_24734);
nor UO_235 (O_235,N_23749,N_23529);
and UO_236 (O_236,N_23756,N_23365);
nand UO_237 (O_237,N_22802,N_24759);
and UO_238 (O_238,N_22569,N_22403);
xnor UO_239 (O_239,N_22622,N_22924);
and UO_240 (O_240,N_24138,N_23053);
nor UO_241 (O_241,N_23727,N_23354);
nor UO_242 (O_242,N_23305,N_23784);
nand UO_243 (O_243,N_24726,N_22730);
nor UO_244 (O_244,N_23119,N_24031);
nor UO_245 (O_245,N_23973,N_23983);
nand UO_246 (O_246,N_24668,N_24434);
and UO_247 (O_247,N_24678,N_24539);
and UO_248 (O_248,N_22430,N_22254);
or UO_249 (O_249,N_23507,N_24421);
or UO_250 (O_250,N_22717,N_23413);
nand UO_251 (O_251,N_24083,N_23280);
and UO_252 (O_252,N_22527,N_23150);
nand UO_253 (O_253,N_23383,N_22454);
nor UO_254 (O_254,N_21992,N_23164);
nor UO_255 (O_255,N_24309,N_22921);
and UO_256 (O_256,N_22485,N_23031);
and UO_257 (O_257,N_23715,N_24382);
xor UO_258 (O_258,N_24857,N_22434);
nor UO_259 (O_259,N_24685,N_23446);
nor UO_260 (O_260,N_22242,N_23371);
nand UO_261 (O_261,N_24201,N_22620);
nand UO_262 (O_262,N_24431,N_23532);
and UO_263 (O_263,N_21897,N_24006);
or UO_264 (O_264,N_24555,N_23068);
or UO_265 (O_265,N_23939,N_24780);
nand UO_266 (O_266,N_22090,N_23112);
nor UO_267 (O_267,N_24358,N_24471);
xor UO_268 (O_268,N_23121,N_23318);
nor UO_269 (O_269,N_23201,N_22250);
nor UO_270 (O_270,N_23613,N_22759);
or UO_271 (O_271,N_24131,N_23257);
and UO_272 (O_272,N_24779,N_24173);
and UO_273 (O_273,N_22718,N_22275);
nand UO_274 (O_274,N_23803,N_22045);
and UO_275 (O_275,N_22538,N_22501);
and UO_276 (O_276,N_22670,N_22324);
nand UO_277 (O_277,N_24920,N_23106);
and UO_278 (O_278,N_24921,N_22400);
xnor UO_279 (O_279,N_22883,N_24597);
or UO_280 (O_280,N_24880,N_24981);
and UO_281 (O_281,N_24760,N_24337);
nand UO_282 (O_282,N_24486,N_24881);
nand UO_283 (O_283,N_24369,N_22722);
nor UO_284 (O_284,N_22998,N_24117);
and UO_285 (O_285,N_24959,N_24196);
or UO_286 (O_286,N_23328,N_22348);
xnor UO_287 (O_287,N_24365,N_24058);
nor UO_288 (O_288,N_23049,N_24914);
or UO_289 (O_289,N_21889,N_22668);
and UO_290 (O_290,N_23994,N_24443);
xnor UO_291 (O_291,N_24312,N_24280);
nor UO_292 (O_292,N_23809,N_24330);
or UO_293 (O_293,N_22841,N_22926);
nor UO_294 (O_294,N_24275,N_23190);
or UO_295 (O_295,N_23479,N_23969);
nor UO_296 (O_296,N_24182,N_23847);
nor UO_297 (O_297,N_24958,N_23865);
nand UO_298 (O_298,N_24219,N_22868);
nor UO_299 (O_299,N_23574,N_22973);
xnor UO_300 (O_300,N_24466,N_23004);
nand UO_301 (O_301,N_23961,N_21892);
or UO_302 (O_302,N_23565,N_24713);
nand UO_303 (O_303,N_24611,N_22760);
nand UO_304 (O_304,N_22936,N_22497);
or UO_305 (O_305,N_24119,N_23437);
nor UO_306 (O_306,N_23521,N_23889);
nor UO_307 (O_307,N_22057,N_23751);
and UO_308 (O_308,N_23951,N_21883);
xnor UO_309 (O_309,N_22375,N_24472);
and UO_310 (O_310,N_24693,N_23722);
nand UO_311 (O_311,N_22644,N_22005);
or UO_312 (O_312,N_24168,N_24752);
xnor UO_313 (O_313,N_22030,N_24268);
and UO_314 (O_314,N_23539,N_23914);
nand UO_315 (O_315,N_24333,N_24964);
nor UO_316 (O_316,N_24553,N_23968);
and UO_317 (O_317,N_22093,N_23949);
or UO_318 (O_318,N_23041,N_24927);
or UO_319 (O_319,N_22922,N_24637);
or UO_320 (O_320,N_22892,N_22828);
nor UO_321 (O_321,N_22975,N_24184);
or UO_322 (O_322,N_24925,N_23266);
nor UO_323 (O_323,N_22424,N_23974);
or UO_324 (O_324,N_24134,N_23852);
nor UO_325 (O_325,N_23608,N_23544);
xor UO_326 (O_326,N_22765,N_24589);
xnor UO_327 (O_327,N_24446,N_24519);
nor UO_328 (O_328,N_24639,N_22263);
and UO_329 (O_329,N_23366,N_24004);
and UO_330 (O_330,N_22831,N_22554);
and UO_331 (O_331,N_22212,N_23227);
and UO_332 (O_332,N_24176,N_21997);
and UO_333 (O_333,N_24436,N_23778);
nand UO_334 (O_334,N_22020,N_24410);
or UO_335 (O_335,N_24242,N_24798);
nand UO_336 (O_336,N_23912,N_22915);
and UO_337 (O_337,N_24822,N_24573);
nor UO_338 (O_338,N_24657,N_22894);
and UO_339 (O_339,N_24025,N_23396);
or UO_340 (O_340,N_23070,N_24430);
or UO_341 (O_341,N_23489,N_23345);
or UO_342 (O_342,N_24442,N_23737);
and UO_343 (O_343,N_24956,N_22756);
xnor UO_344 (O_344,N_22189,N_23731);
or UO_345 (O_345,N_22448,N_22771);
xor UO_346 (O_346,N_23108,N_23927);
or UO_347 (O_347,N_22188,N_23278);
nor UO_348 (O_348,N_22532,N_22415);
nor UO_349 (O_349,N_22092,N_24546);
or UO_350 (O_350,N_22663,N_23460);
nor UO_351 (O_351,N_24730,N_23598);
or UO_352 (O_352,N_22781,N_22713);
or UO_353 (O_353,N_23995,N_23782);
nor UO_354 (O_354,N_22299,N_22276);
and UO_355 (O_355,N_22305,N_24705);
xnor UO_356 (O_356,N_21887,N_24158);
and UO_357 (O_357,N_22941,N_22669);
nor UO_358 (O_358,N_24654,N_21878);
and UO_359 (O_359,N_22297,N_24578);
nor UO_360 (O_360,N_23781,N_22657);
and UO_361 (O_361,N_24147,N_23159);
or UO_362 (O_362,N_23490,N_24960);
nor UO_363 (O_363,N_22694,N_24287);
nand UO_364 (O_364,N_22685,N_23776);
xnor UO_365 (O_365,N_22590,N_23768);
or UO_366 (O_366,N_24924,N_22812);
and UO_367 (O_367,N_24190,N_24045);
nand UO_368 (O_368,N_24207,N_22349);
xnor UO_369 (O_369,N_24349,N_23484);
and UO_370 (O_370,N_22493,N_23235);
xnor UO_371 (O_371,N_22273,N_23370);
xnor UO_372 (O_372,N_21948,N_23836);
nor UO_373 (O_373,N_24237,N_23723);
or UO_374 (O_374,N_22823,N_22416);
nor UO_375 (O_375,N_22682,N_24279);
xor UO_376 (O_376,N_23205,N_23360);
nor UO_377 (O_377,N_24122,N_24978);
xor UO_378 (O_378,N_21974,N_24273);
or UO_379 (O_379,N_24635,N_23829);
or UO_380 (O_380,N_21926,N_24544);
nor UO_381 (O_381,N_24602,N_22721);
nor UO_382 (O_382,N_23247,N_23416);
or UO_383 (O_383,N_21932,N_24977);
xor UO_384 (O_384,N_24229,N_24946);
nor UO_385 (O_385,N_24208,N_21938);
nor UO_386 (O_386,N_24204,N_23424);
and UO_387 (O_387,N_23309,N_22691);
nor UO_388 (O_388,N_24451,N_23214);
nor UO_389 (O_389,N_24586,N_22137);
xor UO_390 (O_390,N_24775,N_22638);
xnor UO_391 (O_391,N_23989,N_23561);
nor UO_392 (O_392,N_23845,N_23285);
and UO_393 (O_393,N_24712,N_23978);
nor UO_394 (O_394,N_23606,N_22140);
and UO_395 (O_395,N_23780,N_24766);
nand UO_396 (O_396,N_24239,N_22292);
and UO_397 (O_397,N_24576,N_24523);
and UO_398 (O_398,N_21900,N_22983);
xnor UO_399 (O_399,N_22982,N_22322);
xnor UO_400 (O_400,N_22897,N_21915);
or UO_401 (O_401,N_24852,N_23153);
and UO_402 (O_402,N_24076,N_22405);
and UO_403 (O_403,N_23146,N_22623);
and UO_404 (O_404,N_22072,N_22022);
nand UO_405 (O_405,N_24088,N_23204);
or UO_406 (O_406,N_24671,N_23943);
or UO_407 (O_407,N_24240,N_24050);
nand UO_408 (O_408,N_23261,N_24743);
nand UO_409 (O_409,N_24347,N_22363);
nand UO_410 (O_410,N_24195,N_24953);
nor UO_411 (O_411,N_22001,N_22857);
nand UO_412 (O_412,N_22775,N_23898);
or UO_413 (O_413,N_22932,N_22645);
and UO_414 (O_414,N_23450,N_23686);
nor UO_415 (O_415,N_22877,N_22080);
nand UO_416 (O_416,N_23807,N_23523);
or UO_417 (O_417,N_22484,N_24912);
nor UO_418 (O_418,N_23406,N_23528);
or UO_419 (O_419,N_22135,N_24097);
and UO_420 (O_420,N_22395,N_22006);
xnor UO_421 (O_421,N_23704,N_23393);
or UO_422 (O_422,N_24728,N_23165);
and UO_423 (O_423,N_22702,N_22651);
xor UO_424 (O_424,N_22996,N_24288);
xnor UO_425 (O_425,N_22147,N_24561);
nor UO_426 (O_426,N_22845,N_23137);
or UO_427 (O_427,N_24433,N_24863);
nor UO_428 (O_428,N_23579,N_24949);
xnor UO_429 (O_429,N_24811,N_23932);
or UO_430 (O_430,N_23903,N_24536);
nand UO_431 (O_431,N_22311,N_24243);
and UO_432 (O_432,N_23981,N_24428);
nand UO_433 (O_433,N_22754,N_24437);
nor UO_434 (O_434,N_24708,N_22585);
nand UO_435 (O_435,N_23331,N_24732);
nor UO_436 (O_436,N_24890,N_24529);
or UO_437 (O_437,N_24310,N_23003);
nand UO_438 (O_438,N_24178,N_24212);
or UO_439 (O_439,N_22846,N_24590);
or UO_440 (O_440,N_24537,N_22824);
xor UO_441 (O_441,N_23619,N_24344);
and UO_442 (O_442,N_23851,N_23913);
and UO_443 (O_443,N_24215,N_24356);
nand UO_444 (O_444,N_24821,N_21919);
and UO_445 (O_445,N_22487,N_21925);
and UO_446 (O_446,N_23526,N_22378);
and UO_447 (O_447,N_24474,N_24815);
nand UO_448 (O_448,N_22655,N_24916);
nor UO_449 (O_449,N_23027,N_22177);
nand UO_450 (O_450,N_24736,N_22918);
nor UO_451 (O_451,N_22432,N_23498);
or UO_452 (O_452,N_24795,N_23026);
or UO_453 (O_453,N_22021,N_22162);
nor UO_454 (O_454,N_24492,N_22104);
nand UO_455 (O_455,N_21943,N_22878);
and UO_456 (O_456,N_22900,N_24620);
nor UO_457 (O_457,N_22666,N_23783);
xor UO_458 (O_458,N_24859,N_22797);
and UO_459 (O_459,N_24963,N_23056);
nor UO_460 (O_460,N_24571,N_23179);
xnor UO_461 (O_461,N_21902,N_22624);
and UO_462 (O_462,N_24982,N_23230);
nand UO_463 (O_463,N_24465,N_22904);
or UO_464 (O_464,N_22673,N_23483);
nor UO_465 (O_465,N_24464,N_24306);
xor UO_466 (O_466,N_23796,N_21891);
nor UO_467 (O_467,N_24481,N_22376);
nor UO_468 (O_468,N_24797,N_22410);
or UO_469 (O_469,N_21888,N_24160);
nor UO_470 (O_470,N_23542,N_22194);
nor UO_471 (O_471,N_23966,N_22393);
nor UO_472 (O_472,N_23626,N_23248);
nand UO_473 (O_473,N_21920,N_24957);
and UO_474 (O_474,N_22643,N_22460);
or UO_475 (O_475,N_22847,N_24662);
nand UO_476 (O_476,N_24901,N_22435);
nor UO_477 (O_477,N_23639,N_24174);
nor UO_478 (O_478,N_24407,N_22495);
or UO_479 (O_479,N_23079,N_22385);
nand UO_480 (O_480,N_24139,N_24129);
and UO_481 (O_481,N_24922,N_23873);
nand UO_482 (O_482,N_24522,N_22965);
nand UO_483 (O_483,N_22370,N_24415);
xnor UO_484 (O_484,N_24033,N_23307);
nor UO_485 (O_485,N_23591,N_24459);
nor UO_486 (O_486,N_24569,N_24367);
and UO_487 (O_487,N_22784,N_24289);
nor UO_488 (O_488,N_22196,N_22099);
nor UO_489 (O_489,N_23602,N_24661);
and UO_490 (O_490,N_23864,N_23110);
nand UO_491 (O_491,N_22171,N_22518);
and UO_492 (O_492,N_22130,N_23802);
nor UO_493 (O_493,N_23511,N_23742);
or UO_494 (O_494,N_23349,N_23118);
nand UO_495 (O_495,N_23198,N_24918);
and UO_496 (O_496,N_24505,N_23568);
and UO_497 (O_497,N_22895,N_24805);
xnor UO_498 (O_498,N_23379,N_24840);
and UO_499 (O_499,N_23551,N_22023);
nor UO_500 (O_500,N_24128,N_22768);
or UO_501 (O_501,N_23792,N_24325);
xnor UO_502 (O_502,N_22499,N_22126);
and UO_503 (O_503,N_24659,N_22558);
nor UO_504 (O_504,N_23047,N_23933);
and UO_505 (O_505,N_24591,N_22058);
xnor UO_506 (O_506,N_24648,N_22640);
and UO_507 (O_507,N_22601,N_23724);
nand UO_508 (O_508,N_23627,N_24809);
and UO_509 (O_509,N_24041,N_22287);
nand UO_510 (O_510,N_24211,N_24404);
nor UO_511 (O_511,N_22455,N_24264);
or UO_512 (O_512,N_23072,N_22611);
or UO_513 (O_513,N_24887,N_24531);
nor UO_514 (O_514,N_23696,N_22182);
nor UO_515 (O_515,N_24320,N_22546);
nor UO_516 (O_516,N_23888,N_23997);
and UO_517 (O_517,N_24944,N_24913);
nand UO_518 (O_518,N_22553,N_21957);
or UO_519 (O_519,N_23274,N_22972);
xnor UO_520 (O_520,N_22085,N_23398);
and UO_521 (O_521,N_22799,N_23545);
nor UO_522 (O_522,N_22226,N_22832);
and UO_523 (O_523,N_24715,N_24048);
nor UO_524 (O_524,N_24691,N_24108);
or UO_525 (O_525,N_23317,N_23559);
nand UO_526 (O_526,N_22256,N_24100);
or UO_527 (O_527,N_24062,N_23999);
or UO_528 (O_528,N_23487,N_24540);
and UO_529 (O_529,N_21998,N_22159);
xor UO_530 (O_530,N_24476,N_22837);
nor UO_531 (O_531,N_23028,N_24092);
nand UO_532 (O_532,N_24619,N_23090);
nand UO_533 (O_533,N_22636,N_23327);
xnor UO_534 (O_534,N_22597,N_23998);
or UO_535 (O_535,N_23452,N_24814);
and UO_536 (O_536,N_24247,N_22555);
or UO_537 (O_537,N_21951,N_23677);
nor UO_538 (O_538,N_23842,N_24077);
nand UO_539 (O_539,N_23812,N_22264);
nand UO_540 (O_540,N_24485,N_23955);
nor UO_541 (O_541,N_24532,N_23367);
or UO_542 (O_542,N_23987,N_23759);
xnor UO_543 (O_543,N_21950,N_22664);
nor UO_544 (O_544,N_24007,N_24298);
nand UO_545 (O_545,N_24600,N_23993);
or UO_546 (O_546,N_22654,N_23604);
nor UO_547 (O_547,N_22979,N_24141);
nand UO_548 (O_548,N_22138,N_24898);
nor UO_549 (O_549,N_24917,N_23060);
nor UO_550 (O_550,N_24362,N_23915);
or UO_551 (O_551,N_22616,N_22959);
nor UO_552 (O_552,N_24063,N_22508);
or UO_553 (O_553,N_21969,N_22821);
and UO_554 (O_554,N_22662,N_23823);
or UO_555 (O_555,N_22383,N_22864);
nand UO_556 (O_556,N_23024,N_22200);
xor UO_557 (O_557,N_24975,N_24094);
nor UO_558 (O_558,N_21955,N_24491);
or UO_559 (O_559,N_23550,N_22255);
and UO_560 (O_560,N_23660,N_23103);
or UO_561 (O_561,N_23646,N_24381);
nand UO_562 (O_562,N_23321,N_22418);
or UO_563 (O_563,N_23258,N_21882);
nand UO_564 (O_564,N_21936,N_24688);
or UO_565 (O_565,N_22631,N_22178);
or UO_566 (O_566,N_24153,N_22066);
nand UO_567 (O_567,N_22908,N_23076);
nor UO_568 (O_568,N_22779,N_23732);
nand UO_569 (O_569,N_22227,N_24820);
nor UO_570 (O_570,N_24057,N_23217);
nor UO_571 (O_571,N_22591,N_24484);
xnor UO_572 (O_572,N_24285,N_23707);
nand UO_573 (O_573,N_24470,N_23980);
nand UO_574 (O_574,N_23376,N_22517);
and UO_575 (O_575,N_24072,N_22548);
and UO_576 (O_576,N_23946,N_23421);
nand UO_577 (O_577,N_24300,N_22388);
and UO_578 (O_578,N_23343,N_22333);
nand UO_579 (O_579,N_24136,N_21956);
nand UO_580 (O_580,N_23211,N_23251);
nand UO_581 (O_581,N_23928,N_24473);
and UO_582 (O_582,N_23455,N_22660);
and UO_583 (O_583,N_23043,N_24879);
nor UO_584 (O_584,N_23329,N_24625);
nand UO_585 (O_585,N_23332,N_24867);
nor UO_586 (O_586,N_23297,N_24023);
and UO_587 (O_587,N_23605,N_22500);
or UO_588 (O_588,N_24810,N_24951);
and UO_589 (O_589,N_24445,N_23797);
and UO_590 (O_590,N_23244,N_22482);
nand UO_591 (O_591,N_22309,N_22352);
nor UO_592 (O_592,N_23656,N_23007);
nor UO_593 (O_593,N_23493,N_22778);
and UO_594 (O_594,N_23044,N_22018);
nor UO_595 (O_595,N_24940,N_24542);
and UO_596 (O_596,N_24377,N_21886);
and UO_597 (O_597,N_24770,N_23081);
nor UO_598 (O_598,N_22787,N_24543);
nand UO_599 (O_599,N_23860,N_23503);
nor UO_600 (O_600,N_22494,N_24938);
or UO_601 (O_601,N_22772,N_22886);
nand UO_602 (O_602,N_23821,N_24236);
xor UO_603 (O_603,N_23287,N_21898);
nand UO_604 (O_604,N_22486,N_24427);
nor UO_605 (O_605,N_22210,N_24010);
xor UO_606 (O_606,N_22002,N_23510);
xor UO_607 (O_607,N_22236,N_22840);
and UO_608 (O_608,N_24520,N_24564);
or UO_609 (O_609,N_23906,N_24487);
nor UO_610 (O_610,N_21953,N_22457);
nand UO_611 (O_611,N_23990,N_23249);
and UO_612 (O_612,N_22929,N_23035);
nor UO_613 (O_613,N_22867,N_23340);
nor UO_614 (O_614,N_22285,N_22592);
nand UO_615 (O_615,N_22397,N_23461);
and UO_616 (O_616,N_23806,N_24545);
and UO_617 (O_617,N_24490,N_22110);
or UO_618 (O_618,N_22444,N_23710);
xnor UO_619 (O_619,N_23353,N_24565);
or UO_620 (O_620,N_24095,N_24768);
xnor UO_621 (O_621,N_23885,N_23911);
and UO_622 (O_622,N_22699,N_23799);
nor UO_623 (O_623,N_22364,N_22562);
nor UO_624 (O_624,N_22084,N_23697);
nor UO_625 (O_625,N_23021,N_23819);
nand UO_626 (O_626,N_24030,N_24191);
nor UO_627 (O_627,N_22814,N_22373);
and UO_628 (O_628,N_23835,N_23554);
or UO_629 (O_629,N_22939,N_24070);
xor UO_630 (O_630,N_23679,N_24856);
or UO_631 (O_631,N_23412,N_24074);
and UO_632 (O_632,N_23269,N_22037);
nand UO_633 (O_633,N_24254,N_24534);
or UO_634 (O_634,N_23846,N_22332);
nand UO_635 (O_635,N_22707,N_22461);
or UO_636 (O_636,N_23923,N_22269);
nand UO_637 (O_637,N_21939,N_22386);
nor UO_638 (O_638,N_22222,N_22291);
and UO_639 (O_639,N_23972,N_23621);
nand UO_640 (O_640,N_21907,N_23861);
nor UO_641 (O_641,N_24373,N_24929);
and UO_642 (O_642,N_22258,N_22858);
and UO_643 (O_643,N_23030,N_24942);
nand UO_644 (O_644,N_22836,N_24655);
and UO_645 (O_645,N_23672,N_22420);
and UO_646 (O_646,N_23405,N_24801);
and UO_647 (O_647,N_23364,N_22522);
nor UO_648 (O_648,N_24653,N_22191);
xor UO_649 (O_649,N_24893,N_23580);
and UO_650 (O_650,N_22523,N_24055);
xor UO_651 (O_651,N_23720,N_23953);
and UO_652 (O_652,N_21980,N_23856);
nand UO_653 (O_653,N_24274,N_23880);
or UO_654 (O_654,N_22903,N_24776);
nor UO_655 (O_655,N_24194,N_24376);
and UO_656 (O_656,N_22671,N_24535);
nor UO_657 (O_657,N_23107,N_23694);
or UO_658 (O_658,N_22214,N_24003);
nor UO_659 (O_659,N_24346,N_23839);
nor UO_660 (O_660,N_22579,N_23838);
nand UO_661 (O_661,N_24757,N_23485);
nor UO_662 (O_662,N_23609,N_23571);
nor UO_663 (O_663,N_23362,N_22598);
and UO_664 (O_664,N_23644,N_24631);
nand UO_665 (O_665,N_24747,N_22075);
nand UO_666 (O_666,N_21896,N_23658);
nand UO_667 (O_667,N_22302,N_24679);
or UO_668 (O_668,N_24013,N_21929);
nand UO_669 (O_669,N_22752,N_22876);
or UO_670 (O_670,N_22168,N_24222);
xor UO_671 (O_671,N_22228,N_23592);
nor UO_672 (O_672,N_24066,N_24021);
nand UO_673 (O_673,N_24501,N_24297);
and UO_674 (O_674,N_22429,N_24355);
nand UO_675 (O_675,N_22407,N_23183);
nor UO_676 (O_676,N_22757,N_24341);
nor UO_677 (O_677,N_24617,N_22785);
and UO_678 (O_678,N_22994,N_23264);
nand UO_679 (O_679,N_22353,N_21977);
or UO_680 (O_680,N_23289,N_24855);
or UO_681 (O_681,N_24164,N_22910);
and UO_682 (O_682,N_22498,N_23262);
or UO_683 (O_683,N_24224,N_23670);
and UO_684 (O_684,N_24644,N_22246);
nor UO_685 (O_685,N_23098,N_24528);
nand UO_686 (O_686,N_23447,N_22989);
xnor UO_687 (O_687,N_23243,N_23895);
nand UO_688 (O_688,N_23163,N_22658);
xor UO_689 (O_689,N_24877,N_24155);
nor UO_690 (O_690,N_24771,N_22221);
nor UO_691 (O_691,N_24278,N_22091);
and UO_692 (O_692,N_23690,N_22039);
nand UO_693 (O_693,N_23541,N_23057);
nor UO_694 (O_694,N_24667,N_22728);
or UO_695 (O_695,N_23603,N_22887);
or UO_696 (O_696,N_21916,N_24379);
xnor UO_697 (O_697,N_24245,N_24252);
or UO_698 (O_698,N_23471,N_22751);
nor UO_699 (O_699,N_23298,N_24674);
nor UO_700 (O_700,N_22116,N_21987);
nor UO_701 (O_701,N_22935,N_23721);
and UO_702 (O_702,N_23698,N_22961);
nor UO_703 (O_703,N_24613,N_24871);
xor UO_704 (O_704,N_23127,N_22893);
and UO_705 (O_705,N_23676,N_22051);
and UO_706 (O_706,N_24731,N_24588);
nor UO_707 (O_707,N_24488,N_22268);
and UO_708 (O_708,N_24169,N_24841);
nor UO_709 (O_709,N_22213,N_22239);
and UO_710 (O_710,N_22036,N_22570);
nand UO_711 (O_711,N_22803,N_24739);
nand UO_712 (O_712,N_23863,N_22040);
and UO_713 (O_713,N_24911,N_23482);
nor UO_714 (O_714,N_24596,N_22436);
nand UO_715 (O_715,N_23138,N_24511);
xor UO_716 (O_716,N_23463,N_24480);
nand UO_717 (O_717,N_23984,N_23929);
and UO_718 (O_718,N_23310,N_22372);
nor UO_719 (O_719,N_22141,N_22272);
or UO_720 (O_720,N_23488,N_23142);
or UO_721 (O_721,N_22835,N_23372);
nor UO_722 (O_722,N_22166,N_21960);
xnor UO_723 (O_723,N_23440,N_23012);
nand UO_724 (O_724,N_22396,N_23363);
and UO_725 (O_725,N_24293,N_21970);
nand UO_726 (O_726,N_22593,N_23985);
nand UO_727 (O_727,N_24995,N_24181);
and UO_728 (O_728,N_22012,N_22186);
nor UO_729 (O_729,N_23996,N_22050);
nor UO_730 (O_730,N_22988,N_22114);
or UO_731 (O_731,N_23653,N_22145);
nand UO_732 (O_732,N_22550,N_23448);
nand UO_733 (O_733,N_22659,N_23143);
and UO_734 (O_734,N_24232,N_23256);
nand UO_735 (O_735,N_23976,N_22113);
and UO_736 (O_736,N_23716,N_24835);
nor UO_737 (O_737,N_23339,N_22838);
nand UO_738 (O_738,N_22792,N_24294);
or UO_739 (O_739,N_23156,N_24039);
or UO_740 (O_740,N_22693,N_24281);
and UO_741 (O_741,N_22849,N_23058);
and UO_742 (O_742,N_24202,N_24990);
xor UO_743 (O_743,N_23161,N_23556);
nor UO_744 (O_744,N_24084,N_21921);
nand UO_745 (O_745,N_22715,N_22575);
and UO_746 (O_746,N_22317,N_22308);
or UO_747 (O_747,N_23664,N_24584);
or UO_748 (O_748,N_22161,N_24858);
and UO_749 (O_749,N_23075,N_22991);
nor UO_750 (O_750,N_23033,N_23590);
and UO_751 (O_751,N_22762,N_24400);
or UO_752 (O_752,N_23548,N_23342);
or UO_753 (O_753,N_23468,N_22776);
xor UO_754 (O_754,N_23225,N_22557);
and UO_755 (O_755,N_24120,N_23435);
and UO_756 (O_756,N_21913,N_24844);
xor UO_757 (O_757,N_23270,N_24514);
nor UO_758 (O_758,N_23395,N_21971);
or UO_759 (O_759,N_22901,N_23169);
nor UO_760 (O_760,N_24848,N_23140);
nand UO_761 (O_761,N_22496,N_24447);
or UO_762 (O_762,N_22428,N_22044);
and UO_763 (O_763,N_22392,N_22028);
nor UO_764 (O_764,N_23671,N_24423);
xor UO_765 (O_765,N_22281,N_24507);
and UO_766 (O_766,N_22478,N_21982);
nor UO_767 (O_767,N_23226,N_21922);
or UO_768 (O_768,N_24015,N_24106);
or UO_769 (O_769,N_22974,N_22714);
or UO_770 (O_770,N_24808,N_24054);
xor UO_771 (O_771,N_24794,N_24646);
or UO_772 (O_772,N_22962,N_22442);
xor UO_773 (O_773,N_24042,N_22150);
or UO_774 (O_774,N_23789,N_22059);
xor UO_775 (O_775,N_23096,N_22103);
nor UO_776 (O_776,N_22026,N_24593);
nor UO_777 (O_777,N_22176,N_23375);
xnor UO_778 (O_778,N_24261,N_23464);
nand UO_779 (O_779,N_22513,N_23457);
or UO_780 (O_780,N_24847,N_22698);
or UO_781 (O_781,N_23006,N_22149);
and UO_782 (O_782,N_22977,N_22933);
nand UO_783 (O_783,N_23157,N_24962);
nor UO_784 (O_784,N_22642,N_22014);
xor UO_785 (O_785,N_24233,N_24800);
or UO_786 (O_786,N_24695,N_24684);
nand UO_787 (O_787,N_23442,N_23095);
and UO_788 (O_788,N_23430,N_23195);
nand UO_789 (O_789,N_23986,N_23736);
or UO_790 (O_790,N_24825,N_22347);
or UO_791 (O_791,N_22489,N_23414);
or UO_792 (O_792,N_23645,N_24142);
xor UO_793 (O_793,N_23422,N_23344);
nand UO_794 (O_794,N_23625,N_22981);
and UO_795 (O_795,N_22984,N_22108);
or UO_796 (O_796,N_22031,N_24284);
nand UO_797 (O_797,N_23196,N_22761);
or UO_798 (O_798,N_22951,N_24322);
or UO_799 (O_799,N_24216,N_24315);
nand UO_800 (O_800,N_22923,N_22992);
or UO_801 (O_801,N_23202,N_24388);
nor UO_802 (O_802,N_23432,N_22199);
and UO_803 (O_803,N_23734,N_24064);
nand UO_804 (O_804,N_23505,N_24116);
and UO_805 (O_805,N_22008,N_22120);
nor UO_806 (O_806,N_23052,N_24581);
xor UO_807 (O_807,N_22764,N_23657);
xor UO_808 (O_808,N_23038,N_22958);
xor UO_809 (O_809,N_22371,N_22745);
and UO_810 (O_810,N_24109,N_23744);
nor UO_811 (O_811,N_22233,N_23386);
and UO_812 (O_812,N_24931,N_24860);
or UO_813 (O_813,N_24143,N_23538);
or UO_814 (O_814,N_22736,N_23689);
nand UO_815 (O_815,N_24993,N_23449);
or UO_816 (O_816,N_23419,N_24889);
nor UO_817 (O_817,N_24826,N_22809);
and UO_818 (O_818,N_24549,N_23001);
and UO_819 (O_819,N_22450,N_23427);
nor UO_820 (O_820,N_24175,N_24575);
nor UO_821 (O_821,N_23937,N_24248);
xor UO_822 (O_822,N_24151,N_22398);
nor UO_823 (O_823,N_22724,N_23133);
or UO_824 (O_824,N_24051,N_22440);
xor UO_825 (O_825,N_23567,N_22795);
nand UO_826 (O_826,N_21935,N_24868);
or UO_827 (O_827,N_23071,N_23010);
or UO_828 (O_828,N_23358,N_23385);
and UO_829 (O_829,N_24689,N_24787);
nand UO_830 (O_830,N_22368,N_23111);
nor UO_831 (O_831,N_24336,N_24513);
nor UO_832 (O_832,N_21918,N_24197);
and UO_833 (O_833,N_21923,N_24035);
nand UO_834 (O_834,N_24908,N_23878);
nor UO_835 (O_835,N_24836,N_22746);
xnor UO_836 (O_836,N_23411,N_23843);
or UO_837 (O_837,N_24516,N_22330);
nor UO_838 (O_838,N_24788,N_22839);
nor UO_839 (O_839,N_22404,N_24256);
or UO_840 (O_840,N_22338,N_22282);
xnor UO_841 (O_841,N_24200,N_24665);
and UO_842 (O_842,N_23125,N_21879);
nand UO_843 (O_843,N_23085,N_23746);
nand UO_844 (O_844,N_24016,N_22594);
and UO_845 (O_845,N_21901,N_23684);
or UO_846 (O_846,N_24267,N_21903);
xnor UO_847 (O_847,N_22231,N_24997);
or UO_848 (O_848,N_24483,N_24071);
or UO_849 (O_849,N_24269,N_24936);
and UO_850 (O_850,N_24947,N_22735);
and UO_851 (O_851,N_22323,N_23682);
and UO_852 (O_852,N_23824,N_23531);
or UO_853 (O_853,N_22024,N_22684);
and UO_854 (O_854,N_21981,N_22146);
nor UO_855 (O_855,N_23337,N_24019);
and UO_856 (O_856,N_22774,N_22571);
or UO_857 (O_857,N_23017,N_22142);
xor UO_858 (O_858,N_24831,N_24526);
or UO_859 (O_859,N_23595,N_24525);
nand UO_860 (O_860,N_23597,N_24983);
and UO_861 (O_861,N_23301,N_22483);
and UO_862 (O_862,N_22198,N_23279);
nand UO_863 (O_863,N_23900,N_22712);
and UO_864 (O_864,N_22969,N_22374);
or UO_865 (O_865,N_21914,N_22033);
nand UO_866 (O_866,N_22909,N_23588);
nand UO_867 (O_867,N_24277,N_24166);
xnor UO_868 (O_868,N_24210,N_22342);
nand UO_869 (O_869,N_24727,N_24681);
or UO_870 (O_870,N_24172,N_24554);
or UO_871 (O_871,N_23166,N_24440);
and UO_872 (O_872,N_22035,N_22381);
nand UO_873 (O_873,N_23229,N_22584);
xor UO_874 (O_874,N_24869,N_24462);
nand UO_875 (O_875,N_23459,N_24509);
or UO_876 (O_876,N_23808,N_21941);
or UO_877 (O_877,N_22480,N_23290);
and UO_878 (O_878,N_22119,N_24038);
or UO_879 (O_879,N_24053,N_24711);
nor UO_880 (O_880,N_24954,N_22475);
or UO_881 (O_881,N_23540,N_24489);
nand UO_882 (O_882,N_24504,N_22252);
and UO_883 (O_883,N_22934,N_23632);
nand UO_884 (O_884,N_22964,N_24781);
nor UO_885 (O_885,N_23445,N_23034);
or UO_886 (O_886,N_21988,N_24950);
nand UO_887 (O_887,N_21991,N_21946);
or UO_888 (O_888,N_22822,N_23586);
xor UO_889 (O_889,N_23576,N_23596);
nand UO_890 (O_890,N_21910,N_22441);
or UO_891 (O_891,N_23695,N_24636);
and UO_892 (O_892,N_22230,N_24295);
xor UO_893 (O_893,N_22459,N_22088);
and UO_894 (O_894,N_24221,N_24926);
and UO_895 (O_895,N_22621,N_24061);
nand UO_896 (O_896,N_23958,N_23947);
and UO_897 (O_897,N_22170,N_22649);
xor UO_898 (O_898,N_24829,N_22833);
and UO_899 (O_899,N_23399,N_23827);
and UO_900 (O_900,N_24351,N_22578);
xnor UO_901 (O_901,N_23917,N_23441);
nor UO_902 (O_902,N_22540,N_22073);
xor UO_903 (O_903,N_23174,N_23314);
xnor UO_904 (O_904,N_24955,N_23563);
nor UO_905 (O_905,N_24078,N_23887);
nand UO_906 (O_906,N_23293,N_23496);
or UO_907 (O_907,N_24391,N_22842);
nand UO_908 (O_908,N_23200,N_21947);
nor UO_909 (O_909,N_23275,N_21881);
nand UO_910 (O_910,N_22117,N_22211);
nor UO_911 (O_911,N_24145,N_22032);
and UO_912 (O_912,N_22382,N_22133);
nor UO_913 (O_913,N_24830,N_23374);
and UO_914 (O_914,N_24939,N_23281);
nor UO_915 (O_915,N_23977,N_23246);
or UO_916 (O_916,N_24786,N_23185);
or UO_917 (O_917,N_23120,N_24263);
nor UO_918 (O_918,N_22843,N_22339);
nand UO_919 (O_919,N_23849,N_24970);
nor UO_920 (O_920,N_23282,N_22976);
xor UO_921 (O_921,N_24179,N_24572);
nand UO_922 (O_922,N_22629,N_23373);
and UO_923 (O_923,N_23086,N_22257);
xnor UO_924 (O_924,N_24510,N_24645);
xor UO_925 (O_925,N_23428,N_23426);
nand UO_926 (O_926,N_24132,N_24580);
and UO_927 (O_927,N_23265,N_22913);
and UO_928 (O_928,N_23073,N_23059);
and UO_929 (O_929,N_22782,N_24570);
nor UO_930 (O_930,N_22905,N_23713);
or UO_931 (O_931,N_22788,N_22087);
nand UO_932 (O_932,N_22326,N_24296);
nor UO_933 (O_933,N_22310,N_22295);
or UO_934 (O_934,N_22356,N_22978);
and UO_935 (O_935,N_23757,N_22466);
or UO_936 (O_936,N_22733,N_24813);
nor UO_937 (O_937,N_23313,N_22101);
and UO_938 (O_938,N_22763,N_24828);
or UO_939 (O_939,N_22247,N_22304);
and UO_940 (O_940,N_22541,N_23131);
or UO_941 (O_941,N_24560,N_23669);
nand UO_942 (O_942,N_22898,N_23276);
xor UO_943 (O_943,N_24541,N_24231);
nor UO_944 (O_944,N_22987,N_22286);
or UO_945 (O_945,N_22401,N_23975);
xnor UO_946 (O_946,N_23477,N_23514);
nor UO_947 (O_947,N_23745,N_24161);
nor UO_948 (O_948,N_24612,N_22874);
and UO_949 (O_949,N_22576,N_23216);
nor UO_950 (O_950,N_23699,N_24652);
or UO_951 (O_951,N_23020,N_22956);
or UO_952 (O_952,N_22465,N_24941);
or UO_953 (O_953,N_24468,N_23239);
xnor UO_954 (O_954,N_23631,N_21911);
or UO_955 (O_955,N_22920,N_23055);
or UO_956 (O_956,N_24370,N_22068);
or UO_957 (O_957,N_21940,N_24371);
or UO_958 (O_958,N_23356,N_23747);
nand UO_959 (O_959,N_23779,N_24738);
nand UO_960 (O_960,N_23311,N_24493);
or UO_961 (O_961,N_24601,N_22298);
and UO_962 (O_962,N_24673,N_22153);
nand UO_963 (O_963,N_23338,N_24253);
and UO_964 (O_964,N_22053,N_23500);
nand UO_965 (O_965,N_24073,N_22603);
nor UO_966 (O_966,N_24363,N_22079);
nand UO_967 (O_967,N_23467,N_23965);
and UO_968 (O_968,N_23794,N_24883);
nand UO_969 (O_969,N_24900,N_24875);
and UO_970 (O_970,N_23470,N_23817);
nand UO_971 (O_971,N_24682,N_24359);
and UO_972 (O_972,N_23323,N_24823);
nor UO_973 (O_973,N_22993,N_22139);
xor UO_974 (O_974,N_23188,N_24937);
and UO_975 (O_975,N_22408,N_23674);
or UO_976 (O_976,N_24521,N_22447);
nor UO_977 (O_977,N_22412,N_24170);
or UO_978 (O_978,N_22206,N_23536);
nor UO_979 (O_979,N_22062,N_22665);
and UO_980 (O_980,N_22617,N_24112);
nor UO_981 (O_981,N_23718,N_22954);
and UO_982 (O_982,N_23738,N_21972);
or UO_983 (O_983,N_22777,N_23930);
nand UO_984 (O_984,N_22948,N_22770);
nor UO_985 (O_985,N_24238,N_22798);
nand UO_986 (O_986,N_22637,N_23242);
or UO_987 (O_987,N_22154,N_21899);
xnor UO_988 (O_988,N_23650,N_24722);
and UO_989 (O_989,N_24567,N_21875);
or UO_990 (O_990,N_22476,N_24783);
xor UO_991 (O_991,N_23703,N_23546);
and UO_992 (O_992,N_24047,N_24686);
and UO_993 (O_993,N_24177,N_24595);
nand UO_994 (O_994,N_22890,N_24985);
or UO_995 (O_995,N_23925,N_23074);
and UO_996 (O_996,N_24966,N_24802);
and UO_997 (O_997,N_24426,N_22202);
nand UO_998 (O_998,N_24101,N_22082);
or UO_999 (O_999,N_22815,N_22474);
nand UO_1000 (O_1000,N_23322,N_23008);
and UO_1001 (O_1001,N_23036,N_22796);
nor UO_1002 (O_1002,N_23032,N_23553);
nor UO_1003 (O_1003,N_24340,N_22912);
and UO_1004 (O_1004,N_23515,N_24755);
nand UO_1005 (O_1005,N_23902,N_23397);
or UO_1006 (O_1006,N_24707,N_23283);
nor UO_1007 (O_1007,N_23350,N_23754);
or UO_1008 (O_1008,N_24699,N_23233);
and UO_1009 (O_1009,N_23862,N_22034);
nor UO_1010 (O_1010,N_22931,N_23312);
nand UO_1011 (O_1011,N_23062,N_23177);
or UO_1012 (O_1012,N_22121,N_22443);
nor UO_1013 (O_1013,N_23578,N_23934);
nor UO_1014 (O_1014,N_21905,N_23410);
nand UO_1015 (O_1015,N_23167,N_23149);
and UO_1016 (O_1016,N_24105,N_24449);
or UO_1017 (O_1017,N_24923,N_22808);
and UO_1018 (O_1018,N_22535,N_24934);
and UO_1019 (O_1019,N_23130,N_24967);
or UO_1020 (O_1020,N_23499,N_22148);
nand UO_1021 (O_1021,N_22791,N_22615);
nand UO_1022 (O_1022,N_24299,N_24251);
or UO_1023 (O_1023,N_22296,N_22144);
nand UO_1024 (O_1024,N_24817,N_24149);
nor UO_1025 (O_1025,N_23922,N_24790);
and UO_1026 (O_1026,N_24675,N_24417);
and UO_1027 (O_1027,N_24717,N_23408);
and UO_1028 (O_1028,N_24012,N_24506);
nand UO_1029 (O_1029,N_24227,N_23800);
nor UO_1030 (O_1030,N_22568,N_24352);
or UO_1031 (O_1031,N_24334,N_22197);
or UO_1032 (O_1032,N_24849,N_22565);
nor UO_1033 (O_1033,N_22300,N_22739);
nand UO_1034 (O_1034,N_23197,N_22521);
xor UO_1035 (O_1035,N_22793,N_24758);
xor UO_1036 (O_1036,N_24387,N_22755);
nor UO_1037 (O_1037,N_24980,N_23700);
and UO_1038 (O_1038,N_22604,N_23502);
or UO_1039 (O_1039,N_23136,N_24789);
and UO_1040 (O_1040,N_23116,N_22700);
or UO_1041 (O_1041,N_24762,N_23189);
xor UO_1042 (O_1042,N_22423,N_24552);
and UO_1043 (O_1043,N_23347,N_24159);
and UO_1044 (O_1044,N_21996,N_24765);
or UO_1045 (O_1045,N_24843,N_22766);
nand UO_1046 (O_1046,N_24988,N_23760);
nand UO_1047 (O_1047,N_23892,N_24819);
nor UO_1048 (O_1048,N_22990,N_24205);
xor UO_1049 (O_1049,N_24649,N_24118);
and UO_1050 (O_1050,N_24518,N_24706);
nor UO_1051 (O_1051,N_24961,N_24872);
nor UO_1052 (O_1052,N_22686,N_24135);
or UO_1053 (O_1053,N_23171,N_22530);
nand UO_1054 (O_1054,N_24996,N_22963);
nor UO_1055 (O_1055,N_22046,N_24399);
nand UO_1056 (O_1056,N_24700,N_23945);
xor UO_1057 (O_1057,N_23109,N_21984);
nor UO_1058 (O_1058,N_24090,N_22284);
nor UO_1059 (O_1059,N_24930,N_24067);
xnor UO_1060 (O_1060,N_22940,N_22217);
nor UO_1061 (O_1061,N_22753,N_21895);
or UO_1062 (O_1062,N_22437,N_22647);
nand UO_1063 (O_1063,N_24517,N_24608);
or UO_1064 (O_1064,N_23859,N_22083);
xnor UO_1065 (O_1065,N_22680,N_24193);
nor UO_1066 (O_1066,N_23320,N_23547);
xnor UO_1067 (O_1067,N_22306,N_22626);
nor UO_1068 (O_1068,N_24140,N_24165);
xnor UO_1069 (O_1069,N_23014,N_24327);
nand UO_1070 (O_1070,N_23387,N_22456);
nor UO_1071 (O_1071,N_24305,N_22224);
or UO_1072 (O_1072,N_22528,N_22580);
nor UO_1073 (O_1073,N_23336,N_21963);
and UO_1074 (O_1074,N_22646,N_23466);
and UO_1075 (O_1075,N_21908,N_22552);
xor UO_1076 (O_1076,N_24187,N_24424);
or UO_1077 (O_1077,N_22744,N_24697);
xor UO_1078 (O_1078,N_22825,N_23206);
and UO_1079 (O_1079,N_24640,N_24246);
nand UO_1080 (O_1080,N_22543,N_22007);
nand UO_1081 (O_1081,N_23099,N_23822);
nor UO_1082 (O_1082,N_23194,N_23614);
nand UO_1083 (O_1083,N_24396,N_23220);
nand UO_1084 (O_1084,N_23991,N_24206);
and UO_1085 (O_1085,N_23067,N_23475);
xor UO_1086 (O_1086,N_23752,N_22380);
or UO_1087 (O_1087,N_24896,N_22789);
or UO_1088 (O_1088,N_23277,N_24989);
nor UO_1089 (O_1089,N_23403,N_24386);
nor UO_1090 (O_1090,N_22054,N_24749);
nand UO_1091 (O_1091,N_23688,N_24672);
xnor UO_1092 (O_1092,N_24332,N_22131);
nor UO_1093 (O_1093,N_22179,N_23790);
nand UO_1094 (O_1094,N_22417,N_21962);
or UO_1095 (O_1095,N_23139,N_23537);
nand UO_1096 (O_1096,N_22634,N_24479);
nand UO_1097 (O_1097,N_22134,N_24146);
and UO_1098 (O_1098,N_24903,N_24374);
nand UO_1099 (O_1099,N_24583,N_23192);
or UO_1100 (O_1100,N_22807,N_23388);
nor UO_1101 (O_1101,N_24861,N_22399);
nor UO_1102 (O_1102,N_21906,N_23764);
nor UO_1103 (O_1103,N_23687,N_22773);
or UO_1104 (O_1104,N_22515,N_23513);
and UO_1105 (O_1105,N_24056,N_22471);
and UO_1106 (O_1106,N_22261,N_22737);
and UO_1107 (O_1107,N_22413,N_22595);
or UO_1108 (O_1108,N_24469,N_22274);
xnor UO_1109 (O_1109,N_24441,N_22360);
nand UO_1110 (O_1110,N_24454,N_24751);
nand UO_1111 (O_1111,N_22881,N_23404);
xnor UO_1112 (O_1112,N_24804,N_22519);
or UO_1113 (O_1113,N_24973,N_24986);
nor UO_1114 (O_1114,N_24767,N_22361);
and UO_1115 (O_1115,N_24965,N_23848);
nand UO_1116 (O_1116,N_22690,N_22015);
nand UO_1117 (O_1117,N_23151,N_24862);
nand UO_1118 (O_1118,N_22692,N_23979);
and UO_1119 (O_1119,N_24725,N_24249);
nand UO_1120 (O_1120,N_23607,N_22180);
nor UO_1121 (O_1121,N_22343,N_24081);
nand UO_1122 (O_1122,N_23692,N_23854);
or UO_1123 (O_1123,N_23088,N_24498);
xor UO_1124 (O_1124,N_22017,N_24928);
nor UO_1125 (O_1125,N_24568,N_24398);
or UO_1126 (O_1126,N_21934,N_24304);
nand UO_1127 (O_1127,N_24380,N_24087);
xnor UO_1128 (O_1128,N_24530,N_23392);
or UO_1129 (O_1129,N_23333,N_23740);
or UO_1130 (O_1130,N_21885,N_24548);
nand UO_1131 (O_1131,N_23952,N_22503);
and UO_1132 (O_1132,N_22960,N_22899);
or UO_1133 (O_1133,N_21952,N_22856);
nor UO_1134 (O_1134,N_24234,N_23208);
nor UO_1135 (O_1135,N_24816,N_22355);
and UO_1136 (O_1136,N_23701,N_23302);
nand UO_1137 (O_1137,N_24080,N_24220);
or UO_1138 (O_1138,N_21945,N_22184);
and UO_1139 (O_1139,N_24152,N_24624);
nor UO_1140 (O_1140,N_23868,N_24812);
nor UO_1141 (O_1141,N_22884,N_22674);
and UO_1142 (O_1142,N_22463,N_23465);
and UO_1143 (O_1143,N_24614,N_23474);
nand UO_1144 (O_1144,N_23755,N_24882);
and UO_1145 (O_1145,N_22786,N_23659);
or UO_1146 (O_1146,N_24796,N_23504);
xor UO_1147 (O_1147,N_24453,N_24460);
nand UO_1148 (O_1148,N_22872,N_23476);
nand UO_1149 (O_1149,N_23325,N_23654);
nor UO_1150 (O_1150,N_24666,N_24874);
or UO_1151 (O_1151,N_22848,N_22608);
nor UO_1152 (O_1152,N_24422,N_23960);
or UO_1153 (O_1153,N_23420,N_23769);
nor UO_1154 (O_1154,N_23402,N_22467);
nand UO_1155 (O_1155,N_22076,N_22695);
and UO_1156 (O_1156,N_22906,N_23982);
nor UO_1157 (O_1157,N_24650,N_23492);
nor UO_1158 (O_1158,N_24904,N_24384);
and UO_1159 (O_1159,N_22192,N_22549);
and UO_1160 (O_1160,N_23791,N_24538);
nor UO_1161 (O_1161,N_23186,N_24034);
nand UO_1162 (O_1162,N_22346,N_23628);
nand UO_1163 (O_1163,N_22237,N_22628);
or UO_1164 (O_1164,N_22740,N_23472);
nor UO_1165 (O_1165,N_22952,N_24036);
nor UO_1166 (O_1166,N_22215,N_24144);
and UO_1167 (O_1167,N_24656,N_23175);
or UO_1168 (O_1168,N_22826,N_23382);
or UO_1169 (O_1169,N_23162,N_22544);
and UO_1170 (O_1170,N_23097,N_24104);
or UO_1171 (O_1171,N_22818,N_23315);
nand UO_1172 (O_1172,N_24972,N_23693);
nand UO_1173 (O_1173,N_24085,N_22387);
nor UO_1174 (O_1174,N_22251,N_24885);
or UO_1175 (O_1175,N_23155,N_22359);
nand UO_1176 (O_1176,N_24551,N_23647);
and UO_1177 (O_1177,N_24343,N_21930);
or UO_1178 (O_1178,N_24527,N_22307);
nor UO_1179 (O_1179,N_24137,N_23286);
and UO_1180 (O_1180,N_24974,N_23144);
xnor UO_1181 (O_1181,N_21968,N_22970);
nand UO_1182 (O_1182,N_22267,N_21961);
xor UO_1183 (O_1183,N_22280,N_23516);
nor UO_1184 (O_1184,N_22468,N_22688);
or UO_1185 (O_1185,N_24566,N_22609);
nor UO_1186 (O_1186,N_24348,N_23509);
nor UO_1187 (O_1187,N_23908,N_23584);
or UO_1188 (O_1188,N_24475,N_22804);
xor UO_1189 (O_1189,N_22098,N_22301);
nand UO_1190 (O_1190,N_22653,N_23706);
and UO_1191 (O_1191,N_24969,N_23436);
nor UO_1192 (O_1192,N_24357,N_22630);
nor UO_1193 (O_1193,N_22452,N_23089);
nand UO_1194 (O_1194,N_23433,N_22827);
and UO_1195 (O_1195,N_22512,N_23152);
nor UO_1196 (O_1196,N_24557,N_23572);
nand UO_1197 (O_1197,N_24414,N_24262);
xnor UO_1198 (O_1198,N_23316,N_22294);
or UO_1199 (O_1199,N_24218,N_24037);
or UO_1200 (O_1200,N_23237,N_23882);
nand UO_1201 (O_1201,N_24626,N_22577);
and UO_1202 (O_1202,N_24192,N_23454);
or UO_1203 (O_1203,N_22502,N_23560);
and UO_1204 (O_1204,N_23431,N_23629);
nor UO_1205 (O_1205,N_23160,N_23901);
and UO_1206 (O_1206,N_22780,N_22889);
or UO_1207 (O_1207,N_24338,N_23828);
nand UO_1208 (O_1208,N_24651,N_24754);
nor UO_1209 (O_1209,N_23303,N_22968);
or UO_1210 (O_1210,N_23907,N_23766);
and UO_1211 (O_1211,N_24512,N_24339);
nand UO_1212 (O_1212,N_22016,N_24126);
xnor UO_1213 (O_1213,N_23618,N_23587);
or UO_1214 (O_1214,N_22676,N_24467);
nor UO_1215 (O_1215,N_22632,N_24413);
or UO_1216 (O_1216,N_22556,N_23113);
nor UO_1217 (O_1217,N_22193,N_22625);
nor UO_1218 (O_1218,N_22574,N_24897);
nand UO_1219 (O_1219,N_22414,N_21954);
and UO_1220 (O_1220,N_23788,N_24029);
nand UO_1221 (O_1221,N_23636,N_22336);
nor UO_1222 (O_1222,N_22861,N_24680);
and UO_1223 (O_1223,N_23444,N_22107);
and UO_1224 (O_1224,N_24283,N_24115);
nand UO_1225 (O_1225,N_23612,N_24850);
nor UO_1226 (O_1226,N_24906,N_23948);
xor UO_1227 (O_1227,N_22949,N_23992);
or UO_1228 (O_1228,N_23570,N_23634);
nand UO_1229 (O_1229,N_22957,N_22516);
or UO_1230 (O_1230,N_23841,N_24558);
nor UO_1231 (O_1231,N_23761,N_23624);
or UO_1232 (O_1232,N_22596,N_24266);
or UO_1233 (O_1233,N_22946,N_24746);
nand UO_1234 (O_1234,N_23228,N_22312);
and UO_1235 (O_1235,N_24598,N_23950);
or UO_1236 (O_1236,N_22271,N_23883);
and UO_1237 (O_1237,N_24641,N_23793);
nor UO_1238 (O_1238,N_22612,N_21877);
nor UO_1239 (O_1239,N_24935,N_21937);
and UO_1240 (O_1240,N_24372,N_24932);
and UO_1241 (O_1241,N_24127,N_21884);
nor UO_1242 (O_1242,N_24272,N_23617);
or UO_1243 (O_1243,N_24845,N_24292);
or UO_1244 (O_1244,N_22425,N_22427);
or UO_1245 (O_1245,N_23919,N_22041);
xnor UO_1246 (O_1246,N_24001,N_23641);
nor UO_1247 (O_1247,N_22743,N_22102);
or UO_1248 (O_1248,N_23931,N_22327);
nor UO_1249 (O_1249,N_23964,N_24354);
nor UO_1250 (O_1250,N_24350,N_24658);
or UO_1251 (O_1251,N_23583,N_23640);
nor UO_1252 (O_1252,N_22995,N_23115);
or UO_1253 (O_1253,N_22462,N_24361);
or UO_1254 (O_1254,N_23763,N_23045);
or UO_1255 (O_1255,N_24079,N_23117);
xnor UO_1256 (O_1256,N_23954,N_23212);
and UO_1257 (O_1257,N_24615,N_23680);
nand UO_1258 (O_1258,N_23558,N_24756);
or UO_1259 (O_1259,N_24075,N_23480);
or UO_1260 (O_1260,N_24217,N_22105);
nand UO_1261 (O_1261,N_22943,N_22687);
or UO_1262 (O_1262,N_22566,N_23124);
xnor UO_1263 (O_1263,N_22156,N_24099);
nor UO_1264 (O_1264,N_22879,N_22409);
or UO_1265 (O_1265,N_22449,N_24603);
or UO_1266 (O_1266,N_22074,N_24133);
nand UO_1267 (O_1267,N_23158,N_22218);
nand UO_1268 (O_1268,N_22262,N_23104);
nor UO_1269 (O_1269,N_23557,N_23599);
and UO_1270 (O_1270,N_22917,N_23905);
nand UO_1271 (O_1271,N_22127,N_24837);
nand UO_1272 (O_1272,N_24157,N_24676);
nor UO_1273 (O_1273,N_22152,N_23122);
nor UO_1274 (O_1274,N_22136,N_22488);
and UO_1275 (O_1275,N_24282,N_24096);
or UO_1276 (O_1276,N_22000,N_23549);
nor UO_1277 (O_1277,N_21976,N_24213);
nand UO_1278 (O_1278,N_21944,N_24383);
xor UO_1279 (O_1279,N_24729,N_22055);
and UO_1280 (O_1280,N_23308,N_22896);
nor UO_1281 (O_1281,N_23346,N_22851);
and UO_1282 (O_1282,N_24302,N_23813);
xnor UO_1283 (O_1283,N_24418,N_22345);
or UO_1284 (O_1284,N_24873,N_23685);
nand UO_1285 (O_1285,N_24317,N_22389);
nand UO_1286 (O_1286,N_23438,N_21894);
or UO_1287 (O_1287,N_23415,N_23879);
or UO_1288 (O_1288,N_23899,N_22860);
and UO_1289 (O_1289,N_22445,N_24082);
xor UO_1290 (O_1290,N_24663,N_23884);
nand UO_1291 (O_1291,N_24891,N_22128);
or UO_1292 (O_1292,N_22064,N_22547);
xnor UO_1293 (O_1293,N_22357,N_23870);
nand UO_1294 (O_1294,N_23091,N_22925);
and UO_1295 (O_1295,N_22869,N_22061);
nor UO_1296 (O_1296,N_24735,N_22278);
nand UO_1297 (O_1297,N_22648,N_21931);
and UO_1298 (O_1298,N_23292,N_22854);
nor UO_1299 (O_1299,N_22203,N_23875);
nor UO_1300 (O_1300,N_23798,N_22369);
or UO_1301 (O_1301,N_24838,N_22875);
and UO_1302 (O_1302,N_23730,N_24102);
nor UO_1303 (O_1303,N_24154,N_23304);
and UO_1304 (O_1304,N_23655,N_24502);
or UO_1305 (O_1305,N_24419,N_23753);
nor UO_1306 (O_1306,N_23361,N_22947);
and UO_1307 (O_1307,N_23811,N_22491);
nand UO_1308 (O_1308,N_24463,N_22747);
nor UO_1309 (O_1309,N_23577,N_24664);
or UO_1310 (O_1310,N_23714,N_21959);
or UO_1311 (O_1311,N_22801,N_23065);
nand UO_1312 (O_1312,N_24291,N_23853);
nor UO_1313 (O_1313,N_22542,N_22422);
or UO_1314 (O_1314,N_23063,N_23128);
or UO_1315 (O_1315,N_22027,N_23181);
and UO_1316 (O_1316,N_22004,N_24610);
nor UO_1317 (O_1317,N_22871,N_23795);
nor UO_1318 (O_1318,N_23193,N_23840);
and UO_1319 (O_1319,N_22481,N_22748);
or UO_1320 (O_1320,N_23029,N_24028);
or UO_1321 (O_1321,N_23589,N_24235);
nor UO_1322 (O_1322,N_22201,N_22850);
or UO_1323 (O_1323,N_22679,N_21993);
nor UO_1324 (O_1324,N_24778,N_22270);
or UO_1325 (O_1325,N_24482,N_24032);
or UO_1326 (O_1326,N_24307,N_21989);
and UO_1327 (O_1327,N_23552,N_24225);
and UO_1328 (O_1328,N_22810,N_22667);
nor UO_1329 (O_1329,N_24366,N_23238);
nand UO_1330 (O_1330,N_22967,N_23355);
nand UO_1331 (O_1331,N_21995,N_24515);
and UO_1332 (O_1332,N_22479,N_24203);
and UO_1333 (O_1333,N_22453,N_23775);
nor UO_1334 (O_1334,N_23725,N_24834);
nand UO_1335 (O_1335,N_24360,N_23083);
and UO_1336 (O_1336,N_22790,N_22696);
nor UO_1337 (O_1337,N_24497,N_24123);
xor UO_1338 (O_1338,N_24892,N_23335);
nor UO_1339 (O_1339,N_24870,N_23494);
or UO_1340 (O_1340,N_22472,N_23207);
nor UO_1341 (O_1341,N_23224,N_22325);
xnor UO_1342 (O_1342,N_22354,N_22132);
or UO_1343 (O_1343,N_23377,N_24563);
nand UO_1344 (O_1344,N_23254,N_24046);
nand UO_1345 (O_1345,N_24329,N_24180);
xor UO_1346 (O_1346,N_24401,N_23093);
nand UO_1347 (O_1347,N_24148,N_22490);
and UO_1348 (O_1348,N_23527,N_22341);
or UO_1349 (O_1349,N_24188,N_24547);
or UO_1350 (O_1350,N_23173,N_22731);
nor UO_1351 (O_1351,N_22042,N_22358);
nor UO_1352 (O_1352,N_22971,N_22321);
and UO_1353 (O_1353,N_22421,N_23064);
nor UO_1354 (O_1354,N_22097,N_23918);
nand UO_1355 (O_1355,N_22029,N_22725);
nand UO_1356 (O_1356,N_24393,N_24508);
nand UO_1357 (O_1357,N_23473,N_22902);
and UO_1358 (O_1358,N_23735,N_24026);
nand UO_1359 (O_1359,N_23296,N_22820);
or UO_1360 (O_1360,N_22350,N_22741);
xor UO_1361 (O_1361,N_24791,N_23245);
nand UO_1362 (O_1362,N_24409,N_22010);
and UO_1363 (O_1363,N_23770,N_23830);
nand UO_1364 (O_1364,N_24110,N_23129);
nand UO_1365 (O_1365,N_24103,N_23562);
nand UO_1366 (O_1366,N_24594,N_22610);
or UO_1367 (O_1367,N_23022,N_22919);
nor UO_1368 (O_1368,N_24326,N_24389);
nor UO_1369 (O_1369,N_24720,N_23341);
xor UO_1370 (O_1370,N_24987,N_23126);
or UO_1371 (O_1371,N_23564,N_23651);
xnor UO_1372 (O_1372,N_24324,N_23077);
nand UO_1373 (O_1373,N_24839,N_23816);
nor UO_1374 (O_1374,N_24345,N_24069);
and UO_1375 (O_1375,N_23712,N_22911);
nand UO_1376 (O_1376,N_22238,N_22391);
or UO_1377 (O_1377,N_22265,N_22477);
or UO_1378 (O_1378,N_21965,N_24171);
nand UO_1379 (O_1379,N_24319,N_24450);
nand UO_1380 (O_1380,N_23959,N_22953);
nor UO_1381 (O_1381,N_23904,N_22340);
xnor UO_1382 (O_1382,N_22870,N_24992);
nand UO_1383 (O_1383,N_23534,N_24000);
xnor UO_1384 (O_1384,N_22563,N_22143);
or UO_1385 (O_1385,N_22581,N_23330);
and UO_1386 (O_1386,N_22431,N_24499);
or UO_1387 (O_1387,N_22852,N_22318);
and UO_1388 (O_1388,N_22277,N_24846);
nand UO_1389 (O_1389,N_24886,N_23519);
nor UO_1390 (O_1390,N_24223,N_22492);
or UO_1391 (O_1391,N_22817,N_24971);
or UO_1392 (O_1392,N_22738,N_24113);
nor UO_1393 (O_1393,N_24660,N_22426);
nand UO_1394 (O_1394,N_22283,N_22710);
or UO_1395 (O_1395,N_22526,N_24721);
and UO_1396 (O_1396,N_23334,N_23804);
or UO_1397 (O_1397,N_23681,N_23637);
and UO_1398 (O_1398,N_22533,N_22172);
nand UO_1399 (O_1399,N_23253,N_23623);
xnor UO_1400 (O_1400,N_23252,N_24605);
or UO_1401 (O_1401,N_24999,N_24316);
and UO_1402 (O_1402,N_22366,N_23675);
and UO_1403 (O_1403,N_24698,N_23635);
and UO_1404 (O_1404,N_24687,N_23967);
nor UO_1405 (O_1405,N_23535,N_24496);
nand UO_1406 (O_1406,N_22507,N_22049);
nand UO_1407 (O_1407,N_24403,N_23092);
or UO_1408 (O_1408,N_24392,N_23478);
nor UO_1409 (O_1409,N_23199,N_22928);
and UO_1410 (O_1410,N_22279,N_23909);
xnor UO_1411 (O_1411,N_24633,N_22118);
nand UO_1412 (O_1412,N_24043,N_22209);
nor UO_1413 (O_1413,N_23921,N_22446);
and UO_1414 (O_1414,N_22365,N_22129);
and UO_1415 (O_1415,N_23005,N_23733);
xor UO_1416 (O_1416,N_24948,N_23891);
or UO_1417 (O_1417,N_24607,N_22510);
nand UO_1418 (O_1418,N_22719,N_22888);
and UO_1419 (O_1419,N_24086,N_22175);
and UO_1420 (O_1420,N_22086,N_22319);
or UO_1421 (O_1421,N_24741,N_24587);
and UO_1422 (O_1422,N_23219,N_22865);
and UO_1423 (O_1423,N_24854,N_23134);
nand UO_1424 (O_1424,N_21983,N_23910);
and UO_1425 (O_1425,N_22613,N_24894);
or UO_1426 (O_1426,N_23691,N_22190);
and UO_1427 (O_1427,N_22052,N_22588);
nor UO_1428 (O_1428,N_22344,N_23456);
and UO_1429 (O_1429,N_22207,N_24461);
or UO_1430 (O_1430,N_24290,N_22313);
nor UO_1431 (O_1431,N_22819,N_24060);
xnor UO_1432 (O_1432,N_23389,N_24432);
and UO_1433 (O_1433,N_22618,N_23622);
and UO_1434 (O_1434,N_22165,N_24390);
nand UO_1435 (O_1435,N_23711,N_23218);
or UO_1436 (O_1436,N_22223,N_23491);
or UO_1437 (O_1437,N_22732,N_22582);
and UO_1438 (O_1438,N_22711,N_23815);
nand UO_1439 (O_1439,N_23673,N_24763);
nor UO_1440 (O_1440,N_23154,N_23453);
or UO_1441 (O_1441,N_23369,N_23957);
and UO_1442 (O_1442,N_22160,N_22635);
nand UO_1443 (O_1443,N_23011,N_22402);
nor UO_1444 (O_1444,N_24718,N_24258);
or UO_1445 (O_1445,N_23876,N_24503);
and UO_1446 (O_1446,N_23051,N_23920);
or UO_1447 (O_1447,N_22095,N_24669);
and UO_1448 (O_1448,N_23040,N_24945);
or UO_1449 (O_1449,N_23777,N_22394);
and UO_1450 (O_1450,N_24121,N_22907);
nor UO_1451 (O_1451,N_22216,N_23581);
and UO_1452 (O_1452,N_23826,N_22701);
nor UO_1453 (O_1453,N_21979,N_22125);
nand UO_1454 (O_1454,N_23890,N_23418);
nand UO_1455 (O_1455,N_23319,N_23530);
nor UO_1456 (O_1456,N_23326,N_22314);
nor UO_1457 (O_1457,N_24186,N_23926);
nor UO_1458 (O_1458,N_22862,N_22720);
nand UO_1459 (O_1459,N_23009,N_24582);
and UO_1460 (O_1460,N_24888,N_23423);
nand UO_1461 (O_1461,N_23443,N_22253);
nor UO_1462 (O_1462,N_21904,N_22916);
and UO_1463 (O_1463,N_22567,N_24049);
nand UO_1464 (O_1464,N_22289,N_23610);
xnor UO_1465 (O_1465,N_23042,N_21973);
or UO_1466 (O_1466,N_21949,N_22855);
or UO_1467 (O_1467,N_23820,N_23683);
or UO_1468 (O_1468,N_22639,N_23600);
nand UO_1469 (O_1469,N_24005,N_23508);
xnor UO_1470 (O_1470,N_24429,N_23765);
nor UO_1471 (O_1471,N_24230,N_22942);
and UO_1472 (O_1472,N_23417,N_22260);
and UO_1473 (O_1473,N_21975,N_22525);
or UO_1474 (O_1474,N_22599,N_23620);
nor UO_1475 (O_1475,N_24710,N_22930);
and UO_1476 (O_1476,N_24183,N_23869);
nand UO_1477 (O_1477,N_23896,N_22109);
xnor UO_1478 (O_1478,N_22181,N_24670);
or UO_1479 (O_1479,N_22769,N_22834);
or UO_1480 (O_1480,N_22469,N_21890);
or UO_1481 (O_1481,N_22806,N_23148);
or UO_1482 (O_1482,N_24876,N_24093);
nand UO_1483 (O_1483,N_23517,N_23834);
nand UO_1484 (O_1484,N_23384,N_23916);
nand UO_1485 (O_1485,N_22729,N_24753);
and UO_1486 (O_1486,N_23709,N_21986);
nand UO_1487 (O_1487,N_23818,N_23767);
and UO_1488 (O_1488,N_22071,N_24130);
xor UO_1489 (O_1489,N_22750,N_23566);
nand UO_1490 (O_1490,N_22163,N_22439);
or UO_1491 (O_1491,N_24604,N_23105);
nor UO_1492 (O_1492,N_24286,N_23630);
nor UO_1493 (O_1493,N_24827,N_24907);
nand UO_1494 (O_1494,N_24408,N_23708);
or UO_1495 (O_1495,N_24323,N_22703);
nor UO_1496 (O_1496,N_22985,N_23069);
nand UO_1497 (O_1497,N_23078,N_22123);
and UO_1498 (O_1498,N_23255,N_24824);
xnor UO_1499 (O_1499,N_22266,N_24550);
or UO_1500 (O_1500,N_24692,N_23743);
nand UO_1501 (O_1501,N_23666,N_24270);
nand UO_1502 (O_1502,N_24562,N_22678);
or UO_1503 (O_1503,N_23187,N_22390);
nand UO_1504 (O_1504,N_21880,N_24579);
or UO_1505 (O_1505,N_22783,N_22627);
or UO_1506 (O_1506,N_22328,N_22315);
and UO_1507 (O_1507,N_22704,N_24574);
nor UO_1508 (O_1508,N_22587,N_23486);
nand UO_1509 (O_1509,N_22767,N_24709);
nand UO_1510 (O_1510,N_23871,N_23874);
nand UO_1511 (O_1511,N_23867,N_23066);
or UO_1512 (O_1512,N_24616,N_22537);
xnor UO_1513 (O_1513,N_23141,N_24899);
or UO_1514 (O_1514,N_23019,N_23380);
or UO_1515 (O_1515,N_23772,N_23359);
or UO_1516 (O_1516,N_23203,N_23963);
nand UO_1517 (O_1517,N_24378,N_22505);
nand UO_1518 (O_1518,N_23633,N_22070);
nor UO_1519 (O_1519,N_22633,N_23501);
and UO_1520 (O_1520,N_24257,N_22811);
and UO_1521 (O_1521,N_22950,N_23025);
and UO_1522 (O_1522,N_22377,N_22362);
or UO_1523 (O_1523,N_22406,N_23702);
nand UO_1524 (O_1524,N_22641,N_22561);
nand UO_1525 (O_1525,N_22115,N_23002);
or UO_1526 (O_1526,N_23215,N_21912);
nand UO_1527 (O_1527,N_23439,N_24909);
nand UO_1528 (O_1528,N_23222,N_24630);
nor UO_1529 (O_1529,N_23866,N_24724);
or UO_1530 (O_1530,N_24818,N_24884);
and UO_1531 (O_1531,N_23401,N_24402);
nand UO_1532 (O_1532,N_23877,N_22288);
and UO_1533 (O_1533,N_23642,N_22794);
nor UO_1534 (O_1534,N_24704,N_24011);
nor UO_1535 (O_1535,N_24638,N_23048);
nor UO_1536 (O_1536,N_24919,N_22473);
xnor UO_1537 (O_1537,N_24311,N_24737);
nand UO_1538 (O_1538,N_22723,N_22650);
xnor UO_1539 (O_1539,N_22320,N_23741);
or UO_1540 (O_1540,N_23750,N_24696);
nand UO_1541 (O_1541,N_23543,N_22564);
nor UO_1542 (O_1542,N_22067,N_21966);
nor UO_1543 (O_1543,N_24335,N_23082);
or UO_1544 (O_1544,N_24059,N_24244);
nand UO_1545 (O_1545,N_24833,N_24878);
and UO_1546 (O_1546,N_24425,N_23145);
and UO_1547 (O_1547,N_23306,N_22955);
nor UO_1548 (O_1548,N_24226,N_23172);
nor UO_1549 (O_1549,N_23080,N_23643);
nand UO_1550 (O_1550,N_23299,N_23294);
or UO_1551 (O_1551,N_24008,N_22096);
nand UO_1552 (O_1552,N_22844,N_23935);
xor UO_1553 (O_1553,N_24495,N_24321);
or UO_1554 (O_1554,N_23263,N_23132);
or UO_1555 (O_1555,N_24643,N_22331);
nor UO_1556 (O_1556,N_24793,N_23894);
nor UO_1557 (O_1557,N_21942,N_23178);
nand UO_1558 (O_1558,N_24368,N_23481);
nand UO_1559 (O_1559,N_23236,N_24524);
nand UO_1560 (O_1560,N_23054,N_24308);
and UO_1561 (O_1561,N_24020,N_21924);
nand UO_1562 (O_1562,N_22011,N_23214);
or UO_1563 (O_1563,N_22267,N_23454);
nand UO_1564 (O_1564,N_22381,N_22774);
nor UO_1565 (O_1565,N_24503,N_22162);
nand UO_1566 (O_1566,N_23559,N_22817);
and UO_1567 (O_1567,N_22367,N_22375);
nor UO_1568 (O_1568,N_23983,N_24490);
or UO_1569 (O_1569,N_23793,N_23441);
nand UO_1570 (O_1570,N_22027,N_23321);
nor UO_1571 (O_1571,N_24371,N_24737);
or UO_1572 (O_1572,N_24051,N_22802);
xor UO_1573 (O_1573,N_22357,N_23915);
nor UO_1574 (O_1574,N_23400,N_22659);
and UO_1575 (O_1575,N_24187,N_23593);
and UO_1576 (O_1576,N_24280,N_22089);
or UO_1577 (O_1577,N_23292,N_22395);
and UO_1578 (O_1578,N_24733,N_24583);
or UO_1579 (O_1579,N_24450,N_23361);
and UO_1580 (O_1580,N_23663,N_23556);
nand UO_1581 (O_1581,N_24319,N_21887);
and UO_1582 (O_1582,N_23457,N_23267);
nor UO_1583 (O_1583,N_23451,N_24865);
nor UO_1584 (O_1584,N_23949,N_24818);
or UO_1585 (O_1585,N_23442,N_23044);
and UO_1586 (O_1586,N_24051,N_21994);
nor UO_1587 (O_1587,N_24539,N_24383);
nand UO_1588 (O_1588,N_23282,N_23746);
nor UO_1589 (O_1589,N_22461,N_23242);
and UO_1590 (O_1590,N_23644,N_22748);
nor UO_1591 (O_1591,N_22068,N_24514);
nor UO_1592 (O_1592,N_24001,N_22771);
nand UO_1593 (O_1593,N_21935,N_22078);
or UO_1594 (O_1594,N_23582,N_24169);
or UO_1595 (O_1595,N_23307,N_22562);
and UO_1596 (O_1596,N_23128,N_23530);
nand UO_1597 (O_1597,N_22621,N_23268);
nor UO_1598 (O_1598,N_23425,N_22848);
nor UO_1599 (O_1599,N_23688,N_22363);
nor UO_1600 (O_1600,N_24290,N_23738);
xnor UO_1601 (O_1601,N_23254,N_24965);
or UO_1602 (O_1602,N_22102,N_24257);
or UO_1603 (O_1603,N_23639,N_23083);
nor UO_1604 (O_1604,N_23149,N_23152);
nor UO_1605 (O_1605,N_22736,N_24192);
and UO_1606 (O_1606,N_22658,N_24429);
nor UO_1607 (O_1607,N_24996,N_22673);
nor UO_1608 (O_1608,N_24001,N_23212);
and UO_1609 (O_1609,N_24030,N_22536);
or UO_1610 (O_1610,N_23428,N_23604);
and UO_1611 (O_1611,N_24580,N_23067);
nand UO_1612 (O_1612,N_22251,N_22021);
nand UO_1613 (O_1613,N_23881,N_24516);
nand UO_1614 (O_1614,N_22116,N_24099);
or UO_1615 (O_1615,N_22916,N_23495);
and UO_1616 (O_1616,N_22862,N_24264);
xnor UO_1617 (O_1617,N_22910,N_22390);
xnor UO_1618 (O_1618,N_22318,N_22730);
nand UO_1619 (O_1619,N_22447,N_24184);
and UO_1620 (O_1620,N_23899,N_23250);
or UO_1621 (O_1621,N_22843,N_22187);
nor UO_1622 (O_1622,N_24674,N_23829);
or UO_1623 (O_1623,N_23870,N_24359);
and UO_1624 (O_1624,N_23142,N_22448);
nor UO_1625 (O_1625,N_24568,N_24043);
or UO_1626 (O_1626,N_21906,N_22264);
and UO_1627 (O_1627,N_22887,N_23480);
or UO_1628 (O_1628,N_24954,N_22463);
nand UO_1629 (O_1629,N_22487,N_22913);
nor UO_1630 (O_1630,N_22886,N_23589);
nand UO_1631 (O_1631,N_22643,N_24063);
xnor UO_1632 (O_1632,N_22315,N_23017);
nand UO_1633 (O_1633,N_24707,N_22020);
nand UO_1634 (O_1634,N_23407,N_24431);
or UO_1635 (O_1635,N_22074,N_22867);
nor UO_1636 (O_1636,N_23847,N_23159);
nand UO_1637 (O_1637,N_23486,N_22478);
and UO_1638 (O_1638,N_22118,N_22545);
xor UO_1639 (O_1639,N_23323,N_24459);
and UO_1640 (O_1640,N_22921,N_24668);
xnor UO_1641 (O_1641,N_22229,N_23197);
nor UO_1642 (O_1642,N_24536,N_23673);
nor UO_1643 (O_1643,N_24614,N_21979);
and UO_1644 (O_1644,N_24758,N_22162);
nor UO_1645 (O_1645,N_24783,N_21911);
nor UO_1646 (O_1646,N_22714,N_23485);
xor UO_1647 (O_1647,N_23853,N_23156);
nand UO_1648 (O_1648,N_24523,N_22193);
nor UO_1649 (O_1649,N_24710,N_24700);
and UO_1650 (O_1650,N_22448,N_22791);
and UO_1651 (O_1651,N_23918,N_22621);
or UO_1652 (O_1652,N_24958,N_23297);
nand UO_1653 (O_1653,N_23320,N_22369);
nor UO_1654 (O_1654,N_24871,N_23646);
nor UO_1655 (O_1655,N_24799,N_24677);
nand UO_1656 (O_1656,N_22693,N_23365);
nor UO_1657 (O_1657,N_24226,N_23318);
or UO_1658 (O_1658,N_22417,N_23707);
and UO_1659 (O_1659,N_23702,N_24157);
nand UO_1660 (O_1660,N_22831,N_23207);
nand UO_1661 (O_1661,N_23903,N_23317);
or UO_1662 (O_1662,N_23570,N_24640);
nand UO_1663 (O_1663,N_24722,N_22792);
or UO_1664 (O_1664,N_24134,N_22787);
and UO_1665 (O_1665,N_24653,N_24364);
or UO_1666 (O_1666,N_23395,N_22860);
or UO_1667 (O_1667,N_22187,N_22269);
or UO_1668 (O_1668,N_23769,N_22116);
or UO_1669 (O_1669,N_24900,N_23871);
xor UO_1670 (O_1670,N_23013,N_24205);
or UO_1671 (O_1671,N_24950,N_23749);
xor UO_1672 (O_1672,N_23344,N_22645);
and UO_1673 (O_1673,N_22074,N_23209);
or UO_1674 (O_1674,N_24659,N_24777);
nor UO_1675 (O_1675,N_23608,N_22035);
xor UO_1676 (O_1676,N_22220,N_24266);
or UO_1677 (O_1677,N_23222,N_24523);
nand UO_1678 (O_1678,N_23742,N_23865);
nand UO_1679 (O_1679,N_23560,N_22120);
nand UO_1680 (O_1680,N_23212,N_23056);
nor UO_1681 (O_1681,N_23927,N_23469);
xnor UO_1682 (O_1682,N_22410,N_21951);
nor UO_1683 (O_1683,N_22229,N_23337);
nor UO_1684 (O_1684,N_21992,N_24985);
and UO_1685 (O_1685,N_22629,N_23413);
and UO_1686 (O_1686,N_23782,N_22757);
nor UO_1687 (O_1687,N_22900,N_23807);
or UO_1688 (O_1688,N_22550,N_23090);
nand UO_1689 (O_1689,N_24343,N_21937);
and UO_1690 (O_1690,N_22083,N_22903);
and UO_1691 (O_1691,N_24326,N_24837);
xor UO_1692 (O_1692,N_24711,N_24868);
nor UO_1693 (O_1693,N_23759,N_24313);
or UO_1694 (O_1694,N_22798,N_23639);
nor UO_1695 (O_1695,N_24944,N_22490);
nand UO_1696 (O_1696,N_23219,N_21959);
nor UO_1697 (O_1697,N_24672,N_23013);
nor UO_1698 (O_1698,N_24943,N_22873);
nand UO_1699 (O_1699,N_24330,N_22948);
nor UO_1700 (O_1700,N_23286,N_23509);
or UO_1701 (O_1701,N_24672,N_22037);
and UO_1702 (O_1702,N_22696,N_24564);
nor UO_1703 (O_1703,N_24425,N_24239);
nor UO_1704 (O_1704,N_22385,N_24336);
nand UO_1705 (O_1705,N_22873,N_22257);
or UO_1706 (O_1706,N_23278,N_23828);
nor UO_1707 (O_1707,N_21951,N_24769);
or UO_1708 (O_1708,N_22718,N_24794);
or UO_1709 (O_1709,N_22005,N_24122);
nor UO_1710 (O_1710,N_22585,N_22550);
or UO_1711 (O_1711,N_23698,N_23303);
or UO_1712 (O_1712,N_23642,N_22109);
and UO_1713 (O_1713,N_23318,N_23597);
and UO_1714 (O_1714,N_24018,N_24774);
and UO_1715 (O_1715,N_22168,N_24185);
nand UO_1716 (O_1716,N_22999,N_24059);
nor UO_1717 (O_1717,N_22184,N_23463);
or UO_1718 (O_1718,N_24987,N_23269);
nor UO_1719 (O_1719,N_22607,N_22149);
or UO_1720 (O_1720,N_22170,N_24943);
nor UO_1721 (O_1721,N_22823,N_22014);
nor UO_1722 (O_1722,N_24629,N_22017);
nor UO_1723 (O_1723,N_24318,N_24375);
or UO_1724 (O_1724,N_24590,N_22409);
nor UO_1725 (O_1725,N_23602,N_24112);
or UO_1726 (O_1726,N_24108,N_22393);
xor UO_1727 (O_1727,N_23822,N_24704);
and UO_1728 (O_1728,N_22185,N_24059);
or UO_1729 (O_1729,N_23773,N_24698);
nor UO_1730 (O_1730,N_23583,N_24765);
and UO_1731 (O_1731,N_21903,N_22444);
nor UO_1732 (O_1732,N_24235,N_24227);
nand UO_1733 (O_1733,N_22665,N_24712);
nand UO_1734 (O_1734,N_24591,N_24371);
or UO_1735 (O_1735,N_24629,N_22663);
or UO_1736 (O_1736,N_24302,N_24175);
and UO_1737 (O_1737,N_23033,N_22419);
nand UO_1738 (O_1738,N_24426,N_23521);
nor UO_1739 (O_1739,N_23319,N_23001);
or UO_1740 (O_1740,N_22759,N_24180);
or UO_1741 (O_1741,N_22985,N_24417);
and UO_1742 (O_1742,N_22136,N_24485);
xnor UO_1743 (O_1743,N_24406,N_23827);
xnor UO_1744 (O_1744,N_21918,N_23513);
nand UO_1745 (O_1745,N_21995,N_23822);
nor UO_1746 (O_1746,N_23625,N_23090);
nand UO_1747 (O_1747,N_24567,N_23198);
xor UO_1748 (O_1748,N_24035,N_23306);
or UO_1749 (O_1749,N_23686,N_23868);
or UO_1750 (O_1750,N_22116,N_24673);
nor UO_1751 (O_1751,N_24888,N_22979);
and UO_1752 (O_1752,N_22798,N_22575);
or UO_1753 (O_1753,N_24260,N_24758);
nor UO_1754 (O_1754,N_23494,N_24546);
or UO_1755 (O_1755,N_23943,N_23122);
xnor UO_1756 (O_1756,N_24242,N_24681);
nor UO_1757 (O_1757,N_24092,N_22979);
and UO_1758 (O_1758,N_21919,N_22014);
or UO_1759 (O_1759,N_23149,N_24457);
xor UO_1760 (O_1760,N_23574,N_23366);
and UO_1761 (O_1761,N_22730,N_23610);
and UO_1762 (O_1762,N_24659,N_23414);
and UO_1763 (O_1763,N_22439,N_23143);
nand UO_1764 (O_1764,N_23827,N_22072);
or UO_1765 (O_1765,N_24137,N_23587);
and UO_1766 (O_1766,N_23611,N_22290);
or UO_1767 (O_1767,N_24847,N_22842);
nand UO_1768 (O_1768,N_23193,N_24386);
or UO_1769 (O_1769,N_23675,N_23278);
nor UO_1770 (O_1770,N_22576,N_23057);
nand UO_1771 (O_1771,N_22387,N_23091);
nand UO_1772 (O_1772,N_22938,N_22697);
nor UO_1773 (O_1773,N_24579,N_22031);
or UO_1774 (O_1774,N_24712,N_24570);
and UO_1775 (O_1775,N_24775,N_23984);
xnor UO_1776 (O_1776,N_24132,N_22741);
nor UO_1777 (O_1777,N_24695,N_23524);
and UO_1778 (O_1778,N_22302,N_22690);
nor UO_1779 (O_1779,N_24302,N_23404);
xnor UO_1780 (O_1780,N_24141,N_22777);
or UO_1781 (O_1781,N_23416,N_23758);
and UO_1782 (O_1782,N_22161,N_22407);
or UO_1783 (O_1783,N_24060,N_24613);
and UO_1784 (O_1784,N_21948,N_24029);
or UO_1785 (O_1785,N_24422,N_23945);
and UO_1786 (O_1786,N_24372,N_23406);
or UO_1787 (O_1787,N_24920,N_22587);
xnor UO_1788 (O_1788,N_23132,N_23076);
nor UO_1789 (O_1789,N_22007,N_23835);
or UO_1790 (O_1790,N_22340,N_22508);
xnor UO_1791 (O_1791,N_24251,N_24260);
and UO_1792 (O_1792,N_24492,N_23657);
and UO_1793 (O_1793,N_23575,N_22725);
and UO_1794 (O_1794,N_23403,N_23499);
nor UO_1795 (O_1795,N_22334,N_24504);
nor UO_1796 (O_1796,N_24316,N_23975);
and UO_1797 (O_1797,N_22167,N_24098);
and UO_1798 (O_1798,N_24053,N_24222);
nand UO_1799 (O_1799,N_22624,N_21896);
and UO_1800 (O_1800,N_21999,N_22202);
nand UO_1801 (O_1801,N_22713,N_22022);
and UO_1802 (O_1802,N_23145,N_24874);
nand UO_1803 (O_1803,N_22153,N_23326);
nand UO_1804 (O_1804,N_22820,N_24718);
xnor UO_1805 (O_1805,N_23956,N_23334);
nor UO_1806 (O_1806,N_23088,N_23386);
and UO_1807 (O_1807,N_22134,N_22254);
and UO_1808 (O_1808,N_24838,N_23658);
and UO_1809 (O_1809,N_23866,N_24186);
and UO_1810 (O_1810,N_23086,N_23781);
nor UO_1811 (O_1811,N_24553,N_24509);
and UO_1812 (O_1812,N_24604,N_22197);
and UO_1813 (O_1813,N_23484,N_23180);
or UO_1814 (O_1814,N_24449,N_22335);
xor UO_1815 (O_1815,N_24404,N_24321);
or UO_1816 (O_1816,N_22209,N_23453);
and UO_1817 (O_1817,N_22186,N_24336);
and UO_1818 (O_1818,N_22126,N_22637);
or UO_1819 (O_1819,N_24285,N_24160);
and UO_1820 (O_1820,N_24376,N_22822);
and UO_1821 (O_1821,N_22086,N_22024);
nand UO_1822 (O_1822,N_23627,N_22921);
nor UO_1823 (O_1823,N_23476,N_22401);
or UO_1824 (O_1824,N_23128,N_22729);
nand UO_1825 (O_1825,N_23540,N_22217);
nand UO_1826 (O_1826,N_22649,N_22302);
or UO_1827 (O_1827,N_24225,N_24282);
or UO_1828 (O_1828,N_24759,N_24138);
or UO_1829 (O_1829,N_22941,N_23939);
or UO_1830 (O_1830,N_23396,N_23960);
nand UO_1831 (O_1831,N_24599,N_22884);
and UO_1832 (O_1832,N_22214,N_23794);
nor UO_1833 (O_1833,N_23942,N_21972);
nor UO_1834 (O_1834,N_24495,N_24976);
or UO_1835 (O_1835,N_23516,N_24453);
nor UO_1836 (O_1836,N_24711,N_23782);
xor UO_1837 (O_1837,N_22145,N_23542);
or UO_1838 (O_1838,N_23061,N_21904);
nand UO_1839 (O_1839,N_23068,N_23732);
and UO_1840 (O_1840,N_23604,N_23158);
nor UO_1841 (O_1841,N_24998,N_23129);
or UO_1842 (O_1842,N_22380,N_23138);
nor UO_1843 (O_1843,N_23283,N_23670);
nand UO_1844 (O_1844,N_23691,N_24029);
and UO_1845 (O_1845,N_22004,N_23656);
and UO_1846 (O_1846,N_24058,N_24736);
nand UO_1847 (O_1847,N_22454,N_22693);
nor UO_1848 (O_1848,N_23985,N_23830);
xor UO_1849 (O_1849,N_23391,N_24096);
nand UO_1850 (O_1850,N_23648,N_24065);
and UO_1851 (O_1851,N_22207,N_22822);
and UO_1852 (O_1852,N_23685,N_23184);
or UO_1853 (O_1853,N_23922,N_23392);
nor UO_1854 (O_1854,N_24343,N_23030);
nand UO_1855 (O_1855,N_22613,N_24646);
xor UO_1856 (O_1856,N_23063,N_22639);
nor UO_1857 (O_1857,N_22247,N_23250);
nor UO_1858 (O_1858,N_23500,N_22182);
nand UO_1859 (O_1859,N_22308,N_22726);
nand UO_1860 (O_1860,N_23739,N_22355);
nor UO_1861 (O_1861,N_23658,N_22468);
nor UO_1862 (O_1862,N_22026,N_21984);
or UO_1863 (O_1863,N_23165,N_24951);
and UO_1864 (O_1864,N_23658,N_21919);
nor UO_1865 (O_1865,N_22405,N_21941);
or UO_1866 (O_1866,N_23248,N_22354);
nor UO_1867 (O_1867,N_24464,N_23451);
and UO_1868 (O_1868,N_24588,N_24199);
nor UO_1869 (O_1869,N_22102,N_23501);
nand UO_1870 (O_1870,N_22183,N_22025);
nor UO_1871 (O_1871,N_22494,N_24813);
nand UO_1872 (O_1872,N_24474,N_21898);
nor UO_1873 (O_1873,N_22492,N_22358);
or UO_1874 (O_1874,N_21933,N_24849);
and UO_1875 (O_1875,N_21946,N_24210);
nor UO_1876 (O_1876,N_23426,N_23166);
and UO_1877 (O_1877,N_22625,N_23952);
nand UO_1878 (O_1878,N_22454,N_23821);
nor UO_1879 (O_1879,N_22875,N_22973);
xnor UO_1880 (O_1880,N_22096,N_22789);
nor UO_1881 (O_1881,N_23906,N_23001);
or UO_1882 (O_1882,N_24505,N_24750);
nand UO_1883 (O_1883,N_22316,N_23822);
nor UO_1884 (O_1884,N_22480,N_22833);
and UO_1885 (O_1885,N_22406,N_22539);
nand UO_1886 (O_1886,N_21887,N_24656);
nor UO_1887 (O_1887,N_22322,N_22095);
and UO_1888 (O_1888,N_24813,N_22177);
and UO_1889 (O_1889,N_22148,N_22903);
nand UO_1890 (O_1890,N_24486,N_24438);
or UO_1891 (O_1891,N_24870,N_23268);
or UO_1892 (O_1892,N_24497,N_21912);
and UO_1893 (O_1893,N_23849,N_22022);
nand UO_1894 (O_1894,N_22408,N_24458);
and UO_1895 (O_1895,N_23091,N_24524);
or UO_1896 (O_1896,N_23489,N_24817);
and UO_1897 (O_1897,N_21986,N_24030);
nand UO_1898 (O_1898,N_24448,N_22703);
xnor UO_1899 (O_1899,N_22473,N_23654);
nand UO_1900 (O_1900,N_22087,N_24326);
nor UO_1901 (O_1901,N_22073,N_23075);
or UO_1902 (O_1902,N_22035,N_23208);
xnor UO_1903 (O_1903,N_24442,N_22228);
or UO_1904 (O_1904,N_24697,N_22009);
nand UO_1905 (O_1905,N_21910,N_23916);
xnor UO_1906 (O_1906,N_23491,N_23723);
or UO_1907 (O_1907,N_24616,N_23913);
xor UO_1908 (O_1908,N_23190,N_24332);
nor UO_1909 (O_1909,N_22550,N_22518);
nor UO_1910 (O_1910,N_22699,N_23036);
xor UO_1911 (O_1911,N_22770,N_23559);
nor UO_1912 (O_1912,N_23205,N_22088);
nand UO_1913 (O_1913,N_23034,N_23042);
and UO_1914 (O_1914,N_24035,N_24488);
and UO_1915 (O_1915,N_23984,N_23719);
or UO_1916 (O_1916,N_22215,N_23250);
nand UO_1917 (O_1917,N_22403,N_22655);
or UO_1918 (O_1918,N_22821,N_24136);
or UO_1919 (O_1919,N_23037,N_24286);
and UO_1920 (O_1920,N_23873,N_24676);
or UO_1921 (O_1921,N_23584,N_22184);
nand UO_1922 (O_1922,N_24928,N_24921);
or UO_1923 (O_1923,N_24508,N_24943);
nor UO_1924 (O_1924,N_24440,N_24965);
nor UO_1925 (O_1925,N_22225,N_23133);
nor UO_1926 (O_1926,N_23005,N_23320);
nand UO_1927 (O_1927,N_22410,N_24142);
nand UO_1928 (O_1928,N_24279,N_24448);
nor UO_1929 (O_1929,N_24948,N_24896);
or UO_1930 (O_1930,N_23003,N_22940);
nand UO_1931 (O_1931,N_22601,N_24812);
nor UO_1932 (O_1932,N_22000,N_22632);
nand UO_1933 (O_1933,N_22325,N_24575);
and UO_1934 (O_1934,N_24551,N_23004);
and UO_1935 (O_1935,N_22300,N_24599);
or UO_1936 (O_1936,N_24673,N_24202);
or UO_1937 (O_1937,N_23416,N_21974);
nor UO_1938 (O_1938,N_22097,N_24754);
nand UO_1939 (O_1939,N_24146,N_22177);
nand UO_1940 (O_1940,N_24840,N_22126);
nor UO_1941 (O_1941,N_23485,N_23691);
nand UO_1942 (O_1942,N_23284,N_24520);
and UO_1943 (O_1943,N_24103,N_24192);
or UO_1944 (O_1944,N_23258,N_23518);
and UO_1945 (O_1945,N_24248,N_23122);
nand UO_1946 (O_1946,N_23394,N_24686);
nand UO_1947 (O_1947,N_21898,N_22161);
xnor UO_1948 (O_1948,N_24033,N_23081);
nor UO_1949 (O_1949,N_22708,N_24824);
nand UO_1950 (O_1950,N_24690,N_22174);
nand UO_1951 (O_1951,N_22334,N_21997);
xor UO_1952 (O_1952,N_24320,N_21899);
nor UO_1953 (O_1953,N_24455,N_22302);
nor UO_1954 (O_1954,N_24276,N_22425);
nor UO_1955 (O_1955,N_23817,N_24469);
nor UO_1956 (O_1956,N_22833,N_24019);
nor UO_1957 (O_1957,N_24689,N_22446);
and UO_1958 (O_1958,N_22745,N_22893);
nor UO_1959 (O_1959,N_24295,N_24294);
and UO_1960 (O_1960,N_23004,N_24939);
nand UO_1961 (O_1961,N_22129,N_22459);
or UO_1962 (O_1962,N_23418,N_23780);
and UO_1963 (O_1963,N_23532,N_22185);
or UO_1964 (O_1964,N_22782,N_23252);
nor UO_1965 (O_1965,N_24937,N_24435);
or UO_1966 (O_1966,N_22377,N_24809);
and UO_1967 (O_1967,N_24938,N_24374);
nor UO_1968 (O_1968,N_24227,N_22682);
or UO_1969 (O_1969,N_22403,N_24580);
or UO_1970 (O_1970,N_22000,N_24630);
nand UO_1971 (O_1971,N_22052,N_24624);
nand UO_1972 (O_1972,N_24725,N_24497);
nor UO_1973 (O_1973,N_24490,N_23556);
or UO_1974 (O_1974,N_24236,N_23800);
or UO_1975 (O_1975,N_23823,N_23503);
and UO_1976 (O_1976,N_22308,N_23240);
xnor UO_1977 (O_1977,N_23914,N_21968);
nand UO_1978 (O_1978,N_24156,N_24532);
nand UO_1979 (O_1979,N_22346,N_22791);
nand UO_1980 (O_1980,N_23164,N_24082);
and UO_1981 (O_1981,N_22590,N_23417);
or UO_1982 (O_1982,N_24413,N_23961);
nand UO_1983 (O_1983,N_24634,N_23273);
and UO_1984 (O_1984,N_24613,N_22131);
and UO_1985 (O_1985,N_24037,N_24177);
nor UO_1986 (O_1986,N_21897,N_24816);
nand UO_1987 (O_1987,N_23098,N_24688);
nor UO_1988 (O_1988,N_24514,N_22887);
and UO_1989 (O_1989,N_22158,N_24512);
or UO_1990 (O_1990,N_23976,N_23303);
or UO_1991 (O_1991,N_23033,N_21989);
or UO_1992 (O_1992,N_24102,N_22067);
and UO_1993 (O_1993,N_23289,N_23198);
nand UO_1994 (O_1994,N_22637,N_24689);
or UO_1995 (O_1995,N_22564,N_22372);
nand UO_1996 (O_1996,N_24152,N_22335);
and UO_1997 (O_1997,N_22645,N_22398);
or UO_1998 (O_1998,N_23469,N_24174);
xnor UO_1999 (O_1999,N_24248,N_23929);
or UO_2000 (O_2000,N_22899,N_23947);
and UO_2001 (O_2001,N_23035,N_22665);
or UO_2002 (O_2002,N_22744,N_23700);
nand UO_2003 (O_2003,N_22199,N_23051);
or UO_2004 (O_2004,N_23026,N_24952);
xnor UO_2005 (O_2005,N_23164,N_22392);
nand UO_2006 (O_2006,N_23420,N_23561);
or UO_2007 (O_2007,N_21915,N_24217);
or UO_2008 (O_2008,N_24475,N_23752);
nor UO_2009 (O_2009,N_23306,N_24645);
nor UO_2010 (O_2010,N_24999,N_22597);
and UO_2011 (O_2011,N_22920,N_24467);
nand UO_2012 (O_2012,N_22011,N_22020);
or UO_2013 (O_2013,N_21953,N_23209);
nor UO_2014 (O_2014,N_23594,N_23414);
nor UO_2015 (O_2015,N_22824,N_23342);
xnor UO_2016 (O_2016,N_23277,N_22238);
nand UO_2017 (O_2017,N_24059,N_22388);
and UO_2018 (O_2018,N_22484,N_24416);
nor UO_2019 (O_2019,N_24706,N_23295);
nand UO_2020 (O_2020,N_22669,N_24318);
and UO_2021 (O_2021,N_23062,N_23706);
nor UO_2022 (O_2022,N_24567,N_23447);
or UO_2023 (O_2023,N_23816,N_23457);
nor UO_2024 (O_2024,N_24694,N_21958);
nor UO_2025 (O_2025,N_24342,N_23979);
nand UO_2026 (O_2026,N_24827,N_22842);
and UO_2027 (O_2027,N_23358,N_22585);
or UO_2028 (O_2028,N_23200,N_22508);
nand UO_2029 (O_2029,N_23819,N_24906);
nor UO_2030 (O_2030,N_23679,N_24238);
xnor UO_2031 (O_2031,N_23364,N_24946);
xor UO_2032 (O_2032,N_24658,N_24816);
nor UO_2033 (O_2033,N_23057,N_23709);
nand UO_2034 (O_2034,N_23335,N_24091);
and UO_2035 (O_2035,N_22483,N_24826);
nor UO_2036 (O_2036,N_21938,N_23316);
or UO_2037 (O_2037,N_23491,N_22124);
nor UO_2038 (O_2038,N_24975,N_24713);
or UO_2039 (O_2039,N_23583,N_23134);
and UO_2040 (O_2040,N_23910,N_22321);
nand UO_2041 (O_2041,N_21908,N_21879);
nand UO_2042 (O_2042,N_24433,N_22551);
xnor UO_2043 (O_2043,N_22996,N_23899);
nor UO_2044 (O_2044,N_23414,N_22870);
and UO_2045 (O_2045,N_23244,N_23075);
nand UO_2046 (O_2046,N_24236,N_23994);
nand UO_2047 (O_2047,N_24962,N_22709);
and UO_2048 (O_2048,N_24581,N_22367);
nor UO_2049 (O_2049,N_23781,N_22338);
nand UO_2050 (O_2050,N_24902,N_23179);
nor UO_2051 (O_2051,N_22244,N_24638);
and UO_2052 (O_2052,N_23812,N_22696);
xnor UO_2053 (O_2053,N_23082,N_23821);
nor UO_2054 (O_2054,N_22807,N_23936);
or UO_2055 (O_2055,N_24502,N_21926);
xor UO_2056 (O_2056,N_23500,N_23630);
nor UO_2057 (O_2057,N_24636,N_23447);
or UO_2058 (O_2058,N_23842,N_23112);
and UO_2059 (O_2059,N_22142,N_24458);
xor UO_2060 (O_2060,N_22689,N_24765);
and UO_2061 (O_2061,N_23114,N_24976);
nor UO_2062 (O_2062,N_23524,N_22241);
or UO_2063 (O_2063,N_22903,N_24609);
and UO_2064 (O_2064,N_24844,N_23259);
or UO_2065 (O_2065,N_24859,N_23185);
and UO_2066 (O_2066,N_23150,N_21893);
nor UO_2067 (O_2067,N_24411,N_24077);
or UO_2068 (O_2068,N_24332,N_23641);
or UO_2069 (O_2069,N_22699,N_23448);
or UO_2070 (O_2070,N_23297,N_24005);
nor UO_2071 (O_2071,N_21999,N_22314);
and UO_2072 (O_2072,N_23006,N_22461);
xor UO_2073 (O_2073,N_24563,N_24510);
nand UO_2074 (O_2074,N_23816,N_24160);
nor UO_2075 (O_2075,N_24274,N_21898);
or UO_2076 (O_2076,N_24741,N_23469);
nor UO_2077 (O_2077,N_23895,N_23713);
or UO_2078 (O_2078,N_23465,N_24868);
xnor UO_2079 (O_2079,N_21959,N_22384);
and UO_2080 (O_2080,N_22942,N_22638);
nand UO_2081 (O_2081,N_24713,N_23419);
nor UO_2082 (O_2082,N_24391,N_22479);
and UO_2083 (O_2083,N_22729,N_22291);
and UO_2084 (O_2084,N_24001,N_23018);
and UO_2085 (O_2085,N_21989,N_23439);
or UO_2086 (O_2086,N_23324,N_23062);
nor UO_2087 (O_2087,N_22013,N_23351);
or UO_2088 (O_2088,N_23323,N_23245);
nand UO_2089 (O_2089,N_24319,N_23288);
nor UO_2090 (O_2090,N_21975,N_24412);
nand UO_2091 (O_2091,N_24233,N_23409);
nor UO_2092 (O_2092,N_23171,N_24962);
nand UO_2093 (O_2093,N_22014,N_24057);
nor UO_2094 (O_2094,N_24702,N_23909);
and UO_2095 (O_2095,N_21884,N_22740);
nor UO_2096 (O_2096,N_24537,N_22214);
and UO_2097 (O_2097,N_22568,N_24704);
nand UO_2098 (O_2098,N_22689,N_24564);
and UO_2099 (O_2099,N_22077,N_24576);
nand UO_2100 (O_2100,N_23982,N_23525);
and UO_2101 (O_2101,N_23893,N_22607);
and UO_2102 (O_2102,N_24262,N_22542);
and UO_2103 (O_2103,N_22264,N_22197);
or UO_2104 (O_2104,N_23114,N_22034);
or UO_2105 (O_2105,N_24956,N_22167);
nor UO_2106 (O_2106,N_24249,N_23989);
nand UO_2107 (O_2107,N_24580,N_22520);
nand UO_2108 (O_2108,N_23766,N_23294);
or UO_2109 (O_2109,N_23229,N_24140);
nor UO_2110 (O_2110,N_22578,N_23732);
xor UO_2111 (O_2111,N_24881,N_23722);
or UO_2112 (O_2112,N_24436,N_24375);
xnor UO_2113 (O_2113,N_24643,N_22155);
or UO_2114 (O_2114,N_22886,N_22310);
nor UO_2115 (O_2115,N_22548,N_24046);
or UO_2116 (O_2116,N_24619,N_23076);
nand UO_2117 (O_2117,N_24879,N_24151);
or UO_2118 (O_2118,N_24125,N_23622);
nand UO_2119 (O_2119,N_24339,N_24763);
nor UO_2120 (O_2120,N_22939,N_23031);
or UO_2121 (O_2121,N_22074,N_24479);
xnor UO_2122 (O_2122,N_24871,N_24635);
or UO_2123 (O_2123,N_24954,N_22515);
nand UO_2124 (O_2124,N_22921,N_24925);
or UO_2125 (O_2125,N_23892,N_22847);
nand UO_2126 (O_2126,N_22057,N_22790);
nor UO_2127 (O_2127,N_24797,N_23857);
nor UO_2128 (O_2128,N_22191,N_23714);
and UO_2129 (O_2129,N_24410,N_22797);
and UO_2130 (O_2130,N_23589,N_22382);
nor UO_2131 (O_2131,N_24429,N_24403);
nor UO_2132 (O_2132,N_22989,N_22658);
nor UO_2133 (O_2133,N_24837,N_22307);
nor UO_2134 (O_2134,N_23955,N_23165);
nor UO_2135 (O_2135,N_23244,N_23677);
or UO_2136 (O_2136,N_23985,N_23982);
nor UO_2137 (O_2137,N_23050,N_23943);
and UO_2138 (O_2138,N_23594,N_22283);
nor UO_2139 (O_2139,N_23955,N_24126);
nor UO_2140 (O_2140,N_24605,N_21935);
and UO_2141 (O_2141,N_23932,N_24655);
xnor UO_2142 (O_2142,N_24302,N_22696);
and UO_2143 (O_2143,N_22228,N_24214);
nand UO_2144 (O_2144,N_24843,N_22203);
nand UO_2145 (O_2145,N_22330,N_23648);
nor UO_2146 (O_2146,N_23525,N_23908);
or UO_2147 (O_2147,N_24827,N_21994);
or UO_2148 (O_2148,N_24193,N_22113);
nand UO_2149 (O_2149,N_24400,N_23763);
nor UO_2150 (O_2150,N_22699,N_24868);
nor UO_2151 (O_2151,N_24591,N_22396);
or UO_2152 (O_2152,N_22135,N_24082);
nand UO_2153 (O_2153,N_22429,N_24476);
xor UO_2154 (O_2154,N_22531,N_23735);
nor UO_2155 (O_2155,N_22635,N_22016);
nor UO_2156 (O_2156,N_22850,N_23767);
xor UO_2157 (O_2157,N_24150,N_23953);
or UO_2158 (O_2158,N_22490,N_22290);
nor UO_2159 (O_2159,N_22446,N_22154);
nor UO_2160 (O_2160,N_21959,N_22626);
and UO_2161 (O_2161,N_23439,N_22024);
and UO_2162 (O_2162,N_24988,N_23133);
and UO_2163 (O_2163,N_23505,N_24613);
and UO_2164 (O_2164,N_22829,N_22679);
and UO_2165 (O_2165,N_22164,N_22127);
and UO_2166 (O_2166,N_23238,N_22805);
nor UO_2167 (O_2167,N_23158,N_22982);
nor UO_2168 (O_2168,N_22222,N_23576);
and UO_2169 (O_2169,N_22714,N_24746);
or UO_2170 (O_2170,N_22427,N_23865);
xnor UO_2171 (O_2171,N_24043,N_24553);
and UO_2172 (O_2172,N_22948,N_24421);
nand UO_2173 (O_2173,N_23456,N_23078);
nand UO_2174 (O_2174,N_23204,N_23897);
nor UO_2175 (O_2175,N_23013,N_24078);
or UO_2176 (O_2176,N_23569,N_22021);
and UO_2177 (O_2177,N_22436,N_22721);
nor UO_2178 (O_2178,N_22003,N_22008);
or UO_2179 (O_2179,N_22039,N_23075);
and UO_2180 (O_2180,N_23536,N_22567);
nor UO_2181 (O_2181,N_24085,N_24999);
or UO_2182 (O_2182,N_23058,N_23502);
xor UO_2183 (O_2183,N_22317,N_23241);
nor UO_2184 (O_2184,N_22848,N_22932);
and UO_2185 (O_2185,N_24425,N_22162);
nor UO_2186 (O_2186,N_22174,N_24079);
and UO_2187 (O_2187,N_22627,N_23682);
xor UO_2188 (O_2188,N_23328,N_22252);
and UO_2189 (O_2189,N_22450,N_23118);
or UO_2190 (O_2190,N_24785,N_22778);
nor UO_2191 (O_2191,N_24886,N_22396);
and UO_2192 (O_2192,N_24077,N_23521);
nor UO_2193 (O_2193,N_24190,N_22867);
or UO_2194 (O_2194,N_22249,N_24120);
nor UO_2195 (O_2195,N_24505,N_24522);
xor UO_2196 (O_2196,N_24868,N_22450);
or UO_2197 (O_2197,N_22611,N_22357);
xnor UO_2198 (O_2198,N_22078,N_22277);
and UO_2199 (O_2199,N_23671,N_23180);
and UO_2200 (O_2200,N_22091,N_22175);
and UO_2201 (O_2201,N_24546,N_21986);
nand UO_2202 (O_2202,N_24037,N_23909);
nor UO_2203 (O_2203,N_22967,N_23276);
nor UO_2204 (O_2204,N_22967,N_23487);
nor UO_2205 (O_2205,N_23439,N_24204);
and UO_2206 (O_2206,N_23570,N_24859);
nand UO_2207 (O_2207,N_22852,N_22974);
nor UO_2208 (O_2208,N_22069,N_23745);
or UO_2209 (O_2209,N_24315,N_22648);
xor UO_2210 (O_2210,N_22096,N_22873);
nor UO_2211 (O_2211,N_23477,N_21956);
and UO_2212 (O_2212,N_23940,N_24260);
nand UO_2213 (O_2213,N_22946,N_22731);
nor UO_2214 (O_2214,N_22979,N_22718);
nor UO_2215 (O_2215,N_23797,N_24938);
or UO_2216 (O_2216,N_23553,N_23101);
or UO_2217 (O_2217,N_23977,N_24320);
and UO_2218 (O_2218,N_24410,N_22187);
nor UO_2219 (O_2219,N_24875,N_23246);
nand UO_2220 (O_2220,N_23004,N_24925);
or UO_2221 (O_2221,N_24457,N_22352);
nor UO_2222 (O_2222,N_22278,N_24194);
or UO_2223 (O_2223,N_24072,N_22139);
or UO_2224 (O_2224,N_22727,N_23298);
or UO_2225 (O_2225,N_24427,N_23368);
nand UO_2226 (O_2226,N_21879,N_23788);
or UO_2227 (O_2227,N_22603,N_23830);
nand UO_2228 (O_2228,N_23234,N_24432);
nor UO_2229 (O_2229,N_23536,N_23485);
xnor UO_2230 (O_2230,N_23783,N_22482);
xnor UO_2231 (O_2231,N_22856,N_22063);
or UO_2232 (O_2232,N_23787,N_23896);
and UO_2233 (O_2233,N_22491,N_23126);
or UO_2234 (O_2234,N_23479,N_24801);
or UO_2235 (O_2235,N_23778,N_23364);
and UO_2236 (O_2236,N_24337,N_23948);
xnor UO_2237 (O_2237,N_24145,N_23719);
and UO_2238 (O_2238,N_23694,N_23189);
or UO_2239 (O_2239,N_24065,N_24693);
nor UO_2240 (O_2240,N_23937,N_23611);
or UO_2241 (O_2241,N_22373,N_22293);
nand UO_2242 (O_2242,N_24839,N_24547);
or UO_2243 (O_2243,N_22769,N_23757);
nor UO_2244 (O_2244,N_24566,N_22011);
and UO_2245 (O_2245,N_23804,N_23280);
nor UO_2246 (O_2246,N_23249,N_22865);
nor UO_2247 (O_2247,N_23750,N_24898);
or UO_2248 (O_2248,N_24689,N_24678);
and UO_2249 (O_2249,N_22869,N_24325);
nor UO_2250 (O_2250,N_24698,N_24300);
or UO_2251 (O_2251,N_24036,N_23669);
nand UO_2252 (O_2252,N_23508,N_23533);
nand UO_2253 (O_2253,N_24869,N_22330);
or UO_2254 (O_2254,N_23227,N_23651);
nor UO_2255 (O_2255,N_23484,N_24023);
nand UO_2256 (O_2256,N_24916,N_23686);
nand UO_2257 (O_2257,N_22247,N_23980);
and UO_2258 (O_2258,N_23623,N_23971);
nor UO_2259 (O_2259,N_24215,N_24183);
and UO_2260 (O_2260,N_23704,N_23474);
and UO_2261 (O_2261,N_22329,N_22910);
and UO_2262 (O_2262,N_22197,N_22515);
and UO_2263 (O_2263,N_23579,N_24958);
or UO_2264 (O_2264,N_22018,N_24065);
xnor UO_2265 (O_2265,N_22882,N_21939);
and UO_2266 (O_2266,N_22113,N_24834);
nor UO_2267 (O_2267,N_24495,N_24755);
nor UO_2268 (O_2268,N_23660,N_24523);
nand UO_2269 (O_2269,N_22093,N_24777);
xnor UO_2270 (O_2270,N_21912,N_24140);
or UO_2271 (O_2271,N_22209,N_23029);
nand UO_2272 (O_2272,N_22350,N_23487);
or UO_2273 (O_2273,N_24951,N_24036);
nand UO_2274 (O_2274,N_22227,N_23382);
or UO_2275 (O_2275,N_22878,N_21890);
nand UO_2276 (O_2276,N_23471,N_22013);
nand UO_2277 (O_2277,N_22564,N_23492);
nor UO_2278 (O_2278,N_22927,N_24192);
nand UO_2279 (O_2279,N_23519,N_23164);
and UO_2280 (O_2280,N_23600,N_23628);
and UO_2281 (O_2281,N_24724,N_23272);
nand UO_2282 (O_2282,N_22888,N_24202);
nor UO_2283 (O_2283,N_22918,N_22459);
nor UO_2284 (O_2284,N_22905,N_23824);
or UO_2285 (O_2285,N_23127,N_22766);
and UO_2286 (O_2286,N_24672,N_21916);
nor UO_2287 (O_2287,N_22451,N_24472);
nand UO_2288 (O_2288,N_22556,N_22672);
xor UO_2289 (O_2289,N_23291,N_22880);
nor UO_2290 (O_2290,N_22615,N_23195);
and UO_2291 (O_2291,N_22191,N_22248);
xnor UO_2292 (O_2292,N_22802,N_22606);
and UO_2293 (O_2293,N_24914,N_24194);
nor UO_2294 (O_2294,N_24006,N_24568);
or UO_2295 (O_2295,N_23237,N_21947);
nor UO_2296 (O_2296,N_24694,N_22930);
or UO_2297 (O_2297,N_23866,N_24437);
or UO_2298 (O_2298,N_24420,N_24221);
or UO_2299 (O_2299,N_24300,N_22333);
and UO_2300 (O_2300,N_24835,N_24253);
nand UO_2301 (O_2301,N_22503,N_23848);
xnor UO_2302 (O_2302,N_24198,N_21968);
and UO_2303 (O_2303,N_22292,N_24720);
nor UO_2304 (O_2304,N_22504,N_23045);
nand UO_2305 (O_2305,N_22230,N_24466);
nand UO_2306 (O_2306,N_24559,N_24788);
nand UO_2307 (O_2307,N_22301,N_24940);
xnor UO_2308 (O_2308,N_23848,N_22160);
nand UO_2309 (O_2309,N_24788,N_23923);
or UO_2310 (O_2310,N_22462,N_23639);
and UO_2311 (O_2311,N_23912,N_23166);
xor UO_2312 (O_2312,N_24823,N_22876);
and UO_2313 (O_2313,N_24875,N_22733);
xnor UO_2314 (O_2314,N_23342,N_23831);
and UO_2315 (O_2315,N_22341,N_22430);
xor UO_2316 (O_2316,N_22681,N_23448);
or UO_2317 (O_2317,N_24057,N_22036);
xnor UO_2318 (O_2318,N_24826,N_24990);
and UO_2319 (O_2319,N_24299,N_23779);
xor UO_2320 (O_2320,N_22807,N_22128);
or UO_2321 (O_2321,N_23474,N_24466);
or UO_2322 (O_2322,N_23479,N_23852);
and UO_2323 (O_2323,N_22583,N_24421);
nor UO_2324 (O_2324,N_23745,N_23235);
and UO_2325 (O_2325,N_22506,N_24748);
nor UO_2326 (O_2326,N_23546,N_24121);
xnor UO_2327 (O_2327,N_23596,N_23307);
nand UO_2328 (O_2328,N_24596,N_24226);
or UO_2329 (O_2329,N_24348,N_24114);
nand UO_2330 (O_2330,N_23145,N_23869);
nand UO_2331 (O_2331,N_24454,N_24197);
nor UO_2332 (O_2332,N_22376,N_22398);
nor UO_2333 (O_2333,N_22146,N_24474);
and UO_2334 (O_2334,N_23948,N_24693);
nor UO_2335 (O_2335,N_24824,N_23581);
nor UO_2336 (O_2336,N_22547,N_23289);
xnor UO_2337 (O_2337,N_23946,N_24073);
nor UO_2338 (O_2338,N_22848,N_22322);
or UO_2339 (O_2339,N_22936,N_22266);
and UO_2340 (O_2340,N_23839,N_24896);
and UO_2341 (O_2341,N_22559,N_23491);
nor UO_2342 (O_2342,N_22505,N_24792);
nor UO_2343 (O_2343,N_23837,N_23196);
and UO_2344 (O_2344,N_22666,N_24779);
and UO_2345 (O_2345,N_22571,N_22304);
nand UO_2346 (O_2346,N_24895,N_24155);
and UO_2347 (O_2347,N_24243,N_24905);
or UO_2348 (O_2348,N_22795,N_22113);
or UO_2349 (O_2349,N_23756,N_22253);
or UO_2350 (O_2350,N_23487,N_24631);
nand UO_2351 (O_2351,N_24066,N_24017);
nor UO_2352 (O_2352,N_23748,N_22231);
or UO_2353 (O_2353,N_23510,N_23237);
xnor UO_2354 (O_2354,N_23468,N_22995);
nor UO_2355 (O_2355,N_22265,N_23232);
nand UO_2356 (O_2356,N_24357,N_24346);
nor UO_2357 (O_2357,N_22051,N_24784);
nor UO_2358 (O_2358,N_24209,N_23346);
and UO_2359 (O_2359,N_22619,N_24745);
nor UO_2360 (O_2360,N_22601,N_22706);
nand UO_2361 (O_2361,N_24459,N_22469);
or UO_2362 (O_2362,N_22895,N_22320);
and UO_2363 (O_2363,N_24040,N_24870);
and UO_2364 (O_2364,N_24583,N_22504);
nand UO_2365 (O_2365,N_22448,N_21998);
or UO_2366 (O_2366,N_23196,N_24912);
and UO_2367 (O_2367,N_23501,N_23419);
nand UO_2368 (O_2368,N_23313,N_22378);
nor UO_2369 (O_2369,N_22160,N_23641);
nand UO_2370 (O_2370,N_24657,N_22358);
xor UO_2371 (O_2371,N_22449,N_24056);
nor UO_2372 (O_2372,N_23818,N_22945);
and UO_2373 (O_2373,N_22965,N_22031);
nand UO_2374 (O_2374,N_23004,N_24619);
and UO_2375 (O_2375,N_24193,N_22646);
nand UO_2376 (O_2376,N_24821,N_22654);
and UO_2377 (O_2377,N_23308,N_22478);
or UO_2378 (O_2378,N_23944,N_24351);
or UO_2379 (O_2379,N_23852,N_23445);
and UO_2380 (O_2380,N_24755,N_23527);
or UO_2381 (O_2381,N_23043,N_24923);
nor UO_2382 (O_2382,N_24848,N_22095);
or UO_2383 (O_2383,N_21953,N_23753);
or UO_2384 (O_2384,N_22711,N_24400);
nand UO_2385 (O_2385,N_24160,N_22706);
or UO_2386 (O_2386,N_22521,N_22576);
or UO_2387 (O_2387,N_22830,N_24926);
and UO_2388 (O_2388,N_22366,N_24864);
and UO_2389 (O_2389,N_24259,N_23176);
nand UO_2390 (O_2390,N_22924,N_24875);
and UO_2391 (O_2391,N_24119,N_23258);
nor UO_2392 (O_2392,N_24070,N_22446);
nor UO_2393 (O_2393,N_24065,N_23610);
nor UO_2394 (O_2394,N_24991,N_23040);
nand UO_2395 (O_2395,N_22523,N_23243);
or UO_2396 (O_2396,N_24987,N_24123);
and UO_2397 (O_2397,N_23808,N_22918);
and UO_2398 (O_2398,N_23713,N_22659);
nor UO_2399 (O_2399,N_22924,N_23922);
nand UO_2400 (O_2400,N_22580,N_24210);
nor UO_2401 (O_2401,N_24955,N_24070);
and UO_2402 (O_2402,N_22904,N_22505);
or UO_2403 (O_2403,N_24283,N_24912);
or UO_2404 (O_2404,N_22457,N_22483);
nand UO_2405 (O_2405,N_22292,N_22877);
or UO_2406 (O_2406,N_23306,N_21987);
or UO_2407 (O_2407,N_22316,N_22499);
xor UO_2408 (O_2408,N_24228,N_24876);
nand UO_2409 (O_2409,N_23484,N_23556);
nand UO_2410 (O_2410,N_23701,N_24618);
nand UO_2411 (O_2411,N_24161,N_22205);
nor UO_2412 (O_2412,N_22898,N_24926);
and UO_2413 (O_2413,N_22736,N_23687);
or UO_2414 (O_2414,N_24904,N_24329);
and UO_2415 (O_2415,N_24840,N_22992);
or UO_2416 (O_2416,N_23973,N_23074);
nand UO_2417 (O_2417,N_22852,N_23024);
and UO_2418 (O_2418,N_22596,N_24191);
nor UO_2419 (O_2419,N_24011,N_22703);
and UO_2420 (O_2420,N_24370,N_24068);
and UO_2421 (O_2421,N_24888,N_21951);
nor UO_2422 (O_2422,N_24516,N_22122);
nor UO_2423 (O_2423,N_23891,N_23335);
nand UO_2424 (O_2424,N_22305,N_23419);
nand UO_2425 (O_2425,N_23786,N_22227);
xor UO_2426 (O_2426,N_23113,N_23427);
nor UO_2427 (O_2427,N_24270,N_22023);
nand UO_2428 (O_2428,N_24734,N_22800);
nor UO_2429 (O_2429,N_21890,N_23690);
or UO_2430 (O_2430,N_22791,N_22366);
nand UO_2431 (O_2431,N_24350,N_24987);
nand UO_2432 (O_2432,N_23405,N_22495);
nor UO_2433 (O_2433,N_22115,N_22876);
nor UO_2434 (O_2434,N_22630,N_22048);
or UO_2435 (O_2435,N_24896,N_23334);
nor UO_2436 (O_2436,N_22691,N_24025);
xor UO_2437 (O_2437,N_22613,N_23123);
nand UO_2438 (O_2438,N_23557,N_23534);
nor UO_2439 (O_2439,N_23143,N_22973);
nand UO_2440 (O_2440,N_22328,N_24794);
nand UO_2441 (O_2441,N_22653,N_21987);
or UO_2442 (O_2442,N_23461,N_23189);
nor UO_2443 (O_2443,N_23193,N_24403);
and UO_2444 (O_2444,N_22815,N_22695);
or UO_2445 (O_2445,N_24294,N_23365);
nor UO_2446 (O_2446,N_24320,N_24486);
or UO_2447 (O_2447,N_24317,N_23557);
nor UO_2448 (O_2448,N_22868,N_23612);
nand UO_2449 (O_2449,N_22629,N_22582);
or UO_2450 (O_2450,N_24424,N_23918);
or UO_2451 (O_2451,N_24458,N_22277);
or UO_2452 (O_2452,N_22773,N_22834);
nor UO_2453 (O_2453,N_22708,N_23042);
nor UO_2454 (O_2454,N_24959,N_23653);
or UO_2455 (O_2455,N_22788,N_22785);
and UO_2456 (O_2456,N_23742,N_23027);
nor UO_2457 (O_2457,N_24753,N_22804);
or UO_2458 (O_2458,N_23837,N_24173);
or UO_2459 (O_2459,N_23472,N_24149);
nor UO_2460 (O_2460,N_22769,N_22626);
nand UO_2461 (O_2461,N_24603,N_21956);
or UO_2462 (O_2462,N_24178,N_23775);
nand UO_2463 (O_2463,N_24545,N_23207);
and UO_2464 (O_2464,N_22953,N_22528);
or UO_2465 (O_2465,N_23025,N_22863);
and UO_2466 (O_2466,N_23131,N_23501);
and UO_2467 (O_2467,N_23770,N_23846);
nor UO_2468 (O_2468,N_22822,N_22017);
and UO_2469 (O_2469,N_22638,N_23627);
xnor UO_2470 (O_2470,N_24427,N_24192);
and UO_2471 (O_2471,N_24402,N_21879);
or UO_2472 (O_2472,N_23240,N_24301);
nor UO_2473 (O_2473,N_22071,N_23668);
and UO_2474 (O_2474,N_23377,N_23917);
or UO_2475 (O_2475,N_24625,N_24136);
nor UO_2476 (O_2476,N_24579,N_23374);
nand UO_2477 (O_2477,N_22218,N_24541);
nand UO_2478 (O_2478,N_24402,N_24733);
nand UO_2479 (O_2479,N_22108,N_23755);
or UO_2480 (O_2480,N_22508,N_24041);
xnor UO_2481 (O_2481,N_23156,N_24241);
and UO_2482 (O_2482,N_23012,N_23798);
nand UO_2483 (O_2483,N_22652,N_22257);
nor UO_2484 (O_2484,N_23695,N_23092);
nor UO_2485 (O_2485,N_22577,N_24301);
xnor UO_2486 (O_2486,N_24105,N_23613);
nor UO_2487 (O_2487,N_23441,N_23836);
nor UO_2488 (O_2488,N_22116,N_23860);
nand UO_2489 (O_2489,N_23923,N_22683);
nand UO_2490 (O_2490,N_24094,N_22451);
and UO_2491 (O_2491,N_22103,N_22618);
xor UO_2492 (O_2492,N_22607,N_22251);
nor UO_2493 (O_2493,N_22653,N_24217);
or UO_2494 (O_2494,N_21957,N_22609);
nand UO_2495 (O_2495,N_23822,N_22374);
nor UO_2496 (O_2496,N_24333,N_23183);
nand UO_2497 (O_2497,N_23257,N_22728);
xnor UO_2498 (O_2498,N_23792,N_24156);
nand UO_2499 (O_2499,N_23966,N_22730);
and UO_2500 (O_2500,N_24737,N_23759);
and UO_2501 (O_2501,N_23272,N_23859);
or UO_2502 (O_2502,N_24142,N_23723);
and UO_2503 (O_2503,N_23598,N_22783);
xor UO_2504 (O_2504,N_24899,N_23130);
or UO_2505 (O_2505,N_22140,N_23493);
or UO_2506 (O_2506,N_23606,N_24854);
and UO_2507 (O_2507,N_24101,N_24541);
nand UO_2508 (O_2508,N_24924,N_23834);
and UO_2509 (O_2509,N_23639,N_24724);
xor UO_2510 (O_2510,N_23941,N_24305);
and UO_2511 (O_2511,N_24694,N_24227);
nand UO_2512 (O_2512,N_23982,N_22023);
nand UO_2513 (O_2513,N_22183,N_23016);
nand UO_2514 (O_2514,N_23784,N_22169);
or UO_2515 (O_2515,N_23916,N_24141);
and UO_2516 (O_2516,N_22616,N_24274);
or UO_2517 (O_2517,N_22377,N_24547);
or UO_2518 (O_2518,N_24176,N_24593);
and UO_2519 (O_2519,N_22945,N_23598);
and UO_2520 (O_2520,N_24570,N_22894);
and UO_2521 (O_2521,N_24436,N_24708);
nor UO_2522 (O_2522,N_24842,N_23965);
and UO_2523 (O_2523,N_22513,N_22729);
and UO_2524 (O_2524,N_23582,N_24413);
nand UO_2525 (O_2525,N_24899,N_23626);
nand UO_2526 (O_2526,N_24886,N_23259);
and UO_2527 (O_2527,N_23294,N_23322);
or UO_2528 (O_2528,N_23978,N_22132);
or UO_2529 (O_2529,N_23871,N_23982);
or UO_2530 (O_2530,N_24234,N_23553);
nand UO_2531 (O_2531,N_23305,N_23582);
nand UO_2532 (O_2532,N_22304,N_23837);
or UO_2533 (O_2533,N_24166,N_23672);
nor UO_2534 (O_2534,N_22692,N_23162);
nor UO_2535 (O_2535,N_23854,N_22153);
or UO_2536 (O_2536,N_23805,N_22699);
nand UO_2537 (O_2537,N_22918,N_22272);
and UO_2538 (O_2538,N_24306,N_23296);
and UO_2539 (O_2539,N_23292,N_24861);
or UO_2540 (O_2540,N_23122,N_22127);
or UO_2541 (O_2541,N_23551,N_24033);
and UO_2542 (O_2542,N_23978,N_22383);
nor UO_2543 (O_2543,N_21900,N_24361);
nor UO_2544 (O_2544,N_23832,N_22973);
nand UO_2545 (O_2545,N_24447,N_22102);
nand UO_2546 (O_2546,N_22749,N_24094);
or UO_2547 (O_2547,N_23316,N_23134);
nor UO_2548 (O_2548,N_23961,N_24324);
nand UO_2549 (O_2549,N_24319,N_22817);
and UO_2550 (O_2550,N_24163,N_24196);
or UO_2551 (O_2551,N_24262,N_23637);
and UO_2552 (O_2552,N_24347,N_22701);
nor UO_2553 (O_2553,N_23867,N_24052);
nand UO_2554 (O_2554,N_23318,N_22980);
and UO_2555 (O_2555,N_21974,N_23490);
or UO_2556 (O_2556,N_22748,N_22835);
nand UO_2557 (O_2557,N_22294,N_23351);
xnor UO_2558 (O_2558,N_22957,N_23605);
nand UO_2559 (O_2559,N_23657,N_24285);
and UO_2560 (O_2560,N_23470,N_21937);
nand UO_2561 (O_2561,N_23713,N_23061);
and UO_2562 (O_2562,N_23398,N_22815);
and UO_2563 (O_2563,N_23341,N_22910);
and UO_2564 (O_2564,N_22819,N_22681);
nand UO_2565 (O_2565,N_23906,N_23909);
xor UO_2566 (O_2566,N_24132,N_22540);
xor UO_2567 (O_2567,N_23955,N_23566);
xor UO_2568 (O_2568,N_21996,N_22760);
nor UO_2569 (O_2569,N_22304,N_23101);
xor UO_2570 (O_2570,N_23737,N_22159);
nor UO_2571 (O_2571,N_23099,N_23146);
nor UO_2572 (O_2572,N_22565,N_23511);
or UO_2573 (O_2573,N_24568,N_22372);
and UO_2574 (O_2574,N_23600,N_23710);
and UO_2575 (O_2575,N_22968,N_24237);
nor UO_2576 (O_2576,N_24897,N_24450);
nor UO_2577 (O_2577,N_23287,N_22992);
nand UO_2578 (O_2578,N_22092,N_23138);
or UO_2579 (O_2579,N_22703,N_22961);
nor UO_2580 (O_2580,N_24719,N_22118);
and UO_2581 (O_2581,N_24691,N_24872);
and UO_2582 (O_2582,N_24952,N_23293);
and UO_2583 (O_2583,N_23430,N_22264);
nor UO_2584 (O_2584,N_24003,N_24186);
or UO_2585 (O_2585,N_24852,N_22188);
and UO_2586 (O_2586,N_23372,N_24361);
nand UO_2587 (O_2587,N_23165,N_24943);
or UO_2588 (O_2588,N_24430,N_22621);
xor UO_2589 (O_2589,N_22710,N_23913);
or UO_2590 (O_2590,N_24419,N_23967);
nor UO_2591 (O_2591,N_22026,N_23766);
nand UO_2592 (O_2592,N_24064,N_24161);
or UO_2593 (O_2593,N_24132,N_23504);
and UO_2594 (O_2594,N_24898,N_24115);
xnor UO_2595 (O_2595,N_24715,N_24376);
nor UO_2596 (O_2596,N_23649,N_23760);
and UO_2597 (O_2597,N_23866,N_22167);
and UO_2598 (O_2598,N_23162,N_24963);
nor UO_2599 (O_2599,N_24913,N_22711);
nand UO_2600 (O_2600,N_22950,N_24477);
nor UO_2601 (O_2601,N_24685,N_22268);
and UO_2602 (O_2602,N_22267,N_22784);
nand UO_2603 (O_2603,N_24444,N_22777);
or UO_2604 (O_2604,N_24867,N_22807);
nand UO_2605 (O_2605,N_22086,N_24317);
nor UO_2606 (O_2606,N_24964,N_23841);
xnor UO_2607 (O_2607,N_22337,N_22453);
or UO_2608 (O_2608,N_22793,N_23673);
nand UO_2609 (O_2609,N_23324,N_22036);
nand UO_2610 (O_2610,N_24165,N_23867);
nand UO_2611 (O_2611,N_23164,N_22311);
nor UO_2612 (O_2612,N_23822,N_22771);
or UO_2613 (O_2613,N_24607,N_24523);
nor UO_2614 (O_2614,N_22069,N_23603);
or UO_2615 (O_2615,N_24893,N_24367);
and UO_2616 (O_2616,N_24987,N_22780);
or UO_2617 (O_2617,N_23975,N_23938);
nand UO_2618 (O_2618,N_21979,N_24681);
nand UO_2619 (O_2619,N_23982,N_23487);
or UO_2620 (O_2620,N_23785,N_22874);
nor UO_2621 (O_2621,N_22372,N_23738);
and UO_2622 (O_2622,N_24826,N_22009);
and UO_2623 (O_2623,N_22209,N_23776);
or UO_2624 (O_2624,N_22050,N_24169);
and UO_2625 (O_2625,N_21959,N_23821);
xor UO_2626 (O_2626,N_22449,N_22483);
or UO_2627 (O_2627,N_23561,N_22382);
xnor UO_2628 (O_2628,N_22716,N_24028);
or UO_2629 (O_2629,N_22966,N_22312);
nand UO_2630 (O_2630,N_23903,N_22918);
nor UO_2631 (O_2631,N_23957,N_22299);
or UO_2632 (O_2632,N_24459,N_22439);
nor UO_2633 (O_2633,N_23203,N_24397);
nand UO_2634 (O_2634,N_24616,N_22823);
and UO_2635 (O_2635,N_23462,N_22309);
nand UO_2636 (O_2636,N_22048,N_23609);
and UO_2637 (O_2637,N_22444,N_23780);
nor UO_2638 (O_2638,N_24742,N_23052);
nor UO_2639 (O_2639,N_22805,N_24930);
nand UO_2640 (O_2640,N_22942,N_22749);
nand UO_2641 (O_2641,N_22556,N_22513);
nor UO_2642 (O_2642,N_24762,N_22498);
and UO_2643 (O_2643,N_22791,N_23670);
and UO_2644 (O_2644,N_22646,N_22319);
and UO_2645 (O_2645,N_23216,N_22172);
or UO_2646 (O_2646,N_22205,N_22383);
nand UO_2647 (O_2647,N_23944,N_23453);
nand UO_2648 (O_2648,N_24159,N_24291);
nand UO_2649 (O_2649,N_23458,N_24624);
or UO_2650 (O_2650,N_24922,N_23407);
and UO_2651 (O_2651,N_23393,N_23785);
and UO_2652 (O_2652,N_22733,N_22452);
nor UO_2653 (O_2653,N_24506,N_24364);
or UO_2654 (O_2654,N_23673,N_22385);
nand UO_2655 (O_2655,N_24570,N_22491);
or UO_2656 (O_2656,N_22843,N_23284);
nand UO_2657 (O_2657,N_22625,N_21905);
or UO_2658 (O_2658,N_23959,N_22322);
nand UO_2659 (O_2659,N_22555,N_24282);
nor UO_2660 (O_2660,N_23139,N_22945);
nor UO_2661 (O_2661,N_22922,N_24185);
and UO_2662 (O_2662,N_21882,N_24527);
nor UO_2663 (O_2663,N_23970,N_24680);
or UO_2664 (O_2664,N_24612,N_23033);
or UO_2665 (O_2665,N_22743,N_23211);
and UO_2666 (O_2666,N_22568,N_23447);
and UO_2667 (O_2667,N_24135,N_21900);
or UO_2668 (O_2668,N_24095,N_22592);
nor UO_2669 (O_2669,N_24299,N_22310);
or UO_2670 (O_2670,N_22517,N_23256);
nor UO_2671 (O_2671,N_22647,N_24571);
and UO_2672 (O_2672,N_22308,N_24149);
xnor UO_2673 (O_2673,N_24272,N_23933);
nor UO_2674 (O_2674,N_24500,N_23630);
xnor UO_2675 (O_2675,N_22060,N_22444);
and UO_2676 (O_2676,N_22305,N_24418);
nand UO_2677 (O_2677,N_23870,N_22722);
nor UO_2678 (O_2678,N_24106,N_24639);
nand UO_2679 (O_2679,N_22065,N_24941);
or UO_2680 (O_2680,N_22153,N_23181);
nand UO_2681 (O_2681,N_24044,N_23903);
nor UO_2682 (O_2682,N_24883,N_23448);
and UO_2683 (O_2683,N_22098,N_22831);
nand UO_2684 (O_2684,N_23544,N_23759);
nand UO_2685 (O_2685,N_23335,N_24517);
and UO_2686 (O_2686,N_23568,N_23266);
or UO_2687 (O_2687,N_22288,N_22202);
nor UO_2688 (O_2688,N_21892,N_22132);
nor UO_2689 (O_2689,N_22755,N_21906);
nand UO_2690 (O_2690,N_22232,N_24219);
xor UO_2691 (O_2691,N_24839,N_23407);
nand UO_2692 (O_2692,N_22867,N_23413);
or UO_2693 (O_2693,N_23075,N_23909);
and UO_2694 (O_2694,N_24724,N_22905);
or UO_2695 (O_2695,N_23631,N_22077);
or UO_2696 (O_2696,N_23111,N_24002);
and UO_2697 (O_2697,N_23806,N_24654);
nand UO_2698 (O_2698,N_23321,N_23678);
nor UO_2699 (O_2699,N_24449,N_24943);
nor UO_2700 (O_2700,N_23950,N_24901);
nand UO_2701 (O_2701,N_23804,N_24534);
or UO_2702 (O_2702,N_23999,N_24373);
and UO_2703 (O_2703,N_23533,N_22224);
xor UO_2704 (O_2704,N_23598,N_24533);
xor UO_2705 (O_2705,N_24673,N_23050);
nor UO_2706 (O_2706,N_23841,N_22451);
nor UO_2707 (O_2707,N_23179,N_22142);
and UO_2708 (O_2708,N_21983,N_24826);
xnor UO_2709 (O_2709,N_24907,N_24697);
nand UO_2710 (O_2710,N_23880,N_22482);
nor UO_2711 (O_2711,N_22205,N_22815);
xor UO_2712 (O_2712,N_22489,N_21944);
and UO_2713 (O_2713,N_23426,N_21883);
and UO_2714 (O_2714,N_24067,N_23948);
and UO_2715 (O_2715,N_24911,N_22423);
nor UO_2716 (O_2716,N_23996,N_24544);
and UO_2717 (O_2717,N_24579,N_22957);
nand UO_2718 (O_2718,N_23838,N_22609);
xor UO_2719 (O_2719,N_22206,N_22992);
or UO_2720 (O_2720,N_22312,N_22886);
or UO_2721 (O_2721,N_24703,N_23964);
nor UO_2722 (O_2722,N_23801,N_23934);
or UO_2723 (O_2723,N_23759,N_24819);
nand UO_2724 (O_2724,N_22219,N_24390);
or UO_2725 (O_2725,N_22240,N_22400);
xnor UO_2726 (O_2726,N_23739,N_23762);
or UO_2727 (O_2727,N_22076,N_24038);
or UO_2728 (O_2728,N_23113,N_23173);
nor UO_2729 (O_2729,N_24321,N_23799);
nor UO_2730 (O_2730,N_22628,N_24811);
or UO_2731 (O_2731,N_23124,N_23205);
and UO_2732 (O_2732,N_23291,N_23949);
xnor UO_2733 (O_2733,N_23936,N_23811);
xnor UO_2734 (O_2734,N_23907,N_23733);
or UO_2735 (O_2735,N_22921,N_23469);
and UO_2736 (O_2736,N_23151,N_24027);
nand UO_2737 (O_2737,N_22068,N_23994);
xor UO_2738 (O_2738,N_23638,N_23931);
and UO_2739 (O_2739,N_24486,N_22747);
xor UO_2740 (O_2740,N_22996,N_24041);
and UO_2741 (O_2741,N_22204,N_21992);
nand UO_2742 (O_2742,N_22238,N_24205);
xor UO_2743 (O_2743,N_24133,N_21929);
nand UO_2744 (O_2744,N_23986,N_24539);
or UO_2745 (O_2745,N_23248,N_24575);
nor UO_2746 (O_2746,N_22653,N_23417);
nor UO_2747 (O_2747,N_23973,N_22952);
and UO_2748 (O_2748,N_23756,N_23887);
and UO_2749 (O_2749,N_23737,N_23089);
and UO_2750 (O_2750,N_23022,N_23786);
nor UO_2751 (O_2751,N_23205,N_23547);
and UO_2752 (O_2752,N_24493,N_23865);
nand UO_2753 (O_2753,N_24356,N_24522);
and UO_2754 (O_2754,N_22550,N_22924);
nor UO_2755 (O_2755,N_22787,N_22879);
nor UO_2756 (O_2756,N_22603,N_23362);
nand UO_2757 (O_2757,N_24937,N_23643);
and UO_2758 (O_2758,N_24684,N_22639);
nand UO_2759 (O_2759,N_23029,N_22027);
or UO_2760 (O_2760,N_22745,N_22033);
nand UO_2761 (O_2761,N_24656,N_22059);
nand UO_2762 (O_2762,N_24413,N_22130);
nand UO_2763 (O_2763,N_24649,N_23563);
and UO_2764 (O_2764,N_22295,N_23316);
nand UO_2765 (O_2765,N_23279,N_23127);
xnor UO_2766 (O_2766,N_22254,N_22417);
or UO_2767 (O_2767,N_22764,N_22288);
and UO_2768 (O_2768,N_22491,N_22501);
or UO_2769 (O_2769,N_23875,N_24721);
nand UO_2770 (O_2770,N_23602,N_24819);
or UO_2771 (O_2771,N_23425,N_24457);
or UO_2772 (O_2772,N_23226,N_24529);
nand UO_2773 (O_2773,N_23054,N_24003);
or UO_2774 (O_2774,N_23137,N_23955);
nor UO_2775 (O_2775,N_24858,N_23237);
nor UO_2776 (O_2776,N_22024,N_23386);
or UO_2777 (O_2777,N_23284,N_22840);
or UO_2778 (O_2778,N_22930,N_24785);
or UO_2779 (O_2779,N_23960,N_23358);
and UO_2780 (O_2780,N_22710,N_22973);
and UO_2781 (O_2781,N_24859,N_23840);
and UO_2782 (O_2782,N_23291,N_23057);
or UO_2783 (O_2783,N_24002,N_23441);
nor UO_2784 (O_2784,N_24401,N_24379);
nor UO_2785 (O_2785,N_24951,N_23539);
or UO_2786 (O_2786,N_24035,N_24981);
or UO_2787 (O_2787,N_22120,N_23765);
and UO_2788 (O_2788,N_23638,N_22746);
nand UO_2789 (O_2789,N_23810,N_23723);
nor UO_2790 (O_2790,N_23908,N_22909);
and UO_2791 (O_2791,N_24137,N_24390);
nor UO_2792 (O_2792,N_24565,N_24458);
nor UO_2793 (O_2793,N_24948,N_23064);
nor UO_2794 (O_2794,N_23521,N_22947);
nand UO_2795 (O_2795,N_23701,N_22510);
and UO_2796 (O_2796,N_23878,N_24276);
and UO_2797 (O_2797,N_23500,N_22896);
or UO_2798 (O_2798,N_23534,N_23332);
and UO_2799 (O_2799,N_23659,N_22305);
and UO_2800 (O_2800,N_22475,N_23302);
and UO_2801 (O_2801,N_22999,N_22678);
nand UO_2802 (O_2802,N_24515,N_22287);
nand UO_2803 (O_2803,N_22399,N_22200);
and UO_2804 (O_2804,N_22146,N_22073);
xnor UO_2805 (O_2805,N_24632,N_22768);
or UO_2806 (O_2806,N_24528,N_22203);
nor UO_2807 (O_2807,N_23339,N_22435);
or UO_2808 (O_2808,N_24106,N_22673);
nor UO_2809 (O_2809,N_24107,N_24265);
or UO_2810 (O_2810,N_24513,N_24921);
or UO_2811 (O_2811,N_22793,N_22552);
nor UO_2812 (O_2812,N_23304,N_23724);
nand UO_2813 (O_2813,N_24117,N_23196);
nor UO_2814 (O_2814,N_23170,N_22748);
xnor UO_2815 (O_2815,N_22986,N_22776);
nand UO_2816 (O_2816,N_22224,N_22922);
or UO_2817 (O_2817,N_23537,N_22427);
nor UO_2818 (O_2818,N_23136,N_22484);
nand UO_2819 (O_2819,N_23491,N_24164);
or UO_2820 (O_2820,N_22491,N_21906);
xor UO_2821 (O_2821,N_22331,N_23372);
xnor UO_2822 (O_2822,N_21917,N_23332);
nor UO_2823 (O_2823,N_22006,N_22772);
or UO_2824 (O_2824,N_24420,N_21883);
or UO_2825 (O_2825,N_23480,N_23245);
nor UO_2826 (O_2826,N_24163,N_23419);
xor UO_2827 (O_2827,N_23206,N_22684);
or UO_2828 (O_2828,N_24806,N_24730);
nor UO_2829 (O_2829,N_22833,N_23584);
nor UO_2830 (O_2830,N_22747,N_24066);
nand UO_2831 (O_2831,N_22115,N_21920);
xnor UO_2832 (O_2832,N_24777,N_24035);
or UO_2833 (O_2833,N_24863,N_22726);
or UO_2834 (O_2834,N_24419,N_23321);
nor UO_2835 (O_2835,N_23538,N_23853);
and UO_2836 (O_2836,N_23152,N_24594);
or UO_2837 (O_2837,N_24555,N_22013);
and UO_2838 (O_2838,N_22398,N_23611);
nand UO_2839 (O_2839,N_23239,N_24321);
nor UO_2840 (O_2840,N_24097,N_23959);
and UO_2841 (O_2841,N_22863,N_24221);
or UO_2842 (O_2842,N_22391,N_23888);
nand UO_2843 (O_2843,N_23986,N_23327);
or UO_2844 (O_2844,N_23448,N_22405);
nor UO_2845 (O_2845,N_24739,N_23622);
and UO_2846 (O_2846,N_21931,N_22664);
and UO_2847 (O_2847,N_24866,N_24006);
and UO_2848 (O_2848,N_23083,N_24035);
nand UO_2849 (O_2849,N_22895,N_23397);
and UO_2850 (O_2850,N_22893,N_22864);
or UO_2851 (O_2851,N_23855,N_23147);
nor UO_2852 (O_2852,N_23066,N_22808);
xnor UO_2853 (O_2853,N_23478,N_22144);
nand UO_2854 (O_2854,N_22076,N_22920);
nand UO_2855 (O_2855,N_24351,N_21990);
nand UO_2856 (O_2856,N_24521,N_23928);
and UO_2857 (O_2857,N_24409,N_24091);
and UO_2858 (O_2858,N_23207,N_24119);
or UO_2859 (O_2859,N_23490,N_24845);
nand UO_2860 (O_2860,N_24247,N_23364);
nand UO_2861 (O_2861,N_24531,N_23500);
nor UO_2862 (O_2862,N_23971,N_22036);
nand UO_2863 (O_2863,N_24183,N_24157);
nor UO_2864 (O_2864,N_22602,N_23987);
nor UO_2865 (O_2865,N_23794,N_24007);
and UO_2866 (O_2866,N_24191,N_23103);
nand UO_2867 (O_2867,N_24180,N_24205);
nor UO_2868 (O_2868,N_23108,N_24282);
xor UO_2869 (O_2869,N_22594,N_22469);
nand UO_2870 (O_2870,N_23726,N_23337);
and UO_2871 (O_2871,N_23689,N_21936);
nand UO_2872 (O_2872,N_21875,N_23007);
and UO_2873 (O_2873,N_21996,N_23778);
and UO_2874 (O_2874,N_22234,N_24084);
nand UO_2875 (O_2875,N_23759,N_23173);
or UO_2876 (O_2876,N_22630,N_22669);
xor UO_2877 (O_2877,N_24672,N_24644);
nand UO_2878 (O_2878,N_24612,N_24756);
and UO_2879 (O_2879,N_24095,N_24292);
nor UO_2880 (O_2880,N_23074,N_23166);
and UO_2881 (O_2881,N_23165,N_23589);
xnor UO_2882 (O_2882,N_21950,N_23409);
and UO_2883 (O_2883,N_24469,N_24922);
and UO_2884 (O_2884,N_24625,N_23433);
nor UO_2885 (O_2885,N_22714,N_23963);
and UO_2886 (O_2886,N_23855,N_22934);
or UO_2887 (O_2887,N_24512,N_24328);
and UO_2888 (O_2888,N_21901,N_22066);
or UO_2889 (O_2889,N_23465,N_24050);
and UO_2890 (O_2890,N_23383,N_22939);
nor UO_2891 (O_2891,N_23480,N_23037);
nor UO_2892 (O_2892,N_24704,N_23505);
xor UO_2893 (O_2893,N_22962,N_23569);
and UO_2894 (O_2894,N_23357,N_23095);
and UO_2895 (O_2895,N_22964,N_24365);
and UO_2896 (O_2896,N_24444,N_22617);
and UO_2897 (O_2897,N_24174,N_24995);
and UO_2898 (O_2898,N_22365,N_24305);
nor UO_2899 (O_2899,N_23710,N_24680);
nor UO_2900 (O_2900,N_23140,N_23718);
or UO_2901 (O_2901,N_21947,N_23346);
and UO_2902 (O_2902,N_23552,N_23063);
and UO_2903 (O_2903,N_24277,N_23708);
nand UO_2904 (O_2904,N_22931,N_22653);
xnor UO_2905 (O_2905,N_22176,N_24915);
or UO_2906 (O_2906,N_22357,N_23156);
xor UO_2907 (O_2907,N_24836,N_22008);
or UO_2908 (O_2908,N_24075,N_23074);
or UO_2909 (O_2909,N_22587,N_24286);
nor UO_2910 (O_2910,N_22207,N_22907);
or UO_2911 (O_2911,N_24650,N_22656);
xnor UO_2912 (O_2912,N_24086,N_22782);
or UO_2913 (O_2913,N_24308,N_24410);
and UO_2914 (O_2914,N_23782,N_23436);
nand UO_2915 (O_2915,N_24997,N_22716);
nand UO_2916 (O_2916,N_22094,N_24938);
and UO_2917 (O_2917,N_24501,N_22255);
or UO_2918 (O_2918,N_23040,N_21997);
or UO_2919 (O_2919,N_23263,N_23098);
nor UO_2920 (O_2920,N_22460,N_24181);
or UO_2921 (O_2921,N_22327,N_23942);
or UO_2922 (O_2922,N_24836,N_22373);
nor UO_2923 (O_2923,N_22403,N_24336);
nor UO_2924 (O_2924,N_23463,N_23997);
or UO_2925 (O_2925,N_23251,N_24340);
nor UO_2926 (O_2926,N_22875,N_24677);
nand UO_2927 (O_2927,N_24848,N_24859);
or UO_2928 (O_2928,N_22542,N_22471);
nand UO_2929 (O_2929,N_23490,N_23954);
or UO_2930 (O_2930,N_23136,N_23573);
nand UO_2931 (O_2931,N_24050,N_22563);
or UO_2932 (O_2932,N_22646,N_24700);
and UO_2933 (O_2933,N_24127,N_22258);
and UO_2934 (O_2934,N_24297,N_23542);
nand UO_2935 (O_2935,N_24605,N_23897);
nand UO_2936 (O_2936,N_23408,N_24831);
nand UO_2937 (O_2937,N_22247,N_24025);
and UO_2938 (O_2938,N_22842,N_24089);
and UO_2939 (O_2939,N_24051,N_24541);
xor UO_2940 (O_2940,N_22237,N_24052);
nor UO_2941 (O_2941,N_22133,N_23584);
nor UO_2942 (O_2942,N_24105,N_23307);
xor UO_2943 (O_2943,N_23551,N_23658);
and UO_2944 (O_2944,N_24572,N_24510);
and UO_2945 (O_2945,N_23621,N_21928);
nor UO_2946 (O_2946,N_22536,N_24570);
or UO_2947 (O_2947,N_22775,N_24026);
and UO_2948 (O_2948,N_23849,N_24329);
or UO_2949 (O_2949,N_22113,N_22135);
nand UO_2950 (O_2950,N_23981,N_22110);
nor UO_2951 (O_2951,N_22608,N_22370);
and UO_2952 (O_2952,N_24413,N_24393);
nand UO_2953 (O_2953,N_24389,N_23655);
nor UO_2954 (O_2954,N_22067,N_22012);
and UO_2955 (O_2955,N_23324,N_23558);
nor UO_2956 (O_2956,N_23846,N_24362);
nand UO_2957 (O_2957,N_23851,N_23763);
nor UO_2958 (O_2958,N_21934,N_24841);
and UO_2959 (O_2959,N_24148,N_23003);
or UO_2960 (O_2960,N_24824,N_23739);
or UO_2961 (O_2961,N_23780,N_22805);
nor UO_2962 (O_2962,N_24290,N_22955);
nand UO_2963 (O_2963,N_22752,N_22275);
nor UO_2964 (O_2964,N_24482,N_22208);
or UO_2965 (O_2965,N_22660,N_21979);
and UO_2966 (O_2966,N_24050,N_22795);
nor UO_2967 (O_2967,N_22629,N_22384);
nor UO_2968 (O_2968,N_24088,N_24269);
nor UO_2969 (O_2969,N_21951,N_23348);
and UO_2970 (O_2970,N_24090,N_23686);
and UO_2971 (O_2971,N_24458,N_22912);
nor UO_2972 (O_2972,N_23699,N_24256);
nor UO_2973 (O_2973,N_22924,N_23399);
nand UO_2974 (O_2974,N_22164,N_22196);
nand UO_2975 (O_2975,N_23193,N_24576);
or UO_2976 (O_2976,N_23265,N_24796);
and UO_2977 (O_2977,N_23816,N_23713);
or UO_2978 (O_2978,N_22938,N_23823);
nand UO_2979 (O_2979,N_23676,N_22654);
and UO_2980 (O_2980,N_22266,N_24970);
xnor UO_2981 (O_2981,N_24264,N_22721);
or UO_2982 (O_2982,N_23143,N_24889);
and UO_2983 (O_2983,N_22456,N_24465);
xor UO_2984 (O_2984,N_23113,N_22352);
nor UO_2985 (O_2985,N_23638,N_24440);
xnor UO_2986 (O_2986,N_23121,N_23721);
nor UO_2987 (O_2987,N_24158,N_24033);
and UO_2988 (O_2988,N_22497,N_24151);
nor UO_2989 (O_2989,N_22028,N_22087);
nor UO_2990 (O_2990,N_22856,N_22592);
nand UO_2991 (O_2991,N_24811,N_23972);
xnor UO_2992 (O_2992,N_22696,N_22672);
or UO_2993 (O_2993,N_23413,N_24085);
or UO_2994 (O_2994,N_24505,N_23065);
nor UO_2995 (O_2995,N_22659,N_23696);
nor UO_2996 (O_2996,N_23637,N_22489);
and UO_2997 (O_2997,N_22162,N_23617);
nand UO_2998 (O_2998,N_22998,N_24865);
xnor UO_2999 (O_2999,N_24478,N_24869);
endmodule