module basic_1500_15000_2000_75_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_833,In_196);
xor U1 (N_1,In_98,In_661);
or U2 (N_2,In_46,In_1148);
nor U3 (N_3,In_633,In_1200);
nor U4 (N_4,In_1096,In_1342);
or U5 (N_5,In_877,In_379);
xor U6 (N_6,In_20,In_9);
or U7 (N_7,In_329,In_368);
xnor U8 (N_8,In_253,In_51);
nor U9 (N_9,In_1431,In_532);
nor U10 (N_10,In_624,In_1032);
nor U11 (N_11,In_1105,In_652);
or U12 (N_12,In_1001,In_945);
xor U13 (N_13,In_545,In_440);
or U14 (N_14,In_421,In_798);
xnor U15 (N_15,In_521,In_836);
nand U16 (N_16,In_1341,In_268);
xor U17 (N_17,In_157,In_892);
xnor U18 (N_18,In_416,In_881);
xnor U19 (N_19,In_817,In_1386);
and U20 (N_20,In_1213,In_1223);
and U21 (N_21,In_968,In_839);
or U22 (N_22,In_535,In_457);
nand U23 (N_23,In_30,In_39);
nand U24 (N_24,In_720,In_1450);
xor U25 (N_25,In_1022,In_310);
and U26 (N_26,In_999,In_623);
and U27 (N_27,In_381,In_461);
xor U28 (N_28,In_1278,In_852);
and U29 (N_29,In_481,In_330);
nor U30 (N_30,In_216,In_608);
or U31 (N_31,In_691,In_832);
nand U32 (N_32,In_269,In_426);
xor U33 (N_33,In_1282,In_478);
nand U34 (N_34,In_1488,In_703);
nor U35 (N_35,In_1272,In_942);
and U36 (N_36,In_1146,In_889);
and U37 (N_37,In_208,In_1322);
and U38 (N_38,In_214,In_24);
and U39 (N_39,In_256,In_1081);
and U40 (N_40,In_921,In_1416);
nor U41 (N_41,In_1215,In_627);
and U42 (N_42,In_843,In_1493);
and U43 (N_43,In_826,In_636);
nand U44 (N_44,In_634,In_1058);
or U45 (N_45,In_1210,In_539);
xnor U46 (N_46,In_513,In_1007);
or U47 (N_47,In_1296,In_89);
and U48 (N_48,In_909,In_940);
and U49 (N_49,In_1233,In_86);
xnor U50 (N_50,In_763,In_1290);
or U51 (N_51,In_1027,In_610);
xor U52 (N_52,In_311,In_1017);
xnor U53 (N_53,In_533,In_371);
xnor U54 (N_54,In_463,In_1126);
or U55 (N_55,In_181,In_854);
or U56 (N_56,In_84,In_960);
xor U57 (N_57,In_584,In_1339);
nor U58 (N_58,In_66,In_471);
nand U59 (N_59,In_516,In_1161);
nor U60 (N_60,In_126,In_737);
xnor U61 (N_61,In_1425,In_849);
nor U62 (N_62,In_825,In_923);
xor U63 (N_63,In_856,In_199);
or U64 (N_64,In_434,In_122);
xnor U65 (N_65,In_615,In_354);
nand U66 (N_66,In_1359,In_308);
and U67 (N_67,In_682,In_1289);
nand U68 (N_68,In_931,In_1042);
nor U69 (N_69,In_99,In_591);
or U70 (N_70,In_15,In_668);
xnor U71 (N_71,In_76,In_569);
and U72 (N_72,In_1206,In_684);
or U73 (N_73,In_997,In_1265);
and U74 (N_74,In_231,In_517);
or U75 (N_75,In_234,In_152);
nor U76 (N_76,In_727,In_777);
or U77 (N_77,In_1098,In_1154);
nor U78 (N_78,In_315,In_272);
nand U79 (N_79,In_1152,In_638);
nor U80 (N_80,In_523,In_343);
or U81 (N_81,In_896,In_1066);
and U82 (N_82,In_1413,In_36);
and U83 (N_83,In_495,In_820);
xor U84 (N_84,In_319,In_698);
nand U85 (N_85,In_904,In_410);
nor U86 (N_86,In_17,In_985);
and U87 (N_87,In_588,In_910);
and U88 (N_88,In_1155,In_241);
and U89 (N_89,In_1417,In_660);
xnor U90 (N_90,In_1079,In_838);
and U91 (N_91,In_948,In_151);
or U92 (N_92,In_304,In_938);
xnor U93 (N_93,In_48,In_1064);
or U94 (N_94,In_642,In_286);
and U95 (N_95,In_1497,In_873);
or U96 (N_96,In_1082,In_753);
xor U97 (N_97,In_185,In_988);
nor U98 (N_98,In_639,In_1074);
xor U99 (N_99,In_518,In_32);
nand U100 (N_100,In_1407,In_472);
xnor U101 (N_101,In_246,In_1216);
and U102 (N_102,In_1016,In_1059);
nand U103 (N_103,In_251,In_82);
or U104 (N_104,In_5,In_977);
and U105 (N_105,In_612,In_946);
xnor U106 (N_106,In_43,In_1006);
or U107 (N_107,In_582,In_869);
nor U108 (N_108,In_1071,In_123);
and U109 (N_109,In_930,In_1327);
nor U110 (N_110,In_823,In_62);
nand U111 (N_111,In_748,In_1004);
and U112 (N_112,In_803,In_834);
or U113 (N_113,In_1185,In_1217);
nand U114 (N_114,In_1255,In_100);
nor U115 (N_115,In_562,In_1034);
xor U116 (N_116,In_1305,In_511);
or U117 (N_117,In_870,In_1326);
and U118 (N_118,In_656,In_769);
nand U119 (N_119,In_38,In_1434);
or U120 (N_120,In_644,In_1468);
or U121 (N_121,In_127,In_927);
nand U122 (N_122,In_73,In_863);
or U123 (N_123,In_822,In_814);
xor U124 (N_124,In_860,In_1372);
and U125 (N_125,In_1276,In_735);
xnor U126 (N_126,In_149,In_439);
and U127 (N_127,In_801,In_150);
nand U128 (N_128,In_1026,In_679);
nand U129 (N_129,In_50,In_1165);
or U130 (N_130,In_141,In_1243);
xnor U131 (N_131,In_235,In_441);
and U132 (N_132,In_1487,In_233);
and U133 (N_133,In_1367,In_1041);
nor U134 (N_134,In_204,In_1020);
or U135 (N_135,In_383,In_594);
xor U136 (N_136,In_1422,In_678);
or U137 (N_137,In_1136,In_508);
xnor U138 (N_138,In_673,In_905);
and U139 (N_139,In_767,In_766);
xor U140 (N_140,In_959,In_68);
nand U141 (N_141,In_363,In_56);
nor U142 (N_142,In_1121,In_366);
and U143 (N_143,In_578,In_292);
or U144 (N_144,In_1212,In_929);
nor U145 (N_145,In_955,In_859);
xor U146 (N_146,In_16,In_374);
or U147 (N_147,In_34,In_1410);
and U148 (N_148,In_1112,In_509);
nand U149 (N_149,In_1402,In_276);
or U150 (N_150,In_590,In_619);
and U151 (N_151,In_281,In_550);
nor U152 (N_152,In_1463,In_1315);
nand U153 (N_153,In_649,In_1308);
xor U154 (N_154,In_317,In_802);
or U155 (N_155,In_220,In_779);
or U156 (N_156,In_617,In_1228);
or U157 (N_157,In_117,In_996);
and U158 (N_158,In_1182,In_771);
xor U159 (N_159,In_773,In_1134);
and U160 (N_160,In_982,In_184);
and U161 (N_161,In_1418,In_1334);
nand U162 (N_162,In_1354,In_707);
xnor U163 (N_163,In_53,In_1335);
nor U164 (N_164,In_925,In_331);
and U165 (N_165,In_1170,In_283);
and U166 (N_166,In_688,In_1370);
xnor U167 (N_167,In_159,In_1403);
xor U168 (N_168,In_190,In_764);
nor U169 (N_169,In_1317,In_294);
and U170 (N_170,In_1333,In_260);
and U171 (N_171,In_1309,In_405);
and U172 (N_172,In_218,In_1441);
nor U173 (N_173,In_719,In_129);
xnor U174 (N_174,In_394,In_212);
xor U175 (N_175,In_29,In_1099);
nand U176 (N_176,In_774,In_525);
nand U177 (N_177,In_812,In_1275);
and U178 (N_178,In_1406,In_756);
nor U179 (N_179,In_64,In_1436);
or U180 (N_180,In_872,In_238);
and U181 (N_181,In_1464,In_1150);
and U182 (N_182,In_307,In_237);
and U183 (N_183,In_1439,In_55);
and U184 (N_184,In_314,In_1107);
xnor U185 (N_185,In_950,In_965);
nor U186 (N_186,In_454,In_37);
and U187 (N_187,In_742,In_671);
or U188 (N_188,In_1473,In_1044);
nand U189 (N_189,In_1222,In_215);
or U190 (N_190,In_1187,In_322);
xor U191 (N_191,In_641,In_344);
or U192 (N_192,In_87,In_1106);
or U193 (N_193,In_288,In_1130);
or U194 (N_194,In_544,In_1125);
nand U195 (N_195,In_1287,In_1415);
or U196 (N_196,In_821,In_447);
or U197 (N_197,In_867,In_674);
or U198 (N_198,In_110,In_918);
or U199 (N_199,In_1189,In_566);
nor U200 (N_200,In_976,In_824);
or U201 (N_201,In_496,In_217);
and U202 (N_202,N_88,In_989);
or U203 (N_203,In_589,N_49);
and U204 (N_204,In_1284,In_738);
and U205 (N_205,In_1094,In_180);
and U206 (N_206,N_146,In_1038);
xnor U207 (N_207,N_89,N_57);
nor U208 (N_208,In_1244,In_599);
and U209 (N_209,In_723,In_1273);
and U210 (N_210,In_1135,In_400);
or U211 (N_211,In_320,In_1252);
nand U212 (N_212,In_1123,In_585);
nor U213 (N_213,In_290,In_1085);
nor U214 (N_214,In_501,In_375);
or U215 (N_215,In_1012,In_210);
xnor U216 (N_216,In_1128,In_351);
nand U217 (N_217,In_1404,In_506);
nor U218 (N_218,In_1344,N_108);
or U219 (N_219,In_983,In_1432);
and U220 (N_220,In_991,In_552);
nor U221 (N_221,In_1390,N_170);
xor U222 (N_222,In_494,In_1226);
nand U223 (N_223,In_1194,In_785);
and U224 (N_224,In_125,In_758);
and U225 (N_225,N_198,In_1000);
and U226 (N_226,In_922,In_411);
and U227 (N_227,In_964,In_898);
and U228 (N_228,In_1171,N_124);
nor U229 (N_229,In_829,In_653);
xnor U230 (N_230,In_476,In_336);
nor U231 (N_231,N_47,In_1264);
nand U232 (N_232,N_55,In_205);
nor U233 (N_233,In_1346,In_1365);
nor U234 (N_234,N_32,N_69);
xor U235 (N_235,In_42,In_791);
and U236 (N_236,In_78,In_681);
and U237 (N_237,N_52,In_1442);
xor U238 (N_238,N_138,N_175);
nor U239 (N_239,N_13,N_65);
xor U240 (N_240,In_359,In_990);
and U241 (N_241,In_160,In_357);
or U242 (N_242,In_1055,In_1286);
nor U243 (N_243,N_172,In_413);
nand U244 (N_244,In_568,In_458);
nand U245 (N_245,In_614,N_6);
and U246 (N_246,In_436,In_685);
nand U247 (N_247,In_1469,In_760);
nor U248 (N_248,In_143,In_1051);
and U249 (N_249,N_16,In_1046);
and U250 (N_250,In_348,In_1191);
nor U251 (N_251,In_1486,In_882);
and U252 (N_252,In_576,In_913);
or U253 (N_253,In_1440,In_1045);
nand U254 (N_254,In_949,In_665);
xor U255 (N_255,N_159,In_72);
nor U256 (N_256,In_1481,In_244);
and U257 (N_257,In_1,In_1225);
and U258 (N_258,In_321,In_1140);
nand U259 (N_259,In_1015,N_51);
nor U260 (N_260,In_1299,N_36);
and U261 (N_261,In_522,In_1092);
xnor U262 (N_262,In_557,In_101);
nand U263 (N_263,In_1307,In_944);
xor U264 (N_264,In_107,N_43);
xnor U265 (N_265,N_41,N_189);
nor U266 (N_266,In_750,N_23);
xnor U267 (N_267,In_1120,In_864);
nor U268 (N_268,In_148,In_986);
nand U269 (N_269,In_1387,In_221);
xnor U270 (N_270,In_1172,In_847);
or U271 (N_271,In_1166,In_1197);
nor U272 (N_272,In_731,In_736);
nand U273 (N_273,In_499,In_1435);
nand U274 (N_274,In_277,N_178);
and U275 (N_275,In_339,In_419);
nand U276 (N_276,In_759,In_880);
xnor U277 (N_277,N_83,In_1461);
and U278 (N_278,In_1274,In_1294);
or U279 (N_279,In_970,In_564);
nor U280 (N_280,In_460,In_118);
nand U281 (N_281,In_486,In_762);
nor U282 (N_282,In_828,In_906);
nand U283 (N_283,In_1376,In_1364);
and U284 (N_284,In_708,In_915);
nor U285 (N_285,In_647,In_271);
nor U286 (N_286,In_560,In_1369);
nand U287 (N_287,In_804,In_1183);
nor U288 (N_288,N_54,In_527);
nor U289 (N_289,In_83,N_179);
nand U290 (N_290,In_692,In_1495);
xor U291 (N_291,In_1269,In_429);
or U292 (N_292,In_1023,In_900);
or U293 (N_293,N_91,In_223);
nand U294 (N_294,N_163,In_939);
nand U295 (N_295,In_592,In_13);
nor U296 (N_296,In_963,In_555);
and U297 (N_297,In_49,In_91);
nand U298 (N_298,In_431,N_106);
xor U299 (N_299,In_728,In_630);
xnor U300 (N_300,In_710,In_360);
nand U301 (N_301,In_1288,In_1428);
nor U302 (N_302,In_395,In_453);
nand U303 (N_303,In_391,In_1355);
or U304 (N_304,In_356,In_729);
nor U305 (N_305,In_23,In_899);
nand U306 (N_306,N_63,In_347);
xor U307 (N_307,N_133,In_1242);
and U308 (N_308,In_380,In_1109);
nor U309 (N_309,In_1408,In_423);
nor U310 (N_310,In_669,In_567);
nor U311 (N_311,In_248,In_755);
nand U312 (N_312,In_175,N_67);
and U313 (N_313,In_1033,In_616);
nand U314 (N_314,N_68,In_409);
or U315 (N_315,N_161,In_561);
nand U316 (N_316,In_4,In_1249);
and U317 (N_317,N_114,In_879);
and U318 (N_318,In_63,In_477);
nand U319 (N_319,In_1283,In_784);
xnor U320 (N_320,In_715,In_444);
or U321 (N_321,In_1202,In_105);
and U322 (N_322,In_1483,In_1449);
or U323 (N_323,In_1360,In_1113);
nor U324 (N_324,In_254,In_730);
nand U325 (N_325,N_66,In_1400);
and U326 (N_326,In_1380,N_0);
and U327 (N_327,In_1313,In_831);
xor U328 (N_328,In_1347,In_1377);
and U329 (N_329,In_1169,In_503);
and U330 (N_330,N_79,In_795);
and U331 (N_331,In_1453,In_245);
nor U332 (N_332,In_1447,In_1235);
nor U333 (N_333,In_919,In_1164);
and U334 (N_334,In_741,In_632);
or U335 (N_335,In_261,In_109);
nand U336 (N_336,N_15,In_933);
nor U337 (N_337,In_1117,In_645);
nand U338 (N_338,In_740,In_1427);
xnor U339 (N_339,In_537,In_240);
nand U340 (N_340,In_775,In_1084);
and U341 (N_341,N_137,In_1195);
and U342 (N_342,N_101,N_153);
nand U343 (N_343,In_743,In_908);
xnor U344 (N_344,In_1070,In_1218);
nor U345 (N_345,In_154,In_607);
nor U346 (N_346,In_524,In_1208);
nand U347 (N_347,N_185,In_298);
or U348 (N_348,N_192,N_145);
nand U349 (N_349,In_1379,In_2);
nand U350 (N_350,In_172,In_74);
xor U351 (N_351,In_41,In_1268);
nand U352 (N_352,In_1230,In_757);
and U353 (N_353,In_280,N_10);
nor U354 (N_354,In_858,In_1102);
or U355 (N_355,In_1303,In_1475);
and U356 (N_356,In_514,In_408);
xor U357 (N_357,In_734,In_818);
nand U358 (N_358,N_31,In_372);
nand U359 (N_359,In_489,In_250);
nor U360 (N_360,In_786,In_425);
nand U361 (N_361,In_1203,In_1156);
nand U362 (N_362,In_1209,N_53);
xnor U363 (N_363,In_1457,In_58);
xor U364 (N_364,In_994,N_197);
xor U365 (N_365,In_1295,N_156);
nor U366 (N_366,In_451,In_378);
nor U367 (N_367,In_1492,In_659);
xnor U368 (N_368,In_1458,In_529);
nor U369 (N_369,N_24,In_512);
and U370 (N_370,In_1131,In_393);
xor U371 (N_371,N_166,In_534);
nand U372 (N_372,In_1076,In_1318);
and U373 (N_373,In_428,In_540);
and U374 (N_374,In_293,In_559);
nand U375 (N_375,In_1314,In_1143);
xor U376 (N_376,In_115,In_211);
xnor U377 (N_377,In_1470,In_497);
nand U378 (N_378,In_403,N_46);
or U379 (N_379,In_266,In_464);
and U380 (N_380,In_800,In_1030);
xnor U381 (N_381,In_222,In_1395);
xnor U382 (N_382,In_365,In_1093);
nor U383 (N_383,In_385,In_1316);
nand U384 (N_384,N_5,In_407);
and U385 (N_385,In_1352,In_156);
nor U386 (N_386,In_850,In_672);
nand U387 (N_387,In_718,In_761);
or U388 (N_388,In_326,N_60);
and U389 (N_389,In_249,In_1139);
and U390 (N_390,In_191,In_1494);
nor U391 (N_391,In_1477,In_848);
and U392 (N_392,In_664,In_427);
xnor U393 (N_393,In_155,In_625);
or U394 (N_394,In_683,N_7);
xor U395 (N_395,In_981,In_1231);
nand U396 (N_396,N_11,In_866);
xnor U397 (N_397,In_136,In_25);
xnor U398 (N_398,In_657,In_8);
nand U399 (N_399,In_780,In_1382);
nand U400 (N_400,In_334,N_56);
nand U401 (N_401,In_163,In_171);
nor U402 (N_402,N_302,In_3);
or U403 (N_403,In_655,In_799);
or U404 (N_404,In_1391,N_385);
nand U405 (N_405,In_954,In_1122);
nor U406 (N_406,In_811,In_1234);
nor U407 (N_407,N_210,In_1411);
nand U408 (N_408,In_333,In_505);
nor U409 (N_409,In_1271,In_714);
or U410 (N_410,In_415,In_1052);
nand U411 (N_411,In_677,N_167);
xor U412 (N_412,N_278,In_328);
nand U413 (N_413,In_270,N_381);
nand U414 (N_414,In_1054,In_169);
nand U415 (N_415,In_937,N_382);
nand U416 (N_416,In_1251,N_109);
and U417 (N_417,N_144,In_79);
nand U418 (N_418,In_1168,In_102);
nor U419 (N_419,N_364,In_556);
nor U420 (N_420,N_240,N_241);
xnor U421 (N_421,N_202,N_86);
or U422 (N_422,N_44,N_366);
or U423 (N_423,In_285,In_1091);
and U424 (N_424,N_256,N_295);
and U425 (N_425,In_739,N_247);
xor U426 (N_426,In_1049,In_170);
nand U427 (N_427,In_548,In_327);
nand U428 (N_428,In_620,In_1104);
or U429 (N_429,In_259,In_133);
xor U430 (N_430,N_64,N_226);
nor U431 (N_431,In_1329,N_254);
and U432 (N_432,In_1392,N_351);
and U433 (N_433,N_150,In_340);
nand U434 (N_434,In_243,In_264);
xor U435 (N_435,N_184,N_76);
or U436 (N_436,N_152,N_18);
or U437 (N_437,In_1456,N_277);
nand U438 (N_438,In_445,In_1285);
and U439 (N_439,In_104,In_805);
xnor U440 (N_440,N_239,In_1336);
nor U441 (N_441,In_1311,In_1111);
nand U442 (N_442,In_456,In_935);
and U443 (N_443,In_1384,In_1138);
and U444 (N_444,In_1389,In_1196);
or U445 (N_445,N_151,In_1201);
nor U446 (N_446,In_751,In_1147);
or U447 (N_447,In_1089,N_50);
xnor U448 (N_448,N_328,In_907);
nor U449 (N_449,In_1351,N_232);
xnor U450 (N_450,N_211,In_1036);
xnor U451 (N_451,In_470,N_314);
nor U452 (N_452,In_891,In_60);
and U453 (N_453,N_111,N_307);
or U454 (N_454,In_1116,In_776);
nand U455 (N_455,N_228,In_928);
xnor U456 (N_456,In_840,N_119);
or U457 (N_457,In_1446,In_377);
or U458 (N_458,In_600,In_93);
nand U459 (N_459,In_1214,N_315);
and U460 (N_460,N_316,In_1124);
xor U461 (N_461,N_289,In_158);
nor U462 (N_462,N_306,In_574);
nor U463 (N_463,In_1388,In_448);
xor U464 (N_464,In_570,In_819);
xor U465 (N_465,In_1338,In_1256);
and U466 (N_466,In_1320,In_1080);
xor U467 (N_467,In_1067,N_168);
or U468 (N_468,In_1060,N_392);
nand U469 (N_469,In_837,In_130);
xnor U470 (N_470,In_1073,In_370);
or U471 (N_471,In_189,N_267);
nand U472 (N_472,In_397,N_107);
nor U473 (N_473,N_213,In_577);
nand U474 (N_474,N_141,N_321);
nand U475 (N_475,In_1173,In_1163);
and U476 (N_476,In_493,In_146);
xor U477 (N_477,In_1366,In_1072);
or U478 (N_478,N_182,N_281);
nand U479 (N_479,In_446,In_345);
nand U480 (N_480,N_73,In_654);
xor U481 (N_481,In_835,In_198);
nor U482 (N_482,In_1438,In_449);
nor U483 (N_483,In_467,In_88);
nand U484 (N_484,In_1363,In_845);
nand U485 (N_485,In_1247,In_565);
nor U486 (N_486,In_161,N_207);
or U487 (N_487,In_596,N_177);
or U488 (N_488,In_1028,In_701);
xnor U489 (N_489,In_178,In_917);
xor U490 (N_490,In_745,In_690);
or U491 (N_491,In_587,N_253);
and U492 (N_492,In_726,In_305);
xor U493 (N_493,In_1399,N_374);
nor U494 (N_494,N_129,N_234);
nand U495 (N_495,N_348,In_901);
xor U496 (N_496,In_40,In_520);
and U497 (N_497,In_1061,N_251);
xnor U498 (N_498,In_1361,N_287);
and U499 (N_499,In_704,In_980);
or U500 (N_500,N_378,N_22);
xnor U501 (N_501,In_1409,In_1184);
nor U502 (N_502,N_263,In_765);
nor U503 (N_503,In_1174,N_48);
nand U504 (N_504,N_359,In_1448);
nand U505 (N_505,In_865,N_78);
or U506 (N_506,In_693,In_1454);
and U507 (N_507,In_1029,N_270);
nor U508 (N_508,N_353,In_984);
nor U509 (N_509,In_1158,In_492);
nand U510 (N_510,In_31,In_422);
and U511 (N_511,In_606,N_12);
xor U512 (N_512,In_466,In_1132);
or U513 (N_513,N_395,N_208);
or U514 (N_514,N_70,In_575);
or U515 (N_515,N_252,In_1095);
and U516 (N_516,In_868,In_116);
nor U517 (N_517,In_287,In_364);
nand U518 (N_518,In_229,N_187);
xnor U519 (N_519,In_810,In_1310);
and U520 (N_520,In_1141,N_221);
nand U521 (N_521,In_10,N_25);
nor U522 (N_522,In_1480,In_603);
xor U523 (N_523,In_924,N_384);
nand U524 (N_524,In_1385,In_1204);
xnor U525 (N_525,N_349,N_126);
nand U526 (N_526,In_367,In_1345);
xnor U527 (N_527,N_99,In_1424);
xor U528 (N_528,In_1035,N_304);
and U529 (N_529,In_111,In_443);
or U530 (N_530,In_97,In_1167);
and U531 (N_531,In_1383,In_618);
xnor U532 (N_532,In_1176,In_173);
nand U533 (N_533,N_199,In_1455);
or U534 (N_534,In_376,In_1025);
xor U535 (N_535,In_1498,In_1292);
xor U536 (N_536,In_504,In_911);
nand U537 (N_537,N_97,In_114);
nand U538 (N_538,In_744,In_61);
xor U539 (N_539,N_193,In_1373);
and U540 (N_540,N_87,In_474);
xor U541 (N_541,N_203,N_265);
or U542 (N_542,In_309,In_551);
nand U543 (N_543,In_1188,In_274);
xor U544 (N_544,N_105,In_1300);
nand U545 (N_545,In_792,In_324);
and U546 (N_546,N_357,N_102);
nor U547 (N_547,N_125,In_815);
and U548 (N_548,In_1332,In_313);
or U549 (N_549,In_1108,N_90);
and U550 (N_550,In_52,In_1484);
nand U551 (N_551,In_262,In_1068);
nand U552 (N_552,In_962,In_549);
xor U553 (N_553,In_770,N_45);
nand U554 (N_554,In_1177,In_113);
and U555 (N_555,N_311,In_119);
and U556 (N_556,N_201,In_1069);
or U557 (N_557,N_93,In_306);
xor U558 (N_558,N_243,In_874);
or U559 (N_559,N_110,N_20);
or U560 (N_560,In_1356,In_1426);
and U561 (N_561,In_793,In_267);
nor U562 (N_562,In_121,In_1261);
nand U563 (N_563,In_601,In_144);
nand U564 (N_564,N_206,In_1293);
or U565 (N_565,In_515,In_1343);
or U566 (N_566,N_338,In_1009);
nand U567 (N_567,N_29,In_1460);
nor U568 (N_568,In_193,In_995);
or U569 (N_569,In_1375,In_887);
xor U570 (N_570,In_1151,In_1083);
and U571 (N_571,N_332,N_370);
nor U572 (N_572,In_44,In_137);
and U573 (N_573,In_510,In_252);
nor U574 (N_574,In_361,N_282);
and U575 (N_575,In_531,N_269);
nor U576 (N_576,In_14,In_482);
xnor U577 (N_577,N_235,In_1393);
and U578 (N_578,In_325,In_1037);
xnor U579 (N_579,In_1014,In_1110);
xor U580 (N_580,In_1419,In_586);
or U581 (N_581,In_85,In_335);
xnor U582 (N_582,N_355,In_1330);
nor U583 (N_583,In_1452,In_1362);
and U584 (N_584,N_297,In_263);
nor U585 (N_585,N_181,N_219);
nand U586 (N_586,In_442,In_622);
and U587 (N_587,In_553,In_862);
nand U588 (N_588,In_1229,In_1118);
and U589 (N_589,N_223,In_164);
and U590 (N_590,In_92,N_292);
nor U591 (N_591,In_203,In_106);
or U592 (N_592,In_711,In_207);
xnor U593 (N_593,N_95,N_339);
xnor U594 (N_594,In_1472,In_1056);
xor U595 (N_595,N_305,In_1266);
xnor U596 (N_596,In_1368,N_323);
or U597 (N_597,In_1465,In_1220);
nor U598 (N_598,In_462,In_1103);
xor U599 (N_599,In_1474,In_490);
xor U600 (N_600,N_276,N_204);
xnor U601 (N_601,In_1405,In_885);
xnor U602 (N_602,In_890,N_38);
xor U603 (N_603,N_429,N_454);
nor U604 (N_604,In_1048,In_593);
nor U605 (N_605,N_231,N_416);
and U606 (N_606,In_1043,N_587);
or U607 (N_607,N_128,N_532);
or U608 (N_608,In_675,In_640);
and U609 (N_609,In_484,N_412);
and U610 (N_610,N_363,In_519);
xnor U611 (N_611,N_431,N_324);
and U612 (N_612,In_967,In_1443);
xnor U613 (N_613,N_434,In_916);
and U614 (N_614,N_75,In_604);
nor U615 (N_615,In_209,N_537);
nand U616 (N_616,In_637,In_816);
nor U617 (N_617,In_279,N_318);
and U618 (N_618,In_1324,N_552);
nor U619 (N_619,In_554,In_1008);
nor U620 (N_620,N_212,In_219);
and U621 (N_621,In_153,N_317);
or U622 (N_622,N_597,N_379);
nand U623 (N_623,N_411,In_1401);
nand U624 (N_624,In_174,In_846);
and U625 (N_625,In_809,N_248);
nand U626 (N_626,In_602,In_778);
or U627 (N_627,N_176,N_42);
and U628 (N_628,N_398,N_346);
and U629 (N_629,N_402,N_9);
xor U630 (N_630,In_28,N_335);
nor U631 (N_631,N_424,In_182);
nor U632 (N_632,N_465,In_81);
and U633 (N_633,N_140,In_851);
nand U634 (N_634,In_747,N_565);
xnor U635 (N_635,In_941,N_471);
xnor U636 (N_636,In_128,N_1);
nor U637 (N_637,In_258,In_1267);
or U638 (N_638,N_116,N_40);
xor U639 (N_639,N_345,In_140);
and U640 (N_640,In_312,In_966);
and U641 (N_641,N_139,N_476);
and U642 (N_642,In_1086,In_236);
nor U643 (N_643,In_488,In_401);
or U644 (N_644,In_571,N_477);
xor U645 (N_645,In_709,N_422);
or U646 (N_646,N_444,N_571);
or U647 (N_647,In_807,In_886);
xor U648 (N_648,N_325,In_1423);
nor U649 (N_649,N_365,N_403);
nor U650 (N_650,In_689,N_290);
or U651 (N_651,N_485,In_580);
nand U652 (N_652,N_122,In_947);
and U653 (N_653,In_168,N_196);
nor U654 (N_654,N_410,N_438);
nand U655 (N_655,N_433,In_1211);
or U656 (N_656,N_469,In_1075);
xnor U657 (N_657,In_583,N_550);
xor U658 (N_658,N_274,In_902);
nor U659 (N_659,N_480,N_200);
nand U660 (N_660,In_1101,N_113);
and U661 (N_661,N_377,N_418);
nand U662 (N_662,In_165,N_4);
and U663 (N_663,N_127,In_643);
and U664 (N_664,N_216,In_404);
and U665 (N_665,In_680,In_275);
and U666 (N_666,In_952,N_442);
xor U667 (N_667,In_781,In_1057);
and U668 (N_668,N_82,In_35);
and U669 (N_669,In_414,In_1021);
nand U670 (N_670,In_943,In_1039);
and U671 (N_671,In_498,N_591);
or U672 (N_672,N_244,In_200);
and U673 (N_673,N_487,In_696);
nor U674 (N_674,In_749,N_132);
xnor U675 (N_675,N_186,N_527);
nor U676 (N_676,In_957,In_808);
and U677 (N_677,N_333,In_871);
nor U678 (N_678,In_398,N_308);
nor U679 (N_679,N_387,In_1321);
nor U680 (N_680,In_1127,In_1437);
xnor U681 (N_681,N_120,N_81);
and U682 (N_682,N_503,N_34);
xnor U683 (N_683,N_559,In_145);
nor U684 (N_684,N_313,N_522);
nor U685 (N_685,In_546,N_458);
or U686 (N_686,In_69,N_507);
nand U687 (N_687,In_430,N_298);
or U688 (N_688,N_59,In_350);
or U689 (N_689,N_233,In_22);
nor U690 (N_690,In_1199,In_491);
nand U691 (N_691,N_589,In_629);
nor U692 (N_692,In_355,N_375);
or U693 (N_693,N_312,In_706);
nand U694 (N_694,N_14,N_104);
or U695 (N_695,In_969,N_330);
nor U696 (N_696,In_438,In_57);
nor U697 (N_697,N_533,N_347);
and U698 (N_698,In_1193,N_356);
and U699 (N_699,N_436,In_628);
nand U700 (N_700,N_94,N_553);
or U701 (N_701,In_1312,N_486);
nor U702 (N_702,N_396,In_558);
nor U703 (N_703,N_386,In_459);
xnor U704 (N_704,In_1398,In_635);
or U705 (N_705,In_224,N_37);
or U706 (N_706,N_100,In_132);
nand U707 (N_707,N_517,N_294);
nand U708 (N_708,N_508,N_275);
or U709 (N_709,N_407,In_697);
or U710 (N_710,N_456,N_563);
nor U711 (N_711,N_92,In_337);
or U712 (N_712,In_399,In_1002);
and U713 (N_713,In_500,In_611);
and U714 (N_714,N_340,In_295);
xor U715 (N_715,In_341,N_582);
xor U716 (N_716,N_147,In_1281);
nand U717 (N_717,In_300,In_861);
and U718 (N_718,N_584,N_336);
or U719 (N_719,In_382,N_404);
nand U720 (N_720,In_1263,In_432);
nor U721 (N_721,In_7,N_462);
xnor U722 (N_722,N_142,N_473);
nand U723 (N_723,In_1018,In_227);
or U724 (N_724,In_1207,In_581);
or U725 (N_725,In_974,In_1331);
xor U726 (N_726,In_598,In_289);
nor U727 (N_727,N_447,N_490);
nor U728 (N_728,N_296,N_540);
nand U729 (N_729,N_390,In_12);
and U730 (N_730,In_406,N_136);
or U731 (N_731,N_326,In_1348);
nand U732 (N_732,N_593,In_541);
xor U733 (N_733,In_1496,N_28);
nor U734 (N_734,N_595,N_470);
nand U735 (N_735,In_1291,In_1259);
nand U736 (N_736,N_393,In_384);
xor U737 (N_737,N_368,N_174);
or U738 (N_738,N_420,N_350);
and U739 (N_739,In_70,N_148);
xor U740 (N_740,In_1232,N_502);
nor U741 (N_741,In_1298,N_521);
xnor U742 (N_742,In_884,In_1178);
nor U743 (N_743,N_195,In_538);
nand U744 (N_744,In_291,In_953);
xnor U745 (N_745,In_1394,In_853);
nand U746 (N_746,In_1471,In_1024);
xor U747 (N_747,In_1414,In_797);
nand U748 (N_748,N_548,N_513);
nor U749 (N_749,In_1397,N_575);
or U750 (N_750,In_255,In_1162);
and U751 (N_751,In_80,In_1159);
nor U752 (N_752,In_876,In_1357);
xnor U753 (N_753,N_115,In_992);
nor U754 (N_754,In_1459,N_288);
nand U755 (N_755,In_1490,In_386);
nand U756 (N_756,In_301,In_1433);
nor U757 (N_757,In_713,In_103);
nand U758 (N_758,N_358,In_303);
xnor U759 (N_759,N_421,N_229);
and U760 (N_760,N_236,In_1062);
nor U761 (N_761,In_687,N_467);
or U762 (N_762,In_1257,N_84);
xnor U763 (N_763,In_1100,N_536);
xor U764 (N_764,In_597,N_529);
nor U765 (N_765,In_1153,N_520);
nand U766 (N_766,N_439,In_694);
and U767 (N_767,In_420,In_782);
nor U768 (N_768,In_502,In_1238);
nor U769 (N_769,In_1482,N_322);
nor U770 (N_770,In_316,In_1180);
and U771 (N_771,N_549,In_646);
or U772 (N_772,In_1491,In_1179);
nand U773 (N_773,In_721,In_183);
or U774 (N_774,In_257,In_507);
nand U775 (N_775,N_169,In_1381);
and U776 (N_776,N_371,N_238);
xnor U777 (N_777,In_27,N_506);
nor U778 (N_778,In_134,N_30);
xnor U779 (N_779,N_405,In_65);
or U780 (N_780,In_1262,In_468);
xnor U781 (N_781,N_117,N_245);
or U782 (N_782,N_310,N_227);
xnor U783 (N_783,In_1476,N_523);
xor U784 (N_784,N_453,N_594);
nand U785 (N_785,In_302,In_914);
nand U786 (N_786,In_1371,In_71);
nor U787 (N_787,In_1478,In_1227);
or U788 (N_788,In_1250,In_1396);
and U789 (N_789,In_389,In_1279);
nor U790 (N_790,N_514,N_441);
and U791 (N_791,In_894,In_936);
xnor U792 (N_792,N_586,N_242);
and U793 (N_793,N_134,In_1078);
or U794 (N_794,N_217,In_700);
xor U795 (N_795,In_225,N_445);
nor U796 (N_796,N_479,In_1219);
nor U797 (N_797,N_261,In_1040);
xor U798 (N_798,In_667,N_33);
nand U799 (N_799,N_448,N_246);
and U800 (N_800,N_376,N_257);
or U801 (N_801,N_214,In_1412);
or U802 (N_802,N_602,N_555);
xor U803 (N_803,N_657,N_629);
or U804 (N_804,In_579,N_743);
or U805 (N_805,In_1149,In_813);
xor U806 (N_806,N_459,N_642);
nor U807 (N_807,In_1306,In_1010);
and U808 (N_808,In_1190,N_720);
nor U809 (N_809,N_215,In_1358);
nor U810 (N_810,N_524,In_433);
nor U811 (N_811,In_201,N_708);
nor U812 (N_812,In_1258,In_1047);
xnor U813 (N_813,In_54,N_249);
xnor U814 (N_814,In_353,N_483);
nand U815 (N_815,N_568,N_783);
nor U816 (N_816,In_338,N_709);
nor U817 (N_817,In_1087,N_573);
and U818 (N_818,N_671,In_956);
xor U819 (N_819,N_621,N_696);
nand U820 (N_820,In_247,In_479);
nor U821 (N_821,N_654,In_1302);
nand U822 (N_822,In_772,N_615);
nand U823 (N_823,N_674,N_640);
nand U824 (N_824,N_676,N_588);
or U825 (N_825,N_601,In_202);
nor U826 (N_826,In_595,N_500);
or U827 (N_827,In_1160,In_1349);
or U828 (N_828,In_732,N_341);
and U829 (N_829,In_895,N_612);
nor U830 (N_830,N_225,In_1142);
and U831 (N_831,N_191,N_303);
nand U832 (N_832,In_1145,In_543);
and U833 (N_833,N_435,N_659);
and U834 (N_834,N_391,N_772);
xnor U835 (N_835,N_272,N_3);
nand U836 (N_836,N_637,In_1420);
and U837 (N_837,In_342,N_693);
and U838 (N_838,N_689,N_534);
nand U839 (N_839,N_598,N_747);
nor U840 (N_840,N_85,In_1175);
or U841 (N_841,In_651,N_285);
nand U842 (N_842,In_166,N_730);
and U843 (N_843,N_634,N_690);
nand U844 (N_844,In_45,N_451);
xor U845 (N_845,N_691,N_526);
nand U846 (N_846,N_596,N_319);
nor U847 (N_847,N_798,N_380);
nand U848 (N_848,In_475,N_17);
and U849 (N_849,In_609,N_577);
nand U850 (N_850,N_599,In_450);
nand U851 (N_851,In_1462,N_103);
and U852 (N_852,N_670,In_768);
and U853 (N_853,In_47,In_1237);
nor U854 (N_854,In_631,N_343);
nand U855 (N_855,In_875,In_487);
or U856 (N_856,N_774,N_130);
or U857 (N_857,N_749,In_77);
and U858 (N_858,In_783,N_286);
and U859 (N_859,In_1224,N_188);
or U860 (N_860,N_682,N_663);
xor U861 (N_861,N_342,In_284);
nor U862 (N_862,In_6,N_781);
xor U863 (N_863,N_677,N_645);
nor U864 (N_864,N_679,N_80);
xnor U865 (N_865,In_396,N_773);
xor U866 (N_866,N_474,In_1144);
nand U867 (N_867,N_644,N_408);
xor U868 (N_868,N_578,N_790);
and U869 (N_869,N_625,N_668);
nand U870 (N_870,N_780,In_1019);
nand U871 (N_871,In_131,N_171);
and U872 (N_872,N_722,N_771);
nand U873 (N_873,In_1236,N_698);
or U874 (N_874,N_320,N_260);
xor U875 (N_875,In_621,N_604);
and U876 (N_876,N_739,In_346);
or U877 (N_877,In_662,N_190);
nand U878 (N_878,In_1319,N_764);
and U879 (N_879,N_543,N_535);
xnor U880 (N_880,N_425,N_516);
nand U881 (N_881,N_766,In_912);
nand U882 (N_882,In_177,In_1489);
or U883 (N_883,In_903,N_583);
nand U884 (N_884,N_58,N_567);
and U885 (N_885,In_722,N_700);
or U886 (N_886,N_501,In_228);
or U887 (N_887,In_323,In_1097);
nand U888 (N_888,In_1466,In_297);
xor U889 (N_889,In_961,In_418);
nand U890 (N_890,In_842,N_717);
xor U891 (N_891,N_760,In_124);
nor U892 (N_892,N_694,In_1114);
or U893 (N_893,N_194,In_716);
or U894 (N_894,In_213,In_613);
nor U895 (N_895,N_482,In_1467);
nor U896 (N_896,N_74,N_8);
and U897 (N_897,In_273,In_1421);
xnor U898 (N_898,In_373,N_788);
xor U899 (N_899,N_660,N_667);
and U900 (N_900,N_778,N_711);
nor U901 (N_901,In_695,In_1137);
and U902 (N_902,N_491,N_160);
nor U903 (N_903,In_855,N_554);
or U904 (N_904,N_389,N_752);
nor U905 (N_905,N_98,N_611);
nor U906 (N_906,In_318,In_1485);
nor U907 (N_907,In_352,In_188);
xnor U908 (N_908,N_273,In_167);
or U909 (N_909,In_232,N_515);
nand U910 (N_910,N_149,In_752);
and U911 (N_911,N_361,N_528);
nor U912 (N_912,N_61,N_712);
or U913 (N_913,In_663,N_455);
xnor U914 (N_914,N_539,N_792);
nor U915 (N_915,N_538,N_754);
xor U916 (N_916,N_409,In_194);
xor U917 (N_917,N_542,N_546);
nor U918 (N_918,N_603,N_279);
or U919 (N_919,N_570,In_1304);
nor U920 (N_920,In_18,N_547);
nand U921 (N_921,In_702,In_195);
nand U922 (N_922,N_489,In_754);
xnor U923 (N_923,N_419,In_978);
nand U924 (N_924,In_1245,N_569);
nor U925 (N_925,N_666,N_770);
and U926 (N_926,In_658,N_96);
and U927 (N_927,In_402,In_705);
nand U928 (N_928,In_21,N_763);
and U929 (N_929,N_449,N_647);
nor U930 (N_930,In_1337,N_796);
nor U931 (N_931,N_544,In_299);
xor U932 (N_932,N_673,In_973);
and U933 (N_933,N_776,N_618);
nand U934 (N_934,In_920,N_481);
xnor U935 (N_935,In_699,In_1328);
nand U936 (N_936,In_1353,N_745);
nand U937 (N_937,N_669,In_1297);
xor U938 (N_938,N_518,In_483);
nor U939 (N_939,N_610,In_437);
xor U940 (N_940,N_750,In_362);
xnor U941 (N_941,N_748,N_639);
nand U942 (N_942,In_278,N_684);
and U943 (N_943,N_545,N_630);
xor U944 (N_944,In_666,N_131);
nor U945 (N_945,N_579,N_427);
and U946 (N_946,In_830,In_1325);
or U947 (N_947,N_291,In_1198);
nor U948 (N_948,In_789,In_605);
or U949 (N_949,In_197,N_672);
xnor U950 (N_950,In_473,In_1280);
and U951 (N_951,N_793,N_707);
xor U952 (N_952,N_664,N_413);
xor U953 (N_953,N_632,N_466);
or U954 (N_954,N_665,N_782);
or U955 (N_955,N_692,N_701);
or U956 (N_956,N_755,N_728);
xnor U957 (N_957,N_255,In_572);
xnor U958 (N_958,In_1088,N_706);
nor U959 (N_959,N_680,N_736);
nor U960 (N_960,N_299,N_746);
xor U961 (N_961,N_562,N_797);
and U962 (N_962,N_705,N_725);
nor U963 (N_963,N_649,In_135);
nand U964 (N_964,N_121,In_1205);
nand U965 (N_965,N_581,N_661);
nand U966 (N_966,N_505,N_271);
or U967 (N_967,N_399,N_498);
or U968 (N_968,N_777,In_998);
nand U969 (N_969,In_230,N_606);
or U970 (N_970,N_572,N_430);
nor U971 (N_971,N_617,N_112);
nor U972 (N_972,In_112,In_526);
xor U973 (N_973,In_1445,N_627);
xor U974 (N_974,In_11,N_230);
and U975 (N_975,In_1374,N_468);
or U976 (N_976,In_670,In_1277);
or U977 (N_977,In_59,In_725);
nand U978 (N_978,N_721,N_283);
nor U979 (N_979,N_354,In_547);
nor U980 (N_980,N_557,N_494);
nand U981 (N_981,N_556,N_638);
or U982 (N_982,N_686,N_662);
nand U983 (N_983,N_608,In_120);
nor U984 (N_984,N_220,N_723);
and U985 (N_985,N_443,In_349);
nand U986 (N_986,In_1133,N_768);
and U987 (N_987,N_264,N_394);
and U988 (N_988,N_687,N_729);
nor U989 (N_989,In_686,In_417);
or U990 (N_990,N_180,In_712);
nand U991 (N_991,In_1115,N_756);
xor U992 (N_992,N_280,N_293);
xor U993 (N_993,N_695,N_735);
and U994 (N_994,N_699,In_387);
nor U995 (N_995,N_704,In_1050);
and U996 (N_996,N_268,N_600);
xor U997 (N_997,N_432,In_465);
nand U998 (N_998,In_844,N_19);
nor U999 (N_999,In_893,In_563);
xor U1000 (N_1000,N_900,In_1429);
nor U1001 (N_1001,N_904,In_926);
and U1002 (N_1002,N_787,In_96);
nand U1003 (N_1003,N_975,N_899);
or U1004 (N_1004,N_968,In_971);
or U1005 (N_1005,N_915,N_903);
or U1006 (N_1006,N_813,N_902);
or U1007 (N_1007,N_834,N_616);
nand U1008 (N_1008,N_224,N_864);
nor U1009 (N_1009,In_1444,In_1378);
or U1010 (N_1010,In_717,N_831);
nor U1011 (N_1011,N_566,N_26);
nand U1012 (N_1012,N_683,N_947);
and U1013 (N_1013,N_825,N_919);
nor U1014 (N_1014,N_35,In_480);
or U1015 (N_1015,N_938,N_803);
nand U1016 (N_1016,N_804,N_950);
xor U1017 (N_1017,N_872,In_1011);
nor U1018 (N_1018,N_809,In_206);
and U1019 (N_1019,N_876,N_964);
nand U1020 (N_1020,N_926,N_525);
nor U1021 (N_1021,N_414,N_258);
and U1022 (N_1022,N_165,N_948);
nand U1023 (N_1023,N_762,N_731);
nor U1024 (N_1024,N_724,N_991);
nand U1025 (N_1025,N_337,In_142);
xor U1026 (N_1026,In_242,N_519);
nor U1027 (N_1027,N_822,N_893);
nand U1028 (N_1028,In_1240,N_646);
nand U1029 (N_1029,N_590,N_811);
xor U1030 (N_1030,N_605,N_561);
nand U1031 (N_1031,N_262,N_967);
xor U1032 (N_1032,N_955,N_732);
nor U1033 (N_1033,N_879,N_984);
or U1034 (N_1034,N_987,N_888);
nand U1035 (N_1035,N_844,In_878);
and U1036 (N_1036,N_388,N_623);
xor U1037 (N_1037,N_937,N_785);
and U1038 (N_1038,N_123,N_440);
xnor U1039 (N_1039,N_767,N_923);
nor U1040 (N_1040,N_958,N_871);
nand U1041 (N_1041,N_758,N_259);
or U1042 (N_1042,In_1479,N_775);
nand U1043 (N_1043,N_877,N_367);
xor U1044 (N_1044,N_656,N_821);
xor U1045 (N_1045,N_607,N_450);
nand U1046 (N_1046,N_940,N_918);
nor U1047 (N_1047,N_817,N_965);
nor U1048 (N_1048,In_75,In_979);
and U1049 (N_1049,N_946,N_914);
nor U1050 (N_1050,N_769,In_67);
nand U1051 (N_1051,N_887,N_913);
xor U1052 (N_1052,N_77,N_928);
nor U1053 (N_1053,N_971,N_2);
xnor U1054 (N_1054,In_573,N_908);
and U1055 (N_1055,N_925,In_1241);
and U1056 (N_1056,N_718,N_805);
nand U1057 (N_1057,N_626,N_753);
and U1058 (N_1058,N_860,N_886);
and U1059 (N_1059,In_746,In_94);
and U1060 (N_1060,N_631,N_905);
nand U1061 (N_1061,N_558,In_1301);
nand U1062 (N_1062,N_868,N_504);
xor U1063 (N_1063,N_855,N_820);
xnor U1064 (N_1064,In_1181,In_724);
or U1065 (N_1065,In_1340,N_154);
or U1066 (N_1066,N_653,N_941);
nand U1067 (N_1067,N_497,N_818);
nor U1068 (N_1068,N_799,In_90);
and U1069 (N_1069,In_1186,N_158);
nor U1070 (N_1070,N_741,N_417);
nor U1071 (N_1071,N_806,N_651);
nor U1072 (N_1072,N_857,N_300);
nor U1073 (N_1073,N_499,N_944);
xnor U1074 (N_1074,In_138,In_435);
and U1075 (N_1075,N_765,N_976);
and U1076 (N_1076,N_585,N_352);
or U1077 (N_1077,N_426,In_626);
nor U1078 (N_1078,N_636,In_1031);
and U1079 (N_1079,N_824,N_716);
nand U1080 (N_1080,N_173,In_1129);
and U1081 (N_1081,N_530,N_878);
and U1082 (N_1082,N_863,N_209);
xor U1083 (N_1083,N_492,In_788);
xnor U1084 (N_1084,N_815,In_186);
nor U1085 (N_1085,In_147,N_833);
xor U1086 (N_1086,N_998,N_344);
or U1087 (N_1087,N_898,N_861);
or U1088 (N_1088,In_187,N_284);
nand U1089 (N_1089,In_424,In_1246);
or U1090 (N_1090,N_845,N_942);
xnor U1091 (N_1091,In_265,N_870);
and U1092 (N_1092,N_423,In_1077);
nand U1093 (N_1093,In_226,N_945);
xnor U1094 (N_1094,N_970,N_164);
nor U1095 (N_1095,N_850,N_463);
nor U1096 (N_1096,N_727,In_841);
and U1097 (N_1097,N_369,N_678);
nand U1098 (N_1098,N_633,N_891);
nor U1099 (N_1099,In_542,N_496);
nand U1100 (N_1100,In_1248,N_966);
xnor U1101 (N_1101,In_536,N_71);
or U1102 (N_1102,N_428,N_560);
xnor U1103 (N_1103,N_960,N_327);
nor U1104 (N_1104,In_1350,In_1013);
xor U1105 (N_1105,N_802,N_744);
nor U1106 (N_1106,N_334,N_962);
nor U1107 (N_1107,N_922,N_801);
and U1108 (N_1108,N_911,N_460);
xnor U1109 (N_1109,N_974,N_874);
or U1110 (N_1110,In_452,In_95);
or U1111 (N_1111,N_954,In_1260);
nand U1112 (N_1112,N_929,N_856);
xnor U1113 (N_1113,In_179,N_866);
or U1114 (N_1114,N_488,N_27);
and U1115 (N_1115,N_851,N_650);
or U1116 (N_1116,N_784,N_383);
and U1117 (N_1117,N_837,N_789);
nand U1118 (N_1118,N_541,N_995);
nor U1119 (N_1119,N_973,N_840);
or U1120 (N_1120,N_959,In_888);
and U1121 (N_1121,In_388,In_390);
xor U1122 (N_1122,N_493,N_400);
xnor U1123 (N_1123,N_935,N_574);
nor U1124 (N_1124,N_619,In_987);
and U1125 (N_1125,N_401,N_972);
nand U1126 (N_1126,In_827,N_183);
xor U1127 (N_1127,N_927,N_862);
xnor U1128 (N_1128,N_823,In_1253);
and U1129 (N_1129,N_266,N_362);
and U1130 (N_1130,N_658,In_192);
xor U1131 (N_1131,N_143,In_932);
nor U1132 (N_1132,N_643,N_884);
or U1133 (N_1133,N_816,N_994);
nand U1134 (N_1134,N_858,N_910);
and U1135 (N_1135,N_511,N_949);
xnor U1136 (N_1136,N_881,N_437);
nand U1137 (N_1137,N_963,In_26);
xor U1138 (N_1138,In_972,N_702);
xor U1139 (N_1139,In_1063,N_807);
nand U1140 (N_1140,N_648,In_790);
nor U1141 (N_1141,N_713,N_810);
nor U1142 (N_1142,N_155,N_992);
xnor U1143 (N_1143,In_650,N_986);
nor U1144 (N_1144,N_484,N_719);
xnor U1145 (N_1145,In_648,N_461);
and U1146 (N_1146,N_932,In_958);
and U1147 (N_1147,N_703,N_685);
xnor U1148 (N_1148,In_296,N_933);
nor U1149 (N_1149,N_835,In_733);
xor U1150 (N_1150,In_806,N_576);
or U1151 (N_1151,In_1221,N_688);
xnor U1152 (N_1152,In_1053,N_641);
nor U1153 (N_1153,N_397,N_978);
nor U1154 (N_1154,In_676,In_332);
and U1155 (N_1155,In_934,In_1499);
nand U1156 (N_1156,N_331,N_512);
xnor U1157 (N_1157,N_714,N_624);
nand U1158 (N_1158,N_808,N_218);
xor U1159 (N_1159,N_988,N_849);
and U1160 (N_1160,N_373,N_620);
nor U1161 (N_1161,N_865,N_62);
nand U1162 (N_1162,N_847,In_528);
nor U1163 (N_1163,N_846,In_951);
nand U1164 (N_1164,N_985,In_993);
nand U1165 (N_1165,N_907,N_889);
or U1166 (N_1166,N_830,N_794);
nand U1167 (N_1167,N_39,N_652);
or U1168 (N_1168,In_1239,N_936);
xor U1169 (N_1169,N_531,N_622);
nor U1170 (N_1170,N_894,N_836);
and U1171 (N_1171,N_890,In_1254);
nand U1172 (N_1172,N_917,N_882);
xor U1173 (N_1173,N_969,N_495);
nor U1174 (N_1174,N_510,In_469);
xor U1175 (N_1175,N_952,N_329);
nor U1176 (N_1176,N_838,In_1270);
or U1177 (N_1177,In_485,In_1451);
nand U1178 (N_1178,N_982,N_989);
xor U1179 (N_1179,N_956,N_843);
and U1180 (N_1180,In_392,N_859);
nand U1181 (N_1181,N_883,N_916);
xnor U1182 (N_1182,N_157,In_794);
xnor U1183 (N_1183,N_839,N_675);
xnor U1184 (N_1184,N_795,N_981);
and U1185 (N_1185,N_759,In_412);
xor U1186 (N_1186,N_909,N_475);
or U1187 (N_1187,N_446,N_997);
or U1188 (N_1188,N_250,N_309);
xor U1189 (N_1189,In_787,N_135);
nor U1190 (N_1190,N_733,N_162);
and U1191 (N_1191,N_920,N_205);
xor U1192 (N_1192,N_360,N_896);
xnor U1193 (N_1193,N_757,N_551);
nor U1194 (N_1194,N_613,N_930);
nand U1195 (N_1195,In_1157,N_738);
or U1196 (N_1196,N_681,N_72);
xor U1197 (N_1197,N_897,N_819);
nand U1198 (N_1198,N_943,N_880);
nor U1199 (N_1199,N_509,N_827);
and U1200 (N_1200,N_1021,N_1044);
or U1201 (N_1201,N_1053,In_1323);
and U1202 (N_1202,N_1048,N_934);
xor U1203 (N_1203,N_800,N_1187);
and U1204 (N_1204,N_1183,N_1022);
and U1205 (N_1205,N_828,N_1151);
or U1206 (N_1206,N_990,N_1118);
and U1207 (N_1207,N_1082,N_372);
nand U1208 (N_1208,N_1156,N_1077);
and U1209 (N_1209,N_951,N_931);
and U1210 (N_1210,N_1078,N_1199);
and U1211 (N_1211,N_1161,N_1164);
nor U1212 (N_1212,N_791,N_726);
nor U1213 (N_1213,N_1035,N_1085);
nor U1214 (N_1214,N_580,N_1195);
nor U1215 (N_1215,In_33,N_875);
nand U1216 (N_1216,N_1065,N_1080);
and U1217 (N_1217,N_957,N_848);
nor U1218 (N_1218,N_1052,N_237);
nand U1219 (N_1219,N_1130,N_1132);
nor U1220 (N_1220,N_779,N_1177);
nor U1221 (N_1221,N_1142,N_1124);
nor U1222 (N_1222,N_895,N_1117);
or U1223 (N_1223,N_980,N_1011);
nand U1224 (N_1224,N_21,N_961);
xnor U1225 (N_1225,N_1042,N_1169);
and U1226 (N_1226,N_841,N_1137);
xnor U1227 (N_1227,N_1185,N_1198);
xor U1228 (N_1228,N_1079,N_814);
xor U1229 (N_1229,N_1040,N_842);
nand U1230 (N_1230,N_1145,N_1134);
or U1231 (N_1231,In_369,N_1066);
nand U1232 (N_1232,N_472,N_1093);
and U1233 (N_1233,N_1112,In_282);
or U1234 (N_1234,N_1092,N_1148);
and U1235 (N_1235,N_1037,N_853);
nand U1236 (N_1236,In_358,N_1060);
xor U1237 (N_1237,In_975,N_628);
or U1238 (N_1238,N_1073,N_1155);
nand U1239 (N_1239,N_1004,N_1197);
nand U1240 (N_1240,N_1122,N_1146);
nand U1241 (N_1241,N_609,N_737);
and U1242 (N_1242,N_832,N_1016);
xor U1243 (N_1243,N_826,N_1116);
nand U1244 (N_1244,In_1119,N_1174);
nand U1245 (N_1245,N_1178,N_1125);
and U1246 (N_1246,In_108,N_1010);
nor U1247 (N_1247,N_740,N_1133);
nand U1248 (N_1248,N_1038,In_1090);
nand U1249 (N_1249,N_1171,N_912);
nor U1250 (N_1250,N_1182,N_1043);
nor U1251 (N_1251,N_1050,N_1184);
xnor U1252 (N_1252,N_1166,N_1167);
and U1253 (N_1253,N_1192,N_1190);
nor U1254 (N_1254,N_1086,N_1108);
nand U1255 (N_1255,N_1153,N_1104);
or U1256 (N_1256,N_1013,N_1031);
xnor U1257 (N_1257,N_1064,N_1149);
nand U1258 (N_1258,N_993,N_1058);
and U1259 (N_1259,N_1030,N_1111);
nand U1260 (N_1260,N_1039,N_1027);
and U1261 (N_1261,N_1121,N_873);
nor U1262 (N_1262,N_1015,N_1101);
and U1263 (N_1263,N_1025,N_1176);
or U1264 (N_1264,N_1006,N_1068);
xnor U1265 (N_1265,N_1000,N_1165);
nand U1266 (N_1266,N_983,In_239);
or U1267 (N_1267,N_1023,N_977);
and U1268 (N_1268,N_1163,N_885);
nand U1269 (N_1269,N_1075,N_924);
xnor U1270 (N_1270,N_415,N_1088);
or U1271 (N_1271,N_761,N_1126);
and U1272 (N_1272,N_1109,N_829);
or U1273 (N_1273,N_939,N_1012);
or U1274 (N_1274,N_592,N_1194);
nand U1275 (N_1275,N_1136,N_901);
nor U1276 (N_1276,N_1172,N_1099);
xor U1277 (N_1277,N_1114,N_1055);
nand U1278 (N_1278,N_1189,N_1150);
nand U1279 (N_1279,N_906,N_1017);
xor U1280 (N_1280,N_1107,N_1056);
or U1281 (N_1281,N_464,N_1138);
xnor U1282 (N_1282,N_715,N_457);
and U1283 (N_1283,N_1123,N_1041);
and U1284 (N_1284,N_1063,N_812);
nand U1285 (N_1285,N_742,N_564);
nor U1286 (N_1286,N_1036,N_118);
nor U1287 (N_1287,N_1143,In_1065);
xnor U1288 (N_1288,N_1019,N_1057);
and U1289 (N_1289,In_139,N_1179);
and U1290 (N_1290,N_999,N_301);
nor U1291 (N_1291,N_1162,N_1110);
nor U1292 (N_1292,N_1129,N_1152);
nand U1293 (N_1293,N_1105,N_1157);
xnor U1294 (N_1294,N_1061,N_1051);
or U1295 (N_1295,In_1003,N_1106);
nor U1296 (N_1296,N_1083,N_1009);
xor U1297 (N_1297,N_1103,In_1005);
nor U1298 (N_1298,N_1090,In_455);
xor U1299 (N_1299,N_867,In_530);
nor U1300 (N_1300,N_1096,N_1084);
xnor U1301 (N_1301,In_883,N_1094);
nor U1302 (N_1302,In_796,N_1029);
xor U1303 (N_1303,N_1071,N_1074);
xor U1304 (N_1304,N_1026,N_1144);
or U1305 (N_1305,N_1139,N_751);
and U1306 (N_1306,N_697,N_222);
nor U1307 (N_1307,N_1135,N_869);
or U1308 (N_1308,In_857,N_1024);
nand U1309 (N_1309,N_1014,N_1119);
and U1310 (N_1310,N_655,N_1140);
nand U1311 (N_1311,N_1070,N_1147);
or U1312 (N_1312,N_635,N_854);
nand U1313 (N_1313,N_1095,In_0);
xor U1314 (N_1314,N_734,N_1181);
nor U1315 (N_1315,N_1100,N_1007);
nor U1316 (N_1316,N_852,N_1072);
and U1317 (N_1317,N_1127,In_1192);
and U1318 (N_1318,N_1003,N_1067);
and U1319 (N_1319,N_1097,N_1032);
or U1320 (N_1320,N_1089,N_1170);
nor U1321 (N_1321,N_892,N_1001);
and U1322 (N_1322,In_897,N_921);
xor U1323 (N_1323,N_710,N_1168);
or U1324 (N_1324,N_1175,N_953);
nand U1325 (N_1325,N_1128,N_1028);
and U1326 (N_1326,N_1091,N_1069);
xor U1327 (N_1327,N_1131,N_478);
or U1328 (N_1328,N_1193,N_786);
nor U1329 (N_1329,N_979,N_1046);
xnor U1330 (N_1330,N_1160,N_1158);
and U1331 (N_1331,In_162,N_406);
and U1332 (N_1332,N_1062,N_1034);
or U1333 (N_1333,N_1018,In_19);
xnor U1334 (N_1334,N_1033,N_1081);
xor U1335 (N_1335,N_1076,N_1115);
and U1336 (N_1336,N_1054,N_1113);
and U1337 (N_1337,N_452,N_1154);
and U1338 (N_1338,N_1159,N_1186);
xor U1339 (N_1339,N_1047,N_996);
and U1340 (N_1340,N_1045,N_614);
or U1341 (N_1341,N_1196,N_1059);
xor U1342 (N_1342,N_1005,In_176);
nor U1343 (N_1343,N_1180,N_1049);
and U1344 (N_1344,N_1008,N_1120);
nor U1345 (N_1345,N_1087,N_1002);
nor U1346 (N_1346,N_1102,In_1430);
xor U1347 (N_1347,N_1098,N_1141);
nor U1348 (N_1348,N_1191,N_1173);
nor U1349 (N_1349,N_1020,N_1188);
xor U1350 (N_1350,N_1000,N_1053);
nand U1351 (N_1351,N_1080,N_1143);
or U1352 (N_1352,N_1081,N_1121);
nand U1353 (N_1353,N_222,N_592);
nor U1354 (N_1354,N_1085,N_1003);
nand U1355 (N_1355,N_848,N_1009);
nor U1356 (N_1356,N_1014,N_1063);
and U1357 (N_1357,N_1015,N_1088);
and U1358 (N_1358,N_1026,N_1107);
or U1359 (N_1359,N_1047,N_828);
nor U1360 (N_1360,N_1193,N_1035);
xor U1361 (N_1361,N_222,N_737);
or U1362 (N_1362,N_1054,N_1023);
and U1363 (N_1363,N_1166,N_1143);
nor U1364 (N_1364,N_1113,N_1060);
nor U1365 (N_1365,N_472,N_1048);
and U1366 (N_1366,N_1028,N_875);
or U1367 (N_1367,N_1163,N_875);
or U1368 (N_1368,N_841,N_869);
or U1369 (N_1369,In_857,N_1042);
xnor U1370 (N_1370,N_1137,N_1143);
nor U1371 (N_1371,In_975,N_1111);
nand U1372 (N_1372,In_176,N_1157);
nor U1373 (N_1373,N_1163,N_980);
nor U1374 (N_1374,N_999,N_1163);
and U1375 (N_1375,N_1080,N_1079);
or U1376 (N_1376,N_592,N_1061);
xnor U1377 (N_1377,N_237,N_812);
and U1378 (N_1378,In_796,N_609);
xnor U1379 (N_1379,N_1125,N_1195);
and U1380 (N_1380,N_1017,N_742);
xor U1381 (N_1381,In_108,N_1046);
and U1382 (N_1382,N_301,N_1167);
nor U1383 (N_1383,N_1156,N_464);
xor U1384 (N_1384,N_609,N_901);
xor U1385 (N_1385,N_1086,N_1078);
or U1386 (N_1386,N_1191,N_1119);
or U1387 (N_1387,N_828,In_139);
nand U1388 (N_1388,N_1197,N_1126);
nor U1389 (N_1389,N_1160,N_1153);
nand U1390 (N_1390,In_1065,N_1028);
nor U1391 (N_1391,N_1174,N_1149);
nor U1392 (N_1392,In_857,N_1155);
and U1393 (N_1393,N_1007,N_1134);
xnor U1394 (N_1394,In_530,N_1088);
or U1395 (N_1395,N_1089,N_1179);
or U1396 (N_1396,In_369,N_1063);
or U1397 (N_1397,N_1193,N_1002);
nor U1398 (N_1398,N_1188,N_1084);
nor U1399 (N_1399,N_912,N_1026);
or U1400 (N_1400,N_1310,N_1366);
or U1401 (N_1401,N_1234,N_1380);
or U1402 (N_1402,N_1384,N_1215);
or U1403 (N_1403,N_1262,N_1323);
xor U1404 (N_1404,N_1396,N_1390);
and U1405 (N_1405,N_1238,N_1256);
nor U1406 (N_1406,N_1317,N_1359);
and U1407 (N_1407,N_1301,N_1247);
nand U1408 (N_1408,N_1309,N_1205);
xor U1409 (N_1409,N_1331,N_1240);
and U1410 (N_1410,N_1299,N_1217);
nor U1411 (N_1411,N_1338,N_1228);
or U1412 (N_1412,N_1298,N_1268);
or U1413 (N_1413,N_1272,N_1330);
and U1414 (N_1414,N_1393,N_1258);
xnor U1415 (N_1415,N_1216,N_1336);
xor U1416 (N_1416,N_1208,N_1209);
xor U1417 (N_1417,N_1388,N_1255);
or U1418 (N_1418,N_1369,N_1252);
nor U1419 (N_1419,N_1232,N_1337);
and U1420 (N_1420,N_1312,N_1230);
xnor U1421 (N_1421,N_1320,N_1253);
xnor U1422 (N_1422,N_1324,N_1377);
nand U1423 (N_1423,N_1294,N_1306);
nand U1424 (N_1424,N_1218,N_1318);
xor U1425 (N_1425,N_1353,N_1308);
nand U1426 (N_1426,N_1328,N_1354);
nand U1427 (N_1427,N_1334,N_1212);
or U1428 (N_1428,N_1361,N_1376);
xnor U1429 (N_1429,N_1292,N_1235);
and U1430 (N_1430,N_1311,N_1300);
and U1431 (N_1431,N_1259,N_1383);
nand U1432 (N_1432,N_1261,N_1305);
or U1433 (N_1433,N_1213,N_1332);
and U1434 (N_1434,N_1281,N_1207);
or U1435 (N_1435,N_1341,N_1274);
or U1436 (N_1436,N_1316,N_1263);
xnor U1437 (N_1437,N_1368,N_1371);
and U1438 (N_1438,N_1276,N_1279);
or U1439 (N_1439,N_1219,N_1282);
nand U1440 (N_1440,N_1201,N_1389);
and U1441 (N_1441,N_1398,N_1271);
xnor U1442 (N_1442,N_1333,N_1357);
nand U1443 (N_1443,N_1254,N_1363);
or U1444 (N_1444,N_1347,N_1378);
xnor U1445 (N_1445,N_1348,N_1260);
and U1446 (N_1446,N_1246,N_1343);
xnor U1447 (N_1447,N_1329,N_1245);
xor U1448 (N_1448,N_1239,N_1285);
nor U1449 (N_1449,N_1322,N_1267);
xnor U1450 (N_1450,N_1237,N_1206);
and U1451 (N_1451,N_1278,N_1373);
and U1452 (N_1452,N_1381,N_1362);
nand U1453 (N_1453,N_1236,N_1257);
xnor U1454 (N_1454,N_1335,N_1284);
xnor U1455 (N_1455,N_1248,N_1287);
nor U1456 (N_1456,N_1210,N_1286);
and U1457 (N_1457,N_1295,N_1293);
nand U1458 (N_1458,N_1244,N_1315);
nand U1459 (N_1459,N_1387,N_1220);
and U1460 (N_1460,N_1374,N_1342);
nand U1461 (N_1461,N_1200,N_1303);
nand U1462 (N_1462,N_1350,N_1379);
nor U1463 (N_1463,N_1325,N_1313);
nand U1464 (N_1464,N_1395,N_1229);
nor U1465 (N_1465,N_1399,N_1211);
nor U1466 (N_1466,N_1202,N_1314);
nand U1467 (N_1467,N_1307,N_1352);
nand U1468 (N_1468,N_1288,N_1227);
or U1469 (N_1469,N_1249,N_1233);
xnor U1470 (N_1470,N_1264,N_1203);
nand U1471 (N_1471,N_1283,N_1226);
or U1472 (N_1472,N_1280,N_1340);
nor U1473 (N_1473,N_1364,N_1297);
and U1474 (N_1474,N_1346,N_1321);
and U1475 (N_1475,N_1385,N_1351);
xor U1476 (N_1476,N_1349,N_1367);
and U1477 (N_1477,N_1214,N_1221);
nor U1478 (N_1478,N_1275,N_1222);
and U1479 (N_1479,N_1345,N_1370);
or U1480 (N_1480,N_1225,N_1223);
xnor U1481 (N_1481,N_1339,N_1392);
xor U1482 (N_1482,N_1243,N_1358);
and U1483 (N_1483,N_1242,N_1386);
nor U1484 (N_1484,N_1290,N_1302);
nand U1485 (N_1485,N_1224,N_1273);
or U1486 (N_1486,N_1391,N_1270);
nor U1487 (N_1487,N_1204,N_1360);
nor U1488 (N_1488,N_1365,N_1356);
and U1489 (N_1489,N_1326,N_1355);
xor U1490 (N_1490,N_1327,N_1382);
nand U1491 (N_1491,N_1251,N_1277);
nand U1492 (N_1492,N_1289,N_1372);
and U1493 (N_1493,N_1394,N_1250);
or U1494 (N_1494,N_1319,N_1296);
or U1495 (N_1495,N_1397,N_1375);
nor U1496 (N_1496,N_1231,N_1269);
xnor U1497 (N_1497,N_1291,N_1241);
and U1498 (N_1498,N_1265,N_1304);
or U1499 (N_1499,N_1266,N_1344);
nor U1500 (N_1500,N_1242,N_1375);
nor U1501 (N_1501,N_1349,N_1233);
nand U1502 (N_1502,N_1351,N_1243);
or U1503 (N_1503,N_1346,N_1327);
xor U1504 (N_1504,N_1390,N_1349);
and U1505 (N_1505,N_1298,N_1379);
nand U1506 (N_1506,N_1349,N_1302);
xor U1507 (N_1507,N_1263,N_1246);
nand U1508 (N_1508,N_1305,N_1278);
and U1509 (N_1509,N_1243,N_1274);
and U1510 (N_1510,N_1241,N_1337);
xor U1511 (N_1511,N_1271,N_1228);
xor U1512 (N_1512,N_1263,N_1243);
and U1513 (N_1513,N_1207,N_1369);
and U1514 (N_1514,N_1350,N_1377);
or U1515 (N_1515,N_1369,N_1312);
nand U1516 (N_1516,N_1200,N_1376);
xor U1517 (N_1517,N_1298,N_1284);
nand U1518 (N_1518,N_1245,N_1397);
or U1519 (N_1519,N_1309,N_1203);
nand U1520 (N_1520,N_1333,N_1201);
nand U1521 (N_1521,N_1227,N_1363);
and U1522 (N_1522,N_1360,N_1248);
and U1523 (N_1523,N_1282,N_1261);
and U1524 (N_1524,N_1260,N_1362);
xor U1525 (N_1525,N_1270,N_1300);
xor U1526 (N_1526,N_1299,N_1225);
or U1527 (N_1527,N_1237,N_1235);
xnor U1528 (N_1528,N_1238,N_1224);
nand U1529 (N_1529,N_1264,N_1295);
or U1530 (N_1530,N_1319,N_1337);
and U1531 (N_1531,N_1322,N_1268);
xnor U1532 (N_1532,N_1213,N_1281);
nor U1533 (N_1533,N_1366,N_1232);
and U1534 (N_1534,N_1220,N_1371);
xnor U1535 (N_1535,N_1377,N_1273);
xor U1536 (N_1536,N_1247,N_1344);
xnor U1537 (N_1537,N_1327,N_1386);
nand U1538 (N_1538,N_1256,N_1272);
nand U1539 (N_1539,N_1363,N_1283);
nand U1540 (N_1540,N_1238,N_1334);
or U1541 (N_1541,N_1324,N_1336);
xnor U1542 (N_1542,N_1224,N_1222);
and U1543 (N_1543,N_1335,N_1383);
nand U1544 (N_1544,N_1337,N_1370);
or U1545 (N_1545,N_1218,N_1351);
or U1546 (N_1546,N_1298,N_1309);
nor U1547 (N_1547,N_1251,N_1311);
nand U1548 (N_1548,N_1398,N_1290);
nand U1549 (N_1549,N_1395,N_1249);
and U1550 (N_1550,N_1377,N_1373);
nor U1551 (N_1551,N_1247,N_1232);
nand U1552 (N_1552,N_1355,N_1200);
and U1553 (N_1553,N_1288,N_1258);
xor U1554 (N_1554,N_1336,N_1355);
and U1555 (N_1555,N_1293,N_1335);
nor U1556 (N_1556,N_1266,N_1230);
and U1557 (N_1557,N_1384,N_1216);
nor U1558 (N_1558,N_1220,N_1393);
nor U1559 (N_1559,N_1343,N_1214);
and U1560 (N_1560,N_1218,N_1375);
and U1561 (N_1561,N_1381,N_1351);
or U1562 (N_1562,N_1307,N_1302);
nor U1563 (N_1563,N_1234,N_1302);
nand U1564 (N_1564,N_1222,N_1241);
nor U1565 (N_1565,N_1352,N_1300);
nand U1566 (N_1566,N_1297,N_1321);
nand U1567 (N_1567,N_1330,N_1354);
or U1568 (N_1568,N_1323,N_1257);
and U1569 (N_1569,N_1276,N_1204);
xnor U1570 (N_1570,N_1210,N_1345);
and U1571 (N_1571,N_1330,N_1276);
nand U1572 (N_1572,N_1378,N_1299);
and U1573 (N_1573,N_1330,N_1377);
nor U1574 (N_1574,N_1329,N_1208);
nand U1575 (N_1575,N_1239,N_1236);
and U1576 (N_1576,N_1355,N_1389);
nand U1577 (N_1577,N_1265,N_1365);
and U1578 (N_1578,N_1330,N_1327);
or U1579 (N_1579,N_1227,N_1297);
nand U1580 (N_1580,N_1231,N_1356);
and U1581 (N_1581,N_1306,N_1384);
nand U1582 (N_1582,N_1353,N_1348);
xor U1583 (N_1583,N_1276,N_1337);
nand U1584 (N_1584,N_1211,N_1229);
and U1585 (N_1585,N_1280,N_1282);
xor U1586 (N_1586,N_1328,N_1378);
nor U1587 (N_1587,N_1334,N_1265);
or U1588 (N_1588,N_1308,N_1251);
nor U1589 (N_1589,N_1376,N_1329);
nand U1590 (N_1590,N_1230,N_1290);
nor U1591 (N_1591,N_1377,N_1227);
xnor U1592 (N_1592,N_1391,N_1343);
nor U1593 (N_1593,N_1339,N_1219);
and U1594 (N_1594,N_1381,N_1397);
and U1595 (N_1595,N_1332,N_1253);
nand U1596 (N_1596,N_1228,N_1353);
nor U1597 (N_1597,N_1257,N_1347);
and U1598 (N_1598,N_1226,N_1239);
nor U1599 (N_1599,N_1390,N_1380);
or U1600 (N_1600,N_1507,N_1576);
or U1601 (N_1601,N_1452,N_1491);
xor U1602 (N_1602,N_1439,N_1537);
xnor U1603 (N_1603,N_1432,N_1423);
nor U1604 (N_1604,N_1467,N_1519);
nor U1605 (N_1605,N_1583,N_1543);
and U1606 (N_1606,N_1506,N_1524);
xnor U1607 (N_1607,N_1413,N_1482);
xor U1608 (N_1608,N_1502,N_1459);
and U1609 (N_1609,N_1446,N_1525);
or U1610 (N_1610,N_1431,N_1566);
or U1611 (N_1611,N_1409,N_1435);
nor U1612 (N_1612,N_1577,N_1593);
xnor U1613 (N_1613,N_1533,N_1441);
nand U1614 (N_1614,N_1487,N_1585);
and U1615 (N_1615,N_1540,N_1480);
or U1616 (N_1616,N_1425,N_1493);
or U1617 (N_1617,N_1461,N_1450);
nor U1618 (N_1618,N_1477,N_1573);
nand U1619 (N_1619,N_1400,N_1410);
or U1620 (N_1620,N_1565,N_1417);
nor U1621 (N_1621,N_1570,N_1440);
or U1622 (N_1622,N_1584,N_1481);
xor U1623 (N_1623,N_1466,N_1515);
nand U1624 (N_1624,N_1445,N_1545);
and U1625 (N_1625,N_1529,N_1516);
or U1626 (N_1626,N_1501,N_1534);
and U1627 (N_1627,N_1427,N_1572);
and U1628 (N_1628,N_1530,N_1532);
xor U1629 (N_1629,N_1541,N_1568);
and U1630 (N_1630,N_1415,N_1483);
nor U1631 (N_1631,N_1528,N_1464);
xor U1632 (N_1632,N_1468,N_1581);
nand U1633 (N_1633,N_1489,N_1598);
nand U1634 (N_1634,N_1421,N_1479);
and U1635 (N_1635,N_1455,N_1562);
or U1636 (N_1636,N_1492,N_1426);
xnor U1637 (N_1637,N_1544,N_1419);
nand U1638 (N_1638,N_1474,N_1592);
nand U1639 (N_1639,N_1438,N_1469);
or U1640 (N_1640,N_1494,N_1485);
nor U1641 (N_1641,N_1520,N_1526);
nand U1642 (N_1642,N_1434,N_1463);
nor U1643 (N_1643,N_1542,N_1538);
nand U1644 (N_1644,N_1476,N_1546);
nand U1645 (N_1645,N_1551,N_1497);
nor U1646 (N_1646,N_1510,N_1559);
xnor U1647 (N_1647,N_1402,N_1509);
xor U1648 (N_1648,N_1561,N_1498);
xor U1649 (N_1649,N_1499,N_1536);
xnor U1650 (N_1650,N_1444,N_1560);
and U1651 (N_1651,N_1454,N_1405);
xnor U1652 (N_1652,N_1420,N_1406);
nand U1653 (N_1653,N_1448,N_1418);
and U1654 (N_1654,N_1578,N_1594);
and U1655 (N_1655,N_1517,N_1587);
and U1656 (N_1656,N_1555,N_1599);
and U1657 (N_1657,N_1401,N_1567);
nor U1658 (N_1658,N_1595,N_1512);
nand U1659 (N_1659,N_1447,N_1552);
nor U1660 (N_1660,N_1486,N_1451);
or U1661 (N_1661,N_1586,N_1407);
or U1662 (N_1662,N_1574,N_1470);
nor U1663 (N_1663,N_1548,N_1535);
and U1664 (N_1664,N_1496,N_1473);
xor U1665 (N_1665,N_1465,N_1557);
nor U1666 (N_1666,N_1508,N_1442);
nand U1667 (N_1667,N_1422,N_1575);
xor U1668 (N_1668,N_1579,N_1504);
nor U1669 (N_1669,N_1456,N_1511);
nor U1670 (N_1670,N_1437,N_1443);
or U1671 (N_1671,N_1564,N_1495);
and U1672 (N_1672,N_1549,N_1582);
and U1673 (N_1673,N_1554,N_1490);
and U1674 (N_1674,N_1488,N_1484);
nor U1675 (N_1675,N_1505,N_1547);
or U1676 (N_1676,N_1460,N_1580);
and U1677 (N_1677,N_1556,N_1500);
nand U1678 (N_1678,N_1563,N_1471);
xor U1679 (N_1679,N_1462,N_1588);
nor U1680 (N_1680,N_1513,N_1408);
xor U1681 (N_1681,N_1458,N_1590);
or U1682 (N_1682,N_1414,N_1430);
or U1683 (N_1683,N_1475,N_1472);
xor U1684 (N_1684,N_1416,N_1596);
and U1685 (N_1685,N_1433,N_1527);
xnor U1686 (N_1686,N_1569,N_1436);
nor U1687 (N_1687,N_1412,N_1429);
nor U1688 (N_1688,N_1531,N_1597);
and U1689 (N_1689,N_1522,N_1550);
or U1690 (N_1690,N_1449,N_1558);
nand U1691 (N_1691,N_1539,N_1403);
xor U1692 (N_1692,N_1514,N_1521);
nor U1693 (N_1693,N_1424,N_1503);
nor U1694 (N_1694,N_1591,N_1589);
and U1695 (N_1695,N_1411,N_1553);
and U1696 (N_1696,N_1457,N_1404);
nor U1697 (N_1697,N_1428,N_1478);
and U1698 (N_1698,N_1453,N_1571);
and U1699 (N_1699,N_1523,N_1518);
and U1700 (N_1700,N_1491,N_1483);
and U1701 (N_1701,N_1475,N_1575);
and U1702 (N_1702,N_1423,N_1411);
or U1703 (N_1703,N_1418,N_1423);
nor U1704 (N_1704,N_1592,N_1463);
xor U1705 (N_1705,N_1585,N_1560);
xnor U1706 (N_1706,N_1525,N_1406);
nand U1707 (N_1707,N_1405,N_1446);
and U1708 (N_1708,N_1413,N_1478);
xor U1709 (N_1709,N_1461,N_1473);
xnor U1710 (N_1710,N_1400,N_1498);
nor U1711 (N_1711,N_1547,N_1574);
nand U1712 (N_1712,N_1474,N_1403);
nand U1713 (N_1713,N_1469,N_1516);
xnor U1714 (N_1714,N_1470,N_1532);
xnor U1715 (N_1715,N_1596,N_1547);
nand U1716 (N_1716,N_1577,N_1470);
or U1717 (N_1717,N_1586,N_1458);
xor U1718 (N_1718,N_1497,N_1428);
xnor U1719 (N_1719,N_1441,N_1588);
and U1720 (N_1720,N_1517,N_1489);
and U1721 (N_1721,N_1478,N_1495);
or U1722 (N_1722,N_1419,N_1429);
xnor U1723 (N_1723,N_1432,N_1556);
or U1724 (N_1724,N_1428,N_1503);
and U1725 (N_1725,N_1461,N_1547);
or U1726 (N_1726,N_1514,N_1530);
xor U1727 (N_1727,N_1516,N_1458);
xnor U1728 (N_1728,N_1568,N_1552);
or U1729 (N_1729,N_1477,N_1560);
nor U1730 (N_1730,N_1510,N_1532);
or U1731 (N_1731,N_1543,N_1491);
xor U1732 (N_1732,N_1450,N_1553);
nor U1733 (N_1733,N_1506,N_1596);
and U1734 (N_1734,N_1476,N_1506);
nand U1735 (N_1735,N_1453,N_1438);
xor U1736 (N_1736,N_1573,N_1543);
or U1737 (N_1737,N_1559,N_1580);
nand U1738 (N_1738,N_1442,N_1467);
nand U1739 (N_1739,N_1495,N_1533);
and U1740 (N_1740,N_1482,N_1406);
nor U1741 (N_1741,N_1561,N_1523);
xnor U1742 (N_1742,N_1451,N_1403);
or U1743 (N_1743,N_1518,N_1509);
or U1744 (N_1744,N_1564,N_1470);
nand U1745 (N_1745,N_1485,N_1564);
or U1746 (N_1746,N_1495,N_1567);
or U1747 (N_1747,N_1542,N_1460);
and U1748 (N_1748,N_1595,N_1410);
or U1749 (N_1749,N_1460,N_1427);
and U1750 (N_1750,N_1548,N_1511);
nor U1751 (N_1751,N_1475,N_1578);
or U1752 (N_1752,N_1401,N_1534);
nand U1753 (N_1753,N_1505,N_1412);
nand U1754 (N_1754,N_1486,N_1423);
xor U1755 (N_1755,N_1420,N_1411);
nor U1756 (N_1756,N_1419,N_1449);
and U1757 (N_1757,N_1442,N_1575);
xnor U1758 (N_1758,N_1567,N_1503);
xor U1759 (N_1759,N_1462,N_1449);
nor U1760 (N_1760,N_1499,N_1449);
and U1761 (N_1761,N_1510,N_1584);
xnor U1762 (N_1762,N_1518,N_1494);
xnor U1763 (N_1763,N_1427,N_1529);
or U1764 (N_1764,N_1558,N_1454);
nand U1765 (N_1765,N_1445,N_1522);
nor U1766 (N_1766,N_1446,N_1514);
nand U1767 (N_1767,N_1453,N_1446);
nand U1768 (N_1768,N_1400,N_1401);
and U1769 (N_1769,N_1556,N_1577);
xnor U1770 (N_1770,N_1439,N_1512);
nor U1771 (N_1771,N_1501,N_1590);
nand U1772 (N_1772,N_1596,N_1473);
nor U1773 (N_1773,N_1522,N_1569);
nand U1774 (N_1774,N_1496,N_1577);
nor U1775 (N_1775,N_1510,N_1542);
nand U1776 (N_1776,N_1524,N_1530);
and U1777 (N_1777,N_1548,N_1517);
nor U1778 (N_1778,N_1421,N_1419);
nor U1779 (N_1779,N_1468,N_1433);
or U1780 (N_1780,N_1589,N_1428);
nor U1781 (N_1781,N_1525,N_1443);
nor U1782 (N_1782,N_1579,N_1490);
or U1783 (N_1783,N_1421,N_1553);
nand U1784 (N_1784,N_1463,N_1473);
nor U1785 (N_1785,N_1509,N_1432);
xnor U1786 (N_1786,N_1488,N_1575);
or U1787 (N_1787,N_1504,N_1527);
and U1788 (N_1788,N_1581,N_1500);
xnor U1789 (N_1789,N_1532,N_1486);
nand U1790 (N_1790,N_1464,N_1552);
and U1791 (N_1791,N_1527,N_1547);
nand U1792 (N_1792,N_1486,N_1419);
nor U1793 (N_1793,N_1563,N_1456);
and U1794 (N_1794,N_1593,N_1440);
xor U1795 (N_1795,N_1490,N_1546);
xnor U1796 (N_1796,N_1534,N_1476);
nor U1797 (N_1797,N_1582,N_1573);
xnor U1798 (N_1798,N_1595,N_1456);
xnor U1799 (N_1799,N_1424,N_1401);
nand U1800 (N_1800,N_1730,N_1693);
and U1801 (N_1801,N_1779,N_1739);
or U1802 (N_1802,N_1774,N_1778);
nor U1803 (N_1803,N_1625,N_1675);
xnor U1804 (N_1804,N_1707,N_1703);
xnor U1805 (N_1805,N_1736,N_1669);
or U1806 (N_1806,N_1666,N_1757);
nor U1807 (N_1807,N_1668,N_1712);
nor U1808 (N_1808,N_1609,N_1754);
or U1809 (N_1809,N_1798,N_1758);
or U1810 (N_1810,N_1610,N_1679);
nand U1811 (N_1811,N_1607,N_1697);
xnor U1812 (N_1812,N_1631,N_1765);
xor U1813 (N_1813,N_1637,N_1680);
nor U1814 (N_1814,N_1717,N_1752);
and U1815 (N_1815,N_1655,N_1664);
nor U1816 (N_1816,N_1600,N_1729);
nor U1817 (N_1817,N_1677,N_1797);
nor U1818 (N_1818,N_1740,N_1769);
nand U1819 (N_1819,N_1792,N_1702);
nor U1820 (N_1820,N_1748,N_1721);
xnor U1821 (N_1821,N_1785,N_1737);
and U1822 (N_1822,N_1762,N_1684);
xor U1823 (N_1823,N_1788,N_1743);
nand U1824 (N_1824,N_1647,N_1648);
nand U1825 (N_1825,N_1636,N_1756);
and U1826 (N_1826,N_1790,N_1761);
nand U1827 (N_1827,N_1651,N_1783);
xor U1828 (N_1828,N_1782,N_1628);
or U1829 (N_1829,N_1724,N_1727);
and U1830 (N_1830,N_1733,N_1700);
and U1831 (N_1831,N_1608,N_1726);
nor U1832 (N_1832,N_1641,N_1686);
xor U1833 (N_1833,N_1674,N_1692);
xnor U1834 (N_1834,N_1618,N_1704);
xor U1835 (N_1835,N_1742,N_1644);
nor U1836 (N_1836,N_1665,N_1716);
nor U1837 (N_1837,N_1683,N_1620);
and U1838 (N_1838,N_1606,N_1614);
and U1839 (N_1839,N_1626,N_1698);
or U1840 (N_1840,N_1670,N_1685);
or U1841 (N_1841,N_1642,N_1766);
and U1842 (N_1842,N_1638,N_1708);
xnor U1843 (N_1843,N_1734,N_1786);
nor U1844 (N_1844,N_1658,N_1767);
and U1845 (N_1845,N_1656,N_1661);
nand U1846 (N_1846,N_1745,N_1643);
nor U1847 (N_1847,N_1612,N_1710);
nor U1848 (N_1848,N_1659,N_1645);
nand U1849 (N_1849,N_1719,N_1671);
nor U1850 (N_1850,N_1689,N_1738);
xor U1851 (N_1851,N_1723,N_1731);
nor U1852 (N_1852,N_1694,N_1696);
xor U1853 (N_1853,N_1649,N_1755);
nand U1854 (N_1854,N_1718,N_1725);
nand U1855 (N_1855,N_1624,N_1793);
and U1856 (N_1856,N_1772,N_1760);
nor U1857 (N_1857,N_1722,N_1690);
nor U1858 (N_1858,N_1640,N_1632);
or U1859 (N_1859,N_1751,N_1775);
or U1860 (N_1860,N_1713,N_1720);
nor U1861 (N_1861,N_1633,N_1747);
nand U1862 (N_1862,N_1771,N_1768);
nand U1863 (N_1863,N_1667,N_1678);
and U1864 (N_1864,N_1750,N_1789);
and U1865 (N_1865,N_1687,N_1654);
and U1866 (N_1866,N_1603,N_1619);
and U1867 (N_1867,N_1617,N_1657);
xnor U1868 (N_1868,N_1630,N_1749);
or U1869 (N_1869,N_1627,N_1759);
nor U1870 (N_1870,N_1602,N_1634);
xor U1871 (N_1871,N_1673,N_1650);
nand U1872 (N_1872,N_1672,N_1646);
and U1873 (N_1873,N_1714,N_1796);
or U1874 (N_1874,N_1635,N_1770);
nand U1875 (N_1875,N_1639,N_1611);
nand U1876 (N_1876,N_1781,N_1753);
xor U1877 (N_1877,N_1791,N_1653);
nand U1878 (N_1878,N_1728,N_1629);
xor U1879 (N_1879,N_1746,N_1621);
nor U1880 (N_1880,N_1763,N_1780);
nand U1881 (N_1881,N_1784,N_1662);
and U1882 (N_1882,N_1706,N_1613);
xor U1883 (N_1883,N_1735,N_1616);
nor U1884 (N_1884,N_1691,N_1695);
xnor U1885 (N_1885,N_1682,N_1663);
nor U1886 (N_1886,N_1744,N_1799);
or U1887 (N_1887,N_1660,N_1676);
nor U1888 (N_1888,N_1652,N_1711);
and U1889 (N_1889,N_1732,N_1705);
or U1890 (N_1890,N_1764,N_1715);
or U1891 (N_1891,N_1699,N_1688);
or U1892 (N_1892,N_1622,N_1794);
nand U1893 (N_1893,N_1604,N_1773);
nand U1894 (N_1894,N_1709,N_1623);
xnor U1895 (N_1895,N_1681,N_1776);
nor U1896 (N_1896,N_1601,N_1615);
nand U1897 (N_1897,N_1787,N_1795);
and U1898 (N_1898,N_1777,N_1741);
nand U1899 (N_1899,N_1605,N_1701);
nor U1900 (N_1900,N_1740,N_1656);
nand U1901 (N_1901,N_1622,N_1641);
nor U1902 (N_1902,N_1692,N_1778);
nand U1903 (N_1903,N_1778,N_1605);
or U1904 (N_1904,N_1757,N_1793);
nor U1905 (N_1905,N_1769,N_1739);
or U1906 (N_1906,N_1779,N_1680);
or U1907 (N_1907,N_1631,N_1794);
xnor U1908 (N_1908,N_1796,N_1605);
or U1909 (N_1909,N_1617,N_1772);
and U1910 (N_1910,N_1747,N_1763);
and U1911 (N_1911,N_1752,N_1799);
xnor U1912 (N_1912,N_1664,N_1795);
nand U1913 (N_1913,N_1646,N_1643);
or U1914 (N_1914,N_1752,N_1659);
nor U1915 (N_1915,N_1710,N_1732);
nand U1916 (N_1916,N_1719,N_1781);
nor U1917 (N_1917,N_1773,N_1734);
xnor U1918 (N_1918,N_1785,N_1696);
nor U1919 (N_1919,N_1788,N_1618);
xor U1920 (N_1920,N_1714,N_1694);
xor U1921 (N_1921,N_1604,N_1643);
xnor U1922 (N_1922,N_1715,N_1794);
and U1923 (N_1923,N_1697,N_1631);
xnor U1924 (N_1924,N_1733,N_1787);
nand U1925 (N_1925,N_1683,N_1626);
or U1926 (N_1926,N_1713,N_1784);
xnor U1927 (N_1927,N_1662,N_1689);
xnor U1928 (N_1928,N_1635,N_1765);
xor U1929 (N_1929,N_1722,N_1776);
nand U1930 (N_1930,N_1765,N_1664);
or U1931 (N_1931,N_1727,N_1768);
nor U1932 (N_1932,N_1705,N_1703);
nor U1933 (N_1933,N_1647,N_1691);
nor U1934 (N_1934,N_1725,N_1760);
or U1935 (N_1935,N_1757,N_1626);
nor U1936 (N_1936,N_1768,N_1619);
nor U1937 (N_1937,N_1728,N_1747);
nor U1938 (N_1938,N_1615,N_1633);
xor U1939 (N_1939,N_1672,N_1794);
or U1940 (N_1940,N_1784,N_1682);
nand U1941 (N_1941,N_1609,N_1735);
nand U1942 (N_1942,N_1735,N_1784);
xor U1943 (N_1943,N_1705,N_1683);
nor U1944 (N_1944,N_1797,N_1657);
xor U1945 (N_1945,N_1709,N_1733);
nor U1946 (N_1946,N_1758,N_1639);
nor U1947 (N_1947,N_1614,N_1722);
nor U1948 (N_1948,N_1725,N_1798);
nand U1949 (N_1949,N_1666,N_1761);
nor U1950 (N_1950,N_1764,N_1672);
or U1951 (N_1951,N_1737,N_1701);
and U1952 (N_1952,N_1654,N_1788);
xnor U1953 (N_1953,N_1663,N_1622);
nand U1954 (N_1954,N_1705,N_1730);
or U1955 (N_1955,N_1664,N_1707);
nor U1956 (N_1956,N_1710,N_1665);
or U1957 (N_1957,N_1773,N_1709);
nor U1958 (N_1958,N_1652,N_1655);
or U1959 (N_1959,N_1736,N_1614);
and U1960 (N_1960,N_1623,N_1760);
nand U1961 (N_1961,N_1791,N_1613);
nor U1962 (N_1962,N_1691,N_1671);
nand U1963 (N_1963,N_1663,N_1609);
nand U1964 (N_1964,N_1607,N_1653);
xnor U1965 (N_1965,N_1611,N_1678);
nand U1966 (N_1966,N_1634,N_1640);
xor U1967 (N_1967,N_1789,N_1793);
xnor U1968 (N_1968,N_1787,N_1633);
xnor U1969 (N_1969,N_1693,N_1657);
nand U1970 (N_1970,N_1709,N_1649);
nor U1971 (N_1971,N_1742,N_1627);
nor U1972 (N_1972,N_1657,N_1741);
nand U1973 (N_1973,N_1771,N_1670);
and U1974 (N_1974,N_1773,N_1764);
xnor U1975 (N_1975,N_1600,N_1617);
and U1976 (N_1976,N_1789,N_1745);
xor U1977 (N_1977,N_1757,N_1704);
xor U1978 (N_1978,N_1732,N_1735);
nor U1979 (N_1979,N_1654,N_1671);
and U1980 (N_1980,N_1692,N_1781);
xnor U1981 (N_1981,N_1602,N_1712);
and U1982 (N_1982,N_1611,N_1781);
or U1983 (N_1983,N_1603,N_1602);
or U1984 (N_1984,N_1695,N_1607);
nand U1985 (N_1985,N_1707,N_1752);
xor U1986 (N_1986,N_1754,N_1720);
or U1987 (N_1987,N_1686,N_1720);
and U1988 (N_1988,N_1785,N_1619);
xor U1989 (N_1989,N_1741,N_1604);
and U1990 (N_1990,N_1648,N_1790);
nand U1991 (N_1991,N_1686,N_1634);
xnor U1992 (N_1992,N_1729,N_1641);
or U1993 (N_1993,N_1682,N_1655);
nand U1994 (N_1994,N_1633,N_1756);
or U1995 (N_1995,N_1720,N_1751);
nand U1996 (N_1996,N_1738,N_1782);
and U1997 (N_1997,N_1692,N_1688);
nand U1998 (N_1998,N_1667,N_1641);
nor U1999 (N_1999,N_1708,N_1735);
or U2000 (N_2000,N_1916,N_1815);
nand U2001 (N_2001,N_1863,N_1821);
or U2002 (N_2002,N_1928,N_1858);
nand U2003 (N_2003,N_1828,N_1989);
xnor U2004 (N_2004,N_1992,N_1820);
xor U2005 (N_2005,N_1999,N_1813);
and U2006 (N_2006,N_1801,N_1852);
and U2007 (N_2007,N_1873,N_1956);
or U2008 (N_2008,N_1908,N_1853);
xor U2009 (N_2009,N_1847,N_1855);
nor U2010 (N_2010,N_1915,N_1874);
or U2011 (N_2011,N_1904,N_1805);
nand U2012 (N_2012,N_1800,N_1802);
or U2013 (N_2013,N_1954,N_1885);
xnor U2014 (N_2014,N_1881,N_1948);
nand U2015 (N_2015,N_1832,N_1955);
nand U2016 (N_2016,N_1930,N_1838);
or U2017 (N_2017,N_1897,N_1834);
xor U2018 (N_2018,N_1899,N_1988);
xor U2019 (N_2019,N_1917,N_1937);
nor U2020 (N_2020,N_1976,N_1825);
and U2021 (N_2021,N_1840,N_1887);
and U2022 (N_2022,N_1934,N_1890);
or U2023 (N_2023,N_1895,N_1923);
and U2024 (N_2024,N_1991,N_1967);
xor U2025 (N_2025,N_1811,N_1851);
nand U2026 (N_2026,N_1869,N_1918);
or U2027 (N_2027,N_1886,N_1819);
and U2028 (N_2028,N_1902,N_1818);
nand U2029 (N_2029,N_1817,N_1835);
or U2030 (N_2030,N_1866,N_1994);
xor U2031 (N_2031,N_1953,N_1803);
nand U2032 (N_2032,N_1868,N_1824);
or U2033 (N_2033,N_1949,N_1943);
and U2034 (N_2034,N_1891,N_1827);
nor U2035 (N_2035,N_1935,N_1946);
nand U2036 (N_2036,N_1939,N_1896);
xnor U2037 (N_2037,N_1972,N_1987);
and U2038 (N_2038,N_1849,N_1965);
and U2039 (N_2039,N_1977,N_1841);
and U2040 (N_2040,N_1839,N_1984);
nor U2041 (N_2041,N_1900,N_1993);
nand U2042 (N_2042,N_1836,N_1812);
nand U2043 (N_2043,N_1964,N_1959);
nand U2044 (N_2044,N_1906,N_1960);
xor U2045 (N_2045,N_1962,N_1971);
and U2046 (N_2046,N_1814,N_1850);
and U2047 (N_2047,N_1951,N_1975);
nor U2048 (N_2048,N_1846,N_1995);
nor U2049 (N_2049,N_1907,N_1912);
nand U2050 (N_2050,N_1926,N_1982);
nand U2051 (N_2051,N_1894,N_1856);
nor U2052 (N_2052,N_1898,N_1878);
or U2053 (N_2053,N_1867,N_1889);
and U2054 (N_2054,N_1997,N_1854);
xnor U2055 (N_2055,N_1986,N_1950);
and U2056 (N_2056,N_1913,N_1882);
xnor U2057 (N_2057,N_1901,N_1978);
nand U2058 (N_2058,N_1870,N_1941);
or U2059 (N_2059,N_1809,N_1826);
nand U2060 (N_2060,N_1998,N_1892);
nor U2061 (N_2061,N_1810,N_1921);
or U2062 (N_2062,N_1961,N_1911);
nand U2063 (N_2063,N_1940,N_1914);
nor U2064 (N_2064,N_1981,N_1958);
or U2065 (N_2065,N_1945,N_1974);
and U2066 (N_2066,N_1859,N_1942);
xnor U2067 (N_2067,N_1936,N_1932);
xor U2068 (N_2068,N_1833,N_1860);
or U2069 (N_2069,N_1876,N_1883);
nor U2070 (N_2070,N_1808,N_1933);
nor U2071 (N_2071,N_1922,N_1944);
or U2072 (N_2072,N_1990,N_1872);
nor U2073 (N_2073,N_1980,N_1862);
nand U2074 (N_2074,N_1848,N_1842);
xor U2075 (N_2075,N_1947,N_1963);
nand U2076 (N_2076,N_1807,N_1816);
xnor U2077 (N_2077,N_1966,N_1925);
xnor U2078 (N_2078,N_1844,N_1970);
nor U2079 (N_2079,N_1893,N_1861);
or U2080 (N_2080,N_1865,N_1831);
and U2081 (N_2081,N_1829,N_1837);
and U2082 (N_2082,N_1938,N_1822);
xor U2083 (N_2083,N_1924,N_1968);
and U2084 (N_2084,N_1843,N_1905);
nor U2085 (N_2085,N_1804,N_1830);
xor U2086 (N_2086,N_1823,N_1920);
and U2087 (N_2087,N_1877,N_1871);
and U2088 (N_2088,N_1879,N_1909);
xnor U2089 (N_2089,N_1919,N_1857);
nor U2090 (N_2090,N_1910,N_1985);
nand U2091 (N_2091,N_1884,N_1979);
xnor U2092 (N_2092,N_1969,N_1929);
xnor U2093 (N_2093,N_1888,N_1880);
nor U2094 (N_2094,N_1875,N_1845);
xnor U2095 (N_2095,N_1864,N_1973);
and U2096 (N_2096,N_1806,N_1903);
and U2097 (N_2097,N_1952,N_1927);
nand U2098 (N_2098,N_1996,N_1983);
and U2099 (N_2099,N_1957,N_1931);
and U2100 (N_2100,N_1994,N_1808);
nand U2101 (N_2101,N_1824,N_1981);
xnor U2102 (N_2102,N_1857,N_1959);
or U2103 (N_2103,N_1870,N_1886);
and U2104 (N_2104,N_1972,N_1901);
or U2105 (N_2105,N_1909,N_1818);
nand U2106 (N_2106,N_1935,N_1841);
nand U2107 (N_2107,N_1972,N_1990);
and U2108 (N_2108,N_1877,N_1813);
nand U2109 (N_2109,N_1871,N_1844);
and U2110 (N_2110,N_1854,N_1971);
xnor U2111 (N_2111,N_1931,N_1960);
and U2112 (N_2112,N_1839,N_1807);
xor U2113 (N_2113,N_1880,N_1969);
xnor U2114 (N_2114,N_1989,N_1907);
and U2115 (N_2115,N_1914,N_1986);
xor U2116 (N_2116,N_1994,N_1908);
xnor U2117 (N_2117,N_1882,N_1824);
or U2118 (N_2118,N_1894,N_1928);
nand U2119 (N_2119,N_1933,N_1957);
nor U2120 (N_2120,N_1924,N_1926);
and U2121 (N_2121,N_1850,N_1940);
nand U2122 (N_2122,N_1860,N_1945);
xnor U2123 (N_2123,N_1821,N_1884);
nor U2124 (N_2124,N_1857,N_1887);
and U2125 (N_2125,N_1843,N_1807);
nor U2126 (N_2126,N_1846,N_1918);
and U2127 (N_2127,N_1807,N_1953);
nor U2128 (N_2128,N_1856,N_1805);
nand U2129 (N_2129,N_1952,N_1894);
nand U2130 (N_2130,N_1991,N_1893);
nand U2131 (N_2131,N_1816,N_1889);
xnor U2132 (N_2132,N_1988,N_1917);
and U2133 (N_2133,N_1856,N_1974);
nand U2134 (N_2134,N_1893,N_1921);
and U2135 (N_2135,N_1924,N_1859);
nand U2136 (N_2136,N_1997,N_1956);
or U2137 (N_2137,N_1830,N_1936);
or U2138 (N_2138,N_1841,N_1947);
nand U2139 (N_2139,N_1814,N_1922);
nand U2140 (N_2140,N_1988,N_1981);
nand U2141 (N_2141,N_1844,N_1815);
or U2142 (N_2142,N_1974,N_1815);
nor U2143 (N_2143,N_1965,N_1919);
and U2144 (N_2144,N_1802,N_1883);
nor U2145 (N_2145,N_1834,N_1908);
nor U2146 (N_2146,N_1853,N_1810);
and U2147 (N_2147,N_1962,N_1923);
or U2148 (N_2148,N_1865,N_1892);
nand U2149 (N_2149,N_1815,N_1910);
xor U2150 (N_2150,N_1842,N_1904);
nor U2151 (N_2151,N_1979,N_1911);
and U2152 (N_2152,N_1800,N_1954);
and U2153 (N_2153,N_1866,N_1968);
and U2154 (N_2154,N_1975,N_1954);
nand U2155 (N_2155,N_1850,N_1921);
or U2156 (N_2156,N_1977,N_1840);
nand U2157 (N_2157,N_1948,N_1831);
nand U2158 (N_2158,N_1886,N_1987);
nand U2159 (N_2159,N_1874,N_1983);
xor U2160 (N_2160,N_1906,N_1812);
nand U2161 (N_2161,N_1976,N_1967);
and U2162 (N_2162,N_1819,N_1945);
xnor U2163 (N_2163,N_1837,N_1834);
or U2164 (N_2164,N_1836,N_1951);
nor U2165 (N_2165,N_1812,N_1913);
xor U2166 (N_2166,N_1909,N_1852);
nor U2167 (N_2167,N_1963,N_1841);
or U2168 (N_2168,N_1863,N_1902);
nand U2169 (N_2169,N_1810,N_1979);
and U2170 (N_2170,N_1922,N_1853);
and U2171 (N_2171,N_1932,N_1856);
nand U2172 (N_2172,N_1901,N_1875);
xor U2173 (N_2173,N_1946,N_1833);
nor U2174 (N_2174,N_1811,N_1973);
or U2175 (N_2175,N_1889,N_1887);
or U2176 (N_2176,N_1897,N_1837);
nor U2177 (N_2177,N_1900,N_1847);
nand U2178 (N_2178,N_1973,N_1962);
nor U2179 (N_2179,N_1835,N_1991);
nor U2180 (N_2180,N_1875,N_1861);
and U2181 (N_2181,N_1960,N_1871);
nand U2182 (N_2182,N_1856,N_1833);
xnor U2183 (N_2183,N_1907,N_1854);
or U2184 (N_2184,N_1939,N_1905);
nor U2185 (N_2185,N_1924,N_1958);
xnor U2186 (N_2186,N_1815,N_1955);
or U2187 (N_2187,N_1837,N_1805);
and U2188 (N_2188,N_1997,N_1839);
xnor U2189 (N_2189,N_1961,N_1945);
nand U2190 (N_2190,N_1970,N_1818);
nand U2191 (N_2191,N_1810,N_1920);
xnor U2192 (N_2192,N_1982,N_1844);
xnor U2193 (N_2193,N_1814,N_1897);
and U2194 (N_2194,N_1875,N_1863);
or U2195 (N_2195,N_1815,N_1973);
or U2196 (N_2196,N_1813,N_1821);
nand U2197 (N_2197,N_1948,N_1955);
nand U2198 (N_2198,N_1989,N_1982);
and U2199 (N_2199,N_1909,N_1943);
xor U2200 (N_2200,N_2128,N_2012);
and U2201 (N_2201,N_2075,N_2073);
nand U2202 (N_2202,N_2107,N_2052);
or U2203 (N_2203,N_2105,N_2114);
nor U2204 (N_2204,N_2069,N_2032);
or U2205 (N_2205,N_2008,N_2002);
and U2206 (N_2206,N_2095,N_2017);
nor U2207 (N_2207,N_2184,N_2005);
and U2208 (N_2208,N_2113,N_2187);
nor U2209 (N_2209,N_2010,N_2104);
nand U2210 (N_2210,N_2155,N_2124);
nand U2211 (N_2211,N_2197,N_2011);
or U2212 (N_2212,N_2083,N_2175);
and U2213 (N_2213,N_2072,N_2021);
xor U2214 (N_2214,N_2089,N_2167);
and U2215 (N_2215,N_2020,N_2037);
xor U2216 (N_2216,N_2051,N_2134);
xnor U2217 (N_2217,N_2192,N_2179);
nor U2218 (N_2218,N_2038,N_2186);
xnor U2219 (N_2219,N_2022,N_2120);
xor U2220 (N_2220,N_2149,N_2042);
or U2221 (N_2221,N_2048,N_2088);
and U2222 (N_2222,N_2090,N_2176);
nand U2223 (N_2223,N_2045,N_2119);
nor U2224 (N_2224,N_2111,N_2106);
and U2225 (N_2225,N_2157,N_2018);
and U2226 (N_2226,N_2071,N_2150);
xor U2227 (N_2227,N_2057,N_2101);
and U2228 (N_2228,N_2188,N_2094);
or U2229 (N_2229,N_2193,N_2076);
xnor U2230 (N_2230,N_2023,N_2098);
nand U2231 (N_2231,N_2161,N_2028);
xor U2232 (N_2232,N_2151,N_2189);
or U2233 (N_2233,N_2046,N_2178);
and U2234 (N_2234,N_2040,N_2183);
or U2235 (N_2235,N_2004,N_2171);
or U2236 (N_2236,N_2116,N_2031);
nor U2237 (N_2237,N_2136,N_2109);
nand U2238 (N_2238,N_2064,N_2047);
and U2239 (N_2239,N_2190,N_2182);
nor U2240 (N_2240,N_2156,N_2198);
or U2241 (N_2241,N_2035,N_2082);
nor U2242 (N_2242,N_2122,N_2146);
xor U2243 (N_2243,N_2180,N_2170);
and U2244 (N_2244,N_2139,N_2079);
nor U2245 (N_2245,N_2063,N_2078);
xor U2246 (N_2246,N_2026,N_2043);
nor U2247 (N_2247,N_2056,N_2177);
xor U2248 (N_2248,N_2027,N_2108);
nand U2249 (N_2249,N_2148,N_2133);
or U2250 (N_2250,N_2129,N_2112);
nand U2251 (N_2251,N_2085,N_2102);
nor U2252 (N_2252,N_2044,N_2121);
and U2253 (N_2253,N_2166,N_2060);
and U2254 (N_2254,N_2172,N_2123);
or U2255 (N_2255,N_2093,N_2066);
or U2256 (N_2256,N_2131,N_2096);
nand U2257 (N_2257,N_2086,N_2194);
or U2258 (N_2258,N_2053,N_2055);
nand U2259 (N_2259,N_2158,N_2103);
and U2260 (N_2260,N_2081,N_2135);
nand U2261 (N_2261,N_2054,N_2185);
xor U2262 (N_2262,N_2117,N_2062);
and U2263 (N_2263,N_2007,N_2145);
or U2264 (N_2264,N_2015,N_2140);
or U2265 (N_2265,N_2169,N_2191);
and U2266 (N_2266,N_2126,N_2065);
nand U2267 (N_2267,N_2195,N_2059);
or U2268 (N_2268,N_2036,N_2009);
and U2269 (N_2269,N_2100,N_2199);
nor U2270 (N_2270,N_2067,N_2118);
xor U2271 (N_2271,N_2013,N_2070);
xnor U2272 (N_2272,N_2153,N_2181);
xor U2273 (N_2273,N_2132,N_2000);
nand U2274 (N_2274,N_2029,N_2001);
nor U2275 (N_2275,N_2003,N_2050);
and U2276 (N_2276,N_2077,N_2039);
nor U2277 (N_2277,N_2041,N_2092);
nand U2278 (N_2278,N_2137,N_2173);
and U2279 (N_2279,N_2061,N_2033);
xnor U2280 (N_2280,N_2142,N_2163);
and U2281 (N_2281,N_2080,N_2141);
nand U2282 (N_2282,N_2196,N_2084);
xor U2283 (N_2283,N_2160,N_2049);
or U2284 (N_2284,N_2068,N_2099);
nand U2285 (N_2285,N_2014,N_2152);
xor U2286 (N_2286,N_2074,N_2144);
nand U2287 (N_2287,N_2034,N_2110);
or U2288 (N_2288,N_2143,N_2165);
or U2289 (N_2289,N_2168,N_2030);
xor U2290 (N_2290,N_2154,N_2025);
and U2291 (N_2291,N_2138,N_2016);
and U2292 (N_2292,N_2091,N_2174);
and U2293 (N_2293,N_2019,N_2162);
or U2294 (N_2294,N_2024,N_2164);
nor U2295 (N_2295,N_2087,N_2115);
nand U2296 (N_2296,N_2147,N_2097);
xnor U2297 (N_2297,N_2159,N_2058);
or U2298 (N_2298,N_2130,N_2125);
nand U2299 (N_2299,N_2006,N_2127);
nor U2300 (N_2300,N_2135,N_2089);
and U2301 (N_2301,N_2195,N_2175);
or U2302 (N_2302,N_2134,N_2132);
and U2303 (N_2303,N_2085,N_2182);
nor U2304 (N_2304,N_2106,N_2182);
xnor U2305 (N_2305,N_2160,N_2046);
nor U2306 (N_2306,N_2050,N_2146);
nor U2307 (N_2307,N_2035,N_2099);
or U2308 (N_2308,N_2028,N_2059);
xor U2309 (N_2309,N_2106,N_2070);
nand U2310 (N_2310,N_2050,N_2099);
xnor U2311 (N_2311,N_2194,N_2136);
xor U2312 (N_2312,N_2170,N_2179);
or U2313 (N_2313,N_2175,N_2015);
nand U2314 (N_2314,N_2144,N_2182);
nor U2315 (N_2315,N_2039,N_2134);
xnor U2316 (N_2316,N_2139,N_2153);
and U2317 (N_2317,N_2151,N_2166);
xnor U2318 (N_2318,N_2138,N_2199);
nand U2319 (N_2319,N_2187,N_2115);
nor U2320 (N_2320,N_2094,N_2179);
or U2321 (N_2321,N_2015,N_2160);
nor U2322 (N_2322,N_2022,N_2121);
nand U2323 (N_2323,N_2120,N_2055);
or U2324 (N_2324,N_2073,N_2142);
nand U2325 (N_2325,N_2114,N_2029);
xor U2326 (N_2326,N_2183,N_2050);
and U2327 (N_2327,N_2198,N_2171);
nor U2328 (N_2328,N_2142,N_2080);
xor U2329 (N_2329,N_2103,N_2062);
and U2330 (N_2330,N_2090,N_2173);
or U2331 (N_2331,N_2042,N_2088);
xnor U2332 (N_2332,N_2121,N_2106);
nor U2333 (N_2333,N_2167,N_2023);
nand U2334 (N_2334,N_2102,N_2026);
or U2335 (N_2335,N_2001,N_2075);
xor U2336 (N_2336,N_2116,N_2152);
nand U2337 (N_2337,N_2086,N_2128);
nor U2338 (N_2338,N_2185,N_2052);
nor U2339 (N_2339,N_2191,N_2116);
or U2340 (N_2340,N_2195,N_2142);
xor U2341 (N_2341,N_2193,N_2188);
and U2342 (N_2342,N_2013,N_2150);
nand U2343 (N_2343,N_2071,N_2026);
xor U2344 (N_2344,N_2002,N_2057);
nand U2345 (N_2345,N_2173,N_2130);
xnor U2346 (N_2346,N_2153,N_2011);
nor U2347 (N_2347,N_2089,N_2104);
nor U2348 (N_2348,N_2093,N_2062);
xor U2349 (N_2349,N_2056,N_2129);
nand U2350 (N_2350,N_2012,N_2182);
xor U2351 (N_2351,N_2129,N_2055);
xor U2352 (N_2352,N_2033,N_2002);
nand U2353 (N_2353,N_2121,N_2078);
and U2354 (N_2354,N_2025,N_2008);
xor U2355 (N_2355,N_2005,N_2031);
nand U2356 (N_2356,N_2061,N_2170);
xnor U2357 (N_2357,N_2043,N_2000);
xnor U2358 (N_2358,N_2100,N_2031);
nor U2359 (N_2359,N_2138,N_2013);
nand U2360 (N_2360,N_2102,N_2076);
nand U2361 (N_2361,N_2023,N_2055);
and U2362 (N_2362,N_2106,N_2016);
and U2363 (N_2363,N_2103,N_2174);
nand U2364 (N_2364,N_2185,N_2105);
nand U2365 (N_2365,N_2025,N_2157);
nand U2366 (N_2366,N_2135,N_2049);
nand U2367 (N_2367,N_2087,N_2192);
or U2368 (N_2368,N_2118,N_2162);
xor U2369 (N_2369,N_2159,N_2190);
nor U2370 (N_2370,N_2156,N_2103);
nand U2371 (N_2371,N_2138,N_2180);
or U2372 (N_2372,N_2039,N_2178);
and U2373 (N_2373,N_2166,N_2020);
and U2374 (N_2374,N_2089,N_2117);
xor U2375 (N_2375,N_2130,N_2191);
nor U2376 (N_2376,N_2059,N_2162);
xor U2377 (N_2377,N_2157,N_2030);
nor U2378 (N_2378,N_2103,N_2189);
nand U2379 (N_2379,N_2045,N_2106);
and U2380 (N_2380,N_2141,N_2122);
or U2381 (N_2381,N_2144,N_2056);
nand U2382 (N_2382,N_2131,N_2021);
xor U2383 (N_2383,N_2076,N_2075);
or U2384 (N_2384,N_2145,N_2121);
and U2385 (N_2385,N_2058,N_2004);
nor U2386 (N_2386,N_2070,N_2095);
and U2387 (N_2387,N_2074,N_2194);
xor U2388 (N_2388,N_2063,N_2089);
or U2389 (N_2389,N_2100,N_2193);
xnor U2390 (N_2390,N_2028,N_2083);
and U2391 (N_2391,N_2184,N_2001);
nor U2392 (N_2392,N_2061,N_2001);
nor U2393 (N_2393,N_2152,N_2017);
and U2394 (N_2394,N_2100,N_2064);
and U2395 (N_2395,N_2111,N_2035);
or U2396 (N_2396,N_2076,N_2156);
xor U2397 (N_2397,N_2120,N_2015);
xnor U2398 (N_2398,N_2037,N_2133);
and U2399 (N_2399,N_2173,N_2077);
xnor U2400 (N_2400,N_2270,N_2344);
nand U2401 (N_2401,N_2259,N_2300);
xnor U2402 (N_2402,N_2252,N_2295);
or U2403 (N_2403,N_2278,N_2366);
nand U2404 (N_2404,N_2392,N_2244);
xor U2405 (N_2405,N_2239,N_2238);
nor U2406 (N_2406,N_2380,N_2387);
xnor U2407 (N_2407,N_2318,N_2216);
or U2408 (N_2408,N_2266,N_2398);
and U2409 (N_2409,N_2315,N_2378);
or U2410 (N_2410,N_2274,N_2210);
and U2411 (N_2411,N_2208,N_2372);
xor U2412 (N_2412,N_2396,N_2258);
nand U2413 (N_2413,N_2303,N_2355);
nand U2414 (N_2414,N_2296,N_2217);
nor U2415 (N_2415,N_2271,N_2334);
or U2416 (N_2416,N_2230,N_2360);
nand U2417 (N_2417,N_2348,N_2291);
nand U2418 (N_2418,N_2337,N_2367);
or U2419 (N_2419,N_2317,N_2322);
xnor U2420 (N_2420,N_2307,N_2316);
nand U2421 (N_2421,N_2356,N_2235);
and U2422 (N_2422,N_2202,N_2393);
xnor U2423 (N_2423,N_2373,N_2394);
nor U2424 (N_2424,N_2286,N_2345);
xnor U2425 (N_2425,N_2326,N_2350);
nand U2426 (N_2426,N_2320,N_2285);
xnor U2427 (N_2427,N_2383,N_2292);
and U2428 (N_2428,N_2395,N_2377);
or U2429 (N_2429,N_2241,N_2282);
nor U2430 (N_2430,N_2375,N_2341);
or U2431 (N_2431,N_2261,N_2243);
or U2432 (N_2432,N_2200,N_2226);
and U2433 (N_2433,N_2294,N_2240);
and U2434 (N_2434,N_2354,N_2343);
nand U2435 (N_2435,N_2263,N_2273);
nand U2436 (N_2436,N_2390,N_2242);
nor U2437 (N_2437,N_2385,N_2249);
xnor U2438 (N_2438,N_2370,N_2301);
nor U2439 (N_2439,N_2359,N_2229);
nand U2440 (N_2440,N_2212,N_2260);
and U2441 (N_2441,N_2201,N_2311);
or U2442 (N_2442,N_2289,N_2265);
xnor U2443 (N_2443,N_2335,N_2379);
xor U2444 (N_2444,N_2330,N_2310);
nor U2445 (N_2445,N_2227,N_2209);
xnor U2446 (N_2446,N_2205,N_2281);
and U2447 (N_2447,N_2299,N_2399);
nor U2448 (N_2448,N_2207,N_2371);
nand U2449 (N_2449,N_2228,N_2336);
or U2450 (N_2450,N_2255,N_2357);
or U2451 (N_2451,N_2369,N_2232);
nor U2452 (N_2452,N_2327,N_2251);
or U2453 (N_2453,N_2352,N_2331);
nor U2454 (N_2454,N_2287,N_2215);
nor U2455 (N_2455,N_2221,N_2256);
and U2456 (N_2456,N_2304,N_2204);
nor U2457 (N_2457,N_2237,N_2213);
and U2458 (N_2458,N_2333,N_2219);
and U2459 (N_2459,N_2342,N_2245);
or U2460 (N_2460,N_2293,N_2262);
or U2461 (N_2461,N_2218,N_2363);
or U2462 (N_2462,N_2314,N_2246);
nand U2463 (N_2463,N_2203,N_2358);
xnor U2464 (N_2464,N_2381,N_2234);
and U2465 (N_2465,N_2211,N_2384);
xnor U2466 (N_2466,N_2306,N_2220);
or U2467 (N_2467,N_2288,N_2298);
or U2468 (N_2468,N_2214,N_2361);
nand U2469 (N_2469,N_2364,N_2386);
nand U2470 (N_2470,N_2225,N_2332);
nand U2471 (N_2471,N_2305,N_2284);
nor U2472 (N_2472,N_2312,N_2276);
and U2473 (N_2473,N_2272,N_2279);
or U2474 (N_2474,N_2323,N_2376);
or U2475 (N_2475,N_2267,N_2338);
nand U2476 (N_2476,N_2297,N_2222);
xor U2477 (N_2477,N_2250,N_2277);
xnor U2478 (N_2478,N_2247,N_2268);
xnor U2479 (N_2479,N_2257,N_2391);
xor U2480 (N_2480,N_2264,N_2302);
nand U2481 (N_2481,N_2321,N_2280);
nand U2482 (N_2482,N_2254,N_2224);
nand U2483 (N_2483,N_2382,N_2236);
xor U2484 (N_2484,N_2324,N_2340);
nand U2485 (N_2485,N_2290,N_2206);
xnor U2486 (N_2486,N_2319,N_2339);
xnor U2487 (N_2487,N_2253,N_2275);
nor U2488 (N_2488,N_2353,N_2389);
and U2489 (N_2489,N_2308,N_2347);
nand U2490 (N_2490,N_2365,N_2325);
xor U2491 (N_2491,N_2223,N_2362);
xnor U2492 (N_2492,N_2388,N_2328);
xnor U2493 (N_2493,N_2349,N_2231);
xnor U2494 (N_2494,N_2248,N_2346);
nand U2495 (N_2495,N_2374,N_2283);
or U2496 (N_2496,N_2329,N_2269);
or U2497 (N_2497,N_2309,N_2313);
nor U2498 (N_2498,N_2351,N_2397);
and U2499 (N_2499,N_2368,N_2233);
or U2500 (N_2500,N_2232,N_2279);
xor U2501 (N_2501,N_2381,N_2244);
or U2502 (N_2502,N_2346,N_2237);
xor U2503 (N_2503,N_2211,N_2374);
nor U2504 (N_2504,N_2240,N_2327);
or U2505 (N_2505,N_2273,N_2250);
xnor U2506 (N_2506,N_2391,N_2204);
and U2507 (N_2507,N_2206,N_2298);
xnor U2508 (N_2508,N_2385,N_2384);
nor U2509 (N_2509,N_2333,N_2324);
nand U2510 (N_2510,N_2339,N_2346);
nor U2511 (N_2511,N_2216,N_2252);
nand U2512 (N_2512,N_2356,N_2368);
nand U2513 (N_2513,N_2336,N_2351);
nand U2514 (N_2514,N_2301,N_2300);
xnor U2515 (N_2515,N_2207,N_2343);
or U2516 (N_2516,N_2325,N_2316);
nor U2517 (N_2517,N_2343,N_2280);
and U2518 (N_2518,N_2385,N_2257);
xnor U2519 (N_2519,N_2318,N_2326);
and U2520 (N_2520,N_2377,N_2356);
nor U2521 (N_2521,N_2259,N_2310);
and U2522 (N_2522,N_2223,N_2352);
nand U2523 (N_2523,N_2267,N_2210);
xnor U2524 (N_2524,N_2233,N_2361);
xor U2525 (N_2525,N_2202,N_2390);
and U2526 (N_2526,N_2336,N_2294);
nor U2527 (N_2527,N_2356,N_2352);
and U2528 (N_2528,N_2380,N_2245);
or U2529 (N_2529,N_2319,N_2353);
xnor U2530 (N_2530,N_2299,N_2363);
and U2531 (N_2531,N_2374,N_2237);
nand U2532 (N_2532,N_2243,N_2226);
nand U2533 (N_2533,N_2290,N_2308);
xnor U2534 (N_2534,N_2253,N_2332);
and U2535 (N_2535,N_2367,N_2320);
and U2536 (N_2536,N_2328,N_2294);
nand U2537 (N_2537,N_2231,N_2253);
xor U2538 (N_2538,N_2238,N_2348);
and U2539 (N_2539,N_2217,N_2344);
and U2540 (N_2540,N_2377,N_2294);
nand U2541 (N_2541,N_2259,N_2333);
and U2542 (N_2542,N_2354,N_2353);
nor U2543 (N_2543,N_2375,N_2310);
nand U2544 (N_2544,N_2384,N_2285);
nand U2545 (N_2545,N_2201,N_2247);
or U2546 (N_2546,N_2258,N_2376);
xor U2547 (N_2547,N_2216,N_2288);
or U2548 (N_2548,N_2205,N_2260);
or U2549 (N_2549,N_2390,N_2223);
nand U2550 (N_2550,N_2231,N_2382);
xor U2551 (N_2551,N_2365,N_2210);
nor U2552 (N_2552,N_2271,N_2354);
nand U2553 (N_2553,N_2233,N_2379);
and U2554 (N_2554,N_2357,N_2350);
nor U2555 (N_2555,N_2206,N_2259);
nand U2556 (N_2556,N_2330,N_2309);
nand U2557 (N_2557,N_2388,N_2272);
nor U2558 (N_2558,N_2246,N_2219);
and U2559 (N_2559,N_2321,N_2371);
xnor U2560 (N_2560,N_2264,N_2337);
nor U2561 (N_2561,N_2246,N_2204);
or U2562 (N_2562,N_2361,N_2339);
nor U2563 (N_2563,N_2321,N_2247);
nand U2564 (N_2564,N_2203,N_2236);
and U2565 (N_2565,N_2360,N_2365);
nor U2566 (N_2566,N_2358,N_2290);
nor U2567 (N_2567,N_2373,N_2254);
nand U2568 (N_2568,N_2291,N_2373);
nand U2569 (N_2569,N_2307,N_2356);
or U2570 (N_2570,N_2350,N_2297);
xor U2571 (N_2571,N_2325,N_2345);
nand U2572 (N_2572,N_2374,N_2342);
nor U2573 (N_2573,N_2264,N_2259);
nand U2574 (N_2574,N_2248,N_2265);
and U2575 (N_2575,N_2391,N_2212);
or U2576 (N_2576,N_2227,N_2291);
xor U2577 (N_2577,N_2336,N_2378);
and U2578 (N_2578,N_2223,N_2300);
nand U2579 (N_2579,N_2228,N_2327);
and U2580 (N_2580,N_2218,N_2289);
xor U2581 (N_2581,N_2388,N_2346);
nor U2582 (N_2582,N_2213,N_2318);
nor U2583 (N_2583,N_2396,N_2382);
nor U2584 (N_2584,N_2311,N_2359);
or U2585 (N_2585,N_2323,N_2304);
xor U2586 (N_2586,N_2393,N_2244);
nor U2587 (N_2587,N_2259,N_2219);
nand U2588 (N_2588,N_2292,N_2225);
xor U2589 (N_2589,N_2377,N_2243);
or U2590 (N_2590,N_2261,N_2270);
nor U2591 (N_2591,N_2347,N_2317);
xor U2592 (N_2592,N_2377,N_2242);
xnor U2593 (N_2593,N_2235,N_2296);
nor U2594 (N_2594,N_2229,N_2246);
nand U2595 (N_2595,N_2393,N_2307);
nor U2596 (N_2596,N_2330,N_2271);
xor U2597 (N_2597,N_2267,N_2373);
nand U2598 (N_2598,N_2201,N_2273);
and U2599 (N_2599,N_2352,N_2314);
nand U2600 (N_2600,N_2592,N_2434);
xnor U2601 (N_2601,N_2491,N_2402);
nand U2602 (N_2602,N_2408,N_2435);
or U2603 (N_2603,N_2578,N_2401);
xor U2604 (N_2604,N_2573,N_2502);
and U2605 (N_2605,N_2597,N_2589);
nor U2606 (N_2606,N_2547,N_2492);
xnor U2607 (N_2607,N_2555,N_2407);
nand U2608 (N_2608,N_2579,N_2413);
nor U2609 (N_2609,N_2419,N_2409);
nor U2610 (N_2610,N_2465,N_2454);
and U2611 (N_2611,N_2554,N_2473);
nor U2612 (N_2612,N_2459,N_2500);
and U2613 (N_2613,N_2405,N_2521);
and U2614 (N_2614,N_2486,N_2525);
and U2615 (N_2615,N_2537,N_2479);
and U2616 (N_2616,N_2545,N_2447);
xor U2617 (N_2617,N_2553,N_2540);
and U2618 (N_2618,N_2508,N_2582);
xor U2619 (N_2619,N_2507,N_2460);
nor U2620 (N_2620,N_2535,N_2478);
and U2621 (N_2621,N_2498,N_2594);
or U2622 (N_2622,N_2511,N_2475);
xor U2623 (N_2623,N_2504,N_2449);
nand U2624 (N_2624,N_2416,N_2559);
or U2625 (N_2625,N_2466,N_2448);
xor U2626 (N_2626,N_2506,N_2562);
nor U2627 (N_2627,N_2595,N_2468);
nor U2628 (N_2628,N_2438,N_2539);
or U2629 (N_2629,N_2489,N_2463);
or U2630 (N_2630,N_2569,N_2563);
and U2631 (N_2631,N_2567,N_2546);
nand U2632 (N_2632,N_2445,N_2565);
nor U2633 (N_2633,N_2484,N_2471);
nor U2634 (N_2634,N_2568,N_2517);
nor U2635 (N_2635,N_2423,N_2404);
nor U2636 (N_2636,N_2572,N_2426);
or U2637 (N_2637,N_2580,N_2499);
and U2638 (N_2638,N_2487,N_2510);
nor U2639 (N_2639,N_2541,N_2431);
xor U2640 (N_2640,N_2470,N_2433);
or U2641 (N_2641,N_2482,N_2485);
nand U2642 (N_2642,N_2450,N_2457);
or U2643 (N_2643,N_2490,N_2526);
and U2644 (N_2644,N_2421,N_2436);
and U2645 (N_2645,N_2406,N_2453);
and U2646 (N_2646,N_2585,N_2509);
nand U2647 (N_2647,N_2429,N_2570);
or U2648 (N_2648,N_2528,N_2420);
xnor U2649 (N_2649,N_2455,N_2557);
nor U2650 (N_2650,N_2560,N_2469);
nor U2651 (N_2651,N_2530,N_2488);
and U2652 (N_2652,N_2503,N_2480);
or U2653 (N_2653,N_2415,N_2496);
and U2654 (N_2654,N_2456,N_2442);
xnor U2655 (N_2655,N_2577,N_2586);
or U2656 (N_2656,N_2495,N_2422);
nor U2657 (N_2657,N_2497,N_2593);
and U2658 (N_2658,N_2538,N_2583);
xor U2659 (N_2659,N_2519,N_2472);
nor U2660 (N_2660,N_2403,N_2516);
and U2661 (N_2661,N_2574,N_2414);
xnor U2662 (N_2662,N_2462,N_2514);
nand U2663 (N_2663,N_2513,N_2417);
or U2664 (N_2664,N_2400,N_2515);
nand U2665 (N_2665,N_2587,N_2552);
nor U2666 (N_2666,N_2461,N_2424);
nand U2667 (N_2667,N_2444,N_2428);
and U2668 (N_2668,N_2432,N_2576);
xnor U2669 (N_2669,N_2533,N_2571);
nand U2670 (N_2670,N_2598,N_2412);
nor U2671 (N_2671,N_2575,N_2590);
and U2672 (N_2672,N_2467,N_2451);
and U2673 (N_2673,N_2474,N_2440);
nand U2674 (N_2674,N_2452,N_2418);
nor U2675 (N_2675,N_2477,N_2561);
xor U2676 (N_2676,N_2476,N_2520);
xor U2677 (N_2677,N_2512,N_2558);
or U2678 (N_2678,N_2534,N_2518);
and U2679 (N_2679,N_2531,N_2548);
or U2680 (N_2680,N_2493,N_2481);
and U2681 (N_2681,N_2523,N_2529);
nor U2682 (N_2682,N_2441,N_2544);
and U2683 (N_2683,N_2501,N_2527);
nand U2684 (N_2684,N_2483,N_2410);
or U2685 (N_2685,N_2411,N_2551);
nor U2686 (N_2686,N_2443,N_2439);
xnor U2687 (N_2687,N_2599,N_2588);
or U2688 (N_2688,N_2542,N_2458);
and U2689 (N_2689,N_2430,N_2549);
nor U2690 (N_2690,N_2596,N_2446);
and U2691 (N_2691,N_2505,N_2532);
nor U2692 (N_2692,N_2494,N_2564);
or U2693 (N_2693,N_2464,N_2584);
nand U2694 (N_2694,N_2427,N_2566);
nand U2695 (N_2695,N_2425,N_2522);
or U2696 (N_2696,N_2524,N_2536);
xor U2697 (N_2697,N_2591,N_2550);
nor U2698 (N_2698,N_2581,N_2437);
and U2699 (N_2699,N_2556,N_2543);
or U2700 (N_2700,N_2504,N_2549);
nor U2701 (N_2701,N_2482,N_2541);
xnor U2702 (N_2702,N_2584,N_2434);
or U2703 (N_2703,N_2519,N_2579);
nand U2704 (N_2704,N_2572,N_2460);
xnor U2705 (N_2705,N_2577,N_2411);
and U2706 (N_2706,N_2523,N_2580);
or U2707 (N_2707,N_2402,N_2444);
nand U2708 (N_2708,N_2514,N_2513);
nand U2709 (N_2709,N_2432,N_2522);
nand U2710 (N_2710,N_2483,N_2528);
nand U2711 (N_2711,N_2484,N_2433);
nand U2712 (N_2712,N_2527,N_2573);
nor U2713 (N_2713,N_2599,N_2411);
and U2714 (N_2714,N_2554,N_2542);
nor U2715 (N_2715,N_2528,N_2422);
or U2716 (N_2716,N_2432,N_2498);
or U2717 (N_2717,N_2456,N_2451);
or U2718 (N_2718,N_2486,N_2448);
nand U2719 (N_2719,N_2547,N_2455);
nand U2720 (N_2720,N_2563,N_2524);
xor U2721 (N_2721,N_2483,N_2458);
nor U2722 (N_2722,N_2492,N_2576);
nor U2723 (N_2723,N_2408,N_2576);
and U2724 (N_2724,N_2417,N_2509);
xnor U2725 (N_2725,N_2595,N_2457);
and U2726 (N_2726,N_2550,N_2494);
nor U2727 (N_2727,N_2519,N_2590);
or U2728 (N_2728,N_2510,N_2486);
xor U2729 (N_2729,N_2451,N_2534);
nor U2730 (N_2730,N_2503,N_2520);
and U2731 (N_2731,N_2541,N_2420);
xor U2732 (N_2732,N_2445,N_2577);
nor U2733 (N_2733,N_2420,N_2521);
or U2734 (N_2734,N_2585,N_2512);
and U2735 (N_2735,N_2579,N_2571);
or U2736 (N_2736,N_2510,N_2437);
nor U2737 (N_2737,N_2529,N_2541);
nor U2738 (N_2738,N_2564,N_2501);
xnor U2739 (N_2739,N_2534,N_2475);
and U2740 (N_2740,N_2495,N_2538);
xnor U2741 (N_2741,N_2478,N_2528);
nor U2742 (N_2742,N_2478,N_2412);
and U2743 (N_2743,N_2484,N_2571);
xnor U2744 (N_2744,N_2489,N_2564);
nor U2745 (N_2745,N_2591,N_2411);
or U2746 (N_2746,N_2449,N_2414);
and U2747 (N_2747,N_2580,N_2571);
nand U2748 (N_2748,N_2491,N_2537);
and U2749 (N_2749,N_2597,N_2433);
and U2750 (N_2750,N_2537,N_2495);
nor U2751 (N_2751,N_2516,N_2527);
nand U2752 (N_2752,N_2581,N_2415);
and U2753 (N_2753,N_2433,N_2535);
xor U2754 (N_2754,N_2588,N_2582);
or U2755 (N_2755,N_2501,N_2480);
and U2756 (N_2756,N_2439,N_2560);
nor U2757 (N_2757,N_2418,N_2442);
nand U2758 (N_2758,N_2514,N_2488);
nand U2759 (N_2759,N_2420,N_2416);
and U2760 (N_2760,N_2436,N_2427);
or U2761 (N_2761,N_2552,N_2573);
or U2762 (N_2762,N_2585,N_2405);
nor U2763 (N_2763,N_2516,N_2487);
xnor U2764 (N_2764,N_2476,N_2589);
nor U2765 (N_2765,N_2491,N_2590);
xnor U2766 (N_2766,N_2560,N_2478);
nor U2767 (N_2767,N_2538,N_2454);
xor U2768 (N_2768,N_2409,N_2515);
or U2769 (N_2769,N_2465,N_2492);
nor U2770 (N_2770,N_2493,N_2438);
and U2771 (N_2771,N_2545,N_2569);
nand U2772 (N_2772,N_2468,N_2425);
nand U2773 (N_2773,N_2585,N_2456);
nor U2774 (N_2774,N_2550,N_2414);
nor U2775 (N_2775,N_2506,N_2503);
nor U2776 (N_2776,N_2560,N_2507);
xnor U2777 (N_2777,N_2455,N_2560);
or U2778 (N_2778,N_2574,N_2556);
or U2779 (N_2779,N_2558,N_2570);
or U2780 (N_2780,N_2559,N_2461);
and U2781 (N_2781,N_2423,N_2469);
xnor U2782 (N_2782,N_2523,N_2450);
nor U2783 (N_2783,N_2522,N_2483);
nand U2784 (N_2784,N_2486,N_2591);
nor U2785 (N_2785,N_2568,N_2580);
nand U2786 (N_2786,N_2524,N_2428);
nor U2787 (N_2787,N_2455,N_2513);
or U2788 (N_2788,N_2509,N_2482);
or U2789 (N_2789,N_2515,N_2565);
xnor U2790 (N_2790,N_2548,N_2412);
or U2791 (N_2791,N_2458,N_2569);
or U2792 (N_2792,N_2429,N_2458);
nand U2793 (N_2793,N_2554,N_2480);
or U2794 (N_2794,N_2590,N_2501);
and U2795 (N_2795,N_2465,N_2573);
xor U2796 (N_2796,N_2537,N_2551);
and U2797 (N_2797,N_2594,N_2402);
nand U2798 (N_2798,N_2583,N_2463);
or U2799 (N_2799,N_2410,N_2458);
xnor U2800 (N_2800,N_2778,N_2612);
xor U2801 (N_2801,N_2611,N_2729);
xnor U2802 (N_2802,N_2639,N_2730);
and U2803 (N_2803,N_2741,N_2796);
and U2804 (N_2804,N_2779,N_2621);
or U2805 (N_2805,N_2676,N_2750);
or U2806 (N_2806,N_2601,N_2638);
and U2807 (N_2807,N_2769,N_2764);
nand U2808 (N_2808,N_2687,N_2681);
and U2809 (N_2809,N_2757,N_2705);
nor U2810 (N_2810,N_2689,N_2618);
and U2811 (N_2811,N_2726,N_2628);
xnor U2812 (N_2812,N_2633,N_2771);
xor U2813 (N_2813,N_2780,N_2731);
and U2814 (N_2814,N_2747,N_2772);
nor U2815 (N_2815,N_2718,N_2746);
and U2816 (N_2816,N_2706,N_2708);
xnor U2817 (N_2817,N_2685,N_2697);
nor U2818 (N_2818,N_2652,N_2775);
nor U2819 (N_2819,N_2738,N_2716);
nand U2820 (N_2820,N_2720,N_2632);
xor U2821 (N_2821,N_2655,N_2784);
or U2822 (N_2822,N_2703,N_2760);
or U2823 (N_2823,N_2653,N_2785);
nor U2824 (N_2824,N_2758,N_2795);
nor U2825 (N_2825,N_2640,N_2677);
nor U2826 (N_2826,N_2651,N_2659);
and U2827 (N_2827,N_2732,N_2691);
or U2828 (N_2828,N_2709,N_2751);
nand U2829 (N_2829,N_2776,N_2641);
xor U2830 (N_2830,N_2695,N_2600);
xor U2831 (N_2831,N_2754,N_2622);
nand U2832 (N_2832,N_2770,N_2717);
xor U2833 (N_2833,N_2781,N_2745);
and U2834 (N_2834,N_2736,N_2635);
or U2835 (N_2835,N_2678,N_2684);
xnor U2836 (N_2836,N_2701,N_2753);
xor U2837 (N_2837,N_2671,N_2783);
nor U2838 (N_2838,N_2749,N_2714);
xor U2839 (N_2839,N_2735,N_2670);
or U2840 (N_2840,N_2723,N_2668);
or U2841 (N_2841,N_2752,N_2774);
nand U2842 (N_2842,N_2629,N_2667);
or U2843 (N_2843,N_2607,N_2767);
and U2844 (N_2844,N_2791,N_2644);
or U2845 (N_2845,N_2634,N_2623);
xnor U2846 (N_2846,N_2742,N_2664);
nor U2847 (N_2847,N_2782,N_2661);
xnor U2848 (N_2848,N_2759,N_2686);
xnor U2849 (N_2849,N_2626,N_2787);
or U2850 (N_2850,N_2704,N_2657);
nor U2851 (N_2851,N_2674,N_2692);
or U2852 (N_2852,N_2707,N_2693);
xnor U2853 (N_2853,N_2615,N_2696);
and U2854 (N_2854,N_2773,N_2762);
nand U2855 (N_2855,N_2719,N_2702);
xnor U2856 (N_2856,N_2700,N_2650);
and U2857 (N_2857,N_2665,N_2636);
nor U2858 (N_2858,N_2630,N_2797);
and U2859 (N_2859,N_2675,N_2649);
and U2860 (N_2860,N_2690,N_2763);
or U2861 (N_2861,N_2673,N_2765);
xnor U2862 (N_2862,N_2608,N_2660);
xnor U2863 (N_2863,N_2625,N_2679);
nand U2864 (N_2864,N_2711,N_2793);
xnor U2865 (N_2865,N_2603,N_2642);
xor U2866 (N_2866,N_2712,N_2799);
xor U2867 (N_2867,N_2604,N_2613);
nand U2868 (N_2868,N_2740,N_2788);
xor U2869 (N_2869,N_2728,N_2722);
xnor U2870 (N_2870,N_2658,N_2755);
nor U2871 (N_2871,N_2609,N_2798);
nand U2872 (N_2872,N_2744,N_2669);
nor U2873 (N_2873,N_2680,N_2683);
and U2874 (N_2874,N_2654,N_2648);
xnor U2875 (N_2875,N_2627,N_2663);
nor U2876 (N_2876,N_2616,N_2792);
nor U2877 (N_2877,N_2694,N_2656);
xor U2878 (N_2878,N_2768,N_2602);
nand U2879 (N_2879,N_2698,N_2624);
nand U2880 (N_2880,N_2733,N_2682);
xnor U2881 (N_2881,N_2614,N_2610);
nand U2882 (N_2882,N_2766,N_2748);
nor U2883 (N_2883,N_2743,N_2721);
nor U2884 (N_2884,N_2643,N_2605);
nand U2885 (N_2885,N_2637,N_2672);
nand U2886 (N_2886,N_2688,N_2646);
and U2887 (N_2887,N_2794,N_2725);
xnor U2888 (N_2888,N_2724,N_2620);
and U2889 (N_2889,N_2756,N_2715);
and U2890 (N_2890,N_2761,N_2727);
and U2891 (N_2891,N_2734,N_2619);
nand U2892 (N_2892,N_2777,N_2662);
and U2893 (N_2893,N_2617,N_2739);
and U2894 (N_2894,N_2713,N_2666);
or U2895 (N_2895,N_2647,N_2790);
or U2896 (N_2896,N_2786,N_2737);
and U2897 (N_2897,N_2631,N_2699);
and U2898 (N_2898,N_2789,N_2645);
or U2899 (N_2899,N_2606,N_2710);
and U2900 (N_2900,N_2619,N_2750);
and U2901 (N_2901,N_2766,N_2757);
or U2902 (N_2902,N_2719,N_2641);
xor U2903 (N_2903,N_2708,N_2681);
nor U2904 (N_2904,N_2771,N_2770);
or U2905 (N_2905,N_2783,N_2622);
or U2906 (N_2906,N_2749,N_2742);
or U2907 (N_2907,N_2713,N_2752);
and U2908 (N_2908,N_2774,N_2668);
xnor U2909 (N_2909,N_2600,N_2602);
and U2910 (N_2910,N_2728,N_2714);
nand U2911 (N_2911,N_2701,N_2731);
nand U2912 (N_2912,N_2603,N_2662);
nand U2913 (N_2913,N_2714,N_2618);
xor U2914 (N_2914,N_2617,N_2781);
and U2915 (N_2915,N_2654,N_2620);
nor U2916 (N_2916,N_2624,N_2783);
or U2917 (N_2917,N_2710,N_2727);
nor U2918 (N_2918,N_2639,N_2748);
or U2919 (N_2919,N_2732,N_2612);
and U2920 (N_2920,N_2601,N_2624);
xnor U2921 (N_2921,N_2645,N_2674);
nor U2922 (N_2922,N_2748,N_2757);
and U2923 (N_2923,N_2708,N_2612);
nand U2924 (N_2924,N_2717,N_2751);
and U2925 (N_2925,N_2755,N_2680);
and U2926 (N_2926,N_2731,N_2657);
xor U2927 (N_2927,N_2779,N_2711);
nor U2928 (N_2928,N_2768,N_2661);
xor U2929 (N_2929,N_2654,N_2605);
and U2930 (N_2930,N_2703,N_2772);
nand U2931 (N_2931,N_2758,N_2761);
nor U2932 (N_2932,N_2779,N_2760);
nor U2933 (N_2933,N_2744,N_2786);
xor U2934 (N_2934,N_2718,N_2623);
and U2935 (N_2935,N_2716,N_2733);
nand U2936 (N_2936,N_2680,N_2664);
xnor U2937 (N_2937,N_2753,N_2773);
xnor U2938 (N_2938,N_2692,N_2687);
or U2939 (N_2939,N_2669,N_2691);
nand U2940 (N_2940,N_2723,N_2601);
and U2941 (N_2941,N_2728,N_2735);
nand U2942 (N_2942,N_2618,N_2747);
nand U2943 (N_2943,N_2744,N_2672);
or U2944 (N_2944,N_2694,N_2689);
xor U2945 (N_2945,N_2754,N_2638);
or U2946 (N_2946,N_2788,N_2628);
and U2947 (N_2947,N_2617,N_2740);
nand U2948 (N_2948,N_2772,N_2651);
or U2949 (N_2949,N_2705,N_2706);
xor U2950 (N_2950,N_2615,N_2737);
nor U2951 (N_2951,N_2796,N_2643);
nor U2952 (N_2952,N_2729,N_2628);
nand U2953 (N_2953,N_2675,N_2742);
xnor U2954 (N_2954,N_2789,N_2673);
or U2955 (N_2955,N_2735,N_2672);
or U2956 (N_2956,N_2600,N_2720);
and U2957 (N_2957,N_2720,N_2631);
nand U2958 (N_2958,N_2757,N_2651);
nor U2959 (N_2959,N_2733,N_2718);
and U2960 (N_2960,N_2679,N_2771);
or U2961 (N_2961,N_2667,N_2793);
and U2962 (N_2962,N_2748,N_2630);
nor U2963 (N_2963,N_2619,N_2606);
nand U2964 (N_2964,N_2610,N_2773);
or U2965 (N_2965,N_2613,N_2628);
nor U2966 (N_2966,N_2657,N_2750);
nand U2967 (N_2967,N_2711,N_2794);
nor U2968 (N_2968,N_2734,N_2683);
and U2969 (N_2969,N_2658,N_2671);
nand U2970 (N_2970,N_2667,N_2733);
and U2971 (N_2971,N_2613,N_2797);
xor U2972 (N_2972,N_2757,N_2698);
or U2973 (N_2973,N_2717,N_2609);
or U2974 (N_2974,N_2678,N_2741);
nor U2975 (N_2975,N_2682,N_2790);
nor U2976 (N_2976,N_2750,N_2760);
or U2977 (N_2977,N_2737,N_2629);
nor U2978 (N_2978,N_2757,N_2704);
nor U2979 (N_2979,N_2628,N_2775);
and U2980 (N_2980,N_2733,N_2754);
xnor U2981 (N_2981,N_2692,N_2649);
or U2982 (N_2982,N_2790,N_2659);
and U2983 (N_2983,N_2668,N_2780);
nor U2984 (N_2984,N_2731,N_2665);
xnor U2985 (N_2985,N_2701,N_2770);
or U2986 (N_2986,N_2769,N_2710);
and U2987 (N_2987,N_2652,N_2690);
nand U2988 (N_2988,N_2688,N_2604);
nand U2989 (N_2989,N_2660,N_2672);
nor U2990 (N_2990,N_2786,N_2713);
or U2991 (N_2991,N_2716,N_2723);
and U2992 (N_2992,N_2699,N_2643);
nand U2993 (N_2993,N_2731,N_2649);
or U2994 (N_2994,N_2618,N_2665);
nor U2995 (N_2995,N_2708,N_2679);
or U2996 (N_2996,N_2641,N_2648);
or U2997 (N_2997,N_2768,N_2610);
or U2998 (N_2998,N_2749,N_2672);
xnor U2999 (N_2999,N_2703,N_2635);
xnor U3000 (N_3000,N_2805,N_2806);
and U3001 (N_3001,N_2931,N_2829);
or U3002 (N_3002,N_2967,N_2828);
or U3003 (N_3003,N_2856,N_2843);
and U3004 (N_3004,N_2968,N_2825);
xor U3005 (N_3005,N_2980,N_2820);
nand U3006 (N_3006,N_2916,N_2917);
xor U3007 (N_3007,N_2874,N_2901);
or U3008 (N_3008,N_2869,N_2817);
nand U3009 (N_3009,N_2850,N_2994);
and U3010 (N_3010,N_2849,N_2953);
nand U3011 (N_3011,N_2937,N_2888);
nand U3012 (N_3012,N_2986,N_2816);
and U3013 (N_3013,N_2815,N_2819);
nand U3014 (N_3014,N_2894,N_2873);
nand U3015 (N_3015,N_2866,N_2952);
nor U3016 (N_3016,N_2867,N_2990);
and U3017 (N_3017,N_2954,N_2960);
nor U3018 (N_3018,N_2851,N_2826);
nor U3019 (N_3019,N_2886,N_2876);
or U3020 (N_3020,N_2922,N_2938);
or U3021 (N_3021,N_2951,N_2904);
nand U3022 (N_3022,N_2844,N_2814);
and U3023 (N_3023,N_2963,N_2924);
or U3024 (N_3024,N_2955,N_2810);
nand U3025 (N_3025,N_2884,N_2897);
and U3026 (N_3026,N_2800,N_2944);
and U3027 (N_3027,N_2847,N_2863);
or U3028 (N_3028,N_2895,N_2973);
nand U3029 (N_3029,N_2977,N_2852);
or U3030 (N_3030,N_2985,N_2911);
nor U3031 (N_3031,N_2949,N_2958);
nor U3032 (N_3032,N_2885,N_2975);
xor U3033 (N_3033,N_2982,N_2839);
and U3034 (N_3034,N_2969,N_2930);
nand U3035 (N_3035,N_2920,N_2932);
nand U3036 (N_3036,N_2864,N_2902);
and U3037 (N_3037,N_2971,N_2890);
nor U3038 (N_3038,N_2919,N_2976);
or U3039 (N_3039,N_2933,N_2870);
nor U3040 (N_3040,N_2972,N_2837);
nor U3041 (N_3041,N_2891,N_2841);
or U3042 (N_3042,N_2823,N_2908);
nand U3043 (N_3043,N_2812,N_2912);
xnor U3044 (N_3044,N_2992,N_2946);
and U3045 (N_3045,N_2991,N_2981);
nor U3046 (N_3046,N_2809,N_2927);
and U3047 (N_3047,N_2880,N_2898);
or U3048 (N_3048,N_2860,N_2840);
or U3049 (N_3049,N_2956,N_2983);
xor U3050 (N_3050,N_2813,N_2964);
or U3051 (N_3051,N_2935,N_2872);
nor U3052 (N_3052,N_2896,N_2878);
nand U3053 (N_3053,N_2934,N_2906);
nor U3054 (N_3054,N_2855,N_2965);
nor U3055 (N_3055,N_2893,N_2865);
xor U3056 (N_3056,N_2995,N_2974);
and U3057 (N_3057,N_2803,N_2808);
or U3058 (N_3058,N_2868,N_2905);
or U3059 (N_3059,N_2802,N_2907);
nor U3060 (N_3060,N_2950,N_2943);
nand U3061 (N_3061,N_2900,N_2853);
xor U3062 (N_3062,N_2899,N_2970);
or U3063 (N_3063,N_2848,N_2989);
xor U3064 (N_3064,N_2961,N_2801);
nand U3065 (N_3065,N_2807,N_2914);
nand U3066 (N_3066,N_2928,N_2940);
nand U3067 (N_3067,N_2913,N_2879);
or U3068 (N_3068,N_2861,N_2832);
nor U3069 (N_3069,N_2835,N_2988);
and U3070 (N_3070,N_2925,N_2877);
nor U3071 (N_3071,N_2836,N_2921);
nand U3072 (N_3072,N_2993,N_2910);
xnor U3073 (N_3073,N_2824,N_2957);
or U3074 (N_3074,N_2915,N_2833);
nor U3075 (N_3075,N_2831,N_2947);
xor U3076 (N_3076,N_2822,N_2942);
nor U3077 (N_3077,N_2984,N_2811);
xnor U3078 (N_3078,N_2834,N_2827);
nand U3079 (N_3079,N_2858,N_2939);
and U3080 (N_3080,N_2842,N_2909);
nand U3081 (N_3081,N_2918,N_2821);
and U3082 (N_3082,N_2998,N_2857);
nor U3083 (N_3083,N_2959,N_2845);
or U3084 (N_3084,N_2941,N_2881);
or U3085 (N_3085,N_2987,N_2887);
nor U3086 (N_3086,N_2996,N_2892);
or U3087 (N_3087,N_2923,N_2830);
or U3088 (N_3088,N_2838,N_2979);
or U3089 (N_3089,N_2945,N_2818);
and U3090 (N_3090,N_2862,N_2882);
xor U3091 (N_3091,N_2978,N_2948);
nand U3092 (N_3092,N_2962,N_2903);
and U3093 (N_3093,N_2883,N_2871);
nor U3094 (N_3094,N_2804,N_2859);
nand U3095 (N_3095,N_2936,N_2875);
nand U3096 (N_3096,N_2929,N_2889);
or U3097 (N_3097,N_2997,N_2846);
xnor U3098 (N_3098,N_2999,N_2966);
nor U3099 (N_3099,N_2926,N_2854);
xor U3100 (N_3100,N_2937,N_2822);
xnor U3101 (N_3101,N_2906,N_2850);
and U3102 (N_3102,N_2982,N_2843);
nand U3103 (N_3103,N_2943,N_2807);
xor U3104 (N_3104,N_2851,N_2968);
and U3105 (N_3105,N_2825,N_2897);
nand U3106 (N_3106,N_2894,N_2905);
and U3107 (N_3107,N_2856,N_2882);
xor U3108 (N_3108,N_2974,N_2989);
and U3109 (N_3109,N_2898,N_2806);
xor U3110 (N_3110,N_2811,N_2919);
and U3111 (N_3111,N_2828,N_2884);
or U3112 (N_3112,N_2804,N_2942);
nand U3113 (N_3113,N_2861,N_2924);
xor U3114 (N_3114,N_2992,N_2834);
xor U3115 (N_3115,N_2947,N_2916);
xnor U3116 (N_3116,N_2907,N_2906);
nor U3117 (N_3117,N_2980,N_2879);
or U3118 (N_3118,N_2944,N_2881);
and U3119 (N_3119,N_2824,N_2928);
and U3120 (N_3120,N_2814,N_2932);
nor U3121 (N_3121,N_2846,N_2837);
and U3122 (N_3122,N_2877,N_2965);
nand U3123 (N_3123,N_2811,N_2875);
and U3124 (N_3124,N_2909,N_2848);
xor U3125 (N_3125,N_2854,N_2810);
nand U3126 (N_3126,N_2828,N_2988);
nor U3127 (N_3127,N_2971,N_2893);
and U3128 (N_3128,N_2893,N_2958);
nor U3129 (N_3129,N_2946,N_2822);
nand U3130 (N_3130,N_2989,N_2898);
and U3131 (N_3131,N_2928,N_2860);
xnor U3132 (N_3132,N_2912,N_2995);
nor U3133 (N_3133,N_2986,N_2847);
xnor U3134 (N_3134,N_2813,N_2853);
and U3135 (N_3135,N_2942,N_2803);
xor U3136 (N_3136,N_2964,N_2877);
and U3137 (N_3137,N_2949,N_2893);
or U3138 (N_3138,N_2847,N_2942);
nor U3139 (N_3139,N_2956,N_2848);
nor U3140 (N_3140,N_2872,N_2918);
nor U3141 (N_3141,N_2929,N_2850);
nand U3142 (N_3142,N_2824,N_2878);
nor U3143 (N_3143,N_2809,N_2916);
and U3144 (N_3144,N_2850,N_2844);
nand U3145 (N_3145,N_2851,N_2876);
nor U3146 (N_3146,N_2884,N_2949);
nand U3147 (N_3147,N_2912,N_2996);
nand U3148 (N_3148,N_2892,N_2861);
xor U3149 (N_3149,N_2886,N_2990);
or U3150 (N_3150,N_2910,N_2850);
nand U3151 (N_3151,N_2823,N_2994);
or U3152 (N_3152,N_2927,N_2825);
xor U3153 (N_3153,N_2870,N_2835);
or U3154 (N_3154,N_2879,N_2807);
or U3155 (N_3155,N_2989,N_2918);
xor U3156 (N_3156,N_2974,N_2896);
xnor U3157 (N_3157,N_2900,N_2939);
or U3158 (N_3158,N_2837,N_2827);
or U3159 (N_3159,N_2964,N_2840);
and U3160 (N_3160,N_2916,N_2999);
and U3161 (N_3161,N_2940,N_2937);
nand U3162 (N_3162,N_2971,N_2977);
xor U3163 (N_3163,N_2868,N_2931);
or U3164 (N_3164,N_2946,N_2845);
and U3165 (N_3165,N_2808,N_2982);
xor U3166 (N_3166,N_2961,N_2842);
nand U3167 (N_3167,N_2971,N_2883);
or U3168 (N_3168,N_2929,N_2991);
nand U3169 (N_3169,N_2926,N_2928);
or U3170 (N_3170,N_2985,N_2922);
nand U3171 (N_3171,N_2834,N_2996);
or U3172 (N_3172,N_2819,N_2952);
xor U3173 (N_3173,N_2875,N_2937);
nor U3174 (N_3174,N_2842,N_2959);
or U3175 (N_3175,N_2944,N_2928);
or U3176 (N_3176,N_2852,N_2855);
or U3177 (N_3177,N_2931,N_2844);
or U3178 (N_3178,N_2991,N_2885);
nand U3179 (N_3179,N_2880,N_2946);
nand U3180 (N_3180,N_2862,N_2936);
and U3181 (N_3181,N_2879,N_2956);
nand U3182 (N_3182,N_2936,N_2866);
xnor U3183 (N_3183,N_2939,N_2888);
nor U3184 (N_3184,N_2984,N_2823);
and U3185 (N_3185,N_2835,N_2974);
nand U3186 (N_3186,N_2844,N_2997);
xor U3187 (N_3187,N_2851,N_2855);
nand U3188 (N_3188,N_2884,N_2899);
nand U3189 (N_3189,N_2881,N_2935);
and U3190 (N_3190,N_2962,N_2997);
nand U3191 (N_3191,N_2819,N_2847);
nor U3192 (N_3192,N_2928,N_2933);
nand U3193 (N_3193,N_2969,N_2909);
and U3194 (N_3194,N_2915,N_2824);
or U3195 (N_3195,N_2871,N_2831);
xnor U3196 (N_3196,N_2812,N_2918);
xnor U3197 (N_3197,N_2983,N_2826);
or U3198 (N_3198,N_2929,N_2843);
xnor U3199 (N_3199,N_2969,N_2985);
nand U3200 (N_3200,N_3187,N_3186);
nand U3201 (N_3201,N_3057,N_3061);
nand U3202 (N_3202,N_3091,N_3063);
and U3203 (N_3203,N_3021,N_3039);
nor U3204 (N_3204,N_3084,N_3006);
nor U3205 (N_3205,N_3035,N_3075);
nand U3206 (N_3206,N_3157,N_3151);
and U3207 (N_3207,N_3053,N_3133);
nand U3208 (N_3208,N_3002,N_3031);
nand U3209 (N_3209,N_3183,N_3062);
xor U3210 (N_3210,N_3016,N_3081);
nand U3211 (N_3211,N_3092,N_3199);
and U3212 (N_3212,N_3146,N_3041);
nor U3213 (N_3213,N_3123,N_3104);
nor U3214 (N_3214,N_3124,N_3093);
or U3215 (N_3215,N_3015,N_3182);
and U3216 (N_3216,N_3070,N_3072);
and U3217 (N_3217,N_3162,N_3149);
nand U3218 (N_3218,N_3000,N_3013);
xnor U3219 (N_3219,N_3109,N_3197);
nand U3220 (N_3220,N_3167,N_3164);
or U3221 (N_3221,N_3023,N_3101);
xor U3222 (N_3222,N_3178,N_3115);
xnor U3223 (N_3223,N_3058,N_3087);
xnor U3224 (N_3224,N_3011,N_3168);
and U3225 (N_3225,N_3066,N_3034);
xor U3226 (N_3226,N_3026,N_3064);
nand U3227 (N_3227,N_3079,N_3147);
and U3228 (N_3228,N_3154,N_3136);
and U3229 (N_3229,N_3180,N_3014);
nand U3230 (N_3230,N_3055,N_3119);
and U3231 (N_3231,N_3161,N_3176);
and U3232 (N_3232,N_3172,N_3027);
nand U3233 (N_3233,N_3043,N_3001);
xnor U3234 (N_3234,N_3165,N_3148);
xor U3235 (N_3235,N_3193,N_3159);
nor U3236 (N_3236,N_3122,N_3113);
nor U3237 (N_3237,N_3007,N_3105);
and U3238 (N_3238,N_3129,N_3181);
nor U3239 (N_3239,N_3071,N_3096);
and U3240 (N_3240,N_3155,N_3012);
nor U3241 (N_3241,N_3005,N_3078);
nor U3242 (N_3242,N_3077,N_3028);
xnor U3243 (N_3243,N_3128,N_3040);
or U3244 (N_3244,N_3117,N_3019);
nor U3245 (N_3245,N_3152,N_3125);
or U3246 (N_3246,N_3051,N_3138);
and U3247 (N_3247,N_3049,N_3107);
nor U3248 (N_3248,N_3065,N_3140);
nand U3249 (N_3249,N_3116,N_3150);
nand U3250 (N_3250,N_3085,N_3024);
nand U3251 (N_3251,N_3097,N_3111);
xor U3252 (N_3252,N_3095,N_3010);
xnor U3253 (N_3253,N_3196,N_3139);
and U3254 (N_3254,N_3134,N_3025);
nand U3255 (N_3255,N_3184,N_3068);
nor U3256 (N_3256,N_3131,N_3163);
nor U3257 (N_3257,N_3177,N_3191);
nor U3258 (N_3258,N_3089,N_3083);
and U3259 (N_3259,N_3108,N_3179);
or U3260 (N_3260,N_3106,N_3100);
xnor U3261 (N_3261,N_3144,N_3073);
or U3262 (N_3262,N_3174,N_3158);
nand U3263 (N_3263,N_3003,N_3036);
nand U3264 (N_3264,N_3120,N_3132);
and U3265 (N_3265,N_3050,N_3088);
and U3266 (N_3266,N_3094,N_3098);
or U3267 (N_3267,N_3195,N_3082);
nor U3268 (N_3268,N_3038,N_3190);
xor U3269 (N_3269,N_3112,N_3074);
or U3270 (N_3270,N_3047,N_3194);
nor U3271 (N_3271,N_3032,N_3052);
nand U3272 (N_3272,N_3102,N_3048);
or U3273 (N_3273,N_3029,N_3046);
nor U3274 (N_3274,N_3110,N_3009);
xnor U3275 (N_3275,N_3017,N_3114);
and U3276 (N_3276,N_3118,N_3188);
or U3277 (N_3277,N_3054,N_3018);
nor U3278 (N_3278,N_3160,N_3126);
nor U3279 (N_3279,N_3137,N_3059);
or U3280 (N_3280,N_3135,N_3080);
xor U3281 (N_3281,N_3060,N_3030);
and U3282 (N_3282,N_3069,N_3130);
nand U3283 (N_3283,N_3004,N_3103);
nand U3284 (N_3284,N_3045,N_3173);
xor U3285 (N_3285,N_3042,N_3169);
and U3286 (N_3286,N_3022,N_3008);
xnor U3287 (N_3287,N_3076,N_3067);
and U3288 (N_3288,N_3189,N_3156);
and U3289 (N_3289,N_3143,N_3141);
and U3290 (N_3290,N_3086,N_3127);
xnor U3291 (N_3291,N_3170,N_3033);
or U3292 (N_3292,N_3171,N_3153);
nand U3293 (N_3293,N_3056,N_3185);
xnor U3294 (N_3294,N_3020,N_3037);
or U3295 (N_3295,N_3175,N_3090);
and U3296 (N_3296,N_3166,N_3099);
nor U3297 (N_3297,N_3044,N_3192);
or U3298 (N_3298,N_3198,N_3142);
and U3299 (N_3299,N_3145,N_3121);
nand U3300 (N_3300,N_3135,N_3169);
and U3301 (N_3301,N_3100,N_3062);
nor U3302 (N_3302,N_3147,N_3080);
xor U3303 (N_3303,N_3073,N_3007);
or U3304 (N_3304,N_3136,N_3066);
xnor U3305 (N_3305,N_3182,N_3044);
or U3306 (N_3306,N_3113,N_3187);
nor U3307 (N_3307,N_3174,N_3147);
nand U3308 (N_3308,N_3167,N_3120);
nor U3309 (N_3309,N_3070,N_3098);
xnor U3310 (N_3310,N_3138,N_3164);
and U3311 (N_3311,N_3175,N_3102);
nor U3312 (N_3312,N_3146,N_3171);
nand U3313 (N_3313,N_3056,N_3188);
xnor U3314 (N_3314,N_3191,N_3150);
nand U3315 (N_3315,N_3060,N_3187);
and U3316 (N_3316,N_3066,N_3048);
or U3317 (N_3317,N_3030,N_3185);
xor U3318 (N_3318,N_3031,N_3147);
nor U3319 (N_3319,N_3086,N_3073);
or U3320 (N_3320,N_3121,N_3177);
nand U3321 (N_3321,N_3134,N_3045);
nor U3322 (N_3322,N_3099,N_3110);
or U3323 (N_3323,N_3144,N_3197);
nand U3324 (N_3324,N_3095,N_3108);
and U3325 (N_3325,N_3149,N_3009);
and U3326 (N_3326,N_3105,N_3146);
xnor U3327 (N_3327,N_3173,N_3011);
xnor U3328 (N_3328,N_3147,N_3197);
nand U3329 (N_3329,N_3010,N_3081);
and U3330 (N_3330,N_3015,N_3162);
or U3331 (N_3331,N_3064,N_3014);
nor U3332 (N_3332,N_3136,N_3021);
nand U3333 (N_3333,N_3145,N_3036);
nand U3334 (N_3334,N_3196,N_3076);
nor U3335 (N_3335,N_3104,N_3155);
and U3336 (N_3336,N_3092,N_3036);
and U3337 (N_3337,N_3088,N_3002);
or U3338 (N_3338,N_3141,N_3001);
or U3339 (N_3339,N_3150,N_3134);
nor U3340 (N_3340,N_3156,N_3103);
xor U3341 (N_3341,N_3153,N_3091);
xor U3342 (N_3342,N_3087,N_3109);
xnor U3343 (N_3343,N_3003,N_3004);
nand U3344 (N_3344,N_3184,N_3188);
xor U3345 (N_3345,N_3088,N_3137);
nor U3346 (N_3346,N_3147,N_3170);
xnor U3347 (N_3347,N_3194,N_3110);
nand U3348 (N_3348,N_3183,N_3175);
or U3349 (N_3349,N_3056,N_3076);
nor U3350 (N_3350,N_3084,N_3025);
xnor U3351 (N_3351,N_3095,N_3085);
nand U3352 (N_3352,N_3051,N_3112);
nor U3353 (N_3353,N_3032,N_3022);
and U3354 (N_3354,N_3186,N_3034);
or U3355 (N_3355,N_3171,N_3106);
nor U3356 (N_3356,N_3093,N_3064);
nor U3357 (N_3357,N_3140,N_3047);
or U3358 (N_3358,N_3096,N_3014);
nand U3359 (N_3359,N_3128,N_3101);
nand U3360 (N_3360,N_3004,N_3173);
or U3361 (N_3361,N_3114,N_3048);
xnor U3362 (N_3362,N_3168,N_3020);
nor U3363 (N_3363,N_3013,N_3093);
or U3364 (N_3364,N_3179,N_3128);
nand U3365 (N_3365,N_3103,N_3187);
nand U3366 (N_3366,N_3004,N_3186);
nor U3367 (N_3367,N_3051,N_3077);
nor U3368 (N_3368,N_3027,N_3150);
or U3369 (N_3369,N_3072,N_3163);
and U3370 (N_3370,N_3111,N_3033);
or U3371 (N_3371,N_3020,N_3153);
and U3372 (N_3372,N_3071,N_3117);
xnor U3373 (N_3373,N_3125,N_3132);
or U3374 (N_3374,N_3153,N_3191);
and U3375 (N_3375,N_3007,N_3078);
xor U3376 (N_3376,N_3150,N_3144);
nand U3377 (N_3377,N_3188,N_3018);
and U3378 (N_3378,N_3079,N_3062);
or U3379 (N_3379,N_3189,N_3143);
xnor U3380 (N_3380,N_3144,N_3007);
nor U3381 (N_3381,N_3070,N_3152);
xor U3382 (N_3382,N_3179,N_3187);
and U3383 (N_3383,N_3025,N_3142);
and U3384 (N_3384,N_3065,N_3146);
and U3385 (N_3385,N_3027,N_3154);
or U3386 (N_3386,N_3155,N_3022);
nand U3387 (N_3387,N_3045,N_3146);
or U3388 (N_3388,N_3049,N_3157);
nand U3389 (N_3389,N_3089,N_3179);
and U3390 (N_3390,N_3157,N_3104);
or U3391 (N_3391,N_3073,N_3166);
xnor U3392 (N_3392,N_3096,N_3010);
nor U3393 (N_3393,N_3087,N_3199);
nor U3394 (N_3394,N_3099,N_3019);
xnor U3395 (N_3395,N_3115,N_3150);
nor U3396 (N_3396,N_3019,N_3151);
nor U3397 (N_3397,N_3172,N_3112);
or U3398 (N_3398,N_3179,N_3159);
or U3399 (N_3399,N_3095,N_3189);
nor U3400 (N_3400,N_3293,N_3355);
nor U3401 (N_3401,N_3350,N_3323);
and U3402 (N_3402,N_3375,N_3295);
nor U3403 (N_3403,N_3238,N_3271);
and U3404 (N_3404,N_3363,N_3342);
and U3405 (N_3405,N_3376,N_3397);
and U3406 (N_3406,N_3287,N_3211);
and U3407 (N_3407,N_3386,N_3345);
xor U3408 (N_3408,N_3255,N_3389);
xor U3409 (N_3409,N_3262,N_3292);
or U3410 (N_3410,N_3398,N_3387);
or U3411 (N_3411,N_3388,N_3351);
or U3412 (N_3412,N_3365,N_3276);
xnor U3413 (N_3413,N_3311,N_3231);
and U3414 (N_3414,N_3368,N_3250);
or U3415 (N_3415,N_3235,N_3393);
nor U3416 (N_3416,N_3358,N_3296);
nor U3417 (N_3417,N_3348,N_3337);
nor U3418 (N_3418,N_3294,N_3267);
or U3419 (N_3419,N_3246,N_3298);
nand U3420 (N_3420,N_3317,N_3218);
xor U3421 (N_3421,N_3214,N_3391);
or U3422 (N_3422,N_3320,N_3374);
nand U3423 (N_3423,N_3257,N_3390);
nor U3424 (N_3424,N_3304,N_3366);
or U3425 (N_3425,N_3349,N_3283);
nand U3426 (N_3426,N_3249,N_3200);
nor U3427 (N_3427,N_3381,N_3360);
or U3428 (N_3428,N_3297,N_3209);
nor U3429 (N_3429,N_3256,N_3384);
nor U3430 (N_3430,N_3290,N_3318);
xnor U3431 (N_3431,N_3341,N_3321);
or U3432 (N_3432,N_3313,N_3286);
or U3433 (N_3433,N_3383,N_3336);
xor U3434 (N_3434,N_3291,N_3319);
and U3435 (N_3435,N_3237,N_3264);
nand U3436 (N_3436,N_3356,N_3334);
or U3437 (N_3437,N_3309,N_3308);
or U3438 (N_3438,N_3251,N_3208);
nor U3439 (N_3439,N_3312,N_3316);
and U3440 (N_3440,N_3277,N_3288);
nand U3441 (N_3441,N_3346,N_3343);
nor U3442 (N_3442,N_3282,N_3289);
and U3443 (N_3443,N_3201,N_3325);
or U3444 (N_3444,N_3362,N_3221);
xnor U3445 (N_3445,N_3258,N_3329);
nor U3446 (N_3446,N_3307,N_3219);
nor U3447 (N_3447,N_3330,N_3380);
or U3448 (N_3448,N_3263,N_3217);
or U3449 (N_3449,N_3284,N_3212);
nor U3450 (N_3450,N_3314,N_3332);
nor U3451 (N_3451,N_3326,N_3339);
and U3452 (N_3452,N_3315,N_3373);
nor U3453 (N_3453,N_3242,N_3302);
and U3454 (N_3454,N_3204,N_3222);
and U3455 (N_3455,N_3370,N_3364);
or U3456 (N_3456,N_3385,N_3279);
or U3457 (N_3457,N_3310,N_3202);
and U3458 (N_3458,N_3253,N_3228);
xor U3459 (N_3459,N_3241,N_3361);
nand U3460 (N_3460,N_3252,N_3275);
xor U3461 (N_3461,N_3239,N_3223);
or U3462 (N_3462,N_3327,N_3224);
xnor U3463 (N_3463,N_3396,N_3216);
nor U3464 (N_3464,N_3331,N_3372);
nand U3465 (N_3465,N_3322,N_3248);
and U3466 (N_3466,N_3301,N_3203);
or U3467 (N_3467,N_3254,N_3280);
nand U3468 (N_3468,N_3395,N_3369);
nor U3469 (N_3469,N_3382,N_3399);
nand U3470 (N_3470,N_3357,N_3265);
nand U3471 (N_3471,N_3226,N_3300);
and U3472 (N_3472,N_3371,N_3394);
nand U3473 (N_3473,N_3340,N_3303);
nand U3474 (N_3474,N_3260,N_3227);
xnor U3475 (N_3475,N_3230,N_3229);
xor U3476 (N_3476,N_3205,N_3367);
or U3477 (N_3477,N_3285,N_3359);
and U3478 (N_3478,N_3234,N_3215);
nor U3479 (N_3479,N_3353,N_3392);
xor U3480 (N_3480,N_3225,N_3273);
nand U3481 (N_3481,N_3379,N_3324);
and U3482 (N_3482,N_3281,N_3210);
or U3483 (N_3483,N_3240,N_3207);
nand U3484 (N_3484,N_3266,N_3377);
and U3485 (N_3485,N_3344,N_3244);
and U3486 (N_3486,N_3268,N_3245);
nor U3487 (N_3487,N_3378,N_3232);
nand U3488 (N_3488,N_3243,N_3306);
nand U3489 (N_3489,N_3272,N_3347);
and U3490 (N_3490,N_3354,N_3206);
and U3491 (N_3491,N_3278,N_3259);
nor U3492 (N_3492,N_3299,N_3220);
nand U3493 (N_3493,N_3335,N_3269);
or U3494 (N_3494,N_3236,N_3328);
or U3495 (N_3495,N_3338,N_3274);
nor U3496 (N_3496,N_3247,N_3333);
nor U3497 (N_3497,N_3213,N_3261);
or U3498 (N_3498,N_3270,N_3352);
nand U3499 (N_3499,N_3233,N_3305);
nand U3500 (N_3500,N_3398,N_3245);
nand U3501 (N_3501,N_3307,N_3318);
and U3502 (N_3502,N_3382,N_3393);
or U3503 (N_3503,N_3283,N_3319);
xnor U3504 (N_3504,N_3381,N_3339);
nor U3505 (N_3505,N_3277,N_3266);
and U3506 (N_3506,N_3366,N_3219);
xnor U3507 (N_3507,N_3390,N_3252);
nand U3508 (N_3508,N_3276,N_3395);
nor U3509 (N_3509,N_3231,N_3259);
nor U3510 (N_3510,N_3241,N_3284);
or U3511 (N_3511,N_3380,N_3366);
nand U3512 (N_3512,N_3304,N_3280);
nor U3513 (N_3513,N_3223,N_3306);
or U3514 (N_3514,N_3248,N_3216);
nand U3515 (N_3515,N_3315,N_3389);
nor U3516 (N_3516,N_3326,N_3329);
xor U3517 (N_3517,N_3326,N_3286);
xnor U3518 (N_3518,N_3264,N_3219);
nand U3519 (N_3519,N_3268,N_3223);
xor U3520 (N_3520,N_3320,N_3244);
or U3521 (N_3521,N_3205,N_3397);
and U3522 (N_3522,N_3358,N_3355);
xnor U3523 (N_3523,N_3203,N_3378);
or U3524 (N_3524,N_3210,N_3329);
nand U3525 (N_3525,N_3205,N_3308);
nor U3526 (N_3526,N_3372,N_3249);
nor U3527 (N_3527,N_3398,N_3399);
nor U3528 (N_3528,N_3206,N_3392);
xnor U3529 (N_3529,N_3246,N_3279);
xnor U3530 (N_3530,N_3259,N_3212);
or U3531 (N_3531,N_3381,N_3390);
xnor U3532 (N_3532,N_3239,N_3231);
and U3533 (N_3533,N_3264,N_3352);
or U3534 (N_3534,N_3337,N_3252);
or U3535 (N_3535,N_3299,N_3295);
nor U3536 (N_3536,N_3282,N_3226);
nand U3537 (N_3537,N_3334,N_3382);
nand U3538 (N_3538,N_3267,N_3306);
and U3539 (N_3539,N_3338,N_3318);
and U3540 (N_3540,N_3292,N_3224);
xor U3541 (N_3541,N_3346,N_3326);
xor U3542 (N_3542,N_3381,N_3283);
nand U3543 (N_3543,N_3325,N_3200);
xnor U3544 (N_3544,N_3395,N_3303);
nand U3545 (N_3545,N_3309,N_3361);
nor U3546 (N_3546,N_3387,N_3322);
xnor U3547 (N_3547,N_3300,N_3318);
and U3548 (N_3548,N_3213,N_3338);
nor U3549 (N_3549,N_3292,N_3321);
nor U3550 (N_3550,N_3221,N_3281);
xor U3551 (N_3551,N_3251,N_3237);
and U3552 (N_3552,N_3340,N_3270);
xnor U3553 (N_3553,N_3376,N_3221);
and U3554 (N_3554,N_3268,N_3269);
and U3555 (N_3555,N_3368,N_3221);
and U3556 (N_3556,N_3228,N_3276);
or U3557 (N_3557,N_3330,N_3373);
xor U3558 (N_3558,N_3277,N_3228);
xor U3559 (N_3559,N_3378,N_3214);
and U3560 (N_3560,N_3273,N_3359);
xor U3561 (N_3561,N_3281,N_3387);
or U3562 (N_3562,N_3240,N_3237);
nor U3563 (N_3563,N_3339,N_3219);
nor U3564 (N_3564,N_3335,N_3292);
or U3565 (N_3565,N_3286,N_3386);
nand U3566 (N_3566,N_3218,N_3299);
nor U3567 (N_3567,N_3353,N_3207);
or U3568 (N_3568,N_3333,N_3338);
nor U3569 (N_3569,N_3337,N_3241);
nor U3570 (N_3570,N_3392,N_3275);
or U3571 (N_3571,N_3254,N_3277);
nand U3572 (N_3572,N_3251,N_3252);
xor U3573 (N_3573,N_3299,N_3319);
xor U3574 (N_3574,N_3278,N_3209);
and U3575 (N_3575,N_3397,N_3341);
nand U3576 (N_3576,N_3222,N_3201);
nor U3577 (N_3577,N_3369,N_3249);
or U3578 (N_3578,N_3395,N_3321);
nand U3579 (N_3579,N_3211,N_3338);
nor U3580 (N_3580,N_3333,N_3224);
or U3581 (N_3581,N_3204,N_3397);
xor U3582 (N_3582,N_3396,N_3381);
or U3583 (N_3583,N_3323,N_3218);
xor U3584 (N_3584,N_3307,N_3209);
nor U3585 (N_3585,N_3279,N_3394);
nor U3586 (N_3586,N_3330,N_3377);
and U3587 (N_3587,N_3394,N_3272);
nor U3588 (N_3588,N_3390,N_3351);
or U3589 (N_3589,N_3217,N_3231);
or U3590 (N_3590,N_3260,N_3337);
xnor U3591 (N_3591,N_3209,N_3328);
nor U3592 (N_3592,N_3232,N_3377);
or U3593 (N_3593,N_3256,N_3207);
and U3594 (N_3594,N_3330,N_3258);
or U3595 (N_3595,N_3295,N_3289);
xor U3596 (N_3596,N_3235,N_3336);
xnor U3597 (N_3597,N_3367,N_3296);
and U3598 (N_3598,N_3274,N_3236);
nand U3599 (N_3599,N_3394,N_3383);
nor U3600 (N_3600,N_3558,N_3596);
xnor U3601 (N_3601,N_3407,N_3590);
and U3602 (N_3602,N_3451,N_3540);
nand U3603 (N_3603,N_3482,N_3573);
or U3604 (N_3604,N_3447,N_3457);
and U3605 (N_3605,N_3585,N_3423);
or U3606 (N_3606,N_3406,N_3592);
and U3607 (N_3607,N_3500,N_3554);
or U3608 (N_3608,N_3545,N_3535);
nor U3609 (N_3609,N_3491,N_3538);
or U3610 (N_3610,N_3452,N_3476);
nand U3611 (N_3611,N_3571,N_3530);
xor U3612 (N_3612,N_3546,N_3487);
nor U3613 (N_3613,N_3485,N_3569);
nor U3614 (N_3614,N_3428,N_3519);
and U3615 (N_3615,N_3562,N_3516);
and U3616 (N_3616,N_3525,N_3414);
xnor U3617 (N_3617,N_3549,N_3479);
nor U3618 (N_3618,N_3495,N_3502);
or U3619 (N_3619,N_3450,N_3578);
or U3620 (N_3620,N_3421,N_3460);
or U3621 (N_3621,N_3597,N_3580);
nor U3622 (N_3622,N_3599,N_3405);
nor U3623 (N_3623,N_3501,N_3449);
xnor U3624 (N_3624,N_3598,N_3470);
nor U3625 (N_3625,N_3453,N_3586);
and U3626 (N_3626,N_3531,N_3413);
and U3627 (N_3627,N_3523,N_3418);
xnor U3628 (N_3628,N_3526,N_3498);
and U3629 (N_3629,N_3567,N_3422);
and U3630 (N_3630,N_3555,N_3572);
nand U3631 (N_3631,N_3468,N_3420);
nor U3632 (N_3632,N_3574,N_3466);
or U3633 (N_3633,N_3544,N_3433);
nor U3634 (N_3634,N_3507,N_3432);
or U3635 (N_3635,N_3489,N_3577);
or U3636 (N_3636,N_3542,N_3575);
and U3637 (N_3637,N_3475,N_3565);
or U3638 (N_3638,N_3529,N_3462);
nor U3639 (N_3639,N_3480,N_3412);
xor U3640 (N_3640,N_3591,N_3430);
nand U3641 (N_3641,N_3439,N_3570);
xnor U3642 (N_3642,N_3589,N_3497);
nor U3643 (N_3643,N_3429,N_3504);
and U3644 (N_3644,N_3513,N_3584);
nand U3645 (N_3645,N_3488,N_3547);
and U3646 (N_3646,N_3438,N_3474);
xor U3647 (N_3647,N_3563,N_3404);
and U3648 (N_3648,N_3403,N_3444);
nor U3649 (N_3649,N_3455,N_3517);
nand U3650 (N_3650,N_3492,N_3566);
and U3651 (N_3651,N_3401,N_3463);
nor U3652 (N_3652,N_3593,N_3582);
and U3653 (N_3653,N_3539,N_3467);
xor U3654 (N_3654,N_3594,N_3494);
nand U3655 (N_3655,N_3541,N_3579);
nand U3656 (N_3656,N_3464,N_3587);
nor U3657 (N_3657,N_3576,N_3459);
nor U3658 (N_3658,N_3508,N_3556);
xnor U3659 (N_3659,N_3561,N_3527);
nor U3660 (N_3660,N_3434,N_3534);
or U3661 (N_3661,N_3499,N_3543);
nor U3662 (N_3662,N_3409,N_3528);
nor U3663 (N_3663,N_3548,N_3581);
nand U3664 (N_3664,N_3445,N_3550);
and U3665 (N_3665,N_3402,N_3496);
nor U3666 (N_3666,N_3552,N_3551);
or U3667 (N_3667,N_3515,N_3559);
nand U3668 (N_3668,N_3419,N_3411);
nor U3669 (N_3669,N_3509,N_3440);
xnor U3670 (N_3670,N_3518,N_3532);
nor U3671 (N_3671,N_3471,N_3533);
or U3672 (N_3672,N_3503,N_3410);
xnor U3673 (N_3673,N_3481,N_3553);
nand U3674 (N_3674,N_3415,N_3416);
nand U3675 (N_3675,N_3537,N_3478);
or U3676 (N_3676,N_3557,N_3469);
and U3677 (N_3677,N_3431,N_3560);
nand U3678 (N_3678,N_3506,N_3595);
xnor U3679 (N_3679,N_3436,N_3521);
or U3680 (N_3680,N_3465,N_3536);
and U3681 (N_3681,N_3417,N_3448);
nand U3682 (N_3682,N_3493,N_3458);
xnor U3683 (N_3683,N_3446,N_3511);
and U3684 (N_3684,N_3424,N_3441);
and U3685 (N_3685,N_3472,N_3588);
xor U3686 (N_3686,N_3426,N_3505);
nor U3687 (N_3687,N_3522,N_3524);
and U3688 (N_3688,N_3490,N_3484);
or U3689 (N_3689,N_3477,N_3456);
or U3690 (N_3690,N_3443,N_3483);
and U3691 (N_3691,N_3514,N_3583);
and U3692 (N_3692,N_3408,N_3512);
nor U3693 (N_3693,N_3454,N_3486);
or U3694 (N_3694,N_3425,N_3564);
nand U3695 (N_3695,N_3461,N_3442);
xor U3696 (N_3696,N_3437,N_3510);
xnor U3697 (N_3697,N_3427,N_3473);
xor U3698 (N_3698,N_3568,N_3520);
and U3699 (N_3699,N_3435,N_3400);
or U3700 (N_3700,N_3421,N_3440);
nand U3701 (N_3701,N_3410,N_3544);
or U3702 (N_3702,N_3446,N_3525);
nor U3703 (N_3703,N_3596,N_3406);
nand U3704 (N_3704,N_3518,N_3470);
xnor U3705 (N_3705,N_3574,N_3478);
and U3706 (N_3706,N_3473,N_3537);
and U3707 (N_3707,N_3452,N_3506);
nand U3708 (N_3708,N_3593,N_3437);
xor U3709 (N_3709,N_3441,N_3547);
or U3710 (N_3710,N_3558,N_3497);
xor U3711 (N_3711,N_3503,N_3587);
and U3712 (N_3712,N_3578,N_3517);
or U3713 (N_3713,N_3597,N_3533);
and U3714 (N_3714,N_3556,N_3402);
xnor U3715 (N_3715,N_3444,N_3499);
or U3716 (N_3716,N_3401,N_3596);
and U3717 (N_3717,N_3574,N_3522);
xnor U3718 (N_3718,N_3479,N_3444);
nand U3719 (N_3719,N_3582,N_3568);
nand U3720 (N_3720,N_3477,N_3497);
or U3721 (N_3721,N_3519,N_3568);
or U3722 (N_3722,N_3590,N_3573);
nor U3723 (N_3723,N_3416,N_3571);
nor U3724 (N_3724,N_3425,N_3411);
nor U3725 (N_3725,N_3554,N_3410);
nand U3726 (N_3726,N_3493,N_3446);
xnor U3727 (N_3727,N_3559,N_3493);
or U3728 (N_3728,N_3540,N_3563);
nor U3729 (N_3729,N_3487,N_3557);
or U3730 (N_3730,N_3537,N_3543);
and U3731 (N_3731,N_3425,N_3417);
xor U3732 (N_3732,N_3429,N_3489);
xor U3733 (N_3733,N_3545,N_3439);
xnor U3734 (N_3734,N_3405,N_3593);
or U3735 (N_3735,N_3431,N_3569);
nor U3736 (N_3736,N_3589,N_3580);
or U3737 (N_3737,N_3414,N_3503);
nor U3738 (N_3738,N_3463,N_3457);
or U3739 (N_3739,N_3422,N_3583);
xor U3740 (N_3740,N_3459,N_3468);
nand U3741 (N_3741,N_3419,N_3428);
and U3742 (N_3742,N_3573,N_3412);
nor U3743 (N_3743,N_3465,N_3476);
xnor U3744 (N_3744,N_3414,N_3576);
or U3745 (N_3745,N_3463,N_3570);
xnor U3746 (N_3746,N_3420,N_3505);
or U3747 (N_3747,N_3416,N_3528);
nor U3748 (N_3748,N_3482,N_3534);
and U3749 (N_3749,N_3579,N_3415);
or U3750 (N_3750,N_3465,N_3579);
and U3751 (N_3751,N_3568,N_3572);
or U3752 (N_3752,N_3547,N_3470);
and U3753 (N_3753,N_3541,N_3521);
and U3754 (N_3754,N_3481,N_3479);
nand U3755 (N_3755,N_3490,N_3590);
xnor U3756 (N_3756,N_3584,N_3493);
and U3757 (N_3757,N_3520,N_3461);
nand U3758 (N_3758,N_3503,N_3519);
xor U3759 (N_3759,N_3574,N_3525);
or U3760 (N_3760,N_3482,N_3429);
nor U3761 (N_3761,N_3464,N_3585);
or U3762 (N_3762,N_3413,N_3496);
xor U3763 (N_3763,N_3445,N_3485);
nor U3764 (N_3764,N_3432,N_3452);
nor U3765 (N_3765,N_3574,N_3515);
xor U3766 (N_3766,N_3452,N_3572);
nor U3767 (N_3767,N_3475,N_3407);
or U3768 (N_3768,N_3463,N_3498);
and U3769 (N_3769,N_3529,N_3566);
and U3770 (N_3770,N_3445,N_3479);
nor U3771 (N_3771,N_3479,N_3462);
nor U3772 (N_3772,N_3554,N_3434);
and U3773 (N_3773,N_3567,N_3468);
nand U3774 (N_3774,N_3540,N_3596);
or U3775 (N_3775,N_3410,N_3412);
or U3776 (N_3776,N_3592,N_3594);
nor U3777 (N_3777,N_3595,N_3556);
or U3778 (N_3778,N_3436,N_3595);
or U3779 (N_3779,N_3452,N_3482);
xor U3780 (N_3780,N_3595,N_3523);
nand U3781 (N_3781,N_3417,N_3410);
xor U3782 (N_3782,N_3427,N_3471);
and U3783 (N_3783,N_3430,N_3510);
xor U3784 (N_3784,N_3446,N_3571);
xor U3785 (N_3785,N_3582,N_3462);
nand U3786 (N_3786,N_3507,N_3502);
nand U3787 (N_3787,N_3500,N_3577);
and U3788 (N_3788,N_3562,N_3416);
nand U3789 (N_3789,N_3436,N_3576);
or U3790 (N_3790,N_3564,N_3545);
nand U3791 (N_3791,N_3486,N_3543);
xor U3792 (N_3792,N_3456,N_3521);
and U3793 (N_3793,N_3512,N_3524);
nor U3794 (N_3794,N_3549,N_3502);
nor U3795 (N_3795,N_3538,N_3567);
nor U3796 (N_3796,N_3522,N_3521);
or U3797 (N_3797,N_3453,N_3429);
and U3798 (N_3798,N_3417,N_3476);
and U3799 (N_3799,N_3410,N_3515);
nor U3800 (N_3800,N_3674,N_3605);
xnor U3801 (N_3801,N_3661,N_3657);
xnor U3802 (N_3802,N_3743,N_3707);
and U3803 (N_3803,N_3662,N_3617);
and U3804 (N_3804,N_3742,N_3749);
xor U3805 (N_3805,N_3640,N_3744);
nor U3806 (N_3806,N_3687,N_3664);
xor U3807 (N_3807,N_3679,N_3761);
or U3808 (N_3808,N_3784,N_3636);
nor U3809 (N_3809,N_3748,N_3633);
xnor U3810 (N_3810,N_3625,N_3634);
and U3811 (N_3811,N_3793,N_3788);
or U3812 (N_3812,N_3705,N_3733);
nand U3813 (N_3813,N_3727,N_3686);
and U3814 (N_3814,N_3663,N_3780);
or U3815 (N_3815,N_3624,N_3692);
nor U3816 (N_3816,N_3650,N_3794);
and U3817 (N_3817,N_3773,N_3714);
nand U3818 (N_3818,N_3741,N_3771);
or U3819 (N_3819,N_3632,N_3729);
or U3820 (N_3820,N_3680,N_3764);
nand U3821 (N_3821,N_3683,N_3607);
nor U3822 (N_3822,N_3765,N_3772);
nand U3823 (N_3823,N_3665,N_3659);
nand U3824 (N_3824,N_3739,N_3647);
nor U3825 (N_3825,N_3658,N_3715);
nand U3826 (N_3826,N_3734,N_3635);
nor U3827 (N_3827,N_3775,N_3668);
or U3828 (N_3828,N_3614,N_3629);
nand U3829 (N_3829,N_3756,N_3768);
nor U3830 (N_3830,N_3783,N_3667);
nor U3831 (N_3831,N_3646,N_3696);
nor U3832 (N_3832,N_3758,N_3796);
or U3833 (N_3833,N_3785,N_3799);
nand U3834 (N_3834,N_3631,N_3701);
nand U3835 (N_3835,N_3601,N_3722);
xnor U3836 (N_3836,N_3672,N_3637);
nor U3837 (N_3837,N_3755,N_3704);
xnor U3838 (N_3838,N_3754,N_3712);
and U3839 (N_3839,N_3612,N_3676);
xor U3840 (N_3840,N_3751,N_3735);
xnor U3841 (N_3841,N_3747,N_3623);
xnor U3842 (N_3842,N_3767,N_3684);
xor U3843 (N_3843,N_3621,N_3675);
and U3844 (N_3844,N_3725,N_3613);
and U3845 (N_3845,N_3738,N_3797);
nand U3846 (N_3846,N_3770,N_3719);
nand U3847 (N_3847,N_3654,N_3723);
nor U3848 (N_3848,N_3746,N_3792);
or U3849 (N_3849,N_3753,N_3721);
nor U3850 (N_3850,N_3626,N_3791);
or U3851 (N_3851,N_3622,N_3651);
nor U3852 (N_3852,N_3777,N_3609);
nor U3853 (N_3853,N_3763,N_3627);
or U3854 (N_3854,N_3685,N_3769);
nand U3855 (N_3855,N_3731,N_3728);
nor U3856 (N_3856,N_3697,N_3699);
nor U3857 (N_3857,N_3611,N_3642);
xnor U3858 (N_3858,N_3736,N_3606);
nor U3859 (N_3859,N_3678,N_3600);
and U3860 (N_3860,N_3610,N_3652);
nor U3861 (N_3861,N_3759,N_3694);
or U3862 (N_3862,N_3762,N_3677);
xor U3863 (N_3863,N_3700,N_3781);
xnor U3864 (N_3864,N_3655,N_3670);
xor U3865 (N_3865,N_3766,N_3776);
nor U3866 (N_3866,N_3724,N_3710);
nor U3867 (N_3867,N_3618,N_3602);
or U3868 (N_3868,N_3778,N_3604);
nand U3869 (N_3869,N_3682,N_3750);
xnor U3870 (N_3870,N_3774,N_3703);
nand U3871 (N_3871,N_3645,N_3666);
or U3872 (N_3872,N_3644,N_3745);
or U3873 (N_3873,N_3691,N_3779);
and U3874 (N_3874,N_3630,N_3620);
xnor U3875 (N_3875,N_3786,N_3681);
nand U3876 (N_3876,N_3671,N_3757);
and U3877 (N_3877,N_3709,N_3732);
or U3878 (N_3878,N_3615,N_3716);
and U3879 (N_3879,N_3737,N_3660);
xnor U3880 (N_3880,N_3713,N_3688);
xor U3881 (N_3881,N_3718,N_3726);
nand U3882 (N_3882,N_3711,N_3690);
nor U3883 (N_3883,N_3603,N_3648);
nand U3884 (N_3884,N_3693,N_3689);
or U3885 (N_3885,N_3717,N_3638);
xnor U3886 (N_3886,N_3619,N_3608);
nand U3887 (N_3887,N_3616,N_3789);
nand U3888 (N_3888,N_3695,N_3643);
or U3889 (N_3889,N_3798,N_3628);
and U3890 (N_3890,N_3653,N_3673);
nand U3891 (N_3891,N_3782,N_3787);
nor U3892 (N_3892,N_3708,N_3730);
nand U3893 (N_3893,N_3760,N_3656);
nand U3894 (N_3894,N_3795,N_3740);
xnor U3895 (N_3895,N_3649,N_3641);
and U3896 (N_3896,N_3639,N_3790);
nand U3897 (N_3897,N_3752,N_3669);
and U3898 (N_3898,N_3702,N_3698);
xor U3899 (N_3899,N_3706,N_3720);
nor U3900 (N_3900,N_3696,N_3670);
or U3901 (N_3901,N_3716,N_3734);
xnor U3902 (N_3902,N_3758,N_3788);
nor U3903 (N_3903,N_3776,N_3616);
and U3904 (N_3904,N_3655,N_3749);
xnor U3905 (N_3905,N_3796,N_3621);
nand U3906 (N_3906,N_3716,N_3626);
or U3907 (N_3907,N_3748,N_3749);
xor U3908 (N_3908,N_3716,N_3612);
xnor U3909 (N_3909,N_3654,N_3660);
nand U3910 (N_3910,N_3602,N_3708);
nor U3911 (N_3911,N_3611,N_3778);
or U3912 (N_3912,N_3646,N_3773);
xnor U3913 (N_3913,N_3678,N_3694);
or U3914 (N_3914,N_3608,N_3673);
nand U3915 (N_3915,N_3615,N_3745);
xor U3916 (N_3916,N_3610,N_3631);
nor U3917 (N_3917,N_3620,N_3609);
or U3918 (N_3918,N_3660,N_3618);
and U3919 (N_3919,N_3791,N_3729);
nand U3920 (N_3920,N_3636,N_3765);
nor U3921 (N_3921,N_3678,N_3740);
or U3922 (N_3922,N_3675,N_3601);
xnor U3923 (N_3923,N_3695,N_3756);
xor U3924 (N_3924,N_3628,N_3609);
and U3925 (N_3925,N_3621,N_3674);
xnor U3926 (N_3926,N_3792,N_3689);
nand U3927 (N_3927,N_3713,N_3654);
or U3928 (N_3928,N_3788,N_3649);
and U3929 (N_3929,N_3775,N_3778);
xnor U3930 (N_3930,N_3716,N_3613);
or U3931 (N_3931,N_3617,N_3668);
nor U3932 (N_3932,N_3739,N_3635);
and U3933 (N_3933,N_3750,N_3745);
nor U3934 (N_3934,N_3759,N_3678);
xnor U3935 (N_3935,N_3608,N_3701);
nor U3936 (N_3936,N_3621,N_3618);
and U3937 (N_3937,N_3715,N_3610);
nand U3938 (N_3938,N_3744,N_3604);
and U3939 (N_3939,N_3665,N_3683);
nand U3940 (N_3940,N_3744,N_3735);
and U3941 (N_3941,N_3679,N_3752);
nand U3942 (N_3942,N_3608,N_3786);
or U3943 (N_3943,N_3782,N_3646);
nand U3944 (N_3944,N_3748,N_3774);
xnor U3945 (N_3945,N_3618,N_3647);
xnor U3946 (N_3946,N_3624,N_3735);
and U3947 (N_3947,N_3722,N_3688);
nand U3948 (N_3948,N_3708,N_3766);
and U3949 (N_3949,N_3772,N_3780);
or U3950 (N_3950,N_3799,N_3708);
nor U3951 (N_3951,N_3778,N_3621);
nand U3952 (N_3952,N_3731,N_3668);
nand U3953 (N_3953,N_3646,N_3612);
xnor U3954 (N_3954,N_3780,N_3728);
nor U3955 (N_3955,N_3719,N_3724);
or U3956 (N_3956,N_3667,N_3606);
xnor U3957 (N_3957,N_3709,N_3666);
or U3958 (N_3958,N_3773,N_3670);
xnor U3959 (N_3959,N_3627,N_3736);
xor U3960 (N_3960,N_3757,N_3680);
and U3961 (N_3961,N_3721,N_3763);
or U3962 (N_3962,N_3662,N_3730);
or U3963 (N_3963,N_3651,N_3797);
and U3964 (N_3964,N_3672,N_3765);
or U3965 (N_3965,N_3634,N_3665);
nor U3966 (N_3966,N_3735,N_3634);
and U3967 (N_3967,N_3629,N_3606);
nor U3968 (N_3968,N_3789,N_3700);
or U3969 (N_3969,N_3796,N_3747);
or U3970 (N_3970,N_3755,N_3762);
and U3971 (N_3971,N_3608,N_3797);
xnor U3972 (N_3972,N_3719,N_3728);
nor U3973 (N_3973,N_3647,N_3781);
xnor U3974 (N_3974,N_3615,N_3620);
nor U3975 (N_3975,N_3669,N_3737);
and U3976 (N_3976,N_3748,N_3609);
xor U3977 (N_3977,N_3620,N_3732);
or U3978 (N_3978,N_3739,N_3617);
or U3979 (N_3979,N_3761,N_3788);
nand U3980 (N_3980,N_3651,N_3778);
or U3981 (N_3981,N_3797,N_3652);
or U3982 (N_3982,N_3653,N_3675);
nor U3983 (N_3983,N_3706,N_3740);
and U3984 (N_3984,N_3729,N_3681);
and U3985 (N_3985,N_3629,N_3715);
nor U3986 (N_3986,N_3716,N_3635);
xnor U3987 (N_3987,N_3622,N_3687);
or U3988 (N_3988,N_3720,N_3740);
and U3989 (N_3989,N_3720,N_3770);
nand U3990 (N_3990,N_3716,N_3737);
or U3991 (N_3991,N_3702,N_3704);
xor U3992 (N_3992,N_3763,N_3698);
nand U3993 (N_3993,N_3727,N_3642);
nand U3994 (N_3994,N_3624,N_3711);
nor U3995 (N_3995,N_3646,N_3627);
xnor U3996 (N_3996,N_3772,N_3674);
or U3997 (N_3997,N_3645,N_3688);
nand U3998 (N_3998,N_3643,N_3670);
xnor U3999 (N_3999,N_3668,N_3664);
nor U4000 (N_4000,N_3809,N_3829);
nor U4001 (N_4001,N_3816,N_3876);
nand U4002 (N_4002,N_3835,N_3971);
xnor U4003 (N_4003,N_3860,N_3975);
xnor U4004 (N_4004,N_3807,N_3909);
nor U4005 (N_4005,N_3950,N_3849);
xor U4006 (N_4006,N_3853,N_3962);
and U4007 (N_4007,N_3918,N_3992);
or U4008 (N_4008,N_3923,N_3899);
xor U4009 (N_4009,N_3877,N_3949);
nor U4010 (N_4010,N_3999,N_3805);
xor U4011 (N_4011,N_3969,N_3940);
or U4012 (N_4012,N_3916,N_3961);
xnor U4013 (N_4013,N_3884,N_3984);
nor U4014 (N_4014,N_3886,N_3904);
nand U4015 (N_4015,N_3836,N_3817);
and U4016 (N_4016,N_3953,N_3878);
nand U4017 (N_4017,N_3910,N_3821);
xor U4018 (N_4018,N_3951,N_3841);
nor U4019 (N_4019,N_3855,N_3881);
nor U4020 (N_4020,N_3943,N_3956);
and U4021 (N_4021,N_3813,N_3926);
nor U4022 (N_4022,N_3939,N_3814);
nor U4023 (N_4023,N_3907,N_3867);
or U4024 (N_4024,N_3968,N_3862);
xnor U4025 (N_4025,N_3919,N_3812);
or U4026 (N_4026,N_3858,N_3942);
and U4027 (N_4027,N_3966,N_3959);
nor U4028 (N_4028,N_3917,N_3868);
nand U4029 (N_4029,N_3838,N_3852);
xnor U4030 (N_4030,N_3839,N_3982);
nor U4031 (N_4031,N_3882,N_3801);
nor U4032 (N_4032,N_3811,N_3911);
and U4033 (N_4033,N_3987,N_3800);
and U4034 (N_4034,N_3879,N_3998);
xnor U4035 (N_4035,N_3818,N_3922);
nand U4036 (N_4036,N_3850,N_3927);
nor U4037 (N_4037,N_3967,N_3955);
and U4038 (N_4038,N_3820,N_3897);
or U4039 (N_4039,N_3828,N_3819);
and U4040 (N_4040,N_3827,N_3833);
nand U4041 (N_4041,N_3986,N_3857);
nor U4042 (N_4042,N_3941,N_3854);
and U4043 (N_4043,N_3823,N_3848);
xor U4044 (N_4044,N_3974,N_3981);
xor U4045 (N_4045,N_3920,N_3834);
or U4046 (N_4046,N_3832,N_3880);
or U4047 (N_4047,N_3865,N_3875);
or U4048 (N_4048,N_3863,N_3985);
xnor U4049 (N_4049,N_3806,N_3895);
nor U4050 (N_4050,N_3997,N_3845);
xnor U4051 (N_4051,N_3869,N_3932);
or U4052 (N_4052,N_3893,N_3891);
nand U4053 (N_4053,N_3996,N_3921);
nor U4054 (N_4054,N_3871,N_3948);
and U4055 (N_4055,N_3808,N_3844);
nor U4056 (N_4056,N_3892,N_3831);
nand U4057 (N_4057,N_3952,N_3973);
xor U4058 (N_4058,N_3933,N_3908);
nand U4059 (N_4059,N_3957,N_3898);
and U4060 (N_4060,N_3914,N_3924);
xor U4061 (N_4061,N_3937,N_3979);
nand U4062 (N_4062,N_3993,N_3815);
and U4063 (N_4063,N_3885,N_3803);
nor U4064 (N_4064,N_3912,N_3837);
nand U4065 (N_4065,N_3847,N_3822);
nor U4066 (N_4066,N_3915,N_3980);
xor U4067 (N_4067,N_3935,N_3954);
nand U4068 (N_4068,N_3965,N_3851);
nand U4069 (N_4069,N_3931,N_3856);
and U4070 (N_4070,N_3874,N_3983);
nor U4071 (N_4071,N_3901,N_3936);
or U4072 (N_4072,N_3970,N_3842);
xnor U4073 (N_4073,N_3896,N_3988);
and U4074 (N_4074,N_3894,N_3846);
or U4075 (N_4075,N_3866,N_3928);
and U4076 (N_4076,N_3903,N_3913);
and U4077 (N_4077,N_3840,N_3978);
nor U4078 (N_4078,N_3989,N_3944);
and U4079 (N_4079,N_3824,N_3964);
nor U4080 (N_4080,N_3990,N_3902);
and U4081 (N_4081,N_3906,N_3900);
xor U4082 (N_4082,N_3883,N_3890);
or U4083 (N_4083,N_3946,N_3930);
nor U4084 (N_4084,N_3960,N_3830);
nor U4085 (N_4085,N_3995,N_3826);
nand U4086 (N_4086,N_3888,N_3934);
nand U4087 (N_4087,N_3872,N_3825);
or U4088 (N_4088,N_3958,N_3889);
or U4089 (N_4089,N_3810,N_3905);
nand U4090 (N_4090,N_3925,N_3864);
and U4091 (N_4091,N_3861,N_3870);
and U4092 (N_4092,N_3977,N_3947);
and U4093 (N_4093,N_3804,N_3802);
or U4094 (N_4094,N_3859,N_3994);
nand U4095 (N_4095,N_3929,N_3938);
and U4096 (N_4096,N_3843,N_3963);
and U4097 (N_4097,N_3873,N_3972);
xnor U4098 (N_4098,N_3991,N_3976);
nor U4099 (N_4099,N_3887,N_3945);
or U4100 (N_4100,N_3885,N_3865);
or U4101 (N_4101,N_3988,N_3940);
or U4102 (N_4102,N_3877,N_3820);
or U4103 (N_4103,N_3904,N_3823);
xnor U4104 (N_4104,N_3815,N_3889);
xnor U4105 (N_4105,N_3978,N_3891);
or U4106 (N_4106,N_3966,N_3991);
xnor U4107 (N_4107,N_3990,N_3888);
nand U4108 (N_4108,N_3926,N_3936);
xnor U4109 (N_4109,N_3867,N_3814);
and U4110 (N_4110,N_3812,N_3842);
or U4111 (N_4111,N_3816,N_3805);
and U4112 (N_4112,N_3887,N_3931);
nand U4113 (N_4113,N_3868,N_3919);
or U4114 (N_4114,N_3822,N_3828);
and U4115 (N_4115,N_3981,N_3836);
and U4116 (N_4116,N_3859,N_3947);
nand U4117 (N_4117,N_3937,N_3838);
nand U4118 (N_4118,N_3949,N_3897);
nor U4119 (N_4119,N_3890,N_3874);
xnor U4120 (N_4120,N_3834,N_3878);
and U4121 (N_4121,N_3808,N_3801);
xor U4122 (N_4122,N_3807,N_3819);
xor U4123 (N_4123,N_3920,N_3845);
and U4124 (N_4124,N_3991,N_3895);
nor U4125 (N_4125,N_3960,N_3981);
or U4126 (N_4126,N_3935,N_3809);
or U4127 (N_4127,N_3943,N_3835);
nor U4128 (N_4128,N_3820,N_3899);
nor U4129 (N_4129,N_3804,N_3903);
xnor U4130 (N_4130,N_3850,N_3859);
or U4131 (N_4131,N_3807,N_3890);
nor U4132 (N_4132,N_3973,N_3819);
and U4133 (N_4133,N_3848,N_3985);
nand U4134 (N_4134,N_3946,N_3962);
xnor U4135 (N_4135,N_3949,N_3936);
nand U4136 (N_4136,N_3912,N_3845);
nand U4137 (N_4137,N_3975,N_3862);
nand U4138 (N_4138,N_3971,N_3975);
nor U4139 (N_4139,N_3804,N_3827);
or U4140 (N_4140,N_3804,N_3885);
nor U4141 (N_4141,N_3869,N_3862);
xor U4142 (N_4142,N_3946,N_3843);
or U4143 (N_4143,N_3838,N_3833);
nor U4144 (N_4144,N_3935,N_3881);
xor U4145 (N_4145,N_3945,N_3912);
xor U4146 (N_4146,N_3837,N_3923);
xor U4147 (N_4147,N_3996,N_3947);
nor U4148 (N_4148,N_3933,N_3939);
nor U4149 (N_4149,N_3812,N_3847);
and U4150 (N_4150,N_3916,N_3969);
and U4151 (N_4151,N_3811,N_3806);
xor U4152 (N_4152,N_3819,N_3843);
xnor U4153 (N_4153,N_3813,N_3954);
and U4154 (N_4154,N_3931,N_3918);
nand U4155 (N_4155,N_3882,N_3973);
nand U4156 (N_4156,N_3896,N_3884);
nand U4157 (N_4157,N_3920,N_3946);
nand U4158 (N_4158,N_3953,N_3927);
and U4159 (N_4159,N_3860,N_3863);
and U4160 (N_4160,N_3852,N_3848);
or U4161 (N_4161,N_3957,N_3845);
xor U4162 (N_4162,N_3936,N_3948);
or U4163 (N_4163,N_3883,N_3993);
nor U4164 (N_4164,N_3841,N_3966);
nand U4165 (N_4165,N_3962,N_3945);
nor U4166 (N_4166,N_3965,N_3898);
and U4167 (N_4167,N_3855,N_3862);
nand U4168 (N_4168,N_3826,N_3914);
nand U4169 (N_4169,N_3975,N_3989);
and U4170 (N_4170,N_3925,N_3830);
or U4171 (N_4171,N_3806,N_3997);
xor U4172 (N_4172,N_3870,N_3912);
and U4173 (N_4173,N_3948,N_3937);
xnor U4174 (N_4174,N_3919,N_3987);
and U4175 (N_4175,N_3876,N_3829);
nand U4176 (N_4176,N_3963,N_3864);
nor U4177 (N_4177,N_3898,N_3977);
nand U4178 (N_4178,N_3971,N_3843);
or U4179 (N_4179,N_3930,N_3847);
or U4180 (N_4180,N_3908,N_3815);
nand U4181 (N_4181,N_3943,N_3863);
xor U4182 (N_4182,N_3962,N_3891);
nor U4183 (N_4183,N_3809,N_3878);
nand U4184 (N_4184,N_3850,N_3809);
nand U4185 (N_4185,N_3969,N_3837);
xor U4186 (N_4186,N_3837,N_3801);
nor U4187 (N_4187,N_3890,N_3840);
xor U4188 (N_4188,N_3951,N_3834);
xor U4189 (N_4189,N_3997,N_3974);
xnor U4190 (N_4190,N_3857,N_3846);
or U4191 (N_4191,N_3987,N_3949);
xor U4192 (N_4192,N_3820,N_3822);
nor U4193 (N_4193,N_3902,N_3853);
and U4194 (N_4194,N_3940,N_3937);
nand U4195 (N_4195,N_3914,N_3886);
nand U4196 (N_4196,N_3865,N_3844);
and U4197 (N_4197,N_3925,N_3944);
xor U4198 (N_4198,N_3851,N_3943);
nor U4199 (N_4199,N_3964,N_3945);
or U4200 (N_4200,N_4160,N_4123);
nand U4201 (N_4201,N_4106,N_4136);
nor U4202 (N_4202,N_4055,N_4194);
or U4203 (N_4203,N_4151,N_4022);
or U4204 (N_4204,N_4139,N_4019);
xor U4205 (N_4205,N_4178,N_4148);
nand U4206 (N_4206,N_4075,N_4078);
nor U4207 (N_4207,N_4095,N_4067);
and U4208 (N_4208,N_4193,N_4119);
or U4209 (N_4209,N_4066,N_4058);
xor U4210 (N_4210,N_4083,N_4175);
nand U4211 (N_4211,N_4086,N_4161);
xnor U4212 (N_4212,N_4018,N_4189);
and U4213 (N_4213,N_4185,N_4147);
and U4214 (N_4214,N_4035,N_4121);
nor U4215 (N_4215,N_4011,N_4001);
xnor U4216 (N_4216,N_4039,N_4124);
nand U4217 (N_4217,N_4113,N_4156);
or U4218 (N_4218,N_4159,N_4199);
or U4219 (N_4219,N_4037,N_4181);
nand U4220 (N_4220,N_4026,N_4004);
nor U4221 (N_4221,N_4056,N_4021);
and U4222 (N_4222,N_4071,N_4168);
nor U4223 (N_4223,N_4182,N_4177);
nor U4224 (N_4224,N_4135,N_4009);
and U4225 (N_4225,N_4081,N_4167);
or U4226 (N_4226,N_4012,N_4120);
or U4227 (N_4227,N_4010,N_4129);
xnor U4228 (N_4228,N_4100,N_4032);
and U4229 (N_4229,N_4154,N_4062);
xnor U4230 (N_4230,N_4079,N_4198);
xnor U4231 (N_4231,N_4112,N_4165);
nor U4232 (N_4232,N_4036,N_4180);
xnor U4233 (N_4233,N_4153,N_4025);
and U4234 (N_4234,N_4184,N_4163);
or U4235 (N_4235,N_4031,N_4104);
and U4236 (N_4236,N_4152,N_4099);
nor U4237 (N_4237,N_4195,N_4146);
nand U4238 (N_4238,N_4110,N_4085);
nand U4239 (N_4239,N_4063,N_4028);
nor U4240 (N_4240,N_4109,N_4057);
nor U4241 (N_4241,N_4142,N_4150);
or U4242 (N_4242,N_4014,N_4125);
nand U4243 (N_4243,N_4131,N_4134);
nand U4244 (N_4244,N_4061,N_4138);
nor U4245 (N_4245,N_4111,N_4137);
or U4246 (N_4246,N_4087,N_4197);
nand U4247 (N_4247,N_4044,N_4164);
and U4248 (N_4248,N_4076,N_4141);
nand U4249 (N_4249,N_4038,N_4192);
or U4250 (N_4250,N_4023,N_4082);
or U4251 (N_4251,N_4068,N_4060);
and U4252 (N_4252,N_4000,N_4027);
and U4253 (N_4253,N_4116,N_4080);
nand U4254 (N_4254,N_4054,N_4126);
and U4255 (N_4255,N_4017,N_4140);
or U4256 (N_4256,N_4097,N_4077);
nor U4257 (N_4257,N_4034,N_4187);
and U4258 (N_4258,N_4145,N_4105);
xnor U4259 (N_4259,N_4162,N_4045);
or U4260 (N_4260,N_4051,N_4002);
nor U4261 (N_4261,N_4093,N_4042);
xnor U4262 (N_4262,N_4172,N_4094);
or U4263 (N_4263,N_4005,N_4128);
and U4264 (N_4264,N_4047,N_4191);
nor U4265 (N_4265,N_4130,N_4174);
nor U4266 (N_4266,N_4101,N_4003);
nand U4267 (N_4267,N_4006,N_4183);
or U4268 (N_4268,N_4170,N_4046);
xor U4269 (N_4269,N_4065,N_4030);
nor U4270 (N_4270,N_4052,N_4020);
xnor U4271 (N_4271,N_4098,N_4158);
nor U4272 (N_4272,N_4029,N_4090);
and U4273 (N_4273,N_4024,N_4016);
nor U4274 (N_4274,N_4049,N_4118);
nor U4275 (N_4275,N_4103,N_4089);
xnor U4276 (N_4276,N_4008,N_4157);
nor U4277 (N_4277,N_4149,N_4173);
nor U4278 (N_4278,N_4007,N_4143);
nand U4279 (N_4279,N_4050,N_4179);
nand U4280 (N_4280,N_4070,N_4186);
nor U4281 (N_4281,N_4048,N_4096);
xnor U4282 (N_4282,N_4074,N_4072);
or U4283 (N_4283,N_4133,N_4132);
xnor U4284 (N_4284,N_4107,N_4069);
nor U4285 (N_4285,N_4190,N_4073);
and U4286 (N_4286,N_4196,N_4084);
or U4287 (N_4287,N_4166,N_4040);
nor U4288 (N_4288,N_4117,N_4092);
and U4289 (N_4289,N_4064,N_4053);
nor U4290 (N_4290,N_4169,N_4043);
and U4291 (N_4291,N_4188,N_4115);
nand U4292 (N_4292,N_4114,N_4091);
xor U4293 (N_4293,N_4013,N_4015);
nand U4294 (N_4294,N_4102,N_4171);
nor U4295 (N_4295,N_4059,N_4108);
and U4296 (N_4296,N_4127,N_4144);
and U4297 (N_4297,N_4033,N_4041);
nand U4298 (N_4298,N_4088,N_4176);
nand U4299 (N_4299,N_4155,N_4122);
or U4300 (N_4300,N_4161,N_4015);
or U4301 (N_4301,N_4192,N_4031);
and U4302 (N_4302,N_4117,N_4134);
nor U4303 (N_4303,N_4012,N_4178);
or U4304 (N_4304,N_4103,N_4149);
nor U4305 (N_4305,N_4053,N_4027);
xnor U4306 (N_4306,N_4187,N_4006);
xor U4307 (N_4307,N_4182,N_4010);
xnor U4308 (N_4308,N_4022,N_4122);
nor U4309 (N_4309,N_4060,N_4138);
nand U4310 (N_4310,N_4176,N_4012);
and U4311 (N_4311,N_4091,N_4163);
nand U4312 (N_4312,N_4029,N_4191);
nor U4313 (N_4313,N_4108,N_4159);
nor U4314 (N_4314,N_4120,N_4148);
xor U4315 (N_4315,N_4169,N_4017);
xnor U4316 (N_4316,N_4170,N_4082);
and U4317 (N_4317,N_4112,N_4013);
nand U4318 (N_4318,N_4141,N_4089);
nor U4319 (N_4319,N_4043,N_4052);
nor U4320 (N_4320,N_4031,N_4160);
or U4321 (N_4321,N_4080,N_4091);
and U4322 (N_4322,N_4049,N_4047);
and U4323 (N_4323,N_4115,N_4111);
or U4324 (N_4324,N_4034,N_4182);
nor U4325 (N_4325,N_4090,N_4015);
or U4326 (N_4326,N_4111,N_4012);
nand U4327 (N_4327,N_4168,N_4179);
nor U4328 (N_4328,N_4016,N_4079);
and U4329 (N_4329,N_4090,N_4096);
or U4330 (N_4330,N_4184,N_4061);
xor U4331 (N_4331,N_4086,N_4011);
nand U4332 (N_4332,N_4030,N_4143);
xnor U4333 (N_4333,N_4149,N_4102);
nor U4334 (N_4334,N_4169,N_4053);
nand U4335 (N_4335,N_4065,N_4117);
or U4336 (N_4336,N_4186,N_4177);
xnor U4337 (N_4337,N_4019,N_4039);
and U4338 (N_4338,N_4025,N_4151);
xor U4339 (N_4339,N_4196,N_4190);
nand U4340 (N_4340,N_4148,N_4019);
nor U4341 (N_4341,N_4128,N_4034);
or U4342 (N_4342,N_4040,N_4130);
nor U4343 (N_4343,N_4194,N_4056);
nor U4344 (N_4344,N_4012,N_4025);
xor U4345 (N_4345,N_4084,N_4162);
nor U4346 (N_4346,N_4192,N_4081);
nor U4347 (N_4347,N_4119,N_4073);
and U4348 (N_4348,N_4196,N_4127);
nor U4349 (N_4349,N_4126,N_4060);
and U4350 (N_4350,N_4047,N_4165);
or U4351 (N_4351,N_4000,N_4176);
xnor U4352 (N_4352,N_4167,N_4139);
or U4353 (N_4353,N_4086,N_4138);
or U4354 (N_4354,N_4015,N_4153);
nor U4355 (N_4355,N_4013,N_4082);
xor U4356 (N_4356,N_4093,N_4175);
nand U4357 (N_4357,N_4115,N_4184);
and U4358 (N_4358,N_4036,N_4081);
or U4359 (N_4359,N_4090,N_4056);
and U4360 (N_4360,N_4102,N_4075);
xor U4361 (N_4361,N_4088,N_4131);
nor U4362 (N_4362,N_4192,N_4170);
nand U4363 (N_4363,N_4181,N_4033);
nand U4364 (N_4364,N_4097,N_4143);
nand U4365 (N_4365,N_4110,N_4186);
and U4366 (N_4366,N_4161,N_4147);
or U4367 (N_4367,N_4195,N_4011);
nand U4368 (N_4368,N_4059,N_4074);
xnor U4369 (N_4369,N_4083,N_4031);
nor U4370 (N_4370,N_4018,N_4106);
nor U4371 (N_4371,N_4040,N_4025);
xnor U4372 (N_4372,N_4149,N_4086);
nand U4373 (N_4373,N_4103,N_4115);
nand U4374 (N_4374,N_4137,N_4107);
nand U4375 (N_4375,N_4015,N_4026);
and U4376 (N_4376,N_4171,N_4084);
nor U4377 (N_4377,N_4125,N_4059);
xor U4378 (N_4378,N_4179,N_4119);
nor U4379 (N_4379,N_4090,N_4105);
or U4380 (N_4380,N_4016,N_4028);
nor U4381 (N_4381,N_4175,N_4098);
nor U4382 (N_4382,N_4018,N_4133);
xnor U4383 (N_4383,N_4023,N_4103);
nand U4384 (N_4384,N_4159,N_4198);
nand U4385 (N_4385,N_4083,N_4136);
or U4386 (N_4386,N_4007,N_4097);
xor U4387 (N_4387,N_4022,N_4137);
nor U4388 (N_4388,N_4035,N_4058);
nand U4389 (N_4389,N_4090,N_4110);
xor U4390 (N_4390,N_4114,N_4141);
or U4391 (N_4391,N_4195,N_4098);
and U4392 (N_4392,N_4130,N_4173);
xnor U4393 (N_4393,N_4176,N_4109);
nor U4394 (N_4394,N_4141,N_4167);
xor U4395 (N_4395,N_4127,N_4026);
nand U4396 (N_4396,N_4122,N_4139);
nor U4397 (N_4397,N_4162,N_4133);
xor U4398 (N_4398,N_4034,N_4004);
nand U4399 (N_4399,N_4023,N_4035);
xor U4400 (N_4400,N_4225,N_4254);
nor U4401 (N_4401,N_4348,N_4280);
nor U4402 (N_4402,N_4204,N_4372);
nor U4403 (N_4403,N_4325,N_4290);
xor U4404 (N_4404,N_4316,N_4217);
nand U4405 (N_4405,N_4265,N_4321);
and U4406 (N_4406,N_4359,N_4271);
and U4407 (N_4407,N_4337,N_4390);
or U4408 (N_4408,N_4212,N_4356);
and U4409 (N_4409,N_4261,N_4329);
or U4410 (N_4410,N_4377,N_4393);
nor U4411 (N_4411,N_4236,N_4209);
nor U4412 (N_4412,N_4244,N_4281);
xor U4413 (N_4413,N_4245,N_4363);
xor U4414 (N_4414,N_4331,N_4397);
and U4415 (N_4415,N_4311,N_4362);
and U4416 (N_4416,N_4333,N_4279);
or U4417 (N_4417,N_4259,N_4350);
or U4418 (N_4418,N_4273,N_4361);
xor U4419 (N_4419,N_4386,N_4205);
and U4420 (N_4420,N_4246,N_4305);
xnor U4421 (N_4421,N_4210,N_4360);
or U4422 (N_4422,N_4213,N_4349);
nor U4423 (N_4423,N_4260,N_4385);
nor U4424 (N_4424,N_4370,N_4282);
xor U4425 (N_4425,N_4297,N_4203);
nand U4426 (N_4426,N_4272,N_4354);
xor U4427 (N_4427,N_4310,N_4382);
xnor U4428 (N_4428,N_4270,N_4286);
and U4429 (N_4429,N_4215,N_4335);
nor U4430 (N_4430,N_4257,N_4275);
or U4431 (N_4431,N_4320,N_4276);
xor U4432 (N_4432,N_4317,N_4231);
or U4433 (N_4433,N_4322,N_4296);
and U4434 (N_4434,N_4375,N_4223);
and U4435 (N_4435,N_4251,N_4303);
xnor U4436 (N_4436,N_4340,N_4330);
xnor U4437 (N_4437,N_4396,N_4389);
xnor U4438 (N_4438,N_4289,N_4339);
nand U4439 (N_4439,N_4332,N_4308);
or U4440 (N_4440,N_4392,N_4307);
nor U4441 (N_4441,N_4237,N_4299);
and U4442 (N_4442,N_4219,N_4274);
nand U4443 (N_4443,N_4327,N_4364);
or U4444 (N_4444,N_4230,N_4222);
or U4445 (N_4445,N_4383,N_4394);
or U4446 (N_4446,N_4374,N_4309);
or U4447 (N_4447,N_4352,N_4224);
xor U4448 (N_4448,N_4267,N_4238);
xnor U4449 (N_4449,N_4234,N_4243);
nand U4450 (N_4450,N_4338,N_4268);
or U4451 (N_4451,N_4201,N_4284);
xnor U4452 (N_4452,N_4253,N_4206);
nor U4453 (N_4453,N_4380,N_4398);
or U4454 (N_4454,N_4241,N_4344);
and U4455 (N_4455,N_4326,N_4301);
nor U4456 (N_4456,N_4221,N_4379);
xnor U4457 (N_4457,N_4287,N_4306);
nand U4458 (N_4458,N_4351,N_4278);
xnor U4459 (N_4459,N_4292,N_4319);
nand U4460 (N_4460,N_4371,N_4358);
xnor U4461 (N_4461,N_4250,N_4249);
or U4462 (N_4462,N_4283,N_4343);
nor U4463 (N_4463,N_4315,N_4388);
and U4464 (N_4464,N_4264,N_4399);
xnor U4465 (N_4465,N_4387,N_4255);
and U4466 (N_4466,N_4247,N_4384);
nand U4467 (N_4467,N_4381,N_4346);
nand U4468 (N_4468,N_4334,N_4300);
and U4469 (N_4469,N_4345,N_4395);
xnor U4470 (N_4470,N_4314,N_4232);
nand U4471 (N_4471,N_4366,N_4336);
xor U4472 (N_4472,N_4207,N_4342);
nand U4473 (N_4473,N_4302,N_4248);
nand U4474 (N_4474,N_4355,N_4240);
xor U4475 (N_4475,N_4298,N_4365);
and U4476 (N_4476,N_4285,N_4256);
xnor U4477 (N_4477,N_4291,N_4214);
nor U4478 (N_4478,N_4220,N_4367);
or U4479 (N_4479,N_4200,N_4239);
xnor U4480 (N_4480,N_4312,N_4328);
nand U4481 (N_4481,N_4226,N_4323);
nand U4482 (N_4482,N_4211,N_4304);
nand U4483 (N_4483,N_4227,N_4252);
nand U4484 (N_4484,N_4347,N_4288);
or U4485 (N_4485,N_4357,N_4208);
xnor U4486 (N_4486,N_4266,N_4294);
nor U4487 (N_4487,N_4258,N_4233);
nor U4488 (N_4488,N_4353,N_4263);
nand U4489 (N_4489,N_4269,N_4313);
nor U4490 (N_4490,N_4228,N_4235);
or U4491 (N_4491,N_4318,N_4341);
xor U4492 (N_4492,N_4373,N_4378);
nor U4493 (N_4493,N_4368,N_4218);
nor U4494 (N_4494,N_4202,N_4293);
or U4495 (N_4495,N_4376,N_4391);
nand U4496 (N_4496,N_4229,N_4324);
xnor U4497 (N_4497,N_4242,N_4369);
nand U4498 (N_4498,N_4295,N_4277);
or U4499 (N_4499,N_4262,N_4216);
nand U4500 (N_4500,N_4282,N_4348);
xor U4501 (N_4501,N_4213,N_4229);
or U4502 (N_4502,N_4340,N_4220);
nand U4503 (N_4503,N_4319,N_4246);
xor U4504 (N_4504,N_4338,N_4264);
xor U4505 (N_4505,N_4321,N_4368);
and U4506 (N_4506,N_4339,N_4323);
and U4507 (N_4507,N_4398,N_4387);
and U4508 (N_4508,N_4356,N_4395);
nor U4509 (N_4509,N_4280,N_4213);
xnor U4510 (N_4510,N_4317,N_4319);
or U4511 (N_4511,N_4392,N_4341);
nor U4512 (N_4512,N_4231,N_4398);
or U4513 (N_4513,N_4206,N_4242);
and U4514 (N_4514,N_4365,N_4296);
nand U4515 (N_4515,N_4321,N_4342);
or U4516 (N_4516,N_4394,N_4366);
or U4517 (N_4517,N_4264,N_4266);
nor U4518 (N_4518,N_4390,N_4306);
nand U4519 (N_4519,N_4228,N_4262);
xor U4520 (N_4520,N_4324,N_4288);
nor U4521 (N_4521,N_4319,N_4327);
xor U4522 (N_4522,N_4314,N_4355);
and U4523 (N_4523,N_4308,N_4276);
nand U4524 (N_4524,N_4331,N_4364);
or U4525 (N_4525,N_4399,N_4284);
nor U4526 (N_4526,N_4230,N_4244);
nor U4527 (N_4527,N_4375,N_4393);
nand U4528 (N_4528,N_4340,N_4390);
or U4529 (N_4529,N_4204,N_4278);
nor U4530 (N_4530,N_4223,N_4248);
and U4531 (N_4531,N_4367,N_4286);
nor U4532 (N_4532,N_4287,N_4254);
nor U4533 (N_4533,N_4213,N_4335);
and U4534 (N_4534,N_4378,N_4225);
or U4535 (N_4535,N_4348,N_4340);
xor U4536 (N_4536,N_4335,N_4334);
and U4537 (N_4537,N_4241,N_4361);
and U4538 (N_4538,N_4321,N_4293);
nand U4539 (N_4539,N_4331,N_4203);
or U4540 (N_4540,N_4205,N_4254);
or U4541 (N_4541,N_4277,N_4203);
nand U4542 (N_4542,N_4222,N_4249);
xnor U4543 (N_4543,N_4290,N_4285);
and U4544 (N_4544,N_4362,N_4211);
nand U4545 (N_4545,N_4262,N_4211);
and U4546 (N_4546,N_4237,N_4277);
nand U4547 (N_4547,N_4220,N_4361);
nand U4548 (N_4548,N_4351,N_4272);
or U4549 (N_4549,N_4332,N_4216);
xnor U4550 (N_4550,N_4291,N_4235);
xor U4551 (N_4551,N_4291,N_4224);
xnor U4552 (N_4552,N_4270,N_4364);
and U4553 (N_4553,N_4213,N_4358);
xor U4554 (N_4554,N_4370,N_4301);
nand U4555 (N_4555,N_4354,N_4393);
or U4556 (N_4556,N_4385,N_4249);
or U4557 (N_4557,N_4275,N_4254);
and U4558 (N_4558,N_4209,N_4329);
or U4559 (N_4559,N_4306,N_4367);
nand U4560 (N_4560,N_4373,N_4259);
xnor U4561 (N_4561,N_4259,N_4258);
xnor U4562 (N_4562,N_4394,N_4340);
or U4563 (N_4563,N_4224,N_4280);
xnor U4564 (N_4564,N_4323,N_4393);
nor U4565 (N_4565,N_4226,N_4270);
nand U4566 (N_4566,N_4365,N_4236);
nand U4567 (N_4567,N_4270,N_4370);
nand U4568 (N_4568,N_4365,N_4331);
xnor U4569 (N_4569,N_4396,N_4286);
and U4570 (N_4570,N_4308,N_4316);
or U4571 (N_4571,N_4248,N_4399);
xor U4572 (N_4572,N_4248,N_4327);
or U4573 (N_4573,N_4202,N_4295);
nor U4574 (N_4574,N_4341,N_4256);
and U4575 (N_4575,N_4360,N_4275);
xnor U4576 (N_4576,N_4390,N_4365);
xnor U4577 (N_4577,N_4379,N_4225);
or U4578 (N_4578,N_4266,N_4313);
nand U4579 (N_4579,N_4266,N_4237);
nand U4580 (N_4580,N_4312,N_4366);
or U4581 (N_4581,N_4285,N_4239);
nor U4582 (N_4582,N_4370,N_4348);
and U4583 (N_4583,N_4205,N_4258);
nor U4584 (N_4584,N_4227,N_4225);
or U4585 (N_4585,N_4332,N_4374);
or U4586 (N_4586,N_4285,N_4221);
or U4587 (N_4587,N_4320,N_4262);
or U4588 (N_4588,N_4397,N_4364);
xnor U4589 (N_4589,N_4263,N_4322);
nand U4590 (N_4590,N_4236,N_4397);
or U4591 (N_4591,N_4375,N_4396);
xnor U4592 (N_4592,N_4250,N_4355);
xor U4593 (N_4593,N_4342,N_4390);
nand U4594 (N_4594,N_4238,N_4265);
and U4595 (N_4595,N_4298,N_4206);
xnor U4596 (N_4596,N_4270,N_4210);
or U4597 (N_4597,N_4399,N_4282);
xnor U4598 (N_4598,N_4283,N_4218);
xnor U4599 (N_4599,N_4294,N_4321);
nor U4600 (N_4600,N_4511,N_4508);
or U4601 (N_4601,N_4524,N_4514);
nand U4602 (N_4602,N_4448,N_4450);
xor U4603 (N_4603,N_4539,N_4517);
nor U4604 (N_4604,N_4500,N_4575);
nor U4605 (N_4605,N_4540,N_4556);
nor U4606 (N_4606,N_4522,N_4446);
or U4607 (N_4607,N_4597,N_4592);
xor U4608 (N_4608,N_4461,N_4553);
and U4609 (N_4609,N_4568,N_4590);
and U4610 (N_4610,N_4585,N_4530);
nand U4611 (N_4611,N_4431,N_4579);
nor U4612 (N_4612,N_4510,N_4596);
and U4613 (N_4613,N_4422,N_4523);
xor U4614 (N_4614,N_4456,N_4440);
xnor U4615 (N_4615,N_4488,N_4407);
and U4616 (N_4616,N_4473,N_4430);
nand U4617 (N_4617,N_4462,N_4416);
and U4618 (N_4618,N_4413,N_4476);
nor U4619 (N_4619,N_4546,N_4464);
xnor U4620 (N_4620,N_4496,N_4576);
or U4621 (N_4621,N_4454,N_4519);
nand U4622 (N_4622,N_4563,N_4435);
nand U4623 (N_4623,N_4534,N_4402);
or U4624 (N_4624,N_4483,N_4509);
and U4625 (N_4625,N_4417,N_4533);
nand U4626 (N_4626,N_4518,N_4437);
nand U4627 (N_4627,N_4588,N_4542);
xnor U4628 (N_4628,N_4529,N_4512);
xnor U4629 (N_4629,N_4506,N_4475);
or U4630 (N_4630,N_4544,N_4598);
nand U4631 (N_4631,N_4498,N_4423);
xor U4632 (N_4632,N_4559,N_4557);
nor U4633 (N_4633,N_4513,N_4482);
or U4634 (N_4634,N_4583,N_4494);
nand U4635 (N_4635,N_4418,N_4425);
xnor U4636 (N_4636,N_4562,N_4504);
nor U4637 (N_4637,N_4507,N_4442);
and U4638 (N_4638,N_4445,N_4554);
nor U4639 (N_4639,N_4444,N_4497);
xnor U4640 (N_4640,N_4502,N_4499);
and U4641 (N_4641,N_4532,N_4481);
nand U4642 (N_4642,N_4451,N_4549);
xnor U4643 (N_4643,N_4552,N_4571);
nand U4644 (N_4644,N_4426,N_4471);
xnor U4645 (N_4645,N_4587,N_4428);
nor U4646 (N_4646,N_4584,N_4538);
and U4647 (N_4647,N_4593,N_4468);
nand U4648 (N_4648,N_4566,N_4467);
or U4649 (N_4649,N_4480,N_4493);
and U4650 (N_4650,N_4531,N_4412);
nor U4651 (N_4651,N_4470,N_4420);
nor U4652 (N_4652,N_4515,N_4479);
xnor U4653 (N_4653,N_4561,N_4409);
and U4654 (N_4654,N_4457,N_4487);
nand U4655 (N_4655,N_4569,N_4536);
xor U4656 (N_4656,N_4453,N_4555);
or U4657 (N_4657,N_4469,N_4429);
xor U4658 (N_4658,N_4574,N_4403);
and U4659 (N_4659,N_4577,N_4564);
nand U4660 (N_4660,N_4406,N_4527);
and U4661 (N_4661,N_4492,N_4433);
and U4662 (N_4662,N_4581,N_4491);
nand U4663 (N_4663,N_4455,N_4572);
or U4664 (N_4664,N_4537,N_4541);
xor U4665 (N_4665,N_4567,N_4505);
xor U4666 (N_4666,N_4432,N_4419);
and U4667 (N_4667,N_4516,N_4438);
and U4668 (N_4668,N_4595,N_4408);
nand U4669 (N_4669,N_4565,N_4551);
xor U4670 (N_4670,N_4421,N_4415);
or U4671 (N_4671,N_4459,N_4452);
and U4672 (N_4672,N_4434,N_4449);
xnor U4673 (N_4673,N_4458,N_4543);
and U4674 (N_4674,N_4490,N_4460);
nor U4675 (N_4675,N_4547,N_4586);
nor U4676 (N_4676,N_4424,N_4526);
nand U4677 (N_4677,N_4443,N_4405);
xnor U4678 (N_4678,N_4580,N_4463);
nand U4679 (N_4679,N_4589,N_4525);
or U4680 (N_4680,N_4495,N_4548);
xor U4681 (N_4681,N_4439,N_4400);
xor U4682 (N_4682,N_4465,N_4472);
nor U4683 (N_4683,N_4521,N_4478);
nand U4684 (N_4684,N_4550,N_4582);
nand U4685 (N_4685,N_4591,N_4447);
or U4686 (N_4686,N_4578,N_4427);
and U4687 (N_4687,N_4436,N_4486);
nor U4688 (N_4688,N_4570,N_4401);
xor U4689 (N_4689,N_4485,N_4404);
nor U4690 (N_4690,N_4594,N_4501);
nand U4691 (N_4691,N_4484,N_4545);
and U4692 (N_4692,N_4520,N_4474);
or U4693 (N_4693,N_4503,N_4477);
nor U4694 (N_4694,N_4558,N_4528);
xor U4695 (N_4695,N_4535,N_4411);
and U4696 (N_4696,N_4441,N_4573);
and U4697 (N_4697,N_4466,N_4410);
xor U4698 (N_4698,N_4560,N_4599);
nand U4699 (N_4699,N_4489,N_4414);
nor U4700 (N_4700,N_4503,N_4507);
nor U4701 (N_4701,N_4517,N_4421);
nand U4702 (N_4702,N_4438,N_4559);
xnor U4703 (N_4703,N_4566,N_4454);
or U4704 (N_4704,N_4459,N_4548);
or U4705 (N_4705,N_4522,N_4496);
and U4706 (N_4706,N_4421,N_4486);
xor U4707 (N_4707,N_4499,N_4469);
nand U4708 (N_4708,N_4451,N_4571);
nand U4709 (N_4709,N_4548,N_4542);
nor U4710 (N_4710,N_4487,N_4465);
or U4711 (N_4711,N_4471,N_4502);
xor U4712 (N_4712,N_4426,N_4516);
or U4713 (N_4713,N_4574,N_4546);
and U4714 (N_4714,N_4411,N_4408);
nor U4715 (N_4715,N_4585,N_4502);
and U4716 (N_4716,N_4403,N_4442);
nand U4717 (N_4717,N_4428,N_4456);
xor U4718 (N_4718,N_4504,N_4436);
xor U4719 (N_4719,N_4426,N_4405);
and U4720 (N_4720,N_4460,N_4411);
or U4721 (N_4721,N_4516,N_4540);
nand U4722 (N_4722,N_4511,N_4464);
and U4723 (N_4723,N_4592,N_4494);
and U4724 (N_4724,N_4582,N_4401);
or U4725 (N_4725,N_4423,N_4410);
or U4726 (N_4726,N_4460,N_4552);
nor U4727 (N_4727,N_4572,N_4573);
nand U4728 (N_4728,N_4516,N_4564);
and U4729 (N_4729,N_4517,N_4503);
or U4730 (N_4730,N_4565,N_4486);
or U4731 (N_4731,N_4480,N_4573);
xor U4732 (N_4732,N_4435,N_4430);
nand U4733 (N_4733,N_4458,N_4487);
nand U4734 (N_4734,N_4589,N_4572);
and U4735 (N_4735,N_4554,N_4407);
and U4736 (N_4736,N_4436,N_4558);
nand U4737 (N_4737,N_4442,N_4436);
xor U4738 (N_4738,N_4526,N_4594);
and U4739 (N_4739,N_4534,N_4509);
xnor U4740 (N_4740,N_4530,N_4535);
and U4741 (N_4741,N_4460,N_4426);
nand U4742 (N_4742,N_4406,N_4452);
or U4743 (N_4743,N_4448,N_4487);
and U4744 (N_4744,N_4407,N_4453);
or U4745 (N_4745,N_4427,N_4400);
or U4746 (N_4746,N_4455,N_4439);
or U4747 (N_4747,N_4506,N_4505);
and U4748 (N_4748,N_4505,N_4410);
nand U4749 (N_4749,N_4553,N_4401);
or U4750 (N_4750,N_4489,N_4528);
and U4751 (N_4751,N_4427,N_4576);
xor U4752 (N_4752,N_4583,N_4417);
or U4753 (N_4753,N_4595,N_4427);
nand U4754 (N_4754,N_4509,N_4482);
nand U4755 (N_4755,N_4545,N_4571);
nor U4756 (N_4756,N_4568,N_4446);
nand U4757 (N_4757,N_4512,N_4489);
nand U4758 (N_4758,N_4501,N_4454);
nor U4759 (N_4759,N_4511,N_4433);
nand U4760 (N_4760,N_4588,N_4405);
nand U4761 (N_4761,N_4516,N_4462);
and U4762 (N_4762,N_4576,N_4545);
or U4763 (N_4763,N_4561,N_4594);
and U4764 (N_4764,N_4557,N_4505);
nor U4765 (N_4765,N_4555,N_4444);
nor U4766 (N_4766,N_4559,N_4479);
or U4767 (N_4767,N_4450,N_4426);
nor U4768 (N_4768,N_4428,N_4454);
nor U4769 (N_4769,N_4461,N_4438);
xnor U4770 (N_4770,N_4498,N_4512);
nand U4771 (N_4771,N_4595,N_4461);
xor U4772 (N_4772,N_4409,N_4590);
nor U4773 (N_4773,N_4485,N_4534);
nor U4774 (N_4774,N_4422,N_4411);
or U4775 (N_4775,N_4589,N_4524);
xor U4776 (N_4776,N_4594,N_4415);
nor U4777 (N_4777,N_4548,N_4577);
xor U4778 (N_4778,N_4528,N_4429);
nand U4779 (N_4779,N_4450,N_4475);
nand U4780 (N_4780,N_4461,N_4455);
nand U4781 (N_4781,N_4536,N_4416);
nand U4782 (N_4782,N_4574,N_4504);
xnor U4783 (N_4783,N_4487,N_4460);
nand U4784 (N_4784,N_4409,N_4430);
nor U4785 (N_4785,N_4578,N_4493);
or U4786 (N_4786,N_4529,N_4568);
xor U4787 (N_4787,N_4423,N_4552);
xor U4788 (N_4788,N_4471,N_4557);
and U4789 (N_4789,N_4427,N_4497);
and U4790 (N_4790,N_4510,N_4566);
nor U4791 (N_4791,N_4480,N_4422);
xnor U4792 (N_4792,N_4481,N_4544);
nor U4793 (N_4793,N_4510,N_4429);
nand U4794 (N_4794,N_4526,N_4522);
nand U4795 (N_4795,N_4583,N_4470);
and U4796 (N_4796,N_4475,N_4468);
and U4797 (N_4797,N_4441,N_4497);
or U4798 (N_4798,N_4587,N_4536);
or U4799 (N_4799,N_4526,N_4575);
or U4800 (N_4800,N_4639,N_4750);
nand U4801 (N_4801,N_4755,N_4737);
nand U4802 (N_4802,N_4766,N_4605);
nand U4803 (N_4803,N_4745,N_4619);
nand U4804 (N_4804,N_4759,N_4618);
and U4805 (N_4805,N_4716,N_4701);
nor U4806 (N_4806,N_4658,N_4747);
nand U4807 (N_4807,N_4652,N_4644);
nor U4808 (N_4808,N_4788,N_4706);
and U4809 (N_4809,N_4783,N_4698);
xor U4810 (N_4810,N_4715,N_4749);
and U4811 (N_4811,N_4743,N_4683);
nand U4812 (N_4812,N_4684,N_4682);
nor U4813 (N_4813,N_4611,N_4738);
nand U4814 (N_4814,N_4751,N_4795);
or U4815 (N_4815,N_4718,N_4625);
nor U4816 (N_4816,N_4774,N_4786);
nor U4817 (N_4817,N_4742,N_4664);
or U4818 (N_4818,N_4662,N_4672);
xor U4819 (N_4819,N_4707,N_4779);
nor U4820 (N_4820,N_4740,N_4656);
nand U4821 (N_4821,N_4635,N_4600);
and U4822 (N_4822,N_4627,N_4709);
nand U4823 (N_4823,N_4669,N_4686);
xnor U4824 (N_4824,N_4660,N_4726);
nor U4825 (N_4825,N_4687,N_4696);
or U4826 (N_4826,N_4612,N_4610);
nor U4827 (N_4827,N_4705,N_4633);
nand U4828 (N_4828,N_4675,N_4735);
and U4829 (N_4829,N_4665,N_4606);
and U4830 (N_4830,N_4704,N_4787);
or U4831 (N_4831,N_4777,N_4729);
or U4832 (N_4832,N_4648,N_4703);
nor U4833 (N_4833,N_4700,N_4650);
nor U4834 (N_4834,N_4799,N_4762);
or U4835 (N_4835,N_4720,N_4732);
nand U4836 (N_4836,N_4756,N_4671);
xor U4837 (N_4837,N_4722,N_4621);
or U4838 (N_4838,N_4632,N_4768);
and U4839 (N_4839,N_4731,N_4666);
or U4840 (N_4840,N_4736,N_4798);
and U4841 (N_4841,N_4630,N_4622);
nor U4842 (N_4842,N_4673,N_4661);
nand U4843 (N_4843,N_4782,N_4676);
xor U4844 (N_4844,N_4769,N_4746);
or U4845 (N_4845,N_4616,N_4670);
and U4846 (N_4846,N_4604,N_4629);
and U4847 (N_4847,N_4748,N_4699);
or U4848 (N_4848,N_4641,N_4636);
and U4849 (N_4849,N_4784,N_4744);
or U4850 (N_4850,N_4690,N_4758);
nor U4851 (N_4851,N_4711,N_4655);
or U4852 (N_4852,N_4695,N_4602);
nor U4853 (N_4853,N_4667,N_4725);
nor U4854 (N_4854,N_4617,N_4753);
nor U4855 (N_4855,N_4772,N_4754);
nand U4856 (N_4856,N_4790,N_4674);
xor U4857 (N_4857,N_4668,N_4789);
nand U4858 (N_4858,N_4717,N_4734);
nor U4859 (N_4859,N_4603,N_4614);
nand U4860 (N_4860,N_4647,N_4776);
nand U4861 (N_4861,N_4792,N_4757);
xnor U4862 (N_4862,N_4767,N_4781);
nand U4863 (N_4863,N_4773,N_4724);
nand U4864 (N_4864,N_4663,N_4733);
xor U4865 (N_4865,N_4728,N_4739);
or U4866 (N_4866,N_4723,N_4638);
and U4867 (N_4867,N_4693,N_4719);
xnor U4868 (N_4868,N_4761,N_4714);
or U4869 (N_4869,N_4626,N_4679);
xnor U4870 (N_4870,N_4691,N_4797);
nand U4871 (N_4871,N_4688,N_4642);
and U4872 (N_4872,N_4609,N_4794);
or U4873 (N_4873,N_4615,N_4624);
and U4874 (N_4874,N_4710,N_4694);
nor U4875 (N_4875,N_4681,N_4791);
xnor U4876 (N_4876,N_4730,N_4763);
nand U4877 (N_4877,N_4771,N_4678);
nand U4878 (N_4878,N_4780,N_4727);
and U4879 (N_4879,N_4640,N_4775);
and U4880 (N_4880,N_4692,N_4637);
and U4881 (N_4881,N_4628,N_4643);
or U4882 (N_4882,N_4631,N_4765);
and U4883 (N_4883,N_4796,N_4741);
nand U4884 (N_4884,N_4601,N_4689);
xor U4885 (N_4885,N_4764,N_4712);
nor U4886 (N_4886,N_4645,N_4634);
nor U4887 (N_4887,N_4651,N_4607);
or U4888 (N_4888,N_4702,N_4653);
and U4889 (N_4889,N_4620,N_4697);
nor U4890 (N_4890,N_4785,N_4654);
nand U4891 (N_4891,N_4760,N_4646);
xnor U4892 (N_4892,N_4778,N_4721);
nor U4893 (N_4893,N_4657,N_4770);
nand U4894 (N_4894,N_4613,N_4793);
xor U4895 (N_4895,N_4713,N_4708);
xnor U4896 (N_4896,N_4608,N_4623);
nor U4897 (N_4897,N_4659,N_4680);
and U4898 (N_4898,N_4752,N_4685);
and U4899 (N_4899,N_4677,N_4649);
and U4900 (N_4900,N_4639,N_4699);
xnor U4901 (N_4901,N_4716,N_4702);
xor U4902 (N_4902,N_4698,N_4776);
nand U4903 (N_4903,N_4627,N_4774);
nand U4904 (N_4904,N_4737,N_4739);
nor U4905 (N_4905,N_4719,N_4705);
xor U4906 (N_4906,N_4655,N_4680);
nand U4907 (N_4907,N_4710,N_4775);
or U4908 (N_4908,N_4787,N_4625);
and U4909 (N_4909,N_4737,N_4793);
nor U4910 (N_4910,N_4697,N_4611);
nand U4911 (N_4911,N_4668,N_4734);
or U4912 (N_4912,N_4736,N_4668);
and U4913 (N_4913,N_4783,N_4786);
and U4914 (N_4914,N_4736,N_4635);
nand U4915 (N_4915,N_4729,N_4738);
nor U4916 (N_4916,N_4763,N_4765);
nor U4917 (N_4917,N_4768,N_4728);
and U4918 (N_4918,N_4665,N_4763);
and U4919 (N_4919,N_4736,N_4715);
nand U4920 (N_4920,N_4643,N_4750);
and U4921 (N_4921,N_4797,N_4710);
xor U4922 (N_4922,N_4732,N_4660);
nand U4923 (N_4923,N_4614,N_4706);
and U4924 (N_4924,N_4707,N_4758);
nor U4925 (N_4925,N_4746,N_4641);
nor U4926 (N_4926,N_4688,N_4681);
xor U4927 (N_4927,N_4714,N_4671);
or U4928 (N_4928,N_4755,N_4638);
and U4929 (N_4929,N_4757,N_4600);
nor U4930 (N_4930,N_4711,N_4606);
or U4931 (N_4931,N_4732,N_4711);
nand U4932 (N_4932,N_4718,N_4775);
xnor U4933 (N_4933,N_4666,N_4732);
and U4934 (N_4934,N_4636,N_4689);
and U4935 (N_4935,N_4734,N_4639);
or U4936 (N_4936,N_4747,N_4702);
and U4937 (N_4937,N_4773,N_4772);
nand U4938 (N_4938,N_4680,N_4698);
xor U4939 (N_4939,N_4786,N_4731);
nor U4940 (N_4940,N_4638,N_4657);
nor U4941 (N_4941,N_4717,N_4792);
xor U4942 (N_4942,N_4652,N_4647);
or U4943 (N_4943,N_4737,N_4649);
or U4944 (N_4944,N_4632,N_4789);
nor U4945 (N_4945,N_4730,N_4665);
and U4946 (N_4946,N_4771,N_4674);
xor U4947 (N_4947,N_4613,N_4674);
and U4948 (N_4948,N_4765,N_4788);
nor U4949 (N_4949,N_4688,N_4620);
nand U4950 (N_4950,N_4701,N_4695);
and U4951 (N_4951,N_4701,N_4730);
nand U4952 (N_4952,N_4770,N_4742);
xor U4953 (N_4953,N_4693,N_4782);
or U4954 (N_4954,N_4643,N_4687);
nand U4955 (N_4955,N_4643,N_4723);
xnor U4956 (N_4956,N_4658,N_4678);
or U4957 (N_4957,N_4785,N_4601);
xnor U4958 (N_4958,N_4707,N_4775);
nor U4959 (N_4959,N_4782,N_4667);
or U4960 (N_4960,N_4637,N_4781);
and U4961 (N_4961,N_4603,N_4711);
and U4962 (N_4962,N_4627,N_4732);
and U4963 (N_4963,N_4775,N_4749);
nor U4964 (N_4964,N_4753,N_4717);
nand U4965 (N_4965,N_4698,N_4613);
or U4966 (N_4966,N_4628,N_4716);
xnor U4967 (N_4967,N_4793,N_4741);
and U4968 (N_4968,N_4679,N_4701);
and U4969 (N_4969,N_4609,N_4783);
xnor U4970 (N_4970,N_4791,N_4700);
nor U4971 (N_4971,N_4663,N_4744);
and U4972 (N_4972,N_4642,N_4691);
or U4973 (N_4973,N_4706,N_4787);
or U4974 (N_4974,N_4774,N_4676);
xnor U4975 (N_4975,N_4703,N_4673);
and U4976 (N_4976,N_4698,N_4630);
xnor U4977 (N_4977,N_4602,N_4606);
or U4978 (N_4978,N_4705,N_4781);
nand U4979 (N_4979,N_4659,N_4628);
xor U4980 (N_4980,N_4608,N_4729);
nand U4981 (N_4981,N_4671,N_4611);
xor U4982 (N_4982,N_4630,N_4636);
xor U4983 (N_4983,N_4680,N_4692);
nor U4984 (N_4984,N_4778,N_4616);
xnor U4985 (N_4985,N_4608,N_4624);
nor U4986 (N_4986,N_4624,N_4720);
nor U4987 (N_4987,N_4735,N_4707);
nor U4988 (N_4988,N_4608,N_4765);
nor U4989 (N_4989,N_4690,N_4789);
nand U4990 (N_4990,N_4681,N_4795);
nand U4991 (N_4991,N_4606,N_4642);
nor U4992 (N_4992,N_4610,N_4782);
or U4993 (N_4993,N_4794,N_4688);
xor U4994 (N_4994,N_4771,N_4689);
nor U4995 (N_4995,N_4647,N_4724);
and U4996 (N_4996,N_4764,N_4732);
nand U4997 (N_4997,N_4624,N_4768);
nand U4998 (N_4998,N_4758,N_4714);
and U4999 (N_4999,N_4710,N_4640);
and U5000 (N_5000,N_4930,N_4989);
and U5001 (N_5001,N_4941,N_4949);
nand U5002 (N_5002,N_4819,N_4999);
or U5003 (N_5003,N_4905,N_4836);
xnor U5004 (N_5004,N_4982,N_4957);
or U5005 (N_5005,N_4943,N_4938);
nand U5006 (N_5006,N_4914,N_4812);
or U5007 (N_5007,N_4968,N_4820);
and U5008 (N_5008,N_4903,N_4811);
nand U5009 (N_5009,N_4961,N_4804);
and U5010 (N_5010,N_4986,N_4893);
and U5011 (N_5011,N_4996,N_4976);
nor U5012 (N_5012,N_4925,N_4880);
xor U5013 (N_5013,N_4921,N_4829);
or U5014 (N_5014,N_4908,N_4975);
nor U5015 (N_5015,N_4869,N_4826);
nand U5016 (N_5016,N_4840,N_4870);
xor U5017 (N_5017,N_4823,N_4853);
nand U5018 (N_5018,N_4966,N_4886);
nor U5019 (N_5019,N_4931,N_4877);
nand U5020 (N_5020,N_4848,N_4808);
and U5021 (N_5021,N_4858,N_4912);
and U5022 (N_5022,N_4841,N_4906);
xor U5023 (N_5023,N_4810,N_4958);
and U5024 (N_5024,N_4834,N_4932);
xor U5025 (N_5025,N_4860,N_4969);
nor U5026 (N_5026,N_4970,N_4828);
and U5027 (N_5027,N_4872,N_4951);
and U5028 (N_5028,N_4851,N_4861);
nand U5029 (N_5029,N_4990,N_4801);
xor U5030 (N_5030,N_4881,N_4822);
nand U5031 (N_5031,N_4807,N_4991);
and U5032 (N_5032,N_4824,N_4890);
or U5033 (N_5033,N_4821,N_4850);
nor U5034 (N_5034,N_4902,N_4898);
nand U5035 (N_5035,N_4907,N_4948);
xnor U5036 (N_5036,N_4887,N_4827);
nand U5037 (N_5037,N_4899,N_4981);
nor U5038 (N_5038,N_4814,N_4998);
or U5039 (N_5039,N_4967,N_4972);
nor U5040 (N_5040,N_4945,N_4875);
xnor U5041 (N_5041,N_4842,N_4947);
or U5042 (N_5042,N_4847,N_4953);
xor U5043 (N_5043,N_4960,N_4876);
or U5044 (N_5044,N_4984,N_4865);
nor U5045 (N_5045,N_4816,N_4964);
nand U5046 (N_5046,N_4918,N_4885);
or U5047 (N_5047,N_4985,N_4963);
xnor U5048 (N_5048,N_4825,N_4916);
nor U5049 (N_5049,N_4896,N_4855);
or U5050 (N_5050,N_4874,N_4978);
xor U5051 (N_5051,N_4956,N_4959);
nand U5052 (N_5052,N_4838,N_4813);
and U5053 (N_5053,N_4944,N_4864);
nand U5054 (N_5054,N_4892,N_4927);
nor U5055 (N_5055,N_4913,N_4936);
and U5056 (N_5056,N_4909,N_4805);
and U5057 (N_5057,N_4974,N_4849);
xor U5058 (N_5058,N_4950,N_4800);
nor U5059 (N_5059,N_4915,N_4933);
or U5060 (N_5060,N_4809,N_4929);
nor U5061 (N_5061,N_4983,N_4926);
nor U5062 (N_5062,N_4979,N_4866);
nor U5063 (N_5063,N_4854,N_4802);
xnor U5064 (N_5064,N_4894,N_4862);
nor U5065 (N_5065,N_4856,N_4987);
xor U5066 (N_5066,N_4837,N_4901);
and U5067 (N_5067,N_4844,N_4971);
or U5068 (N_5068,N_4928,N_4859);
nor U5069 (N_5069,N_4965,N_4817);
and U5070 (N_5070,N_4884,N_4845);
and U5071 (N_5071,N_4911,N_4993);
and U5072 (N_5072,N_4883,N_4934);
nor U5073 (N_5073,N_4833,N_4910);
nand U5074 (N_5074,N_4839,N_4803);
xor U5075 (N_5075,N_4924,N_4873);
and U5076 (N_5076,N_4846,N_4857);
nand U5077 (N_5077,N_4806,N_4878);
or U5078 (N_5078,N_4897,N_4900);
or U5079 (N_5079,N_4852,N_4888);
nor U5080 (N_5080,N_4917,N_4997);
nand U5081 (N_5081,N_4843,N_4994);
nand U5082 (N_5082,N_4992,N_4835);
or U5083 (N_5083,N_4879,N_4923);
nor U5084 (N_5084,N_4935,N_4863);
or U5085 (N_5085,N_4868,N_4871);
nand U5086 (N_5086,N_4973,N_4920);
nor U5087 (N_5087,N_4940,N_4988);
and U5088 (N_5088,N_4831,N_4946);
xor U5089 (N_5089,N_4937,N_4818);
xor U5090 (N_5090,N_4995,N_4939);
or U5091 (N_5091,N_4832,N_4895);
or U5092 (N_5092,N_4952,N_4922);
and U5093 (N_5093,N_4980,N_4962);
and U5094 (N_5094,N_4942,N_4889);
or U5095 (N_5095,N_4867,N_4891);
or U5096 (N_5096,N_4954,N_4815);
xor U5097 (N_5097,N_4882,N_4955);
nand U5098 (N_5098,N_4919,N_4830);
or U5099 (N_5099,N_4977,N_4904);
xor U5100 (N_5100,N_4929,N_4919);
and U5101 (N_5101,N_4867,N_4808);
or U5102 (N_5102,N_4831,N_4820);
nand U5103 (N_5103,N_4844,N_4847);
nor U5104 (N_5104,N_4880,N_4989);
nor U5105 (N_5105,N_4903,N_4931);
xor U5106 (N_5106,N_4952,N_4921);
or U5107 (N_5107,N_4946,N_4852);
or U5108 (N_5108,N_4815,N_4973);
nand U5109 (N_5109,N_4860,N_4989);
and U5110 (N_5110,N_4837,N_4806);
xnor U5111 (N_5111,N_4908,N_4946);
and U5112 (N_5112,N_4834,N_4805);
or U5113 (N_5113,N_4817,N_4885);
xnor U5114 (N_5114,N_4914,N_4830);
and U5115 (N_5115,N_4813,N_4823);
nor U5116 (N_5116,N_4800,N_4905);
and U5117 (N_5117,N_4940,N_4879);
and U5118 (N_5118,N_4811,N_4992);
xor U5119 (N_5119,N_4875,N_4963);
xnor U5120 (N_5120,N_4805,N_4986);
or U5121 (N_5121,N_4903,N_4999);
nand U5122 (N_5122,N_4968,N_4840);
nor U5123 (N_5123,N_4908,N_4907);
nand U5124 (N_5124,N_4810,N_4970);
nor U5125 (N_5125,N_4993,N_4964);
nand U5126 (N_5126,N_4919,N_4913);
xnor U5127 (N_5127,N_4994,N_4803);
or U5128 (N_5128,N_4941,N_4972);
nand U5129 (N_5129,N_4970,N_4808);
nor U5130 (N_5130,N_4961,N_4946);
nand U5131 (N_5131,N_4902,N_4886);
xor U5132 (N_5132,N_4860,N_4818);
xnor U5133 (N_5133,N_4972,N_4813);
and U5134 (N_5134,N_4846,N_4901);
nand U5135 (N_5135,N_4895,N_4811);
xor U5136 (N_5136,N_4952,N_4888);
and U5137 (N_5137,N_4817,N_4922);
nand U5138 (N_5138,N_4937,N_4944);
nor U5139 (N_5139,N_4808,N_4922);
xor U5140 (N_5140,N_4922,N_4893);
and U5141 (N_5141,N_4844,N_4988);
nor U5142 (N_5142,N_4866,N_4801);
xnor U5143 (N_5143,N_4984,N_4814);
nor U5144 (N_5144,N_4854,N_4839);
or U5145 (N_5145,N_4883,N_4991);
or U5146 (N_5146,N_4867,N_4890);
and U5147 (N_5147,N_4996,N_4901);
nor U5148 (N_5148,N_4922,N_4906);
nor U5149 (N_5149,N_4921,N_4869);
xnor U5150 (N_5150,N_4955,N_4874);
or U5151 (N_5151,N_4835,N_4975);
and U5152 (N_5152,N_4961,N_4864);
and U5153 (N_5153,N_4895,N_4817);
and U5154 (N_5154,N_4963,N_4836);
nand U5155 (N_5155,N_4875,N_4865);
nand U5156 (N_5156,N_4906,N_4961);
or U5157 (N_5157,N_4833,N_4951);
nor U5158 (N_5158,N_4972,N_4832);
or U5159 (N_5159,N_4843,N_4887);
and U5160 (N_5160,N_4948,N_4979);
nor U5161 (N_5161,N_4800,N_4856);
or U5162 (N_5162,N_4852,N_4816);
and U5163 (N_5163,N_4968,N_4828);
nand U5164 (N_5164,N_4922,N_4899);
or U5165 (N_5165,N_4838,N_4870);
and U5166 (N_5166,N_4883,N_4846);
nor U5167 (N_5167,N_4841,N_4947);
nor U5168 (N_5168,N_4836,N_4840);
nand U5169 (N_5169,N_4853,N_4935);
nand U5170 (N_5170,N_4929,N_4942);
nor U5171 (N_5171,N_4854,N_4908);
xnor U5172 (N_5172,N_4937,N_4819);
xnor U5173 (N_5173,N_4883,N_4881);
or U5174 (N_5174,N_4949,N_4984);
xnor U5175 (N_5175,N_4874,N_4998);
nand U5176 (N_5176,N_4922,N_4835);
nor U5177 (N_5177,N_4820,N_4971);
or U5178 (N_5178,N_4938,N_4961);
nand U5179 (N_5179,N_4905,N_4810);
and U5180 (N_5180,N_4927,N_4893);
xor U5181 (N_5181,N_4939,N_4893);
xnor U5182 (N_5182,N_4859,N_4851);
and U5183 (N_5183,N_4835,N_4801);
xor U5184 (N_5184,N_4994,N_4955);
or U5185 (N_5185,N_4833,N_4911);
or U5186 (N_5186,N_4812,N_4889);
xnor U5187 (N_5187,N_4867,N_4970);
xor U5188 (N_5188,N_4858,N_4902);
or U5189 (N_5189,N_4851,N_4941);
xnor U5190 (N_5190,N_4810,N_4800);
nor U5191 (N_5191,N_4892,N_4876);
nor U5192 (N_5192,N_4953,N_4996);
nor U5193 (N_5193,N_4921,N_4839);
and U5194 (N_5194,N_4914,N_4833);
xor U5195 (N_5195,N_4848,N_4917);
nor U5196 (N_5196,N_4942,N_4947);
nand U5197 (N_5197,N_4846,N_4899);
xnor U5198 (N_5198,N_4891,N_4935);
and U5199 (N_5199,N_4808,N_4991);
and U5200 (N_5200,N_5116,N_5068);
and U5201 (N_5201,N_5158,N_5033);
and U5202 (N_5202,N_5041,N_5069);
nand U5203 (N_5203,N_5059,N_5018);
nand U5204 (N_5204,N_5067,N_5038);
or U5205 (N_5205,N_5137,N_5133);
and U5206 (N_5206,N_5156,N_5026);
nand U5207 (N_5207,N_5003,N_5019);
xnor U5208 (N_5208,N_5085,N_5110);
and U5209 (N_5209,N_5090,N_5170);
nor U5210 (N_5210,N_5095,N_5056);
and U5211 (N_5211,N_5187,N_5050);
or U5212 (N_5212,N_5124,N_5051);
xnor U5213 (N_5213,N_5125,N_5005);
nor U5214 (N_5214,N_5149,N_5055);
nor U5215 (N_5215,N_5064,N_5163);
and U5216 (N_5216,N_5081,N_5130);
or U5217 (N_5217,N_5189,N_5101);
and U5218 (N_5218,N_5084,N_5058);
and U5219 (N_5219,N_5103,N_5034);
or U5220 (N_5220,N_5045,N_5159);
nor U5221 (N_5221,N_5169,N_5086);
and U5222 (N_5222,N_5111,N_5177);
and U5223 (N_5223,N_5166,N_5148);
nand U5224 (N_5224,N_5127,N_5009);
xnor U5225 (N_5225,N_5087,N_5185);
nor U5226 (N_5226,N_5001,N_5036);
and U5227 (N_5227,N_5126,N_5021);
nor U5228 (N_5228,N_5164,N_5198);
nor U5229 (N_5229,N_5151,N_5175);
xnor U5230 (N_5230,N_5176,N_5165);
and U5231 (N_5231,N_5012,N_5117);
nor U5232 (N_5232,N_5154,N_5102);
and U5233 (N_5233,N_5020,N_5048);
nand U5234 (N_5234,N_5007,N_5061);
nor U5235 (N_5235,N_5071,N_5035);
nand U5236 (N_5236,N_5023,N_5104);
and U5237 (N_5237,N_5186,N_5112);
or U5238 (N_5238,N_5161,N_5171);
nand U5239 (N_5239,N_5053,N_5062);
nand U5240 (N_5240,N_5047,N_5132);
nor U5241 (N_5241,N_5180,N_5093);
nand U5242 (N_5242,N_5178,N_5162);
xnor U5243 (N_5243,N_5192,N_5140);
nor U5244 (N_5244,N_5190,N_5022);
or U5245 (N_5245,N_5136,N_5076);
and U5246 (N_5246,N_5083,N_5088);
nor U5247 (N_5247,N_5197,N_5098);
nand U5248 (N_5248,N_5160,N_5072);
xnor U5249 (N_5249,N_5194,N_5153);
nand U5250 (N_5250,N_5031,N_5167);
nor U5251 (N_5251,N_5078,N_5075);
or U5252 (N_5252,N_5006,N_5029);
xnor U5253 (N_5253,N_5129,N_5106);
xnor U5254 (N_5254,N_5183,N_5040);
or U5255 (N_5255,N_5131,N_5115);
xor U5256 (N_5256,N_5063,N_5042);
or U5257 (N_5257,N_5191,N_5077);
and U5258 (N_5258,N_5168,N_5016);
nor U5259 (N_5259,N_5173,N_5179);
and U5260 (N_5260,N_5028,N_5066);
or U5261 (N_5261,N_5139,N_5013);
or U5262 (N_5262,N_5172,N_5134);
and U5263 (N_5263,N_5123,N_5024);
nand U5264 (N_5264,N_5120,N_5025);
xor U5265 (N_5265,N_5152,N_5195);
nand U5266 (N_5266,N_5017,N_5182);
and U5267 (N_5267,N_5119,N_5004);
nand U5268 (N_5268,N_5135,N_5054);
nand U5269 (N_5269,N_5107,N_5030);
xnor U5270 (N_5270,N_5089,N_5015);
or U5271 (N_5271,N_5144,N_5188);
xnor U5272 (N_5272,N_5027,N_5060);
or U5273 (N_5273,N_5150,N_5097);
or U5274 (N_5274,N_5109,N_5141);
nor U5275 (N_5275,N_5091,N_5199);
and U5276 (N_5276,N_5002,N_5128);
xnor U5277 (N_5277,N_5157,N_5065);
or U5278 (N_5278,N_5105,N_5184);
nand U5279 (N_5279,N_5147,N_5108);
xnor U5280 (N_5280,N_5174,N_5080);
nand U5281 (N_5281,N_5014,N_5049);
and U5282 (N_5282,N_5196,N_5092);
and U5283 (N_5283,N_5057,N_5011);
and U5284 (N_5284,N_5113,N_5138);
nor U5285 (N_5285,N_5046,N_5073);
nand U5286 (N_5286,N_5043,N_5037);
nand U5287 (N_5287,N_5099,N_5082);
nand U5288 (N_5288,N_5070,N_5118);
nor U5289 (N_5289,N_5143,N_5096);
and U5290 (N_5290,N_5079,N_5142);
nand U5291 (N_5291,N_5155,N_5008);
nor U5292 (N_5292,N_5193,N_5052);
or U5293 (N_5293,N_5094,N_5074);
xor U5294 (N_5294,N_5181,N_5010);
nor U5295 (N_5295,N_5044,N_5039);
nand U5296 (N_5296,N_5146,N_5114);
nor U5297 (N_5297,N_5121,N_5032);
and U5298 (N_5298,N_5000,N_5100);
xor U5299 (N_5299,N_5145,N_5122);
nand U5300 (N_5300,N_5046,N_5103);
and U5301 (N_5301,N_5184,N_5194);
nor U5302 (N_5302,N_5117,N_5045);
nor U5303 (N_5303,N_5100,N_5056);
or U5304 (N_5304,N_5086,N_5107);
and U5305 (N_5305,N_5047,N_5126);
or U5306 (N_5306,N_5131,N_5055);
and U5307 (N_5307,N_5066,N_5152);
or U5308 (N_5308,N_5158,N_5078);
xnor U5309 (N_5309,N_5078,N_5195);
xor U5310 (N_5310,N_5062,N_5105);
nand U5311 (N_5311,N_5088,N_5058);
and U5312 (N_5312,N_5081,N_5146);
or U5313 (N_5313,N_5050,N_5126);
and U5314 (N_5314,N_5057,N_5135);
or U5315 (N_5315,N_5059,N_5185);
nand U5316 (N_5316,N_5106,N_5171);
xnor U5317 (N_5317,N_5090,N_5087);
xor U5318 (N_5318,N_5078,N_5197);
or U5319 (N_5319,N_5168,N_5174);
or U5320 (N_5320,N_5168,N_5031);
and U5321 (N_5321,N_5120,N_5170);
nor U5322 (N_5322,N_5137,N_5169);
xnor U5323 (N_5323,N_5066,N_5149);
or U5324 (N_5324,N_5169,N_5185);
and U5325 (N_5325,N_5092,N_5138);
or U5326 (N_5326,N_5148,N_5103);
xor U5327 (N_5327,N_5172,N_5033);
nor U5328 (N_5328,N_5053,N_5035);
and U5329 (N_5329,N_5019,N_5121);
nand U5330 (N_5330,N_5174,N_5114);
xnor U5331 (N_5331,N_5055,N_5198);
or U5332 (N_5332,N_5016,N_5158);
nor U5333 (N_5333,N_5199,N_5195);
nor U5334 (N_5334,N_5160,N_5099);
and U5335 (N_5335,N_5108,N_5120);
and U5336 (N_5336,N_5173,N_5079);
nor U5337 (N_5337,N_5051,N_5022);
nor U5338 (N_5338,N_5101,N_5055);
xor U5339 (N_5339,N_5076,N_5120);
xnor U5340 (N_5340,N_5038,N_5045);
xor U5341 (N_5341,N_5163,N_5052);
xor U5342 (N_5342,N_5073,N_5189);
nor U5343 (N_5343,N_5113,N_5055);
xnor U5344 (N_5344,N_5166,N_5178);
nor U5345 (N_5345,N_5118,N_5007);
or U5346 (N_5346,N_5081,N_5127);
and U5347 (N_5347,N_5065,N_5003);
or U5348 (N_5348,N_5095,N_5082);
xnor U5349 (N_5349,N_5108,N_5151);
or U5350 (N_5350,N_5061,N_5067);
and U5351 (N_5351,N_5065,N_5025);
nor U5352 (N_5352,N_5188,N_5184);
nand U5353 (N_5353,N_5044,N_5046);
xnor U5354 (N_5354,N_5045,N_5198);
and U5355 (N_5355,N_5052,N_5140);
and U5356 (N_5356,N_5195,N_5052);
and U5357 (N_5357,N_5049,N_5031);
nand U5358 (N_5358,N_5169,N_5112);
and U5359 (N_5359,N_5137,N_5184);
and U5360 (N_5360,N_5062,N_5006);
xor U5361 (N_5361,N_5016,N_5061);
or U5362 (N_5362,N_5056,N_5027);
nor U5363 (N_5363,N_5076,N_5132);
nand U5364 (N_5364,N_5188,N_5164);
nand U5365 (N_5365,N_5088,N_5077);
xor U5366 (N_5366,N_5126,N_5057);
or U5367 (N_5367,N_5100,N_5151);
nor U5368 (N_5368,N_5065,N_5060);
nand U5369 (N_5369,N_5183,N_5029);
nand U5370 (N_5370,N_5043,N_5054);
and U5371 (N_5371,N_5092,N_5014);
and U5372 (N_5372,N_5092,N_5100);
or U5373 (N_5373,N_5108,N_5095);
xnor U5374 (N_5374,N_5024,N_5197);
xor U5375 (N_5375,N_5109,N_5000);
xnor U5376 (N_5376,N_5052,N_5018);
and U5377 (N_5377,N_5064,N_5113);
nand U5378 (N_5378,N_5095,N_5077);
and U5379 (N_5379,N_5098,N_5015);
xnor U5380 (N_5380,N_5011,N_5141);
and U5381 (N_5381,N_5126,N_5124);
and U5382 (N_5382,N_5189,N_5143);
nand U5383 (N_5383,N_5120,N_5107);
nor U5384 (N_5384,N_5122,N_5030);
and U5385 (N_5385,N_5057,N_5075);
xor U5386 (N_5386,N_5131,N_5192);
and U5387 (N_5387,N_5073,N_5178);
xor U5388 (N_5388,N_5066,N_5164);
nor U5389 (N_5389,N_5019,N_5105);
xnor U5390 (N_5390,N_5093,N_5142);
or U5391 (N_5391,N_5001,N_5045);
or U5392 (N_5392,N_5052,N_5016);
nor U5393 (N_5393,N_5031,N_5033);
or U5394 (N_5394,N_5161,N_5053);
or U5395 (N_5395,N_5178,N_5159);
and U5396 (N_5396,N_5049,N_5165);
and U5397 (N_5397,N_5041,N_5159);
xnor U5398 (N_5398,N_5123,N_5036);
nor U5399 (N_5399,N_5033,N_5117);
nor U5400 (N_5400,N_5245,N_5264);
nor U5401 (N_5401,N_5395,N_5385);
or U5402 (N_5402,N_5361,N_5282);
xnor U5403 (N_5403,N_5301,N_5340);
nand U5404 (N_5404,N_5311,N_5278);
xor U5405 (N_5405,N_5242,N_5371);
xor U5406 (N_5406,N_5201,N_5397);
xor U5407 (N_5407,N_5271,N_5359);
nand U5408 (N_5408,N_5347,N_5336);
and U5409 (N_5409,N_5226,N_5374);
xnor U5410 (N_5410,N_5341,N_5253);
nor U5411 (N_5411,N_5356,N_5383);
xnor U5412 (N_5412,N_5288,N_5273);
and U5413 (N_5413,N_5332,N_5258);
xor U5414 (N_5414,N_5286,N_5346);
xnor U5415 (N_5415,N_5318,N_5276);
nand U5416 (N_5416,N_5297,N_5229);
xor U5417 (N_5417,N_5367,N_5215);
or U5418 (N_5418,N_5207,N_5339);
or U5419 (N_5419,N_5211,N_5390);
xor U5420 (N_5420,N_5254,N_5274);
and U5421 (N_5421,N_5335,N_5302);
or U5422 (N_5422,N_5261,N_5265);
xnor U5423 (N_5423,N_5272,N_5322);
nand U5424 (N_5424,N_5376,N_5369);
nor U5425 (N_5425,N_5257,N_5355);
xor U5426 (N_5426,N_5352,N_5398);
and U5427 (N_5427,N_5219,N_5364);
and U5428 (N_5428,N_5217,N_5260);
xnor U5429 (N_5429,N_5357,N_5218);
or U5430 (N_5430,N_5314,N_5263);
nor U5431 (N_5431,N_5391,N_5227);
xnor U5432 (N_5432,N_5238,N_5377);
nand U5433 (N_5433,N_5360,N_5208);
xnor U5434 (N_5434,N_5350,N_5247);
or U5435 (N_5435,N_5354,N_5331);
nand U5436 (N_5436,N_5380,N_5241);
nor U5437 (N_5437,N_5204,N_5329);
nand U5438 (N_5438,N_5303,N_5366);
or U5439 (N_5439,N_5345,N_5285);
nand U5440 (N_5440,N_5333,N_5232);
nand U5441 (N_5441,N_5269,N_5216);
nor U5442 (N_5442,N_5221,N_5293);
nand U5443 (N_5443,N_5225,N_5389);
nand U5444 (N_5444,N_5328,N_5384);
nor U5445 (N_5445,N_5239,N_5231);
and U5446 (N_5446,N_5393,N_5290);
xnor U5447 (N_5447,N_5316,N_5262);
nor U5448 (N_5448,N_5246,N_5396);
or U5449 (N_5449,N_5373,N_5266);
nand U5450 (N_5450,N_5324,N_5375);
nand U5451 (N_5451,N_5243,N_5342);
nand U5452 (N_5452,N_5202,N_5280);
or U5453 (N_5453,N_5315,N_5228);
nand U5454 (N_5454,N_5382,N_5283);
xnor U5455 (N_5455,N_5281,N_5305);
xor U5456 (N_5456,N_5267,N_5252);
or U5457 (N_5457,N_5330,N_5224);
xor U5458 (N_5458,N_5277,N_5378);
nand U5459 (N_5459,N_5388,N_5323);
nand U5460 (N_5460,N_5312,N_5353);
xnor U5461 (N_5461,N_5300,N_5304);
or U5462 (N_5462,N_5368,N_5279);
or U5463 (N_5463,N_5292,N_5210);
or U5464 (N_5464,N_5365,N_5370);
xor U5465 (N_5465,N_5348,N_5206);
nand U5466 (N_5466,N_5205,N_5310);
nor U5467 (N_5467,N_5306,N_5259);
nand U5468 (N_5468,N_5327,N_5299);
and U5469 (N_5469,N_5326,N_5351);
nand U5470 (N_5470,N_5392,N_5394);
nor U5471 (N_5471,N_5250,N_5237);
nor U5472 (N_5472,N_5363,N_5308);
or U5473 (N_5473,N_5338,N_5399);
or U5474 (N_5474,N_5358,N_5270);
xor U5475 (N_5475,N_5319,N_5317);
nand U5476 (N_5476,N_5203,N_5214);
xnor U5477 (N_5477,N_5255,N_5234);
and U5478 (N_5478,N_5372,N_5291);
nand U5479 (N_5479,N_5309,N_5362);
or U5480 (N_5480,N_5244,N_5223);
or U5481 (N_5481,N_5298,N_5337);
xnor U5482 (N_5482,N_5343,N_5349);
nor U5483 (N_5483,N_5230,N_5287);
or U5484 (N_5484,N_5296,N_5248);
and U5485 (N_5485,N_5381,N_5387);
nand U5486 (N_5486,N_5313,N_5268);
nor U5487 (N_5487,N_5222,N_5213);
and U5488 (N_5488,N_5236,N_5209);
or U5489 (N_5489,N_5320,N_5275);
or U5490 (N_5490,N_5212,N_5321);
nor U5491 (N_5491,N_5307,N_5294);
xnor U5492 (N_5492,N_5240,N_5334);
nand U5493 (N_5493,N_5220,N_5233);
and U5494 (N_5494,N_5251,N_5295);
or U5495 (N_5495,N_5200,N_5325);
nand U5496 (N_5496,N_5256,N_5344);
nand U5497 (N_5497,N_5379,N_5235);
xor U5498 (N_5498,N_5249,N_5284);
xnor U5499 (N_5499,N_5386,N_5289);
nor U5500 (N_5500,N_5359,N_5261);
or U5501 (N_5501,N_5215,N_5351);
nor U5502 (N_5502,N_5262,N_5257);
and U5503 (N_5503,N_5336,N_5278);
or U5504 (N_5504,N_5259,N_5277);
nand U5505 (N_5505,N_5225,N_5337);
nand U5506 (N_5506,N_5216,N_5306);
nor U5507 (N_5507,N_5397,N_5355);
or U5508 (N_5508,N_5277,N_5209);
and U5509 (N_5509,N_5277,N_5226);
nand U5510 (N_5510,N_5373,N_5370);
nand U5511 (N_5511,N_5363,N_5350);
nor U5512 (N_5512,N_5322,N_5275);
nand U5513 (N_5513,N_5332,N_5383);
nor U5514 (N_5514,N_5327,N_5301);
nand U5515 (N_5515,N_5240,N_5208);
and U5516 (N_5516,N_5352,N_5271);
or U5517 (N_5517,N_5308,N_5353);
nor U5518 (N_5518,N_5348,N_5350);
or U5519 (N_5519,N_5295,N_5260);
nor U5520 (N_5520,N_5236,N_5327);
or U5521 (N_5521,N_5297,N_5220);
nand U5522 (N_5522,N_5232,N_5377);
or U5523 (N_5523,N_5225,N_5280);
nand U5524 (N_5524,N_5278,N_5240);
and U5525 (N_5525,N_5342,N_5308);
nand U5526 (N_5526,N_5296,N_5313);
nor U5527 (N_5527,N_5354,N_5377);
nand U5528 (N_5528,N_5296,N_5226);
and U5529 (N_5529,N_5229,N_5223);
and U5530 (N_5530,N_5311,N_5359);
and U5531 (N_5531,N_5333,N_5205);
and U5532 (N_5532,N_5274,N_5256);
and U5533 (N_5533,N_5205,N_5227);
xnor U5534 (N_5534,N_5318,N_5254);
xor U5535 (N_5535,N_5382,N_5257);
or U5536 (N_5536,N_5219,N_5360);
or U5537 (N_5537,N_5399,N_5391);
nor U5538 (N_5538,N_5329,N_5338);
nor U5539 (N_5539,N_5240,N_5311);
and U5540 (N_5540,N_5374,N_5376);
xnor U5541 (N_5541,N_5314,N_5285);
and U5542 (N_5542,N_5220,N_5307);
nor U5543 (N_5543,N_5277,N_5266);
xor U5544 (N_5544,N_5261,N_5201);
or U5545 (N_5545,N_5269,N_5310);
xnor U5546 (N_5546,N_5304,N_5326);
nor U5547 (N_5547,N_5275,N_5295);
nor U5548 (N_5548,N_5386,N_5261);
nor U5549 (N_5549,N_5326,N_5208);
nand U5550 (N_5550,N_5320,N_5306);
or U5551 (N_5551,N_5223,N_5352);
xor U5552 (N_5552,N_5297,N_5325);
or U5553 (N_5553,N_5294,N_5368);
xor U5554 (N_5554,N_5365,N_5383);
nor U5555 (N_5555,N_5263,N_5306);
and U5556 (N_5556,N_5379,N_5319);
nand U5557 (N_5557,N_5393,N_5361);
nor U5558 (N_5558,N_5347,N_5373);
and U5559 (N_5559,N_5388,N_5226);
or U5560 (N_5560,N_5202,N_5326);
nor U5561 (N_5561,N_5265,N_5275);
or U5562 (N_5562,N_5297,N_5315);
xor U5563 (N_5563,N_5281,N_5399);
nor U5564 (N_5564,N_5383,N_5260);
nand U5565 (N_5565,N_5262,N_5226);
nor U5566 (N_5566,N_5259,N_5242);
and U5567 (N_5567,N_5351,N_5312);
xnor U5568 (N_5568,N_5365,N_5318);
or U5569 (N_5569,N_5354,N_5317);
or U5570 (N_5570,N_5383,N_5276);
nor U5571 (N_5571,N_5298,N_5280);
nand U5572 (N_5572,N_5273,N_5243);
and U5573 (N_5573,N_5231,N_5395);
xnor U5574 (N_5574,N_5234,N_5357);
xor U5575 (N_5575,N_5399,N_5245);
or U5576 (N_5576,N_5309,N_5327);
or U5577 (N_5577,N_5240,N_5261);
and U5578 (N_5578,N_5202,N_5367);
or U5579 (N_5579,N_5249,N_5379);
nand U5580 (N_5580,N_5328,N_5218);
and U5581 (N_5581,N_5288,N_5290);
nor U5582 (N_5582,N_5214,N_5337);
xnor U5583 (N_5583,N_5291,N_5315);
nand U5584 (N_5584,N_5327,N_5312);
nor U5585 (N_5585,N_5261,N_5362);
xor U5586 (N_5586,N_5395,N_5225);
nor U5587 (N_5587,N_5257,N_5267);
and U5588 (N_5588,N_5336,N_5388);
and U5589 (N_5589,N_5272,N_5240);
xnor U5590 (N_5590,N_5380,N_5219);
xor U5591 (N_5591,N_5203,N_5299);
nor U5592 (N_5592,N_5258,N_5356);
nor U5593 (N_5593,N_5353,N_5263);
nor U5594 (N_5594,N_5311,N_5318);
nor U5595 (N_5595,N_5354,N_5387);
and U5596 (N_5596,N_5213,N_5243);
or U5597 (N_5597,N_5285,N_5385);
xnor U5598 (N_5598,N_5242,N_5332);
xor U5599 (N_5599,N_5283,N_5259);
xor U5600 (N_5600,N_5416,N_5485);
nand U5601 (N_5601,N_5465,N_5582);
xor U5602 (N_5602,N_5529,N_5594);
nor U5603 (N_5603,N_5576,N_5404);
xnor U5604 (N_5604,N_5454,N_5461);
nand U5605 (N_5605,N_5561,N_5500);
nor U5606 (N_5606,N_5541,N_5460);
xor U5607 (N_5607,N_5532,N_5421);
nor U5608 (N_5608,N_5528,N_5525);
nor U5609 (N_5609,N_5572,N_5507);
nand U5610 (N_5610,N_5508,N_5456);
nand U5611 (N_5611,N_5530,N_5544);
nand U5612 (N_5612,N_5567,N_5433);
nor U5613 (N_5613,N_5554,N_5592);
or U5614 (N_5614,N_5584,N_5571);
and U5615 (N_5615,N_5440,N_5523);
and U5616 (N_5616,N_5546,N_5463);
xor U5617 (N_5617,N_5423,N_5549);
and U5618 (N_5618,N_5413,N_5574);
nor U5619 (N_5619,N_5451,N_5406);
nand U5620 (N_5620,N_5462,N_5402);
nand U5621 (N_5621,N_5470,N_5459);
xnor U5622 (N_5622,N_5597,N_5579);
nor U5623 (N_5623,N_5498,N_5448);
xnor U5624 (N_5624,N_5452,N_5563);
and U5625 (N_5625,N_5457,N_5506);
and U5626 (N_5626,N_5480,N_5518);
nor U5627 (N_5627,N_5581,N_5401);
nand U5628 (N_5628,N_5533,N_5495);
nand U5629 (N_5629,N_5468,N_5443);
or U5630 (N_5630,N_5512,N_5573);
or U5631 (N_5631,N_5475,N_5479);
xor U5632 (N_5632,N_5441,N_5472);
and U5633 (N_5633,N_5474,N_5410);
nor U5634 (N_5634,N_5545,N_5531);
nand U5635 (N_5635,N_5434,N_5471);
xnor U5636 (N_5636,N_5431,N_5504);
nand U5637 (N_5637,N_5478,N_5509);
or U5638 (N_5638,N_5464,N_5400);
or U5639 (N_5639,N_5537,N_5599);
and U5640 (N_5640,N_5578,N_5503);
or U5641 (N_5641,N_5477,N_5420);
and U5642 (N_5642,N_5505,N_5522);
nor U5643 (N_5643,N_5535,N_5487);
or U5644 (N_5644,N_5499,N_5435);
and U5645 (N_5645,N_5557,N_5534);
and U5646 (N_5646,N_5515,N_5419);
xor U5647 (N_5647,N_5483,N_5439);
or U5648 (N_5648,N_5412,N_5590);
nor U5649 (N_5649,N_5447,N_5488);
xnor U5650 (N_5650,N_5540,N_5445);
nor U5651 (N_5651,N_5565,N_5497);
and U5652 (N_5652,N_5559,N_5493);
nand U5653 (N_5653,N_5438,N_5444);
nor U5654 (N_5654,N_5494,N_5586);
and U5655 (N_5655,N_5539,N_5418);
or U5656 (N_5656,N_5442,N_5536);
nand U5657 (N_5657,N_5517,N_5467);
nor U5658 (N_5658,N_5486,N_5575);
xor U5659 (N_5659,N_5593,N_5427);
nor U5660 (N_5660,N_5405,N_5548);
and U5661 (N_5661,N_5436,N_5414);
nor U5662 (N_5662,N_5564,N_5473);
nand U5663 (N_5663,N_5511,N_5526);
xor U5664 (N_5664,N_5492,N_5422);
xor U5665 (N_5665,N_5569,N_5550);
or U5666 (N_5666,N_5596,N_5481);
nor U5667 (N_5667,N_5450,N_5484);
nor U5668 (N_5668,N_5408,N_5598);
xor U5669 (N_5669,N_5556,N_5424);
nor U5670 (N_5670,N_5551,N_5562);
xnor U5671 (N_5671,N_5458,N_5403);
and U5672 (N_5672,N_5510,N_5589);
or U5673 (N_5673,N_5437,N_5519);
nand U5674 (N_5674,N_5585,N_5583);
nand U5675 (N_5675,N_5560,N_5566);
nand U5676 (N_5676,N_5489,N_5580);
nor U5677 (N_5677,N_5568,N_5587);
nand U5678 (N_5678,N_5521,N_5516);
nand U5679 (N_5679,N_5552,N_5527);
nand U5680 (N_5680,N_5547,N_5491);
nor U5681 (N_5681,N_5417,N_5409);
nor U5682 (N_5682,N_5453,N_5558);
nand U5683 (N_5683,N_5425,N_5555);
or U5684 (N_5684,N_5501,N_5469);
nand U5685 (N_5685,N_5428,N_5430);
nand U5686 (N_5686,N_5407,N_5595);
nand U5687 (N_5687,N_5513,N_5588);
xor U5688 (N_5688,N_5446,N_5426);
nor U5689 (N_5689,N_5524,N_5591);
nor U5690 (N_5690,N_5429,N_5482);
xnor U5691 (N_5691,N_5496,N_5432);
and U5692 (N_5692,N_5455,N_5502);
xnor U5693 (N_5693,N_5476,N_5570);
nor U5694 (N_5694,N_5553,N_5415);
nand U5695 (N_5695,N_5542,N_5577);
and U5696 (N_5696,N_5538,N_5543);
xor U5697 (N_5697,N_5490,N_5411);
or U5698 (N_5698,N_5449,N_5466);
and U5699 (N_5699,N_5514,N_5520);
xor U5700 (N_5700,N_5518,N_5586);
nor U5701 (N_5701,N_5406,N_5570);
nand U5702 (N_5702,N_5532,N_5562);
nor U5703 (N_5703,N_5406,N_5441);
and U5704 (N_5704,N_5580,N_5544);
or U5705 (N_5705,N_5545,N_5550);
nor U5706 (N_5706,N_5573,N_5407);
nand U5707 (N_5707,N_5546,N_5572);
nor U5708 (N_5708,N_5564,N_5408);
nand U5709 (N_5709,N_5583,N_5420);
or U5710 (N_5710,N_5406,N_5517);
xor U5711 (N_5711,N_5510,N_5493);
nand U5712 (N_5712,N_5421,N_5585);
and U5713 (N_5713,N_5492,N_5521);
nor U5714 (N_5714,N_5416,N_5432);
or U5715 (N_5715,N_5432,N_5595);
nand U5716 (N_5716,N_5552,N_5568);
and U5717 (N_5717,N_5450,N_5447);
xor U5718 (N_5718,N_5480,N_5439);
nor U5719 (N_5719,N_5445,N_5509);
or U5720 (N_5720,N_5521,N_5559);
or U5721 (N_5721,N_5520,N_5404);
or U5722 (N_5722,N_5507,N_5425);
and U5723 (N_5723,N_5558,N_5414);
nor U5724 (N_5724,N_5534,N_5506);
nor U5725 (N_5725,N_5463,N_5507);
and U5726 (N_5726,N_5477,N_5505);
nor U5727 (N_5727,N_5526,N_5402);
or U5728 (N_5728,N_5532,N_5450);
nor U5729 (N_5729,N_5422,N_5586);
and U5730 (N_5730,N_5433,N_5416);
and U5731 (N_5731,N_5534,N_5575);
nor U5732 (N_5732,N_5413,N_5560);
and U5733 (N_5733,N_5497,N_5477);
or U5734 (N_5734,N_5400,N_5587);
xnor U5735 (N_5735,N_5419,N_5423);
xnor U5736 (N_5736,N_5487,N_5485);
xnor U5737 (N_5737,N_5504,N_5414);
nand U5738 (N_5738,N_5494,N_5598);
nor U5739 (N_5739,N_5484,N_5557);
nor U5740 (N_5740,N_5431,N_5548);
nor U5741 (N_5741,N_5461,N_5553);
nor U5742 (N_5742,N_5573,N_5422);
nor U5743 (N_5743,N_5577,N_5508);
xnor U5744 (N_5744,N_5530,N_5409);
or U5745 (N_5745,N_5532,N_5494);
and U5746 (N_5746,N_5579,N_5458);
and U5747 (N_5747,N_5434,N_5476);
or U5748 (N_5748,N_5587,N_5539);
and U5749 (N_5749,N_5421,N_5408);
or U5750 (N_5750,N_5483,N_5574);
xor U5751 (N_5751,N_5430,N_5429);
nor U5752 (N_5752,N_5510,N_5401);
and U5753 (N_5753,N_5422,N_5599);
and U5754 (N_5754,N_5550,N_5571);
nor U5755 (N_5755,N_5443,N_5519);
or U5756 (N_5756,N_5598,N_5458);
or U5757 (N_5757,N_5426,N_5511);
nor U5758 (N_5758,N_5562,N_5594);
nor U5759 (N_5759,N_5516,N_5405);
or U5760 (N_5760,N_5512,N_5412);
or U5761 (N_5761,N_5576,N_5442);
nand U5762 (N_5762,N_5588,N_5409);
nor U5763 (N_5763,N_5523,N_5501);
xnor U5764 (N_5764,N_5519,N_5550);
nor U5765 (N_5765,N_5535,N_5405);
xnor U5766 (N_5766,N_5497,N_5547);
and U5767 (N_5767,N_5570,N_5428);
xnor U5768 (N_5768,N_5445,N_5438);
nor U5769 (N_5769,N_5567,N_5589);
or U5770 (N_5770,N_5558,N_5507);
nor U5771 (N_5771,N_5497,N_5437);
xor U5772 (N_5772,N_5437,N_5439);
or U5773 (N_5773,N_5560,N_5537);
and U5774 (N_5774,N_5515,N_5441);
nand U5775 (N_5775,N_5528,N_5592);
nand U5776 (N_5776,N_5417,N_5477);
and U5777 (N_5777,N_5431,N_5463);
nand U5778 (N_5778,N_5592,N_5430);
nor U5779 (N_5779,N_5415,N_5411);
nor U5780 (N_5780,N_5566,N_5435);
xor U5781 (N_5781,N_5415,N_5426);
or U5782 (N_5782,N_5450,N_5513);
and U5783 (N_5783,N_5508,N_5454);
nor U5784 (N_5784,N_5403,N_5499);
xor U5785 (N_5785,N_5591,N_5531);
xnor U5786 (N_5786,N_5544,N_5570);
and U5787 (N_5787,N_5429,N_5599);
nand U5788 (N_5788,N_5566,N_5467);
xor U5789 (N_5789,N_5448,N_5577);
and U5790 (N_5790,N_5464,N_5569);
and U5791 (N_5791,N_5543,N_5442);
or U5792 (N_5792,N_5595,N_5456);
nand U5793 (N_5793,N_5535,N_5590);
nor U5794 (N_5794,N_5449,N_5426);
and U5795 (N_5795,N_5505,N_5443);
nand U5796 (N_5796,N_5523,N_5571);
and U5797 (N_5797,N_5560,N_5586);
xnor U5798 (N_5798,N_5478,N_5465);
nand U5799 (N_5799,N_5581,N_5516);
or U5800 (N_5800,N_5619,N_5614);
nor U5801 (N_5801,N_5749,N_5687);
and U5802 (N_5802,N_5617,N_5618);
nand U5803 (N_5803,N_5611,N_5643);
nand U5804 (N_5804,N_5650,N_5606);
or U5805 (N_5805,N_5775,N_5753);
nor U5806 (N_5806,N_5750,N_5710);
nand U5807 (N_5807,N_5686,N_5625);
and U5808 (N_5808,N_5731,N_5740);
xor U5809 (N_5809,N_5665,N_5676);
nand U5810 (N_5810,N_5719,N_5738);
nor U5811 (N_5811,N_5766,N_5636);
xnor U5812 (N_5812,N_5799,N_5670);
nand U5813 (N_5813,N_5605,N_5760);
and U5814 (N_5814,N_5716,N_5737);
and U5815 (N_5815,N_5717,N_5616);
xnor U5816 (N_5816,N_5721,N_5627);
nor U5817 (N_5817,N_5767,N_5600);
or U5818 (N_5818,N_5725,N_5756);
and U5819 (N_5819,N_5777,N_5692);
nand U5820 (N_5820,N_5714,N_5680);
nor U5821 (N_5821,N_5651,N_5628);
nor U5822 (N_5822,N_5615,N_5701);
nand U5823 (N_5823,N_5654,N_5792);
nor U5824 (N_5824,N_5757,N_5720);
xnor U5825 (N_5825,N_5679,N_5640);
or U5826 (N_5826,N_5659,N_5764);
and U5827 (N_5827,N_5695,N_5662);
xor U5828 (N_5828,N_5786,N_5704);
nor U5829 (N_5829,N_5774,N_5706);
xnor U5830 (N_5830,N_5747,N_5648);
nand U5831 (N_5831,N_5794,N_5655);
nand U5832 (N_5832,N_5769,N_5700);
nor U5833 (N_5833,N_5796,N_5736);
nor U5834 (N_5834,N_5663,N_5660);
nor U5835 (N_5835,N_5694,N_5730);
xnor U5836 (N_5836,N_5782,N_5669);
xor U5837 (N_5837,N_5772,N_5728);
and U5838 (N_5838,N_5644,N_5798);
xnor U5839 (N_5839,N_5675,N_5791);
xnor U5840 (N_5840,N_5751,N_5672);
nor U5841 (N_5841,N_5607,N_5733);
xnor U5842 (N_5842,N_5682,N_5781);
nand U5843 (N_5843,N_5661,N_5678);
nand U5844 (N_5844,N_5604,N_5688);
and U5845 (N_5845,N_5624,N_5601);
or U5846 (N_5846,N_5784,N_5696);
and U5847 (N_5847,N_5797,N_5629);
xor U5848 (N_5848,N_5621,N_5674);
and U5849 (N_5849,N_5633,N_5709);
or U5850 (N_5850,N_5787,N_5745);
nor U5851 (N_5851,N_5683,N_5761);
nand U5852 (N_5852,N_5759,N_5609);
xnor U5853 (N_5853,N_5681,N_5713);
and U5854 (N_5854,N_5754,N_5622);
or U5855 (N_5855,N_5705,N_5723);
or U5856 (N_5856,N_5652,N_5697);
or U5857 (N_5857,N_5726,N_5645);
nand U5858 (N_5858,N_5620,N_5789);
or U5859 (N_5859,N_5765,N_5715);
and U5860 (N_5860,N_5758,N_5780);
xor U5861 (N_5861,N_5752,N_5613);
or U5862 (N_5862,N_5763,N_5668);
xnor U5863 (N_5863,N_5666,N_5641);
and U5864 (N_5864,N_5691,N_5690);
nand U5865 (N_5865,N_5795,N_5707);
xnor U5866 (N_5866,N_5649,N_5646);
xnor U5867 (N_5867,N_5739,N_5667);
and U5868 (N_5868,N_5742,N_5639);
xnor U5869 (N_5869,N_5638,N_5664);
nor U5870 (N_5870,N_5727,N_5693);
and U5871 (N_5871,N_5722,N_5741);
nor U5872 (N_5872,N_5642,N_5702);
and U5873 (N_5873,N_5788,N_5608);
or U5874 (N_5874,N_5623,N_5703);
and U5875 (N_5875,N_5743,N_5724);
or U5876 (N_5876,N_5712,N_5783);
nor U5877 (N_5877,N_5612,N_5734);
nand U5878 (N_5878,N_5793,N_5632);
and U5879 (N_5879,N_5647,N_5729);
and U5880 (N_5880,N_5778,N_5785);
and U5881 (N_5881,N_5653,N_5762);
and U5882 (N_5882,N_5657,N_5626);
nor U5883 (N_5883,N_5698,N_5602);
or U5884 (N_5884,N_5779,N_5630);
nor U5885 (N_5885,N_5634,N_5673);
nor U5886 (N_5886,N_5755,N_5658);
and U5887 (N_5887,N_5637,N_5631);
nor U5888 (N_5888,N_5603,N_5771);
and U5889 (N_5889,N_5684,N_5744);
xor U5890 (N_5890,N_5770,N_5732);
xnor U5891 (N_5891,N_5610,N_5708);
and U5892 (N_5892,N_5735,N_5656);
xnor U5893 (N_5893,N_5748,N_5746);
nand U5894 (N_5894,N_5635,N_5711);
or U5895 (N_5895,N_5768,N_5677);
nor U5896 (N_5896,N_5790,N_5671);
nor U5897 (N_5897,N_5773,N_5699);
nor U5898 (N_5898,N_5776,N_5685);
or U5899 (N_5899,N_5718,N_5689);
nand U5900 (N_5900,N_5670,N_5711);
and U5901 (N_5901,N_5651,N_5700);
and U5902 (N_5902,N_5717,N_5697);
nor U5903 (N_5903,N_5711,N_5634);
xnor U5904 (N_5904,N_5623,N_5790);
xnor U5905 (N_5905,N_5724,N_5680);
nand U5906 (N_5906,N_5752,N_5631);
nand U5907 (N_5907,N_5753,N_5740);
and U5908 (N_5908,N_5614,N_5644);
xnor U5909 (N_5909,N_5769,N_5753);
nand U5910 (N_5910,N_5758,N_5643);
xor U5911 (N_5911,N_5675,N_5634);
nor U5912 (N_5912,N_5658,N_5770);
or U5913 (N_5913,N_5651,N_5600);
xnor U5914 (N_5914,N_5684,N_5604);
nor U5915 (N_5915,N_5727,N_5707);
and U5916 (N_5916,N_5748,N_5740);
and U5917 (N_5917,N_5779,N_5744);
xor U5918 (N_5918,N_5719,N_5604);
xnor U5919 (N_5919,N_5778,N_5733);
nand U5920 (N_5920,N_5632,N_5648);
and U5921 (N_5921,N_5793,N_5630);
nand U5922 (N_5922,N_5690,N_5622);
nor U5923 (N_5923,N_5677,N_5682);
nand U5924 (N_5924,N_5716,N_5637);
nand U5925 (N_5925,N_5714,N_5760);
and U5926 (N_5926,N_5788,N_5724);
and U5927 (N_5927,N_5610,N_5601);
or U5928 (N_5928,N_5626,N_5764);
nor U5929 (N_5929,N_5624,N_5713);
xor U5930 (N_5930,N_5719,N_5725);
nor U5931 (N_5931,N_5667,N_5724);
and U5932 (N_5932,N_5610,N_5750);
nand U5933 (N_5933,N_5652,N_5605);
nand U5934 (N_5934,N_5715,N_5759);
nor U5935 (N_5935,N_5730,N_5791);
nor U5936 (N_5936,N_5678,N_5700);
xnor U5937 (N_5937,N_5669,N_5616);
xor U5938 (N_5938,N_5650,N_5697);
nand U5939 (N_5939,N_5682,N_5752);
and U5940 (N_5940,N_5692,N_5763);
nand U5941 (N_5941,N_5768,N_5625);
nor U5942 (N_5942,N_5600,N_5670);
nor U5943 (N_5943,N_5718,N_5642);
nor U5944 (N_5944,N_5628,N_5754);
nor U5945 (N_5945,N_5774,N_5641);
xor U5946 (N_5946,N_5682,N_5687);
nor U5947 (N_5947,N_5710,N_5720);
nand U5948 (N_5948,N_5739,N_5631);
xnor U5949 (N_5949,N_5769,N_5793);
and U5950 (N_5950,N_5698,N_5656);
and U5951 (N_5951,N_5653,N_5655);
xnor U5952 (N_5952,N_5610,N_5628);
nor U5953 (N_5953,N_5735,N_5799);
nand U5954 (N_5954,N_5766,N_5784);
nor U5955 (N_5955,N_5751,N_5733);
and U5956 (N_5956,N_5706,N_5628);
or U5957 (N_5957,N_5773,N_5650);
or U5958 (N_5958,N_5691,N_5617);
nand U5959 (N_5959,N_5625,N_5687);
xor U5960 (N_5960,N_5721,N_5795);
nand U5961 (N_5961,N_5624,N_5761);
and U5962 (N_5962,N_5750,N_5735);
nor U5963 (N_5963,N_5783,N_5700);
nand U5964 (N_5964,N_5644,N_5725);
and U5965 (N_5965,N_5771,N_5701);
nor U5966 (N_5966,N_5691,N_5692);
or U5967 (N_5967,N_5774,N_5744);
nand U5968 (N_5968,N_5675,N_5692);
and U5969 (N_5969,N_5743,N_5635);
or U5970 (N_5970,N_5680,N_5659);
or U5971 (N_5971,N_5769,N_5738);
xnor U5972 (N_5972,N_5764,N_5635);
xor U5973 (N_5973,N_5604,N_5747);
xnor U5974 (N_5974,N_5675,N_5773);
nor U5975 (N_5975,N_5636,N_5798);
nor U5976 (N_5976,N_5702,N_5608);
or U5977 (N_5977,N_5779,N_5702);
and U5978 (N_5978,N_5605,N_5700);
and U5979 (N_5979,N_5796,N_5620);
xor U5980 (N_5980,N_5623,N_5675);
nor U5981 (N_5981,N_5621,N_5660);
nand U5982 (N_5982,N_5660,N_5798);
xnor U5983 (N_5983,N_5701,N_5694);
nor U5984 (N_5984,N_5772,N_5734);
or U5985 (N_5985,N_5769,N_5748);
nor U5986 (N_5986,N_5713,N_5771);
xor U5987 (N_5987,N_5754,N_5652);
nand U5988 (N_5988,N_5664,N_5778);
xnor U5989 (N_5989,N_5610,N_5797);
nor U5990 (N_5990,N_5767,N_5601);
and U5991 (N_5991,N_5631,N_5618);
nand U5992 (N_5992,N_5638,N_5704);
or U5993 (N_5993,N_5649,N_5757);
nand U5994 (N_5994,N_5776,N_5617);
nor U5995 (N_5995,N_5663,N_5643);
nand U5996 (N_5996,N_5668,N_5736);
nor U5997 (N_5997,N_5680,N_5725);
xnor U5998 (N_5998,N_5651,N_5781);
or U5999 (N_5999,N_5721,N_5646);
or U6000 (N_6000,N_5840,N_5892);
nand U6001 (N_6001,N_5990,N_5866);
nand U6002 (N_6002,N_5880,N_5810);
and U6003 (N_6003,N_5912,N_5996);
nand U6004 (N_6004,N_5975,N_5909);
nor U6005 (N_6005,N_5964,N_5906);
or U6006 (N_6006,N_5986,N_5901);
nand U6007 (N_6007,N_5828,N_5848);
or U6008 (N_6008,N_5876,N_5968);
or U6009 (N_6009,N_5830,N_5920);
xor U6010 (N_6010,N_5800,N_5854);
or U6011 (N_6011,N_5963,N_5823);
nand U6012 (N_6012,N_5818,N_5918);
xnor U6013 (N_6013,N_5845,N_5937);
or U6014 (N_6014,N_5944,N_5821);
nor U6015 (N_6015,N_5811,N_5939);
nor U6016 (N_6016,N_5951,N_5860);
or U6017 (N_6017,N_5988,N_5857);
nand U6018 (N_6018,N_5908,N_5980);
nor U6019 (N_6019,N_5837,N_5997);
xnor U6020 (N_6020,N_5977,N_5868);
nor U6021 (N_6021,N_5842,N_5970);
or U6022 (N_6022,N_5923,N_5894);
nand U6023 (N_6023,N_5819,N_5808);
or U6024 (N_6024,N_5905,N_5884);
xnor U6025 (N_6025,N_5881,N_5993);
nor U6026 (N_6026,N_5816,N_5917);
nor U6027 (N_6027,N_5915,N_5979);
and U6028 (N_6028,N_5889,N_5853);
nor U6029 (N_6029,N_5947,N_5803);
or U6030 (N_6030,N_5882,N_5812);
xor U6031 (N_6031,N_5833,N_5844);
xnor U6032 (N_6032,N_5954,N_5832);
nor U6033 (N_6033,N_5888,N_5934);
nor U6034 (N_6034,N_5813,N_5836);
nor U6035 (N_6035,N_5814,N_5924);
xnor U6036 (N_6036,N_5862,N_5942);
nor U6037 (N_6037,N_5815,N_5929);
xor U6038 (N_6038,N_5843,N_5855);
nand U6039 (N_6039,N_5981,N_5935);
xnor U6040 (N_6040,N_5956,N_5941);
or U6041 (N_6041,N_5802,N_5886);
nand U6042 (N_6042,N_5958,N_5846);
and U6043 (N_6043,N_5926,N_5829);
nand U6044 (N_6044,N_5932,N_5982);
xnor U6045 (N_6045,N_5839,N_5870);
xnor U6046 (N_6046,N_5893,N_5885);
and U6047 (N_6047,N_5946,N_5807);
xnor U6048 (N_6048,N_5835,N_5873);
or U6049 (N_6049,N_5838,N_5994);
nor U6050 (N_6050,N_5971,N_5927);
nor U6051 (N_6051,N_5867,N_5989);
or U6052 (N_6052,N_5865,N_5938);
or U6053 (N_6053,N_5902,N_5953);
nand U6054 (N_6054,N_5972,N_5921);
nand U6055 (N_6055,N_5841,N_5897);
and U6056 (N_6056,N_5883,N_5851);
or U6057 (N_6057,N_5900,N_5962);
or U6058 (N_6058,N_5861,N_5945);
and U6059 (N_6059,N_5991,N_5878);
nand U6060 (N_6060,N_5933,N_5890);
or U6061 (N_6061,N_5976,N_5858);
or U6062 (N_6062,N_5913,N_5859);
nor U6063 (N_6063,N_5914,N_5872);
nand U6064 (N_6064,N_5899,N_5974);
xor U6065 (N_6065,N_5864,N_5983);
or U6066 (N_6066,N_5925,N_5804);
and U6067 (N_6067,N_5978,N_5984);
and U6068 (N_6068,N_5961,N_5992);
or U6069 (N_6069,N_5831,N_5911);
and U6070 (N_6070,N_5949,N_5966);
nand U6071 (N_6071,N_5904,N_5849);
xnor U6072 (N_6072,N_5903,N_5957);
or U6073 (N_6073,N_5936,N_5931);
and U6074 (N_6074,N_5801,N_5995);
or U6075 (N_6075,N_5959,N_5910);
and U6076 (N_6076,N_5948,N_5874);
and U6077 (N_6077,N_5998,N_5869);
or U6078 (N_6078,N_5826,N_5930);
nor U6079 (N_6079,N_5825,N_5852);
or U6080 (N_6080,N_5875,N_5820);
or U6081 (N_6081,N_5887,N_5907);
or U6082 (N_6082,N_5898,N_5965);
and U6083 (N_6083,N_5856,N_5916);
nor U6084 (N_6084,N_5834,N_5863);
xor U6085 (N_6085,N_5827,N_5806);
nand U6086 (N_6086,N_5805,N_5969);
nor U6087 (N_6087,N_5943,N_5952);
nor U6088 (N_6088,N_5822,N_5879);
nor U6089 (N_6089,N_5891,N_5960);
or U6090 (N_6090,N_5985,N_5955);
and U6091 (N_6091,N_5973,N_5847);
nand U6092 (N_6092,N_5950,N_5850);
and U6093 (N_6093,N_5877,N_5817);
nor U6094 (N_6094,N_5895,N_5871);
and U6095 (N_6095,N_5928,N_5824);
and U6096 (N_6096,N_5919,N_5940);
nor U6097 (N_6097,N_5999,N_5967);
or U6098 (N_6098,N_5922,N_5809);
xor U6099 (N_6099,N_5896,N_5987);
nand U6100 (N_6100,N_5818,N_5914);
nand U6101 (N_6101,N_5906,N_5970);
nand U6102 (N_6102,N_5878,N_5801);
and U6103 (N_6103,N_5835,N_5807);
nor U6104 (N_6104,N_5826,N_5918);
nor U6105 (N_6105,N_5989,N_5956);
nor U6106 (N_6106,N_5815,N_5936);
or U6107 (N_6107,N_5973,N_5807);
xor U6108 (N_6108,N_5890,N_5985);
nor U6109 (N_6109,N_5891,N_5975);
nand U6110 (N_6110,N_5807,N_5849);
nand U6111 (N_6111,N_5972,N_5849);
nand U6112 (N_6112,N_5949,N_5807);
xnor U6113 (N_6113,N_5818,N_5876);
nor U6114 (N_6114,N_5991,N_5967);
and U6115 (N_6115,N_5865,N_5819);
nand U6116 (N_6116,N_5902,N_5883);
nand U6117 (N_6117,N_5888,N_5906);
or U6118 (N_6118,N_5837,N_5985);
xor U6119 (N_6119,N_5948,N_5888);
and U6120 (N_6120,N_5837,N_5876);
nor U6121 (N_6121,N_5811,N_5917);
nand U6122 (N_6122,N_5942,N_5988);
nor U6123 (N_6123,N_5825,N_5921);
xor U6124 (N_6124,N_5937,N_5992);
xor U6125 (N_6125,N_5943,N_5962);
and U6126 (N_6126,N_5995,N_5975);
nor U6127 (N_6127,N_5803,N_5887);
or U6128 (N_6128,N_5959,N_5919);
or U6129 (N_6129,N_5813,N_5932);
or U6130 (N_6130,N_5984,N_5890);
xnor U6131 (N_6131,N_5898,N_5836);
xor U6132 (N_6132,N_5949,N_5997);
and U6133 (N_6133,N_5973,N_5828);
or U6134 (N_6134,N_5968,N_5928);
xnor U6135 (N_6135,N_5930,N_5897);
xnor U6136 (N_6136,N_5980,N_5910);
and U6137 (N_6137,N_5843,N_5842);
xnor U6138 (N_6138,N_5817,N_5864);
nand U6139 (N_6139,N_5995,N_5878);
and U6140 (N_6140,N_5946,N_5928);
or U6141 (N_6141,N_5801,N_5888);
or U6142 (N_6142,N_5862,N_5803);
xor U6143 (N_6143,N_5958,N_5941);
nand U6144 (N_6144,N_5956,N_5948);
nand U6145 (N_6145,N_5817,N_5838);
and U6146 (N_6146,N_5875,N_5923);
or U6147 (N_6147,N_5845,N_5901);
xor U6148 (N_6148,N_5904,N_5826);
nand U6149 (N_6149,N_5828,N_5903);
nor U6150 (N_6150,N_5842,N_5915);
or U6151 (N_6151,N_5949,N_5935);
and U6152 (N_6152,N_5868,N_5952);
and U6153 (N_6153,N_5901,N_5991);
nand U6154 (N_6154,N_5943,N_5826);
xor U6155 (N_6155,N_5922,N_5977);
or U6156 (N_6156,N_5990,N_5892);
or U6157 (N_6157,N_5962,N_5985);
and U6158 (N_6158,N_5864,N_5919);
nand U6159 (N_6159,N_5835,N_5859);
and U6160 (N_6160,N_5901,N_5926);
or U6161 (N_6161,N_5907,N_5807);
xnor U6162 (N_6162,N_5879,N_5980);
and U6163 (N_6163,N_5858,N_5925);
nand U6164 (N_6164,N_5833,N_5829);
or U6165 (N_6165,N_5985,N_5913);
or U6166 (N_6166,N_5942,N_5911);
nand U6167 (N_6167,N_5895,N_5959);
xnor U6168 (N_6168,N_5989,N_5947);
and U6169 (N_6169,N_5824,N_5894);
nor U6170 (N_6170,N_5864,N_5972);
nor U6171 (N_6171,N_5885,N_5806);
nor U6172 (N_6172,N_5843,N_5924);
or U6173 (N_6173,N_5909,N_5833);
xnor U6174 (N_6174,N_5863,N_5889);
nor U6175 (N_6175,N_5913,N_5956);
nor U6176 (N_6176,N_5951,N_5884);
xnor U6177 (N_6177,N_5988,N_5811);
and U6178 (N_6178,N_5885,N_5997);
or U6179 (N_6179,N_5800,N_5830);
xor U6180 (N_6180,N_5866,N_5965);
and U6181 (N_6181,N_5841,N_5955);
xor U6182 (N_6182,N_5819,N_5942);
or U6183 (N_6183,N_5883,N_5880);
and U6184 (N_6184,N_5917,N_5868);
nor U6185 (N_6185,N_5890,N_5877);
xor U6186 (N_6186,N_5857,N_5894);
nand U6187 (N_6187,N_5874,N_5982);
nor U6188 (N_6188,N_5962,N_5850);
xor U6189 (N_6189,N_5904,N_5888);
and U6190 (N_6190,N_5924,N_5972);
xor U6191 (N_6191,N_5852,N_5863);
nor U6192 (N_6192,N_5965,N_5873);
nand U6193 (N_6193,N_5834,N_5822);
nand U6194 (N_6194,N_5898,N_5806);
nor U6195 (N_6195,N_5988,N_5915);
nor U6196 (N_6196,N_5845,N_5967);
nand U6197 (N_6197,N_5844,N_5933);
and U6198 (N_6198,N_5855,N_5879);
nor U6199 (N_6199,N_5972,N_5949);
nand U6200 (N_6200,N_6072,N_6098);
nor U6201 (N_6201,N_6000,N_6183);
nor U6202 (N_6202,N_6125,N_6101);
xnor U6203 (N_6203,N_6026,N_6134);
and U6204 (N_6204,N_6150,N_6010);
or U6205 (N_6205,N_6067,N_6196);
or U6206 (N_6206,N_6038,N_6024);
nand U6207 (N_6207,N_6062,N_6083);
nand U6208 (N_6208,N_6020,N_6016);
and U6209 (N_6209,N_6191,N_6061);
nor U6210 (N_6210,N_6058,N_6055);
or U6211 (N_6211,N_6066,N_6109);
xor U6212 (N_6212,N_6132,N_6019);
nand U6213 (N_6213,N_6043,N_6131);
nand U6214 (N_6214,N_6141,N_6140);
or U6215 (N_6215,N_6057,N_6156);
or U6216 (N_6216,N_6040,N_6165);
nand U6217 (N_6217,N_6113,N_6112);
nor U6218 (N_6218,N_6130,N_6099);
nand U6219 (N_6219,N_6079,N_6135);
xnor U6220 (N_6220,N_6158,N_6092);
nand U6221 (N_6221,N_6153,N_6009);
and U6222 (N_6222,N_6106,N_6031);
nand U6223 (N_6223,N_6159,N_6189);
and U6224 (N_6224,N_6033,N_6044);
nand U6225 (N_6225,N_6021,N_6186);
xor U6226 (N_6226,N_6170,N_6075);
and U6227 (N_6227,N_6136,N_6126);
or U6228 (N_6228,N_6195,N_6184);
and U6229 (N_6229,N_6078,N_6198);
or U6230 (N_6230,N_6074,N_6197);
xor U6231 (N_6231,N_6137,N_6168);
xnor U6232 (N_6232,N_6121,N_6048);
nand U6233 (N_6233,N_6084,N_6080);
nor U6234 (N_6234,N_6146,N_6111);
nand U6235 (N_6235,N_6169,N_6088);
nand U6236 (N_6236,N_6172,N_6097);
nor U6237 (N_6237,N_6108,N_6178);
nor U6238 (N_6238,N_6037,N_6171);
or U6239 (N_6239,N_6003,N_6138);
nand U6240 (N_6240,N_6185,N_6139);
nand U6241 (N_6241,N_6029,N_6103);
nand U6242 (N_6242,N_6179,N_6176);
nor U6243 (N_6243,N_6081,N_6152);
nor U6244 (N_6244,N_6091,N_6071);
and U6245 (N_6245,N_6046,N_6012);
and U6246 (N_6246,N_6180,N_6114);
xor U6247 (N_6247,N_6073,N_6022);
nand U6248 (N_6248,N_6151,N_6070);
or U6249 (N_6249,N_6090,N_6059);
nand U6250 (N_6250,N_6045,N_6086);
nand U6251 (N_6251,N_6007,N_6036);
nand U6252 (N_6252,N_6120,N_6032);
nor U6253 (N_6253,N_6157,N_6006);
nand U6254 (N_6254,N_6077,N_6105);
and U6255 (N_6255,N_6142,N_6117);
and U6256 (N_6256,N_6161,N_6123);
nand U6257 (N_6257,N_6051,N_6085);
xnor U6258 (N_6258,N_6160,N_6144);
nand U6259 (N_6259,N_6047,N_6014);
and U6260 (N_6260,N_6148,N_6050);
nand U6261 (N_6261,N_6049,N_6052);
xor U6262 (N_6262,N_6053,N_6005);
nor U6263 (N_6263,N_6069,N_6166);
xor U6264 (N_6264,N_6192,N_6008);
xor U6265 (N_6265,N_6025,N_6182);
and U6266 (N_6266,N_6063,N_6174);
nand U6267 (N_6267,N_6133,N_6181);
nand U6268 (N_6268,N_6149,N_6102);
or U6269 (N_6269,N_6199,N_6147);
and U6270 (N_6270,N_6023,N_6128);
or U6271 (N_6271,N_6193,N_6145);
or U6272 (N_6272,N_6096,N_6162);
xnor U6273 (N_6273,N_6035,N_6030);
or U6274 (N_6274,N_6175,N_6104);
xor U6275 (N_6275,N_6002,N_6177);
nor U6276 (N_6276,N_6013,N_6187);
xnor U6277 (N_6277,N_6095,N_6100);
and U6278 (N_6278,N_6076,N_6018);
nand U6279 (N_6279,N_6118,N_6064);
and U6280 (N_6280,N_6154,N_6094);
or U6281 (N_6281,N_6119,N_6163);
and U6282 (N_6282,N_6034,N_6039);
or U6283 (N_6283,N_6011,N_6190);
and U6284 (N_6284,N_6087,N_6082);
xor U6285 (N_6285,N_6127,N_6041);
and U6286 (N_6286,N_6188,N_6089);
nand U6287 (N_6287,N_6068,N_6056);
nand U6288 (N_6288,N_6004,N_6042);
nor U6289 (N_6289,N_6107,N_6060);
nor U6290 (N_6290,N_6054,N_6093);
or U6291 (N_6291,N_6167,N_6001);
nand U6292 (N_6292,N_6017,N_6015);
and U6293 (N_6293,N_6028,N_6115);
xor U6294 (N_6294,N_6027,N_6194);
and U6295 (N_6295,N_6122,N_6116);
nor U6296 (N_6296,N_6129,N_6124);
nand U6297 (N_6297,N_6065,N_6143);
nand U6298 (N_6298,N_6164,N_6173);
and U6299 (N_6299,N_6110,N_6155);
or U6300 (N_6300,N_6186,N_6190);
or U6301 (N_6301,N_6063,N_6108);
xor U6302 (N_6302,N_6084,N_6180);
nand U6303 (N_6303,N_6135,N_6085);
nand U6304 (N_6304,N_6168,N_6148);
nor U6305 (N_6305,N_6032,N_6164);
nand U6306 (N_6306,N_6169,N_6147);
xor U6307 (N_6307,N_6062,N_6031);
nor U6308 (N_6308,N_6162,N_6134);
xor U6309 (N_6309,N_6092,N_6164);
and U6310 (N_6310,N_6159,N_6062);
nand U6311 (N_6311,N_6132,N_6101);
nand U6312 (N_6312,N_6195,N_6140);
and U6313 (N_6313,N_6172,N_6122);
nand U6314 (N_6314,N_6035,N_6192);
and U6315 (N_6315,N_6108,N_6175);
and U6316 (N_6316,N_6059,N_6148);
nor U6317 (N_6317,N_6195,N_6120);
and U6318 (N_6318,N_6063,N_6079);
nand U6319 (N_6319,N_6098,N_6033);
nor U6320 (N_6320,N_6145,N_6137);
nand U6321 (N_6321,N_6198,N_6172);
or U6322 (N_6322,N_6144,N_6151);
xnor U6323 (N_6323,N_6042,N_6112);
or U6324 (N_6324,N_6002,N_6173);
nand U6325 (N_6325,N_6046,N_6175);
xnor U6326 (N_6326,N_6132,N_6068);
nand U6327 (N_6327,N_6020,N_6010);
nor U6328 (N_6328,N_6039,N_6004);
xor U6329 (N_6329,N_6007,N_6098);
or U6330 (N_6330,N_6180,N_6063);
or U6331 (N_6331,N_6037,N_6194);
and U6332 (N_6332,N_6071,N_6012);
nor U6333 (N_6333,N_6107,N_6156);
xnor U6334 (N_6334,N_6186,N_6001);
or U6335 (N_6335,N_6087,N_6189);
xnor U6336 (N_6336,N_6064,N_6171);
and U6337 (N_6337,N_6001,N_6047);
nor U6338 (N_6338,N_6065,N_6030);
or U6339 (N_6339,N_6041,N_6182);
or U6340 (N_6340,N_6118,N_6177);
nand U6341 (N_6341,N_6148,N_6014);
nor U6342 (N_6342,N_6132,N_6141);
or U6343 (N_6343,N_6152,N_6042);
nor U6344 (N_6344,N_6129,N_6087);
xor U6345 (N_6345,N_6056,N_6148);
and U6346 (N_6346,N_6109,N_6191);
and U6347 (N_6347,N_6010,N_6144);
xor U6348 (N_6348,N_6174,N_6027);
nand U6349 (N_6349,N_6158,N_6140);
nor U6350 (N_6350,N_6084,N_6024);
and U6351 (N_6351,N_6192,N_6037);
xor U6352 (N_6352,N_6025,N_6067);
nor U6353 (N_6353,N_6048,N_6174);
xor U6354 (N_6354,N_6028,N_6076);
xor U6355 (N_6355,N_6090,N_6055);
nand U6356 (N_6356,N_6192,N_6069);
nor U6357 (N_6357,N_6012,N_6061);
nand U6358 (N_6358,N_6110,N_6184);
nor U6359 (N_6359,N_6077,N_6012);
nor U6360 (N_6360,N_6146,N_6135);
or U6361 (N_6361,N_6197,N_6064);
or U6362 (N_6362,N_6153,N_6152);
nor U6363 (N_6363,N_6075,N_6099);
nand U6364 (N_6364,N_6142,N_6156);
or U6365 (N_6365,N_6105,N_6154);
and U6366 (N_6366,N_6068,N_6004);
or U6367 (N_6367,N_6049,N_6082);
nand U6368 (N_6368,N_6069,N_6093);
nor U6369 (N_6369,N_6118,N_6055);
nand U6370 (N_6370,N_6100,N_6004);
xnor U6371 (N_6371,N_6081,N_6004);
or U6372 (N_6372,N_6009,N_6102);
or U6373 (N_6373,N_6174,N_6178);
nor U6374 (N_6374,N_6021,N_6081);
nand U6375 (N_6375,N_6057,N_6000);
and U6376 (N_6376,N_6120,N_6188);
or U6377 (N_6377,N_6186,N_6139);
nor U6378 (N_6378,N_6147,N_6135);
nor U6379 (N_6379,N_6087,N_6118);
and U6380 (N_6380,N_6106,N_6118);
and U6381 (N_6381,N_6030,N_6098);
nand U6382 (N_6382,N_6133,N_6191);
nor U6383 (N_6383,N_6169,N_6036);
or U6384 (N_6384,N_6137,N_6117);
or U6385 (N_6385,N_6088,N_6187);
nor U6386 (N_6386,N_6101,N_6109);
or U6387 (N_6387,N_6119,N_6103);
xnor U6388 (N_6388,N_6091,N_6129);
nor U6389 (N_6389,N_6184,N_6040);
nand U6390 (N_6390,N_6181,N_6051);
and U6391 (N_6391,N_6121,N_6041);
or U6392 (N_6392,N_6032,N_6178);
and U6393 (N_6393,N_6185,N_6129);
nand U6394 (N_6394,N_6054,N_6191);
and U6395 (N_6395,N_6015,N_6186);
xnor U6396 (N_6396,N_6053,N_6036);
nor U6397 (N_6397,N_6143,N_6163);
and U6398 (N_6398,N_6112,N_6055);
nor U6399 (N_6399,N_6043,N_6084);
nand U6400 (N_6400,N_6261,N_6301);
nand U6401 (N_6401,N_6264,N_6255);
nand U6402 (N_6402,N_6394,N_6342);
and U6403 (N_6403,N_6215,N_6380);
or U6404 (N_6404,N_6220,N_6396);
and U6405 (N_6405,N_6209,N_6218);
and U6406 (N_6406,N_6293,N_6249);
nor U6407 (N_6407,N_6327,N_6307);
and U6408 (N_6408,N_6360,N_6270);
nor U6409 (N_6409,N_6251,N_6388);
xnor U6410 (N_6410,N_6253,N_6393);
and U6411 (N_6411,N_6282,N_6354);
nand U6412 (N_6412,N_6239,N_6226);
nor U6413 (N_6413,N_6359,N_6305);
xor U6414 (N_6414,N_6240,N_6335);
or U6415 (N_6415,N_6281,N_6244);
nor U6416 (N_6416,N_6292,N_6367);
xor U6417 (N_6417,N_6263,N_6374);
xor U6418 (N_6418,N_6241,N_6274);
or U6419 (N_6419,N_6280,N_6213);
nand U6420 (N_6420,N_6375,N_6217);
or U6421 (N_6421,N_6331,N_6325);
or U6422 (N_6422,N_6236,N_6296);
or U6423 (N_6423,N_6302,N_6347);
and U6424 (N_6424,N_6372,N_6324);
nand U6425 (N_6425,N_6210,N_6288);
nand U6426 (N_6426,N_6246,N_6295);
and U6427 (N_6427,N_6221,N_6228);
nor U6428 (N_6428,N_6219,N_6227);
and U6429 (N_6429,N_6351,N_6285);
nand U6430 (N_6430,N_6259,N_6385);
and U6431 (N_6431,N_6297,N_6308);
and U6432 (N_6432,N_6387,N_6377);
and U6433 (N_6433,N_6334,N_6339);
nand U6434 (N_6434,N_6231,N_6304);
nor U6435 (N_6435,N_6318,N_6311);
and U6436 (N_6436,N_6328,N_6323);
or U6437 (N_6437,N_6294,N_6317);
or U6438 (N_6438,N_6370,N_6322);
and U6439 (N_6439,N_6383,N_6272);
xnor U6440 (N_6440,N_6376,N_6379);
nand U6441 (N_6441,N_6338,N_6271);
nand U6442 (N_6442,N_6230,N_6278);
nor U6443 (N_6443,N_6309,N_6232);
nand U6444 (N_6444,N_6348,N_6316);
and U6445 (N_6445,N_6345,N_6204);
nand U6446 (N_6446,N_6306,N_6229);
and U6447 (N_6447,N_6257,N_6279);
or U6448 (N_6448,N_6373,N_6265);
and U6449 (N_6449,N_6343,N_6398);
or U6450 (N_6450,N_6395,N_6299);
and U6451 (N_6451,N_6365,N_6289);
and U6452 (N_6452,N_6346,N_6397);
nor U6453 (N_6453,N_6252,N_6386);
xnor U6454 (N_6454,N_6399,N_6378);
xor U6455 (N_6455,N_6237,N_6314);
nor U6456 (N_6456,N_6303,N_6208);
nand U6457 (N_6457,N_6313,N_6256);
and U6458 (N_6458,N_6200,N_6382);
nor U6459 (N_6459,N_6312,N_6258);
or U6460 (N_6460,N_6262,N_6389);
nand U6461 (N_6461,N_6284,N_6207);
nor U6462 (N_6462,N_6315,N_6390);
and U6463 (N_6463,N_6287,N_6260);
and U6464 (N_6464,N_6267,N_6277);
xnor U6465 (N_6465,N_6212,N_6235);
and U6466 (N_6466,N_6326,N_6333);
or U6467 (N_6467,N_6310,N_6254);
nor U6468 (N_6468,N_6222,N_6330);
or U6469 (N_6469,N_6363,N_6321);
xor U6470 (N_6470,N_6224,N_6369);
nor U6471 (N_6471,N_6211,N_6214);
xnor U6472 (N_6472,N_6336,N_6245);
xor U6473 (N_6473,N_6250,N_6206);
or U6474 (N_6474,N_6356,N_6216);
xor U6475 (N_6475,N_6353,N_6298);
nor U6476 (N_6476,N_6341,N_6391);
xor U6477 (N_6477,N_6381,N_6269);
xnor U6478 (N_6478,N_6337,N_6273);
and U6479 (N_6479,N_6233,N_6266);
and U6480 (N_6480,N_6268,N_6300);
nand U6481 (N_6481,N_6329,N_6350);
or U6482 (N_6482,N_6349,N_6205);
nand U6483 (N_6483,N_6248,N_6291);
xor U6484 (N_6484,N_6223,N_6243);
and U6485 (N_6485,N_6371,N_6358);
and U6486 (N_6486,N_6361,N_6352);
and U6487 (N_6487,N_6242,N_6384);
nand U6488 (N_6488,N_6319,N_6234);
xor U6489 (N_6489,N_6202,N_6366);
and U6490 (N_6490,N_6392,N_6225);
xor U6491 (N_6491,N_6247,N_6290);
nor U6492 (N_6492,N_6275,N_6286);
and U6493 (N_6493,N_6276,N_6201);
nand U6494 (N_6494,N_6355,N_6357);
and U6495 (N_6495,N_6320,N_6344);
xnor U6496 (N_6496,N_6340,N_6362);
nor U6497 (N_6497,N_6368,N_6203);
and U6498 (N_6498,N_6332,N_6238);
xnor U6499 (N_6499,N_6364,N_6283);
and U6500 (N_6500,N_6391,N_6274);
and U6501 (N_6501,N_6350,N_6389);
or U6502 (N_6502,N_6205,N_6398);
or U6503 (N_6503,N_6394,N_6234);
nor U6504 (N_6504,N_6269,N_6275);
or U6505 (N_6505,N_6228,N_6207);
xor U6506 (N_6506,N_6200,N_6340);
nand U6507 (N_6507,N_6210,N_6326);
xnor U6508 (N_6508,N_6360,N_6281);
xor U6509 (N_6509,N_6219,N_6392);
or U6510 (N_6510,N_6296,N_6213);
nand U6511 (N_6511,N_6342,N_6237);
or U6512 (N_6512,N_6391,N_6347);
nand U6513 (N_6513,N_6255,N_6364);
and U6514 (N_6514,N_6332,N_6209);
xor U6515 (N_6515,N_6332,N_6367);
and U6516 (N_6516,N_6269,N_6272);
and U6517 (N_6517,N_6247,N_6397);
nor U6518 (N_6518,N_6207,N_6260);
or U6519 (N_6519,N_6246,N_6327);
nand U6520 (N_6520,N_6256,N_6241);
or U6521 (N_6521,N_6248,N_6222);
nor U6522 (N_6522,N_6288,N_6375);
xor U6523 (N_6523,N_6296,N_6376);
nand U6524 (N_6524,N_6230,N_6332);
or U6525 (N_6525,N_6333,N_6266);
xnor U6526 (N_6526,N_6250,N_6265);
or U6527 (N_6527,N_6295,N_6300);
xnor U6528 (N_6528,N_6398,N_6299);
and U6529 (N_6529,N_6201,N_6332);
nand U6530 (N_6530,N_6347,N_6392);
nor U6531 (N_6531,N_6258,N_6350);
nand U6532 (N_6532,N_6344,N_6385);
xor U6533 (N_6533,N_6250,N_6398);
nand U6534 (N_6534,N_6300,N_6338);
nor U6535 (N_6535,N_6303,N_6242);
nor U6536 (N_6536,N_6395,N_6377);
nand U6537 (N_6537,N_6386,N_6342);
nor U6538 (N_6538,N_6243,N_6216);
nor U6539 (N_6539,N_6371,N_6211);
and U6540 (N_6540,N_6339,N_6274);
nand U6541 (N_6541,N_6286,N_6278);
or U6542 (N_6542,N_6270,N_6277);
xnor U6543 (N_6543,N_6331,N_6379);
nand U6544 (N_6544,N_6307,N_6368);
and U6545 (N_6545,N_6288,N_6326);
nor U6546 (N_6546,N_6278,N_6242);
or U6547 (N_6547,N_6211,N_6375);
nor U6548 (N_6548,N_6226,N_6314);
nor U6549 (N_6549,N_6211,N_6252);
and U6550 (N_6550,N_6322,N_6232);
nor U6551 (N_6551,N_6316,N_6210);
or U6552 (N_6552,N_6271,N_6333);
nand U6553 (N_6553,N_6375,N_6381);
or U6554 (N_6554,N_6309,N_6301);
or U6555 (N_6555,N_6399,N_6221);
or U6556 (N_6556,N_6306,N_6211);
nand U6557 (N_6557,N_6202,N_6266);
or U6558 (N_6558,N_6268,N_6277);
xor U6559 (N_6559,N_6278,N_6244);
nand U6560 (N_6560,N_6284,N_6300);
xnor U6561 (N_6561,N_6337,N_6263);
xor U6562 (N_6562,N_6234,N_6203);
and U6563 (N_6563,N_6225,N_6307);
xor U6564 (N_6564,N_6306,N_6256);
or U6565 (N_6565,N_6297,N_6282);
nor U6566 (N_6566,N_6246,N_6384);
nor U6567 (N_6567,N_6216,N_6211);
xor U6568 (N_6568,N_6256,N_6275);
and U6569 (N_6569,N_6253,N_6379);
nor U6570 (N_6570,N_6293,N_6291);
xnor U6571 (N_6571,N_6302,N_6228);
nand U6572 (N_6572,N_6235,N_6363);
or U6573 (N_6573,N_6247,N_6274);
and U6574 (N_6574,N_6392,N_6331);
nor U6575 (N_6575,N_6234,N_6351);
xnor U6576 (N_6576,N_6395,N_6371);
nand U6577 (N_6577,N_6399,N_6282);
or U6578 (N_6578,N_6338,N_6282);
nand U6579 (N_6579,N_6226,N_6341);
nand U6580 (N_6580,N_6374,N_6290);
nor U6581 (N_6581,N_6312,N_6241);
or U6582 (N_6582,N_6249,N_6303);
nor U6583 (N_6583,N_6246,N_6396);
and U6584 (N_6584,N_6382,N_6230);
nand U6585 (N_6585,N_6216,N_6380);
and U6586 (N_6586,N_6220,N_6229);
and U6587 (N_6587,N_6277,N_6346);
xor U6588 (N_6588,N_6217,N_6289);
nor U6589 (N_6589,N_6234,N_6395);
nor U6590 (N_6590,N_6293,N_6300);
nand U6591 (N_6591,N_6303,N_6387);
nor U6592 (N_6592,N_6349,N_6240);
xnor U6593 (N_6593,N_6219,N_6262);
or U6594 (N_6594,N_6395,N_6275);
nor U6595 (N_6595,N_6248,N_6236);
xor U6596 (N_6596,N_6273,N_6346);
nand U6597 (N_6597,N_6351,N_6204);
and U6598 (N_6598,N_6373,N_6290);
or U6599 (N_6599,N_6240,N_6362);
and U6600 (N_6600,N_6587,N_6559);
and U6601 (N_6601,N_6598,N_6539);
xor U6602 (N_6602,N_6405,N_6540);
xnor U6603 (N_6603,N_6527,N_6415);
nor U6604 (N_6604,N_6400,N_6445);
nand U6605 (N_6605,N_6463,N_6434);
and U6606 (N_6606,N_6562,N_6537);
or U6607 (N_6607,N_6556,N_6536);
or U6608 (N_6608,N_6471,N_6594);
nor U6609 (N_6609,N_6501,N_6582);
and U6610 (N_6610,N_6494,N_6591);
and U6611 (N_6611,N_6596,N_6451);
nor U6612 (N_6612,N_6488,N_6454);
xor U6613 (N_6613,N_6499,N_6408);
and U6614 (N_6614,N_6507,N_6535);
xnor U6615 (N_6615,N_6517,N_6567);
and U6616 (N_6616,N_6578,N_6418);
nor U6617 (N_6617,N_6541,N_6545);
xnor U6618 (N_6618,N_6424,N_6576);
nor U6619 (N_6619,N_6520,N_6504);
xnor U6620 (N_6620,N_6563,N_6534);
xnor U6621 (N_6621,N_6533,N_6475);
nor U6622 (N_6622,N_6413,N_6416);
or U6623 (N_6623,N_6558,N_6577);
nand U6624 (N_6624,N_6476,N_6436);
or U6625 (N_6625,N_6467,N_6433);
xnor U6626 (N_6626,N_6555,N_6589);
xor U6627 (N_6627,N_6443,N_6538);
nand U6628 (N_6628,N_6457,N_6410);
nand U6629 (N_6629,N_6455,N_6524);
xnor U6630 (N_6630,N_6491,N_6414);
or U6631 (N_6631,N_6561,N_6525);
nor U6632 (N_6632,N_6502,N_6560);
nor U6633 (N_6633,N_6486,N_6490);
or U6634 (N_6634,N_6466,N_6513);
and U6635 (N_6635,N_6484,N_6459);
nor U6636 (N_6636,N_6464,N_6511);
and U6637 (N_6637,N_6532,N_6554);
nor U6638 (N_6638,N_6522,N_6425);
or U6639 (N_6639,N_6575,N_6581);
or U6640 (N_6640,N_6530,N_6421);
or U6641 (N_6641,N_6461,N_6462);
xor U6642 (N_6642,N_6430,N_6429);
nor U6643 (N_6643,N_6487,N_6586);
nand U6644 (N_6644,N_6569,N_6518);
and U6645 (N_6645,N_6460,N_6407);
xor U6646 (N_6646,N_6495,N_6431);
xor U6647 (N_6647,N_6441,N_6428);
nand U6648 (N_6648,N_6550,N_6565);
xor U6649 (N_6649,N_6516,N_6446);
nand U6650 (N_6650,N_6544,N_6588);
or U6651 (N_6651,N_6468,N_6510);
and U6652 (N_6652,N_6478,N_6584);
nor U6653 (N_6653,N_6572,N_6564);
or U6654 (N_6654,N_6595,N_6528);
or U6655 (N_6655,N_6503,N_6523);
nand U6656 (N_6656,N_6448,N_6531);
nor U6657 (N_6657,N_6546,N_6474);
xor U6658 (N_6658,N_6492,N_6482);
nor U6659 (N_6659,N_6479,N_6422);
nor U6660 (N_6660,N_6447,N_6449);
nand U6661 (N_6661,N_6442,N_6401);
nor U6662 (N_6662,N_6472,N_6548);
or U6663 (N_6663,N_6493,N_6549);
xor U6664 (N_6664,N_6409,N_6438);
nor U6665 (N_6665,N_6453,N_6489);
xnor U6666 (N_6666,N_6417,N_6435);
and U6667 (N_6667,N_6406,N_6480);
nand U6668 (N_6668,N_6411,N_6521);
xor U6669 (N_6669,N_6483,N_6485);
nor U6670 (N_6670,N_6426,N_6465);
or U6671 (N_6671,N_6498,N_6571);
xnor U6672 (N_6672,N_6423,N_6419);
and U6673 (N_6673,N_6439,N_6508);
or U6674 (N_6674,N_6512,N_6580);
or U6675 (N_6675,N_6514,N_6568);
xnor U6676 (N_6676,N_6497,N_6402);
or U6677 (N_6677,N_6543,N_6509);
and U6678 (N_6678,N_6566,N_6452);
nor U6679 (N_6679,N_6553,N_6574);
or U6680 (N_6680,N_6579,N_6557);
xor U6681 (N_6681,N_6506,N_6552);
and U6682 (N_6682,N_6420,N_6458);
nand U6683 (N_6683,N_6597,N_6403);
xor U6684 (N_6684,N_6444,N_6500);
xor U6685 (N_6685,N_6481,N_6456);
and U6686 (N_6686,N_6469,N_6440);
xnor U6687 (N_6687,N_6496,N_6551);
or U6688 (N_6688,N_6542,N_6573);
nand U6689 (N_6689,N_6593,N_6412);
nor U6690 (N_6690,N_6515,N_6470);
and U6691 (N_6691,N_6547,N_6590);
or U6692 (N_6692,N_6570,N_6583);
nand U6693 (N_6693,N_6526,N_6519);
and U6694 (N_6694,N_6450,N_6529);
xnor U6695 (N_6695,N_6592,N_6473);
nor U6696 (N_6696,N_6427,N_6437);
nand U6697 (N_6697,N_6432,N_6585);
nor U6698 (N_6698,N_6505,N_6477);
or U6699 (N_6699,N_6599,N_6404);
nor U6700 (N_6700,N_6565,N_6415);
and U6701 (N_6701,N_6491,N_6489);
nor U6702 (N_6702,N_6452,N_6475);
nand U6703 (N_6703,N_6548,N_6509);
xor U6704 (N_6704,N_6584,N_6530);
xor U6705 (N_6705,N_6430,N_6594);
nand U6706 (N_6706,N_6532,N_6455);
xnor U6707 (N_6707,N_6483,N_6596);
nand U6708 (N_6708,N_6575,N_6515);
nand U6709 (N_6709,N_6494,N_6517);
nor U6710 (N_6710,N_6598,N_6584);
and U6711 (N_6711,N_6428,N_6589);
and U6712 (N_6712,N_6405,N_6456);
xnor U6713 (N_6713,N_6582,N_6444);
nand U6714 (N_6714,N_6501,N_6560);
nand U6715 (N_6715,N_6518,N_6540);
xnor U6716 (N_6716,N_6475,N_6574);
xnor U6717 (N_6717,N_6437,N_6538);
xor U6718 (N_6718,N_6443,N_6542);
or U6719 (N_6719,N_6501,N_6492);
nor U6720 (N_6720,N_6512,N_6585);
or U6721 (N_6721,N_6577,N_6556);
nor U6722 (N_6722,N_6418,N_6447);
and U6723 (N_6723,N_6420,N_6452);
or U6724 (N_6724,N_6450,N_6407);
xor U6725 (N_6725,N_6481,N_6542);
xnor U6726 (N_6726,N_6528,N_6477);
nand U6727 (N_6727,N_6561,N_6565);
xnor U6728 (N_6728,N_6591,N_6586);
xnor U6729 (N_6729,N_6408,N_6578);
xor U6730 (N_6730,N_6493,N_6529);
or U6731 (N_6731,N_6567,N_6530);
xor U6732 (N_6732,N_6518,N_6495);
xor U6733 (N_6733,N_6441,N_6545);
and U6734 (N_6734,N_6575,N_6409);
nand U6735 (N_6735,N_6510,N_6444);
nand U6736 (N_6736,N_6432,N_6435);
nor U6737 (N_6737,N_6561,N_6506);
nor U6738 (N_6738,N_6489,N_6492);
and U6739 (N_6739,N_6401,N_6412);
nor U6740 (N_6740,N_6537,N_6563);
xnor U6741 (N_6741,N_6436,N_6561);
and U6742 (N_6742,N_6467,N_6436);
or U6743 (N_6743,N_6508,N_6481);
xnor U6744 (N_6744,N_6409,N_6437);
and U6745 (N_6745,N_6422,N_6438);
xor U6746 (N_6746,N_6483,N_6423);
nor U6747 (N_6747,N_6465,N_6492);
and U6748 (N_6748,N_6461,N_6427);
xnor U6749 (N_6749,N_6444,N_6559);
nor U6750 (N_6750,N_6516,N_6561);
nor U6751 (N_6751,N_6433,N_6566);
xor U6752 (N_6752,N_6595,N_6550);
nand U6753 (N_6753,N_6442,N_6536);
and U6754 (N_6754,N_6485,N_6448);
nand U6755 (N_6755,N_6405,N_6555);
nand U6756 (N_6756,N_6495,N_6566);
or U6757 (N_6757,N_6443,N_6522);
nand U6758 (N_6758,N_6572,N_6489);
or U6759 (N_6759,N_6455,N_6409);
nor U6760 (N_6760,N_6491,N_6594);
and U6761 (N_6761,N_6416,N_6467);
or U6762 (N_6762,N_6444,N_6455);
nand U6763 (N_6763,N_6547,N_6484);
nand U6764 (N_6764,N_6464,N_6424);
nor U6765 (N_6765,N_6511,N_6526);
xnor U6766 (N_6766,N_6595,N_6479);
xor U6767 (N_6767,N_6447,N_6468);
nand U6768 (N_6768,N_6504,N_6424);
and U6769 (N_6769,N_6454,N_6541);
xnor U6770 (N_6770,N_6429,N_6589);
or U6771 (N_6771,N_6406,N_6440);
or U6772 (N_6772,N_6571,N_6429);
and U6773 (N_6773,N_6494,N_6598);
xor U6774 (N_6774,N_6490,N_6521);
nor U6775 (N_6775,N_6514,N_6471);
and U6776 (N_6776,N_6548,N_6455);
nor U6777 (N_6777,N_6581,N_6454);
or U6778 (N_6778,N_6531,N_6579);
or U6779 (N_6779,N_6576,N_6590);
or U6780 (N_6780,N_6487,N_6445);
and U6781 (N_6781,N_6491,N_6512);
and U6782 (N_6782,N_6521,N_6423);
or U6783 (N_6783,N_6434,N_6493);
nand U6784 (N_6784,N_6474,N_6534);
or U6785 (N_6785,N_6537,N_6531);
nor U6786 (N_6786,N_6439,N_6454);
or U6787 (N_6787,N_6511,N_6587);
nand U6788 (N_6788,N_6557,N_6440);
xnor U6789 (N_6789,N_6518,N_6496);
nor U6790 (N_6790,N_6583,N_6448);
xor U6791 (N_6791,N_6544,N_6585);
xor U6792 (N_6792,N_6537,N_6525);
xor U6793 (N_6793,N_6589,N_6511);
or U6794 (N_6794,N_6491,N_6502);
or U6795 (N_6795,N_6435,N_6530);
xor U6796 (N_6796,N_6424,N_6457);
xor U6797 (N_6797,N_6403,N_6537);
xor U6798 (N_6798,N_6414,N_6550);
xor U6799 (N_6799,N_6475,N_6494);
and U6800 (N_6800,N_6688,N_6656);
or U6801 (N_6801,N_6611,N_6632);
and U6802 (N_6802,N_6753,N_6742);
xor U6803 (N_6803,N_6678,N_6710);
nor U6804 (N_6804,N_6712,N_6795);
nand U6805 (N_6805,N_6727,N_6648);
nand U6806 (N_6806,N_6629,N_6711);
xnor U6807 (N_6807,N_6660,N_6713);
nor U6808 (N_6808,N_6769,N_6676);
xnor U6809 (N_6809,N_6681,N_6770);
or U6810 (N_6810,N_6690,N_6621);
or U6811 (N_6811,N_6636,N_6793);
or U6812 (N_6812,N_6798,N_6761);
or U6813 (N_6813,N_6731,N_6708);
xor U6814 (N_6814,N_6689,N_6759);
nor U6815 (N_6815,N_6651,N_6745);
xor U6816 (N_6816,N_6679,N_6624);
xor U6817 (N_6817,N_6645,N_6669);
xnor U6818 (N_6818,N_6735,N_6718);
nand U6819 (N_6819,N_6622,N_6715);
xor U6820 (N_6820,N_6744,N_6788);
nand U6821 (N_6821,N_6685,N_6606);
xor U6822 (N_6822,N_6767,N_6739);
and U6823 (N_6823,N_6796,N_6618);
nand U6824 (N_6824,N_6625,N_6650);
xor U6825 (N_6825,N_6641,N_6702);
and U6826 (N_6826,N_6655,N_6757);
and U6827 (N_6827,N_6719,N_6644);
and U6828 (N_6828,N_6671,N_6703);
nor U6829 (N_6829,N_6756,N_6608);
nor U6830 (N_6830,N_6609,N_6615);
nor U6831 (N_6831,N_6764,N_6605);
nand U6832 (N_6832,N_6643,N_6707);
or U6833 (N_6833,N_6649,N_6630);
xor U6834 (N_6834,N_6682,N_6777);
and U6835 (N_6835,N_6674,N_6693);
or U6836 (N_6836,N_6728,N_6602);
nor U6837 (N_6837,N_6662,N_6696);
xnor U6838 (N_6838,N_6684,N_6746);
or U6839 (N_6839,N_6705,N_6738);
nand U6840 (N_6840,N_6677,N_6785);
or U6841 (N_6841,N_6610,N_6781);
and U6842 (N_6842,N_6659,N_6663);
or U6843 (N_6843,N_6638,N_6613);
nor U6844 (N_6844,N_6791,N_6751);
or U6845 (N_6845,N_6646,N_6619);
nor U6846 (N_6846,N_6779,N_6792);
nor U6847 (N_6847,N_6771,N_6760);
or U6848 (N_6848,N_6640,N_6787);
nand U6849 (N_6849,N_6763,N_6635);
xnor U6850 (N_6850,N_6673,N_6725);
nand U6851 (N_6851,N_6691,N_6672);
xor U6852 (N_6852,N_6747,N_6698);
xnor U6853 (N_6853,N_6786,N_6748);
nand U6854 (N_6854,N_6607,N_6637);
nand U6855 (N_6855,N_6680,N_6752);
or U6856 (N_6856,N_6765,N_6775);
and U6857 (N_6857,N_6692,N_6667);
nor U6858 (N_6858,N_6665,N_6749);
nor U6859 (N_6859,N_6634,N_6780);
or U6860 (N_6860,N_6612,N_6776);
xnor U6861 (N_6861,N_6716,N_6603);
and U6862 (N_6862,N_6784,N_6697);
or U6863 (N_6863,N_6620,N_6730);
or U6864 (N_6864,N_6714,N_6750);
xor U6865 (N_6865,N_6670,N_6709);
nand U6866 (N_6866,N_6726,N_6724);
nand U6867 (N_6867,N_6687,N_6740);
or U6868 (N_6868,N_6623,N_6661);
or U6869 (N_6869,N_6686,N_6627);
nor U6870 (N_6870,N_6732,N_6658);
nand U6871 (N_6871,N_6754,N_6699);
nor U6872 (N_6872,N_6729,N_6652);
or U6873 (N_6873,N_6675,N_6668);
and U6874 (N_6874,N_6664,N_6666);
and U6875 (N_6875,N_6789,N_6701);
or U6876 (N_6876,N_6799,N_6723);
or U6877 (N_6877,N_6790,N_6794);
nor U6878 (N_6878,N_6633,N_6741);
xor U6879 (N_6879,N_6720,N_6683);
or U6880 (N_6880,N_6774,N_6654);
nor U6881 (N_6881,N_6736,N_6604);
nand U6882 (N_6882,N_6700,N_6766);
xor U6883 (N_6883,N_6755,N_6642);
nor U6884 (N_6884,N_6617,N_6783);
nand U6885 (N_6885,N_6778,N_6600);
nor U6886 (N_6886,N_6782,N_6628);
nand U6887 (N_6887,N_6639,N_6743);
or U6888 (N_6888,N_6737,N_6797);
and U6889 (N_6889,N_6694,N_6758);
nor U6890 (N_6890,N_6601,N_6704);
nor U6891 (N_6891,N_6657,N_6722);
or U6892 (N_6892,N_6647,N_6614);
and U6893 (N_6893,N_6631,N_6773);
and U6894 (N_6894,N_6706,N_6717);
and U6895 (N_6895,N_6695,N_6733);
nor U6896 (N_6896,N_6768,N_6772);
nor U6897 (N_6897,N_6626,N_6616);
xnor U6898 (N_6898,N_6721,N_6734);
xnor U6899 (N_6899,N_6762,N_6653);
and U6900 (N_6900,N_6749,N_6727);
or U6901 (N_6901,N_6664,N_6727);
nand U6902 (N_6902,N_6718,N_6741);
nand U6903 (N_6903,N_6646,N_6601);
nor U6904 (N_6904,N_6630,N_6692);
or U6905 (N_6905,N_6797,N_6789);
or U6906 (N_6906,N_6690,N_6649);
nand U6907 (N_6907,N_6600,N_6744);
and U6908 (N_6908,N_6694,N_6628);
nand U6909 (N_6909,N_6650,N_6728);
xor U6910 (N_6910,N_6611,N_6656);
or U6911 (N_6911,N_6739,N_6635);
nor U6912 (N_6912,N_6760,N_6744);
and U6913 (N_6913,N_6791,N_6692);
and U6914 (N_6914,N_6671,N_6799);
and U6915 (N_6915,N_6613,N_6772);
and U6916 (N_6916,N_6657,N_6689);
nor U6917 (N_6917,N_6629,N_6654);
or U6918 (N_6918,N_6611,N_6718);
and U6919 (N_6919,N_6777,N_6675);
and U6920 (N_6920,N_6630,N_6686);
xor U6921 (N_6921,N_6688,N_6682);
xnor U6922 (N_6922,N_6627,N_6697);
or U6923 (N_6923,N_6785,N_6669);
xor U6924 (N_6924,N_6696,N_6604);
or U6925 (N_6925,N_6695,N_6603);
xor U6926 (N_6926,N_6765,N_6645);
nand U6927 (N_6927,N_6638,N_6672);
and U6928 (N_6928,N_6698,N_6651);
nor U6929 (N_6929,N_6635,N_6657);
nand U6930 (N_6930,N_6671,N_6733);
nand U6931 (N_6931,N_6660,N_6718);
nand U6932 (N_6932,N_6799,N_6701);
nor U6933 (N_6933,N_6613,N_6706);
nor U6934 (N_6934,N_6794,N_6771);
nand U6935 (N_6935,N_6683,N_6633);
xor U6936 (N_6936,N_6793,N_6641);
nor U6937 (N_6937,N_6713,N_6714);
nor U6938 (N_6938,N_6652,N_6622);
nand U6939 (N_6939,N_6704,N_6738);
nand U6940 (N_6940,N_6734,N_6784);
xor U6941 (N_6941,N_6775,N_6691);
nand U6942 (N_6942,N_6790,N_6609);
and U6943 (N_6943,N_6757,N_6618);
nor U6944 (N_6944,N_6739,N_6738);
nor U6945 (N_6945,N_6623,N_6645);
nand U6946 (N_6946,N_6646,N_6778);
nor U6947 (N_6947,N_6692,N_6684);
nor U6948 (N_6948,N_6753,N_6663);
or U6949 (N_6949,N_6640,N_6608);
or U6950 (N_6950,N_6675,N_6658);
or U6951 (N_6951,N_6772,N_6698);
xor U6952 (N_6952,N_6791,N_6760);
and U6953 (N_6953,N_6780,N_6744);
nor U6954 (N_6954,N_6645,N_6694);
and U6955 (N_6955,N_6665,N_6795);
or U6956 (N_6956,N_6622,N_6692);
nand U6957 (N_6957,N_6642,N_6677);
nor U6958 (N_6958,N_6799,N_6734);
xor U6959 (N_6959,N_6765,N_6700);
nor U6960 (N_6960,N_6781,N_6668);
nor U6961 (N_6961,N_6786,N_6780);
nand U6962 (N_6962,N_6786,N_6652);
or U6963 (N_6963,N_6630,N_6659);
nand U6964 (N_6964,N_6747,N_6708);
or U6965 (N_6965,N_6697,N_6667);
xor U6966 (N_6966,N_6643,N_6691);
or U6967 (N_6967,N_6719,N_6782);
or U6968 (N_6968,N_6755,N_6713);
nand U6969 (N_6969,N_6661,N_6625);
xor U6970 (N_6970,N_6713,N_6722);
xor U6971 (N_6971,N_6739,N_6608);
nor U6972 (N_6972,N_6747,N_6714);
or U6973 (N_6973,N_6732,N_6726);
nand U6974 (N_6974,N_6660,N_6641);
nand U6975 (N_6975,N_6742,N_6610);
xor U6976 (N_6976,N_6706,N_6657);
xor U6977 (N_6977,N_6686,N_6682);
or U6978 (N_6978,N_6612,N_6621);
or U6979 (N_6979,N_6650,N_6744);
xnor U6980 (N_6980,N_6774,N_6749);
xor U6981 (N_6981,N_6673,N_6778);
or U6982 (N_6982,N_6648,N_6623);
nand U6983 (N_6983,N_6777,N_6678);
and U6984 (N_6984,N_6735,N_6643);
nand U6985 (N_6985,N_6756,N_6715);
or U6986 (N_6986,N_6636,N_6619);
xnor U6987 (N_6987,N_6773,N_6692);
xnor U6988 (N_6988,N_6628,N_6673);
nand U6989 (N_6989,N_6615,N_6658);
and U6990 (N_6990,N_6695,N_6797);
nor U6991 (N_6991,N_6771,N_6676);
nand U6992 (N_6992,N_6635,N_6670);
nand U6993 (N_6993,N_6651,N_6798);
nand U6994 (N_6994,N_6677,N_6703);
and U6995 (N_6995,N_6725,N_6606);
nand U6996 (N_6996,N_6715,N_6709);
nor U6997 (N_6997,N_6719,N_6759);
and U6998 (N_6998,N_6768,N_6777);
nor U6999 (N_6999,N_6723,N_6615);
nor U7000 (N_7000,N_6880,N_6952);
or U7001 (N_7001,N_6827,N_6822);
xnor U7002 (N_7002,N_6962,N_6966);
xnor U7003 (N_7003,N_6959,N_6879);
and U7004 (N_7004,N_6918,N_6988);
xnor U7005 (N_7005,N_6850,N_6979);
nand U7006 (N_7006,N_6964,N_6810);
and U7007 (N_7007,N_6924,N_6968);
xnor U7008 (N_7008,N_6895,N_6838);
nand U7009 (N_7009,N_6896,N_6871);
xnor U7010 (N_7010,N_6837,N_6969);
and U7011 (N_7011,N_6889,N_6870);
nor U7012 (N_7012,N_6956,N_6971);
nand U7013 (N_7013,N_6851,N_6843);
nor U7014 (N_7014,N_6912,N_6967);
or U7015 (N_7015,N_6937,N_6861);
or U7016 (N_7016,N_6940,N_6991);
nand U7017 (N_7017,N_6925,N_6834);
or U7018 (N_7018,N_6887,N_6831);
or U7019 (N_7019,N_6905,N_6929);
or U7020 (N_7020,N_6856,N_6865);
nand U7021 (N_7021,N_6938,N_6902);
and U7022 (N_7022,N_6922,N_6854);
nor U7023 (N_7023,N_6826,N_6839);
nor U7024 (N_7024,N_6898,N_6953);
and U7025 (N_7025,N_6951,N_6867);
or U7026 (N_7026,N_6993,N_6919);
xor U7027 (N_7027,N_6981,N_6985);
nor U7028 (N_7028,N_6913,N_6823);
and U7029 (N_7029,N_6897,N_6803);
and U7030 (N_7030,N_6946,N_6933);
xnor U7031 (N_7031,N_6884,N_6936);
or U7032 (N_7032,N_6890,N_6868);
xnor U7033 (N_7033,N_6947,N_6883);
nand U7034 (N_7034,N_6930,N_6894);
or U7035 (N_7035,N_6802,N_6833);
and U7036 (N_7036,N_6804,N_6998);
nor U7037 (N_7037,N_6961,N_6858);
or U7038 (N_7038,N_6876,N_6806);
nand U7039 (N_7039,N_6965,N_6943);
xor U7040 (N_7040,N_6974,N_6888);
and U7041 (N_7041,N_6832,N_6800);
and U7042 (N_7042,N_6877,N_6817);
nor U7043 (N_7043,N_6927,N_6801);
and U7044 (N_7044,N_6916,N_6881);
nor U7045 (N_7045,N_6960,N_6875);
or U7046 (N_7046,N_6992,N_6885);
nand U7047 (N_7047,N_6983,N_6907);
and U7048 (N_7048,N_6954,N_6848);
nor U7049 (N_7049,N_6915,N_6872);
nand U7050 (N_7050,N_6909,N_6892);
nor U7051 (N_7051,N_6824,N_6805);
and U7052 (N_7052,N_6821,N_6977);
and U7053 (N_7053,N_6852,N_6809);
xor U7054 (N_7054,N_6814,N_6934);
nand U7055 (N_7055,N_6862,N_6980);
nor U7056 (N_7056,N_6939,N_6944);
nand U7057 (N_7057,N_6845,N_6941);
xor U7058 (N_7058,N_6928,N_6926);
nand U7059 (N_7059,N_6853,N_6982);
and U7060 (N_7060,N_6948,N_6958);
or U7061 (N_7061,N_6835,N_6878);
nor U7062 (N_7062,N_6857,N_6931);
and U7063 (N_7063,N_6950,N_6893);
xor U7064 (N_7064,N_6975,N_6906);
nand U7065 (N_7065,N_6828,N_6808);
or U7066 (N_7066,N_6997,N_6874);
and U7067 (N_7067,N_6914,N_6904);
nand U7068 (N_7068,N_6999,N_6844);
nor U7069 (N_7069,N_6990,N_6860);
nand U7070 (N_7070,N_6842,N_6847);
xor U7071 (N_7071,N_6996,N_6841);
and U7072 (N_7072,N_6923,N_6942);
nor U7073 (N_7073,N_6970,N_6811);
xnor U7074 (N_7074,N_6989,N_6921);
or U7075 (N_7075,N_6978,N_6816);
and U7076 (N_7076,N_6866,N_6908);
xor U7077 (N_7077,N_6987,N_6899);
nand U7078 (N_7078,N_6869,N_6829);
or U7079 (N_7079,N_6986,N_6955);
nand U7080 (N_7080,N_6818,N_6886);
xor U7081 (N_7081,N_6836,N_6945);
or U7082 (N_7082,N_6932,N_6846);
or U7083 (N_7083,N_6995,N_6949);
or U7084 (N_7084,N_6920,N_6864);
or U7085 (N_7085,N_6807,N_6900);
xnor U7086 (N_7086,N_6830,N_6882);
nor U7087 (N_7087,N_6820,N_6910);
nor U7088 (N_7088,N_6973,N_6957);
xnor U7089 (N_7089,N_6891,N_6859);
nand U7090 (N_7090,N_6849,N_6917);
and U7091 (N_7091,N_6972,N_6825);
xor U7092 (N_7092,N_6963,N_6911);
or U7093 (N_7093,N_6873,N_6935);
nand U7094 (N_7094,N_6855,N_6813);
xor U7095 (N_7095,N_6840,N_6994);
xor U7096 (N_7096,N_6815,N_6819);
or U7097 (N_7097,N_6976,N_6812);
nor U7098 (N_7098,N_6863,N_6901);
and U7099 (N_7099,N_6903,N_6984);
and U7100 (N_7100,N_6863,N_6946);
or U7101 (N_7101,N_6982,N_6911);
nand U7102 (N_7102,N_6828,N_6823);
or U7103 (N_7103,N_6954,N_6946);
and U7104 (N_7104,N_6875,N_6818);
and U7105 (N_7105,N_6876,N_6872);
or U7106 (N_7106,N_6836,N_6833);
and U7107 (N_7107,N_6996,N_6957);
xnor U7108 (N_7108,N_6985,N_6871);
and U7109 (N_7109,N_6827,N_6955);
or U7110 (N_7110,N_6817,N_6972);
and U7111 (N_7111,N_6926,N_6894);
nor U7112 (N_7112,N_6867,N_6826);
xnor U7113 (N_7113,N_6930,N_6933);
and U7114 (N_7114,N_6976,N_6888);
and U7115 (N_7115,N_6901,N_6992);
nand U7116 (N_7116,N_6869,N_6951);
and U7117 (N_7117,N_6831,N_6886);
or U7118 (N_7118,N_6833,N_6831);
nor U7119 (N_7119,N_6840,N_6918);
and U7120 (N_7120,N_6893,N_6818);
and U7121 (N_7121,N_6929,N_6945);
or U7122 (N_7122,N_6989,N_6932);
nor U7123 (N_7123,N_6983,N_6908);
nor U7124 (N_7124,N_6841,N_6882);
or U7125 (N_7125,N_6934,N_6988);
nand U7126 (N_7126,N_6860,N_6994);
nand U7127 (N_7127,N_6933,N_6869);
nor U7128 (N_7128,N_6990,N_6998);
xor U7129 (N_7129,N_6988,N_6933);
and U7130 (N_7130,N_6966,N_6922);
or U7131 (N_7131,N_6966,N_6970);
nor U7132 (N_7132,N_6972,N_6983);
nor U7133 (N_7133,N_6989,N_6999);
nor U7134 (N_7134,N_6936,N_6916);
or U7135 (N_7135,N_6920,N_6917);
and U7136 (N_7136,N_6878,N_6952);
nor U7137 (N_7137,N_6803,N_6900);
nor U7138 (N_7138,N_6888,N_6883);
or U7139 (N_7139,N_6841,N_6820);
nor U7140 (N_7140,N_6957,N_6944);
and U7141 (N_7141,N_6893,N_6857);
nor U7142 (N_7142,N_6899,N_6849);
xnor U7143 (N_7143,N_6877,N_6963);
xor U7144 (N_7144,N_6930,N_6809);
nor U7145 (N_7145,N_6866,N_6934);
nor U7146 (N_7146,N_6870,N_6806);
xnor U7147 (N_7147,N_6854,N_6907);
xnor U7148 (N_7148,N_6992,N_6953);
nand U7149 (N_7149,N_6859,N_6990);
nand U7150 (N_7150,N_6942,N_6843);
xnor U7151 (N_7151,N_6897,N_6804);
or U7152 (N_7152,N_6984,N_6870);
nand U7153 (N_7153,N_6864,N_6899);
nand U7154 (N_7154,N_6907,N_6874);
or U7155 (N_7155,N_6819,N_6984);
or U7156 (N_7156,N_6879,N_6976);
xnor U7157 (N_7157,N_6900,N_6933);
xnor U7158 (N_7158,N_6907,N_6895);
nor U7159 (N_7159,N_6840,N_6806);
and U7160 (N_7160,N_6913,N_6874);
nand U7161 (N_7161,N_6876,N_6854);
nor U7162 (N_7162,N_6904,N_6919);
and U7163 (N_7163,N_6919,N_6966);
xnor U7164 (N_7164,N_6918,N_6822);
nand U7165 (N_7165,N_6950,N_6998);
xnor U7166 (N_7166,N_6893,N_6961);
nor U7167 (N_7167,N_6849,N_6832);
nand U7168 (N_7168,N_6822,N_6800);
and U7169 (N_7169,N_6962,N_6939);
or U7170 (N_7170,N_6954,N_6888);
nand U7171 (N_7171,N_6896,N_6843);
xor U7172 (N_7172,N_6956,N_6936);
nand U7173 (N_7173,N_6953,N_6981);
nor U7174 (N_7174,N_6910,N_6848);
or U7175 (N_7175,N_6831,N_6815);
or U7176 (N_7176,N_6984,N_6947);
and U7177 (N_7177,N_6811,N_6979);
nand U7178 (N_7178,N_6906,N_6832);
nand U7179 (N_7179,N_6823,N_6948);
xor U7180 (N_7180,N_6806,N_6970);
or U7181 (N_7181,N_6846,N_6844);
nor U7182 (N_7182,N_6843,N_6845);
and U7183 (N_7183,N_6965,N_6914);
or U7184 (N_7184,N_6842,N_6935);
or U7185 (N_7185,N_6912,N_6945);
nor U7186 (N_7186,N_6915,N_6908);
nor U7187 (N_7187,N_6848,N_6836);
nor U7188 (N_7188,N_6936,N_6890);
nor U7189 (N_7189,N_6993,N_6915);
nor U7190 (N_7190,N_6816,N_6906);
nor U7191 (N_7191,N_6987,N_6960);
and U7192 (N_7192,N_6826,N_6963);
xor U7193 (N_7193,N_6826,N_6964);
nor U7194 (N_7194,N_6928,N_6809);
nor U7195 (N_7195,N_6864,N_6871);
nand U7196 (N_7196,N_6974,N_6876);
or U7197 (N_7197,N_6891,N_6960);
xnor U7198 (N_7198,N_6875,N_6985);
and U7199 (N_7199,N_6919,N_6935);
nor U7200 (N_7200,N_7133,N_7021);
or U7201 (N_7201,N_7125,N_7178);
or U7202 (N_7202,N_7175,N_7012);
xnor U7203 (N_7203,N_7101,N_7093);
or U7204 (N_7204,N_7030,N_7186);
nand U7205 (N_7205,N_7142,N_7194);
and U7206 (N_7206,N_7090,N_7141);
xor U7207 (N_7207,N_7193,N_7097);
nand U7208 (N_7208,N_7129,N_7183);
or U7209 (N_7209,N_7026,N_7004);
nand U7210 (N_7210,N_7076,N_7058);
or U7211 (N_7211,N_7078,N_7050);
nand U7212 (N_7212,N_7109,N_7065);
and U7213 (N_7213,N_7046,N_7198);
xnor U7214 (N_7214,N_7054,N_7002);
and U7215 (N_7215,N_7067,N_7185);
xor U7216 (N_7216,N_7039,N_7092);
or U7217 (N_7217,N_7044,N_7195);
xor U7218 (N_7218,N_7075,N_7149);
xor U7219 (N_7219,N_7118,N_7098);
nand U7220 (N_7220,N_7094,N_7061);
or U7221 (N_7221,N_7174,N_7048);
nand U7222 (N_7222,N_7182,N_7152);
xnor U7223 (N_7223,N_7187,N_7196);
xor U7224 (N_7224,N_7055,N_7188);
or U7225 (N_7225,N_7057,N_7199);
or U7226 (N_7226,N_7104,N_7132);
and U7227 (N_7227,N_7147,N_7031);
nor U7228 (N_7228,N_7179,N_7045);
nor U7229 (N_7229,N_7120,N_7121);
or U7230 (N_7230,N_7167,N_7116);
xnor U7231 (N_7231,N_7134,N_7144);
and U7232 (N_7232,N_7003,N_7018);
nor U7233 (N_7233,N_7153,N_7115);
and U7234 (N_7234,N_7009,N_7056);
or U7235 (N_7235,N_7191,N_7114);
nor U7236 (N_7236,N_7001,N_7105);
xor U7237 (N_7237,N_7190,N_7034);
and U7238 (N_7238,N_7015,N_7166);
nor U7239 (N_7239,N_7028,N_7165);
nor U7240 (N_7240,N_7017,N_7135);
nand U7241 (N_7241,N_7137,N_7177);
and U7242 (N_7242,N_7029,N_7108);
or U7243 (N_7243,N_7027,N_7111);
nand U7244 (N_7244,N_7085,N_7041);
nand U7245 (N_7245,N_7163,N_7047);
nor U7246 (N_7246,N_7155,N_7019);
xnor U7247 (N_7247,N_7042,N_7176);
and U7248 (N_7248,N_7084,N_7119);
nand U7249 (N_7249,N_7036,N_7126);
nand U7250 (N_7250,N_7145,N_7130);
xnor U7251 (N_7251,N_7032,N_7140);
and U7252 (N_7252,N_7181,N_7184);
and U7253 (N_7253,N_7071,N_7136);
nor U7254 (N_7254,N_7005,N_7049);
and U7255 (N_7255,N_7106,N_7095);
and U7256 (N_7256,N_7102,N_7148);
xor U7257 (N_7257,N_7197,N_7007);
nor U7258 (N_7258,N_7087,N_7025);
nor U7259 (N_7259,N_7127,N_7171);
nand U7260 (N_7260,N_7100,N_7173);
and U7261 (N_7261,N_7096,N_7023);
xor U7262 (N_7262,N_7051,N_7022);
nand U7263 (N_7263,N_7064,N_7008);
nor U7264 (N_7264,N_7037,N_7124);
and U7265 (N_7265,N_7086,N_7052);
and U7266 (N_7266,N_7139,N_7162);
nor U7267 (N_7267,N_7103,N_7151);
and U7268 (N_7268,N_7082,N_7013);
or U7269 (N_7269,N_7169,N_7156);
or U7270 (N_7270,N_7099,N_7040);
nand U7271 (N_7271,N_7157,N_7160);
nor U7272 (N_7272,N_7035,N_7158);
nand U7273 (N_7273,N_7091,N_7168);
xnor U7274 (N_7274,N_7062,N_7146);
and U7275 (N_7275,N_7110,N_7117);
xor U7276 (N_7276,N_7006,N_7072);
or U7277 (N_7277,N_7066,N_7107);
nor U7278 (N_7278,N_7159,N_7138);
xor U7279 (N_7279,N_7189,N_7123);
xor U7280 (N_7280,N_7070,N_7077);
xor U7281 (N_7281,N_7073,N_7088);
or U7282 (N_7282,N_7128,N_7081);
or U7283 (N_7283,N_7113,N_7011);
nand U7284 (N_7284,N_7080,N_7000);
or U7285 (N_7285,N_7164,N_7014);
and U7286 (N_7286,N_7038,N_7079);
and U7287 (N_7287,N_7154,N_7172);
or U7288 (N_7288,N_7059,N_7143);
xor U7289 (N_7289,N_7161,N_7010);
and U7290 (N_7290,N_7016,N_7083);
xor U7291 (N_7291,N_7033,N_7170);
or U7292 (N_7292,N_7063,N_7043);
nor U7293 (N_7293,N_7180,N_7053);
and U7294 (N_7294,N_7024,N_7069);
nand U7295 (N_7295,N_7192,N_7060);
xor U7296 (N_7296,N_7020,N_7131);
and U7297 (N_7297,N_7150,N_7068);
or U7298 (N_7298,N_7112,N_7089);
nand U7299 (N_7299,N_7074,N_7122);
nor U7300 (N_7300,N_7068,N_7174);
and U7301 (N_7301,N_7190,N_7097);
nand U7302 (N_7302,N_7055,N_7176);
or U7303 (N_7303,N_7035,N_7152);
xor U7304 (N_7304,N_7040,N_7130);
nor U7305 (N_7305,N_7046,N_7098);
nand U7306 (N_7306,N_7021,N_7064);
and U7307 (N_7307,N_7035,N_7098);
or U7308 (N_7308,N_7089,N_7165);
nor U7309 (N_7309,N_7113,N_7047);
nor U7310 (N_7310,N_7125,N_7061);
and U7311 (N_7311,N_7080,N_7052);
nand U7312 (N_7312,N_7024,N_7085);
xor U7313 (N_7313,N_7001,N_7041);
nor U7314 (N_7314,N_7040,N_7092);
nand U7315 (N_7315,N_7099,N_7043);
and U7316 (N_7316,N_7114,N_7148);
and U7317 (N_7317,N_7087,N_7172);
nor U7318 (N_7318,N_7006,N_7035);
xnor U7319 (N_7319,N_7011,N_7025);
xnor U7320 (N_7320,N_7114,N_7093);
and U7321 (N_7321,N_7194,N_7051);
and U7322 (N_7322,N_7049,N_7110);
nor U7323 (N_7323,N_7152,N_7015);
nand U7324 (N_7324,N_7198,N_7192);
nand U7325 (N_7325,N_7180,N_7014);
nand U7326 (N_7326,N_7048,N_7030);
or U7327 (N_7327,N_7108,N_7198);
nand U7328 (N_7328,N_7192,N_7170);
and U7329 (N_7329,N_7023,N_7136);
or U7330 (N_7330,N_7179,N_7149);
and U7331 (N_7331,N_7117,N_7084);
or U7332 (N_7332,N_7083,N_7145);
xnor U7333 (N_7333,N_7108,N_7025);
nor U7334 (N_7334,N_7166,N_7092);
xnor U7335 (N_7335,N_7034,N_7151);
nand U7336 (N_7336,N_7125,N_7113);
and U7337 (N_7337,N_7041,N_7178);
and U7338 (N_7338,N_7005,N_7092);
nor U7339 (N_7339,N_7094,N_7085);
xor U7340 (N_7340,N_7145,N_7154);
and U7341 (N_7341,N_7148,N_7146);
or U7342 (N_7342,N_7017,N_7037);
and U7343 (N_7343,N_7004,N_7139);
nand U7344 (N_7344,N_7192,N_7059);
nand U7345 (N_7345,N_7052,N_7061);
nand U7346 (N_7346,N_7116,N_7071);
and U7347 (N_7347,N_7168,N_7113);
nor U7348 (N_7348,N_7108,N_7169);
xor U7349 (N_7349,N_7120,N_7140);
xnor U7350 (N_7350,N_7111,N_7007);
or U7351 (N_7351,N_7050,N_7092);
or U7352 (N_7352,N_7189,N_7178);
nor U7353 (N_7353,N_7174,N_7028);
and U7354 (N_7354,N_7165,N_7035);
nand U7355 (N_7355,N_7067,N_7156);
or U7356 (N_7356,N_7014,N_7026);
xor U7357 (N_7357,N_7049,N_7000);
and U7358 (N_7358,N_7099,N_7147);
nor U7359 (N_7359,N_7199,N_7106);
and U7360 (N_7360,N_7177,N_7087);
and U7361 (N_7361,N_7109,N_7040);
or U7362 (N_7362,N_7154,N_7059);
xor U7363 (N_7363,N_7134,N_7140);
xor U7364 (N_7364,N_7126,N_7079);
nand U7365 (N_7365,N_7091,N_7145);
nor U7366 (N_7366,N_7030,N_7111);
and U7367 (N_7367,N_7142,N_7137);
nand U7368 (N_7368,N_7038,N_7066);
nand U7369 (N_7369,N_7086,N_7024);
and U7370 (N_7370,N_7004,N_7064);
nor U7371 (N_7371,N_7004,N_7045);
nand U7372 (N_7372,N_7069,N_7142);
or U7373 (N_7373,N_7106,N_7124);
nand U7374 (N_7374,N_7086,N_7034);
or U7375 (N_7375,N_7055,N_7042);
nand U7376 (N_7376,N_7067,N_7184);
nand U7377 (N_7377,N_7090,N_7027);
or U7378 (N_7378,N_7141,N_7112);
nand U7379 (N_7379,N_7165,N_7154);
or U7380 (N_7380,N_7076,N_7189);
xor U7381 (N_7381,N_7100,N_7028);
xor U7382 (N_7382,N_7074,N_7108);
nor U7383 (N_7383,N_7099,N_7093);
nor U7384 (N_7384,N_7117,N_7061);
and U7385 (N_7385,N_7027,N_7001);
and U7386 (N_7386,N_7083,N_7126);
xnor U7387 (N_7387,N_7164,N_7066);
nand U7388 (N_7388,N_7093,N_7102);
nand U7389 (N_7389,N_7077,N_7050);
xor U7390 (N_7390,N_7193,N_7094);
xor U7391 (N_7391,N_7101,N_7167);
and U7392 (N_7392,N_7199,N_7091);
nor U7393 (N_7393,N_7183,N_7105);
nand U7394 (N_7394,N_7057,N_7049);
xnor U7395 (N_7395,N_7044,N_7052);
and U7396 (N_7396,N_7193,N_7120);
nand U7397 (N_7397,N_7030,N_7026);
nor U7398 (N_7398,N_7048,N_7084);
nand U7399 (N_7399,N_7010,N_7121);
and U7400 (N_7400,N_7276,N_7274);
xor U7401 (N_7401,N_7325,N_7214);
and U7402 (N_7402,N_7388,N_7207);
and U7403 (N_7403,N_7370,N_7350);
and U7404 (N_7404,N_7314,N_7260);
or U7405 (N_7405,N_7375,N_7342);
xnor U7406 (N_7406,N_7265,N_7258);
or U7407 (N_7407,N_7262,N_7346);
nand U7408 (N_7408,N_7241,N_7226);
xor U7409 (N_7409,N_7334,N_7252);
nor U7410 (N_7410,N_7316,N_7259);
xor U7411 (N_7411,N_7392,N_7237);
nand U7412 (N_7412,N_7284,N_7385);
xor U7413 (N_7413,N_7233,N_7387);
xnor U7414 (N_7414,N_7249,N_7285);
xor U7415 (N_7415,N_7315,N_7320);
and U7416 (N_7416,N_7381,N_7277);
and U7417 (N_7417,N_7264,N_7205);
and U7418 (N_7418,N_7296,N_7273);
nand U7419 (N_7419,N_7253,N_7229);
nor U7420 (N_7420,N_7337,N_7328);
or U7421 (N_7421,N_7246,N_7291);
xor U7422 (N_7422,N_7224,N_7216);
nand U7423 (N_7423,N_7394,N_7228);
nand U7424 (N_7424,N_7357,N_7335);
xnor U7425 (N_7425,N_7303,N_7365);
xor U7426 (N_7426,N_7343,N_7242);
nand U7427 (N_7427,N_7379,N_7297);
or U7428 (N_7428,N_7222,N_7359);
or U7429 (N_7429,N_7283,N_7338);
nor U7430 (N_7430,N_7321,N_7332);
nand U7431 (N_7431,N_7386,N_7256);
and U7432 (N_7432,N_7368,N_7373);
xnor U7433 (N_7433,N_7355,N_7358);
or U7434 (N_7434,N_7352,N_7298);
or U7435 (N_7435,N_7268,N_7353);
xor U7436 (N_7436,N_7254,N_7371);
or U7437 (N_7437,N_7272,N_7391);
nand U7438 (N_7438,N_7289,N_7309);
nand U7439 (N_7439,N_7200,N_7356);
or U7440 (N_7440,N_7317,N_7263);
nand U7441 (N_7441,N_7323,N_7267);
nand U7442 (N_7442,N_7327,N_7305);
xor U7443 (N_7443,N_7251,N_7248);
or U7444 (N_7444,N_7279,N_7225);
and U7445 (N_7445,N_7302,N_7329);
xnor U7446 (N_7446,N_7390,N_7333);
and U7447 (N_7447,N_7310,N_7270);
nand U7448 (N_7448,N_7372,N_7217);
xnor U7449 (N_7449,N_7301,N_7257);
nor U7450 (N_7450,N_7243,N_7290);
or U7451 (N_7451,N_7378,N_7347);
nor U7452 (N_7452,N_7396,N_7326);
xnor U7453 (N_7453,N_7204,N_7322);
nand U7454 (N_7454,N_7215,N_7245);
nor U7455 (N_7455,N_7269,N_7398);
or U7456 (N_7456,N_7354,N_7219);
xor U7457 (N_7457,N_7397,N_7348);
nand U7458 (N_7458,N_7367,N_7300);
xnor U7459 (N_7459,N_7203,N_7230);
xor U7460 (N_7460,N_7295,N_7306);
or U7461 (N_7461,N_7223,N_7282);
nor U7462 (N_7462,N_7374,N_7210);
and U7463 (N_7463,N_7221,N_7255);
and U7464 (N_7464,N_7362,N_7336);
and U7465 (N_7465,N_7324,N_7287);
or U7466 (N_7466,N_7201,N_7312);
nor U7467 (N_7467,N_7232,N_7363);
or U7468 (N_7468,N_7384,N_7345);
nand U7469 (N_7469,N_7280,N_7308);
nor U7470 (N_7470,N_7261,N_7208);
nor U7471 (N_7471,N_7202,N_7244);
nand U7472 (N_7472,N_7318,N_7393);
nor U7473 (N_7473,N_7389,N_7220);
nand U7474 (N_7474,N_7213,N_7351);
and U7475 (N_7475,N_7319,N_7341);
or U7476 (N_7476,N_7369,N_7271);
nor U7477 (N_7477,N_7231,N_7218);
and U7478 (N_7478,N_7364,N_7304);
nor U7479 (N_7479,N_7206,N_7236);
nand U7480 (N_7480,N_7307,N_7240);
or U7481 (N_7481,N_7382,N_7361);
xnor U7482 (N_7482,N_7349,N_7235);
xor U7483 (N_7483,N_7227,N_7380);
and U7484 (N_7484,N_7399,N_7340);
nand U7485 (N_7485,N_7281,N_7360);
xnor U7486 (N_7486,N_7376,N_7278);
and U7487 (N_7487,N_7211,N_7250);
nand U7488 (N_7488,N_7330,N_7331);
and U7489 (N_7489,N_7344,N_7383);
nor U7490 (N_7490,N_7239,N_7366);
or U7491 (N_7491,N_7313,N_7293);
xnor U7492 (N_7492,N_7292,N_7234);
and U7493 (N_7493,N_7247,N_7266);
xor U7494 (N_7494,N_7311,N_7275);
and U7495 (N_7495,N_7286,N_7288);
and U7496 (N_7496,N_7395,N_7299);
or U7497 (N_7497,N_7294,N_7339);
nor U7498 (N_7498,N_7209,N_7238);
xor U7499 (N_7499,N_7212,N_7377);
nand U7500 (N_7500,N_7298,N_7201);
xnor U7501 (N_7501,N_7293,N_7344);
nand U7502 (N_7502,N_7391,N_7300);
nand U7503 (N_7503,N_7327,N_7211);
or U7504 (N_7504,N_7284,N_7201);
or U7505 (N_7505,N_7336,N_7385);
or U7506 (N_7506,N_7306,N_7262);
nand U7507 (N_7507,N_7270,N_7364);
nor U7508 (N_7508,N_7212,N_7242);
xnor U7509 (N_7509,N_7318,N_7216);
xnor U7510 (N_7510,N_7212,N_7395);
nor U7511 (N_7511,N_7389,N_7261);
xnor U7512 (N_7512,N_7374,N_7301);
or U7513 (N_7513,N_7213,N_7364);
xnor U7514 (N_7514,N_7237,N_7318);
nand U7515 (N_7515,N_7228,N_7279);
nor U7516 (N_7516,N_7382,N_7328);
nor U7517 (N_7517,N_7364,N_7293);
nand U7518 (N_7518,N_7216,N_7238);
nand U7519 (N_7519,N_7260,N_7381);
nor U7520 (N_7520,N_7244,N_7283);
xnor U7521 (N_7521,N_7257,N_7208);
nor U7522 (N_7522,N_7205,N_7293);
xor U7523 (N_7523,N_7398,N_7328);
and U7524 (N_7524,N_7328,N_7358);
and U7525 (N_7525,N_7274,N_7372);
nand U7526 (N_7526,N_7341,N_7396);
or U7527 (N_7527,N_7263,N_7217);
nor U7528 (N_7528,N_7336,N_7299);
xor U7529 (N_7529,N_7258,N_7366);
nand U7530 (N_7530,N_7358,N_7246);
and U7531 (N_7531,N_7224,N_7327);
nor U7532 (N_7532,N_7304,N_7357);
xor U7533 (N_7533,N_7329,N_7304);
or U7534 (N_7534,N_7244,N_7200);
nor U7535 (N_7535,N_7338,N_7225);
and U7536 (N_7536,N_7243,N_7386);
nand U7537 (N_7537,N_7296,N_7362);
or U7538 (N_7538,N_7259,N_7360);
and U7539 (N_7539,N_7326,N_7276);
or U7540 (N_7540,N_7201,N_7347);
xnor U7541 (N_7541,N_7261,N_7246);
nor U7542 (N_7542,N_7276,N_7308);
nand U7543 (N_7543,N_7304,N_7355);
nor U7544 (N_7544,N_7233,N_7393);
and U7545 (N_7545,N_7287,N_7271);
or U7546 (N_7546,N_7231,N_7249);
or U7547 (N_7547,N_7220,N_7334);
nor U7548 (N_7548,N_7340,N_7349);
nor U7549 (N_7549,N_7343,N_7248);
nor U7550 (N_7550,N_7296,N_7377);
or U7551 (N_7551,N_7223,N_7330);
or U7552 (N_7552,N_7383,N_7380);
xnor U7553 (N_7553,N_7215,N_7239);
nor U7554 (N_7554,N_7391,N_7367);
nor U7555 (N_7555,N_7300,N_7313);
or U7556 (N_7556,N_7266,N_7212);
or U7557 (N_7557,N_7207,N_7394);
nor U7558 (N_7558,N_7211,N_7337);
xor U7559 (N_7559,N_7317,N_7245);
nand U7560 (N_7560,N_7223,N_7314);
nand U7561 (N_7561,N_7268,N_7221);
and U7562 (N_7562,N_7240,N_7312);
and U7563 (N_7563,N_7387,N_7388);
xnor U7564 (N_7564,N_7335,N_7234);
or U7565 (N_7565,N_7206,N_7268);
nand U7566 (N_7566,N_7336,N_7276);
xor U7567 (N_7567,N_7378,N_7248);
and U7568 (N_7568,N_7271,N_7251);
xor U7569 (N_7569,N_7318,N_7397);
or U7570 (N_7570,N_7327,N_7390);
and U7571 (N_7571,N_7275,N_7372);
and U7572 (N_7572,N_7357,N_7364);
nand U7573 (N_7573,N_7377,N_7322);
xor U7574 (N_7574,N_7319,N_7388);
or U7575 (N_7575,N_7291,N_7372);
nand U7576 (N_7576,N_7275,N_7230);
and U7577 (N_7577,N_7244,N_7237);
xor U7578 (N_7578,N_7358,N_7210);
nor U7579 (N_7579,N_7320,N_7309);
and U7580 (N_7580,N_7237,N_7272);
nor U7581 (N_7581,N_7233,N_7365);
nor U7582 (N_7582,N_7315,N_7331);
nand U7583 (N_7583,N_7280,N_7251);
and U7584 (N_7584,N_7323,N_7215);
xor U7585 (N_7585,N_7373,N_7246);
and U7586 (N_7586,N_7311,N_7305);
or U7587 (N_7587,N_7246,N_7337);
nand U7588 (N_7588,N_7290,N_7360);
or U7589 (N_7589,N_7303,N_7211);
xnor U7590 (N_7590,N_7203,N_7392);
or U7591 (N_7591,N_7363,N_7372);
nor U7592 (N_7592,N_7382,N_7315);
xor U7593 (N_7593,N_7355,N_7283);
and U7594 (N_7594,N_7342,N_7241);
or U7595 (N_7595,N_7290,N_7285);
nand U7596 (N_7596,N_7384,N_7276);
nand U7597 (N_7597,N_7245,N_7283);
nand U7598 (N_7598,N_7329,N_7222);
nand U7599 (N_7599,N_7297,N_7282);
and U7600 (N_7600,N_7468,N_7530);
xnor U7601 (N_7601,N_7418,N_7598);
or U7602 (N_7602,N_7557,N_7507);
xnor U7603 (N_7603,N_7432,N_7475);
and U7604 (N_7604,N_7479,N_7473);
nor U7605 (N_7605,N_7596,N_7455);
xnor U7606 (N_7606,N_7477,N_7595);
xor U7607 (N_7607,N_7489,N_7599);
xor U7608 (N_7608,N_7581,N_7487);
and U7609 (N_7609,N_7533,N_7420);
xnor U7610 (N_7610,N_7532,N_7521);
nor U7611 (N_7611,N_7560,N_7571);
nor U7612 (N_7612,N_7400,N_7409);
nor U7613 (N_7613,N_7508,N_7478);
or U7614 (N_7614,N_7590,N_7461);
and U7615 (N_7615,N_7594,N_7421);
nand U7616 (N_7616,N_7417,N_7405);
xnor U7617 (N_7617,N_7579,N_7584);
nor U7618 (N_7618,N_7585,N_7469);
nand U7619 (N_7619,N_7516,N_7467);
nor U7620 (N_7620,N_7518,N_7591);
and U7621 (N_7621,N_7460,N_7506);
nand U7622 (N_7622,N_7412,N_7535);
and U7623 (N_7623,N_7422,N_7553);
or U7624 (N_7624,N_7534,N_7483);
and U7625 (N_7625,N_7463,N_7407);
nor U7626 (N_7626,N_7472,N_7424);
xnor U7627 (N_7627,N_7522,N_7428);
or U7628 (N_7628,N_7569,N_7576);
nand U7629 (N_7629,N_7561,N_7451);
and U7630 (N_7630,N_7491,N_7416);
nor U7631 (N_7631,N_7514,N_7520);
or U7632 (N_7632,N_7493,N_7558);
nand U7633 (N_7633,N_7525,N_7565);
and U7634 (N_7634,N_7515,N_7583);
nand U7635 (N_7635,N_7582,N_7457);
or U7636 (N_7636,N_7509,N_7524);
or U7637 (N_7637,N_7410,N_7430);
nor U7638 (N_7638,N_7448,N_7470);
xor U7639 (N_7639,N_7554,N_7438);
or U7640 (N_7640,N_7434,N_7513);
xor U7641 (N_7641,N_7486,N_7465);
nor U7642 (N_7642,N_7503,N_7415);
nor U7643 (N_7643,N_7556,N_7593);
and U7644 (N_7644,N_7541,N_7481);
nand U7645 (N_7645,N_7484,N_7462);
xnor U7646 (N_7646,N_7511,N_7456);
and U7647 (N_7647,N_7549,N_7490);
and U7648 (N_7648,N_7439,N_7435);
or U7649 (N_7649,N_7458,N_7589);
xnor U7650 (N_7650,N_7464,N_7552);
or U7651 (N_7651,N_7537,N_7496);
or U7652 (N_7652,N_7406,N_7423);
nor U7653 (N_7653,N_7504,N_7586);
nand U7654 (N_7654,N_7447,N_7414);
or U7655 (N_7655,N_7495,N_7544);
nor U7656 (N_7656,N_7476,N_7551);
and U7657 (N_7657,N_7403,N_7572);
nor U7658 (N_7658,N_7546,N_7574);
xor U7659 (N_7659,N_7443,N_7426);
nand U7660 (N_7660,N_7563,N_7531);
or U7661 (N_7661,N_7411,N_7452);
nor U7662 (N_7662,N_7597,N_7440);
xnor U7663 (N_7663,N_7545,N_7529);
or U7664 (N_7664,N_7431,N_7459);
nand U7665 (N_7665,N_7575,N_7485);
or U7666 (N_7666,N_7425,N_7570);
or U7667 (N_7667,N_7567,N_7527);
or U7668 (N_7668,N_7429,N_7550);
and U7669 (N_7669,N_7528,N_7419);
nand U7670 (N_7670,N_7499,N_7450);
xor U7671 (N_7671,N_7562,N_7488);
or U7672 (N_7672,N_7539,N_7592);
nor U7673 (N_7673,N_7519,N_7444);
xor U7674 (N_7674,N_7404,N_7466);
nand U7675 (N_7675,N_7427,N_7454);
nor U7676 (N_7676,N_7433,N_7587);
nand U7677 (N_7677,N_7523,N_7442);
xor U7678 (N_7678,N_7517,N_7577);
xnor U7679 (N_7679,N_7474,N_7580);
and U7680 (N_7680,N_7555,N_7494);
nand U7681 (N_7681,N_7441,N_7480);
nand U7682 (N_7682,N_7498,N_7437);
and U7683 (N_7683,N_7413,N_7548);
xor U7684 (N_7684,N_7471,N_7501);
and U7685 (N_7685,N_7449,N_7497);
xnor U7686 (N_7686,N_7401,N_7538);
nand U7687 (N_7687,N_7502,N_7436);
and U7688 (N_7688,N_7453,N_7500);
xnor U7689 (N_7689,N_7578,N_7492);
or U7690 (N_7690,N_7536,N_7566);
or U7691 (N_7691,N_7408,N_7445);
or U7692 (N_7692,N_7564,N_7542);
and U7693 (N_7693,N_7568,N_7402);
and U7694 (N_7694,N_7510,N_7482);
nor U7695 (N_7695,N_7559,N_7543);
or U7696 (N_7696,N_7588,N_7446);
xnor U7697 (N_7697,N_7526,N_7547);
nor U7698 (N_7698,N_7573,N_7540);
nand U7699 (N_7699,N_7512,N_7505);
nand U7700 (N_7700,N_7588,N_7533);
xor U7701 (N_7701,N_7492,N_7541);
xnor U7702 (N_7702,N_7414,N_7546);
or U7703 (N_7703,N_7502,N_7535);
or U7704 (N_7704,N_7517,N_7401);
xor U7705 (N_7705,N_7526,N_7472);
nand U7706 (N_7706,N_7489,N_7457);
nor U7707 (N_7707,N_7508,N_7506);
nor U7708 (N_7708,N_7583,N_7523);
xor U7709 (N_7709,N_7482,N_7447);
nor U7710 (N_7710,N_7575,N_7497);
nor U7711 (N_7711,N_7435,N_7466);
nor U7712 (N_7712,N_7485,N_7403);
xor U7713 (N_7713,N_7425,N_7596);
or U7714 (N_7714,N_7423,N_7475);
and U7715 (N_7715,N_7583,N_7567);
or U7716 (N_7716,N_7449,N_7499);
nand U7717 (N_7717,N_7409,N_7560);
nor U7718 (N_7718,N_7451,N_7482);
xor U7719 (N_7719,N_7599,N_7426);
nand U7720 (N_7720,N_7405,N_7571);
xnor U7721 (N_7721,N_7417,N_7519);
xnor U7722 (N_7722,N_7418,N_7462);
nand U7723 (N_7723,N_7456,N_7598);
nor U7724 (N_7724,N_7411,N_7485);
xor U7725 (N_7725,N_7442,N_7526);
or U7726 (N_7726,N_7515,N_7521);
or U7727 (N_7727,N_7521,N_7480);
nand U7728 (N_7728,N_7554,N_7471);
nor U7729 (N_7729,N_7574,N_7582);
nor U7730 (N_7730,N_7433,N_7575);
nor U7731 (N_7731,N_7458,N_7420);
nor U7732 (N_7732,N_7446,N_7480);
and U7733 (N_7733,N_7460,N_7425);
nor U7734 (N_7734,N_7536,N_7429);
nor U7735 (N_7735,N_7476,N_7502);
xor U7736 (N_7736,N_7444,N_7574);
or U7737 (N_7737,N_7574,N_7450);
nand U7738 (N_7738,N_7445,N_7480);
nor U7739 (N_7739,N_7529,N_7594);
and U7740 (N_7740,N_7410,N_7526);
or U7741 (N_7741,N_7542,N_7510);
nor U7742 (N_7742,N_7422,N_7487);
and U7743 (N_7743,N_7404,N_7591);
nor U7744 (N_7744,N_7471,N_7411);
and U7745 (N_7745,N_7553,N_7588);
nor U7746 (N_7746,N_7405,N_7539);
and U7747 (N_7747,N_7476,N_7477);
xor U7748 (N_7748,N_7451,N_7501);
nand U7749 (N_7749,N_7508,N_7420);
and U7750 (N_7750,N_7419,N_7425);
and U7751 (N_7751,N_7565,N_7491);
nand U7752 (N_7752,N_7435,N_7418);
nor U7753 (N_7753,N_7562,N_7507);
nor U7754 (N_7754,N_7575,N_7531);
nor U7755 (N_7755,N_7447,N_7411);
nand U7756 (N_7756,N_7471,N_7558);
or U7757 (N_7757,N_7576,N_7571);
nand U7758 (N_7758,N_7519,N_7433);
nand U7759 (N_7759,N_7530,N_7447);
xor U7760 (N_7760,N_7540,N_7448);
or U7761 (N_7761,N_7511,N_7439);
nand U7762 (N_7762,N_7570,N_7432);
and U7763 (N_7763,N_7525,N_7555);
xnor U7764 (N_7764,N_7435,N_7588);
nand U7765 (N_7765,N_7442,N_7513);
nor U7766 (N_7766,N_7476,N_7509);
xnor U7767 (N_7767,N_7437,N_7453);
nand U7768 (N_7768,N_7455,N_7506);
nor U7769 (N_7769,N_7477,N_7586);
nor U7770 (N_7770,N_7472,N_7488);
nand U7771 (N_7771,N_7582,N_7558);
and U7772 (N_7772,N_7552,N_7590);
nand U7773 (N_7773,N_7502,N_7403);
nand U7774 (N_7774,N_7567,N_7475);
xnor U7775 (N_7775,N_7522,N_7473);
nor U7776 (N_7776,N_7413,N_7581);
nor U7777 (N_7777,N_7582,N_7437);
xnor U7778 (N_7778,N_7555,N_7476);
nand U7779 (N_7779,N_7451,N_7591);
and U7780 (N_7780,N_7408,N_7457);
xnor U7781 (N_7781,N_7533,N_7563);
and U7782 (N_7782,N_7581,N_7422);
or U7783 (N_7783,N_7498,N_7497);
nand U7784 (N_7784,N_7427,N_7521);
nor U7785 (N_7785,N_7575,N_7411);
nand U7786 (N_7786,N_7474,N_7560);
nand U7787 (N_7787,N_7577,N_7500);
xor U7788 (N_7788,N_7577,N_7455);
and U7789 (N_7789,N_7471,N_7567);
nor U7790 (N_7790,N_7592,N_7503);
xor U7791 (N_7791,N_7496,N_7556);
or U7792 (N_7792,N_7495,N_7589);
nand U7793 (N_7793,N_7504,N_7484);
or U7794 (N_7794,N_7594,N_7430);
nand U7795 (N_7795,N_7488,N_7461);
and U7796 (N_7796,N_7418,N_7471);
or U7797 (N_7797,N_7511,N_7545);
nand U7798 (N_7798,N_7514,N_7412);
nor U7799 (N_7799,N_7588,N_7493);
and U7800 (N_7800,N_7786,N_7748);
or U7801 (N_7801,N_7626,N_7675);
xnor U7802 (N_7802,N_7751,N_7799);
nand U7803 (N_7803,N_7616,N_7636);
nand U7804 (N_7804,N_7776,N_7721);
or U7805 (N_7805,N_7634,N_7619);
nand U7806 (N_7806,N_7775,N_7651);
nor U7807 (N_7807,N_7796,N_7701);
nor U7808 (N_7808,N_7793,N_7627);
or U7809 (N_7809,N_7784,N_7767);
nand U7810 (N_7810,N_7709,N_7690);
and U7811 (N_7811,N_7719,N_7705);
or U7812 (N_7812,N_7630,N_7696);
nand U7813 (N_7813,N_7687,N_7669);
or U7814 (N_7814,N_7743,N_7672);
nand U7815 (N_7815,N_7695,N_7694);
and U7816 (N_7816,N_7649,N_7684);
and U7817 (N_7817,N_7632,N_7720);
and U7818 (N_7818,N_7702,N_7657);
and U7819 (N_7819,N_7740,N_7755);
and U7820 (N_7820,N_7679,N_7662);
xor U7821 (N_7821,N_7797,N_7635);
and U7822 (N_7822,N_7756,N_7710);
xnor U7823 (N_7823,N_7673,N_7678);
xor U7824 (N_7824,N_7728,N_7700);
or U7825 (N_7825,N_7724,N_7771);
or U7826 (N_7826,N_7715,N_7692);
or U7827 (N_7827,N_7752,N_7666);
and U7828 (N_7828,N_7622,N_7762);
and U7829 (N_7829,N_7647,N_7613);
xor U7830 (N_7830,N_7749,N_7688);
nor U7831 (N_7831,N_7708,N_7711);
nand U7832 (N_7832,N_7660,N_7792);
nand U7833 (N_7833,N_7686,N_7631);
nor U7834 (N_7834,N_7791,N_7620);
xnor U7835 (N_7835,N_7712,N_7645);
nor U7836 (N_7836,N_7727,N_7766);
nor U7837 (N_7837,N_7779,N_7656);
nand U7838 (N_7838,N_7644,N_7606);
nor U7839 (N_7839,N_7670,N_7639);
nand U7840 (N_7840,N_7787,N_7729);
nor U7841 (N_7841,N_7614,N_7783);
nor U7842 (N_7842,N_7621,N_7768);
nor U7843 (N_7843,N_7680,N_7650);
and U7844 (N_7844,N_7612,N_7716);
or U7845 (N_7845,N_7753,N_7658);
nor U7846 (N_7846,N_7667,N_7661);
nand U7847 (N_7847,N_7785,N_7625);
nand U7848 (N_7848,N_7600,N_7698);
xnor U7849 (N_7849,N_7782,N_7604);
or U7850 (N_7850,N_7742,N_7774);
nand U7851 (N_7851,N_7747,N_7788);
xnor U7852 (N_7852,N_7739,N_7664);
nand U7853 (N_7853,N_7717,N_7769);
or U7854 (N_7854,N_7737,N_7736);
and U7855 (N_7855,N_7611,N_7772);
or U7856 (N_7856,N_7781,N_7759);
or U7857 (N_7857,N_7780,N_7628);
or U7858 (N_7858,N_7629,N_7726);
nand U7859 (N_7859,N_7677,N_7730);
nor U7860 (N_7860,N_7643,N_7641);
nor U7861 (N_7861,N_7750,N_7757);
or U7862 (N_7862,N_7741,N_7633);
nor U7863 (N_7863,N_7608,N_7795);
and U7864 (N_7864,N_7682,N_7734);
or U7865 (N_7865,N_7723,N_7655);
nand U7866 (N_7866,N_7623,N_7699);
and U7867 (N_7867,N_7703,N_7754);
nand U7868 (N_7868,N_7689,N_7648);
and U7869 (N_7869,N_7763,N_7764);
and U7870 (N_7870,N_7615,N_7731);
or U7871 (N_7871,N_7618,N_7642);
xnor U7872 (N_7872,N_7637,N_7610);
and U7873 (N_7873,N_7638,N_7609);
nand U7874 (N_7874,N_7773,N_7760);
xor U7875 (N_7875,N_7691,N_7659);
xor U7876 (N_7876,N_7607,N_7778);
nand U7877 (N_7877,N_7707,N_7697);
and U7878 (N_7878,N_7665,N_7676);
nor U7879 (N_7879,N_7765,N_7777);
or U7880 (N_7880,N_7722,N_7761);
nand U7881 (N_7881,N_7770,N_7738);
nand U7882 (N_7882,N_7733,N_7790);
nand U7883 (N_7883,N_7735,N_7758);
nor U7884 (N_7884,N_7746,N_7714);
nor U7885 (N_7885,N_7798,N_7794);
xor U7886 (N_7886,N_7646,N_7671);
nand U7887 (N_7887,N_7617,N_7789);
nand U7888 (N_7888,N_7725,N_7654);
or U7889 (N_7889,N_7624,N_7718);
and U7890 (N_7890,N_7683,N_7653);
nand U7891 (N_7891,N_7681,N_7602);
or U7892 (N_7892,N_7706,N_7605);
and U7893 (N_7893,N_7704,N_7732);
nor U7894 (N_7894,N_7640,N_7603);
nand U7895 (N_7895,N_7652,N_7668);
nor U7896 (N_7896,N_7744,N_7663);
or U7897 (N_7897,N_7745,N_7713);
nand U7898 (N_7898,N_7685,N_7693);
and U7899 (N_7899,N_7674,N_7601);
or U7900 (N_7900,N_7781,N_7705);
xnor U7901 (N_7901,N_7644,N_7641);
or U7902 (N_7902,N_7736,N_7685);
xnor U7903 (N_7903,N_7742,N_7697);
nor U7904 (N_7904,N_7712,N_7615);
xnor U7905 (N_7905,N_7670,N_7705);
nor U7906 (N_7906,N_7677,N_7612);
xor U7907 (N_7907,N_7715,N_7659);
and U7908 (N_7908,N_7748,N_7747);
nor U7909 (N_7909,N_7682,N_7700);
or U7910 (N_7910,N_7655,N_7687);
nand U7911 (N_7911,N_7613,N_7602);
or U7912 (N_7912,N_7701,N_7755);
nor U7913 (N_7913,N_7761,N_7663);
nand U7914 (N_7914,N_7698,N_7777);
and U7915 (N_7915,N_7666,N_7656);
nor U7916 (N_7916,N_7737,N_7769);
and U7917 (N_7917,N_7734,N_7767);
nor U7918 (N_7918,N_7726,N_7776);
or U7919 (N_7919,N_7762,N_7612);
nand U7920 (N_7920,N_7670,N_7653);
and U7921 (N_7921,N_7622,N_7692);
nor U7922 (N_7922,N_7796,N_7666);
nor U7923 (N_7923,N_7673,N_7616);
nand U7924 (N_7924,N_7715,N_7773);
nand U7925 (N_7925,N_7710,N_7770);
xor U7926 (N_7926,N_7774,N_7702);
nand U7927 (N_7927,N_7705,N_7730);
nand U7928 (N_7928,N_7798,N_7600);
or U7929 (N_7929,N_7766,N_7630);
xnor U7930 (N_7930,N_7754,N_7617);
or U7931 (N_7931,N_7734,N_7760);
nor U7932 (N_7932,N_7642,N_7690);
or U7933 (N_7933,N_7604,N_7763);
xor U7934 (N_7934,N_7751,N_7705);
xor U7935 (N_7935,N_7628,N_7752);
or U7936 (N_7936,N_7764,N_7774);
nand U7937 (N_7937,N_7753,N_7780);
and U7938 (N_7938,N_7763,N_7796);
nand U7939 (N_7939,N_7624,N_7769);
or U7940 (N_7940,N_7600,N_7659);
and U7941 (N_7941,N_7789,N_7790);
or U7942 (N_7942,N_7640,N_7649);
nand U7943 (N_7943,N_7775,N_7614);
or U7944 (N_7944,N_7709,N_7753);
nor U7945 (N_7945,N_7753,N_7712);
nor U7946 (N_7946,N_7631,N_7680);
and U7947 (N_7947,N_7607,N_7691);
xnor U7948 (N_7948,N_7728,N_7605);
or U7949 (N_7949,N_7658,N_7775);
nand U7950 (N_7950,N_7778,N_7773);
and U7951 (N_7951,N_7614,N_7639);
or U7952 (N_7952,N_7611,N_7609);
nand U7953 (N_7953,N_7744,N_7660);
nor U7954 (N_7954,N_7787,N_7777);
nor U7955 (N_7955,N_7668,N_7628);
and U7956 (N_7956,N_7754,N_7603);
and U7957 (N_7957,N_7619,N_7731);
xor U7958 (N_7958,N_7626,N_7601);
and U7959 (N_7959,N_7698,N_7616);
xor U7960 (N_7960,N_7746,N_7772);
xnor U7961 (N_7961,N_7777,N_7739);
and U7962 (N_7962,N_7732,N_7621);
nand U7963 (N_7963,N_7650,N_7653);
xnor U7964 (N_7964,N_7681,N_7655);
and U7965 (N_7965,N_7755,N_7605);
nor U7966 (N_7966,N_7689,N_7674);
nand U7967 (N_7967,N_7748,N_7688);
nand U7968 (N_7968,N_7651,N_7616);
or U7969 (N_7969,N_7648,N_7766);
nor U7970 (N_7970,N_7767,N_7604);
and U7971 (N_7971,N_7614,N_7690);
and U7972 (N_7972,N_7620,N_7762);
nor U7973 (N_7973,N_7770,N_7766);
and U7974 (N_7974,N_7684,N_7664);
nor U7975 (N_7975,N_7655,N_7716);
and U7976 (N_7976,N_7643,N_7637);
xnor U7977 (N_7977,N_7771,N_7749);
or U7978 (N_7978,N_7660,N_7742);
xnor U7979 (N_7979,N_7728,N_7776);
nand U7980 (N_7980,N_7600,N_7636);
and U7981 (N_7981,N_7708,N_7643);
or U7982 (N_7982,N_7623,N_7618);
or U7983 (N_7983,N_7794,N_7626);
and U7984 (N_7984,N_7649,N_7788);
and U7985 (N_7985,N_7645,N_7735);
xor U7986 (N_7986,N_7719,N_7713);
and U7987 (N_7987,N_7695,N_7728);
xnor U7988 (N_7988,N_7629,N_7782);
xnor U7989 (N_7989,N_7725,N_7688);
nand U7990 (N_7990,N_7632,N_7626);
nand U7991 (N_7991,N_7627,N_7632);
nand U7992 (N_7992,N_7669,N_7758);
and U7993 (N_7993,N_7689,N_7739);
nand U7994 (N_7994,N_7741,N_7699);
and U7995 (N_7995,N_7625,N_7670);
xnor U7996 (N_7996,N_7656,N_7693);
xnor U7997 (N_7997,N_7679,N_7666);
nand U7998 (N_7998,N_7764,N_7670);
and U7999 (N_7999,N_7751,N_7732);
or U8000 (N_8000,N_7956,N_7817);
nor U8001 (N_8001,N_7950,N_7862);
or U8002 (N_8002,N_7988,N_7873);
or U8003 (N_8003,N_7847,N_7997);
or U8004 (N_8004,N_7899,N_7803);
and U8005 (N_8005,N_7981,N_7937);
or U8006 (N_8006,N_7841,N_7916);
or U8007 (N_8007,N_7869,N_7824);
xnor U8008 (N_8008,N_7801,N_7819);
nand U8009 (N_8009,N_7829,N_7933);
nor U8010 (N_8010,N_7804,N_7864);
nand U8011 (N_8011,N_7823,N_7892);
nand U8012 (N_8012,N_7963,N_7918);
and U8013 (N_8013,N_7993,N_7964);
and U8014 (N_8014,N_7839,N_7930);
or U8015 (N_8015,N_7860,N_7811);
nand U8016 (N_8016,N_7805,N_7912);
xnor U8017 (N_8017,N_7902,N_7896);
nor U8018 (N_8018,N_7851,N_7877);
xor U8019 (N_8019,N_7812,N_7837);
xnor U8020 (N_8020,N_7833,N_7913);
xor U8021 (N_8021,N_7849,N_7921);
or U8022 (N_8022,N_7931,N_7999);
and U8023 (N_8023,N_7955,N_7818);
nor U8024 (N_8024,N_7935,N_7983);
xnor U8025 (N_8025,N_7848,N_7890);
nand U8026 (N_8026,N_7802,N_7843);
xnor U8027 (N_8027,N_7946,N_7966);
nor U8028 (N_8028,N_7826,N_7904);
nor U8029 (N_8029,N_7910,N_7962);
nand U8030 (N_8030,N_7857,N_7920);
xnor U8031 (N_8031,N_7952,N_7954);
nor U8032 (N_8032,N_7936,N_7868);
nor U8033 (N_8033,N_7980,N_7940);
nor U8034 (N_8034,N_7828,N_7926);
and U8035 (N_8035,N_7925,N_7845);
and U8036 (N_8036,N_7942,N_7907);
nor U8037 (N_8037,N_7941,N_7995);
nand U8038 (N_8038,N_7850,N_7915);
or U8039 (N_8039,N_7827,N_7957);
xor U8040 (N_8040,N_7970,N_7893);
nand U8041 (N_8041,N_7932,N_7987);
and U8042 (N_8042,N_7872,N_7919);
nor U8043 (N_8043,N_7886,N_7986);
xor U8044 (N_8044,N_7853,N_7985);
or U8045 (N_8045,N_7943,N_7881);
or U8046 (N_8046,N_7840,N_7992);
nor U8047 (N_8047,N_7800,N_7882);
and U8048 (N_8048,N_7888,N_7809);
nor U8049 (N_8049,N_7855,N_7908);
nand U8050 (N_8050,N_7852,N_7994);
nor U8051 (N_8051,N_7863,N_7879);
nand U8052 (N_8052,N_7923,N_7889);
and U8053 (N_8053,N_7967,N_7885);
nand U8054 (N_8054,N_7901,N_7815);
and U8055 (N_8055,N_7825,N_7835);
nand U8056 (N_8056,N_7807,N_7858);
xnor U8057 (N_8057,N_7810,N_7979);
nand U8058 (N_8058,N_7866,N_7928);
xnor U8059 (N_8059,N_7822,N_7816);
and U8060 (N_8060,N_7968,N_7914);
xor U8061 (N_8061,N_7973,N_7934);
and U8062 (N_8062,N_7838,N_7834);
or U8063 (N_8063,N_7960,N_7927);
nor U8064 (N_8064,N_7965,N_7938);
xnor U8065 (N_8065,N_7831,N_7990);
xor U8066 (N_8066,N_7876,N_7974);
or U8067 (N_8067,N_7984,N_7909);
xor U8068 (N_8068,N_7903,N_7975);
nand U8069 (N_8069,N_7917,N_7959);
nand U8070 (N_8070,N_7953,N_7898);
nor U8071 (N_8071,N_7976,N_7806);
xor U8072 (N_8072,N_7891,N_7883);
xor U8073 (N_8073,N_7887,N_7948);
and U8074 (N_8074,N_7874,N_7996);
or U8075 (N_8075,N_7989,N_7958);
or U8076 (N_8076,N_7884,N_7836);
xor U8077 (N_8077,N_7871,N_7880);
and U8078 (N_8078,N_7972,N_7870);
and U8079 (N_8079,N_7894,N_7969);
or U8080 (N_8080,N_7897,N_7961);
or U8081 (N_8081,N_7929,N_7875);
or U8082 (N_8082,N_7820,N_7854);
nor U8083 (N_8083,N_7808,N_7878);
nand U8084 (N_8084,N_7944,N_7844);
nor U8085 (N_8085,N_7861,N_7982);
or U8086 (N_8086,N_7832,N_7846);
and U8087 (N_8087,N_7939,N_7865);
nor U8088 (N_8088,N_7949,N_7867);
nand U8089 (N_8089,N_7895,N_7945);
and U8090 (N_8090,N_7971,N_7813);
xnor U8091 (N_8091,N_7906,N_7859);
and U8092 (N_8092,N_7856,N_7922);
and U8093 (N_8093,N_7830,N_7842);
and U8094 (N_8094,N_7900,N_7905);
xor U8095 (N_8095,N_7978,N_7951);
nor U8096 (N_8096,N_7911,N_7821);
or U8097 (N_8097,N_7998,N_7991);
nor U8098 (N_8098,N_7924,N_7947);
or U8099 (N_8099,N_7977,N_7814);
xnor U8100 (N_8100,N_7855,N_7806);
nand U8101 (N_8101,N_7907,N_7933);
or U8102 (N_8102,N_7840,N_7827);
nand U8103 (N_8103,N_7849,N_7834);
nor U8104 (N_8104,N_7902,N_7887);
or U8105 (N_8105,N_7873,N_7950);
nor U8106 (N_8106,N_7915,N_7805);
or U8107 (N_8107,N_7995,N_7872);
nand U8108 (N_8108,N_7979,N_7905);
xor U8109 (N_8109,N_7928,N_7852);
nand U8110 (N_8110,N_7826,N_7940);
xnor U8111 (N_8111,N_7867,N_7847);
nor U8112 (N_8112,N_7906,N_7884);
or U8113 (N_8113,N_7848,N_7828);
nor U8114 (N_8114,N_7924,N_7819);
nor U8115 (N_8115,N_7967,N_7867);
and U8116 (N_8116,N_7935,N_7982);
nand U8117 (N_8117,N_7833,N_7993);
or U8118 (N_8118,N_7906,N_7866);
and U8119 (N_8119,N_7846,N_7930);
xnor U8120 (N_8120,N_7888,N_7812);
or U8121 (N_8121,N_7959,N_7824);
nand U8122 (N_8122,N_7966,N_7917);
nand U8123 (N_8123,N_7991,N_7901);
nand U8124 (N_8124,N_7833,N_7839);
or U8125 (N_8125,N_7810,N_7883);
or U8126 (N_8126,N_7875,N_7823);
xnor U8127 (N_8127,N_7883,N_7863);
xor U8128 (N_8128,N_7916,N_7806);
nand U8129 (N_8129,N_7948,N_7814);
or U8130 (N_8130,N_7981,N_7978);
and U8131 (N_8131,N_7989,N_7831);
xor U8132 (N_8132,N_7953,N_7950);
nor U8133 (N_8133,N_7968,N_7814);
and U8134 (N_8134,N_7891,N_7815);
and U8135 (N_8135,N_7911,N_7921);
and U8136 (N_8136,N_7996,N_7984);
nand U8137 (N_8137,N_7888,N_7821);
nor U8138 (N_8138,N_7927,N_7995);
nand U8139 (N_8139,N_7865,N_7877);
or U8140 (N_8140,N_7982,N_7974);
nor U8141 (N_8141,N_7889,N_7924);
nor U8142 (N_8142,N_7948,N_7904);
or U8143 (N_8143,N_7979,N_7943);
nor U8144 (N_8144,N_7937,N_7934);
xor U8145 (N_8145,N_7895,N_7870);
xnor U8146 (N_8146,N_7801,N_7985);
nand U8147 (N_8147,N_7809,N_7876);
xor U8148 (N_8148,N_7882,N_7837);
and U8149 (N_8149,N_7874,N_7877);
or U8150 (N_8150,N_7819,N_7880);
nand U8151 (N_8151,N_7801,N_7991);
or U8152 (N_8152,N_7994,N_7825);
nor U8153 (N_8153,N_7969,N_7912);
nor U8154 (N_8154,N_7830,N_7963);
xnor U8155 (N_8155,N_7865,N_7937);
xnor U8156 (N_8156,N_7916,N_7885);
or U8157 (N_8157,N_7988,N_7811);
nand U8158 (N_8158,N_7980,N_7997);
or U8159 (N_8159,N_7899,N_7912);
and U8160 (N_8160,N_7873,N_7852);
and U8161 (N_8161,N_7839,N_7953);
and U8162 (N_8162,N_7974,N_7819);
or U8163 (N_8163,N_7818,N_7821);
or U8164 (N_8164,N_7870,N_7852);
or U8165 (N_8165,N_7971,N_7840);
nor U8166 (N_8166,N_7996,N_7951);
nor U8167 (N_8167,N_7960,N_7973);
xnor U8168 (N_8168,N_7833,N_7849);
or U8169 (N_8169,N_7930,N_7960);
nand U8170 (N_8170,N_7847,N_7832);
xor U8171 (N_8171,N_7957,N_7924);
and U8172 (N_8172,N_7947,N_7925);
xnor U8173 (N_8173,N_7900,N_7922);
or U8174 (N_8174,N_7931,N_7854);
nor U8175 (N_8175,N_7996,N_7865);
nor U8176 (N_8176,N_7807,N_7868);
or U8177 (N_8177,N_7917,N_7869);
xor U8178 (N_8178,N_7811,N_7835);
xor U8179 (N_8179,N_7962,N_7804);
nor U8180 (N_8180,N_7858,N_7956);
nor U8181 (N_8181,N_7879,N_7958);
nand U8182 (N_8182,N_7884,N_7997);
xnor U8183 (N_8183,N_7984,N_7828);
xor U8184 (N_8184,N_7928,N_7951);
and U8185 (N_8185,N_7829,N_7942);
nand U8186 (N_8186,N_7955,N_7949);
or U8187 (N_8187,N_7827,N_7986);
nand U8188 (N_8188,N_7835,N_7977);
nor U8189 (N_8189,N_7884,N_7846);
and U8190 (N_8190,N_7915,N_7995);
nor U8191 (N_8191,N_7929,N_7975);
nand U8192 (N_8192,N_7851,N_7917);
nand U8193 (N_8193,N_7973,N_7897);
xor U8194 (N_8194,N_7988,N_7945);
nand U8195 (N_8195,N_7806,N_7814);
or U8196 (N_8196,N_7866,N_7860);
and U8197 (N_8197,N_7889,N_7965);
nor U8198 (N_8198,N_7971,N_7816);
or U8199 (N_8199,N_7870,N_7967);
nand U8200 (N_8200,N_8175,N_8139);
xor U8201 (N_8201,N_8080,N_8008);
and U8202 (N_8202,N_8012,N_8166);
xor U8203 (N_8203,N_8143,N_8018);
xor U8204 (N_8204,N_8160,N_8006);
nand U8205 (N_8205,N_8088,N_8067);
xnor U8206 (N_8206,N_8159,N_8199);
nand U8207 (N_8207,N_8141,N_8074);
nor U8208 (N_8208,N_8157,N_8109);
or U8209 (N_8209,N_8033,N_8148);
xnor U8210 (N_8210,N_8097,N_8104);
xor U8211 (N_8211,N_8077,N_8186);
nor U8212 (N_8212,N_8150,N_8130);
and U8213 (N_8213,N_8021,N_8196);
or U8214 (N_8214,N_8154,N_8071);
xnor U8215 (N_8215,N_8189,N_8123);
nand U8216 (N_8216,N_8176,N_8180);
or U8217 (N_8217,N_8023,N_8016);
nand U8218 (N_8218,N_8087,N_8124);
nand U8219 (N_8219,N_8015,N_8064);
nand U8220 (N_8220,N_8062,N_8173);
or U8221 (N_8221,N_8136,N_8164);
or U8222 (N_8222,N_8032,N_8045);
and U8223 (N_8223,N_8039,N_8085);
or U8224 (N_8224,N_8086,N_8098);
xor U8225 (N_8225,N_8151,N_8028);
nand U8226 (N_8226,N_8065,N_8115);
nand U8227 (N_8227,N_8082,N_8131);
xnor U8228 (N_8228,N_8184,N_8044);
xor U8229 (N_8229,N_8041,N_8034);
nor U8230 (N_8230,N_8003,N_8043);
nand U8231 (N_8231,N_8185,N_8038);
nand U8232 (N_8232,N_8122,N_8084);
nor U8233 (N_8233,N_8101,N_8168);
xnor U8234 (N_8234,N_8155,N_8000);
xor U8235 (N_8235,N_8153,N_8096);
and U8236 (N_8236,N_8025,N_8052);
nor U8237 (N_8237,N_8026,N_8050);
and U8238 (N_8238,N_8187,N_8127);
nor U8239 (N_8239,N_8194,N_8110);
xor U8240 (N_8240,N_8061,N_8040);
xor U8241 (N_8241,N_8126,N_8027);
nor U8242 (N_8242,N_8002,N_8056);
xor U8243 (N_8243,N_8068,N_8142);
xor U8244 (N_8244,N_8152,N_8001);
or U8245 (N_8245,N_8073,N_8135);
or U8246 (N_8246,N_8197,N_8113);
nor U8247 (N_8247,N_8193,N_8182);
xor U8248 (N_8248,N_8125,N_8019);
or U8249 (N_8249,N_8095,N_8158);
or U8250 (N_8250,N_8069,N_8047);
and U8251 (N_8251,N_8066,N_8192);
or U8252 (N_8252,N_8133,N_8112);
nor U8253 (N_8253,N_8170,N_8024);
nand U8254 (N_8254,N_8013,N_8055);
nor U8255 (N_8255,N_8083,N_8051);
and U8256 (N_8256,N_8099,N_8029);
or U8257 (N_8257,N_8020,N_8114);
nor U8258 (N_8258,N_8090,N_8165);
or U8259 (N_8259,N_8145,N_8011);
or U8260 (N_8260,N_8146,N_8030);
nand U8261 (N_8261,N_8037,N_8121);
nor U8262 (N_8262,N_8177,N_8134);
nand U8263 (N_8263,N_8035,N_8005);
and U8264 (N_8264,N_8076,N_8053);
nor U8265 (N_8265,N_8129,N_8102);
and U8266 (N_8266,N_8179,N_8118);
nor U8267 (N_8267,N_8119,N_8132);
and U8268 (N_8268,N_8105,N_8078);
and U8269 (N_8269,N_8036,N_8181);
xnor U8270 (N_8270,N_8171,N_8190);
nand U8271 (N_8271,N_8106,N_8049);
nor U8272 (N_8272,N_8111,N_8169);
and U8273 (N_8273,N_8017,N_8014);
nand U8274 (N_8274,N_8009,N_8167);
and U8275 (N_8275,N_8163,N_8094);
and U8276 (N_8276,N_8178,N_8091);
and U8277 (N_8277,N_8031,N_8162);
nand U8278 (N_8278,N_8188,N_8103);
nand U8279 (N_8279,N_8198,N_8144);
and U8280 (N_8280,N_8054,N_8075);
and U8281 (N_8281,N_8108,N_8195);
xor U8282 (N_8282,N_8089,N_8057);
and U8283 (N_8283,N_8058,N_8147);
nor U8284 (N_8284,N_8174,N_8070);
nor U8285 (N_8285,N_8128,N_8063);
and U8286 (N_8286,N_8100,N_8092);
nand U8287 (N_8287,N_8116,N_8117);
or U8288 (N_8288,N_8059,N_8149);
xor U8289 (N_8289,N_8191,N_8010);
nor U8290 (N_8290,N_8156,N_8183);
or U8291 (N_8291,N_8093,N_8022);
nand U8292 (N_8292,N_8079,N_8161);
and U8293 (N_8293,N_8137,N_8138);
nand U8294 (N_8294,N_8042,N_8120);
nand U8295 (N_8295,N_8007,N_8140);
xnor U8296 (N_8296,N_8081,N_8046);
nor U8297 (N_8297,N_8172,N_8060);
xnor U8298 (N_8298,N_8072,N_8048);
nand U8299 (N_8299,N_8107,N_8004);
nor U8300 (N_8300,N_8172,N_8138);
nor U8301 (N_8301,N_8006,N_8054);
xor U8302 (N_8302,N_8171,N_8115);
xnor U8303 (N_8303,N_8141,N_8059);
or U8304 (N_8304,N_8190,N_8037);
xor U8305 (N_8305,N_8164,N_8003);
xor U8306 (N_8306,N_8017,N_8190);
and U8307 (N_8307,N_8093,N_8028);
nor U8308 (N_8308,N_8135,N_8136);
and U8309 (N_8309,N_8135,N_8096);
and U8310 (N_8310,N_8010,N_8085);
and U8311 (N_8311,N_8180,N_8142);
nand U8312 (N_8312,N_8173,N_8157);
nand U8313 (N_8313,N_8012,N_8111);
xnor U8314 (N_8314,N_8083,N_8064);
and U8315 (N_8315,N_8184,N_8137);
and U8316 (N_8316,N_8062,N_8154);
and U8317 (N_8317,N_8086,N_8139);
and U8318 (N_8318,N_8067,N_8185);
nor U8319 (N_8319,N_8142,N_8191);
xor U8320 (N_8320,N_8044,N_8010);
and U8321 (N_8321,N_8118,N_8057);
nor U8322 (N_8322,N_8152,N_8182);
nand U8323 (N_8323,N_8125,N_8177);
and U8324 (N_8324,N_8124,N_8194);
and U8325 (N_8325,N_8082,N_8092);
xor U8326 (N_8326,N_8176,N_8117);
xnor U8327 (N_8327,N_8073,N_8150);
nor U8328 (N_8328,N_8035,N_8120);
xor U8329 (N_8329,N_8147,N_8080);
nand U8330 (N_8330,N_8088,N_8144);
xnor U8331 (N_8331,N_8043,N_8153);
xnor U8332 (N_8332,N_8106,N_8189);
and U8333 (N_8333,N_8032,N_8132);
or U8334 (N_8334,N_8013,N_8006);
xor U8335 (N_8335,N_8189,N_8099);
nand U8336 (N_8336,N_8046,N_8166);
nand U8337 (N_8337,N_8164,N_8138);
xnor U8338 (N_8338,N_8148,N_8084);
xnor U8339 (N_8339,N_8040,N_8073);
nand U8340 (N_8340,N_8143,N_8129);
and U8341 (N_8341,N_8041,N_8195);
xor U8342 (N_8342,N_8194,N_8094);
xor U8343 (N_8343,N_8079,N_8095);
or U8344 (N_8344,N_8032,N_8107);
or U8345 (N_8345,N_8178,N_8135);
or U8346 (N_8346,N_8114,N_8057);
and U8347 (N_8347,N_8137,N_8191);
nor U8348 (N_8348,N_8080,N_8023);
xor U8349 (N_8349,N_8094,N_8173);
nand U8350 (N_8350,N_8093,N_8133);
or U8351 (N_8351,N_8129,N_8194);
or U8352 (N_8352,N_8015,N_8166);
xnor U8353 (N_8353,N_8187,N_8065);
xnor U8354 (N_8354,N_8115,N_8121);
and U8355 (N_8355,N_8173,N_8067);
or U8356 (N_8356,N_8023,N_8175);
nor U8357 (N_8357,N_8163,N_8196);
xnor U8358 (N_8358,N_8122,N_8004);
nor U8359 (N_8359,N_8097,N_8163);
or U8360 (N_8360,N_8164,N_8044);
or U8361 (N_8361,N_8007,N_8148);
xnor U8362 (N_8362,N_8008,N_8159);
or U8363 (N_8363,N_8083,N_8025);
nand U8364 (N_8364,N_8011,N_8128);
nor U8365 (N_8365,N_8114,N_8014);
and U8366 (N_8366,N_8009,N_8056);
nand U8367 (N_8367,N_8036,N_8078);
xnor U8368 (N_8368,N_8035,N_8066);
nand U8369 (N_8369,N_8091,N_8123);
and U8370 (N_8370,N_8098,N_8124);
xnor U8371 (N_8371,N_8145,N_8177);
nor U8372 (N_8372,N_8171,N_8083);
or U8373 (N_8373,N_8082,N_8079);
nor U8374 (N_8374,N_8035,N_8086);
and U8375 (N_8375,N_8006,N_8031);
and U8376 (N_8376,N_8051,N_8008);
nand U8377 (N_8377,N_8135,N_8092);
nor U8378 (N_8378,N_8094,N_8098);
nor U8379 (N_8379,N_8168,N_8164);
nor U8380 (N_8380,N_8182,N_8058);
nand U8381 (N_8381,N_8154,N_8078);
xor U8382 (N_8382,N_8179,N_8056);
and U8383 (N_8383,N_8048,N_8111);
nor U8384 (N_8384,N_8148,N_8145);
or U8385 (N_8385,N_8045,N_8150);
and U8386 (N_8386,N_8080,N_8102);
nand U8387 (N_8387,N_8047,N_8074);
and U8388 (N_8388,N_8195,N_8081);
nor U8389 (N_8389,N_8090,N_8065);
nor U8390 (N_8390,N_8152,N_8100);
nor U8391 (N_8391,N_8106,N_8146);
nand U8392 (N_8392,N_8033,N_8185);
or U8393 (N_8393,N_8132,N_8190);
nand U8394 (N_8394,N_8162,N_8158);
and U8395 (N_8395,N_8023,N_8125);
xnor U8396 (N_8396,N_8164,N_8052);
and U8397 (N_8397,N_8105,N_8092);
or U8398 (N_8398,N_8036,N_8169);
nor U8399 (N_8399,N_8038,N_8068);
nand U8400 (N_8400,N_8387,N_8361);
or U8401 (N_8401,N_8376,N_8274);
nor U8402 (N_8402,N_8377,N_8260);
xnor U8403 (N_8403,N_8251,N_8305);
and U8404 (N_8404,N_8389,N_8399);
nand U8405 (N_8405,N_8241,N_8285);
nand U8406 (N_8406,N_8353,N_8335);
and U8407 (N_8407,N_8224,N_8299);
and U8408 (N_8408,N_8238,N_8282);
nand U8409 (N_8409,N_8379,N_8232);
nand U8410 (N_8410,N_8268,N_8243);
nor U8411 (N_8411,N_8388,N_8356);
nor U8412 (N_8412,N_8225,N_8203);
xor U8413 (N_8413,N_8247,N_8393);
nor U8414 (N_8414,N_8206,N_8242);
and U8415 (N_8415,N_8372,N_8200);
nand U8416 (N_8416,N_8339,N_8217);
nand U8417 (N_8417,N_8332,N_8294);
nand U8418 (N_8418,N_8363,N_8236);
xor U8419 (N_8419,N_8213,N_8337);
or U8420 (N_8420,N_8325,N_8338);
nand U8421 (N_8421,N_8216,N_8343);
nand U8422 (N_8422,N_8221,N_8229);
or U8423 (N_8423,N_8380,N_8306);
or U8424 (N_8424,N_8227,N_8248);
or U8425 (N_8425,N_8258,N_8261);
xnor U8426 (N_8426,N_8344,N_8239);
or U8427 (N_8427,N_8250,N_8202);
nand U8428 (N_8428,N_8280,N_8381);
or U8429 (N_8429,N_8215,N_8375);
nand U8430 (N_8430,N_8291,N_8340);
or U8431 (N_8431,N_8271,N_8228);
and U8432 (N_8432,N_8336,N_8312);
nor U8433 (N_8433,N_8275,N_8330);
nor U8434 (N_8434,N_8214,N_8277);
and U8435 (N_8435,N_8212,N_8326);
xnor U8436 (N_8436,N_8257,N_8392);
nand U8437 (N_8437,N_8226,N_8378);
and U8438 (N_8438,N_8234,N_8310);
xor U8439 (N_8439,N_8374,N_8347);
nor U8440 (N_8440,N_8255,N_8290);
or U8441 (N_8441,N_8231,N_8266);
nand U8442 (N_8442,N_8262,N_8289);
or U8443 (N_8443,N_8360,N_8279);
or U8444 (N_8444,N_8373,N_8395);
or U8445 (N_8445,N_8253,N_8256);
and U8446 (N_8446,N_8342,N_8295);
or U8447 (N_8447,N_8288,N_8309);
nand U8448 (N_8448,N_8396,N_8328);
xor U8449 (N_8449,N_8303,N_8259);
or U8450 (N_8450,N_8201,N_8394);
nor U8451 (N_8451,N_8313,N_8320);
and U8452 (N_8452,N_8252,N_8298);
or U8453 (N_8453,N_8246,N_8317);
or U8454 (N_8454,N_8207,N_8324);
or U8455 (N_8455,N_8235,N_8254);
or U8456 (N_8456,N_8245,N_8286);
nand U8457 (N_8457,N_8244,N_8319);
and U8458 (N_8458,N_8367,N_8210);
nor U8459 (N_8459,N_8351,N_8348);
xnor U8460 (N_8460,N_8314,N_8265);
or U8461 (N_8461,N_8223,N_8352);
nor U8462 (N_8462,N_8267,N_8263);
and U8463 (N_8463,N_8384,N_8222);
nand U8464 (N_8464,N_8269,N_8321);
and U8465 (N_8465,N_8331,N_8370);
nand U8466 (N_8466,N_8365,N_8398);
nor U8467 (N_8467,N_8390,N_8362);
and U8468 (N_8468,N_8296,N_8386);
and U8469 (N_8469,N_8345,N_8327);
nand U8470 (N_8470,N_8209,N_8264);
nand U8471 (N_8471,N_8211,N_8284);
nand U8472 (N_8472,N_8341,N_8368);
or U8473 (N_8473,N_8297,N_8300);
and U8474 (N_8474,N_8391,N_8204);
nand U8475 (N_8475,N_8302,N_8287);
and U8476 (N_8476,N_8278,N_8233);
xor U8477 (N_8477,N_8322,N_8354);
and U8478 (N_8478,N_8316,N_8369);
or U8479 (N_8479,N_8293,N_8208);
or U8480 (N_8480,N_8307,N_8346);
nand U8481 (N_8481,N_8359,N_8240);
and U8482 (N_8482,N_8397,N_8323);
nor U8483 (N_8483,N_8308,N_8329);
and U8484 (N_8484,N_8371,N_8219);
xnor U8485 (N_8485,N_8292,N_8283);
nand U8486 (N_8486,N_8382,N_8205);
nand U8487 (N_8487,N_8272,N_8273);
or U8488 (N_8488,N_8276,N_8318);
xnor U8489 (N_8489,N_8304,N_8237);
xor U8490 (N_8490,N_8230,N_8385);
xnor U8491 (N_8491,N_8218,N_8301);
xnor U8492 (N_8492,N_8270,N_8357);
and U8493 (N_8493,N_8333,N_8349);
or U8494 (N_8494,N_8334,N_8220);
and U8495 (N_8495,N_8355,N_8281);
xor U8496 (N_8496,N_8311,N_8315);
and U8497 (N_8497,N_8383,N_8366);
nand U8498 (N_8498,N_8358,N_8249);
and U8499 (N_8499,N_8364,N_8350);
and U8500 (N_8500,N_8270,N_8210);
nand U8501 (N_8501,N_8383,N_8209);
and U8502 (N_8502,N_8269,N_8351);
and U8503 (N_8503,N_8316,N_8310);
xor U8504 (N_8504,N_8388,N_8346);
nand U8505 (N_8505,N_8259,N_8250);
and U8506 (N_8506,N_8296,N_8369);
xnor U8507 (N_8507,N_8294,N_8221);
xor U8508 (N_8508,N_8293,N_8228);
or U8509 (N_8509,N_8343,N_8247);
xnor U8510 (N_8510,N_8320,N_8364);
xnor U8511 (N_8511,N_8300,N_8365);
nor U8512 (N_8512,N_8346,N_8249);
and U8513 (N_8513,N_8373,N_8389);
or U8514 (N_8514,N_8304,N_8246);
nand U8515 (N_8515,N_8274,N_8216);
or U8516 (N_8516,N_8338,N_8367);
or U8517 (N_8517,N_8351,N_8304);
nor U8518 (N_8518,N_8375,N_8205);
xnor U8519 (N_8519,N_8352,N_8353);
and U8520 (N_8520,N_8388,N_8342);
or U8521 (N_8521,N_8265,N_8385);
xnor U8522 (N_8522,N_8251,N_8378);
nor U8523 (N_8523,N_8348,N_8398);
and U8524 (N_8524,N_8202,N_8253);
or U8525 (N_8525,N_8343,N_8393);
nor U8526 (N_8526,N_8304,N_8303);
nor U8527 (N_8527,N_8290,N_8389);
or U8528 (N_8528,N_8311,N_8301);
or U8529 (N_8529,N_8322,N_8363);
xor U8530 (N_8530,N_8218,N_8211);
nor U8531 (N_8531,N_8354,N_8338);
and U8532 (N_8532,N_8217,N_8238);
or U8533 (N_8533,N_8225,N_8263);
nor U8534 (N_8534,N_8362,N_8288);
nand U8535 (N_8535,N_8356,N_8273);
nand U8536 (N_8536,N_8387,N_8328);
xor U8537 (N_8537,N_8356,N_8223);
and U8538 (N_8538,N_8232,N_8387);
xnor U8539 (N_8539,N_8247,N_8270);
nor U8540 (N_8540,N_8274,N_8335);
xnor U8541 (N_8541,N_8281,N_8313);
xor U8542 (N_8542,N_8335,N_8367);
xor U8543 (N_8543,N_8300,N_8394);
xnor U8544 (N_8544,N_8362,N_8238);
nor U8545 (N_8545,N_8279,N_8322);
xor U8546 (N_8546,N_8250,N_8227);
xnor U8547 (N_8547,N_8295,N_8284);
nor U8548 (N_8548,N_8211,N_8225);
nor U8549 (N_8549,N_8205,N_8313);
xnor U8550 (N_8550,N_8395,N_8302);
and U8551 (N_8551,N_8242,N_8304);
xnor U8552 (N_8552,N_8243,N_8351);
nor U8553 (N_8553,N_8384,N_8211);
and U8554 (N_8554,N_8223,N_8254);
nor U8555 (N_8555,N_8371,N_8230);
xor U8556 (N_8556,N_8332,N_8366);
or U8557 (N_8557,N_8225,N_8247);
or U8558 (N_8558,N_8333,N_8295);
nand U8559 (N_8559,N_8391,N_8356);
nand U8560 (N_8560,N_8258,N_8292);
or U8561 (N_8561,N_8396,N_8203);
or U8562 (N_8562,N_8203,N_8266);
and U8563 (N_8563,N_8281,N_8308);
or U8564 (N_8564,N_8287,N_8216);
nor U8565 (N_8565,N_8206,N_8208);
nor U8566 (N_8566,N_8362,N_8370);
nor U8567 (N_8567,N_8388,N_8282);
nor U8568 (N_8568,N_8348,N_8248);
or U8569 (N_8569,N_8337,N_8397);
nor U8570 (N_8570,N_8397,N_8350);
or U8571 (N_8571,N_8265,N_8219);
nor U8572 (N_8572,N_8336,N_8261);
and U8573 (N_8573,N_8298,N_8323);
or U8574 (N_8574,N_8368,N_8276);
and U8575 (N_8575,N_8369,N_8300);
and U8576 (N_8576,N_8305,N_8270);
or U8577 (N_8577,N_8334,N_8303);
or U8578 (N_8578,N_8232,N_8244);
xnor U8579 (N_8579,N_8270,N_8216);
nand U8580 (N_8580,N_8370,N_8291);
nor U8581 (N_8581,N_8392,N_8271);
or U8582 (N_8582,N_8360,N_8248);
and U8583 (N_8583,N_8349,N_8297);
and U8584 (N_8584,N_8343,N_8296);
nand U8585 (N_8585,N_8228,N_8301);
nor U8586 (N_8586,N_8262,N_8227);
nand U8587 (N_8587,N_8232,N_8313);
or U8588 (N_8588,N_8307,N_8276);
and U8589 (N_8589,N_8371,N_8314);
nor U8590 (N_8590,N_8381,N_8291);
nand U8591 (N_8591,N_8293,N_8359);
xor U8592 (N_8592,N_8272,N_8202);
xor U8593 (N_8593,N_8277,N_8350);
nand U8594 (N_8594,N_8268,N_8324);
nand U8595 (N_8595,N_8250,N_8261);
and U8596 (N_8596,N_8210,N_8310);
nand U8597 (N_8597,N_8317,N_8284);
nand U8598 (N_8598,N_8312,N_8374);
or U8599 (N_8599,N_8360,N_8245);
nand U8600 (N_8600,N_8483,N_8431);
or U8601 (N_8601,N_8430,N_8475);
nand U8602 (N_8602,N_8452,N_8444);
and U8603 (N_8603,N_8491,N_8594);
nor U8604 (N_8604,N_8480,N_8423);
nand U8605 (N_8605,N_8525,N_8409);
nand U8606 (N_8606,N_8599,N_8554);
xor U8607 (N_8607,N_8546,N_8582);
and U8608 (N_8608,N_8580,N_8528);
xor U8609 (N_8609,N_8569,N_8521);
or U8610 (N_8610,N_8576,N_8403);
nor U8611 (N_8611,N_8587,N_8417);
nand U8612 (N_8612,N_8541,N_8413);
nor U8613 (N_8613,N_8435,N_8468);
nor U8614 (N_8614,N_8451,N_8448);
or U8615 (N_8615,N_8586,N_8552);
or U8616 (N_8616,N_8459,N_8527);
or U8617 (N_8617,N_8426,N_8505);
and U8618 (N_8618,N_8581,N_8490);
nor U8619 (N_8619,N_8593,N_8519);
nor U8620 (N_8620,N_8537,N_8410);
nand U8621 (N_8621,N_8566,N_8415);
xnor U8622 (N_8622,N_8400,N_8469);
or U8623 (N_8623,N_8463,N_8484);
and U8624 (N_8624,N_8447,N_8588);
nor U8625 (N_8625,N_8590,N_8473);
nor U8626 (N_8626,N_8474,N_8460);
nor U8627 (N_8627,N_8511,N_8557);
xor U8628 (N_8628,N_8532,N_8436);
and U8629 (N_8629,N_8579,N_8573);
xnor U8630 (N_8630,N_8553,N_8407);
nor U8631 (N_8631,N_8536,N_8467);
or U8632 (N_8632,N_8524,N_8405);
or U8633 (N_8633,N_8424,N_8425);
nor U8634 (N_8634,N_8501,N_8560);
or U8635 (N_8635,N_8564,N_8476);
and U8636 (N_8636,N_8558,N_8438);
and U8637 (N_8637,N_8464,N_8496);
or U8638 (N_8638,N_8535,N_8517);
nand U8639 (N_8639,N_8455,N_8445);
nor U8640 (N_8640,N_8465,N_8562);
and U8641 (N_8641,N_8595,N_8515);
or U8642 (N_8642,N_8548,N_8457);
or U8643 (N_8643,N_8478,N_8578);
xor U8644 (N_8644,N_8518,N_8549);
and U8645 (N_8645,N_8495,N_8477);
nor U8646 (N_8646,N_8509,N_8555);
or U8647 (N_8647,N_8456,N_8513);
nor U8648 (N_8648,N_8493,N_8497);
or U8649 (N_8649,N_8449,N_8544);
xor U8650 (N_8650,N_8499,N_8563);
nand U8651 (N_8651,N_8494,N_8520);
and U8652 (N_8652,N_8500,N_8462);
or U8653 (N_8653,N_8487,N_8538);
xnor U8654 (N_8654,N_8433,N_8547);
nor U8655 (N_8655,N_8550,N_8420);
nand U8656 (N_8656,N_8440,N_8577);
or U8657 (N_8657,N_8418,N_8437);
xor U8658 (N_8658,N_8523,N_8529);
or U8659 (N_8659,N_8568,N_8543);
or U8660 (N_8660,N_8488,N_8504);
nor U8661 (N_8661,N_8453,N_8570);
nand U8662 (N_8662,N_8598,N_8416);
nor U8663 (N_8663,N_8470,N_8565);
nand U8664 (N_8664,N_8571,N_8506);
nand U8665 (N_8665,N_8402,N_8585);
nor U8666 (N_8666,N_8439,N_8510);
nor U8667 (N_8667,N_8572,N_8592);
nor U8668 (N_8668,N_8406,N_8419);
and U8669 (N_8669,N_8472,N_8404);
nand U8670 (N_8670,N_8533,N_8486);
nor U8671 (N_8671,N_8530,N_8503);
nor U8672 (N_8672,N_8498,N_8561);
xor U8673 (N_8673,N_8461,N_8584);
nand U8674 (N_8674,N_8454,N_8507);
xnor U8675 (N_8675,N_8539,N_8591);
and U8676 (N_8676,N_8575,N_8485);
nor U8677 (N_8677,N_8567,N_8422);
xor U8678 (N_8678,N_8512,N_8442);
and U8679 (N_8679,N_8482,N_8551);
or U8680 (N_8680,N_8489,N_8421);
or U8681 (N_8681,N_8556,N_8574);
nor U8682 (N_8682,N_8545,N_8589);
xnor U8683 (N_8683,N_8412,N_8434);
and U8684 (N_8684,N_8427,N_8479);
and U8685 (N_8685,N_8471,N_8542);
and U8686 (N_8686,N_8559,N_8583);
nand U8687 (N_8687,N_8514,N_8596);
or U8688 (N_8688,N_8414,N_8441);
xor U8689 (N_8689,N_8446,N_8481);
nor U8690 (N_8690,N_8443,N_8597);
and U8691 (N_8691,N_8531,N_8411);
or U8692 (N_8692,N_8540,N_8508);
or U8693 (N_8693,N_8429,N_8502);
nand U8694 (N_8694,N_8458,N_8401);
nand U8695 (N_8695,N_8432,N_8516);
nand U8696 (N_8696,N_8526,N_8534);
xor U8697 (N_8697,N_8408,N_8450);
nand U8698 (N_8698,N_8522,N_8466);
and U8699 (N_8699,N_8492,N_8428);
nor U8700 (N_8700,N_8598,N_8542);
and U8701 (N_8701,N_8571,N_8429);
nor U8702 (N_8702,N_8538,N_8457);
nor U8703 (N_8703,N_8567,N_8531);
nor U8704 (N_8704,N_8586,N_8590);
nor U8705 (N_8705,N_8570,N_8585);
and U8706 (N_8706,N_8431,N_8478);
or U8707 (N_8707,N_8470,N_8532);
nand U8708 (N_8708,N_8410,N_8418);
nor U8709 (N_8709,N_8429,N_8587);
xnor U8710 (N_8710,N_8472,N_8402);
or U8711 (N_8711,N_8557,N_8500);
nand U8712 (N_8712,N_8559,N_8495);
nor U8713 (N_8713,N_8459,N_8437);
and U8714 (N_8714,N_8463,N_8593);
and U8715 (N_8715,N_8588,N_8489);
xnor U8716 (N_8716,N_8535,N_8468);
or U8717 (N_8717,N_8530,N_8565);
and U8718 (N_8718,N_8401,N_8421);
nand U8719 (N_8719,N_8475,N_8549);
or U8720 (N_8720,N_8497,N_8563);
and U8721 (N_8721,N_8596,N_8413);
and U8722 (N_8722,N_8443,N_8578);
or U8723 (N_8723,N_8505,N_8461);
and U8724 (N_8724,N_8416,N_8439);
xor U8725 (N_8725,N_8504,N_8579);
nand U8726 (N_8726,N_8564,N_8557);
and U8727 (N_8727,N_8508,N_8453);
nor U8728 (N_8728,N_8403,N_8416);
xor U8729 (N_8729,N_8574,N_8485);
and U8730 (N_8730,N_8432,N_8501);
nand U8731 (N_8731,N_8562,N_8565);
and U8732 (N_8732,N_8594,N_8575);
and U8733 (N_8733,N_8569,N_8545);
or U8734 (N_8734,N_8494,N_8435);
nor U8735 (N_8735,N_8423,N_8545);
nand U8736 (N_8736,N_8493,N_8500);
or U8737 (N_8737,N_8559,N_8568);
nor U8738 (N_8738,N_8576,N_8593);
nand U8739 (N_8739,N_8489,N_8425);
and U8740 (N_8740,N_8418,N_8594);
or U8741 (N_8741,N_8511,N_8403);
nand U8742 (N_8742,N_8540,N_8529);
or U8743 (N_8743,N_8567,N_8421);
xor U8744 (N_8744,N_8569,N_8537);
nor U8745 (N_8745,N_8522,N_8545);
nand U8746 (N_8746,N_8479,N_8556);
nand U8747 (N_8747,N_8428,N_8511);
or U8748 (N_8748,N_8420,N_8541);
nor U8749 (N_8749,N_8546,N_8419);
or U8750 (N_8750,N_8580,N_8530);
nor U8751 (N_8751,N_8458,N_8495);
nand U8752 (N_8752,N_8542,N_8447);
nor U8753 (N_8753,N_8483,N_8468);
and U8754 (N_8754,N_8407,N_8550);
xor U8755 (N_8755,N_8465,N_8596);
nand U8756 (N_8756,N_8426,N_8434);
and U8757 (N_8757,N_8583,N_8488);
or U8758 (N_8758,N_8422,N_8536);
or U8759 (N_8759,N_8585,N_8546);
or U8760 (N_8760,N_8455,N_8430);
and U8761 (N_8761,N_8447,N_8493);
nand U8762 (N_8762,N_8518,N_8501);
xnor U8763 (N_8763,N_8509,N_8437);
nor U8764 (N_8764,N_8547,N_8508);
nand U8765 (N_8765,N_8551,N_8517);
xnor U8766 (N_8766,N_8480,N_8485);
nand U8767 (N_8767,N_8460,N_8419);
or U8768 (N_8768,N_8489,N_8420);
nor U8769 (N_8769,N_8478,N_8523);
xor U8770 (N_8770,N_8538,N_8479);
xor U8771 (N_8771,N_8506,N_8561);
nor U8772 (N_8772,N_8485,N_8532);
nand U8773 (N_8773,N_8531,N_8585);
nand U8774 (N_8774,N_8557,N_8527);
xnor U8775 (N_8775,N_8410,N_8541);
xor U8776 (N_8776,N_8587,N_8461);
and U8777 (N_8777,N_8479,N_8428);
and U8778 (N_8778,N_8504,N_8511);
xnor U8779 (N_8779,N_8445,N_8426);
and U8780 (N_8780,N_8531,N_8501);
and U8781 (N_8781,N_8484,N_8410);
nand U8782 (N_8782,N_8433,N_8466);
xnor U8783 (N_8783,N_8525,N_8564);
and U8784 (N_8784,N_8471,N_8598);
xor U8785 (N_8785,N_8566,N_8594);
or U8786 (N_8786,N_8420,N_8414);
xor U8787 (N_8787,N_8581,N_8536);
xor U8788 (N_8788,N_8511,N_8524);
and U8789 (N_8789,N_8579,N_8475);
nand U8790 (N_8790,N_8489,N_8579);
nand U8791 (N_8791,N_8592,N_8473);
or U8792 (N_8792,N_8475,N_8584);
nand U8793 (N_8793,N_8448,N_8427);
nand U8794 (N_8794,N_8433,N_8501);
or U8795 (N_8795,N_8466,N_8515);
or U8796 (N_8796,N_8562,N_8409);
nand U8797 (N_8797,N_8548,N_8404);
nand U8798 (N_8798,N_8521,N_8461);
or U8799 (N_8799,N_8550,N_8524);
or U8800 (N_8800,N_8689,N_8693);
nor U8801 (N_8801,N_8764,N_8673);
nand U8802 (N_8802,N_8615,N_8712);
nand U8803 (N_8803,N_8748,N_8601);
nand U8804 (N_8804,N_8684,N_8759);
nand U8805 (N_8805,N_8702,N_8637);
or U8806 (N_8806,N_8705,N_8682);
nand U8807 (N_8807,N_8762,N_8799);
and U8808 (N_8808,N_8715,N_8600);
nand U8809 (N_8809,N_8686,N_8633);
xnor U8810 (N_8810,N_8641,N_8758);
nor U8811 (N_8811,N_8740,N_8630);
and U8812 (N_8812,N_8605,N_8646);
and U8813 (N_8813,N_8781,N_8683);
xor U8814 (N_8814,N_8717,N_8798);
nand U8815 (N_8815,N_8733,N_8794);
and U8816 (N_8816,N_8716,N_8743);
xor U8817 (N_8817,N_8729,N_8738);
nor U8818 (N_8818,N_8626,N_8661);
and U8819 (N_8819,N_8741,N_8776);
nand U8820 (N_8820,N_8709,N_8778);
nor U8821 (N_8821,N_8644,N_8657);
and U8822 (N_8822,N_8660,N_8621);
nor U8823 (N_8823,N_8666,N_8674);
xnor U8824 (N_8824,N_8791,N_8779);
or U8825 (N_8825,N_8728,N_8749);
nand U8826 (N_8826,N_8632,N_8659);
nor U8827 (N_8827,N_8730,N_8732);
and U8828 (N_8828,N_8676,N_8628);
nand U8829 (N_8829,N_8649,N_8651);
and U8830 (N_8830,N_8670,N_8752);
or U8831 (N_8831,N_8763,N_8648);
xor U8832 (N_8832,N_8701,N_8620);
and U8833 (N_8833,N_8707,N_8662);
or U8834 (N_8834,N_8720,N_8747);
nand U8835 (N_8835,N_8796,N_8671);
or U8836 (N_8836,N_8681,N_8767);
nor U8837 (N_8837,N_8669,N_8617);
or U8838 (N_8838,N_8777,N_8607);
xnor U8839 (N_8839,N_8770,N_8640);
or U8840 (N_8840,N_8725,N_8692);
and U8841 (N_8841,N_8766,N_8606);
or U8842 (N_8842,N_8624,N_8687);
and U8843 (N_8843,N_8698,N_8695);
or U8844 (N_8844,N_8751,N_8718);
nand U8845 (N_8845,N_8629,N_8634);
and U8846 (N_8846,N_8723,N_8727);
and U8847 (N_8847,N_8616,N_8719);
nand U8848 (N_8848,N_8688,N_8735);
nand U8849 (N_8849,N_8639,N_8614);
and U8850 (N_8850,N_8775,N_8699);
and U8851 (N_8851,N_8754,N_8736);
nand U8852 (N_8852,N_8773,N_8619);
xor U8853 (N_8853,N_8787,N_8610);
and U8854 (N_8854,N_8772,N_8788);
nor U8855 (N_8855,N_8726,N_8677);
or U8856 (N_8856,N_8782,N_8653);
xnor U8857 (N_8857,N_8746,N_8643);
or U8858 (N_8858,N_8737,N_8608);
xnor U8859 (N_8859,N_8724,N_8745);
or U8860 (N_8860,N_8645,N_8647);
nor U8861 (N_8861,N_8721,N_8734);
nand U8862 (N_8862,N_8706,N_8714);
nand U8863 (N_8863,N_8622,N_8690);
xnor U8864 (N_8864,N_8700,N_8786);
nor U8865 (N_8865,N_8631,N_8769);
xnor U8866 (N_8866,N_8744,N_8672);
xor U8867 (N_8867,N_8783,N_8656);
nand U8868 (N_8868,N_8755,N_8685);
and U8869 (N_8869,N_8792,N_8774);
nor U8870 (N_8870,N_8710,N_8795);
nor U8871 (N_8871,N_8625,N_8739);
nand U8872 (N_8872,N_8635,N_8636);
and U8873 (N_8873,N_8785,N_8678);
or U8874 (N_8874,N_8658,N_8731);
xor U8875 (N_8875,N_8703,N_8768);
nand U8876 (N_8876,N_8765,N_8722);
or U8877 (N_8877,N_8789,N_8694);
nor U8878 (N_8878,N_8753,N_8623);
nand U8879 (N_8879,N_8680,N_8771);
nand U8880 (N_8880,N_8790,N_8613);
or U8881 (N_8881,N_8655,N_8611);
and U8882 (N_8882,N_8609,N_8760);
or U8883 (N_8883,N_8704,N_8652);
xor U8884 (N_8884,N_8627,N_8780);
or U8885 (N_8885,N_8654,N_8793);
nor U8886 (N_8886,N_8642,N_8602);
xor U8887 (N_8887,N_8797,N_8742);
nor U8888 (N_8888,N_8713,N_8679);
xnor U8889 (N_8889,N_8756,N_8604);
xor U8890 (N_8890,N_8750,N_8664);
or U8891 (N_8891,N_8603,N_8697);
and U8892 (N_8892,N_8757,N_8668);
and U8893 (N_8893,N_8784,N_8711);
nand U8894 (N_8894,N_8691,N_8665);
or U8895 (N_8895,N_8618,N_8708);
nand U8896 (N_8896,N_8675,N_8761);
nor U8897 (N_8897,N_8612,N_8650);
xor U8898 (N_8898,N_8696,N_8638);
or U8899 (N_8899,N_8663,N_8667);
xnor U8900 (N_8900,N_8797,N_8619);
or U8901 (N_8901,N_8696,N_8775);
nand U8902 (N_8902,N_8677,N_8723);
nor U8903 (N_8903,N_8675,N_8731);
nor U8904 (N_8904,N_8749,N_8740);
nand U8905 (N_8905,N_8671,N_8700);
or U8906 (N_8906,N_8765,N_8785);
or U8907 (N_8907,N_8622,N_8792);
nand U8908 (N_8908,N_8719,N_8611);
xor U8909 (N_8909,N_8783,N_8639);
or U8910 (N_8910,N_8714,N_8735);
xor U8911 (N_8911,N_8722,N_8662);
nor U8912 (N_8912,N_8660,N_8735);
nand U8913 (N_8913,N_8754,N_8638);
xnor U8914 (N_8914,N_8707,N_8639);
or U8915 (N_8915,N_8742,N_8697);
xor U8916 (N_8916,N_8689,N_8799);
and U8917 (N_8917,N_8726,N_8681);
or U8918 (N_8918,N_8744,N_8789);
nand U8919 (N_8919,N_8635,N_8662);
and U8920 (N_8920,N_8796,N_8795);
or U8921 (N_8921,N_8773,N_8797);
and U8922 (N_8922,N_8631,N_8652);
nand U8923 (N_8923,N_8614,N_8613);
nand U8924 (N_8924,N_8703,N_8677);
and U8925 (N_8925,N_8720,N_8670);
and U8926 (N_8926,N_8725,N_8691);
or U8927 (N_8927,N_8656,N_8799);
nor U8928 (N_8928,N_8637,N_8707);
xor U8929 (N_8929,N_8795,N_8686);
nand U8930 (N_8930,N_8788,N_8621);
and U8931 (N_8931,N_8631,N_8634);
and U8932 (N_8932,N_8752,N_8716);
nor U8933 (N_8933,N_8647,N_8794);
nor U8934 (N_8934,N_8685,N_8746);
nor U8935 (N_8935,N_8701,N_8728);
or U8936 (N_8936,N_8788,N_8704);
and U8937 (N_8937,N_8636,N_8714);
xor U8938 (N_8938,N_8713,N_8674);
xnor U8939 (N_8939,N_8619,N_8783);
nand U8940 (N_8940,N_8693,N_8798);
and U8941 (N_8941,N_8674,N_8623);
nor U8942 (N_8942,N_8702,N_8602);
or U8943 (N_8943,N_8611,N_8630);
nand U8944 (N_8944,N_8727,N_8600);
xnor U8945 (N_8945,N_8690,N_8686);
xnor U8946 (N_8946,N_8715,N_8669);
or U8947 (N_8947,N_8784,N_8616);
nand U8948 (N_8948,N_8667,N_8711);
xnor U8949 (N_8949,N_8747,N_8783);
nor U8950 (N_8950,N_8762,N_8781);
nand U8951 (N_8951,N_8793,N_8635);
xor U8952 (N_8952,N_8733,N_8751);
xor U8953 (N_8953,N_8755,N_8674);
xor U8954 (N_8954,N_8754,N_8664);
or U8955 (N_8955,N_8678,N_8740);
or U8956 (N_8956,N_8763,N_8711);
or U8957 (N_8957,N_8740,N_8719);
and U8958 (N_8958,N_8601,N_8610);
xor U8959 (N_8959,N_8654,N_8743);
nor U8960 (N_8960,N_8769,N_8609);
or U8961 (N_8961,N_8771,N_8763);
and U8962 (N_8962,N_8689,N_8716);
xnor U8963 (N_8963,N_8653,N_8658);
nand U8964 (N_8964,N_8735,N_8629);
or U8965 (N_8965,N_8633,N_8740);
and U8966 (N_8966,N_8636,N_8661);
or U8967 (N_8967,N_8655,N_8728);
nand U8968 (N_8968,N_8780,N_8657);
nor U8969 (N_8969,N_8782,N_8771);
nand U8970 (N_8970,N_8669,N_8659);
nand U8971 (N_8971,N_8607,N_8705);
nor U8972 (N_8972,N_8709,N_8649);
xor U8973 (N_8973,N_8731,N_8683);
or U8974 (N_8974,N_8795,N_8702);
or U8975 (N_8975,N_8722,N_8644);
or U8976 (N_8976,N_8693,N_8692);
and U8977 (N_8977,N_8693,N_8794);
xor U8978 (N_8978,N_8605,N_8691);
and U8979 (N_8979,N_8670,N_8757);
xor U8980 (N_8980,N_8714,N_8716);
and U8981 (N_8981,N_8601,N_8621);
nor U8982 (N_8982,N_8695,N_8791);
nand U8983 (N_8983,N_8684,N_8738);
xor U8984 (N_8984,N_8631,N_8645);
and U8985 (N_8985,N_8769,N_8727);
and U8986 (N_8986,N_8611,N_8746);
xnor U8987 (N_8987,N_8714,N_8749);
nand U8988 (N_8988,N_8609,N_8671);
and U8989 (N_8989,N_8787,N_8635);
xnor U8990 (N_8990,N_8622,N_8764);
nor U8991 (N_8991,N_8792,N_8768);
and U8992 (N_8992,N_8688,N_8604);
or U8993 (N_8993,N_8683,N_8672);
nor U8994 (N_8994,N_8650,N_8648);
xnor U8995 (N_8995,N_8701,N_8708);
or U8996 (N_8996,N_8721,N_8603);
nand U8997 (N_8997,N_8647,N_8774);
nor U8998 (N_8998,N_8795,N_8667);
nor U8999 (N_8999,N_8700,N_8645);
nor U9000 (N_9000,N_8997,N_8991);
xor U9001 (N_9001,N_8969,N_8871);
xnor U9002 (N_9002,N_8821,N_8957);
xnor U9003 (N_9003,N_8942,N_8899);
nand U9004 (N_9004,N_8838,N_8956);
and U9005 (N_9005,N_8849,N_8861);
nor U9006 (N_9006,N_8823,N_8912);
and U9007 (N_9007,N_8965,N_8852);
xor U9008 (N_9008,N_8843,N_8968);
nand U9009 (N_9009,N_8934,N_8963);
and U9010 (N_9010,N_8937,N_8847);
xor U9011 (N_9011,N_8954,N_8946);
or U9012 (N_9012,N_8911,N_8818);
and U9013 (N_9013,N_8864,N_8866);
or U9014 (N_9014,N_8862,N_8945);
nor U9015 (N_9015,N_8828,N_8897);
nor U9016 (N_9016,N_8887,N_8802);
and U9017 (N_9017,N_8856,N_8995);
or U9018 (N_9018,N_8872,N_8986);
and U9019 (N_9019,N_8851,N_8905);
and U9020 (N_9020,N_8984,N_8920);
or U9021 (N_9021,N_8904,N_8848);
xor U9022 (N_9022,N_8931,N_8839);
nor U9023 (N_9023,N_8830,N_8987);
or U9024 (N_9024,N_8967,N_8982);
nor U9025 (N_9025,N_8894,N_8827);
and U9026 (N_9026,N_8998,N_8898);
xnor U9027 (N_9027,N_8890,N_8816);
and U9028 (N_9028,N_8907,N_8961);
nand U9029 (N_9029,N_8921,N_8855);
or U9030 (N_9030,N_8959,N_8836);
nor U9031 (N_9031,N_8869,N_8914);
or U9032 (N_9032,N_8973,N_8810);
or U9033 (N_9033,N_8814,N_8983);
nor U9034 (N_9034,N_8908,N_8892);
or U9035 (N_9035,N_8901,N_8875);
and U9036 (N_9036,N_8845,N_8955);
nand U9037 (N_9037,N_8903,N_8980);
nand U9038 (N_9038,N_8859,N_8835);
or U9039 (N_9039,N_8943,N_8803);
nor U9040 (N_9040,N_8981,N_8972);
xor U9041 (N_9041,N_8841,N_8886);
nor U9042 (N_9042,N_8840,N_8906);
nor U9043 (N_9043,N_8976,N_8993);
nand U9044 (N_9044,N_8999,N_8868);
or U9045 (N_9045,N_8834,N_8878);
nand U9046 (N_9046,N_8933,N_8979);
or U9047 (N_9047,N_8917,N_8985);
or U9048 (N_9048,N_8817,N_8910);
nor U9049 (N_9049,N_8923,N_8815);
and U9050 (N_9050,N_8889,N_8813);
nor U9051 (N_9051,N_8974,N_8831);
xor U9052 (N_9052,N_8951,N_8927);
nand U9053 (N_9053,N_8833,N_8873);
xnor U9054 (N_9054,N_8950,N_8806);
xor U9055 (N_9055,N_8844,N_8884);
xnor U9056 (N_9056,N_8807,N_8900);
nor U9057 (N_9057,N_8800,N_8918);
xnor U9058 (N_9058,N_8883,N_8978);
nor U9059 (N_9059,N_8885,N_8936);
nand U9060 (N_9060,N_8867,N_8819);
and U9061 (N_9061,N_8895,N_8826);
or U9062 (N_9062,N_8915,N_8822);
nor U9063 (N_9063,N_8939,N_8928);
nand U9064 (N_9064,N_8857,N_8870);
xnor U9065 (N_9065,N_8820,N_8876);
and U9066 (N_9066,N_8854,N_8925);
nand U9067 (N_9067,N_8804,N_8811);
nor U9068 (N_9068,N_8891,N_8874);
nand U9069 (N_9069,N_8846,N_8926);
xor U9070 (N_9070,N_8958,N_8953);
and U9071 (N_9071,N_8832,N_8948);
and U9072 (N_9072,N_8808,N_8938);
nand U9073 (N_9073,N_8909,N_8941);
xnor U9074 (N_9074,N_8922,N_8971);
and U9075 (N_9075,N_8829,N_8805);
xor U9076 (N_9076,N_8837,N_8994);
and U9077 (N_9077,N_8977,N_8880);
and U9078 (N_9078,N_8893,N_8932);
xor U9079 (N_9079,N_8970,N_8850);
xor U9080 (N_9080,N_8992,N_8988);
and U9081 (N_9081,N_8881,N_8919);
and U9082 (N_9082,N_8949,N_8975);
nand U9083 (N_9083,N_8842,N_8877);
nor U9084 (N_9084,N_8809,N_8888);
nand U9085 (N_9085,N_8962,N_8929);
or U9086 (N_9086,N_8916,N_8947);
and U9087 (N_9087,N_8902,N_8940);
nor U9088 (N_9088,N_8930,N_8812);
or U9089 (N_9089,N_8879,N_8853);
xor U9090 (N_9090,N_8960,N_8824);
nor U9091 (N_9091,N_8924,N_8913);
xor U9092 (N_9092,N_8935,N_8964);
xor U9093 (N_9093,N_8882,N_8865);
and U9094 (N_9094,N_8944,N_8863);
or U9095 (N_9095,N_8860,N_8989);
xor U9096 (N_9096,N_8996,N_8858);
nor U9097 (N_9097,N_8990,N_8825);
xnor U9098 (N_9098,N_8801,N_8896);
and U9099 (N_9099,N_8966,N_8952);
nand U9100 (N_9100,N_8831,N_8816);
or U9101 (N_9101,N_8857,N_8959);
xnor U9102 (N_9102,N_8887,N_8979);
xnor U9103 (N_9103,N_8839,N_8882);
xnor U9104 (N_9104,N_8911,N_8868);
xnor U9105 (N_9105,N_8997,N_8940);
nor U9106 (N_9106,N_8884,N_8980);
xnor U9107 (N_9107,N_8849,N_8923);
or U9108 (N_9108,N_8898,N_8839);
and U9109 (N_9109,N_8925,N_8832);
nor U9110 (N_9110,N_8882,N_8978);
nand U9111 (N_9111,N_8979,N_8828);
and U9112 (N_9112,N_8852,N_8921);
or U9113 (N_9113,N_8892,N_8857);
xor U9114 (N_9114,N_8885,N_8827);
xor U9115 (N_9115,N_8896,N_8853);
xnor U9116 (N_9116,N_8985,N_8992);
nor U9117 (N_9117,N_8836,N_8872);
or U9118 (N_9118,N_8850,N_8847);
or U9119 (N_9119,N_8870,N_8841);
or U9120 (N_9120,N_8911,N_8816);
or U9121 (N_9121,N_8855,N_8968);
nor U9122 (N_9122,N_8964,N_8884);
and U9123 (N_9123,N_8803,N_8862);
nand U9124 (N_9124,N_8834,N_8868);
and U9125 (N_9125,N_8855,N_8876);
nand U9126 (N_9126,N_8829,N_8828);
nor U9127 (N_9127,N_8875,N_8933);
xor U9128 (N_9128,N_8873,N_8904);
and U9129 (N_9129,N_8965,N_8976);
or U9130 (N_9130,N_8875,N_8909);
or U9131 (N_9131,N_8824,N_8987);
xor U9132 (N_9132,N_8867,N_8938);
xnor U9133 (N_9133,N_8861,N_8969);
and U9134 (N_9134,N_8919,N_8859);
xnor U9135 (N_9135,N_8841,N_8882);
or U9136 (N_9136,N_8899,N_8964);
and U9137 (N_9137,N_8862,N_8886);
and U9138 (N_9138,N_8946,N_8909);
or U9139 (N_9139,N_8936,N_8813);
or U9140 (N_9140,N_8997,N_8944);
nand U9141 (N_9141,N_8956,N_8831);
nor U9142 (N_9142,N_8938,N_8837);
and U9143 (N_9143,N_8993,N_8848);
xnor U9144 (N_9144,N_8832,N_8909);
or U9145 (N_9145,N_8854,N_8957);
nand U9146 (N_9146,N_8870,N_8934);
nand U9147 (N_9147,N_8861,N_8996);
nand U9148 (N_9148,N_8962,N_8807);
nor U9149 (N_9149,N_8912,N_8966);
nand U9150 (N_9150,N_8949,N_8947);
nand U9151 (N_9151,N_8988,N_8840);
nor U9152 (N_9152,N_8870,N_8901);
xnor U9153 (N_9153,N_8970,N_8995);
xnor U9154 (N_9154,N_8974,N_8878);
nor U9155 (N_9155,N_8981,N_8967);
xor U9156 (N_9156,N_8830,N_8900);
nor U9157 (N_9157,N_8977,N_8920);
or U9158 (N_9158,N_8863,N_8823);
and U9159 (N_9159,N_8917,N_8824);
xor U9160 (N_9160,N_8937,N_8832);
nor U9161 (N_9161,N_8964,N_8828);
and U9162 (N_9162,N_8872,N_8929);
nand U9163 (N_9163,N_8830,N_8961);
and U9164 (N_9164,N_8882,N_8971);
nor U9165 (N_9165,N_8863,N_8800);
xor U9166 (N_9166,N_8833,N_8923);
or U9167 (N_9167,N_8813,N_8958);
or U9168 (N_9168,N_8864,N_8985);
xnor U9169 (N_9169,N_8933,N_8906);
xnor U9170 (N_9170,N_8934,N_8863);
nor U9171 (N_9171,N_8829,N_8979);
nand U9172 (N_9172,N_8854,N_8901);
and U9173 (N_9173,N_8960,N_8951);
nor U9174 (N_9174,N_8991,N_8949);
nand U9175 (N_9175,N_8913,N_8956);
nor U9176 (N_9176,N_8903,N_8833);
nand U9177 (N_9177,N_8903,N_8808);
nand U9178 (N_9178,N_8919,N_8802);
xor U9179 (N_9179,N_8977,N_8961);
nand U9180 (N_9180,N_8933,N_8805);
xnor U9181 (N_9181,N_8810,N_8979);
and U9182 (N_9182,N_8943,N_8915);
nand U9183 (N_9183,N_8946,N_8920);
nand U9184 (N_9184,N_8987,N_8921);
nor U9185 (N_9185,N_8864,N_8825);
xor U9186 (N_9186,N_8973,N_8907);
xnor U9187 (N_9187,N_8977,N_8936);
nand U9188 (N_9188,N_8941,N_8973);
and U9189 (N_9189,N_8828,N_8937);
xnor U9190 (N_9190,N_8849,N_8807);
xor U9191 (N_9191,N_8864,N_8859);
xor U9192 (N_9192,N_8889,N_8841);
or U9193 (N_9193,N_8891,N_8957);
or U9194 (N_9194,N_8827,N_8981);
nand U9195 (N_9195,N_8991,N_8921);
nor U9196 (N_9196,N_8854,N_8919);
nor U9197 (N_9197,N_8814,N_8942);
nand U9198 (N_9198,N_8902,N_8877);
and U9199 (N_9199,N_8963,N_8843);
nor U9200 (N_9200,N_9190,N_9155);
and U9201 (N_9201,N_9153,N_9067);
and U9202 (N_9202,N_9139,N_9183);
and U9203 (N_9203,N_9162,N_9115);
or U9204 (N_9204,N_9171,N_9077);
nor U9205 (N_9205,N_9130,N_9187);
nand U9206 (N_9206,N_9140,N_9091);
and U9207 (N_9207,N_9147,N_9109);
nand U9208 (N_9208,N_9020,N_9009);
and U9209 (N_9209,N_9176,N_9111);
and U9210 (N_9210,N_9074,N_9006);
nand U9211 (N_9211,N_9041,N_9141);
xnor U9212 (N_9212,N_9144,N_9088);
nor U9213 (N_9213,N_9035,N_9075);
and U9214 (N_9214,N_9045,N_9094);
xor U9215 (N_9215,N_9184,N_9134);
nand U9216 (N_9216,N_9182,N_9008);
and U9217 (N_9217,N_9096,N_9166);
and U9218 (N_9218,N_9178,N_9122);
nor U9219 (N_9219,N_9072,N_9159);
or U9220 (N_9220,N_9033,N_9031);
nand U9221 (N_9221,N_9185,N_9191);
or U9222 (N_9222,N_9152,N_9127);
nor U9223 (N_9223,N_9047,N_9012);
nor U9224 (N_9224,N_9118,N_9112);
nand U9225 (N_9225,N_9099,N_9108);
and U9226 (N_9226,N_9186,N_9192);
or U9227 (N_9227,N_9022,N_9005);
xnor U9228 (N_9228,N_9036,N_9040);
nor U9229 (N_9229,N_9063,N_9143);
nor U9230 (N_9230,N_9048,N_9053);
nand U9231 (N_9231,N_9007,N_9131);
or U9232 (N_9232,N_9049,N_9104);
and U9233 (N_9233,N_9093,N_9142);
and U9234 (N_9234,N_9170,N_9116);
xnor U9235 (N_9235,N_9055,N_9086);
or U9236 (N_9236,N_9107,N_9196);
nand U9237 (N_9237,N_9149,N_9117);
or U9238 (N_9238,N_9168,N_9114);
xnor U9239 (N_9239,N_9023,N_9061);
nand U9240 (N_9240,N_9081,N_9193);
xor U9241 (N_9241,N_9068,N_9058);
xnor U9242 (N_9242,N_9025,N_9100);
nor U9243 (N_9243,N_9121,N_9194);
and U9244 (N_9244,N_9199,N_9028);
xnor U9245 (N_9245,N_9060,N_9004);
xor U9246 (N_9246,N_9054,N_9129);
or U9247 (N_9247,N_9092,N_9039);
xor U9248 (N_9248,N_9137,N_9198);
nand U9249 (N_9249,N_9146,N_9034);
nand U9250 (N_9250,N_9135,N_9078);
nand U9251 (N_9251,N_9042,N_9110);
nand U9252 (N_9252,N_9064,N_9000);
nor U9253 (N_9253,N_9195,N_9043);
and U9254 (N_9254,N_9105,N_9090);
and U9255 (N_9255,N_9181,N_9026);
or U9256 (N_9256,N_9082,N_9016);
nor U9257 (N_9257,N_9103,N_9080);
nor U9258 (N_9258,N_9119,N_9002);
xnor U9259 (N_9259,N_9079,N_9070);
nand U9260 (N_9260,N_9057,N_9165);
nand U9261 (N_9261,N_9010,N_9133);
nand U9262 (N_9262,N_9017,N_9172);
nor U9263 (N_9263,N_9164,N_9138);
nor U9264 (N_9264,N_9071,N_9065);
and U9265 (N_9265,N_9052,N_9136);
or U9266 (N_9266,N_9106,N_9013);
or U9267 (N_9267,N_9145,N_9148);
and U9268 (N_9268,N_9128,N_9151);
xor U9269 (N_9269,N_9001,N_9188);
nand U9270 (N_9270,N_9156,N_9098);
xor U9271 (N_9271,N_9097,N_9024);
or U9272 (N_9272,N_9123,N_9180);
nor U9273 (N_9273,N_9038,N_9179);
or U9274 (N_9274,N_9037,N_9113);
nand U9275 (N_9275,N_9173,N_9021);
xor U9276 (N_9276,N_9101,N_9163);
xor U9277 (N_9277,N_9032,N_9158);
nand U9278 (N_9278,N_9083,N_9174);
or U9279 (N_9279,N_9167,N_9089);
nand U9280 (N_9280,N_9197,N_9069);
and U9281 (N_9281,N_9160,N_9169);
nand U9282 (N_9282,N_9014,N_9124);
and U9283 (N_9283,N_9003,N_9150);
nor U9284 (N_9284,N_9154,N_9015);
nor U9285 (N_9285,N_9019,N_9018);
or U9286 (N_9286,N_9050,N_9046);
or U9287 (N_9287,N_9161,N_9062);
and U9288 (N_9288,N_9087,N_9085);
xnor U9289 (N_9289,N_9044,N_9102);
xnor U9290 (N_9290,N_9029,N_9084);
nand U9291 (N_9291,N_9095,N_9177);
or U9292 (N_9292,N_9073,N_9189);
and U9293 (N_9293,N_9059,N_9120);
nor U9294 (N_9294,N_9157,N_9027);
nor U9295 (N_9295,N_9125,N_9056);
nor U9296 (N_9296,N_9126,N_9030);
or U9297 (N_9297,N_9051,N_9011);
xnor U9298 (N_9298,N_9066,N_9132);
or U9299 (N_9299,N_9076,N_9175);
xnor U9300 (N_9300,N_9139,N_9188);
or U9301 (N_9301,N_9141,N_9199);
and U9302 (N_9302,N_9108,N_9195);
nor U9303 (N_9303,N_9125,N_9122);
and U9304 (N_9304,N_9019,N_9051);
nor U9305 (N_9305,N_9000,N_9070);
or U9306 (N_9306,N_9157,N_9083);
nor U9307 (N_9307,N_9000,N_9096);
nor U9308 (N_9308,N_9080,N_9099);
nand U9309 (N_9309,N_9182,N_9101);
nand U9310 (N_9310,N_9141,N_9080);
nand U9311 (N_9311,N_9038,N_9147);
or U9312 (N_9312,N_9102,N_9053);
nand U9313 (N_9313,N_9130,N_9172);
nand U9314 (N_9314,N_9123,N_9046);
nor U9315 (N_9315,N_9025,N_9172);
nand U9316 (N_9316,N_9071,N_9114);
xor U9317 (N_9317,N_9082,N_9193);
nor U9318 (N_9318,N_9016,N_9182);
xor U9319 (N_9319,N_9093,N_9195);
and U9320 (N_9320,N_9172,N_9121);
or U9321 (N_9321,N_9199,N_9100);
nor U9322 (N_9322,N_9192,N_9181);
and U9323 (N_9323,N_9171,N_9031);
and U9324 (N_9324,N_9189,N_9065);
nor U9325 (N_9325,N_9024,N_9080);
nor U9326 (N_9326,N_9103,N_9025);
nor U9327 (N_9327,N_9196,N_9051);
nand U9328 (N_9328,N_9081,N_9149);
and U9329 (N_9329,N_9123,N_9027);
xor U9330 (N_9330,N_9145,N_9186);
or U9331 (N_9331,N_9086,N_9075);
xnor U9332 (N_9332,N_9037,N_9169);
xnor U9333 (N_9333,N_9005,N_9050);
or U9334 (N_9334,N_9104,N_9057);
or U9335 (N_9335,N_9086,N_9169);
nor U9336 (N_9336,N_9181,N_9024);
xor U9337 (N_9337,N_9072,N_9130);
or U9338 (N_9338,N_9197,N_9024);
xor U9339 (N_9339,N_9177,N_9014);
or U9340 (N_9340,N_9151,N_9184);
xnor U9341 (N_9341,N_9168,N_9126);
nand U9342 (N_9342,N_9128,N_9036);
xor U9343 (N_9343,N_9179,N_9044);
xnor U9344 (N_9344,N_9172,N_9101);
and U9345 (N_9345,N_9081,N_9128);
nor U9346 (N_9346,N_9126,N_9175);
xor U9347 (N_9347,N_9161,N_9050);
and U9348 (N_9348,N_9155,N_9168);
nand U9349 (N_9349,N_9057,N_9026);
nand U9350 (N_9350,N_9124,N_9065);
or U9351 (N_9351,N_9118,N_9170);
nor U9352 (N_9352,N_9103,N_9125);
nor U9353 (N_9353,N_9089,N_9005);
nor U9354 (N_9354,N_9073,N_9122);
or U9355 (N_9355,N_9012,N_9041);
nand U9356 (N_9356,N_9025,N_9053);
nand U9357 (N_9357,N_9120,N_9196);
xnor U9358 (N_9358,N_9033,N_9093);
nand U9359 (N_9359,N_9152,N_9131);
nor U9360 (N_9360,N_9081,N_9124);
nand U9361 (N_9361,N_9001,N_9096);
xnor U9362 (N_9362,N_9128,N_9078);
nand U9363 (N_9363,N_9042,N_9189);
or U9364 (N_9364,N_9141,N_9187);
xnor U9365 (N_9365,N_9049,N_9078);
or U9366 (N_9366,N_9001,N_9048);
and U9367 (N_9367,N_9118,N_9013);
nand U9368 (N_9368,N_9114,N_9081);
or U9369 (N_9369,N_9028,N_9153);
or U9370 (N_9370,N_9143,N_9100);
nand U9371 (N_9371,N_9110,N_9176);
and U9372 (N_9372,N_9140,N_9103);
nand U9373 (N_9373,N_9144,N_9155);
xnor U9374 (N_9374,N_9023,N_9152);
xor U9375 (N_9375,N_9090,N_9155);
or U9376 (N_9376,N_9118,N_9033);
nand U9377 (N_9377,N_9195,N_9055);
xor U9378 (N_9378,N_9024,N_9116);
xor U9379 (N_9379,N_9117,N_9089);
nor U9380 (N_9380,N_9083,N_9084);
nor U9381 (N_9381,N_9182,N_9163);
or U9382 (N_9382,N_9114,N_9162);
nor U9383 (N_9383,N_9071,N_9056);
nor U9384 (N_9384,N_9023,N_9022);
xnor U9385 (N_9385,N_9075,N_9128);
xnor U9386 (N_9386,N_9003,N_9156);
or U9387 (N_9387,N_9020,N_9179);
nor U9388 (N_9388,N_9199,N_9064);
xnor U9389 (N_9389,N_9054,N_9095);
or U9390 (N_9390,N_9056,N_9166);
nor U9391 (N_9391,N_9038,N_9033);
nand U9392 (N_9392,N_9112,N_9079);
nand U9393 (N_9393,N_9008,N_9031);
nand U9394 (N_9394,N_9086,N_9033);
nor U9395 (N_9395,N_9077,N_9109);
xor U9396 (N_9396,N_9163,N_9028);
xor U9397 (N_9397,N_9022,N_9099);
nand U9398 (N_9398,N_9168,N_9081);
and U9399 (N_9399,N_9185,N_9160);
nand U9400 (N_9400,N_9316,N_9381);
and U9401 (N_9401,N_9226,N_9367);
or U9402 (N_9402,N_9273,N_9286);
or U9403 (N_9403,N_9233,N_9338);
nand U9404 (N_9404,N_9205,N_9228);
or U9405 (N_9405,N_9330,N_9351);
and U9406 (N_9406,N_9312,N_9289);
xnor U9407 (N_9407,N_9325,N_9239);
nor U9408 (N_9408,N_9269,N_9274);
nand U9409 (N_9409,N_9279,N_9272);
and U9410 (N_9410,N_9232,N_9308);
or U9411 (N_9411,N_9378,N_9212);
nor U9412 (N_9412,N_9314,N_9298);
xor U9413 (N_9413,N_9215,N_9379);
and U9414 (N_9414,N_9359,N_9322);
and U9415 (N_9415,N_9280,N_9302);
xnor U9416 (N_9416,N_9277,N_9253);
xor U9417 (N_9417,N_9393,N_9240);
xor U9418 (N_9418,N_9229,N_9305);
nand U9419 (N_9419,N_9341,N_9368);
xnor U9420 (N_9420,N_9246,N_9385);
or U9421 (N_9421,N_9377,N_9252);
xnor U9422 (N_9422,N_9324,N_9363);
nor U9423 (N_9423,N_9315,N_9353);
xor U9424 (N_9424,N_9225,N_9260);
nand U9425 (N_9425,N_9294,N_9394);
and U9426 (N_9426,N_9356,N_9321);
nor U9427 (N_9427,N_9237,N_9210);
nor U9428 (N_9428,N_9222,N_9398);
nor U9429 (N_9429,N_9275,N_9238);
or U9430 (N_9430,N_9329,N_9248);
nor U9431 (N_9431,N_9297,N_9370);
or U9432 (N_9432,N_9211,N_9366);
nor U9433 (N_9433,N_9290,N_9317);
xor U9434 (N_9434,N_9261,N_9310);
xor U9435 (N_9435,N_9219,N_9247);
nand U9436 (N_9436,N_9267,N_9373);
and U9437 (N_9437,N_9235,N_9397);
nand U9438 (N_9438,N_9258,N_9284);
or U9439 (N_9439,N_9296,N_9372);
nor U9440 (N_9440,N_9395,N_9250);
and U9441 (N_9441,N_9311,N_9388);
and U9442 (N_9442,N_9245,N_9342);
and U9443 (N_9443,N_9304,N_9241);
or U9444 (N_9444,N_9291,N_9399);
and U9445 (N_9445,N_9282,N_9251);
and U9446 (N_9446,N_9216,N_9278);
nor U9447 (N_9447,N_9365,N_9357);
nor U9448 (N_9448,N_9257,N_9262);
nand U9449 (N_9449,N_9214,N_9391);
or U9450 (N_9450,N_9345,N_9354);
or U9451 (N_9451,N_9333,N_9348);
xnor U9452 (N_9452,N_9332,N_9319);
nor U9453 (N_9453,N_9364,N_9306);
nand U9454 (N_9454,N_9346,N_9328);
nor U9455 (N_9455,N_9334,N_9283);
or U9456 (N_9456,N_9371,N_9323);
nand U9457 (N_9457,N_9361,N_9380);
nor U9458 (N_9458,N_9369,N_9307);
nand U9459 (N_9459,N_9281,N_9360);
nor U9460 (N_9460,N_9220,N_9200);
xnor U9461 (N_9461,N_9344,N_9352);
or U9462 (N_9462,N_9271,N_9227);
nor U9463 (N_9463,N_9203,N_9209);
nand U9464 (N_9464,N_9347,N_9374);
xnor U9465 (N_9465,N_9213,N_9263);
nor U9466 (N_9466,N_9288,N_9218);
xnor U9467 (N_9467,N_9202,N_9206);
nor U9468 (N_9468,N_9201,N_9335);
xnor U9469 (N_9469,N_9336,N_9318);
and U9470 (N_9470,N_9221,N_9349);
xnor U9471 (N_9471,N_9383,N_9254);
nand U9472 (N_9472,N_9293,N_9249);
or U9473 (N_9473,N_9327,N_9309);
nand U9474 (N_9474,N_9243,N_9376);
nand U9475 (N_9475,N_9265,N_9355);
and U9476 (N_9476,N_9340,N_9337);
nor U9477 (N_9477,N_9208,N_9313);
or U9478 (N_9478,N_9303,N_9292);
xnor U9479 (N_9479,N_9266,N_9259);
nor U9480 (N_9480,N_9236,N_9285);
nor U9481 (N_9481,N_9207,N_9276);
nor U9482 (N_9482,N_9350,N_9230);
nor U9483 (N_9483,N_9270,N_9204);
nand U9484 (N_9484,N_9343,N_9234);
xnor U9485 (N_9485,N_9326,N_9287);
nand U9486 (N_9486,N_9299,N_9264);
nor U9487 (N_9487,N_9392,N_9396);
xnor U9488 (N_9488,N_9244,N_9320);
nor U9489 (N_9489,N_9256,N_9268);
and U9490 (N_9490,N_9223,N_9242);
or U9491 (N_9491,N_9217,N_9255);
xnor U9492 (N_9492,N_9375,N_9300);
nor U9493 (N_9493,N_9301,N_9339);
xnor U9494 (N_9494,N_9231,N_9390);
nor U9495 (N_9495,N_9224,N_9382);
xor U9496 (N_9496,N_9387,N_9331);
nor U9497 (N_9497,N_9295,N_9384);
or U9498 (N_9498,N_9358,N_9362);
or U9499 (N_9499,N_9386,N_9389);
nor U9500 (N_9500,N_9240,N_9392);
and U9501 (N_9501,N_9324,N_9251);
nor U9502 (N_9502,N_9321,N_9337);
xor U9503 (N_9503,N_9270,N_9350);
and U9504 (N_9504,N_9215,N_9395);
or U9505 (N_9505,N_9215,N_9323);
or U9506 (N_9506,N_9246,N_9221);
xnor U9507 (N_9507,N_9278,N_9283);
xor U9508 (N_9508,N_9276,N_9397);
xor U9509 (N_9509,N_9253,N_9293);
xnor U9510 (N_9510,N_9389,N_9215);
and U9511 (N_9511,N_9311,N_9229);
xor U9512 (N_9512,N_9321,N_9390);
and U9513 (N_9513,N_9290,N_9334);
or U9514 (N_9514,N_9334,N_9282);
nor U9515 (N_9515,N_9322,N_9284);
or U9516 (N_9516,N_9302,N_9315);
nand U9517 (N_9517,N_9291,N_9374);
xnor U9518 (N_9518,N_9268,N_9314);
and U9519 (N_9519,N_9235,N_9381);
nand U9520 (N_9520,N_9366,N_9393);
xnor U9521 (N_9521,N_9363,N_9399);
nor U9522 (N_9522,N_9262,N_9377);
and U9523 (N_9523,N_9276,N_9360);
nand U9524 (N_9524,N_9239,N_9358);
xor U9525 (N_9525,N_9383,N_9306);
nand U9526 (N_9526,N_9321,N_9372);
nand U9527 (N_9527,N_9345,N_9219);
nor U9528 (N_9528,N_9320,N_9375);
nor U9529 (N_9529,N_9353,N_9283);
xor U9530 (N_9530,N_9361,N_9210);
and U9531 (N_9531,N_9390,N_9256);
xor U9532 (N_9532,N_9388,N_9219);
xor U9533 (N_9533,N_9214,N_9273);
xor U9534 (N_9534,N_9333,N_9384);
nor U9535 (N_9535,N_9264,N_9306);
and U9536 (N_9536,N_9339,N_9318);
and U9537 (N_9537,N_9296,N_9228);
nor U9538 (N_9538,N_9205,N_9312);
xor U9539 (N_9539,N_9290,N_9339);
and U9540 (N_9540,N_9369,N_9335);
and U9541 (N_9541,N_9314,N_9264);
and U9542 (N_9542,N_9332,N_9222);
nand U9543 (N_9543,N_9389,N_9397);
xor U9544 (N_9544,N_9328,N_9209);
or U9545 (N_9545,N_9386,N_9221);
and U9546 (N_9546,N_9270,N_9342);
and U9547 (N_9547,N_9209,N_9254);
and U9548 (N_9548,N_9365,N_9349);
and U9549 (N_9549,N_9343,N_9227);
or U9550 (N_9550,N_9332,N_9367);
nand U9551 (N_9551,N_9295,N_9342);
nor U9552 (N_9552,N_9201,N_9325);
and U9553 (N_9553,N_9334,N_9348);
nand U9554 (N_9554,N_9258,N_9288);
and U9555 (N_9555,N_9290,N_9374);
or U9556 (N_9556,N_9279,N_9257);
nand U9557 (N_9557,N_9253,N_9329);
nor U9558 (N_9558,N_9245,N_9259);
and U9559 (N_9559,N_9218,N_9302);
xor U9560 (N_9560,N_9268,N_9387);
nand U9561 (N_9561,N_9370,N_9265);
xor U9562 (N_9562,N_9341,N_9322);
nor U9563 (N_9563,N_9211,N_9288);
nor U9564 (N_9564,N_9222,N_9243);
xnor U9565 (N_9565,N_9381,N_9305);
and U9566 (N_9566,N_9245,N_9388);
and U9567 (N_9567,N_9232,N_9282);
nand U9568 (N_9568,N_9335,N_9266);
nand U9569 (N_9569,N_9383,N_9381);
nand U9570 (N_9570,N_9213,N_9218);
nor U9571 (N_9571,N_9224,N_9346);
nand U9572 (N_9572,N_9264,N_9262);
xor U9573 (N_9573,N_9209,N_9287);
xor U9574 (N_9574,N_9211,N_9337);
and U9575 (N_9575,N_9364,N_9348);
and U9576 (N_9576,N_9356,N_9367);
nand U9577 (N_9577,N_9331,N_9382);
nor U9578 (N_9578,N_9200,N_9323);
and U9579 (N_9579,N_9322,N_9204);
or U9580 (N_9580,N_9288,N_9351);
and U9581 (N_9581,N_9216,N_9369);
or U9582 (N_9582,N_9249,N_9238);
or U9583 (N_9583,N_9251,N_9231);
or U9584 (N_9584,N_9289,N_9250);
and U9585 (N_9585,N_9297,N_9292);
or U9586 (N_9586,N_9327,N_9265);
nor U9587 (N_9587,N_9329,N_9299);
xor U9588 (N_9588,N_9205,N_9242);
or U9589 (N_9589,N_9280,N_9290);
and U9590 (N_9590,N_9335,N_9331);
and U9591 (N_9591,N_9205,N_9360);
and U9592 (N_9592,N_9387,N_9374);
or U9593 (N_9593,N_9330,N_9311);
or U9594 (N_9594,N_9238,N_9301);
xnor U9595 (N_9595,N_9358,N_9202);
or U9596 (N_9596,N_9243,N_9307);
or U9597 (N_9597,N_9275,N_9382);
and U9598 (N_9598,N_9292,N_9228);
and U9599 (N_9599,N_9373,N_9228);
nor U9600 (N_9600,N_9483,N_9551);
and U9601 (N_9601,N_9432,N_9412);
xnor U9602 (N_9602,N_9542,N_9478);
and U9603 (N_9603,N_9490,N_9586);
nor U9604 (N_9604,N_9489,N_9539);
xor U9605 (N_9605,N_9596,N_9544);
xor U9606 (N_9606,N_9552,N_9429);
xor U9607 (N_9607,N_9431,N_9567);
nand U9608 (N_9608,N_9435,N_9532);
nor U9609 (N_9609,N_9529,N_9500);
nor U9610 (N_9610,N_9447,N_9506);
or U9611 (N_9611,N_9495,N_9585);
nor U9612 (N_9612,N_9442,N_9418);
or U9613 (N_9613,N_9592,N_9556);
or U9614 (N_9614,N_9501,N_9488);
xnor U9615 (N_9615,N_9548,N_9494);
nor U9616 (N_9616,N_9424,N_9496);
and U9617 (N_9617,N_9474,N_9599);
nand U9618 (N_9618,N_9512,N_9545);
and U9619 (N_9619,N_9504,N_9470);
or U9620 (N_9620,N_9425,N_9519);
or U9621 (N_9621,N_9491,N_9427);
nor U9622 (N_9622,N_9402,N_9514);
or U9623 (N_9623,N_9463,N_9400);
xnor U9624 (N_9624,N_9466,N_9449);
or U9625 (N_9625,N_9428,N_9517);
nor U9626 (N_9626,N_9538,N_9420);
nor U9627 (N_9627,N_9575,N_9485);
xor U9628 (N_9628,N_9439,N_9422);
nand U9629 (N_9629,N_9595,N_9597);
xnor U9630 (N_9630,N_9508,N_9405);
nand U9631 (N_9631,N_9593,N_9416);
nor U9632 (N_9632,N_9453,N_9587);
or U9633 (N_9633,N_9481,N_9577);
xnor U9634 (N_9634,N_9456,N_9584);
nor U9635 (N_9635,N_9445,N_9473);
and U9636 (N_9636,N_9594,N_9476);
and U9637 (N_9637,N_9580,N_9417);
or U9638 (N_9638,N_9541,N_9415);
and U9639 (N_9639,N_9461,N_9434);
nor U9640 (N_9640,N_9547,N_9446);
and U9641 (N_9641,N_9563,N_9492);
or U9642 (N_9642,N_9515,N_9540);
or U9643 (N_9643,N_9468,N_9465);
xnor U9644 (N_9644,N_9559,N_9458);
and U9645 (N_9645,N_9561,N_9406);
and U9646 (N_9646,N_9497,N_9480);
nor U9647 (N_9647,N_9578,N_9413);
nand U9648 (N_9648,N_9414,N_9507);
xnor U9649 (N_9649,N_9457,N_9404);
and U9650 (N_9650,N_9516,N_9471);
and U9651 (N_9651,N_9591,N_9460);
xnor U9652 (N_9652,N_9576,N_9581);
nand U9653 (N_9653,N_9523,N_9467);
and U9654 (N_9654,N_9564,N_9430);
xor U9655 (N_9655,N_9574,N_9569);
and U9656 (N_9656,N_9536,N_9543);
xnor U9657 (N_9657,N_9423,N_9560);
or U9658 (N_9658,N_9568,N_9499);
xor U9659 (N_9659,N_9444,N_9503);
nor U9660 (N_9660,N_9472,N_9451);
xor U9661 (N_9661,N_9498,N_9419);
nor U9662 (N_9662,N_9572,N_9403);
nand U9663 (N_9663,N_9486,N_9450);
or U9664 (N_9664,N_9550,N_9479);
nor U9665 (N_9665,N_9558,N_9493);
and U9666 (N_9666,N_9452,N_9527);
nand U9667 (N_9667,N_9462,N_9553);
or U9668 (N_9668,N_9583,N_9421);
nor U9669 (N_9669,N_9436,N_9510);
xor U9670 (N_9670,N_9518,N_9571);
nand U9671 (N_9671,N_9440,N_9573);
xnor U9672 (N_9672,N_9531,N_9566);
and U9673 (N_9673,N_9554,N_9570);
and U9674 (N_9674,N_9509,N_9408);
and U9675 (N_9675,N_9528,N_9505);
nand U9676 (N_9676,N_9590,N_9433);
nand U9677 (N_9677,N_9526,N_9459);
nor U9678 (N_9678,N_9555,N_9546);
xor U9679 (N_9679,N_9582,N_9562);
or U9680 (N_9680,N_9533,N_9521);
nor U9681 (N_9681,N_9438,N_9589);
or U9682 (N_9682,N_9410,N_9535);
or U9683 (N_9683,N_9475,N_9565);
nor U9684 (N_9684,N_9522,N_9524);
nor U9685 (N_9685,N_9448,N_9525);
xor U9686 (N_9686,N_9464,N_9534);
nor U9687 (N_9687,N_9588,N_9537);
nand U9688 (N_9688,N_9426,N_9484);
or U9689 (N_9689,N_9437,N_9598);
nand U9690 (N_9690,N_9454,N_9513);
nand U9691 (N_9691,N_9549,N_9409);
nand U9692 (N_9692,N_9455,N_9407);
xnor U9693 (N_9693,N_9530,N_9477);
nor U9694 (N_9694,N_9401,N_9469);
xnor U9695 (N_9695,N_9511,N_9411);
xor U9696 (N_9696,N_9487,N_9557);
xnor U9697 (N_9697,N_9441,N_9579);
nand U9698 (N_9698,N_9482,N_9502);
and U9699 (N_9699,N_9443,N_9520);
xnor U9700 (N_9700,N_9446,N_9567);
or U9701 (N_9701,N_9545,N_9487);
xor U9702 (N_9702,N_9484,N_9413);
or U9703 (N_9703,N_9447,N_9429);
xnor U9704 (N_9704,N_9500,N_9554);
or U9705 (N_9705,N_9560,N_9471);
or U9706 (N_9706,N_9446,N_9545);
nand U9707 (N_9707,N_9517,N_9498);
nor U9708 (N_9708,N_9531,N_9499);
or U9709 (N_9709,N_9402,N_9523);
or U9710 (N_9710,N_9536,N_9459);
and U9711 (N_9711,N_9405,N_9571);
or U9712 (N_9712,N_9403,N_9436);
and U9713 (N_9713,N_9441,N_9560);
nand U9714 (N_9714,N_9500,N_9432);
or U9715 (N_9715,N_9540,N_9439);
or U9716 (N_9716,N_9400,N_9418);
nor U9717 (N_9717,N_9468,N_9413);
and U9718 (N_9718,N_9406,N_9492);
and U9719 (N_9719,N_9580,N_9575);
nand U9720 (N_9720,N_9570,N_9413);
nand U9721 (N_9721,N_9430,N_9416);
nor U9722 (N_9722,N_9517,N_9487);
nand U9723 (N_9723,N_9443,N_9545);
and U9724 (N_9724,N_9494,N_9454);
and U9725 (N_9725,N_9547,N_9523);
nor U9726 (N_9726,N_9446,N_9570);
nor U9727 (N_9727,N_9413,N_9404);
nor U9728 (N_9728,N_9549,N_9462);
and U9729 (N_9729,N_9593,N_9420);
xnor U9730 (N_9730,N_9518,N_9572);
xnor U9731 (N_9731,N_9548,N_9551);
xnor U9732 (N_9732,N_9537,N_9470);
xnor U9733 (N_9733,N_9439,N_9427);
nor U9734 (N_9734,N_9553,N_9443);
nand U9735 (N_9735,N_9496,N_9455);
and U9736 (N_9736,N_9415,N_9414);
nand U9737 (N_9737,N_9524,N_9564);
xnor U9738 (N_9738,N_9522,N_9483);
nor U9739 (N_9739,N_9512,N_9428);
nand U9740 (N_9740,N_9550,N_9456);
nand U9741 (N_9741,N_9545,N_9499);
nand U9742 (N_9742,N_9508,N_9579);
nand U9743 (N_9743,N_9434,N_9426);
nor U9744 (N_9744,N_9483,N_9508);
xnor U9745 (N_9745,N_9478,N_9422);
nand U9746 (N_9746,N_9412,N_9498);
xnor U9747 (N_9747,N_9499,N_9470);
xor U9748 (N_9748,N_9424,N_9567);
nand U9749 (N_9749,N_9481,N_9467);
xnor U9750 (N_9750,N_9565,N_9522);
and U9751 (N_9751,N_9557,N_9451);
and U9752 (N_9752,N_9435,N_9512);
nand U9753 (N_9753,N_9547,N_9525);
xor U9754 (N_9754,N_9463,N_9492);
nand U9755 (N_9755,N_9537,N_9462);
nor U9756 (N_9756,N_9472,N_9545);
nand U9757 (N_9757,N_9462,N_9496);
xnor U9758 (N_9758,N_9415,N_9462);
or U9759 (N_9759,N_9511,N_9485);
and U9760 (N_9760,N_9453,N_9591);
xnor U9761 (N_9761,N_9587,N_9566);
nand U9762 (N_9762,N_9572,N_9552);
nand U9763 (N_9763,N_9572,N_9488);
nor U9764 (N_9764,N_9587,N_9530);
nand U9765 (N_9765,N_9451,N_9485);
nand U9766 (N_9766,N_9431,N_9536);
nand U9767 (N_9767,N_9440,N_9418);
nor U9768 (N_9768,N_9586,N_9421);
and U9769 (N_9769,N_9543,N_9465);
or U9770 (N_9770,N_9589,N_9428);
and U9771 (N_9771,N_9561,N_9490);
and U9772 (N_9772,N_9596,N_9558);
and U9773 (N_9773,N_9513,N_9595);
nand U9774 (N_9774,N_9467,N_9486);
nand U9775 (N_9775,N_9503,N_9501);
xor U9776 (N_9776,N_9478,N_9585);
and U9777 (N_9777,N_9574,N_9458);
nor U9778 (N_9778,N_9545,N_9523);
and U9779 (N_9779,N_9556,N_9459);
xnor U9780 (N_9780,N_9462,N_9460);
and U9781 (N_9781,N_9499,N_9436);
nor U9782 (N_9782,N_9459,N_9572);
nor U9783 (N_9783,N_9550,N_9571);
nand U9784 (N_9784,N_9535,N_9462);
nor U9785 (N_9785,N_9442,N_9544);
nand U9786 (N_9786,N_9570,N_9400);
and U9787 (N_9787,N_9552,N_9419);
nand U9788 (N_9788,N_9489,N_9461);
nand U9789 (N_9789,N_9468,N_9490);
or U9790 (N_9790,N_9412,N_9468);
or U9791 (N_9791,N_9441,N_9450);
or U9792 (N_9792,N_9515,N_9575);
nor U9793 (N_9793,N_9492,N_9405);
and U9794 (N_9794,N_9479,N_9566);
xnor U9795 (N_9795,N_9443,N_9462);
or U9796 (N_9796,N_9440,N_9587);
nand U9797 (N_9797,N_9590,N_9538);
nand U9798 (N_9798,N_9532,N_9440);
or U9799 (N_9799,N_9466,N_9589);
xnor U9800 (N_9800,N_9767,N_9720);
nor U9801 (N_9801,N_9619,N_9650);
nand U9802 (N_9802,N_9693,N_9746);
xor U9803 (N_9803,N_9731,N_9612);
xnor U9804 (N_9804,N_9714,N_9761);
or U9805 (N_9805,N_9604,N_9637);
and U9806 (N_9806,N_9797,N_9705);
and U9807 (N_9807,N_9671,N_9739);
or U9808 (N_9808,N_9744,N_9799);
xor U9809 (N_9809,N_9747,N_9796);
and U9810 (N_9810,N_9707,N_9770);
xnor U9811 (N_9811,N_9755,N_9723);
and U9812 (N_9812,N_9732,N_9643);
or U9813 (N_9813,N_9751,N_9765);
nand U9814 (N_9814,N_9678,N_9789);
or U9815 (N_9815,N_9614,N_9759);
nor U9816 (N_9816,N_9780,N_9683);
xnor U9817 (N_9817,N_9657,N_9795);
and U9818 (N_9818,N_9631,N_9729);
nor U9819 (N_9819,N_9745,N_9769);
nor U9820 (N_9820,N_9613,N_9749);
nand U9821 (N_9821,N_9622,N_9697);
xor U9822 (N_9822,N_9728,N_9708);
nor U9823 (N_9823,N_9783,N_9641);
nor U9824 (N_9824,N_9764,N_9758);
xor U9825 (N_9825,N_9648,N_9609);
and U9826 (N_9826,N_9735,N_9675);
nor U9827 (N_9827,N_9768,N_9689);
nor U9828 (N_9828,N_9711,N_9667);
nor U9829 (N_9829,N_9670,N_9696);
nor U9830 (N_9830,N_9709,N_9702);
or U9831 (N_9831,N_9794,N_9607);
nor U9832 (N_9832,N_9793,N_9791);
nand U9833 (N_9833,N_9659,N_9685);
nor U9834 (N_9834,N_9664,N_9647);
and U9835 (N_9835,N_9725,N_9640);
or U9836 (N_9836,N_9632,N_9730);
or U9837 (N_9837,N_9651,N_9782);
or U9838 (N_9838,N_9762,N_9716);
nor U9839 (N_9839,N_9736,N_9676);
xor U9840 (N_9840,N_9602,N_9628);
or U9841 (N_9841,N_9771,N_9621);
nand U9842 (N_9842,N_9649,N_9691);
or U9843 (N_9843,N_9625,N_9772);
xor U9844 (N_9844,N_9753,N_9653);
xor U9845 (N_9845,N_9715,N_9630);
nand U9846 (N_9846,N_9655,N_9668);
or U9847 (N_9847,N_9710,N_9712);
xor U9848 (N_9848,N_9665,N_9741);
nor U9849 (N_9849,N_9658,N_9713);
nor U9850 (N_9850,N_9600,N_9666);
and U9851 (N_9851,N_9626,N_9788);
nor U9852 (N_9852,N_9692,N_9679);
and U9853 (N_9853,N_9617,N_9686);
nand U9854 (N_9854,N_9760,N_9662);
and U9855 (N_9855,N_9724,N_9790);
xnor U9856 (N_9856,N_9669,N_9606);
or U9857 (N_9857,N_9611,N_9784);
or U9858 (N_9858,N_9719,N_9726);
or U9859 (N_9859,N_9656,N_9639);
xnor U9860 (N_9860,N_9703,N_9785);
and U9861 (N_9861,N_9698,N_9774);
or U9862 (N_9862,N_9636,N_9798);
nor U9863 (N_9863,N_9734,N_9629);
and U9864 (N_9864,N_9700,N_9766);
xnor U9865 (N_9865,N_9627,N_9684);
nor U9866 (N_9866,N_9695,N_9633);
or U9867 (N_9867,N_9740,N_9763);
xnor U9868 (N_9868,N_9661,N_9756);
nand U9869 (N_9869,N_9638,N_9687);
xor U9870 (N_9870,N_9601,N_9603);
and U9871 (N_9871,N_9660,N_9645);
nand U9872 (N_9872,N_9717,N_9681);
or U9873 (N_9873,N_9786,N_9738);
and U9874 (N_9874,N_9750,N_9605);
or U9875 (N_9875,N_9642,N_9616);
nor U9876 (N_9876,N_9704,N_9754);
nand U9877 (N_9877,N_9701,N_9654);
nand U9878 (N_9878,N_9677,N_9674);
nand U9879 (N_9879,N_9644,N_9776);
nand U9880 (N_9880,N_9682,N_9742);
xor U9881 (N_9881,N_9663,N_9680);
nor U9882 (N_9882,N_9775,N_9623);
nor U9883 (N_9883,N_9620,N_9792);
nand U9884 (N_9884,N_9652,N_9748);
and U9885 (N_9885,N_9781,N_9646);
nand U9886 (N_9886,N_9624,N_9699);
xnor U9887 (N_9887,N_9635,N_9727);
xnor U9888 (N_9888,N_9690,N_9706);
xor U9889 (N_9889,N_9722,N_9787);
xor U9890 (N_9890,N_9779,N_9694);
xnor U9891 (N_9891,N_9721,N_9757);
xnor U9892 (N_9892,N_9718,N_9752);
nor U9893 (N_9893,N_9673,N_9733);
nor U9894 (N_9894,N_9743,N_9608);
xnor U9895 (N_9895,N_9615,N_9610);
xnor U9896 (N_9896,N_9777,N_9773);
nor U9897 (N_9897,N_9688,N_9737);
nor U9898 (N_9898,N_9672,N_9618);
and U9899 (N_9899,N_9634,N_9778);
nand U9900 (N_9900,N_9600,N_9695);
nor U9901 (N_9901,N_9764,N_9777);
nor U9902 (N_9902,N_9682,N_9790);
or U9903 (N_9903,N_9641,N_9619);
nor U9904 (N_9904,N_9626,N_9698);
xor U9905 (N_9905,N_9749,N_9617);
nand U9906 (N_9906,N_9685,N_9673);
and U9907 (N_9907,N_9631,N_9769);
and U9908 (N_9908,N_9715,N_9605);
nor U9909 (N_9909,N_9694,N_9664);
nor U9910 (N_9910,N_9679,N_9739);
or U9911 (N_9911,N_9787,N_9721);
and U9912 (N_9912,N_9739,N_9600);
xor U9913 (N_9913,N_9623,N_9724);
or U9914 (N_9914,N_9730,N_9665);
or U9915 (N_9915,N_9734,N_9658);
nor U9916 (N_9916,N_9774,N_9687);
or U9917 (N_9917,N_9792,N_9621);
xnor U9918 (N_9918,N_9705,N_9703);
nand U9919 (N_9919,N_9637,N_9618);
nor U9920 (N_9920,N_9619,N_9697);
nand U9921 (N_9921,N_9732,N_9620);
nor U9922 (N_9922,N_9696,N_9647);
xnor U9923 (N_9923,N_9795,N_9687);
and U9924 (N_9924,N_9676,N_9602);
nor U9925 (N_9925,N_9659,N_9646);
or U9926 (N_9926,N_9749,N_9748);
nor U9927 (N_9927,N_9756,N_9702);
xnor U9928 (N_9928,N_9762,N_9677);
nand U9929 (N_9929,N_9767,N_9610);
xnor U9930 (N_9930,N_9726,N_9785);
nor U9931 (N_9931,N_9614,N_9798);
or U9932 (N_9932,N_9627,N_9650);
or U9933 (N_9933,N_9733,N_9622);
nand U9934 (N_9934,N_9672,N_9738);
or U9935 (N_9935,N_9776,N_9740);
xor U9936 (N_9936,N_9638,N_9660);
nand U9937 (N_9937,N_9781,N_9670);
nor U9938 (N_9938,N_9708,N_9656);
or U9939 (N_9939,N_9628,N_9770);
xor U9940 (N_9940,N_9759,N_9702);
and U9941 (N_9941,N_9736,N_9776);
and U9942 (N_9942,N_9795,N_9621);
xor U9943 (N_9943,N_9768,N_9711);
nor U9944 (N_9944,N_9730,N_9742);
nand U9945 (N_9945,N_9719,N_9702);
and U9946 (N_9946,N_9773,N_9648);
or U9947 (N_9947,N_9637,N_9641);
or U9948 (N_9948,N_9713,N_9785);
and U9949 (N_9949,N_9619,N_9704);
nand U9950 (N_9950,N_9651,N_9637);
and U9951 (N_9951,N_9783,N_9700);
nand U9952 (N_9952,N_9662,N_9637);
xnor U9953 (N_9953,N_9635,N_9682);
and U9954 (N_9954,N_9616,N_9747);
or U9955 (N_9955,N_9736,N_9612);
nor U9956 (N_9956,N_9656,N_9741);
nor U9957 (N_9957,N_9680,N_9616);
nor U9958 (N_9958,N_9736,N_9741);
xor U9959 (N_9959,N_9684,N_9685);
xnor U9960 (N_9960,N_9797,N_9608);
nand U9961 (N_9961,N_9746,N_9601);
nor U9962 (N_9962,N_9602,N_9687);
and U9963 (N_9963,N_9735,N_9610);
nor U9964 (N_9964,N_9770,N_9754);
xor U9965 (N_9965,N_9746,N_9779);
xor U9966 (N_9966,N_9788,N_9620);
nand U9967 (N_9967,N_9766,N_9774);
nor U9968 (N_9968,N_9705,N_9794);
nor U9969 (N_9969,N_9784,N_9632);
xnor U9970 (N_9970,N_9672,N_9774);
nand U9971 (N_9971,N_9668,N_9751);
nor U9972 (N_9972,N_9676,N_9686);
nand U9973 (N_9973,N_9756,N_9626);
or U9974 (N_9974,N_9674,N_9624);
and U9975 (N_9975,N_9717,N_9680);
nor U9976 (N_9976,N_9639,N_9710);
nand U9977 (N_9977,N_9725,N_9721);
and U9978 (N_9978,N_9678,N_9773);
xor U9979 (N_9979,N_9695,N_9678);
or U9980 (N_9980,N_9783,N_9624);
or U9981 (N_9981,N_9650,N_9714);
and U9982 (N_9982,N_9701,N_9638);
or U9983 (N_9983,N_9639,N_9766);
or U9984 (N_9984,N_9664,N_9751);
or U9985 (N_9985,N_9735,N_9769);
and U9986 (N_9986,N_9758,N_9714);
nor U9987 (N_9987,N_9611,N_9662);
xnor U9988 (N_9988,N_9789,N_9774);
nor U9989 (N_9989,N_9619,N_9780);
xnor U9990 (N_9990,N_9617,N_9708);
nor U9991 (N_9991,N_9759,N_9766);
nor U9992 (N_9992,N_9714,N_9743);
or U9993 (N_9993,N_9746,N_9664);
and U9994 (N_9994,N_9616,N_9649);
nor U9995 (N_9995,N_9721,N_9755);
or U9996 (N_9996,N_9726,N_9661);
or U9997 (N_9997,N_9768,N_9766);
xnor U9998 (N_9998,N_9781,N_9707);
or U9999 (N_9999,N_9759,N_9756);
and U10000 (N_10000,N_9890,N_9806);
nand U10001 (N_10001,N_9830,N_9978);
nand U10002 (N_10002,N_9996,N_9828);
and U10003 (N_10003,N_9993,N_9907);
nor U10004 (N_10004,N_9833,N_9955);
and U10005 (N_10005,N_9898,N_9886);
or U10006 (N_10006,N_9903,N_9845);
and U10007 (N_10007,N_9933,N_9877);
or U10008 (N_10008,N_9817,N_9910);
or U10009 (N_10009,N_9867,N_9836);
xnor U10010 (N_10010,N_9965,N_9875);
and U10011 (N_10011,N_9974,N_9994);
nand U10012 (N_10012,N_9827,N_9963);
or U10013 (N_10013,N_9949,N_9872);
nor U10014 (N_10014,N_9863,N_9945);
and U10015 (N_10015,N_9834,N_9981);
and U10016 (N_10016,N_9913,N_9970);
or U10017 (N_10017,N_9900,N_9813);
nor U10018 (N_10018,N_9849,N_9892);
xor U10019 (N_10019,N_9995,N_9987);
xor U10020 (N_10020,N_9921,N_9808);
nand U10021 (N_10021,N_9878,N_9825);
nor U10022 (N_10022,N_9804,N_9810);
or U10023 (N_10023,N_9893,N_9926);
or U10024 (N_10024,N_9811,N_9944);
and U10025 (N_10025,N_9835,N_9881);
or U10026 (N_10026,N_9832,N_9909);
nand U10027 (N_10027,N_9858,N_9820);
xnor U10028 (N_10028,N_9936,N_9873);
nand U10029 (N_10029,N_9826,N_9988);
xnor U10030 (N_10030,N_9906,N_9896);
nand U10031 (N_10031,N_9976,N_9853);
nor U10032 (N_10032,N_9989,N_9807);
nor U10033 (N_10033,N_9865,N_9980);
and U10034 (N_10034,N_9862,N_9802);
nand U10035 (N_10035,N_9948,N_9962);
xnor U10036 (N_10036,N_9971,N_9801);
and U10037 (N_10037,N_9837,N_9895);
and U10038 (N_10038,N_9992,N_9956);
nor U10039 (N_10039,N_9957,N_9883);
nor U10040 (N_10040,N_9928,N_9940);
or U10041 (N_10041,N_9983,N_9979);
and U10042 (N_10042,N_9879,N_9904);
or U10043 (N_10043,N_9916,N_9998);
nand U10044 (N_10044,N_9953,N_9943);
xor U10045 (N_10045,N_9931,N_9800);
and U10046 (N_10046,N_9860,N_9973);
or U10047 (N_10047,N_9990,N_9871);
nand U10048 (N_10048,N_9961,N_9999);
nor U10049 (N_10049,N_9888,N_9821);
or U10050 (N_10050,N_9912,N_9809);
or U10051 (N_10051,N_9869,N_9950);
nand U10052 (N_10052,N_9920,N_9805);
or U10053 (N_10053,N_9816,N_9841);
or U10054 (N_10054,N_9831,N_9942);
nand U10055 (N_10055,N_9847,N_9818);
nor U10056 (N_10056,N_9925,N_9911);
or U10057 (N_10057,N_9991,N_9859);
or U10058 (N_10058,N_9864,N_9885);
and U10059 (N_10059,N_9952,N_9848);
nand U10060 (N_10060,N_9824,N_9838);
nor U10061 (N_10061,N_9856,N_9897);
and U10062 (N_10062,N_9922,N_9964);
nand U10063 (N_10063,N_9803,N_9814);
or U10064 (N_10064,N_9839,N_9972);
nor U10065 (N_10065,N_9946,N_9868);
or U10066 (N_10066,N_9889,N_9919);
nor U10067 (N_10067,N_9894,N_9924);
and U10068 (N_10068,N_9959,N_9908);
and U10069 (N_10069,N_9861,N_9882);
or U10070 (N_10070,N_9941,N_9899);
and U10071 (N_10071,N_9823,N_9984);
xor U10072 (N_10072,N_9901,N_9935);
nand U10073 (N_10073,N_9937,N_9854);
nand U10074 (N_10074,N_9915,N_9954);
nor U10075 (N_10075,N_9930,N_9874);
nor U10076 (N_10076,N_9884,N_9812);
and U10077 (N_10077,N_9917,N_9844);
nor U10078 (N_10078,N_9932,N_9985);
xnor U10079 (N_10079,N_9967,N_9843);
nand U10080 (N_10080,N_9966,N_9829);
or U10081 (N_10081,N_9947,N_9902);
and U10082 (N_10082,N_9986,N_9997);
nand U10083 (N_10083,N_9977,N_9929);
and U10084 (N_10084,N_9958,N_9934);
nand U10085 (N_10085,N_9846,N_9850);
xnor U10086 (N_10086,N_9960,N_9923);
xor U10087 (N_10087,N_9887,N_9927);
or U10088 (N_10088,N_9968,N_9982);
xor U10089 (N_10089,N_9938,N_9891);
or U10090 (N_10090,N_9905,N_9840);
nand U10091 (N_10091,N_9918,N_9857);
or U10092 (N_10092,N_9851,N_9819);
and U10093 (N_10093,N_9822,N_9870);
nand U10094 (N_10094,N_9969,N_9914);
nor U10095 (N_10095,N_9951,N_9842);
or U10096 (N_10096,N_9866,N_9876);
nor U10097 (N_10097,N_9880,N_9975);
nand U10098 (N_10098,N_9855,N_9852);
or U10099 (N_10099,N_9815,N_9939);
and U10100 (N_10100,N_9875,N_9969);
or U10101 (N_10101,N_9827,N_9940);
and U10102 (N_10102,N_9951,N_9855);
xor U10103 (N_10103,N_9940,N_9866);
and U10104 (N_10104,N_9925,N_9953);
or U10105 (N_10105,N_9919,N_9850);
or U10106 (N_10106,N_9948,N_9889);
xnor U10107 (N_10107,N_9895,N_9970);
nor U10108 (N_10108,N_9864,N_9830);
nor U10109 (N_10109,N_9948,N_9837);
nor U10110 (N_10110,N_9826,N_9864);
nand U10111 (N_10111,N_9850,N_9820);
and U10112 (N_10112,N_9829,N_9935);
xor U10113 (N_10113,N_9821,N_9941);
or U10114 (N_10114,N_9952,N_9808);
nor U10115 (N_10115,N_9904,N_9910);
and U10116 (N_10116,N_9933,N_9845);
nand U10117 (N_10117,N_9903,N_9948);
or U10118 (N_10118,N_9916,N_9962);
nor U10119 (N_10119,N_9957,N_9844);
nor U10120 (N_10120,N_9990,N_9897);
xnor U10121 (N_10121,N_9922,N_9960);
or U10122 (N_10122,N_9832,N_9857);
nor U10123 (N_10123,N_9967,N_9929);
or U10124 (N_10124,N_9814,N_9821);
xor U10125 (N_10125,N_9830,N_9982);
nand U10126 (N_10126,N_9985,N_9853);
nand U10127 (N_10127,N_9941,N_9933);
and U10128 (N_10128,N_9999,N_9856);
and U10129 (N_10129,N_9915,N_9964);
or U10130 (N_10130,N_9883,N_9859);
nor U10131 (N_10131,N_9986,N_9956);
nand U10132 (N_10132,N_9823,N_9982);
or U10133 (N_10133,N_9855,N_9856);
nor U10134 (N_10134,N_9835,N_9840);
or U10135 (N_10135,N_9872,N_9979);
or U10136 (N_10136,N_9891,N_9904);
or U10137 (N_10137,N_9821,N_9987);
xnor U10138 (N_10138,N_9808,N_9996);
or U10139 (N_10139,N_9960,N_9905);
nand U10140 (N_10140,N_9910,N_9869);
nand U10141 (N_10141,N_9942,N_9945);
nor U10142 (N_10142,N_9910,N_9996);
nor U10143 (N_10143,N_9818,N_9903);
xnor U10144 (N_10144,N_9973,N_9955);
and U10145 (N_10145,N_9952,N_9903);
nand U10146 (N_10146,N_9866,N_9961);
and U10147 (N_10147,N_9928,N_9898);
nor U10148 (N_10148,N_9809,N_9842);
nor U10149 (N_10149,N_9954,N_9851);
xnor U10150 (N_10150,N_9917,N_9839);
nand U10151 (N_10151,N_9885,N_9927);
nor U10152 (N_10152,N_9858,N_9955);
or U10153 (N_10153,N_9817,N_9955);
nor U10154 (N_10154,N_9999,N_9831);
nand U10155 (N_10155,N_9840,N_9958);
nor U10156 (N_10156,N_9942,N_9958);
xor U10157 (N_10157,N_9898,N_9831);
xor U10158 (N_10158,N_9943,N_9944);
nor U10159 (N_10159,N_9929,N_9909);
nor U10160 (N_10160,N_9835,N_9920);
xnor U10161 (N_10161,N_9835,N_9965);
nor U10162 (N_10162,N_9897,N_9851);
xnor U10163 (N_10163,N_9825,N_9830);
and U10164 (N_10164,N_9873,N_9953);
and U10165 (N_10165,N_9977,N_9868);
xor U10166 (N_10166,N_9975,N_9813);
nand U10167 (N_10167,N_9911,N_9946);
nor U10168 (N_10168,N_9955,N_9946);
or U10169 (N_10169,N_9853,N_9813);
or U10170 (N_10170,N_9910,N_9822);
and U10171 (N_10171,N_9882,N_9833);
and U10172 (N_10172,N_9943,N_9841);
and U10173 (N_10173,N_9822,N_9804);
or U10174 (N_10174,N_9864,N_9917);
and U10175 (N_10175,N_9923,N_9843);
xnor U10176 (N_10176,N_9964,N_9850);
and U10177 (N_10177,N_9871,N_9956);
nor U10178 (N_10178,N_9931,N_9849);
or U10179 (N_10179,N_9980,N_9867);
nand U10180 (N_10180,N_9862,N_9974);
and U10181 (N_10181,N_9982,N_9855);
and U10182 (N_10182,N_9826,N_9952);
or U10183 (N_10183,N_9837,N_9870);
or U10184 (N_10184,N_9886,N_9955);
or U10185 (N_10185,N_9852,N_9998);
xor U10186 (N_10186,N_9856,N_9823);
and U10187 (N_10187,N_9856,N_9851);
and U10188 (N_10188,N_9837,N_9842);
or U10189 (N_10189,N_9869,N_9852);
or U10190 (N_10190,N_9985,N_9837);
nand U10191 (N_10191,N_9955,N_9959);
nand U10192 (N_10192,N_9882,N_9819);
and U10193 (N_10193,N_9998,N_9877);
xor U10194 (N_10194,N_9881,N_9852);
nor U10195 (N_10195,N_9954,N_9820);
or U10196 (N_10196,N_9837,N_9914);
or U10197 (N_10197,N_9874,N_9834);
nand U10198 (N_10198,N_9853,N_9885);
or U10199 (N_10199,N_9947,N_9839);
and U10200 (N_10200,N_10001,N_10186);
or U10201 (N_10201,N_10126,N_10006);
nand U10202 (N_10202,N_10175,N_10029);
or U10203 (N_10203,N_10194,N_10061);
nand U10204 (N_10204,N_10073,N_10071);
nand U10205 (N_10205,N_10191,N_10151);
xnor U10206 (N_10206,N_10162,N_10127);
or U10207 (N_10207,N_10050,N_10051);
and U10208 (N_10208,N_10136,N_10036);
nor U10209 (N_10209,N_10097,N_10022);
nand U10210 (N_10210,N_10133,N_10172);
and U10211 (N_10211,N_10026,N_10159);
or U10212 (N_10212,N_10177,N_10105);
or U10213 (N_10213,N_10042,N_10009);
or U10214 (N_10214,N_10109,N_10081);
and U10215 (N_10215,N_10132,N_10053);
nand U10216 (N_10216,N_10016,N_10007);
nor U10217 (N_10217,N_10149,N_10135);
nor U10218 (N_10218,N_10044,N_10092);
xor U10219 (N_10219,N_10069,N_10064);
or U10220 (N_10220,N_10140,N_10005);
and U10221 (N_10221,N_10055,N_10032);
nor U10222 (N_10222,N_10020,N_10114);
nand U10223 (N_10223,N_10013,N_10146);
nand U10224 (N_10224,N_10106,N_10008);
and U10225 (N_10225,N_10028,N_10078);
or U10226 (N_10226,N_10014,N_10163);
xor U10227 (N_10227,N_10040,N_10089);
or U10228 (N_10228,N_10080,N_10104);
and U10229 (N_10229,N_10103,N_10045);
and U10230 (N_10230,N_10118,N_10077);
and U10231 (N_10231,N_10138,N_10056);
nor U10232 (N_10232,N_10184,N_10166);
or U10233 (N_10233,N_10173,N_10147);
nand U10234 (N_10234,N_10130,N_10030);
nand U10235 (N_10235,N_10068,N_10094);
xor U10236 (N_10236,N_10131,N_10119);
nor U10237 (N_10237,N_10122,N_10171);
nor U10238 (N_10238,N_10190,N_10060);
xor U10239 (N_10239,N_10164,N_10093);
nand U10240 (N_10240,N_10063,N_10052);
or U10241 (N_10241,N_10128,N_10110);
xor U10242 (N_10242,N_10012,N_10150);
or U10243 (N_10243,N_10003,N_10041);
and U10244 (N_10244,N_10199,N_10074);
or U10245 (N_10245,N_10117,N_10141);
xnor U10246 (N_10246,N_10098,N_10174);
and U10247 (N_10247,N_10048,N_10062);
nand U10248 (N_10248,N_10099,N_10185);
nor U10249 (N_10249,N_10176,N_10155);
xnor U10250 (N_10250,N_10083,N_10082);
xnor U10251 (N_10251,N_10156,N_10058);
and U10252 (N_10252,N_10115,N_10129);
nand U10253 (N_10253,N_10154,N_10066);
xnor U10254 (N_10254,N_10102,N_10086);
and U10255 (N_10255,N_10000,N_10160);
or U10256 (N_10256,N_10027,N_10090);
nand U10257 (N_10257,N_10017,N_10076);
and U10258 (N_10258,N_10145,N_10059);
or U10259 (N_10259,N_10011,N_10095);
xor U10260 (N_10260,N_10101,N_10180);
xor U10261 (N_10261,N_10072,N_10113);
or U10262 (N_10262,N_10165,N_10183);
xnor U10263 (N_10263,N_10142,N_10021);
xor U10264 (N_10264,N_10157,N_10168);
nand U10265 (N_10265,N_10004,N_10144);
and U10266 (N_10266,N_10137,N_10169);
nor U10267 (N_10267,N_10182,N_10070);
xnor U10268 (N_10268,N_10010,N_10112);
or U10269 (N_10269,N_10084,N_10170);
xnor U10270 (N_10270,N_10189,N_10198);
nor U10271 (N_10271,N_10167,N_10031);
nand U10272 (N_10272,N_10038,N_10187);
or U10273 (N_10273,N_10023,N_10121);
nand U10274 (N_10274,N_10123,N_10188);
xnor U10275 (N_10275,N_10193,N_10035);
nand U10276 (N_10276,N_10158,N_10037);
xnor U10277 (N_10277,N_10057,N_10152);
nand U10278 (N_10278,N_10153,N_10065);
and U10279 (N_10279,N_10019,N_10046);
and U10280 (N_10280,N_10197,N_10024);
xnor U10281 (N_10281,N_10125,N_10124);
and U10282 (N_10282,N_10139,N_10116);
nor U10283 (N_10283,N_10181,N_10091);
nand U10284 (N_10284,N_10087,N_10195);
nand U10285 (N_10285,N_10088,N_10018);
or U10286 (N_10286,N_10047,N_10043);
xor U10287 (N_10287,N_10054,N_10148);
or U10288 (N_10288,N_10096,N_10049);
or U10289 (N_10289,N_10192,N_10108);
nor U10290 (N_10290,N_10111,N_10015);
and U10291 (N_10291,N_10034,N_10067);
and U10292 (N_10292,N_10161,N_10079);
nor U10293 (N_10293,N_10025,N_10039);
nand U10294 (N_10294,N_10143,N_10002);
and U10295 (N_10295,N_10085,N_10100);
nand U10296 (N_10296,N_10196,N_10178);
xnor U10297 (N_10297,N_10107,N_10179);
xnor U10298 (N_10298,N_10134,N_10120);
nand U10299 (N_10299,N_10075,N_10033);
and U10300 (N_10300,N_10057,N_10197);
and U10301 (N_10301,N_10062,N_10097);
xor U10302 (N_10302,N_10196,N_10095);
nor U10303 (N_10303,N_10148,N_10139);
nand U10304 (N_10304,N_10052,N_10163);
or U10305 (N_10305,N_10184,N_10187);
and U10306 (N_10306,N_10026,N_10040);
xor U10307 (N_10307,N_10026,N_10075);
xor U10308 (N_10308,N_10129,N_10033);
nand U10309 (N_10309,N_10105,N_10076);
and U10310 (N_10310,N_10126,N_10071);
nor U10311 (N_10311,N_10154,N_10180);
nor U10312 (N_10312,N_10146,N_10046);
and U10313 (N_10313,N_10004,N_10100);
or U10314 (N_10314,N_10024,N_10174);
xor U10315 (N_10315,N_10079,N_10075);
nand U10316 (N_10316,N_10147,N_10047);
and U10317 (N_10317,N_10032,N_10086);
xnor U10318 (N_10318,N_10080,N_10167);
nand U10319 (N_10319,N_10198,N_10064);
xnor U10320 (N_10320,N_10136,N_10028);
or U10321 (N_10321,N_10121,N_10125);
nand U10322 (N_10322,N_10026,N_10056);
nand U10323 (N_10323,N_10121,N_10086);
or U10324 (N_10324,N_10160,N_10109);
nor U10325 (N_10325,N_10122,N_10013);
and U10326 (N_10326,N_10094,N_10001);
xnor U10327 (N_10327,N_10115,N_10029);
or U10328 (N_10328,N_10074,N_10000);
and U10329 (N_10329,N_10080,N_10100);
xnor U10330 (N_10330,N_10183,N_10084);
nand U10331 (N_10331,N_10115,N_10083);
and U10332 (N_10332,N_10129,N_10044);
xor U10333 (N_10333,N_10091,N_10108);
nand U10334 (N_10334,N_10037,N_10174);
nand U10335 (N_10335,N_10074,N_10025);
or U10336 (N_10336,N_10166,N_10101);
or U10337 (N_10337,N_10107,N_10133);
nand U10338 (N_10338,N_10169,N_10061);
nand U10339 (N_10339,N_10060,N_10192);
or U10340 (N_10340,N_10139,N_10047);
and U10341 (N_10341,N_10195,N_10126);
nor U10342 (N_10342,N_10196,N_10106);
or U10343 (N_10343,N_10041,N_10100);
nor U10344 (N_10344,N_10160,N_10048);
nor U10345 (N_10345,N_10090,N_10006);
nor U10346 (N_10346,N_10026,N_10097);
xor U10347 (N_10347,N_10063,N_10090);
nand U10348 (N_10348,N_10064,N_10189);
nand U10349 (N_10349,N_10038,N_10013);
or U10350 (N_10350,N_10175,N_10135);
xor U10351 (N_10351,N_10116,N_10083);
xor U10352 (N_10352,N_10154,N_10017);
nand U10353 (N_10353,N_10075,N_10115);
nor U10354 (N_10354,N_10158,N_10115);
xnor U10355 (N_10355,N_10034,N_10017);
or U10356 (N_10356,N_10145,N_10107);
nor U10357 (N_10357,N_10148,N_10107);
or U10358 (N_10358,N_10175,N_10076);
and U10359 (N_10359,N_10121,N_10028);
xor U10360 (N_10360,N_10114,N_10152);
xor U10361 (N_10361,N_10066,N_10093);
nand U10362 (N_10362,N_10028,N_10125);
nor U10363 (N_10363,N_10138,N_10157);
and U10364 (N_10364,N_10145,N_10080);
nand U10365 (N_10365,N_10047,N_10031);
nor U10366 (N_10366,N_10040,N_10199);
nor U10367 (N_10367,N_10136,N_10032);
xor U10368 (N_10368,N_10101,N_10116);
or U10369 (N_10369,N_10061,N_10090);
nor U10370 (N_10370,N_10007,N_10114);
nand U10371 (N_10371,N_10038,N_10050);
nand U10372 (N_10372,N_10114,N_10165);
nand U10373 (N_10373,N_10031,N_10077);
xor U10374 (N_10374,N_10137,N_10170);
and U10375 (N_10375,N_10057,N_10070);
or U10376 (N_10376,N_10154,N_10008);
nor U10377 (N_10377,N_10176,N_10066);
and U10378 (N_10378,N_10144,N_10105);
nand U10379 (N_10379,N_10167,N_10025);
and U10380 (N_10380,N_10003,N_10076);
or U10381 (N_10381,N_10116,N_10144);
or U10382 (N_10382,N_10004,N_10184);
and U10383 (N_10383,N_10017,N_10110);
nand U10384 (N_10384,N_10047,N_10070);
and U10385 (N_10385,N_10110,N_10050);
xor U10386 (N_10386,N_10187,N_10001);
and U10387 (N_10387,N_10140,N_10041);
nor U10388 (N_10388,N_10149,N_10066);
or U10389 (N_10389,N_10162,N_10153);
or U10390 (N_10390,N_10194,N_10006);
nor U10391 (N_10391,N_10055,N_10161);
or U10392 (N_10392,N_10196,N_10066);
nand U10393 (N_10393,N_10057,N_10050);
nor U10394 (N_10394,N_10022,N_10110);
nor U10395 (N_10395,N_10119,N_10002);
nor U10396 (N_10396,N_10133,N_10181);
nor U10397 (N_10397,N_10103,N_10167);
nor U10398 (N_10398,N_10181,N_10023);
xnor U10399 (N_10399,N_10062,N_10128);
xor U10400 (N_10400,N_10218,N_10239);
nor U10401 (N_10401,N_10376,N_10341);
nand U10402 (N_10402,N_10396,N_10367);
nand U10403 (N_10403,N_10304,N_10289);
nand U10404 (N_10404,N_10221,N_10342);
nand U10405 (N_10405,N_10276,N_10270);
xor U10406 (N_10406,N_10348,N_10273);
xor U10407 (N_10407,N_10216,N_10345);
or U10408 (N_10408,N_10312,N_10208);
nand U10409 (N_10409,N_10334,N_10328);
or U10410 (N_10410,N_10384,N_10308);
or U10411 (N_10411,N_10288,N_10251);
nor U10412 (N_10412,N_10354,N_10359);
and U10413 (N_10413,N_10352,N_10329);
nor U10414 (N_10414,N_10387,N_10390);
xnor U10415 (N_10415,N_10351,N_10379);
or U10416 (N_10416,N_10202,N_10219);
and U10417 (N_10417,N_10398,N_10287);
nand U10418 (N_10418,N_10325,N_10200);
nor U10419 (N_10419,N_10301,N_10211);
or U10420 (N_10420,N_10245,N_10350);
nor U10421 (N_10421,N_10344,N_10298);
or U10422 (N_10422,N_10294,N_10243);
or U10423 (N_10423,N_10231,N_10306);
nand U10424 (N_10424,N_10386,N_10282);
xnor U10425 (N_10425,N_10284,N_10347);
and U10426 (N_10426,N_10353,N_10206);
xnor U10427 (N_10427,N_10349,N_10322);
and U10428 (N_10428,N_10346,N_10389);
and U10429 (N_10429,N_10255,N_10337);
and U10430 (N_10430,N_10254,N_10336);
nor U10431 (N_10431,N_10233,N_10210);
xor U10432 (N_10432,N_10280,N_10357);
nand U10433 (N_10433,N_10368,N_10331);
nand U10434 (N_10434,N_10295,N_10375);
or U10435 (N_10435,N_10303,N_10373);
nor U10436 (N_10436,N_10316,N_10319);
and U10437 (N_10437,N_10340,N_10235);
xnor U10438 (N_10438,N_10205,N_10247);
or U10439 (N_10439,N_10281,N_10394);
nand U10440 (N_10440,N_10260,N_10266);
nor U10441 (N_10441,N_10279,N_10381);
nand U10442 (N_10442,N_10309,N_10310);
or U10443 (N_10443,N_10225,N_10238);
nand U10444 (N_10444,N_10227,N_10307);
and U10445 (N_10445,N_10364,N_10201);
and U10446 (N_10446,N_10203,N_10356);
nor U10447 (N_10447,N_10326,N_10321);
nor U10448 (N_10448,N_10229,N_10237);
and U10449 (N_10449,N_10391,N_10212);
nor U10450 (N_10450,N_10256,N_10278);
nor U10451 (N_10451,N_10338,N_10392);
and U10452 (N_10452,N_10242,N_10264);
nor U10453 (N_10453,N_10220,N_10314);
and U10454 (N_10454,N_10230,N_10269);
and U10455 (N_10455,N_10234,N_10343);
xor U10456 (N_10456,N_10332,N_10267);
or U10457 (N_10457,N_10265,N_10313);
nand U10458 (N_10458,N_10222,N_10397);
nand U10459 (N_10459,N_10380,N_10371);
and U10460 (N_10460,N_10365,N_10204);
nand U10461 (N_10461,N_10291,N_10305);
and U10462 (N_10462,N_10393,N_10293);
and U10463 (N_10463,N_10207,N_10330);
xnor U10464 (N_10464,N_10296,N_10299);
or U10465 (N_10465,N_10327,N_10333);
or U10466 (N_10466,N_10209,N_10277);
nand U10467 (N_10467,N_10374,N_10317);
xor U10468 (N_10468,N_10388,N_10335);
nor U10469 (N_10469,N_10241,N_10372);
nand U10470 (N_10470,N_10360,N_10318);
or U10471 (N_10471,N_10369,N_10215);
xnor U10472 (N_10472,N_10385,N_10263);
nor U10473 (N_10473,N_10323,N_10226);
nand U10474 (N_10474,N_10274,N_10362);
xnor U10475 (N_10475,N_10223,N_10324);
and U10476 (N_10476,N_10258,N_10283);
and U10477 (N_10477,N_10224,N_10395);
xnor U10478 (N_10478,N_10302,N_10275);
xor U10479 (N_10479,N_10300,N_10297);
xor U10480 (N_10480,N_10236,N_10232);
and U10481 (N_10481,N_10290,N_10271);
xor U10482 (N_10482,N_10246,N_10315);
xnor U10483 (N_10483,N_10399,N_10272);
xnor U10484 (N_10484,N_10228,N_10240);
nand U10485 (N_10485,N_10286,N_10250);
or U10486 (N_10486,N_10366,N_10378);
nor U10487 (N_10487,N_10311,N_10377);
nand U10488 (N_10488,N_10382,N_10257);
xnor U10489 (N_10489,N_10292,N_10244);
and U10490 (N_10490,N_10358,N_10249);
and U10491 (N_10491,N_10285,N_10253);
nand U10492 (N_10492,N_10248,N_10213);
xnor U10493 (N_10493,N_10370,N_10339);
nand U10494 (N_10494,N_10383,N_10259);
and U10495 (N_10495,N_10261,N_10217);
and U10496 (N_10496,N_10252,N_10363);
xnor U10497 (N_10497,N_10268,N_10214);
or U10498 (N_10498,N_10355,N_10320);
nand U10499 (N_10499,N_10361,N_10262);
and U10500 (N_10500,N_10299,N_10352);
and U10501 (N_10501,N_10240,N_10222);
and U10502 (N_10502,N_10244,N_10253);
nor U10503 (N_10503,N_10308,N_10253);
or U10504 (N_10504,N_10215,N_10241);
nor U10505 (N_10505,N_10328,N_10318);
nor U10506 (N_10506,N_10254,N_10390);
and U10507 (N_10507,N_10304,N_10211);
and U10508 (N_10508,N_10225,N_10239);
nor U10509 (N_10509,N_10344,N_10361);
nand U10510 (N_10510,N_10368,N_10343);
nand U10511 (N_10511,N_10276,N_10261);
nor U10512 (N_10512,N_10200,N_10338);
nor U10513 (N_10513,N_10209,N_10331);
and U10514 (N_10514,N_10359,N_10250);
xnor U10515 (N_10515,N_10210,N_10246);
and U10516 (N_10516,N_10377,N_10388);
nor U10517 (N_10517,N_10357,N_10247);
nor U10518 (N_10518,N_10377,N_10259);
xnor U10519 (N_10519,N_10301,N_10277);
or U10520 (N_10520,N_10255,N_10311);
or U10521 (N_10521,N_10330,N_10323);
and U10522 (N_10522,N_10226,N_10347);
or U10523 (N_10523,N_10240,N_10241);
and U10524 (N_10524,N_10391,N_10257);
or U10525 (N_10525,N_10283,N_10213);
nand U10526 (N_10526,N_10343,N_10299);
or U10527 (N_10527,N_10375,N_10275);
and U10528 (N_10528,N_10274,N_10324);
nor U10529 (N_10529,N_10372,N_10319);
nand U10530 (N_10530,N_10201,N_10308);
nor U10531 (N_10531,N_10296,N_10261);
or U10532 (N_10532,N_10389,N_10310);
and U10533 (N_10533,N_10252,N_10368);
and U10534 (N_10534,N_10372,N_10388);
nand U10535 (N_10535,N_10270,N_10226);
xor U10536 (N_10536,N_10276,N_10324);
or U10537 (N_10537,N_10343,N_10388);
nand U10538 (N_10538,N_10363,N_10379);
nor U10539 (N_10539,N_10285,N_10245);
xnor U10540 (N_10540,N_10275,N_10333);
or U10541 (N_10541,N_10259,N_10295);
xor U10542 (N_10542,N_10361,N_10250);
xnor U10543 (N_10543,N_10364,N_10238);
and U10544 (N_10544,N_10321,N_10268);
xnor U10545 (N_10545,N_10254,N_10265);
and U10546 (N_10546,N_10273,N_10280);
xnor U10547 (N_10547,N_10367,N_10378);
and U10548 (N_10548,N_10242,N_10256);
xnor U10549 (N_10549,N_10324,N_10235);
xnor U10550 (N_10550,N_10349,N_10208);
nor U10551 (N_10551,N_10293,N_10398);
and U10552 (N_10552,N_10318,N_10239);
and U10553 (N_10553,N_10252,N_10333);
nor U10554 (N_10554,N_10380,N_10378);
and U10555 (N_10555,N_10353,N_10336);
xnor U10556 (N_10556,N_10378,N_10233);
nor U10557 (N_10557,N_10323,N_10390);
nand U10558 (N_10558,N_10389,N_10321);
and U10559 (N_10559,N_10238,N_10287);
or U10560 (N_10560,N_10369,N_10310);
and U10561 (N_10561,N_10318,N_10386);
nand U10562 (N_10562,N_10361,N_10205);
xnor U10563 (N_10563,N_10226,N_10300);
or U10564 (N_10564,N_10383,N_10267);
xnor U10565 (N_10565,N_10259,N_10249);
or U10566 (N_10566,N_10314,N_10254);
nand U10567 (N_10567,N_10399,N_10237);
xor U10568 (N_10568,N_10366,N_10238);
and U10569 (N_10569,N_10222,N_10358);
nand U10570 (N_10570,N_10357,N_10285);
or U10571 (N_10571,N_10205,N_10377);
or U10572 (N_10572,N_10369,N_10303);
xor U10573 (N_10573,N_10339,N_10349);
or U10574 (N_10574,N_10219,N_10324);
nand U10575 (N_10575,N_10252,N_10262);
and U10576 (N_10576,N_10356,N_10330);
and U10577 (N_10577,N_10243,N_10389);
nand U10578 (N_10578,N_10269,N_10202);
nand U10579 (N_10579,N_10280,N_10287);
nor U10580 (N_10580,N_10225,N_10360);
and U10581 (N_10581,N_10280,N_10343);
and U10582 (N_10582,N_10340,N_10368);
nor U10583 (N_10583,N_10274,N_10307);
nand U10584 (N_10584,N_10293,N_10277);
or U10585 (N_10585,N_10350,N_10308);
and U10586 (N_10586,N_10381,N_10253);
nor U10587 (N_10587,N_10304,N_10311);
nor U10588 (N_10588,N_10294,N_10374);
nand U10589 (N_10589,N_10323,N_10346);
xnor U10590 (N_10590,N_10249,N_10304);
and U10591 (N_10591,N_10323,N_10305);
or U10592 (N_10592,N_10254,N_10338);
or U10593 (N_10593,N_10218,N_10383);
or U10594 (N_10594,N_10244,N_10393);
xor U10595 (N_10595,N_10362,N_10396);
nor U10596 (N_10596,N_10334,N_10222);
or U10597 (N_10597,N_10358,N_10229);
nand U10598 (N_10598,N_10245,N_10249);
xnor U10599 (N_10599,N_10221,N_10362);
nand U10600 (N_10600,N_10522,N_10550);
nand U10601 (N_10601,N_10485,N_10532);
nand U10602 (N_10602,N_10432,N_10442);
or U10603 (N_10603,N_10533,N_10409);
or U10604 (N_10604,N_10407,N_10555);
nand U10605 (N_10605,N_10448,N_10521);
nor U10606 (N_10606,N_10591,N_10567);
or U10607 (N_10607,N_10437,N_10509);
or U10608 (N_10608,N_10411,N_10510);
or U10609 (N_10609,N_10529,N_10462);
nand U10610 (N_10610,N_10464,N_10401);
xor U10611 (N_10611,N_10421,N_10547);
and U10612 (N_10612,N_10424,N_10497);
xnor U10613 (N_10613,N_10447,N_10428);
and U10614 (N_10614,N_10441,N_10508);
xnor U10615 (N_10615,N_10470,N_10518);
xor U10616 (N_10616,N_10570,N_10520);
nor U10617 (N_10617,N_10513,N_10561);
and U10618 (N_10618,N_10495,N_10572);
and U10619 (N_10619,N_10482,N_10478);
nand U10620 (N_10620,N_10549,N_10526);
or U10621 (N_10621,N_10493,N_10562);
and U10622 (N_10622,N_10468,N_10425);
nor U10623 (N_10623,N_10423,N_10492);
and U10624 (N_10624,N_10575,N_10466);
and U10625 (N_10625,N_10435,N_10461);
or U10626 (N_10626,N_10429,N_10576);
nand U10627 (N_10627,N_10552,N_10494);
or U10628 (N_10628,N_10586,N_10587);
nand U10629 (N_10629,N_10525,N_10571);
xnor U10630 (N_10630,N_10515,N_10419);
nor U10631 (N_10631,N_10457,N_10582);
and U10632 (N_10632,N_10475,N_10481);
xnor U10633 (N_10633,N_10476,N_10438);
or U10634 (N_10634,N_10463,N_10584);
nand U10635 (N_10635,N_10431,N_10566);
nor U10636 (N_10636,N_10498,N_10543);
xnor U10637 (N_10637,N_10568,N_10544);
and U10638 (N_10638,N_10472,N_10455);
nor U10639 (N_10639,N_10454,N_10404);
xnor U10640 (N_10640,N_10487,N_10592);
and U10641 (N_10641,N_10413,N_10405);
or U10642 (N_10642,N_10579,N_10528);
and U10643 (N_10643,N_10519,N_10469);
or U10644 (N_10644,N_10406,N_10593);
nor U10645 (N_10645,N_10563,N_10542);
nand U10646 (N_10646,N_10574,N_10598);
nor U10647 (N_10647,N_10569,N_10556);
xor U10648 (N_10648,N_10449,N_10506);
xor U10649 (N_10649,N_10430,N_10443);
xnor U10650 (N_10650,N_10459,N_10588);
and U10651 (N_10651,N_10467,N_10565);
nand U10652 (N_10652,N_10536,N_10530);
nor U10653 (N_10653,N_10436,N_10512);
xnor U10654 (N_10654,N_10440,N_10502);
nor U10655 (N_10655,N_10573,N_10417);
nand U10656 (N_10656,N_10581,N_10460);
nor U10657 (N_10657,N_10484,N_10596);
and U10658 (N_10658,N_10585,N_10595);
nand U10659 (N_10659,N_10465,N_10445);
nor U10660 (N_10660,N_10444,N_10402);
xor U10661 (N_10661,N_10546,N_10516);
xor U10662 (N_10662,N_10558,N_10505);
xor U10663 (N_10663,N_10496,N_10499);
nand U10664 (N_10664,N_10408,N_10523);
or U10665 (N_10665,N_10415,N_10527);
and U10666 (N_10666,N_10486,N_10450);
xor U10667 (N_10667,N_10507,N_10531);
xor U10668 (N_10668,N_10557,N_10534);
nand U10669 (N_10669,N_10500,N_10540);
nor U10670 (N_10670,N_10560,N_10427);
nor U10671 (N_10671,N_10451,N_10577);
and U10672 (N_10672,N_10412,N_10594);
nand U10673 (N_10673,N_10599,N_10418);
xor U10674 (N_10674,N_10473,N_10410);
nand U10675 (N_10675,N_10535,N_10564);
and U10676 (N_10676,N_10483,N_10553);
nor U10677 (N_10677,N_10479,N_10578);
or U10678 (N_10678,N_10400,N_10490);
and U10679 (N_10679,N_10583,N_10501);
nand U10680 (N_10680,N_10580,N_10511);
xnor U10681 (N_10681,N_10589,N_10597);
nand U10682 (N_10682,N_10474,N_10446);
and U10683 (N_10683,N_10538,N_10403);
xnor U10684 (N_10684,N_10503,N_10545);
and U10685 (N_10685,N_10414,N_10524);
and U10686 (N_10686,N_10539,N_10541);
nor U10687 (N_10687,N_10477,N_10452);
or U10688 (N_10688,N_10517,N_10439);
or U10689 (N_10689,N_10453,N_10434);
and U10690 (N_10690,N_10416,N_10590);
xnor U10691 (N_10691,N_10420,N_10504);
xnor U10692 (N_10692,N_10491,N_10489);
nor U10693 (N_10693,N_10559,N_10480);
and U10694 (N_10694,N_10433,N_10456);
nor U10695 (N_10695,N_10537,N_10458);
nor U10696 (N_10696,N_10471,N_10514);
and U10697 (N_10697,N_10426,N_10488);
or U10698 (N_10698,N_10551,N_10422);
or U10699 (N_10699,N_10554,N_10548);
nor U10700 (N_10700,N_10434,N_10512);
nor U10701 (N_10701,N_10504,N_10598);
or U10702 (N_10702,N_10594,N_10588);
nor U10703 (N_10703,N_10588,N_10530);
nand U10704 (N_10704,N_10438,N_10493);
or U10705 (N_10705,N_10597,N_10493);
nand U10706 (N_10706,N_10561,N_10552);
or U10707 (N_10707,N_10594,N_10543);
and U10708 (N_10708,N_10544,N_10539);
and U10709 (N_10709,N_10496,N_10517);
nor U10710 (N_10710,N_10431,N_10475);
and U10711 (N_10711,N_10484,N_10529);
or U10712 (N_10712,N_10594,N_10464);
nor U10713 (N_10713,N_10488,N_10547);
or U10714 (N_10714,N_10536,N_10541);
or U10715 (N_10715,N_10523,N_10497);
nand U10716 (N_10716,N_10502,N_10535);
or U10717 (N_10717,N_10477,N_10529);
and U10718 (N_10718,N_10556,N_10456);
or U10719 (N_10719,N_10525,N_10488);
nor U10720 (N_10720,N_10559,N_10562);
xor U10721 (N_10721,N_10486,N_10446);
nor U10722 (N_10722,N_10428,N_10426);
and U10723 (N_10723,N_10458,N_10464);
nor U10724 (N_10724,N_10549,N_10405);
and U10725 (N_10725,N_10506,N_10529);
nor U10726 (N_10726,N_10545,N_10557);
nor U10727 (N_10727,N_10507,N_10501);
xor U10728 (N_10728,N_10525,N_10541);
and U10729 (N_10729,N_10447,N_10546);
or U10730 (N_10730,N_10501,N_10486);
and U10731 (N_10731,N_10401,N_10532);
or U10732 (N_10732,N_10565,N_10478);
xnor U10733 (N_10733,N_10412,N_10564);
or U10734 (N_10734,N_10410,N_10553);
and U10735 (N_10735,N_10476,N_10477);
or U10736 (N_10736,N_10463,N_10466);
or U10737 (N_10737,N_10457,N_10558);
nor U10738 (N_10738,N_10583,N_10448);
and U10739 (N_10739,N_10465,N_10428);
or U10740 (N_10740,N_10449,N_10510);
xnor U10741 (N_10741,N_10443,N_10503);
nor U10742 (N_10742,N_10526,N_10508);
nand U10743 (N_10743,N_10591,N_10574);
or U10744 (N_10744,N_10474,N_10528);
nor U10745 (N_10745,N_10578,N_10434);
nand U10746 (N_10746,N_10433,N_10565);
nor U10747 (N_10747,N_10414,N_10424);
xnor U10748 (N_10748,N_10549,N_10522);
and U10749 (N_10749,N_10401,N_10544);
nor U10750 (N_10750,N_10475,N_10439);
and U10751 (N_10751,N_10473,N_10586);
or U10752 (N_10752,N_10550,N_10590);
and U10753 (N_10753,N_10543,N_10475);
nor U10754 (N_10754,N_10579,N_10486);
nor U10755 (N_10755,N_10440,N_10443);
xnor U10756 (N_10756,N_10402,N_10416);
and U10757 (N_10757,N_10520,N_10423);
and U10758 (N_10758,N_10574,N_10551);
and U10759 (N_10759,N_10431,N_10491);
or U10760 (N_10760,N_10534,N_10435);
nand U10761 (N_10761,N_10474,N_10511);
or U10762 (N_10762,N_10421,N_10540);
nand U10763 (N_10763,N_10425,N_10421);
and U10764 (N_10764,N_10504,N_10442);
and U10765 (N_10765,N_10437,N_10404);
nor U10766 (N_10766,N_10573,N_10519);
nor U10767 (N_10767,N_10442,N_10457);
nor U10768 (N_10768,N_10551,N_10569);
nor U10769 (N_10769,N_10424,N_10588);
and U10770 (N_10770,N_10565,N_10535);
xor U10771 (N_10771,N_10500,N_10459);
or U10772 (N_10772,N_10555,N_10451);
xor U10773 (N_10773,N_10538,N_10429);
or U10774 (N_10774,N_10478,N_10548);
and U10775 (N_10775,N_10577,N_10523);
xor U10776 (N_10776,N_10408,N_10502);
nor U10777 (N_10777,N_10552,N_10474);
xnor U10778 (N_10778,N_10516,N_10587);
nand U10779 (N_10779,N_10415,N_10549);
and U10780 (N_10780,N_10572,N_10540);
or U10781 (N_10781,N_10467,N_10560);
xor U10782 (N_10782,N_10501,N_10408);
and U10783 (N_10783,N_10501,N_10481);
xnor U10784 (N_10784,N_10557,N_10537);
or U10785 (N_10785,N_10481,N_10429);
or U10786 (N_10786,N_10402,N_10520);
or U10787 (N_10787,N_10573,N_10496);
xor U10788 (N_10788,N_10526,N_10524);
xnor U10789 (N_10789,N_10559,N_10409);
and U10790 (N_10790,N_10413,N_10545);
xnor U10791 (N_10791,N_10490,N_10418);
and U10792 (N_10792,N_10466,N_10493);
or U10793 (N_10793,N_10576,N_10580);
xnor U10794 (N_10794,N_10427,N_10461);
nor U10795 (N_10795,N_10489,N_10573);
and U10796 (N_10796,N_10551,N_10496);
nand U10797 (N_10797,N_10435,N_10535);
and U10798 (N_10798,N_10407,N_10595);
nor U10799 (N_10799,N_10593,N_10453);
xor U10800 (N_10800,N_10622,N_10754);
nor U10801 (N_10801,N_10660,N_10667);
xor U10802 (N_10802,N_10774,N_10605);
nand U10803 (N_10803,N_10656,N_10785);
xor U10804 (N_10804,N_10649,N_10752);
xnor U10805 (N_10805,N_10628,N_10681);
nand U10806 (N_10806,N_10790,N_10697);
nand U10807 (N_10807,N_10627,N_10609);
xnor U10808 (N_10808,N_10648,N_10778);
or U10809 (N_10809,N_10693,N_10750);
nand U10810 (N_10810,N_10712,N_10773);
and U10811 (N_10811,N_10634,N_10621);
and U10812 (N_10812,N_10736,N_10714);
nor U10813 (N_10813,N_10610,N_10601);
nor U10814 (N_10814,N_10682,N_10705);
nand U10815 (N_10815,N_10767,N_10701);
nand U10816 (N_10816,N_10633,N_10607);
xnor U10817 (N_10817,N_10685,N_10661);
nand U10818 (N_10818,N_10738,N_10798);
and U10819 (N_10819,N_10692,N_10613);
nor U10820 (N_10820,N_10637,N_10710);
nand U10821 (N_10821,N_10762,N_10679);
or U10822 (N_10822,N_10741,N_10706);
nor U10823 (N_10823,N_10620,N_10703);
xnor U10824 (N_10824,N_10603,N_10678);
and U10825 (N_10825,N_10626,N_10787);
and U10826 (N_10826,N_10675,N_10641);
nand U10827 (N_10827,N_10658,N_10683);
and U10828 (N_10828,N_10746,N_10642);
and U10829 (N_10829,N_10791,N_10756);
or U10830 (N_10830,N_10770,N_10629);
or U10831 (N_10831,N_10696,N_10611);
or U10832 (N_10832,N_10740,N_10698);
or U10833 (N_10833,N_10725,N_10733);
xnor U10834 (N_10834,N_10751,N_10650);
nor U10835 (N_10835,N_10639,N_10781);
nor U10836 (N_10836,N_10619,N_10772);
nand U10837 (N_10837,N_10753,N_10764);
xnor U10838 (N_10838,N_10795,N_10794);
nand U10839 (N_10839,N_10666,N_10789);
or U10840 (N_10840,N_10635,N_10769);
nor U10841 (N_10841,N_10677,N_10744);
or U10842 (N_10842,N_10797,N_10689);
nor U10843 (N_10843,N_10732,N_10748);
nor U10844 (N_10844,N_10788,N_10676);
and U10845 (N_10845,N_10796,N_10686);
or U10846 (N_10846,N_10652,N_10721);
nor U10847 (N_10847,N_10600,N_10776);
and U10848 (N_10848,N_10799,N_10779);
and U10849 (N_10849,N_10631,N_10640);
or U10850 (N_10850,N_10690,N_10674);
xnor U10851 (N_10851,N_10657,N_10636);
and U10852 (N_10852,N_10731,N_10763);
nand U10853 (N_10853,N_10694,N_10688);
nor U10854 (N_10854,N_10726,N_10782);
nor U10855 (N_10855,N_10735,N_10654);
or U10856 (N_10856,N_10616,N_10625);
nor U10857 (N_10857,N_10644,N_10711);
xor U10858 (N_10858,N_10671,N_10687);
or U10859 (N_10859,N_10715,N_10624);
nand U10860 (N_10860,N_10783,N_10646);
nand U10861 (N_10861,N_10665,N_10647);
or U10862 (N_10862,N_10713,N_10775);
nand U10863 (N_10863,N_10645,N_10655);
nand U10864 (N_10864,N_10691,N_10618);
xnor U10865 (N_10865,N_10632,N_10670);
xor U10866 (N_10866,N_10760,N_10716);
or U10867 (N_10867,N_10730,N_10662);
xnor U10868 (N_10868,N_10630,N_10668);
and U10869 (N_10869,N_10793,N_10722);
and U10870 (N_10870,N_10784,N_10758);
nand U10871 (N_10871,N_10673,N_10765);
nor U10872 (N_10872,N_10608,N_10612);
nand U10873 (N_10873,N_10695,N_10743);
nor U10874 (N_10874,N_10720,N_10709);
nand U10875 (N_10875,N_10728,N_10606);
nor U10876 (N_10876,N_10729,N_10604);
nor U10877 (N_10877,N_10704,N_10643);
or U10878 (N_10878,N_10602,N_10653);
nand U10879 (N_10879,N_10702,N_10700);
nor U10880 (N_10880,N_10663,N_10734);
nand U10881 (N_10881,N_10615,N_10766);
and U10882 (N_10882,N_10718,N_10672);
nand U10883 (N_10883,N_10717,N_10680);
nor U10884 (N_10884,N_10708,N_10786);
nand U10885 (N_10885,N_10761,N_10707);
and U10886 (N_10886,N_10623,N_10759);
nand U10887 (N_10887,N_10768,N_10727);
nor U10888 (N_10888,N_10719,N_10777);
nor U10889 (N_10889,N_10724,N_10723);
xor U10890 (N_10890,N_10780,N_10669);
or U10891 (N_10891,N_10664,N_10651);
or U10892 (N_10892,N_10771,N_10742);
nand U10893 (N_10893,N_10745,N_10739);
nand U10894 (N_10894,N_10749,N_10757);
and U10895 (N_10895,N_10659,N_10747);
nor U10896 (N_10896,N_10699,N_10684);
or U10897 (N_10897,N_10617,N_10737);
nand U10898 (N_10898,N_10792,N_10638);
nand U10899 (N_10899,N_10755,N_10614);
xor U10900 (N_10900,N_10712,N_10754);
xor U10901 (N_10901,N_10725,N_10636);
nor U10902 (N_10902,N_10705,N_10657);
xor U10903 (N_10903,N_10747,N_10633);
or U10904 (N_10904,N_10729,N_10703);
and U10905 (N_10905,N_10671,N_10736);
nand U10906 (N_10906,N_10775,N_10679);
or U10907 (N_10907,N_10644,N_10721);
nand U10908 (N_10908,N_10647,N_10781);
nor U10909 (N_10909,N_10677,N_10622);
xor U10910 (N_10910,N_10797,N_10637);
or U10911 (N_10911,N_10765,N_10637);
nand U10912 (N_10912,N_10754,N_10645);
and U10913 (N_10913,N_10626,N_10638);
and U10914 (N_10914,N_10646,N_10727);
and U10915 (N_10915,N_10693,N_10651);
and U10916 (N_10916,N_10722,N_10730);
and U10917 (N_10917,N_10607,N_10737);
nor U10918 (N_10918,N_10691,N_10798);
nand U10919 (N_10919,N_10672,N_10739);
xor U10920 (N_10920,N_10625,N_10784);
xnor U10921 (N_10921,N_10754,N_10781);
or U10922 (N_10922,N_10653,N_10697);
or U10923 (N_10923,N_10645,N_10661);
nor U10924 (N_10924,N_10749,N_10787);
or U10925 (N_10925,N_10667,N_10676);
and U10926 (N_10926,N_10774,N_10682);
and U10927 (N_10927,N_10732,N_10686);
xor U10928 (N_10928,N_10685,N_10606);
or U10929 (N_10929,N_10760,N_10656);
nor U10930 (N_10930,N_10663,N_10792);
and U10931 (N_10931,N_10726,N_10715);
nand U10932 (N_10932,N_10636,N_10702);
nand U10933 (N_10933,N_10737,N_10794);
xor U10934 (N_10934,N_10740,N_10659);
or U10935 (N_10935,N_10600,N_10744);
and U10936 (N_10936,N_10621,N_10765);
nand U10937 (N_10937,N_10748,N_10659);
and U10938 (N_10938,N_10732,N_10689);
or U10939 (N_10939,N_10785,N_10639);
nor U10940 (N_10940,N_10696,N_10666);
nand U10941 (N_10941,N_10616,N_10797);
xnor U10942 (N_10942,N_10627,N_10734);
xnor U10943 (N_10943,N_10715,N_10605);
nor U10944 (N_10944,N_10688,N_10619);
nor U10945 (N_10945,N_10628,N_10715);
xor U10946 (N_10946,N_10692,N_10663);
or U10947 (N_10947,N_10618,N_10658);
nor U10948 (N_10948,N_10703,N_10765);
nor U10949 (N_10949,N_10798,N_10635);
and U10950 (N_10950,N_10730,N_10622);
nor U10951 (N_10951,N_10787,N_10602);
and U10952 (N_10952,N_10670,N_10658);
or U10953 (N_10953,N_10634,N_10700);
xnor U10954 (N_10954,N_10631,N_10646);
and U10955 (N_10955,N_10707,N_10733);
and U10956 (N_10956,N_10734,N_10794);
nand U10957 (N_10957,N_10612,N_10755);
and U10958 (N_10958,N_10688,N_10615);
or U10959 (N_10959,N_10785,N_10629);
xor U10960 (N_10960,N_10619,N_10643);
xor U10961 (N_10961,N_10702,N_10685);
xor U10962 (N_10962,N_10776,N_10645);
and U10963 (N_10963,N_10749,N_10763);
nand U10964 (N_10964,N_10797,N_10719);
or U10965 (N_10965,N_10614,N_10612);
and U10966 (N_10966,N_10671,N_10727);
and U10967 (N_10967,N_10641,N_10629);
nor U10968 (N_10968,N_10757,N_10785);
or U10969 (N_10969,N_10689,N_10601);
and U10970 (N_10970,N_10765,N_10653);
and U10971 (N_10971,N_10668,N_10690);
nor U10972 (N_10972,N_10632,N_10680);
nand U10973 (N_10973,N_10662,N_10710);
nand U10974 (N_10974,N_10652,N_10678);
xnor U10975 (N_10975,N_10768,N_10777);
or U10976 (N_10976,N_10703,N_10617);
nand U10977 (N_10977,N_10774,N_10723);
or U10978 (N_10978,N_10611,N_10601);
nor U10979 (N_10979,N_10667,N_10611);
xnor U10980 (N_10980,N_10732,N_10624);
nand U10981 (N_10981,N_10620,N_10723);
xnor U10982 (N_10982,N_10616,N_10609);
xor U10983 (N_10983,N_10719,N_10735);
xor U10984 (N_10984,N_10603,N_10697);
or U10985 (N_10985,N_10797,N_10623);
nor U10986 (N_10986,N_10640,N_10714);
nand U10987 (N_10987,N_10786,N_10626);
nand U10988 (N_10988,N_10733,N_10772);
or U10989 (N_10989,N_10778,N_10797);
and U10990 (N_10990,N_10665,N_10602);
xor U10991 (N_10991,N_10651,N_10729);
nand U10992 (N_10992,N_10622,N_10698);
nor U10993 (N_10993,N_10663,N_10758);
nor U10994 (N_10994,N_10650,N_10790);
or U10995 (N_10995,N_10741,N_10724);
xor U10996 (N_10996,N_10787,N_10663);
and U10997 (N_10997,N_10797,N_10701);
xnor U10998 (N_10998,N_10643,N_10768);
or U10999 (N_10999,N_10745,N_10603);
nor U11000 (N_11000,N_10927,N_10954);
nor U11001 (N_11001,N_10864,N_10949);
or U11002 (N_11002,N_10856,N_10943);
xor U11003 (N_11003,N_10879,N_10939);
or U11004 (N_11004,N_10809,N_10999);
xnor U11005 (N_11005,N_10937,N_10898);
nand U11006 (N_11006,N_10946,N_10851);
nand U11007 (N_11007,N_10912,N_10974);
or U11008 (N_11008,N_10890,N_10828);
nor U11009 (N_11009,N_10995,N_10867);
or U11010 (N_11010,N_10883,N_10846);
nor U11011 (N_11011,N_10819,N_10972);
nand U11012 (N_11012,N_10895,N_10905);
or U11013 (N_11013,N_10909,N_10823);
or U11014 (N_11014,N_10947,N_10904);
or U11015 (N_11015,N_10994,N_10929);
xnor U11016 (N_11016,N_10858,N_10922);
nor U11017 (N_11017,N_10991,N_10936);
nand U11018 (N_11018,N_10810,N_10825);
xnor U11019 (N_11019,N_10873,N_10827);
or U11020 (N_11020,N_10934,N_10921);
and U11021 (N_11021,N_10812,N_10985);
and U11022 (N_11022,N_10884,N_10888);
nor U11023 (N_11023,N_10913,N_10882);
xnor U11024 (N_11024,N_10981,N_10896);
nand U11025 (N_11025,N_10847,N_10822);
nand U11026 (N_11026,N_10990,N_10925);
and U11027 (N_11027,N_10992,N_10915);
nand U11028 (N_11028,N_10801,N_10857);
or U11029 (N_11029,N_10916,N_10861);
and U11030 (N_11030,N_10869,N_10868);
and U11031 (N_11031,N_10901,N_10848);
nor U11032 (N_11032,N_10983,N_10806);
xnor U11033 (N_11033,N_10963,N_10826);
and U11034 (N_11034,N_10850,N_10986);
or U11035 (N_11035,N_10807,N_10887);
and U11036 (N_11036,N_10821,N_10804);
or U11037 (N_11037,N_10930,N_10965);
xor U11038 (N_11038,N_10892,N_10978);
nand U11039 (N_11039,N_10933,N_10811);
xnor U11040 (N_11040,N_10914,N_10897);
nand U11041 (N_11041,N_10871,N_10935);
xnor U11042 (N_11042,N_10956,N_10942);
nor U11043 (N_11043,N_10923,N_10958);
xnor U11044 (N_11044,N_10960,N_10932);
nor U11045 (N_11045,N_10808,N_10803);
xor U11046 (N_11046,N_10950,N_10989);
xor U11047 (N_11047,N_10993,N_10967);
nor U11048 (N_11048,N_10820,N_10906);
nand U11049 (N_11049,N_10813,N_10860);
or U11050 (N_11050,N_10957,N_10816);
nand U11051 (N_11051,N_10900,N_10845);
or U11052 (N_11052,N_10945,N_10910);
or U11053 (N_11053,N_10908,N_10969);
nor U11054 (N_11054,N_10870,N_10815);
xnor U11055 (N_11055,N_10829,N_10959);
and U11056 (N_11056,N_10878,N_10842);
nor U11057 (N_11057,N_10885,N_10970);
xor U11058 (N_11058,N_10824,N_10832);
nor U11059 (N_11059,N_10952,N_10982);
or U11060 (N_11060,N_10891,N_10971);
nand U11061 (N_11061,N_10893,N_10940);
nor U11062 (N_11062,N_10944,N_10839);
xor U11063 (N_11063,N_10968,N_10997);
or U11064 (N_11064,N_10902,N_10840);
nand U11065 (N_11065,N_10931,N_10966);
nor U11066 (N_11066,N_10855,N_10838);
or U11067 (N_11067,N_10862,N_10903);
nand U11068 (N_11068,N_10833,N_10876);
or U11069 (N_11069,N_10941,N_10863);
and U11070 (N_11070,N_10889,N_10928);
and U11071 (N_11071,N_10874,N_10911);
nor U11072 (N_11072,N_10805,N_10853);
nand U11073 (N_11073,N_10854,N_10852);
xnor U11074 (N_11074,N_10975,N_10899);
and U11075 (N_11075,N_10918,N_10977);
nand U11076 (N_11076,N_10955,N_10938);
nand U11077 (N_11077,N_10881,N_10830);
nand U11078 (N_11078,N_10987,N_10926);
nor U11079 (N_11079,N_10831,N_10817);
xor U11080 (N_11080,N_10872,N_10800);
xnor U11081 (N_11081,N_10973,N_10841);
xor U11082 (N_11082,N_10961,N_10907);
or U11083 (N_11083,N_10951,N_10976);
and U11084 (N_11084,N_10920,N_10866);
or U11085 (N_11085,N_10844,N_10877);
nand U11086 (N_11086,N_10948,N_10886);
nor U11087 (N_11087,N_10835,N_10849);
nor U11088 (N_11088,N_10924,N_10880);
nand U11089 (N_11089,N_10962,N_10953);
or U11090 (N_11090,N_10834,N_10802);
nand U11091 (N_11091,N_10980,N_10984);
xor U11092 (N_11092,N_10843,N_10998);
nor U11093 (N_11093,N_10836,N_10875);
nor U11094 (N_11094,N_10859,N_10964);
nor U11095 (N_11095,N_10865,N_10919);
or U11096 (N_11096,N_10894,N_10996);
nor U11097 (N_11097,N_10979,N_10837);
and U11098 (N_11098,N_10818,N_10988);
nand U11099 (N_11099,N_10814,N_10917);
xor U11100 (N_11100,N_10949,N_10839);
nand U11101 (N_11101,N_10976,N_10947);
xor U11102 (N_11102,N_10900,N_10858);
or U11103 (N_11103,N_10969,N_10976);
and U11104 (N_11104,N_10981,N_10872);
nor U11105 (N_11105,N_10935,N_10916);
nand U11106 (N_11106,N_10847,N_10930);
nand U11107 (N_11107,N_10858,N_10812);
and U11108 (N_11108,N_10912,N_10854);
and U11109 (N_11109,N_10958,N_10843);
and U11110 (N_11110,N_10928,N_10999);
xnor U11111 (N_11111,N_10955,N_10859);
nor U11112 (N_11112,N_10873,N_10941);
nor U11113 (N_11113,N_10844,N_10949);
and U11114 (N_11114,N_10847,N_10977);
nor U11115 (N_11115,N_10826,N_10880);
or U11116 (N_11116,N_10856,N_10928);
nand U11117 (N_11117,N_10903,N_10941);
xnor U11118 (N_11118,N_10893,N_10886);
and U11119 (N_11119,N_10985,N_10873);
nor U11120 (N_11120,N_10870,N_10832);
and U11121 (N_11121,N_10934,N_10813);
nand U11122 (N_11122,N_10817,N_10967);
nor U11123 (N_11123,N_10972,N_10913);
and U11124 (N_11124,N_10825,N_10808);
nand U11125 (N_11125,N_10968,N_10949);
or U11126 (N_11126,N_10900,N_10954);
xor U11127 (N_11127,N_10891,N_10981);
nor U11128 (N_11128,N_10801,N_10865);
xnor U11129 (N_11129,N_10999,N_10968);
and U11130 (N_11130,N_10937,N_10954);
nor U11131 (N_11131,N_10807,N_10935);
and U11132 (N_11132,N_10835,N_10937);
xor U11133 (N_11133,N_10840,N_10826);
or U11134 (N_11134,N_10923,N_10885);
or U11135 (N_11135,N_10827,N_10993);
or U11136 (N_11136,N_10956,N_10843);
nor U11137 (N_11137,N_10852,N_10805);
xnor U11138 (N_11138,N_10868,N_10828);
nor U11139 (N_11139,N_10845,N_10967);
and U11140 (N_11140,N_10856,N_10974);
and U11141 (N_11141,N_10807,N_10896);
nor U11142 (N_11142,N_10901,N_10950);
xnor U11143 (N_11143,N_10980,N_10879);
or U11144 (N_11144,N_10903,N_10908);
xnor U11145 (N_11145,N_10849,N_10886);
xnor U11146 (N_11146,N_10992,N_10849);
nand U11147 (N_11147,N_10889,N_10932);
nor U11148 (N_11148,N_10875,N_10975);
and U11149 (N_11149,N_10803,N_10967);
and U11150 (N_11150,N_10865,N_10982);
and U11151 (N_11151,N_10886,N_10836);
nor U11152 (N_11152,N_10875,N_10849);
and U11153 (N_11153,N_10978,N_10835);
nor U11154 (N_11154,N_10824,N_10944);
and U11155 (N_11155,N_10878,N_10893);
xnor U11156 (N_11156,N_10861,N_10906);
xnor U11157 (N_11157,N_10977,N_10941);
xnor U11158 (N_11158,N_10875,N_10915);
nand U11159 (N_11159,N_10914,N_10995);
nor U11160 (N_11160,N_10926,N_10914);
or U11161 (N_11161,N_10845,N_10906);
xnor U11162 (N_11162,N_10978,N_10937);
and U11163 (N_11163,N_10899,N_10937);
and U11164 (N_11164,N_10806,N_10823);
or U11165 (N_11165,N_10815,N_10918);
nand U11166 (N_11166,N_10936,N_10807);
nor U11167 (N_11167,N_10890,N_10959);
nor U11168 (N_11168,N_10816,N_10907);
or U11169 (N_11169,N_10962,N_10983);
nor U11170 (N_11170,N_10999,N_10882);
or U11171 (N_11171,N_10849,N_10862);
or U11172 (N_11172,N_10921,N_10826);
and U11173 (N_11173,N_10933,N_10944);
or U11174 (N_11174,N_10930,N_10830);
or U11175 (N_11175,N_10830,N_10835);
and U11176 (N_11176,N_10914,N_10990);
and U11177 (N_11177,N_10869,N_10938);
xor U11178 (N_11178,N_10856,N_10848);
or U11179 (N_11179,N_10885,N_10940);
or U11180 (N_11180,N_10873,N_10935);
nand U11181 (N_11181,N_10849,N_10851);
nor U11182 (N_11182,N_10966,N_10971);
nand U11183 (N_11183,N_10898,N_10854);
xor U11184 (N_11184,N_10884,N_10860);
nor U11185 (N_11185,N_10971,N_10821);
nor U11186 (N_11186,N_10827,N_10924);
xnor U11187 (N_11187,N_10873,N_10895);
xnor U11188 (N_11188,N_10878,N_10925);
nor U11189 (N_11189,N_10976,N_10850);
and U11190 (N_11190,N_10870,N_10908);
and U11191 (N_11191,N_10945,N_10986);
xnor U11192 (N_11192,N_10847,N_10964);
xor U11193 (N_11193,N_10897,N_10990);
and U11194 (N_11194,N_10895,N_10953);
xnor U11195 (N_11195,N_10922,N_10964);
or U11196 (N_11196,N_10891,N_10933);
or U11197 (N_11197,N_10920,N_10967);
and U11198 (N_11198,N_10812,N_10883);
or U11199 (N_11199,N_10978,N_10934);
or U11200 (N_11200,N_11151,N_11091);
nand U11201 (N_11201,N_11053,N_11132);
nand U11202 (N_11202,N_11167,N_11075);
nand U11203 (N_11203,N_11142,N_11152);
nor U11204 (N_11204,N_11035,N_11155);
xor U11205 (N_11205,N_11044,N_11186);
xnor U11206 (N_11206,N_11040,N_11008);
and U11207 (N_11207,N_11062,N_11139);
nand U11208 (N_11208,N_11052,N_11161);
nand U11209 (N_11209,N_11140,N_11016);
or U11210 (N_11210,N_11094,N_11189);
or U11211 (N_11211,N_11169,N_11111);
nor U11212 (N_11212,N_11104,N_11148);
xnor U11213 (N_11213,N_11196,N_11117);
and U11214 (N_11214,N_11036,N_11128);
and U11215 (N_11215,N_11156,N_11168);
xnor U11216 (N_11216,N_11071,N_11194);
xnor U11217 (N_11217,N_11033,N_11149);
and U11218 (N_11218,N_11125,N_11025);
nor U11219 (N_11219,N_11059,N_11137);
nor U11220 (N_11220,N_11076,N_11184);
or U11221 (N_11221,N_11002,N_11090);
nand U11222 (N_11222,N_11085,N_11120);
nand U11223 (N_11223,N_11038,N_11046);
or U11224 (N_11224,N_11154,N_11123);
and U11225 (N_11225,N_11078,N_11057);
nor U11226 (N_11226,N_11107,N_11012);
and U11227 (N_11227,N_11014,N_11180);
nand U11228 (N_11228,N_11031,N_11182);
nand U11229 (N_11229,N_11150,N_11121);
or U11230 (N_11230,N_11037,N_11082);
and U11231 (N_11231,N_11122,N_11171);
nand U11232 (N_11232,N_11157,N_11198);
xor U11233 (N_11233,N_11141,N_11098);
xnor U11234 (N_11234,N_11131,N_11110);
xnor U11235 (N_11235,N_11118,N_11146);
xnor U11236 (N_11236,N_11106,N_11181);
nand U11237 (N_11237,N_11084,N_11160);
nand U11238 (N_11238,N_11003,N_11004);
or U11239 (N_11239,N_11048,N_11129);
xnor U11240 (N_11240,N_11089,N_11060);
nor U11241 (N_11241,N_11086,N_11105);
xor U11242 (N_11242,N_11135,N_11097);
xnor U11243 (N_11243,N_11049,N_11145);
nor U11244 (N_11244,N_11095,N_11092);
nor U11245 (N_11245,N_11026,N_11073);
or U11246 (N_11246,N_11176,N_11159);
xor U11247 (N_11247,N_11115,N_11191);
nand U11248 (N_11248,N_11051,N_11028);
or U11249 (N_11249,N_11039,N_11158);
nor U11250 (N_11250,N_11022,N_11018);
or U11251 (N_11251,N_11101,N_11127);
nand U11252 (N_11252,N_11175,N_11006);
nand U11253 (N_11253,N_11005,N_11056);
and U11254 (N_11254,N_11023,N_11077);
or U11255 (N_11255,N_11143,N_11126);
nor U11256 (N_11256,N_11010,N_11093);
nand U11257 (N_11257,N_11001,N_11047);
or U11258 (N_11258,N_11088,N_11113);
xor U11259 (N_11259,N_11083,N_11166);
or U11260 (N_11260,N_11177,N_11066);
or U11261 (N_11261,N_11183,N_11190);
nor U11262 (N_11262,N_11058,N_11015);
nand U11263 (N_11263,N_11112,N_11080);
and U11264 (N_11264,N_11055,N_11102);
nand U11265 (N_11265,N_11165,N_11050);
nor U11266 (N_11266,N_11172,N_11124);
nor U11267 (N_11267,N_11032,N_11069);
or U11268 (N_11268,N_11054,N_11199);
or U11269 (N_11269,N_11079,N_11087);
and U11270 (N_11270,N_11174,N_11109);
and U11271 (N_11271,N_11153,N_11013);
or U11272 (N_11272,N_11081,N_11133);
nor U11273 (N_11273,N_11136,N_11179);
nor U11274 (N_11274,N_11147,N_11063);
nand U11275 (N_11275,N_11188,N_11138);
nand U11276 (N_11276,N_11162,N_11011);
nand U11277 (N_11277,N_11185,N_11029);
or U11278 (N_11278,N_11187,N_11099);
nand U11279 (N_11279,N_11197,N_11034);
or U11280 (N_11280,N_11068,N_11192);
nand U11281 (N_11281,N_11114,N_11067);
and U11282 (N_11282,N_11024,N_11021);
nand U11283 (N_11283,N_11070,N_11027);
or U11284 (N_11284,N_11041,N_11061);
nor U11285 (N_11285,N_11009,N_11042);
nor U11286 (N_11286,N_11170,N_11108);
or U11287 (N_11287,N_11019,N_11072);
nor U11288 (N_11288,N_11178,N_11017);
nor U11289 (N_11289,N_11045,N_11096);
nor U11290 (N_11290,N_11130,N_11134);
nand U11291 (N_11291,N_11103,N_11030);
nand U11292 (N_11292,N_11119,N_11100);
nor U11293 (N_11293,N_11116,N_11193);
and U11294 (N_11294,N_11007,N_11144);
xnor U11295 (N_11295,N_11043,N_11000);
nor U11296 (N_11296,N_11164,N_11064);
nand U11297 (N_11297,N_11173,N_11163);
xnor U11298 (N_11298,N_11065,N_11020);
and U11299 (N_11299,N_11074,N_11195);
nand U11300 (N_11300,N_11167,N_11086);
nand U11301 (N_11301,N_11133,N_11089);
or U11302 (N_11302,N_11158,N_11174);
and U11303 (N_11303,N_11156,N_11047);
and U11304 (N_11304,N_11115,N_11197);
or U11305 (N_11305,N_11032,N_11064);
or U11306 (N_11306,N_11174,N_11057);
nand U11307 (N_11307,N_11090,N_11176);
nand U11308 (N_11308,N_11056,N_11126);
nor U11309 (N_11309,N_11191,N_11192);
xnor U11310 (N_11310,N_11076,N_11039);
or U11311 (N_11311,N_11057,N_11162);
or U11312 (N_11312,N_11098,N_11111);
or U11313 (N_11313,N_11057,N_11077);
nor U11314 (N_11314,N_11103,N_11150);
and U11315 (N_11315,N_11177,N_11040);
nor U11316 (N_11316,N_11062,N_11030);
and U11317 (N_11317,N_11074,N_11027);
or U11318 (N_11318,N_11015,N_11162);
or U11319 (N_11319,N_11132,N_11160);
and U11320 (N_11320,N_11071,N_11086);
nor U11321 (N_11321,N_11123,N_11078);
and U11322 (N_11322,N_11017,N_11104);
and U11323 (N_11323,N_11029,N_11155);
xnor U11324 (N_11324,N_11162,N_11140);
nor U11325 (N_11325,N_11160,N_11130);
or U11326 (N_11326,N_11118,N_11187);
nor U11327 (N_11327,N_11001,N_11161);
and U11328 (N_11328,N_11028,N_11129);
and U11329 (N_11329,N_11112,N_11186);
nor U11330 (N_11330,N_11195,N_11059);
and U11331 (N_11331,N_11060,N_11127);
and U11332 (N_11332,N_11000,N_11169);
nor U11333 (N_11333,N_11080,N_11175);
xor U11334 (N_11334,N_11081,N_11183);
or U11335 (N_11335,N_11172,N_11007);
xnor U11336 (N_11336,N_11167,N_11144);
nand U11337 (N_11337,N_11161,N_11008);
nor U11338 (N_11338,N_11163,N_11156);
xor U11339 (N_11339,N_11165,N_11024);
nand U11340 (N_11340,N_11027,N_11147);
nand U11341 (N_11341,N_11148,N_11026);
or U11342 (N_11342,N_11132,N_11042);
and U11343 (N_11343,N_11057,N_11119);
nand U11344 (N_11344,N_11182,N_11124);
nand U11345 (N_11345,N_11191,N_11159);
xnor U11346 (N_11346,N_11156,N_11029);
and U11347 (N_11347,N_11154,N_11190);
nor U11348 (N_11348,N_11167,N_11187);
nand U11349 (N_11349,N_11016,N_11006);
xnor U11350 (N_11350,N_11065,N_11090);
or U11351 (N_11351,N_11096,N_11123);
nand U11352 (N_11352,N_11126,N_11115);
xor U11353 (N_11353,N_11144,N_11057);
xnor U11354 (N_11354,N_11098,N_11156);
nand U11355 (N_11355,N_11020,N_11036);
or U11356 (N_11356,N_11173,N_11081);
nand U11357 (N_11357,N_11153,N_11105);
nand U11358 (N_11358,N_11007,N_11095);
and U11359 (N_11359,N_11018,N_11152);
or U11360 (N_11360,N_11059,N_11163);
and U11361 (N_11361,N_11023,N_11042);
and U11362 (N_11362,N_11043,N_11155);
xor U11363 (N_11363,N_11082,N_11161);
xnor U11364 (N_11364,N_11152,N_11194);
and U11365 (N_11365,N_11030,N_11198);
or U11366 (N_11366,N_11030,N_11157);
nor U11367 (N_11367,N_11020,N_11104);
or U11368 (N_11368,N_11116,N_11104);
or U11369 (N_11369,N_11179,N_11108);
xnor U11370 (N_11370,N_11135,N_11065);
nor U11371 (N_11371,N_11151,N_11188);
xor U11372 (N_11372,N_11056,N_11149);
and U11373 (N_11373,N_11015,N_11013);
xnor U11374 (N_11374,N_11116,N_11105);
and U11375 (N_11375,N_11076,N_11084);
nor U11376 (N_11376,N_11080,N_11083);
nand U11377 (N_11377,N_11097,N_11089);
and U11378 (N_11378,N_11150,N_11173);
or U11379 (N_11379,N_11143,N_11137);
xor U11380 (N_11380,N_11103,N_11121);
or U11381 (N_11381,N_11027,N_11014);
xor U11382 (N_11382,N_11027,N_11053);
and U11383 (N_11383,N_11024,N_11025);
nand U11384 (N_11384,N_11001,N_11167);
xor U11385 (N_11385,N_11020,N_11147);
xor U11386 (N_11386,N_11171,N_11199);
or U11387 (N_11387,N_11027,N_11037);
nor U11388 (N_11388,N_11162,N_11078);
xor U11389 (N_11389,N_11071,N_11054);
and U11390 (N_11390,N_11104,N_11143);
xnor U11391 (N_11391,N_11029,N_11082);
nand U11392 (N_11392,N_11009,N_11045);
xor U11393 (N_11393,N_11048,N_11135);
xnor U11394 (N_11394,N_11001,N_11063);
or U11395 (N_11395,N_11109,N_11018);
xor U11396 (N_11396,N_11172,N_11114);
and U11397 (N_11397,N_11168,N_11085);
xor U11398 (N_11398,N_11077,N_11105);
xor U11399 (N_11399,N_11024,N_11195);
or U11400 (N_11400,N_11211,N_11221);
nand U11401 (N_11401,N_11368,N_11225);
nor U11402 (N_11402,N_11207,N_11367);
and U11403 (N_11403,N_11360,N_11359);
or U11404 (N_11404,N_11245,N_11285);
nand U11405 (N_11405,N_11301,N_11380);
nor U11406 (N_11406,N_11340,N_11217);
nand U11407 (N_11407,N_11286,N_11348);
xor U11408 (N_11408,N_11292,N_11370);
xnor U11409 (N_11409,N_11297,N_11320);
nand U11410 (N_11410,N_11253,N_11226);
xnor U11411 (N_11411,N_11229,N_11357);
nand U11412 (N_11412,N_11298,N_11398);
nor U11413 (N_11413,N_11248,N_11239);
nand U11414 (N_11414,N_11377,N_11387);
nor U11415 (N_11415,N_11223,N_11375);
or U11416 (N_11416,N_11332,N_11278);
or U11417 (N_11417,N_11265,N_11318);
nor U11418 (N_11418,N_11201,N_11353);
nor U11419 (N_11419,N_11215,N_11382);
or U11420 (N_11420,N_11337,N_11365);
and U11421 (N_11421,N_11203,N_11271);
xnor U11422 (N_11422,N_11338,N_11334);
nor U11423 (N_11423,N_11237,N_11331);
and U11424 (N_11424,N_11287,N_11305);
nor U11425 (N_11425,N_11213,N_11327);
nand U11426 (N_11426,N_11308,N_11291);
nor U11427 (N_11427,N_11210,N_11351);
nor U11428 (N_11428,N_11220,N_11234);
nor U11429 (N_11429,N_11397,N_11324);
nor U11430 (N_11430,N_11208,N_11310);
nor U11431 (N_11431,N_11326,N_11346);
or U11432 (N_11432,N_11264,N_11312);
nand U11433 (N_11433,N_11344,N_11335);
or U11434 (N_11434,N_11243,N_11391);
xnor U11435 (N_11435,N_11394,N_11247);
nand U11436 (N_11436,N_11385,N_11222);
or U11437 (N_11437,N_11272,N_11325);
xor U11438 (N_11438,N_11249,N_11304);
xnor U11439 (N_11439,N_11206,N_11352);
nor U11440 (N_11440,N_11302,N_11289);
or U11441 (N_11441,N_11283,N_11315);
and U11442 (N_11442,N_11322,N_11300);
nor U11443 (N_11443,N_11233,N_11230);
or U11444 (N_11444,N_11293,N_11350);
nor U11445 (N_11445,N_11381,N_11356);
nand U11446 (N_11446,N_11307,N_11232);
nor U11447 (N_11447,N_11366,N_11294);
nand U11448 (N_11448,N_11258,N_11240);
nand U11449 (N_11449,N_11260,N_11259);
xnor U11450 (N_11450,N_11273,N_11309);
nor U11451 (N_11451,N_11256,N_11373);
nand U11452 (N_11452,N_11378,N_11333);
xor U11453 (N_11453,N_11376,N_11390);
nor U11454 (N_11454,N_11343,N_11262);
xnor U11455 (N_11455,N_11371,N_11379);
and U11456 (N_11456,N_11386,N_11336);
xor U11457 (N_11457,N_11363,N_11339);
xor U11458 (N_11458,N_11364,N_11284);
nand U11459 (N_11459,N_11231,N_11244);
and U11460 (N_11460,N_11321,N_11296);
or U11461 (N_11461,N_11374,N_11341);
xor U11462 (N_11462,N_11218,N_11227);
xor U11463 (N_11463,N_11295,N_11319);
xnor U11464 (N_11464,N_11276,N_11399);
and U11465 (N_11465,N_11242,N_11254);
xor U11466 (N_11466,N_11288,N_11358);
nand U11467 (N_11467,N_11212,N_11290);
or U11468 (N_11468,N_11268,N_11299);
nand U11469 (N_11469,N_11228,N_11257);
nor U11470 (N_11470,N_11269,N_11347);
or U11471 (N_11471,N_11349,N_11280);
xnor U11472 (N_11472,N_11388,N_11270);
nand U11473 (N_11473,N_11383,N_11219);
nor U11474 (N_11474,N_11345,N_11250);
and U11475 (N_11475,N_11252,N_11263);
or U11476 (N_11476,N_11266,N_11255);
nand U11477 (N_11477,N_11323,N_11251);
nor U11478 (N_11478,N_11204,N_11396);
and U11479 (N_11479,N_11395,N_11236);
and U11480 (N_11480,N_11361,N_11209);
and U11481 (N_11481,N_11214,N_11311);
or U11482 (N_11482,N_11216,N_11384);
and U11483 (N_11483,N_11238,N_11282);
and U11484 (N_11484,N_11275,N_11205);
nor U11485 (N_11485,N_11330,N_11328);
nor U11486 (N_11486,N_11279,N_11274);
nor U11487 (N_11487,N_11281,N_11329);
nand U11488 (N_11488,N_11200,N_11261);
xor U11489 (N_11489,N_11369,N_11277);
xnor U11490 (N_11490,N_11393,N_11313);
xnor U11491 (N_11491,N_11354,N_11392);
nor U11492 (N_11492,N_11317,N_11342);
xor U11493 (N_11493,N_11314,N_11303);
nor U11494 (N_11494,N_11316,N_11235);
nand U11495 (N_11495,N_11246,N_11267);
or U11496 (N_11496,N_11202,N_11372);
nand U11497 (N_11497,N_11362,N_11389);
nor U11498 (N_11498,N_11355,N_11306);
xor U11499 (N_11499,N_11224,N_11241);
and U11500 (N_11500,N_11262,N_11242);
nand U11501 (N_11501,N_11272,N_11210);
and U11502 (N_11502,N_11206,N_11224);
xor U11503 (N_11503,N_11387,N_11394);
and U11504 (N_11504,N_11204,N_11293);
and U11505 (N_11505,N_11288,N_11386);
and U11506 (N_11506,N_11373,N_11205);
xnor U11507 (N_11507,N_11349,N_11200);
xor U11508 (N_11508,N_11232,N_11282);
or U11509 (N_11509,N_11351,N_11310);
and U11510 (N_11510,N_11207,N_11321);
nand U11511 (N_11511,N_11358,N_11329);
or U11512 (N_11512,N_11289,N_11276);
xnor U11513 (N_11513,N_11217,N_11310);
xor U11514 (N_11514,N_11204,N_11241);
or U11515 (N_11515,N_11382,N_11260);
or U11516 (N_11516,N_11211,N_11316);
and U11517 (N_11517,N_11249,N_11203);
xnor U11518 (N_11518,N_11290,N_11331);
and U11519 (N_11519,N_11386,N_11310);
nand U11520 (N_11520,N_11314,N_11288);
or U11521 (N_11521,N_11272,N_11378);
nand U11522 (N_11522,N_11279,N_11379);
xnor U11523 (N_11523,N_11277,N_11221);
nor U11524 (N_11524,N_11256,N_11217);
and U11525 (N_11525,N_11358,N_11285);
nor U11526 (N_11526,N_11327,N_11324);
and U11527 (N_11527,N_11272,N_11285);
xor U11528 (N_11528,N_11320,N_11369);
or U11529 (N_11529,N_11259,N_11378);
or U11530 (N_11530,N_11271,N_11321);
and U11531 (N_11531,N_11315,N_11237);
xnor U11532 (N_11532,N_11354,N_11230);
nor U11533 (N_11533,N_11363,N_11359);
nand U11534 (N_11534,N_11393,N_11364);
nand U11535 (N_11535,N_11305,N_11306);
nor U11536 (N_11536,N_11318,N_11333);
nand U11537 (N_11537,N_11293,N_11385);
xnor U11538 (N_11538,N_11253,N_11228);
nand U11539 (N_11539,N_11253,N_11376);
nor U11540 (N_11540,N_11365,N_11263);
nor U11541 (N_11541,N_11215,N_11228);
and U11542 (N_11542,N_11332,N_11300);
nor U11543 (N_11543,N_11328,N_11293);
nor U11544 (N_11544,N_11364,N_11312);
nand U11545 (N_11545,N_11352,N_11245);
nor U11546 (N_11546,N_11312,N_11299);
and U11547 (N_11547,N_11354,N_11210);
xnor U11548 (N_11548,N_11316,N_11261);
and U11549 (N_11549,N_11377,N_11355);
or U11550 (N_11550,N_11258,N_11278);
nor U11551 (N_11551,N_11271,N_11380);
or U11552 (N_11552,N_11308,N_11219);
or U11553 (N_11553,N_11307,N_11224);
nor U11554 (N_11554,N_11336,N_11275);
or U11555 (N_11555,N_11231,N_11366);
and U11556 (N_11556,N_11313,N_11227);
nand U11557 (N_11557,N_11344,N_11383);
nor U11558 (N_11558,N_11290,N_11348);
and U11559 (N_11559,N_11200,N_11385);
nor U11560 (N_11560,N_11399,N_11327);
nor U11561 (N_11561,N_11279,N_11211);
nand U11562 (N_11562,N_11351,N_11307);
nand U11563 (N_11563,N_11321,N_11369);
nand U11564 (N_11564,N_11371,N_11206);
nor U11565 (N_11565,N_11346,N_11347);
and U11566 (N_11566,N_11397,N_11245);
nand U11567 (N_11567,N_11377,N_11228);
or U11568 (N_11568,N_11369,N_11377);
and U11569 (N_11569,N_11394,N_11348);
xor U11570 (N_11570,N_11301,N_11313);
or U11571 (N_11571,N_11226,N_11232);
nand U11572 (N_11572,N_11327,N_11344);
nand U11573 (N_11573,N_11326,N_11290);
xor U11574 (N_11574,N_11342,N_11325);
xor U11575 (N_11575,N_11357,N_11206);
and U11576 (N_11576,N_11379,N_11331);
xnor U11577 (N_11577,N_11315,N_11219);
and U11578 (N_11578,N_11392,N_11320);
or U11579 (N_11579,N_11355,N_11234);
and U11580 (N_11580,N_11354,N_11393);
nor U11581 (N_11581,N_11239,N_11316);
nor U11582 (N_11582,N_11308,N_11244);
or U11583 (N_11583,N_11283,N_11306);
nor U11584 (N_11584,N_11210,N_11279);
nor U11585 (N_11585,N_11264,N_11228);
or U11586 (N_11586,N_11290,N_11280);
nor U11587 (N_11587,N_11338,N_11328);
and U11588 (N_11588,N_11253,N_11316);
nor U11589 (N_11589,N_11271,N_11208);
nand U11590 (N_11590,N_11377,N_11223);
xnor U11591 (N_11591,N_11380,N_11240);
nand U11592 (N_11592,N_11216,N_11283);
or U11593 (N_11593,N_11269,N_11341);
nor U11594 (N_11594,N_11322,N_11364);
and U11595 (N_11595,N_11211,N_11385);
xor U11596 (N_11596,N_11357,N_11395);
nor U11597 (N_11597,N_11242,N_11300);
nand U11598 (N_11598,N_11244,N_11259);
nor U11599 (N_11599,N_11289,N_11382);
nand U11600 (N_11600,N_11517,N_11438);
nand U11601 (N_11601,N_11422,N_11544);
nor U11602 (N_11602,N_11597,N_11410);
nand U11603 (N_11603,N_11482,N_11546);
or U11604 (N_11604,N_11501,N_11463);
nor U11605 (N_11605,N_11508,N_11515);
nand U11606 (N_11606,N_11450,N_11568);
and U11607 (N_11607,N_11426,N_11586);
xor U11608 (N_11608,N_11486,N_11555);
nand U11609 (N_11609,N_11488,N_11441);
or U11610 (N_11610,N_11485,N_11582);
nor U11611 (N_11611,N_11417,N_11403);
and U11612 (N_11612,N_11460,N_11554);
nor U11613 (N_11613,N_11400,N_11559);
nand U11614 (N_11614,N_11551,N_11467);
nand U11615 (N_11615,N_11520,N_11500);
nor U11616 (N_11616,N_11470,N_11581);
nand U11617 (N_11617,N_11527,N_11459);
nor U11618 (N_11618,N_11475,N_11569);
nor U11619 (N_11619,N_11491,N_11447);
and U11620 (N_11620,N_11409,N_11519);
xor U11621 (N_11621,N_11537,N_11415);
nand U11622 (N_11622,N_11507,N_11522);
and U11623 (N_11623,N_11576,N_11561);
or U11624 (N_11624,N_11572,N_11549);
xor U11625 (N_11625,N_11487,N_11540);
nand U11626 (N_11626,N_11499,N_11425);
nor U11627 (N_11627,N_11436,N_11532);
xor U11628 (N_11628,N_11479,N_11404);
and U11629 (N_11629,N_11531,N_11589);
and U11630 (N_11630,N_11545,N_11455);
nor U11631 (N_11631,N_11406,N_11408);
or U11632 (N_11632,N_11502,N_11402);
or U11633 (N_11633,N_11553,N_11526);
xor U11634 (N_11634,N_11439,N_11542);
or U11635 (N_11635,N_11558,N_11543);
and U11636 (N_11636,N_11474,N_11456);
and U11637 (N_11637,N_11509,N_11413);
xor U11638 (N_11638,N_11453,N_11560);
and U11639 (N_11639,N_11483,N_11427);
nand U11640 (N_11640,N_11583,N_11504);
xor U11641 (N_11641,N_11466,N_11564);
nand U11642 (N_11642,N_11514,N_11451);
nor U11643 (N_11643,N_11433,N_11566);
or U11644 (N_11644,N_11557,N_11446);
nor U11645 (N_11645,N_11452,N_11428);
and U11646 (N_11646,N_11443,N_11496);
nor U11647 (N_11647,N_11442,N_11461);
nor U11648 (N_11648,N_11407,N_11573);
or U11649 (N_11649,N_11506,N_11574);
and U11650 (N_11650,N_11525,N_11440);
or U11651 (N_11651,N_11579,N_11599);
nor U11652 (N_11652,N_11437,N_11493);
xor U11653 (N_11653,N_11444,N_11431);
or U11654 (N_11654,N_11434,N_11510);
nor U11655 (N_11655,N_11505,N_11590);
xnor U11656 (N_11656,N_11587,N_11518);
nand U11657 (N_11657,N_11420,N_11416);
nor U11658 (N_11658,N_11480,N_11454);
and U11659 (N_11659,N_11534,N_11535);
nor U11660 (N_11660,N_11512,N_11458);
and U11661 (N_11661,N_11571,N_11412);
nor U11662 (N_11662,N_11498,N_11492);
nand U11663 (N_11663,N_11468,N_11424);
xor U11664 (N_11664,N_11473,N_11476);
and U11665 (N_11665,N_11598,N_11575);
or U11666 (N_11666,N_11414,N_11533);
nand U11667 (N_11667,N_11567,N_11464);
nand U11668 (N_11668,N_11591,N_11423);
xor U11669 (N_11669,N_11562,N_11477);
and U11670 (N_11670,N_11538,N_11578);
and U11671 (N_11671,N_11419,N_11595);
nor U11672 (N_11672,N_11580,N_11462);
and U11673 (N_11673,N_11565,N_11471);
nor U11674 (N_11674,N_11411,N_11472);
nor U11675 (N_11675,N_11405,N_11523);
nand U11676 (N_11676,N_11552,N_11490);
xnor U11677 (N_11677,N_11539,N_11593);
nor U11678 (N_11678,N_11530,N_11432);
and U11679 (N_11679,N_11541,N_11521);
or U11680 (N_11680,N_11584,N_11401);
nand U11681 (N_11681,N_11548,N_11449);
nor U11682 (N_11682,N_11516,N_11577);
or U11683 (N_11683,N_11550,N_11511);
or U11684 (N_11684,N_11497,N_11563);
xor U11685 (N_11685,N_11445,N_11457);
nand U11686 (N_11686,N_11556,N_11503);
nand U11687 (N_11687,N_11547,N_11421);
nor U11688 (N_11688,N_11478,N_11594);
or U11689 (N_11689,N_11448,N_11528);
xnor U11690 (N_11690,N_11592,N_11481);
xnor U11691 (N_11691,N_11585,N_11435);
or U11692 (N_11692,N_11570,N_11469);
and U11693 (N_11693,N_11484,N_11513);
nand U11694 (N_11694,N_11495,N_11465);
xnor U11695 (N_11695,N_11596,N_11524);
nor U11696 (N_11696,N_11430,N_11536);
nand U11697 (N_11697,N_11489,N_11588);
xnor U11698 (N_11698,N_11418,N_11429);
nor U11699 (N_11699,N_11529,N_11494);
xnor U11700 (N_11700,N_11544,N_11500);
nor U11701 (N_11701,N_11420,N_11498);
and U11702 (N_11702,N_11460,N_11472);
or U11703 (N_11703,N_11585,N_11551);
nor U11704 (N_11704,N_11583,N_11485);
or U11705 (N_11705,N_11584,N_11495);
and U11706 (N_11706,N_11502,N_11542);
and U11707 (N_11707,N_11516,N_11578);
nand U11708 (N_11708,N_11501,N_11409);
nor U11709 (N_11709,N_11515,N_11539);
or U11710 (N_11710,N_11503,N_11446);
nor U11711 (N_11711,N_11470,N_11534);
xor U11712 (N_11712,N_11552,N_11590);
nand U11713 (N_11713,N_11440,N_11452);
or U11714 (N_11714,N_11495,N_11570);
nand U11715 (N_11715,N_11585,N_11439);
nand U11716 (N_11716,N_11575,N_11538);
nand U11717 (N_11717,N_11477,N_11474);
or U11718 (N_11718,N_11496,N_11545);
nand U11719 (N_11719,N_11416,N_11508);
nand U11720 (N_11720,N_11404,N_11418);
or U11721 (N_11721,N_11520,N_11499);
nor U11722 (N_11722,N_11463,N_11478);
nor U11723 (N_11723,N_11442,N_11416);
nor U11724 (N_11724,N_11414,N_11566);
nor U11725 (N_11725,N_11565,N_11544);
nand U11726 (N_11726,N_11456,N_11531);
xor U11727 (N_11727,N_11429,N_11558);
or U11728 (N_11728,N_11534,N_11492);
nand U11729 (N_11729,N_11521,N_11554);
nand U11730 (N_11730,N_11491,N_11426);
and U11731 (N_11731,N_11410,N_11492);
and U11732 (N_11732,N_11571,N_11480);
and U11733 (N_11733,N_11538,N_11570);
and U11734 (N_11734,N_11419,N_11541);
nor U11735 (N_11735,N_11556,N_11432);
xnor U11736 (N_11736,N_11422,N_11484);
xnor U11737 (N_11737,N_11455,N_11436);
or U11738 (N_11738,N_11586,N_11441);
and U11739 (N_11739,N_11421,N_11453);
and U11740 (N_11740,N_11408,N_11508);
nor U11741 (N_11741,N_11434,N_11414);
and U11742 (N_11742,N_11550,N_11555);
nor U11743 (N_11743,N_11572,N_11543);
nand U11744 (N_11744,N_11547,N_11585);
xnor U11745 (N_11745,N_11451,N_11512);
nand U11746 (N_11746,N_11509,N_11516);
xor U11747 (N_11747,N_11428,N_11569);
or U11748 (N_11748,N_11597,N_11590);
and U11749 (N_11749,N_11561,N_11550);
nor U11750 (N_11750,N_11585,N_11517);
nor U11751 (N_11751,N_11447,N_11511);
nand U11752 (N_11752,N_11471,N_11508);
nor U11753 (N_11753,N_11405,N_11541);
xnor U11754 (N_11754,N_11503,N_11573);
nor U11755 (N_11755,N_11553,N_11444);
nand U11756 (N_11756,N_11574,N_11428);
xor U11757 (N_11757,N_11541,N_11555);
nor U11758 (N_11758,N_11437,N_11503);
nand U11759 (N_11759,N_11560,N_11521);
nand U11760 (N_11760,N_11484,N_11429);
nand U11761 (N_11761,N_11574,N_11473);
xnor U11762 (N_11762,N_11460,N_11487);
and U11763 (N_11763,N_11414,N_11471);
and U11764 (N_11764,N_11536,N_11441);
xor U11765 (N_11765,N_11567,N_11599);
or U11766 (N_11766,N_11549,N_11494);
and U11767 (N_11767,N_11597,N_11432);
xor U11768 (N_11768,N_11545,N_11498);
nand U11769 (N_11769,N_11589,N_11452);
xor U11770 (N_11770,N_11510,N_11516);
xor U11771 (N_11771,N_11581,N_11446);
or U11772 (N_11772,N_11562,N_11587);
xnor U11773 (N_11773,N_11489,N_11443);
and U11774 (N_11774,N_11433,N_11486);
nand U11775 (N_11775,N_11528,N_11596);
nand U11776 (N_11776,N_11481,N_11513);
nor U11777 (N_11777,N_11504,N_11505);
or U11778 (N_11778,N_11568,N_11589);
or U11779 (N_11779,N_11414,N_11458);
and U11780 (N_11780,N_11506,N_11534);
nor U11781 (N_11781,N_11585,N_11446);
nand U11782 (N_11782,N_11495,N_11446);
nand U11783 (N_11783,N_11517,N_11507);
or U11784 (N_11784,N_11479,N_11533);
and U11785 (N_11785,N_11410,N_11592);
nand U11786 (N_11786,N_11433,N_11569);
nand U11787 (N_11787,N_11477,N_11583);
or U11788 (N_11788,N_11512,N_11438);
or U11789 (N_11789,N_11488,N_11480);
and U11790 (N_11790,N_11591,N_11528);
xor U11791 (N_11791,N_11472,N_11437);
or U11792 (N_11792,N_11544,N_11444);
or U11793 (N_11793,N_11542,N_11511);
nor U11794 (N_11794,N_11568,N_11530);
nor U11795 (N_11795,N_11480,N_11436);
nor U11796 (N_11796,N_11488,N_11498);
or U11797 (N_11797,N_11431,N_11509);
and U11798 (N_11798,N_11403,N_11455);
and U11799 (N_11799,N_11574,N_11522);
xnor U11800 (N_11800,N_11785,N_11641);
or U11801 (N_11801,N_11625,N_11653);
and U11802 (N_11802,N_11766,N_11637);
xor U11803 (N_11803,N_11611,N_11779);
xor U11804 (N_11804,N_11697,N_11683);
xor U11805 (N_11805,N_11722,N_11782);
nor U11806 (N_11806,N_11772,N_11712);
nand U11807 (N_11807,N_11634,N_11791);
and U11808 (N_11808,N_11643,N_11601);
xnor U11809 (N_11809,N_11681,N_11620);
nand U11810 (N_11810,N_11719,N_11740);
or U11811 (N_11811,N_11796,N_11684);
and U11812 (N_11812,N_11616,N_11699);
nor U11813 (N_11813,N_11713,N_11656);
nor U11814 (N_11814,N_11728,N_11604);
and U11815 (N_11815,N_11667,N_11645);
xnor U11816 (N_11816,N_11638,N_11642);
xor U11817 (N_11817,N_11792,N_11655);
nand U11818 (N_11818,N_11778,N_11622);
or U11819 (N_11819,N_11650,N_11769);
or U11820 (N_11820,N_11659,N_11762);
nand U11821 (N_11821,N_11748,N_11703);
and U11822 (N_11822,N_11786,N_11639);
xor U11823 (N_11823,N_11714,N_11617);
or U11824 (N_11824,N_11755,N_11636);
or U11825 (N_11825,N_11709,N_11716);
nand U11826 (N_11826,N_11630,N_11672);
xor U11827 (N_11827,N_11674,N_11742);
nand U11828 (N_11828,N_11627,N_11675);
nor U11829 (N_11829,N_11759,N_11652);
nor U11830 (N_11830,N_11633,N_11734);
nand U11831 (N_11831,N_11774,N_11662);
nor U11832 (N_11832,N_11776,N_11640);
nor U11833 (N_11833,N_11665,N_11793);
nand U11834 (N_11834,N_11606,N_11790);
or U11835 (N_11835,N_11666,N_11745);
or U11836 (N_11836,N_11795,N_11789);
nand U11837 (N_11837,N_11692,N_11738);
nand U11838 (N_11838,N_11760,N_11679);
or U11839 (N_11839,N_11696,N_11600);
nand U11840 (N_11840,N_11732,N_11715);
nor U11841 (N_11841,N_11718,N_11731);
nand U11842 (N_11842,N_11635,N_11677);
or U11843 (N_11843,N_11670,N_11673);
nand U11844 (N_11844,N_11610,N_11686);
nor U11845 (N_11845,N_11767,N_11676);
and U11846 (N_11846,N_11725,N_11694);
nor U11847 (N_11847,N_11602,N_11775);
nor U11848 (N_11848,N_11629,N_11710);
nor U11849 (N_11849,N_11743,N_11626);
and U11850 (N_11850,N_11624,N_11691);
or U11851 (N_11851,N_11723,N_11729);
xnor U11852 (N_11852,N_11733,N_11707);
or U11853 (N_11853,N_11682,N_11648);
xor U11854 (N_11854,N_11680,N_11708);
and U11855 (N_11855,N_11765,N_11784);
or U11856 (N_11856,N_11720,N_11690);
nor U11857 (N_11857,N_11763,N_11717);
nor U11858 (N_11858,N_11798,N_11705);
nor U11859 (N_11859,N_11730,N_11746);
or U11860 (N_11860,N_11654,N_11615);
and U11861 (N_11861,N_11664,N_11685);
xnor U11862 (N_11862,N_11721,N_11688);
or U11863 (N_11863,N_11706,N_11661);
nor U11864 (N_11864,N_11704,N_11632);
and U11865 (N_11865,N_11618,N_11663);
or U11866 (N_11866,N_11757,N_11781);
and U11867 (N_11867,N_11770,N_11773);
or U11868 (N_11868,N_11741,N_11687);
or U11869 (N_11869,N_11711,N_11669);
xor U11870 (N_11870,N_11614,N_11780);
nor U11871 (N_11871,N_11612,N_11689);
or U11872 (N_11872,N_11644,N_11736);
nor U11873 (N_11873,N_11693,N_11651);
xnor U11874 (N_11874,N_11668,N_11701);
nand U11875 (N_11875,N_11724,N_11727);
or U11876 (N_11876,N_11756,N_11783);
nor U11877 (N_11877,N_11647,N_11771);
nor U11878 (N_11878,N_11628,N_11761);
nand U11879 (N_11879,N_11749,N_11613);
nor U11880 (N_11880,N_11764,N_11605);
nand U11881 (N_11881,N_11660,N_11754);
xnor U11882 (N_11882,N_11671,N_11768);
nor U11883 (N_11883,N_11608,N_11794);
xor U11884 (N_11884,N_11657,N_11698);
or U11885 (N_11885,N_11700,N_11726);
and U11886 (N_11886,N_11739,N_11788);
nor U11887 (N_11887,N_11737,N_11747);
and U11888 (N_11888,N_11695,N_11621);
nand U11889 (N_11889,N_11609,N_11735);
or U11890 (N_11890,N_11744,N_11619);
nor U11891 (N_11891,N_11777,N_11623);
and U11892 (N_11892,N_11799,N_11750);
and U11893 (N_11893,N_11607,N_11649);
nand U11894 (N_11894,N_11646,N_11702);
or U11895 (N_11895,N_11658,N_11631);
nor U11896 (N_11896,N_11758,N_11752);
xor U11897 (N_11897,N_11753,N_11678);
nand U11898 (N_11898,N_11751,N_11797);
or U11899 (N_11899,N_11603,N_11787);
nor U11900 (N_11900,N_11615,N_11732);
nand U11901 (N_11901,N_11635,N_11797);
xnor U11902 (N_11902,N_11672,N_11712);
or U11903 (N_11903,N_11705,N_11708);
nor U11904 (N_11904,N_11668,N_11717);
or U11905 (N_11905,N_11692,N_11753);
and U11906 (N_11906,N_11784,N_11706);
xnor U11907 (N_11907,N_11671,N_11641);
xnor U11908 (N_11908,N_11719,N_11672);
xnor U11909 (N_11909,N_11643,N_11711);
xor U11910 (N_11910,N_11653,N_11638);
and U11911 (N_11911,N_11778,N_11715);
and U11912 (N_11912,N_11733,N_11763);
xor U11913 (N_11913,N_11636,N_11746);
xor U11914 (N_11914,N_11793,N_11679);
nor U11915 (N_11915,N_11624,N_11672);
nand U11916 (N_11916,N_11739,N_11763);
xnor U11917 (N_11917,N_11643,N_11671);
xor U11918 (N_11918,N_11701,N_11698);
nand U11919 (N_11919,N_11699,N_11628);
xnor U11920 (N_11920,N_11634,N_11709);
nor U11921 (N_11921,N_11636,N_11641);
xnor U11922 (N_11922,N_11770,N_11727);
xor U11923 (N_11923,N_11609,N_11775);
or U11924 (N_11924,N_11626,N_11701);
and U11925 (N_11925,N_11712,N_11739);
and U11926 (N_11926,N_11654,N_11744);
or U11927 (N_11927,N_11632,N_11764);
nand U11928 (N_11928,N_11777,N_11736);
or U11929 (N_11929,N_11724,N_11638);
xor U11930 (N_11930,N_11770,N_11683);
xor U11931 (N_11931,N_11735,N_11785);
xor U11932 (N_11932,N_11602,N_11796);
or U11933 (N_11933,N_11644,N_11715);
xnor U11934 (N_11934,N_11621,N_11733);
and U11935 (N_11935,N_11773,N_11748);
nand U11936 (N_11936,N_11783,N_11624);
nor U11937 (N_11937,N_11622,N_11698);
xor U11938 (N_11938,N_11711,N_11739);
nor U11939 (N_11939,N_11614,N_11625);
xnor U11940 (N_11940,N_11670,N_11769);
xnor U11941 (N_11941,N_11788,N_11702);
xor U11942 (N_11942,N_11689,N_11604);
and U11943 (N_11943,N_11640,N_11628);
nor U11944 (N_11944,N_11656,N_11620);
or U11945 (N_11945,N_11618,N_11726);
and U11946 (N_11946,N_11668,N_11731);
or U11947 (N_11947,N_11740,N_11601);
or U11948 (N_11948,N_11616,N_11629);
and U11949 (N_11949,N_11694,N_11646);
xnor U11950 (N_11950,N_11765,N_11645);
nor U11951 (N_11951,N_11635,N_11642);
or U11952 (N_11952,N_11779,N_11769);
or U11953 (N_11953,N_11682,N_11696);
and U11954 (N_11954,N_11639,N_11712);
and U11955 (N_11955,N_11628,N_11614);
and U11956 (N_11956,N_11706,N_11683);
xor U11957 (N_11957,N_11726,N_11617);
and U11958 (N_11958,N_11625,N_11684);
or U11959 (N_11959,N_11632,N_11774);
xor U11960 (N_11960,N_11783,N_11627);
nor U11961 (N_11961,N_11764,N_11684);
or U11962 (N_11962,N_11600,N_11798);
nor U11963 (N_11963,N_11790,N_11622);
or U11964 (N_11964,N_11760,N_11660);
nor U11965 (N_11965,N_11667,N_11760);
and U11966 (N_11966,N_11636,N_11784);
nor U11967 (N_11967,N_11684,N_11731);
or U11968 (N_11968,N_11671,N_11793);
nor U11969 (N_11969,N_11740,N_11684);
xnor U11970 (N_11970,N_11754,N_11665);
nand U11971 (N_11971,N_11740,N_11698);
nor U11972 (N_11972,N_11659,N_11785);
xor U11973 (N_11973,N_11734,N_11636);
nand U11974 (N_11974,N_11682,N_11764);
nor U11975 (N_11975,N_11771,N_11748);
nor U11976 (N_11976,N_11607,N_11601);
or U11977 (N_11977,N_11757,N_11643);
or U11978 (N_11978,N_11616,N_11680);
and U11979 (N_11979,N_11798,N_11759);
nand U11980 (N_11980,N_11727,N_11607);
and U11981 (N_11981,N_11640,N_11704);
xor U11982 (N_11982,N_11672,N_11701);
nand U11983 (N_11983,N_11646,N_11745);
and U11984 (N_11984,N_11656,N_11714);
or U11985 (N_11985,N_11754,N_11702);
nor U11986 (N_11986,N_11676,N_11763);
xnor U11987 (N_11987,N_11709,N_11672);
and U11988 (N_11988,N_11687,N_11762);
nand U11989 (N_11989,N_11759,N_11621);
nand U11990 (N_11990,N_11718,N_11651);
nand U11991 (N_11991,N_11700,N_11703);
xor U11992 (N_11992,N_11666,N_11610);
and U11993 (N_11993,N_11619,N_11638);
nor U11994 (N_11994,N_11786,N_11743);
or U11995 (N_11995,N_11612,N_11749);
or U11996 (N_11996,N_11746,N_11760);
and U11997 (N_11997,N_11613,N_11737);
xor U11998 (N_11998,N_11689,N_11628);
or U11999 (N_11999,N_11681,N_11739);
and U12000 (N_12000,N_11943,N_11976);
nor U12001 (N_12001,N_11892,N_11858);
and U12002 (N_12002,N_11940,N_11837);
and U12003 (N_12003,N_11930,N_11872);
and U12004 (N_12004,N_11832,N_11951);
nand U12005 (N_12005,N_11908,N_11923);
nand U12006 (N_12006,N_11949,N_11914);
and U12007 (N_12007,N_11843,N_11932);
or U12008 (N_12008,N_11901,N_11912);
or U12009 (N_12009,N_11888,N_11896);
nor U12010 (N_12010,N_11829,N_11931);
nand U12011 (N_12011,N_11885,N_11835);
and U12012 (N_12012,N_11977,N_11897);
and U12013 (N_12013,N_11946,N_11957);
nand U12014 (N_12014,N_11898,N_11844);
nand U12015 (N_12015,N_11988,N_11907);
nor U12016 (N_12016,N_11864,N_11834);
and U12017 (N_12017,N_11811,N_11941);
and U12018 (N_12018,N_11814,N_11839);
nor U12019 (N_12019,N_11920,N_11953);
nor U12020 (N_12020,N_11995,N_11973);
nand U12021 (N_12021,N_11918,N_11978);
or U12022 (N_12022,N_11805,N_11960);
nor U12023 (N_12023,N_11983,N_11956);
or U12024 (N_12024,N_11803,N_11893);
nand U12025 (N_12025,N_11948,N_11827);
xor U12026 (N_12026,N_11911,N_11828);
xor U12027 (N_12027,N_11919,N_11873);
nand U12028 (N_12028,N_11959,N_11987);
nor U12029 (N_12029,N_11944,N_11821);
nand U12030 (N_12030,N_11804,N_11891);
nor U12031 (N_12031,N_11965,N_11991);
and U12032 (N_12032,N_11916,N_11840);
nand U12033 (N_12033,N_11863,N_11866);
or U12034 (N_12034,N_11871,N_11922);
xor U12035 (N_12035,N_11879,N_11971);
and U12036 (N_12036,N_11942,N_11870);
xnor U12037 (N_12037,N_11802,N_11853);
nor U12038 (N_12038,N_11842,N_11939);
nor U12039 (N_12039,N_11993,N_11927);
xor U12040 (N_12040,N_11909,N_11921);
and U12041 (N_12041,N_11851,N_11867);
nand U12042 (N_12042,N_11868,N_11852);
and U12043 (N_12043,N_11928,N_11833);
and U12044 (N_12044,N_11929,N_11817);
and U12045 (N_12045,N_11850,N_11878);
xor U12046 (N_12046,N_11859,N_11979);
nand U12047 (N_12047,N_11816,N_11974);
xor U12048 (N_12048,N_11831,N_11904);
or U12049 (N_12049,N_11876,N_11855);
nand U12050 (N_12050,N_11982,N_11926);
or U12051 (N_12051,N_11925,N_11886);
or U12052 (N_12052,N_11937,N_11854);
xnor U12053 (N_12053,N_11980,N_11913);
nand U12054 (N_12054,N_11963,N_11848);
and U12055 (N_12055,N_11985,N_11915);
nand U12056 (N_12056,N_11954,N_11883);
nand U12057 (N_12057,N_11857,N_11862);
and U12058 (N_12058,N_11836,N_11812);
nor U12059 (N_12059,N_11820,N_11903);
xor U12060 (N_12060,N_11964,N_11996);
nand U12061 (N_12061,N_11905,N_11823);
nand U12062 (N_12062,N_11967,N_11826);
xor U12063 (N_12063,N_11813,N_11970);
nor U12064 (N_12064,N_11860,N_11874);
nor U12065 (N_12065,N_11910,N_11899);
xnor U12066 (N_12066,N_11972,N_11825);
and U12067 (N_12067,N_11989,N_11845);
xor U12068 (N_12068,N_11894,N_11958);
nor U12069 (N_12069,N_11966,N_11924);
or U12070 (N_12070,N_11984,N_11881);
nor U12071 (N_12071,N_11986,N_11819);
xor U12072 (N_12072,N_11815,N_11981);
and U12073 (N_12073,N_11968,N_11887);
nand U12074 (N_12074,N_11818,N_11994);
nor U12075 (N_12075,N_11955,N_11830);
nand U12076 (N_12076,N_11869,N_11809);
or U12077 (N_12077,N_11875,N_11998);
or U12078 (N_12078,N_11841,N_11938);
and U12079 (N_12079,N_11861,N_11808);
and U12080 (N_12080,N_11952,N_11997);
xnor U12081 (N_12081,N_11884,N_11807);
or U12082 (N_12082,N_11822,N_11902);
nand U12083 (N_12083,N_11900,N_11810);
nand U12084 (N_12084,N_11849,N_11933);
nor U12085 (N_12085,N_11975,N_11877);
and U12086 (N_12086,N_11969,N_11865);
nor U12087 (N_12087,N_11846,N_11895);
or U12088 (N_12088,N_11999,N_11935);
or U12089 (N_12089,N_11882,N_11838);
nand U12090 (N_12090,N_11990,N_11806);
or U12091 (N_12091,N_11934,N_11950);
xnor U12092 (N_12092,N_11936,N_11947);
and U12093 (N_12093,N_11889,N_11906);
or U12094 (N_12094,N_11824,N_11800);
or U12095 (N_12095,N_11962,N_11847);
xor U12096 (N_12096,N_11801,N_11880);
xor U12097 (N_12097,N_11890,N_11961);
or U12098 (N_12098,N_11917,N_11992);
xor U12099 (N_12099,N_11856,N_11945);
xor U12100 (N_12100,N_11889,N_11802);
nor U12101 (N_12101,N_11915,N_11858);
nor U12102 (N_12102,N_11834,N_11987);
nor U12103 (N_12103,N_11977,N_11908);
nand U12104 (N_12104,N_11913,N_11886);
and U12105 (N_12105,N_11872,N_11889);
xor U12106 (N_12106,N_11824,N_11972);
nand U12107 (N_12107,N_11800,N_11980);
and U12108 (N_12108,N_11889,N_11927);
nor U12109 (N_12109,N_11801,N_11851);
nor U12110 (N_12110,N_11908,N_11915);
nand U12111 (N_12111,N_11889,N_11820);
and U12112 (N_12112,N_11987,N_11864);
or U12113 (N_12113,N_11855,N_11916);
and U12114 (N_12114,N_11993,N_11998);
nor U12115 (N_12115,N_11824,N_11842);
and U12116 (N_12116,N_11899,N_11813);
or U12117 (N_12117,N_11839,N_11976);
nand U12118 (N_12118,N_11922,N_11937);
xnor U12119 (N_12119,N_11938,N_11845);
nor U12120 (N_12120,N_11898,N_11880);
and U12121 (N_12121,N_11950,N_11889);
xor U12122 (N_12122,N_11976,N_11954);
nand U12123 (N_12123,N_11910,N_11941);
and U12124 (N_12124,N_11828,N_11926);
and U12125 (N_12125,N_11868,N_11910);
xor U12126 (N_12126,N_11809,N_11831);
or U12127 (N_12127,N_11986,N_11949);
xnor U12128 (N_12128,N_11885,N_11807);
or U12129 (N_12129,N_11858,N_11881);
nor U12130 (N_12130,N_11968,N_11877);
and U12131 (N_12131,N_11907,N_11894);
nand U12132 (N_12132,N_11971,N_11985);
and U12133 (N_12133,N_11813,N_11841);
and U12134 (N_12134,N_11817,N_11941);
xor U12135 (N_12135,N_11959,N_11878);
xor U12136 (N_12136,N_11804,N_11834);
nand U12137 (N_12137,N_11972,N_11935);
or U12138 (N_12138,N_11956,N_11917);
nand U12139 (N_12139,N_11892,N_11977);
or U12140 (N_12140,N_11931,N_11839);
nor U12141 (N_12141,N_11933,N_11996);
nor U12142 (N_12142,N_11875,N_11952);
or U12143 (N_12143,N_11959,N_11912);
nor U12144 (N_12144,N_11849,N_11870);
and U12145 (N_12145,N_11992,N_11974);
xnor U12146 (N_12146,N_11957,N_11997);
xor U12147 (N_12147,N_11816,N_11822);
nor U12148 (N_12148,N_11960,N_11935);
xnor U12149 (N_12149,N_11997,N_11919);
xnor U12150 (N_12150,N_11821,N_11990);
xnor U12151 (N_12151,N_11981,N_11946);
nand U12152 (N_12152,N_11875,N_11904);
nand U12153 (N_12153,N_11999,N_11879);
xnor U12154 (N_12154,N_11918,N_11931);
and U12155 (N_12155,N_11929,N_11855);
or U12156 (N_12156,N_11980,N_11928);
nor U12157 (N_12157,N_11819,N_11961);
nand U12158 (N_12158,N_11846,N_11809);
xnor U12159 (N_12159,N_11888,N_11881);
or U12160 (N_12160,N_11964,N_11909);
nor U12161 (N_12161,N_11928,N_11853);
xor U12162 (N_12162,N_11826,N_11985);
or U12163 (N_12163,N_11863,N_11893);
or U12164 (N_12164,N_11851,N_11885);
or U12165 (N_12165,N_11876,N_11877);
and U12166 (N_12166,N_11824,N_11969);
nand U12167 (N_12167,N_11960,N_11892);
and U12168 (N_12168,N_11921,N_11868);
nor U12169 (N_12169,N_11941,N_11931);
nor U12170 (N_12170,N_11800,N_11953);
xnor U12171 (N_12171,N_11804,N_11920);
xnor U12172 (N_12172,N_11998,N_11810);
nand U12173 (N_12173,N_11861,N_11823);
or U12174 (N_12174,N_11961,N_11971);
or U12175 (N_12175,N_11969,N_11971);
nand U12176 (N_12176,N_11866,N_11824);
nor U12177 (N_12177,N_11884,N_11816);
and U12178 (N_12178,N_11956,N_11958);
nand U12179 (N_12179,N_11898,N_11913);
and U12180 (N_12180,N_11982,N_11814);
or U12181 (N_12181,N_11872,N_11870);
nor U12182 (N_12182,N_11963,N_11937);
nor U12183 (N_12183,N_11894,N_11984);
or U12184 (N_12184,N_11928,N_11911);
and U12185 (N_12185,N_11881,N_11882);
and U12186 (N_12186,N_11902,N_11881);
or U12187 (N_12187,N_11878,N_11967);
and U12188 (N_12188,N_11842,N_11846);
or U12189 (N_12189,N_11963,N_11928);
xnor U12190 (N_12190,N_11900,N_11975);
or U12191 (N_12191,N_11926,N_11943);
or U12192 (N_12192,N_11966,N_11800);
or U12193 (N_12193,N_11982,N_11818);
xnor U12194 (N_12194,N_11800,N_11979);
and U12195 (N_12195,N_11978,N_11931);
nor U12196 (N_12196,N_11831,N_11882);
and U12197 (N_12197,N_11863,N_11977);
and U12198 (N_12198,N_11870,N_11805);
and U12199 (N_12199,N_11850,N_11920);
and U12200 (N_12200,N_12011,N_12036);
nand U12201 (N_12201,N_12168,N_12024);
and U12202 (N_12202,N_12062,N_12006);
xnor U12203 (N_12203,N_12100,N_12161);
nand U12204 (N_12204,N_12003,N_12194);
or U12205 (N_12205,N_12061,N_12163);
nand U12206 (N_12206,N_12067,N_12107);
xor U12207 (N_12207,N_12099,N_12090);
nand U12208 (N_12208,N_12127,N_12010);
or U12209 (N_12209,N_12129,N_12094);
or U12210 (N_12210,N_12130,N_12178);
nand U12211 (N_12211,N_12095,N_12116);
or U12212 (N_12212,N_12073,N_12049);
or U12213 (N_12213,N_12113,N_12064);
nand U12214 (N_12214,N_12088,N_12172);
nand U12215 (N_12215,N_12066,N_12187);
nand U12216 (N_12216,N_12111,N_12158);
and U12217 (N_12217,N_12152,N_12193);
and U12218 (N_12218,N_12125,N_12176);
nor U12219 (N_12219,N_12023,N_12124);
nand U12220 (N_12220,N_12189,N_12026);
xnor U12221 (N_12221,N_12145,N_12171);
xnor U12222 (N_12222,N_12005,N_12004);
or U12223 (N_12223,N_12001,N_12119);
nand U12224 (N_12224,N_12112,N_12179);
nor U12225 (N_12225,N_12008,N_12195);
nor U12226 (N_12226,N_12013,N_12177);
xor U12227 (N_12227,N_12173,N_12136);
and U12228 (N_12228,N_12051,N_12022);
nand U12229 (N_12229,N_12123,N_12019);
nor U12230 (N_12230,N_12121,N_12105);
or U12231 (N_12231,N_12078,N_12033);
nand U12232 (N_12232,N_12184,N_12077);
and U12233 (N_12233,N_12043,N_12052);
nor U12234 (N_12234,N_12082,N_12079);
nand U12235 (N_12235,N_12159,N_12138);
nand U12236 (N_12236,N_12012,N_12057);
nor U12237 (N_12237,N_12154,N_12035);
xor U12238 (N_12238,N_12137,N_12044);
nand U12239 (N_12239,N_12092,N_12083);
xor U12240 (N_12240,N_12086,N_12118);
and U12241 (N_12241,N_12048,N_12128);
xnor U12242 (N_12242,N_12115,N_12108);
nor U12243 (N_12243,N_12150,N_12147);
nor U12244 (N_12244,N_12030,N_12196);
nand U12245 (N_12245,N_12153,N_12096);
and U12246 (N_12246,N_12198,N_12183);
and U12247 (N_12247,N_12149,N_12175);
nor U12248 (N_12248,N_12182,N_12007);
nand U12249 (N_12249,N_12072,N_12143);
nor U12250 (N_12250,N_12018,N_12160);
nand U12251 (N_12251,N_12188,N_12040);
or U12252 (N_12252,N_12055,N_12089);
nand U12253 (N_12253,N_12166,N_12041);
or U12254 (N_12254,N_12032,N_12144);
and U12255 (N_12255,N_12038,N_12191);
and U12256 (N_12256,N_12091,N_12098);
nand U12257 (N_12257,N_12148,N_12065);
nand U12258 (N_12258,N_12021,N_12039);
nor U12259 (N_12259,N_12131,N_12157);
xor U12260 (N_12260,N_12053,N_12027);
nand U12261 (N_12261,N_12047,N_12106);
or U12262 (N_12262,N_12142,N_12190);
or U12263 (N_12263,N_12110,N_12000);
and U12264 (N_12264,N_12059,N_12063);
nor U12265 (N_12265,N_12139,N_12014);
and U12266 (N_12266,N_12084,N_12164);
or U12267 (N_12267,N_12141,N_12122);
or U12268 (N_12268,N_12140,N_12169);
and U12269 (N_12269,N_12034,N_12133);
or U12270 (N_12270,N_12080,N_12103);
nor U12271 (N_12271,N_12134,N_12146);
or U12272 (N_12272,N_12085,N_12156);
nand U12273 (N_12273,N_12025,N_12031);
nor U12274 (N_12274,N_12028,N_12015);
nor U12275 (N_12275,N_12155,N_12069);
and U12276 (N_12276,N_12017,N_12132);
nor U12277 (N_12277,N_12037,N_12104);
or U12278 (N_12278,N_12093,N_12185);
xnor U12279 (N_12279,N_12109,N_12135);
and U12280 (N_12280,N_12192,N_12002);
or U12281 (N_12281,N_12174,N_12101);
xnor U12282 (N_12282,N_12058,N_12102);
and U12283 (N_12283,N_12199,N_12197);
and U12284 (N_12284,N_12170,N_12070);
nand U12285 (N_12285,N_12009,N_12056);
xor U12286 (N_12286,N_12120,N_12126);
or U12287 (N_12287,N_12162,N_12114);
nand U12288 (N_12288,N_12165,N_12087);
xor U12289 (N_12289,N_12097,N_12071);
xnor U12290 (N_12290,N_12151,N_12186);
xnor U12291 (N_12291,N_12180,N_12181);
and U12292 (N_12292,N_12060,N_12117);
nand U12293 (N_12293,N_12020,N_12167);
nor U12294 (N_12294,N_12054,N_12050);
and U12295 (N_12295,N_12029,N_12046);
nor U12296 (N_12296,N_12074,N_12076);
xnor U12297 (N_12297,N_12042,N_12075);
or U12298 (N_12298,N_12045,N_12016);
nand U12299 (N_12299,N_12081,N_12068);
nand U12300 (N_12300,N_12184,N_12036);
or U12301 (N_12301,N_12009,N_12042);
xor U12302 (N_12302,N_12115,N_12039);
or U12303 (N_12303,N_12049,N_12006);
nor U12304 (N_12304,N_12073,N_12199);
or U12305 (N_12305,N_12064,N_12162);
nor U12306 (N_12306,N_12080,N_12038);
and U12307 (N_12307,N_12084,N_12064);
xnor U12308 (N_12308,N_12009,N_12023);
and U12309 (N_12309,N_12077,N_12100);
nor U12310 (N_12310,N_12090,N_12045);
nand U12311 (N_12311,N_12074,N_12090);
xnor U12312 (N_12312,N_12197,N_12163);
xor U12313 (N_12313,N_12079,N_12100);
nor U12314 (N_12314,N_12059,N_12000);
or U12315 (N_12315,N_12092,N_12068);
and U12316 (N_12316,N_12066,N_12189);
nand U12317 (N_12317,N_12199,N_12084);
and U12318 (N_12318,N_12054,N_12040);
nand U12319 (N_12319,N_12056,N_12125);
nand U12320 (N_12320,N_12056,N_12005);
xnor U12321 (N_12321,N_12063,N_12144);
or U12322 (N_12322,N_12072,N_12175);
or U12323 (N_12323,N_12107,N_12098);
nand U12324 (N_12324,N_12038,N_12066);
and U12325 (N_12325,N_12145,N_12009);
and U12326 (N_12326,N_12160,N_12012);
nand U12327 (N_12327,N_12089,N_12194);
xnor U12328 (N_12328,N_12103,N_12160);
xor U12329 (N_12329,N_12141,N_12124);
nand U12330 (N_12330,N_12069,N_12138);
nor U12331 (N_12331,N_12121,N_12195);
and U12332 (N_12332,N_12062,N_12031);
nor U12333 (N_12333,N_12153,N_12165);
nand U12334 (N_12334,N_12024,N_12016);
or U12335 (N_12335,N_12188,N_12004);
and U12336 (N_12336,N_12148,N_12163);
or U12337 (N_12337,N_12045,N_12014);
nor U12338 (N_12338,N_12094,N_12078);
nor U12339 (N_12339,N_12136,N_12094);
nand U12340 (N_12340,N_12077,N_12008);
nand U12341 (N_12341,N_12052,N_12166);
or U12342 (N_12342,N_12099,N_12170);
nor U12343 (N_12343,N_12100,N_12011);
nand U12344 (N_12344,N_12092,N_12091);
and U12345 (N_12345,N_12124,N_12047);
or U12346 (N_12346,N_12003,N_12100);
nand U12347 (N_12347,N_12085,N_12192);
nor U12348 (N_12348,N_12181,N_12040);
or U12349 (N_12349,N_12193,N_12067);
nor U12350 (N_12350,N_12144,N_12080);
xor U12351 (N_12351,N_12148,N_12081);
nand U12352 (N_12352,N_12094,N_12159);
or U12353 (N_12353,N_12111,N_12094);
nor U12354 (N_12354,N_12166,N_12118);
nor U12355 (N_12355,N_12112,N_12049);
nor U12356 (N_12356,N_12077,N_12119);
nor U12357 (N_12357,N_12024,N_12000);
nor U12358 (N_12358,N_12004,N_12055);
and U12359 (N_12359,N_12092,N_12163);
nand U12360 (N_12360,N_12114,N_12168);
nor U12361 (N_12361,N_12005,N_12026);
nor U12362 (N_12362,N_12021,N_12185);
xnor U12363 (N_12363,N_12145,N_12051);
xor U12364 (N_12364,N_12154,N_12087);
and U12365 (N_12365,N_12085,N_12009);
nor U12366 (N_12366,N_12145,N_12113);
nand U12367 (N_12367,N_12067,N_12018);
or U12368 (N_12368,N_12190,N_12179);
and U12369 (N_12369,N_12004,N_12135);
nor U12370 (N_12370,N_12133,N_12171);
or U12371 (N_12371,N_12162,N_12072);
and U12372 (N_12372,N_12047,N_12064);
nor U12373 (N_12373,N_12053,N_12077);
xnor U12374 (N_12374,N_12137,N_12049);
or U12375 (N_12375,N_12015,N_12170);
and U12376 (N_12376,N_12014,N_12195);
nand U12377 (N_12377,N_12027,N_12052);
or U12378 (N_12378,N_12114,N_12090);
or U12379 (N_12379,N_12116,N_12014);
nor U12380 (N_12380,N_12072,N_12166);
and U12381 (N_12381,N_12159,N_12019);
nor U12382 (N_12382,N_12095,N_12114);
or U12383 (N_12383,N_12040,N_12094);
xor U12384 (N_12384,N_12010,N_12068);
xor U12385 (N_12385,N_12037,N_12135);
nand U12386 (N_12386,N_12021,N_12150);
and U12387 (N_12387,N_12129,N_12032);
nand U12388 (N_12388,N_12149,N_12189);
nand U12389 (N_12389,N_12187,N_12064);
nor U12390 (N_12390,N_12119,N_12097);
or U12391 (N_12391,N_12180,N_12169);
and U12392 (N_12392,N_12036,N_12177);
nor U12393 (N_12393,N_12050,N_12191);
xor U12394 (N_12394,N_12096,N_12024);
nor U12395 (N_12395,N_12181,N_12013);
and U12396 (N_12396,N_12016,N_12144);
nor U12397 (N_12397,N_12141,N_12144);
or U12398 (N_12398,N_12041,N_12175);
nor U12399 (N_12399,N_12189,N_12085);
and U12400 (N_12400,N_12342,N_12202);
nor U12401 (N_12401,N_12244,N_12363);
nor U12402 (N_12402,N_12323,N_12224);
and U12403 (N_12403,N_12227,N_12313);
nand U12404 (N_12404,N_12294,N_12357);
nand U12405 (N_12405,N_12246,N_12365);
nor U12406 (N_12406,N_12254,N_12325);
or U12407 (N_12407,N_12364,N_12328);
nor U12408 (N_12408,N_12374,N_12265);
xnor U12409 (N_12409,N_12211,N_12281);
nor U12410 (N_12410,N_12303,N_12214);
nor U12411 (N_12411,N_12308,N_12274);
nor U12412 (N_12412,N_12355,N_12228);
nand U12413 (N_12413,N_12330,N_12384);
or U12414 (N_12414,N_12215,N_12208);
or U12415 (N_12415,N_12286,N_12379);
nor U12416 (N_12416,N_12229,N_12234);
or U12417 (N_12417,N_12306,N_12268);
nor U12418 (N_12418,N_12368,N_12337);
or U12419 (N_12419,N_12247,N_12322);
and U12420 (N_12420,N_12235,N_12280);
xor U12421 (N_12421,N_12329,N_12387);
nand U12422 (N_12422,N_12319,N_12372);
and U12423 (N_12423,N_12282,N_12395);
nor U12424 (N_12424,N_12257,N_12315);
xor U12425 (N_12425,N_12200,N_12207);
nand U12426 (N_12426,N_12255,N_12333);
or U12427 (N_12427,N_12301,N_12361);
xnor U12428 (N_12428,N_12290,N_12292);
nand U12429 (N_12429,N_12339,N_12230);
or U12430 (N_12430,N_12375,N_12206);
nor U12431 (N_12431,N_12344,N_12204);
nand U12432 (N_12432,N_12307,N_12237);
xnor U12433 (N_12433,N_12213,N_12334);
nand U12434 (N_12434,N_12277,N_12356);
nand U12435 (N_12435,N_12284,N_12381);
or U12436 (N_12436,N_12219,N_12296);
xnor U12437 (N_12437,N_12350,N_12391);
and U12438 (N_12438,N_12271,N_12270);
nand U12439 (N_12439,N_12222,N_12242);
and U12440 (N_12440,N_12351,N_12305);
nand U12441 (N_12441,N_12309,N_12348);
or U12442 (N_12442,N_12226,N_12248);
or U12443 (N_12443,N_12253,N_12297);
xor U12444 (N_12444,N_12311,N_12392);
xnor U12445 (N_12445,N_12338,N_12203);
and U12446 (N_12446,N_12373,N_12288);
and U12447 (N_12447,N_12335,N_12295);
or U12448 (N_12448,N_12376,N_12209);
or U12449 (N_12449,N_12367,N_12398);
or U12450 (N_12450,N_12359,N_12336);
xor U12451 (N_12451,N_12318,N_12261);
nand U12452 (N_12452,N_12287,N_12302);
nor U12453 (N_12453,N_12217,N_12304);
nor U12454 (N_12454,N_12279,N_12238);
nand U12455 (N_12455,N_12298,N_12272);
or U12456 (N_12456,N_12347,N_12201);
or U12457 (N_12457,N_12377,N_12331);
xor U12458 (N_12458,N_12273,N_12251);
nand U12459 (N_12459,N_12397,N_12383);
nand U12460 (N_12460,N_12324,N_12386);
xnor U12461 (N_12461,N_12220,N_12316);
or U12462 (N_12462,N_12341,N_12378);
nor U12463 (N_12463,N_12266,N_12314);
nand U12464 (N_12464,N_12396,N_12276);
and U12465 (N_12465,N_12382,N_12267);
nor U12466 (N_12466,N_12216,N_12249);
or U12467 (N_12467,N_12326,N_12252);
xor U12468 (N_12468,N_12346,N_12293);
nor U12469 (N_12469,N_12320,N_12299);
xnor U12470 (N_12470,N_12380,N_12362);
or U12471 (N_12471,N_12232,N_12218);
and U12472 (N_12472,N_12240,N_12260);
and U12473 (N_12473,N_12370,N_12353);
xnor U12474 (N_12474,N_12256,N_12394);
nor U12475 (N_12475,N_12236,N_12233);
nand U12476 (N_12476,N_12262,N_12289);
nand U12477 (N_12477,N_12221,N_12366);
and U12478 (N_12478,N_12278,N_12352);
xor U12479 (N_12479,N_12345,N_12285);
nand U12480 (N_12480,N_12239,N_12358);
xnor U12481 (N_12481,N_12317,N_12321);
or U12482 (N_12482,N_12263,N_12332);
xor U12483 (N_12483,N_12369,N_12360);
xor U12484 (N_12484,N_12310,N_12399);
and U12485 (N_12485,N_12388,N_12212);
xor U12486 (N_12486,N_12259,N_12258);
xnor U12487 (N_12487,N_12371,N_12340);
and U12488 (N_12488,N_12245,N_12225);
or U12489 (N_12489,N_12205,N_12354);
and U12490 (N_12490,N_12243,N_12291);
nor U12491 (N_12491,N_12264,N_12393);
nor U12492 (N_12492,N_12343,N_12385);
nand U12493 (N_12493,N_12349,N_12250);
xnor U12494 (N_12494,N_12390,N_12327);
nand U12495 (N_12495,N_12283,N_12300);
and U12496 (N_12496,N_12223,N_12389);
and U12497 (N_12497,N_12269,N_12312);
xnor U12498 (N_12498,N_12241,N_12231);
xor U12499 (N_12499,N_12210,N_12275);
and U12500 (N_12500,N_12350,N_12332);
and U12501 (N_12501,N_12279,N_12347);
xor U12502 (N_12502,N_12216,N_12259);
and U12503 (N_12503,N_12377,N_12394);
xnor U12504 (N_12504,N_12252,N_12254);
or U12505 (N_12505,N_12217,N_12254);
xnor U12506 (N_12506,N_12335,N_12286);
nor U12507 (N_12507,N_12395,N_12292);
nor U12508 (N_12508,N_12389,N_12307);
and U12509 (N_12509,N_12227,N_12339);
nand U12510 (N_12510,N_12340,N_12329);
nor U12511 (N_12511,N_12305,N_12304);
nand U12512 (N_12512,N_12286,N_12337);
xor U12513 (N_12513,N_12362,N_12363);
nor U12514 (N_12514,N_12234,N_12300);
nor U12515 (N_12515,N_12283,N_12252);
or U12516 (N_12516,N_12329,N_12242);
xor U12517 (N_12517,N_12320,N_12343);
or U12518 (N_12518,N_12362,N_12285);
or U12519 (N_12519,N_12266,N_12303);
or U12520 (N_12520,N_12367,N_12375);
or U12521 (N_12521,N_12364,N_12296);
and U12522 (N_12522,N_12375,N_12326);
xnor U12523 (N_12523,N_12349,N_12395);
nand U12524 (N_12524,N_12382,N_12346);
xor U12525 (N_12525,N_12364,N_12331);
nand U12526 (N_12526,N_12224,N_12221);
nand U12527 (N_12527,N_12245,N_12381);
xor U12528 (N_12528,N_12399,N_12376);
and U12529 (N_12529,N_12236,N_12322);
xnor U12530 (N_12530,N_12339,N_12374);
nor U12531 (N_12531,N_12398,N_12357);
xnor U12532 (N_12532,N_12323,N_12381);
nor U12533 (N_12533,N_12309,N_12326);
and U12534 (N_12534,N_12364,N_12345);
nor U12535 (N_12535,N_12251,N_12399);
xnor U12536 (N_12536,N_12383,N_12385);
nor U12537 (N_12537,N_12243,N_12275);
nor U12538 (N_12538,N_12366,N_12392);
xnor U12539 (N_12539,N_12308,N_12271);
or U12540 (N_12540,N_12235,N_12396);
or U12541 (N_12541,N_12366,N_12214);
and U12542 (N_12542,N_12344,N_12374);
or U12543 (N_12543,N_12238,N_12240);
nor U12544 (N_12544,N_12375,N_12351);
nand U12545 (N_12545,N_12349,N_12234);
nand U12546 (N_12546,N_12258,N_12215);
nand U12547 (N_12547,N_12319,N_12320);
or U12548 (N_12548,N_12236,N_12303);
nor U12549 (N_12549,N_12303,N_12356);
and U12550 (N_12550,N_12233,N_12222);
and U12551 (N_12551,N_12387,N_12374);
and U12552 (N_12552,N_12323,N_12341);
nand U12553 (N_12553,N_12354,N_12345);
nand U12554 (N_12554,N_12265,N_12395);
or U12555 (N_12555,N_12324,N_12319);
xor U12556 (N_12556,N_12344,N_12360);
nor U12557 (N_12557,N_12316,N_12318);
nand U12558 (N_12558,N_12317,N_12339);
or U12559 (N_12559,N_12211,N_12341);
and U12560 (N_12560,N_12286,N_12361);
or U12561 (N_12561,N_12387,N_12305);
or U12562 (N_12562,N_12314,N_12221);
nand U12563 (N_12563,N_12344,N_12244);
nand U12564 (N_12564,N_12375,N_12317);
nor U12565 (N_12565,N_12225,N_12293);
nor U12566 (N_12566,N_12350,N_12235);
nor U12567 (N_12567,N_12336,N_12253);
and U12568 (N_12568,N_12271,N_12322);
nand U12569 (N_12569,N_12399,N_12345);
or U12570 (N_12570,N_12347,N_12283);
and U12571 (N_12571,N_12256,N_12288);
and U12572 (N_12572,N_12220,N_12318);
xor U12573 (N_12573,N_12381,N_12318);
nand U12574 (N_12574,N_12217,N_12353);
and U12575 (N_12575,N_12274,N_12255);
nand U12576 (N_12576,N_12340,N_12207);
and U12577 (N_12577,N_12384,N_12236);
and U12578 (N_12578,N_12288,N_12215);
nor U12579 (N_12579,N_12264,N_12243);
or U12580 (N_12580,N_12289,N_12274);
and U12581 (N_12581,N_12360,N_12308);
and U12582 (N_12582,N_12383,N_12245);
and U12583 (N_12583,N_12212,N_12312);
xnor U12584 (N_12584,N_12214,N_12388);
and U12585 (N_12585,N_12367,N_12258);
nand U12586 (N_12586,N_12390,N_12310);
xor U12587 (N_12587,N_12258,N_12395);
or U12588 (N_12588,N_12305,N_12346);
and U12589 (N_12589,N_12363,N_12257);
xnor U12590 (N_12590,N_12207,N_12360);
or U12591 (N_12591,N_12336,N_12301);
nor U12592 (N_12592,N_12381,N_12340);
nor U12593 (N_12593,N_12366,N_12243);
or U12594 (N_12594,N_12364,N_12313);
and U12595 (N_12595,N_12369,N_12390);
nand U12596 (N_12596,N_12302,N_12325);
nor U12597 (N_12597,N_12349,N_12289);
xor U12598 (N_12598,N_12270,N_12220);
nor U12599 (N_12599,N_12336,N_12270);
and U12600 (N_12600,N_12571,N_12542);
xor U12601 (N_12601,N_12451,N_12434);
and U12602 (N_12602,N_12465,N_12579);
nand U12603 (N_12603,N_12507,N_12510);
and U12604 (N_12604,N_12461,N_12544);
and U12605 (N_12605,N_12456,N_12531);
nand U12606 (N_12606,N_12538,N_12404);
nand U12607 (N_12607,N_12508,N_12445);
nand U12608 (N_12608,N_12532,N_12432);
xnor U12609 (N_12609,N_12592,N_12479);
or U12610 (N_12610,N_12554,N_12535);
xnor U12611 (N_12611,N_12526,N_12567);
nand U12612 (N_12612,N_12521,N_12541);
nor U12613 (N_12613,N_12599,N_12488);
or U12614 (N_12614,N_12486,N_12517);
nor U12615 (N_12615,N_12509,N_12444);
nor U12616 (N_12616,N_12454,N_12401);
nor U12617 (N_12617,N_12413,N_12522);
xnor U12618 (N_12618,N_12437,N_12481);
or U12619 (N_12619,N_12424,N_12408);
nor U12620 (N_12620,N_12406,N_12566);
or U12621 (N_12621,N_12573,N_12426);
nand U12622 (N_12622,N_12474,N_12411);
nand U12623 (N_12623,N_12559,N_12588);
nand U12624 (N_12624,N_12466,N_12568);
nand U12625 (N_12625,N_12598,N_12491);
nand U12626 (N_12626,N_12419,N_12484);
xor U12627 (N_12627,N_12500,N_12405);
and U12628 (N_12628,N_12492,N_12436);
and U12629 (N_12629,N_12540,N_12476);
xnor U12630 (N_12630,N_12543,N_12412);
nand U12631 (N_12631,N_12525,N_12447);
or U12632 (N_12632,N_12504,N_12418);
or U12633 (N_12633,N_12572,N_12511);
nand U12634 (N_12634,N_12414,N_12530);
nor U12635 (N_12635,N_12452,N_12450);
nor U12636 (N_12636,N_12443,N_12410);
or U12637 (N_12637,N_12528,N_12519);
or U12638 (N_12638,N_12583,N_12478);
and U12639 (N_12639,N_12514,N_12428);
or U12640 (N_12640,N_12417,N_12503);
nor U12641 (N_12641,N_12487,N_12576);
and U12642 (N_12642,N_12471,N_12529);
nor U12643 (N_12643,N_12427,N_12597);
or U12644 (N_12644,N_12595,N_12473);
and U12645 (N_12645,N_12455,N_12558);
nand U12646 (N_12646,N_12497,N_12448);
and U12647 (N_12647,N_12552,N_12470);
nor U12648 (N_12648,N_12520,N_12593);
or U12649 (N_12649,N_12489,N_12555);
nor U12650 (N_12650,N_12537,N_12464);
nor U12651 (N_12651,N_12581,N_12490);
nand U12652 (N_12652,N_12409,N_12459);
nor U12653 (N_12653,N_12446,N_12533);
and U12654 (N_12654,N_12400,N_12547);
nor U12655 (N_12655,N_12578,N_12524);
nor U12656 (N_12656,N_12506,N_12560);
nand U12657 (N_12657,N_12498,N_12587);
or U12658 (N_12658,N_12527,N_12402);
and U12659 (N_12659,N_12562,N_12467);
or U12660 (N_12660,N_12591,N_12403);
nand U12661 (N_12661,N_12539,N_12439);
xor U12662 (N_12662,N_12570,N_12416);
and U12663 (N_12663,N_12512,N_12423);
xnor U12664 (N_12664,N_12556,N_12441);
and U12665 (N_12665,N_12457,N_12546);
nand U12666 (N_12666,N_12548,N_12574);
xor U12667 (N_12667,N_12516,N_12577);
and U12668 (N_12668,N_12586,N_12545);
xor U12669 (N_12669,N_12483,N_12569);
or U12670 (N_12670,N_12429,N_12433);
and U12671 (N_12671,N_12463,N_12553);
nor U12672 (N_12672,N_12590,N_12458);
xor U12673 (N_12673,N_12496,N_12442);
or U12674 (N_12674,N_12440,N_12420);
or U12675 (N_12675,N_12523,N_12563);
or U12676 (N_12676,N_12493,N_12462);
and U12677 (N_12677,N_12460,N_12580);
xor U12678 (N_12678,N_12449,N_12515);
or U12679 (N_12679,N_12584,N_12551);
or U12680 (N_12680,N_12453,N_12407);
or U12681 (N_12681,N_12485,N_12534);
and U12682 (N_12682,N_12518,N_12477);
xor U12683 (N_12683,N_12575,N_12425);
or U12684 (N_12684,N_12589,N_12501);
or U12685 (N_12685,N_12438,N_12505);
and U12686 (N_12686,N_12582,N_12585);
and U12687 (N_12687,N_12561,N_12430);
or U12688 (N_12688,N_12536,N_12565);
xnor U12689 (N_12689,N_12594,N_12469);
nand U12690 (N_12690,N_12468,N_12431);
nand U12691 (N_12691,N_12494,N_12472);
and U12692 (N_12692,N_12513,N_12482);
and U12693 (N_12693,N_12564,N_12549);
nor U12694 (N_12694,N_12502,N_12415);
nor U12695 (N_12695,N_12475,N_12435);
or U12696 (N_12696,N_12421,N_12550);
nand U12697 (N_12697,N_12480,N_12422);
nand U12698 (N_12698,N_12557,N_12495);
nor U12699 (N_12699,N_12499,N_12596);
nand U12700 (N_12700,N_12440,N_12407);
nor U12701 (N_12701,N_12448,N_12502);
and U12702 (N_12702,N_12549,N_12583);
and U12703 (N_12703,N_12469,N_12426);
nand U12704 (N_12704,N_12598,N_12507);
nor U12705 (N_12705,N_12581,N_12428);
nand U12706 (N_12706,N_12490,N_12551);
and U12707 (N_12707,N_12561,N_12470);
xor U12708 (N_12708,N_12546,N_12420);
xor U12709 (N_12709,N_12546,N_12411);
nand U12710 (N_12710,N_12583,N_12537);
and U12711 (N_12711,N_12580,N_12437);
nor U12712 (N_12712,N_12409,N_12515);
nor U12713 (N_12713,N_12558,N_12487);
or U12714 (N_12714,N_12516,N_12401);
nor U12715 (N_12715,N_12454,N_12403);
and U12716 (N_12716,N_12433,N_12589);
or U12717 (N_12717,N_12590,N_12574);
or U12718 (N_12718,N_12447,N_12464);
and U12719 (N_12719,N_12576,N_12409);
or U12720 (N_12720,N_12519,N_12475);
and U12721 (N_12721,N_12474,N_12470);
nand U12722 (N_12722,N_12494,N_12508);
xnor U12723 (N_12723,N_12505,N_12428);
or U12724 (N_12724,N_12503,N_12500);
xor U12725 (N_12725,N_12427,N_12562);
and U12726 (N_12726,N_12448,N_12473);
and U12727 (N_12727,N_12427,N_12430);
nor U12728 (N_12728,N_12555,N_12564);
or U12729 (N_12729,N_12442,N_12521);
and U12730 (N_12730,N_12598,N_12590);
and U12731 (N_12731,N_12449,N_12498);
and U12732 (N_12732,N_12481,N_12579);
nand U12733 (N_12733,N_12472,N_12420);
or U12734 (N_12734,N_12555,N_12401);
xnor U12735 (N_12735,N_12510,N_12500);
xnor U12736 (N_12736,N_12422,N_12471);
or U12737 (N_12737,N_12459,N_12577);
nand U12738 (N_12738,N_12505,N_12500);
and U12739 (N_12739,N_12469,N_12401);
and U12740 (N_12740,N_12448,N_12508);
xnor U12741 (N_12741,N_12564,N_12544);
or U12742 (N_12742,N_12504,N_12498);
xor U12743 (N_12743,N_12448,N_12451);
nor U12744 (N_12744,N_12592,N_12551);
nor U12745 (N_12745,N_12522,N_12458);
nor U12746 (N_12746,N_12584,N_12496);
nor U12747 (N_12747,N_12526,N_12599);
and U12748 (N_12748,N_12447,N_12433);
nand U12749 (N_12749,N_12429,N_12565);
or U12750 (N_12750,N_12514,N_12498);
xnor U12751 (N_12751,N_12430,N_12412);
nor U12752 (N_12752,N_12450,N_12444);
or U12753 (N_12753,N_12418,N_12422);
xnor U12754 (N_12754,N_12503,N_12493);
xnor U12755 (N_12755,N_12530,N_12534);
and U12756 (N_12756,N_12442,N_12569);
xnor U12757 (N_12757,N_12430,N_12506);
xor U12758 (N_12758,N_12531,N_12493);
xnor U12759 (N_12759,N_12407,N_12481);
or U12760 (N_12760,N_12493,N_12582);
xor U12761 (N_12761,N_12557,N_12597);
and U12762 (N_12762,N_12500,N_12508);
xor U12763 (N_12763,N_12593,N_12430);
xnor U12764 (N_12764,N_12536,N_12593);
xnor U12765 (N_12765,N_12477,N_12428);
xnor U12766 (N_12766,N_12572,N_12514);
nor U12767 (N_12767,N_12449,N_12517);
xor U12768 (N_12768,N_12516,N_12419);
and U12769 (N_12769,N_12476,N_12534);
nand U12770 (N_12770,N_12419,N_12503);
or U12771 (N_12771,N_12553,N_12485);
and U12772 (N_12772,N_12522,N_12516);
or U12773 (N_12773,N_12538,N_12428);
or U12774 (N_12774,N_12583,N_12429);
nor U12775 (N_12775,N_12577,N_12569);
nand U12776 (N_12776,N_12545,N_12477);
and U12777 (N_12777,N_12575,N_12522);
nor U12778 (N_12778,N_12519,N_12400);
and U12779 (N_12779,N_12509,N_12461);
xor U12780 (N_12780,N_12561,N_12567);
nand U12781 (N_12781,N_12465,N_12433);
nand U12782 (N_12782,N_12424,N_12504);
xor U12783 (N_12783,N_12575,N_12544);
and U12784 (N_12784,N_12562,N_12465);
or U12785 (N_12785,N_12464,N_12555);
or U12786 (N_12786,N_12536,N_12578);
xor U12787 (N_12787,N_12522,N_12523);
and U12788 (N_12788,N_12473,N_12507);
or U12789 (N_12789,N_12420,N_12417);
and U12790 (N_12790,N_12593,N_12560);
nor U12791 (N_12791,N_12556,N_12422);
nor U12792 (N_12792,N_12482,N_12406);
xnor U12793 (N_12793,N_12498,N_12437);
nor U12794 (N_12794,N_12509,N_12563);
or U12795 (N_12795,N_12576,N_12527);
xnor U12796 (N_12796,N_12571,N_12589);
or U12797 (N_12797,N_12465,N_12595);
xnor U12798 (N_12798,N_12445,N_12439);
nor U12799 (N_12799,N_12550,N_12469);
and U12800 (N_12800,N_12671,N_12773);
nand U12801 (N_12801,N_12790,N_12645);
xor U12802 (N_12802,N_12661,N_12759);
xnor U12803 (N_12803,N_12735,N_12750);
or U12804 (N_12804,N_12670,N_12751);
nor U12805 (N_12805,N_12799,N_12611);
and U12806 (N_12806,N_12730,N_12682);
and U12807 (N_12807,N_12641,N_12777);
and U12808 (N_12808,N_12640,N_12795);
nor U12809 (N_12809,N_12711,N_12692);
nor U12810 (N_12810,N_12685,N_12679);
nor U12811 (N_12811,N_12728,N_12787);
or U12812 (N_12812,N_12717,N_12713);
nand U12813 (N_12813,N_12697,N_12747);
nor U12814 (N_12814,N_12667,N_12631);
nand U12815 (N_12815,N_12740,N_12690);
xor U12816 (N_12816,N_12616,N_12742);
nor U12817 (N_12817,N_12792,N_12624);
xor U12818 (N_12818,N_12648,N_12786);
or U12819 (N_12819,N_12788,N_12673);
nand U12820 (N_12820,N_12691,N_12714);
nor U12821 (N_12821,N_12638,N_12783);
nor U12822 (N_12822,N_12748,N_12703);
xor U12823 (N_12823,N_12652,N_12604);
nor U12824 (N_12824,N_12789,N_12676);
nand U12825 (N_12825,N_12665,N_12681);
xor U12826 (N_12826,N_12608,N_12791);
nor U12827 (N_12827,N_12776,N_12694);
nor U12828 (N_12828,N_12708,N_12724);
or U12829 (N_12829,N_12601,N_12774);
and U12830 (N_12830,N_12672,N_12757);
xor U12831 (N_12831,N_12745,N_12693);
nand U12832 (N_12832,N_12636,N_12744);
xnor U12833 (N_12833,N_12705,N_12754);
xnor U12834 (N_12834,N_12619,N_12736);
and U12835 (N_12835,N_12621,N_12687);
xor U12836 (N_12836,N_12626,N_12769);
or U12837 (N_12837,N_12796,N_12606);
nor U12838 (N_12838,N_12746,N_12635);
nor U12839 (N_12839,N_12675,N_12605);
or U12840 (N_12840,N_12674,N_12755);
nor U12841 (N_12841,N_12770,N_12763);
nor U12842 (N_12842,N_12775,N_12729);
nor U12843 (N_12843,N_12739,N_12700);
or U12844 (N_12844,N_12753,N_12632);
and U12845 (N_12845,N_12732,N_12756);
or U12846 (N_12846,N_12743,N_12686);
xnor U12847 (N_12847,N_12722,N_12761);
and U12848 (N_12848,N_12760,N_12678);
or U12849 (N_12849,N_12710,N_12752);
xor U12850 (N_12850,N_12680,N_12643);
and U12851 (N_12851,N_12781,N_12651);
and U12852 (N_12852,N_12649,N_12704);
nand U12853 (N_12853,N_12749,N_12771);
and U12854 (N_12854,N_12772,N_12620);
xnor U12855 (N_12855,N_12656,N_12737);
and U12856 (N_12856,N_12660,N_12603);
nand U12857 (N_12857,N_12662,N_12612);
and U12858 (N_12858,N_12706,N_12718);
nand U12859 (N_12859,N_12764,N_12684);
nor U12860 (N_12860,N_12609,N_12627);
or U12861 (N_12861,N_12758,N_12654);
nor U12862 (N_12862,N_12666,N_12699);
or U12863 (N_12863,N_12600,N_12629);
and U12864 (N_12864,N_12653,N_12785);
or U12865 (N_12865,N_12625,N_12634);
nand U12866 (N_12866,N_12657,N_12683);
and U12867 (N_12867,N_12793,N_12655);
nor U12868 (N_12868,N_12765,N_12669);
nand U12869 (N_12869,N_12779,N_12727);
nand U12870 (N_12870,N_12628,N_12695);
and U12871 (N_12871,N_12658,N_12659);
xor U12872 (N_12872,N_12668,N_12702);
xor U12873 (N_12873,N_12725,N_12613);
nor U12874 (N_12874,N_12782,N_12610);
nor U12875 (N_12875,N_12707,N_12650);
or U12876 (N_12876,N_12794,N_12698);
nor U12877 (N_12877,N_12642,N_12623);
nor U12878 (N_12878,N_12639,N_12721);
nand U12879 (N_12879,N_12712,N_12738);
nor U12880 (N_12880,N_12646,N_12630);
xnor U12881 (N_12881,N_12715,N_12647);
xor U12882 (N_12882,N_12726,N_12677);
or U12883 (N_12883,N_12766,N_12767);
xor U12884 (N_12884,N_12696,N_12720);
and U12885 (N_12885,N_12797,N_12731);
nor U12886 (N_12886,N_12633,N_12637);
nor U12887 (N_12887,N_12784,N_12618);
nand U12888 (N_12888,N_12688,N_12768);
and U12889 (N_12889,N_12664,N_12622);
and U12890 (N_12890,N_12607,N_12614);
nor U12891 (N_12891,N_12762,N_12709);
nand U12892 (N_12892,N_12716,N_12798);
nor U12893 (N_12893,N_12723,N_12701);
and U12894 (N_12894,N_12741,N_12602);
nor U12895 (N_12895,N_12615,N_12778);
nand U12896 (N_12896,N_12644,N_12780);
xor U12897 (N_12897,N_12663,N_12689);
or U12898 (N_12898,N_12719,N_12734);
or U12899 (N_12899,N_12733,N_12617);
nand U12900 (N_12900,N_12733,N_12721);
and U12901 (N_12901,N_12749,N_12730);
xor U12902 (N_12902,N_12766,N_12776);
nand U12903 (N_12903,N_12795,N_12645);
nand U12904 (N_12904,N_12719,N_12644);
and U12905 (N_12905,N_12747,N_12795);
or U12906 (N_12906,N_12666,N_12601);
nand U12907 (N_12907,N_12712,N_12614);
or U12908 (N_12908,N_12648,N_12701);
xnor U12909 (N_12909,N_12777,N_12620);
xnor U12910 (N_12910,N_12751,N_12720);
nor U12911 (N_12911,N_12617,N_12773);
xnor U12912 (N_12912,N_12674,N_12611);
xnor U12913 (N_12913,N_12703,N_12754);
and U12914 (N_12914,N_12726,N_12670);
nand U12915 (N_12915,N_12663,N_12798);
or U12916 (N_12916,N_12683,N_12637);
and U12917 (N_12917,N_12650,N_12796);
nand U12918 (N_12918,N_12763,N_12725);
xnor U12919 (N_12919,N_12743,N_12670);
nand U12920 (N_12920,N_12759,N_12650);
nand U12921 (N_12921,N_12639,N_12650);
nand U12922 (N_12922,N_12736,N_12655);
xnor U12923 (N_12923,N_12640,N_12722);
or U12924 (N_12924,N_12776,N_12789);
nand U12925 (N_12925,N_12629,N_12731);
nor U12926 (N_12926,N_12697,N_12675);
nor U12927 (N_12927,N_12657,N_12679);
nor U12928 (N_12928,N_12734,N_12601);
and U12929 (N_12929,N_12785,N_12637);
nor U12930 (N_12930,N_12795,N_12699);
and U12931 (N_12931,N_12694,N_12770);
and U12932 (N_12932,N_12661,N_12608);
or U12933 (N_12933,N_12675,N_12754);
nand U12934 (N_12934,N_12677,N_12651);
and U12935 (N_12935,N_12792,N_12649);
nand U12936 (N_12936,N_12640,N_12775);
and U12937 (N_12937,N_12645,N_12763);
nand U12938 (N_12938,N_12795,N_12694);
or U12939 (N_12939,N_12713,N_12663);
and U12940 (N_12940,N_12683,N_12628);
xor U12941 (N_12941,N_12646,N_12652);
and U12942 (N_12942,N_12776,N_12780);
nor U12943 (N_12943,N_12743,N_12620);
nand U12944 (N_12944,N_12766,N_12659);
and U12945 (N_12945,N_12761,N_12673);
xor U12946 (N_12946,N_12714,N_12776);
nor U12947 (N_12947,N_12607,N_12620);
or U12948 (N_12948,N_12747,N_12631);
and U12949 (N_12949,N_12615,N_12765);
xor U12950 (N_12950,N_12600,N_12704);
nor U12951 (N_12951,N_12775,N_12711);
xor U12952 (N_12952,N_12799,N_12692);
and U12953 (N_12953,N_12786,N_12711);
xnor U12954 (N_12954,N_12764,N_12786);
nand U12955 (N_12955,N_12616,N_12782);
nor U12956 (N_12956,N_12629,N_12640);
nor U12957 (N_12957,N_12660,N_12677);
or U12958 (N_12958,N_12609,N_12732);
nand U12959 (N_12959,N_12674,N_12793);
or U12960 (N_12960,N_12789,N_12748);
nand U12961 (N_12961,N_12727,N_12624);
and U12962 (N_12962,N_12662,N_12614);
or U12963 (N_12963,N_12777,N_12665);
nand U12964 (N_12964,N_12761,N_12671);
or U12965 (N_12965,N_12619,N_12727);
nor U12966 (N_12966,N_12651,N_12730);
xor U12967 (N_12967,N_12644,N_12726);
or U12968 (N_12968,N_12682,N_12792);
or U12969 (N_12969,N_12661,N_12760);
and U12970 (N_12970,N_12789,N_12651);
and U12971 (N_12971,N_12767,N_12605);
or U12972 (N_12972,N_12764,N_12667);
nand U12973 (N_12973,N_12668,N_12628);
or U12974 (N_12974,N_12701,N_12782);
and U12975 (N_12975,N_12625,N_12797);
xnor U12976 (N_12976,N_12635,N_12780);
and U12977 (N_12977,N_12798,N_12747);
or U12978 (N_12978,N_12712,N_12743);
or U12979 (N_12979,N_12658,N_12643);
and U12980 (N_12980,N_12646,N_12775);
nor U12981 (N_12981,N_12795,N_12622);
xnor U12982 (N_12982,N_12650,N_12636);
nor U12983 (N_12983,N_12697,N_12737);
xnor U12984 (N_12984,N_12638,N_12671);
and U12985 (N_12985,N_12755,N_12702);
and U12986 (N_12986,N_12746,N_12696);
or U12987 (N_12987,N_12719,N_12689);
nor U12988 (N_12988,N_12707,N_12663);
nand U12989 (N_12989,N_12683,N_12631);
xor U12990 (N_12990,N_12757,N_12743);
nor U12991 (N_12991,N_12794,N_12676);
nand U12992 (N_12992,N_12615,N_12777);
or U12993 (N_12993,N_12613,N_12732);
and U12994 (N_12994,N_12699,N_12698);
and U12995 (N_12995,N_12738,N_12700);
xor U12996 (N_12996,N_12657,N_12694);
nand U12997 (N_12997,N_12686,N_12737);
or U12998 (N_12998,N_12684,N_12689);
and U12999 (N_12999,N_12730,N_12741);
and U13000 (N_13000,N_12907,N_12997);
nor U13001 (N_13001,N_12949,N_12956);
xor U13002 (N_13002,N_12849,N_12817);
nand U13003 (N_13003,N_12958,N_12940);
or U13004 (N_13004,N_12923,N_12964);
nand U13005 (N_13005,N_12827,N_12912);
or U13006 (N_13006,N_12843,N_12976);
and U13007 (N_13007,N_12813,N_12806);
nand U13008 (N_13008,N_12820,N_12910);
nor U13009 (N_13009,N_12874,N_12993);
and U13010 (N_13010,N_12946,N_12819);
and U13011 (N_13011,N_12848,N_12953);
nor U13012 (N_13012,N_12800,N_12971);
nand U13013 (N_13013,N_12860,N_12870);
and U13014 (N_13014,N_12954,N_12866);
xor U13015 (N_13015,N_12879,N_12886);
and U13016 (N_13016,N_12965,N_12995);
or U13017 (N_13017,N_12810,N_12927);
or U13018 (N_13018,N_12939,N_12852);
nand U13019 (N_13019,N_12893,N_12994);
nand U13020 (N_13020,N_12839,N_12804);
and U13021 (N_13021,N_12890,N_12805);
nand U13022 (N_13022,N_12877,N_12983);
nand U13023 (N_13023,N_12845,N_12826);
xnor U13024 (N_13024,N_12986,N_12957);
xor U13025 (N_13025,N_12926,N_12815);
nand U13026 (N_13026,N_12811,N_12873);
nor U13027 (N_13027,N_12809,N_12967);
and U13028 (N_13028,N_12865,N_12854);
and U13029 (N_13029,N_12981,N_12841);
and U13030 (N_13030,N_12937,N_12867);
nand U13031 (N_13031,N_12858,N_12833);
and U13032 (N_13032,N_12821,N_12931);
xor U13033 (N_13033,N_12896,N_12835);
and U13034 (N_13034,N_12919,N_12970);
xnor U13035 (N_13035,N_12978,N_12934);
nand U13036 (N_13036,N_12960,N_12948);
and U13037 (N_13037,N_12984,N_12911);
or U13038 (N_13038,N_12928,N_12853);
or U13039 (N_13039,N_12807,N_12880);
and U13040 (N_13040,N_12812,N_12889);
nand U13041 (N_13041,N_12938,N_12961);
and U13042 (N_13042,N_12876,N_12972);
nor U13043 (N_13043,N_12918,N_12840);
nor U13044 (N_13044,N_12851,N_12861);
nor U13045 (N_13045,N_12917,N_12908);
nand U13046 (N_13046,N_12905,N_12999);
or U13047 (N_13047,N_12888,N_12823);
and U13048 (N_13048,N_12900,N_12902);
and U13049 (N_13049,N_12882,N_12885);
xor U13050 (N_13050,N_12904,N_12925);
nand U13051 (N_13051,N_12901,N_12950);
xnor U13052 (N_13052,N_12977,N_12913);
or U13053 (N_13053,N_12868,N_12871);
or U13054 (N_13054,N_12844,N_12996);
xnor U13055 (N_13055,N_12990,N_12929);
xnor U13056 (N_13056,N_12836,N_12824);
nand U13057 (N_13057,N_12920,N_12822);
or U13058 (N_13058,N_12985,N_12982);
and U13059 (N_13059,N_12899,N_12855);
nor U13060 (N_13060,N_12837,N_12859);
or U13061 (N_13061,N_12872,N_12969);
xnor U13062 (N_13062,N_12916,N_12869);
and U13063 (N_13063,N_12915,N_12959);
nor U13064 (N_13064,N_12987,N_12862);
and U13065 (N_13065,N_12830,N_12942);
xor U13066 (N_13066,N_12979,N_12856);
and U13067 (N_13067,N_12975,N_12850);
nor U13068 (N_13068,N_12814,N_12903);
or U13069 (N_13069,N_12842,N_12992);
and U13070 (N_13070,N_12966,N_12947);
nor U13071 (N_13071,N_12943,N_12921);
or U13072 (N_13072,N_12924,N_12909);
nand U13073 (N_13073,N_12828,N_12933);
nor U13074 (N_13074,N_12895,N_12825);
xnor U13075 (N_13075,N_12930,N_12831);
and U13076 (N_13076,N_12898,N_12952);
and U13077 (N_13077,N_12936,N_12878);
xor U13078 (N_13078,N_12801,N_12832);
nor U13079 (N_13079,N_12847,N_12881);
nor U13080 (N_13080,N_12891,N_12818);
and U13081 (N_13081,N_12991,N_12864);
nand U13082 (N_13082,N_12973,N_12884);
or U13083 (N_13083,N_12894,N_12951);
and U13084 (N_13084,N_12829,N_12892);
and U13085 (N_13085,N_12980,N_12955);
xor U13086 (N_13086,N_12846,N_12887);
or U13087 (N_13087,N_12963,N_12883);
nor U13088 (N_13088,N_12857,N_12914);
nor U13089 (N_13089,N_12998,N_12906);
xor U13090 (N_13090,N_12803,N_12922);
xor U13091 (N_13091,N_12875,N_12932);
and U13092 (N_13092,N_12802,N_12944);
or U13093 (N_13093,N_12863,N_12834);
or U13094 (N_13094,N_12962,N_12935);
and U13095 (N_13095,N_12816,N_12974);
or U13096 (N_13096,N_12989,N_12838);
nor U13097 (N_13097,N_12945,N_12808);
or U13098 (N_13098,N_12968,N_12988);
xor U13099 (N_13099,N_12897,N_12941);
xnor U13100 (N_13100,N_12911,N_12924);
and U13101 (N_13101,N_12987,N_12893);
nand U13102 (N_13102,N_12841,N_12859);
and U13103 (N_13103,N_12923,N_12984);
nor U13104 (N_13104,N_12812,N_12893);
xnor U13105 (N_13105,N_12911,N_12801);
or U13106 (N_13106,N_12896,N_12894);
nand U13107 (N_13107,N_12826,N_12931);
xnor U13108 (N_13108,N_12947,N_12990);
nor U13109 (N_13109,N_12952,N_12957);
nand U13110 (N_13110,N_12932,N_12953);
and U13111 (N_13111,N_12807,N_12822);
and U13112 (N_13112,N_12963,N_12801);
xnor U13113 (N_13113,N_12914,N_12957);
nor U13114 (N_13114,N_12992,N_12803);
xnor U13115 (N_13115,N_12807,N_12892);
xor U13116 (N_13116,N_12875,N_12985);
nor U13117 (N_13117,N_12914,N_12900);
nor U13118 (N_13118,N_12945,N_12817);
xnor U13119 (N_13119,N_12963,N_12856);
or U13120 (N_13120,N_12945,N_12871);
xor U13121 (N_13121,N_12880,N_12988);
nand U13122 (N_13122,N_12952,N_12949);
or U13123 (N_13123,N_12891,N_12811);
and U13124 (N_13124,N_12824,N_12829);
nand U13125 (N_13125,N_12819,N_12907);
or U13126 (N_13126,N_12905,N_12980);
and U13127 (N_13127,N_12837,N_12913);
nor U13128 (N_13128,N_12847,N_12831);
nor U13129 (N_13129,N_12910,N_12998);
nor U13130 (N_13130,N_12962,N_12864);
nor U13131 (N_13131,N_12806,N_12953);
or U13132 (N_13132,N_12932,N_12945);
xnor U13133 (N_13133,N_12927,N_12944);
or U13134 (N_13134,N_12968,N_12972);
and U13135 (N_13135,N_12933,N_12835);
nor U13136 (N_13136,N_12819,N_12961);
nor U13137 (N_13137,N_12935,N_12937);
xnor U13138 (N_13138,N_12988,N_12838);
and U13139 (N_13139,N_12948,N_12900);
nand U13140 (N_13140,N_12893,N_12899);
nand U13141 (N_13141,N_12854,N_12931);
and U13142 (N_13142,N_12904,N_12895);
nand U13143 (N_13143,N_12861,N_12887);
nand U13144 (N_13144,N_12935,N_12914);
xnor U13145 (N_13145,N_12999,N_12959);
and U13146 (N_13146,N_12822,N_12884);
xnor U13147 (N_13147,N_12908,N_12901);
or U13148 (N_13148,N_12859,N_12930);
nor U13149 (N_13149,N_12866,N_12895);
or U13150 (N_13150,N_12838,N_12987);
or U13151 (N_13151,N_12863,N_12812);
or U13152 (N_13152,N_12978,N_12809);
nand U13153 (N_13153,N_12903,N_12921);
and U13154 (N_13154,N_12899,N_12863);
xnor U13155 (N_13155,N_12893,N_12859);
nand U13156 (N_13156,N_12938,N_12823);
xnor U13157 (N_13157,N_12815,N_12937);
xor U13158 (N_13158,N_12942,N_12950);
nor U13159 (N_13159,N_12827,N_12987);
and U13160 (N_13160,N_12868,N_12846);
nand U13161 (N_13161,N_12921,N_12938);
xnor U13162 (N_13162,N_12912,N_12908);
nor U13163 (N_13163,N_12883,N_12958);
xnor U13164 (N_13164,N_12978,N_12922);
and U13165 (N_13165,N_12805,N_12853);
nand U13166 (N_13166,N_12990,N_12820);
or U13167 (N_13167,N_12900,N_12907);
and U13168 (N_13168,N_12813,N_12881);
and U13169 (N_13169,N_12996,N_12801);
and U13170 (N_13170,N_12830,N_12996);
nand U13171 (N_13171,N_12932,N_12994);
nor U13172 (N_13172,N_12916,N_12881);
xnor U13173 (N_13173,N_12819,N_12854);
and U13174 (N_13174,N_12825,N_12858);
xnor U13175 (N_13175,N_12846,N_12922);
and U13176 (N_13176,N_12923,N_12845);
or U13177 (N_13177,N_12981,N_12902);
or U13178 (N_13178,N_12982,N_12986);
and U13179 (N_13179,N_12949,N_12928);
and U13180 (N_13180,N_12897,N_12994);
or U13181 (N_13181,N_12878,N_12822);
and U13182 (N_13182,N_12944,N_12961);
or U13183 (N_13183,N_12984,N_12838);
or U13184 (N_13184,N_12813,N_12872);
xor U13185 (N_13185,N_12828,N_12923);
nand U13186 (N_13186,N_12807,N_12928);
or U13187 (N_13187,N_12906,N_12956);
nand U13188 (N_13188,N_12929,N_12849);
nand U13189 (N_13189,N_12856,N_12968);
nor U13190 (N_13190,N_12946,N_12955);
or U13191 (N_13191,N_12937,N_12981);
or U13192 (N_13192,N_12964,N_12867);
and U13193 (N_13193,N_12933,N_12802);
xor U13194 (N_13194,N_12833,N_12975);
xnor U13195 (N_13195,N_12965,N_12876);
xnor U13196 (N_13196,N_12994,N_12813);
nor U13197 (N_13197,N_12865,N_12809);
and U13198 (N_13198,N_12808,N_12995);
or U13199 (N_13199,N_12956,N_12802);
xnor U13200 (N_13200,N_13169,N_13140);
xor U13201 (N_13201,N_13133,N_13021);
and U13202 (N_13202,N_13058,N_13009);
nand U13203 (N_13203,N_13109,N_13024);
and U13204 (N_13204,N_13172,N_13026);
or U13205 (N_13205,N_13086,N_13182);
nor U13206 (N_13206,N_13114,N_13106);
nand U13207 (N_13207,N_13118,N_13078);
xnor U13208 (N_13208,N_13127,N_13096);
nand U13209 (N_13209,N_13197,N_13089);
nand U13210 (N_13210,N_13038,N_13168);
or U13211 (N_13211,N_13023,N_13069);
and U13212 (N_13212,N_13068,N_13156);
nor U13213 (N_13213,N_13130,N_13084);
xnor U13214 (N_13214,N_13049,N_13035);
and U13215 (N_13215,N_13176,N_13150);
nor U13216 (N_13216,N_13159,N_13076);
nand U13217 (N_13217,N_13022,N_13187);
nor U13218 (N_13218,N_13161,N_13011);
and U13219 (N_13219,N_13020,N_13042);
or U13220 (N_13220,N_13163,N_13093);
and U13221 (N_13221,N_13134,N_13074);
xor U13222 (N_13222,N_13046,N_13015);
or U13223 (N_13223,N_13010,N_13087);
and U13224 (N_13224,N_13094,N_13122);
and U13225 (N_13225,N_13029,N_13157);
xnor U13226 (N_13226,N_13119,N_13128);
nor U13227 (N_13227,N_13132,N_13162);
and U13228 (N_13228,N_13097,N_13018);
and U13229 (N_13229,N_13137,N_13085);
nor U13230 (N_13230,N_13057,N_13198);
nor U13231 (N_13231,N_13177,N_13174);
xnor U13232 (N_13232,N_13158,N_13129);
nor U13233 (N_13233,N_13194,N_13185);
nand U13234 (N_13234,N_13007,N_13017);
xnor U13235 (N_13235,N_13062,N_13103);
and U13236 (N_13236,N_13091,N_13173);
xor U13237 (N_13237,N_13070,N_13110);
or U13238 (N_13238,N_13165,N_13080);
nand U13239 (N_13239,N_13193,N_13039);
nand U13240 (N_13240,N_13120,N_13148);
and U13241 (N_13241,N_13167,N_13183);
nand U13242 (N_13242,N_13008,N_13092);
nand U13243 (N_13243,N_13048,N_13044);
nand U13244 (N_13244,N_13190,N_13065);
nand U13245 (N_13245,N_13144,N_13051);
nand U13246 (N_13246,N_13012,N_13112);
and U13247 (N_13247,N_13082,N_13151);
or U13248 (N_13248,N_13045,N_13164);
nor U13249 (N_13249,N_13126,N_13125);
nand U13250 (N_13250,N_13003,N_13180);
or U13251 (N_13251,N_13145,N_13079);
nand U13252 (N_13252,N_13066,N_13032);
nand U13253 (N_13253,N_13095,N_13027);
xor U13254 (N_13254,N_13013,N_13090);
nor U13255 (N_13255,N_13192,N_13104);
and U13256 (N_13256,N_13107,N_13199);
xnor U13257 (N_13257,N_13131,N_13072);
and U13258 (N_13258,N_13178,N_13195);
xor U13259 (N_13259,N_13153,N_13138);
xor U13260 (N_13260,N_13099,N_13041);
nor U13261 (N_13261,N_13077,N_13073);
or U13262 (N_13262,N_13191,N_13031);
nor U13263 (N_13263,N_13054,N_13184);
nor U13264 (N_13264,N_13100,N_13111);
nor U13265 (N_13265,N_13047,N_13083);
nand U13266 (N_13266,N_13059,N_13034);
and U13267 (N_13267,N_13124,N_13101);
or U13268 (N_13268,N_13037,N_13115);
or U13269 (N_13269,N_13141,N_13006);
nand U13270 (N_13270,N_13102,N_13116);
nor U13271 (N_13271,N_13188,N_13001);
or U13272 (N_13272,N_13067,N_13075);
nor U13273 (N_13273,N_13108,N_13033);
nand U13274 (N_13274,N_13117,N_13060);
nand U13275 (N_13275,N_13028,N_13146);
and U13276 (N_13276,N_13189,N_13170);
or U13277 (N_13277,N_13071,N_13136);
and U13278 (N_13278,N_13030,N_13000);
or U13279 (N_13279,N_13121,N_13105);
or U13280 (N_13280,N_13181,N_13142);
xnor U13281 (N_13281,N_13186,N_13160);
and U13282 (N_13282,N_13043,N_13004);
nand U13283 (N_13283,N_13016,N_13061);
or U13284 (N_13284,N_13149,N_13139);
xnor U13285 (N_13285,N_13053,N_13175);
nand U13286 (N_13286,N_13196,N_13040);
nand U13287 (N_13287,N_13147,N_13171);
or U13288 (N_13288,N_13052,N_13154);
nand U13289 (N_13289,N_13056,N_13135);
and U13290 (N_13290,N_13019,N_13064);
nor U13291 (N_13291,N_13025,N_13179);
and U13292 (N_13292,N_13050,N_13063);
or U13293 (N_13293,N_13143,N_13166);
or U13294 (N_13294,N_13081,N_13002);
and U13295 (N_13295,N_13155,N_13005);
nand U13296 (N_13296,N_13088,N_13113);
xor U13297 (N_13297,N_13036,N_13152);
nor U13298 (N_13298,N_13123,N_13014);
nor U13299 (N_13299,N_13098,N_13055);
xor U13300 (N_13300,N_13187,N_13095);
xor U13301 (N_13301,N_13002,N_13155);
and U13302 (N_13302,N_13191,N_13148);
and U13303 (N_13303,N_13174,N_13028);
nor U13304 (N_13304,N_13164,N_13097);
or U13305 (N_13305,N_13022,N_13166);
nand U13306 (N_13306,N_13059,N_13136);
and U13307 (N_13307,N_13089,N_13069);
or U13308 (N_13308,N_13177,N_13019);
nor U13309 (N_13309,N_13182,N_13090);
nand U13310 (N_13310,N_13148,N_13144);
xor U13311 (N_13311,N_13086,N_13063);
nand U13312 (N_13312,N_13163,N_13092);
nand U13313 (N_13313,N_13110,N_13094);
and U13314 (N_13314,N_13140,N_13087);
nand U13315 (N_13315,N_13110,N_13018);
and U13316 (N_13316,N_13162,N_13049);
and U13317 (N_13317,N_13025,N_13045);
xor U13318 (N_13318,N_13011,N_13038);
nor U13319 (N_13319,N_13198,N_13144);
or U13320 (N_13320,N_13161,N_13125);
or U13321 (N_13321,N_13168,N_13193);
and U13322 (N_13322,N_13059,N_13026);
xnor U13323 (N_13323,N_13095,N_13086);
nor U13324 (N_13324,N_13039,N_13029);
and U13325 (N_13325,N_13122,N_13120);
xor U13326 (N_13326,N_13169,N_13092);
nor U13327 (N_13327,N_13121,N_13181);
nand U13328 (N_13328,N_13127,N_13116);
or U13329 (N_13329,N_13194,N_13084);
and U13330 (N_13330,N_13110,N_13051);
or U13331 (N_13331,N_13052,N_13112);
nor U13332 (N_13332,N_13013,N_13020);
and U13333 (N_13333,N_13039,N_13189);
xnor U13334 (N_13334,N_13007,N_13091);
xor U13335 (N_13335,N_13096,N_13027);
xnor U13336 (N_13336,N_13067,N_13101);
nor U13337 (N_13337,N_13085,N_13111);
nor U13338 (N_13338,N_13025,N_13060);
nand U13339 (N_13339,N_13037,N_13103);
xor U13340 (N_13340,N_13128,N_13057);
or U13341 (N_13341,N_13161,N_13140);
or U13342 (N_13342,N_13073,N_13057);
and U13343 (N_13343,N_13000,N_13002);
xor U13344 (N_13344,N_13167,N_13059);
nand U13345 (N_13345,N_13164,N_13165);
and U13346 (N_13346,N_13160,N_13001);
and U13347 (N_13347,N_13060,N_13026);
and U13348 (N_13348,N_13112,N_13186);
or U13349 (N_13349,N_13193,N_13159);
xnor U13350 (N_13350,N_13052,N_13166);
or U13351 (N_13351,N_13003,N_13094);
and U13352 (N_13352,N_13179,N_13189);
nand U13353 (N_13353,N_13147,N_13044);
or U13354 (N_13354,N_13190,N_13040);
xor U13355 (N_13355,N_13128,N_13079);
nor U13356 (N_13356,N_13063,N_13037);
or U13357 (N_13357,N_13189,N_13135);
nor U13358 (N_13358,N_13011,N_13107);
nand U13359 (N_13359,N_13145,N_13102);
nor U13360 (N_13360,N_13157,N_13011);
xor U13361 (N_13361,N_13117,N_13058);
xnor U13362 (N_13362,N_13141,N_13170);
or U13363 (N_13363,N_13080,N_13060);
xor U13364 (N_13364,N_13096,N_13098);
xor U13365 (N_13365,N_13099,N_13169);
xor U13366 (N_13366,N_13118,N_13189);
and U13367 (N_13367,N_13095,N_13117);
nor U13368 (N_13368,N_13013,N_13102);
and U13369 (N_13369,N_13104,N_13019);
and U13370 (N_13370,N_13116,N_13122);
and U13371 (N_13371,N_13071,N_13023);
and U13372 (N_13372,N_13090,N_13065);
or U13373 (N_13373,N_13019,N_13005);
xor U13374 (N_13374,N_13059,N_13070);
or U13375 (N_13375,N_13025,N_13192);
or U13376 (N_13376,N_13139,N_13032);
and U13377 (N_13377,N_13172,N_13004);
nor U13378 (N_13378,N_13165,N_13117);
xor U13379 (N_13379,N_13071,N_13041);
xor U13380 (N_13380,N_13190,N_13055);
nand U13381 (N_13381,N_13151,N_13101);
or U13382 (N_13382,N_13110,N_13005);
and U13383 (N_13383,N_13064,N_13131);
nor U13384 (N_13384,N_13084,N_13020);
and U13385 (N_13385,N_13059,N_13189);
or U13386 (N_13386,N_13091,N_13131);
or U13387 (N_13387,N_13128,N_13078);
or U13388 (N_13388,N_13142,N_13127);
nor U13389 (N_13389,N_13120,N_13024);
or U13390 (N_13390,N_13174,N_13156);
and U13391 (N_13391,N_13190,N_13184);
or U13392 (N_13392,N_13123,N_13187);
xor U13393 (N_13393,N_13127,N_13186);
nand U13394 (N_13394,N_13034,N_13150);
and U13395 (N_13395,N_13152,N_13031);
and U13396 (N_13396,N_13177,N_13071);
xnor U13397 (N_13397,N_13011,N_13110);
nand U13398 (N_13398,N_13111,N_13078);
nor U13399 (N_13399,N_13106,N_13134);
and U13400 (N_13400,N_13319,N_13378);
xnor U13401 (N_13401,N_13222,N_13354);
xnor U13402 (N_13402,N_13274,N_13334);
and U13403 (N_13403,N_13280,N_13208);
nand U13404 (N_13404,N_13376,N_13295);
or U13405 (N_13405,N_13273,N_13324);
nand U13406 (N_13406,N_13327,N_13322);
nand U13407 (N_13407,N_13344,N_13369);
xnor U13408 (N_13408,N_13336,N_13359);
and U13409 (N_13409,N_13333,N_13220);
nand U13410 (N_13410,N_13391,N_13394);
nand U13411 (N_13411,N_13240,N_13297);
nand U13412 (N_13412,N_13370,N_13247);
nand U13413 (N_13413,N_13216,N_13340);
or U13414 (N_13414,N_13356,N_13395);
xnor U13415 (N_13415,N_13380,N_13321);
and U13416 (N_13416,N_13218,N_13215);
nor U13417 (N_13417,N_13304,N_13225);
and U13418 (N_13418,N_13294,N_13347);
and U13419 (N_13419,N_13363,N_13313);
nor U13420 (N_13420,N_13349,N_13352);
xnor U13421 (N_13421,N_13228,N_13379);
nand U13422 (N_13422,N_13383,N_13207);
nand U13423 (N_13423,N_13371,N_13350);
nand U13424 (N_13424,N_13296,N_13287);
nand U13425 (N_13425,N_13377,N_13246);
nand U13426 (N_13426,N_13390,N_13248);
nor U13427 (N_13427,N_13263,N_13374);
xnor U13428 (N_13428,N_13397,N_13241);
or U13429 (N_13429,N_13353,N_13223);
xor U13430 (N_13430,N_13357,N_13330);
nor U13431 (N_13431,N_13221,N_13205);
nor U13432 (N_13432,N_13341,N_13236);
nor U13433 (N_13433,N_13314,N_13217);
or U13434 (N_13434,N_13277,N_13250);
nand U13435 (N_13435,N_13312,N_13213);
or U13436 (N_13436,N_13283,N_13366);
xnor U13437 (N_13437,N_13358,N_13345);
and U13438 (N_13438,N_13282,N_13257);
xnor U13439 (N_13439,N_13329,N_13372);
or U13440 (N_13440,N_13230,N_13275);
nand U13441 (N_13441,N_13293,N_13320);
nor U13442 (N_13442,N_13261,N_13242);
nor U13443 (N_13443,N_13231,N_13335);
nor U13444 (N_13444,N_13239,N_13318);
xnor U13445 (N_13445,N_13233,N_13393);
or U13446 (N_13446,N_13251,N_13386);
and U13447 (N_13447,N_13337,N_13206);
nand U13448 (N_13448,N_13285,N_13382);
or U13449 (N_13449,N_13388,N_13266);
xor U13450 (N_13450,N_13291,N_13278);
and U13451 (N_13451,N_13323,N_13302);
nor U13452 (N_13452,N_13385,N_13332);
or U13453 (N_13453,N_13203,N_13226);
and U13454 (N_13454,N_13219,N_13362);
nand U13455 (N_13455,N_13384,N_13237);
xnor U13456 (N_13456,N_13316,N_13256);
nand U13457 (N_13457,N_13212,N_13286);
nor U13458 (N_13458,N_13298,N_13300);
or U13459 (N_13459,N_13326,N_13209);
nand U13460 (N_13460,N_13214,N_13346);
and U13461 (N_13461,N_13365,N_13305);
nor U13462 (N_13462,N_13254,N_13325);
xor U13463 (N_13463,N_13202,N_13367);
xnor U13464 (N_13464,N_13392,N_13338);
nand U13465 (N_13465,N_13301,N_13328);
nand U13466 (N_13466,N_13309,N_13201);
and U13467 (N_13467,N_13299,N_13258);
or U13468 (N_13468,N_13317,N_13292);
and U13469 (N_13469,N_13368,N_13269);
nor U13470 (N_13470,N_13315,N_13262);
or U13471 (N_13471,N_13264,N_13204);
or U13472 (N_13472,N_13267,N_13310);
nand U13473 (N_13473,N_13270,N_13339);
and U13474 (N_13474,N_13245,N_13381);
nor U13475 (N_13475,N_13252,N_13234);
xnor U13476 (N_13476,N_13279,N_13244);
nor U13477 (N_13477,N_13268,N_13348);
nand U13478 (N_13478,N_13224,N_13272);
nand U13479 (N_13479,N_13306,N_13229);
nor U13480 (N_13480,N_13276,N_13308);
nand U13481 (N_13481,N_13200,N_13271);
and U13482 (N_13482,N_13331,N_13311);
xor U13483 (N_13483,N_13389,N_13211);
or U13484 (N_13484,N_13396,N_13232);
xor U13485 (N_13485,N_13361,N_13243);
nor U13486 (N_13486,N_13235,N_13281);
xor U13487 (N_13487,N_13355,N_13343);
nor U13488 (N_13488,N_13289,N_13307);
and U13489 (N_13489,N_13360,N_13288);
and U13490 (N_13490,N_13373,N_13259);
nand U13491 (N_13491,N_13227,N_13260);
nor U13492 (N_13492,N_13342,N_13238);
xor U13493 (N_13493,N_13265,N_13210);
xnor U13494 (N_13494,N_13351,N_13255);
nand U13495 (N_13495,N_13399,N_13364);
nor U13496 (N_13496,N_13253,N_13375);
and U13497 (N_13497,N_13398,N_13249);
and U13498 (N_13498,N_13284,N_13303);
nor U13499 (N_13499,N_13387,N_13290);
or U13500 (N_13500,N_13283,N_13319);
nor U13501 (N_13501,N_13248,N_13368);
nand U13502 (N_13502,N_13273,N_13251);
nand U13503 (N_13503,N_13288,N_13253);
nor U13504 (N_13504,N_13326,N_13200);
nor U13505 (N_13505,N_13242,N_13394);
and U13506 (N_13506,N_13276,N_13314);
nor U13507 (N_13507,N_13232,N_13315);
nor U13508 (N_13508,N_13258,N_13358);
xor U13509 (N_13509,N_13370,N_13316);
or U13510 (N_13510,N_13325,N_13313);
xnor U13511 (N_13511,N_13284,N_13371);
nor U13512 (N_13512,N_13239,N_13214);
nand U13513 (N_13513,N_13226,N_13364);
and U13514 (N_13514,N_13373,N_13216);
or U13515 (N_13515,N_13355,N_13224);
xor U13516 (N_13516,N_13354,N_13389);
and U13517 (N_13517,N_13391,N_13217);
nor U13518 (N_13518,N_13296,N_13379);
nor U13519 (N_13519,N_13313,N_13271);
nor U13520 (N_13520,N_13234,N_13321);
or U13521 (N_13521,N_13354,N_13233);
xor U13522 (N_13522,N_13264,N_13394);
or U13523 (N_13523,N_13384,N_13271);
and U13524 (N_13524,N_13331,N_13283);
nand U13525 (N_13525,N_13288,N_13283);
xnor U13526 (N_13526,N_13326,N_13248);
and U13527 (N_13527,N_13268,N_13385);
nand U13528 (N_13528,N_13215,N_13333);
and U13529 (N_13529,N_13376,N_13214);
xnor U13530 (N_13530,N_13360,N_13317);
nand U13531 (N_13531,N_13233,N_13222);
or U13532 (N_13532,N_13256,N_13318);
nand U13533 (N_13533,N_13202,N_13269);
and U13534 (N_13534,N_13380,N_13207);
nand U13535 (N_13535,N_13325,N_13302);
and U13536 (N_13536,N_13360,N_13361);
or U13537 (N_13537,N_13370,N_13310);
and U13538 (N_13538,N_13360,N_13228);
and U13539 (N_13539,N_13356,N_13342);
nor U13540 (N_13540,N_13387,N_13204);
nand U13541 (N_13541,N_13318,N_13262);
nor U13542 (N_13542,N_13229,N_13300);
or U13543 (N_13543,N_13247,N_13260);
or U13544 (N_13544,N_13381,N_13282);
or U13545 (N_13545,N_13366,N_13278);
xor U13546 (N_13546,N_13374,N_13339);
and U13547 (N_13547,N_13274,N_13248);
xor U13548 (N_13548,N_13342,N_13217);
or U13549 (N_13549,N_13244,N_13206);
nand U13550 (N_13550,N_13312,N_13225);
and U13551 (N_13551,N_13298,N_13345);
and U13552 (N_13552,N_13332,N_13245);
nand U13553 (N_13553,N_13332,N_13269);
nand U13554 (N_13554,N_13348,N_13221);
xor U13555 (N_13555,N_13295,N_13310);
and U13556 (N_13556,N_13224,N_13203);
or U13557 (N_13557,N_13212,N_13320);
nand U13558 (N_13558,N_13202,N_13240);
or U13559 (N_13559,N_13374,N_13216);
nand U13560 (N_13560,N_13368,N_13291);
or U13561 (N_13561,N_13304,N_13336);
and U13562 (N_13562,N_13372,N_13351);
xor U13563 (N_13563,N_13250,N_13278);
nor U13564 (N_13564,N_13317,N_13274);
and U13565 (N_13565,N_13214,N_13258);
and U13566 (N_13566,N_13346,N_13206);
xor U13567 (N_13567,N_13330,N_13342);
nor U13568 (N_13568,N_13240,N_13392);
xor U13569 (N_13569,N_13223,N_13219);
nor U13570 (N_13570,N_13228,N_13212);
and U13571 (N_13571,N_13225,N_13340);
and U13572 (N_13572,N_13290,N_13259);
xor U13573 (N_13573,N_13270,N_13337);
or U13574 (N_13574,N_13364,N_13230);
nand U13575 (N_13575,N_13243,N_13296);
and U13576 (N_13576,N_13205,N_13330);
and U13577 (N_13577,N_13394,N_13393);
and U13578 (N_13578,N_13312,N_13361);
and U13579 (N_13579,N_13215,N_13212);
or U13580 (N_13580,N_13233,N_13359);
xnor U13581 (N_13581,N_13201,N_13386);
nor U13582 (N_13582,N_13373,N_13351);
xor U13583 (N_13583,N_13322,N_13395);
and U13584 (N_13584,N_13366,N_13393);
and U13585 (N_13585,N_13331,N_13392);
or U13586 (N_13586,N_13328,N_13205);
or U13587 (N_13587,N_13324,N_13304);
or U13588 (N_13588,N_13256,N_13357);
and U13589 (N_13589,N_13288,N_13313);
nand U13590 (N_13590,N_13327,N_13381);
nand U13591 (N_13591,N_13398,N_13284);
xor U13592 (N_13592,N_13350,N_13226);
and U13593 (N_13593,N_13377,N_13316);
and U13594 (N_13594,N_13275,N_13358);
and U13595 (N_13595,N_13335,N_13200);
nand U13596 (N_13596,N_13329,N_13229);
nand U13597 (N_13597,N_13230,N_13283);
or U13598 (N_13598,N_13208,N_13387);
nand U13599 (N_13599,N_13280,N_13229);
or U13600 (N_13600,N_13464,N_13557);
or U13601 (N_13601,N_13441,N_13517);
and U13602 (N_13602,N_13522,N_13487);
nand U13603 (N_13603,N_13577,N_13429);
xor U13604 (N_13604,N_13593,N_13574);
nand U13605 (N_13605,N_13542,N_13415);
xnor U13606 (N_13606,N_13446,N_13523);
nand U13607 (N_13607,N_13581,N_13416);
and U13608 (N_13608,N_13536,N_13481);
xor U13609 (N_13609,N_13453,N_13566);
and U13610 (N_13610,N_13412,N_13496);
xor U13611 (N_13611,N_13587,N_13569);
or U13612 (N_13612,N_13562,N_13485);
or U13613 (N_13613,N_13514,N_13451);
nor U13614 (N_13614,N_13466,N_13431);
or U13615 (N_13615,N_13424,N_13433);
nor U13616 (N_13616,N_13545,N_13571);
and U13617 (N_13617,N_13544,N_13539);
or U13618 (N_13618,N_13478,N_13530);
and U13619 (N_13619,N_13471,N_13546);
nand U13620 (N_13620,N_13499,N_13426);
nand U13621 (N_13621,N_13472,N_13452);
nor U13622 (N_13622,N_13435,N_13457);
and U13623 (N_13623,N_13537,N_13510);
and U13624 (N_13624,N_13505,N_13428);
nor U13625 (N_13625,N_13506,N_13486);
and U13626 (N_13626,N_13404,N_13576);
nand U13627 (N_13627,N_13443,N_13520);
or U13628 (N_13628,N_13526,N_13449);
nand U13629 (N_13629,N_13531,N_13425);
xor U13630 (N_13630,N_13475,N_13589);
nor U13631 (N_13631,N_13403,N_13518);
and U13632 (N_13632,N_13543,N_13463);
or U13633 (N_13633,N_13555,N_13417);
or U13634 (N_13634,N_13549,N_13553);
nand U13635 (N_13635,N_13405,N_13447);
and U13636 (N_13636,N_13459,N_13411);
nor U13637 (N_13637,N_13439,N_13473);
nor U13638 (N_13638,N_13568,N_13401);
and U13639 (N_13639,N_13570,N_13525);
and U13640 (N_13640,N_13504,N_13594);
and U13641 (N_13641,N_13414,N_13437);
nor U13642 (N_13642,N_13560,N_13507);
nor U13643 (N_13643,N_13552,N_13434);
nor U13644 (N_13644,N_13400,N_13407);
xnor U13645 (N_13645,N_13578,N_13529);
or U13646 (N_13646,N_13567,N_13575);
nand U13647 (N_13647,N_13524,N_13460);
xnor U13648 (N_13648,N_13468,N_13572);
nand U13649 (N_13649,N_13590,N_13527);
nor U13650 (N_13650,N_13503,N_13558);
and U13651 (N_13651,N_13516,N_13551);
nand U13652 (N_13652,N_13461,N_13595);
nor U13653 (N_13653,N_13588,N_13479);
nor U13654 (N_13654,N_13535,N_13584);
nand U13655 (N_13655,N_13440,N_13597);
nor U13656 (N_13656,N_13580,N_13501);
nand U13657 (N_13657,N_13563,N_13483);
and U13658 (N_13658,N_13533,N_13469);
or U13659 (N_13659,N_13476,N_13474);
xnor U13660 (N_13660,N_13482,N_13515);
nand U13661 (N_13661,N_13421,N_13458);
or U13662 (N_13662,N_13427,N_13491);
and U13663 (N_13663,N_13502,N_13493);
nor U13664 (N_13664,N_13534,N_13423);
nor U13665 (N_13665,N_13492,N_13442);
nor U13666 (N_13666,N_13490,N_13556);
nor U13667 (N_13667,N_13489,N_13559);
xor U13668 (N_13668,N_13432,N_13436);
xor U13669 (N_13669,N_13418,N_13430);
nand U13670 (N_13670,N_13444,N_13513);
nand U13671 (N_13671,N_13438,N_13410);
or U13672 (N_13672,N_13413,N_13409);
nand U13673 (N_13673,N_13500,N_13406);
or U13674 (N_13674,N_13511,N_13512);
or U13675 (N_13675,N_13494,N_13547);
and U13676 (N_13676,N_13455,N_13448);
and U13677 (N_13677,N_13598,N_13599);
or U13678 (N_13678,N_13521,N_13585);
xor U13679 (N_13679,N_13538,N_13561);
nand U13680 (N_13680,N_13419,N_13591);
or U13681 (N_13681,N_13497,N_13554);
or U13682 (N_13682,N_13454,N_13519);
nor U13683 (N_13683,N_13422,N_13509);
or U13684 (N_13684,N_13484,N_13420);
xnor U13685 (N_13685,N_13541,N_13564);
or U13686 (N_13686,N_13586,N_13582);
or U13687 (N_13687,N_13532,N_13508);
nor U13688 (N_13688,N_13550,N_13596);
or U13689 (N_13689,N_13470,N_13528);
nand U13690 (N_13690,N_13462,N_13445);
nor U13691 (N_13691,N_13402,N_13548);
nor U13692 (N_13692,N_13540,N_13467);
nand U13693 (N_13693,N_13579,N_13565);
xor U13694 (N_13694,N_13592,N_13465);
nand U13695 (N_13695,N_13456,N_13477);
nand U13696 (N_13696,N_13450,N_13408);
nor U13697 (N_13697,N_13583,N_13573);
and U13698 (N_13698,N_13498,N_13495);
and U13699 (N_13699,N_13480,N_13488);
nand U13700 (N_13700,N_13565,N_13514);
and U13701 (N_13701,N_13503,N_13591);
and U13702 (N_13702,N_13442,N_13553);
xor U13703 (N_13703,N_13559,N_13496);
or U13704 (N_13704,N_13553,N_13515);
or U13705 (N_13705,N_13553,N_13537);
or U13706 (N_13706,N_13482,N_13525);
and U13707 (N_13707,N_13413,N_13578);
nand U13708 (N_13708,N_13543,N_13589);
or U13709 (N_13709,N_13563,N_13471);
nand U13710 (N_13710,N_13539,N_13533);
or U13711 (N_13711,N_13416,N_13439);
and U13712 (N_13712,N_13534,N_13571);
or U13713 (N_13713,N_13571,N_13566);
and U13714 (N_13714,N_13425,N_13595);
and U13715 (N_13715,N_13455,N_13427);
and U13716 (N_13716,N_13514,N_13558);
and U13717 (N_13717,N_13431,N_13561);
or U13718 (N_13718,N_13496,N_13480);
nor U13719 (N_13719,N_13400,N_13459);
nor U13720 (N_13720,N_13593,N_13407);
or U13721 (N_13721,N_13468,N_13579);
and U13722 (N_13722,N_13516,N_13575);
and U13723 (N_13723,N_13492,N_13581);
and U13724 (N_13724,N_13559,N_13526);
and U13725 (N_13725,N_13462,N_13584);
xor U13726 (N_13726,N_13527,N_13430);
xnor U13727 (N_13727,N_13513,N_13462);
or U13728 (N_13728,N_13429,N_13416);
or U13729 (N_13729,N_13449,N_13487);
nor U13730 (N_13730,N_13440,N_13452);
or U13731 (N_13731,N_13550,N_13441);
and U13732 (N_13732,N_13432,N_13510);
or U13733 (N_13733,N_13459,N_13480);
or U13734 (N_13734,N_13558,N_13536);
or U13735 (N_13735,N_13565,N_13590);
and U13736 (N_13736,N_13480,N_13579);
xnor U13737 (N_13737,N_13482,N_13585);
or U13738 (N_13738,N_13498,N_13434);
nor U13739 (N_13739,N_13575,N_13416);
nand U13740 (N_13740,N_13413,N_13437);
nor U13741 (N_13741,N_13555,N_13432);
nor U13742 (N_13742,N_13485,N_13412);
nor U13743 (N_13743,N_13478,N_13538);
nor U13744 (N_13744,N_13533,N_13566);
nor U13745 (N_13745,N_13475,N_13543);
xnor U13746 (N_13746,N_13446,N_13447);
nor U13747 (N_13747,N_13565,N_13523);
nor U13748 (N_13748,N_13518,N_13580);
nor U13749 (N_13749,N_13587,N_13555);
xor U13750 (N_13750,N_13462,N_13438);
xnor U13751 (N_13751,N_13422,N_13572);
nor U13752 (N_13752,N_13582,N_13526);
or U13753 (N_13753,N_13541,N_13474);
or U13754 (N_13754,N_13464,N_13478);
xor U13755 (N_13755,N_13424,N_13453);
nor U13756 (N_13756,N_13478,N_13585);
nor U13757 (N_13757,N_13532,N_13585);
and U13758 (N_13758,N_13494,N_13576);
xor U13759 (N_13759,N_13473,N_13488);
or U13760 (N_13760,N_13583,N_13442);
and U13761 (N_13761,N_13582,N_13574);
nand U13762 (N_13762,N_13500,N_13583);
nor U13763 (N_13763,N_13421,N_13598);
or U13764 (N_13764,N_13541,N_13486);
and U13765 (N_13765,N_13596,N_13499);
nor U13766 (N_13766,N_13529,N_13509);
nor U13767 (N_13767,N_13485,N_13538);
or U13768 (N_13768,N_13563,N_13514);
nand U13769 (N_13769,N_13443,N_13433);
and U13770 (N_13770,N_13502,N_13562);
or U13771 (N_13771,N_13432,N_13485);
nor U13772 (N_13772,N_13570,N_13514);
or U13773 (N_13773,N_13519,N_13598);
nor U13774 (N_13774,N_13496,N_13418);
and U13775 (N_13775,N_13466,N_13561);
or U13776 (N_13776,N_13427,N_13544);
nor U13777 (N_13777,N_13460,N_13479);
nand U13778 (N_13778,N_13578,N_13451);
nor U13779 (N_13779,N_13595,N_13558);
or U13780 (N_13780,N_13429,N_13404);
or U13781 (N_13781,N_13478,N_13421);
or U13782 (N_13782,N_13446,N_13512);
and U13783 (N_13783,N_13412,N_13492);
nor U13784 (N_13784,N_13502,N_13489);
or U13785 (N_13785,N_13478,N_13486);
nand U13786 (N_13786,N_13477,N_13544);
and U13787 (N_13787,N_13599,N_13542);
and U13788 (N_13788,N_13560,N_13482);
and U13789 (N_13789,N_13415,N_13431);
nand U13790 (N_13790,N_13480,N_13484);
or U13791 (N_13791,N_13479,N_13403);
or U13792 (N_13792,N_13415,N_13416);
nor U13793 (N_13793,N_13594,N_13518);
xnor U13794 (N_13794,N_13584,N_13511);
nor U13795 (N_13795,N_13502,N_13582);
and U13796 (N_13796,N_13416,N_13485);
nand U13797 (N_13797,N_13513,N_13405);
nor U13798 (N_13798,N_13463,N_13580);
xor U13799 (N_13799,N_13416,N_13515);
and U13800 (N_13800,N_13673,N_13631);
and U13801 (N_13801,N_13761,N_13708);
nor U13802 (N_13802,N_13689,N_13753);
and U13803 (N_13803,N_13735,N_13739);
nor U13804 (N_13804,N_13626,N_13718);
or U13805 (N_13805,N_13773,N_13712);
or U13806 (N_13806,N_13664,N_13792);
nand U13807 (N_13807,N_13774,N_13662);
or U13808 (N_13808,N_13757,N_13674);
nor U13809 (N_13809,N_13747,N_13691);
and U13810 (N_13810,N_13690,N_13607);
and U13811 (N_13811,N_13786,N_13637);
and U13812 (N_13812,N_13639,N_13726);
or U13813 (N_13813,N_13759,N_13738);
nand U13814 (N_13814,N_13781,N_13653);
nand U13815 (N_13815,N_13789,N_13630);
and U13816 (N_13816,N_13658,N_13633);
and U13817 (N_13817,N_13788,N_13696);
nand U13818 (N_13818,N_13778,N_13672);
xnor U13819 (N_13819,N_13681,N_13769);
or U13820 (N_13820,N_13706,N_13733);
xor U13821 (N_13821,N_13725,N_13799);
and U13822 (N_13822,N_13621,N_13755);
and U13823 (N_13823,N_13635,N_13750);
nor U13824 (N_13824,N_13765,N_13790);
nand U13825 (N_13825,N_13685,N_13612);
nor U13826 (N_13826,N_13628,N_13796);
nand U13827 (N_13827,N_13716,N_13693);
xnor U13828 (N_13828,N_13697,N_13665);
nand U13829 (N_13829,N_13652,N_13627);
xnor U13830 (N_13830,N_13709,N_13734);
nand U13831 (N_13831,N_13701,N_13651);
and U13832 (N_13832,N_13636,N_13794);
and U13833 (N_13833,N_13613,N_13704);
nor U13834 (N_13834,N_13719,N_13772);
and U13835 (N_13835,N_13643,N_13713);
or U13836 (N_13836,N_13618,N_13604);
or U13837 (N_13837,N_13638,N_13793);
nor U13838 (N_13838,N_13608,N_13655);
xnor U13839 (N_13839,N_13752,N_13629);
and U13840 (N_13840,N_13707,N_13710);
xor U13841 (N_13841,N_13601,N_13732);
and U13842 (N_13842,N_13632,N_13714);
or U13843 (N_13843,N_13666,N_13650);
or U13844 (N_13844,N_13740,N_13670);
and U13845 (N_13845,N_13727,N_13785);
nor U13846 (N_13846,N_13657,N_13768);
or U13847 (N_13847,N_13600,N_13787);
or U13848 (N_13848,N_13663,N_13620);
and U13849 (N_13849,N_13784,N_13602);
nor U13850 (N_13850,N_13671,N_13659);
nor U13851 (N_13851,N_13642,N_13669);
nand U13852 (N_13852,N_13783,N_13688);
xor U13853 (N_13853,N_13743,N_13634);
nor U13854 (N_13854,N_13703,N_13700);
nor U13855 (N_13855,N_13728,N_13647);
xor U13856 (N_13856,N_13623,N_13646);
nor U13857 (N_13857,N_13782,N_13771);
or U13858 (N_13858,N_13722,N_13721);
nand U13859 (N_13859,N_13680,N_13683);
xnor U13860 (N_13860,N_13731,N_13737);
nand U13861 (N_13861,N_13758,N_13711);
nor U13862 (N_13862,N_13742,N_13684);
nor U13863 (N_13863,N_13695,N_13617);
xnor U13864 (N_13864,N_13641,N_13741);
and U13865 (N_13865,N_13720,N_13748);
nand U13866 (N_13866,N_13640,N_13756);
nand U13867 (N_13867,N_13744,N_13677);
xor U13868 (N_13868,N_13678,N_13609);
xnor U13869 (N_13869,N_13699,N_13798);
nor U13870 (N_13870,N_13687,N_13698);
and U13871 (N_13871,N_13705,N_13780);
or U13872 (N_13872,N_13729,N_13745);
nand U13873 (N_13873,N_13749,N_13625);
or U13874 (N_13874,N_13797,N_13676);
xnor U13875 (N_13875,N_13692,N_13622);
and U13876 (N_13876,N_13645,N_13616);
xor U13877 (N_13877,N_13715,N_13770);
nand U13878 (N_13878,N_13606,N_13679);
and U13879 (N_13879,N_13614,N_13754);
or U13880 (N_13880,N_13654,N_13694);
and U13881 (N_13881,N_13675,N_13615);
nand U13882 (N_13882,N_13779,N_13777);
and U13883 (N_13883,N_13776,N_13751);
xnor U13884 (N_13884,N_13775,N_13648);
or U13885 (N_13885,N_13760,N_13649);
and U13886 (N_13886,N_13746,N_13605);
nor U13887 (N_13887,N_13660,N_13702);
nor U13888 (N_13888,N_13661,N_13791);
or U13889 (N_13889,N_13724,N_13624);
or U13890 (N_13890,N_13656,N_13795);
nand U13891 (N_13891,N_13611,N_13667);
or U13892 (N_13892,N_13764,N_13644);
and U13893 (N_13893,N_13723,N_13766);
or U13894 (N_13894,N_13717,N_13668);
xnor U13895 (N_13895,N_13730,N_13686);
and U13896 (N_13896,N_13763,N_13762);
or U13897 (N_13897,N_13767,N_13682);
or U13898 (N_13898,N_13610,N_13736);
nand U13899 (N_13899,N_13603,N_13619);
nand U13900 (N_13900,N_13627,N_13772);
and U13901 (N_13901,N_13695,N_13716);
nor U13902 (N_13902,N_13745,N_13686);
nand U13903 (N_13903,N_13762,N_13759);
or U13904 (N_13904,N_13618,N_13796);
and U13905 (N_13905,N_13626,N_13600);
and U13906 (N_13906,N_13610,N_13686);
xnor U13907 (N_13907,N_13743,N_13639);
and U13908 (N_13908,N_13728,N_13627);
or U13909 (N_13909,N_13781,N_13790);
nand U13910 (N_13910,N_13734,N_13635);
xnor U13911 (N_13911,N_13715,N_13755);
or U13912 (N_13912,N_13634,N_13650);
or U13913 (N_13913,N_13766,N_13751);
and U13914 (N_13914,N_13687,N_13643);
nor U13915 (N_13915,N_13627,N_13614);
or U13916 (N_13916,N_13705,N_13748);
and U13917 (N_13917,N_13624,N_13674);
or U13918 (N_13918,N_13651,N_13664);
nor U13919 (N_13919,N_13752,N_13769);
and U13920 (N_13920,N_13789,N_13681);
nand U13921 (N_13921,N_13724,N_13788);
or U13922 (N_13922,N_13636,N_13642);
and U13923 (N_13923,N_13643,N_13650);
or U13924 (N_13924,N_13625,N_13636);
and U13925 (N_13925,N_13703,N_13775);
or U13926 (N_13926,N_13704,N_13621);
and U13927 (N_13927,N_13780,N_13702);
and U13928 (N_13928,N_13750,N_13796);
and U13929 (N_13929,N_13747,N_13782);
nand U13930 (N_13930,N_13725,N_13787);
or U13931 (N_13931,N_13706,N_13707);
nor U13932 (N_13932,N_13679,N_13653);
nand U13933 (N_13933,N_13793,N_13681);
xor U13934 (N_13934,N_13729,N_13667);
nor U13935 (N_13935,N_13702,N_13740);
xor U13936 (N_13936,N_13631,N_13619);
nand U13937 (N_13937,N_13653,N_13638);
and U13938 (N_13938,N_13788,N_13630);
nor U13939 (N_13939,N_13766,N_13621);
nand U13940 (N_13940,N_13625,N_13779);
or U13941 (N_13941,N_13715,N_13663);
or U13942 (N_13942,N_13662,N_13683);
nand U13943 (N_13943,N_13668,N_13736);
nand U13944 (N_13944,N_13680,N_13777);
or U13945 (N_13945,N_13719,N_13618);
or U13946 (N_13946,N_13621,N_13694);
nor U13947 (N_13947,N_13770,N_13705);
nor U13948 (N_13948,N_13709,N_13728);
nand U13949 (N_13949,N_13657,N_13771);
and U13950 (N_13950,N_13787,N_13679);
xor U13951 (N_13951,N_13788,N_13623);
nand U13952 (N_13952,N_13775,N_13791);
nor U13953 (N_13953,N_13667,N_13759);
or U13954 (N_13954,N_13744,N_13650);
xor U13955 (N_13955,N_13739,N_13650);
and U13956 (N_13956,N_13795,N_13668);
or U13957 (N_13957,N_13719,N_13653);
nor U13958 (N_13958,N_13761,N_13741);
xor U13959 (N_13959,N_13649,N_13609);
and U13960 (N_13960,N_13629,N_13700);
or U13961 (N_13961,N_13798,N_13737);
nand U13962 (N_13962,N_13783,N_13656);
nor U13963 (N_13963,N_13614,N_13700);
xor U13964 (N_13964,N_13742,N_13703);
and U13965 (N_13965,N_13725,N_13749);
and U13966 (N_13966,N_13744,N_13757);
xor U13967 (N_13967,N_13700,N_13757);
nand U13968 (N_13968,N_13640,N_13671);
nor U13969 (N_13969,N_13603,N_13768);
or U13970 (N_13970,N_13609,N_13625);
xnor U13971 (N_13971,N_13741,N_13721);
and U13972 (N_13972,N_13768,N_13690);
or U13973 (N_13973,N_13636,N_13600);
xor U13974 (N_13974,N_13793,N_13706);
xor U13975 (N_13975,N_13628,N_13777);
and U13976 (N_13976,N_13789,N_13687);
and U13977 (N_13977,N_13601,N_13665);
nor U13978 (N_13978,N_13664,N_13711);
or U13979 (N_13979,N_13635,N_13610);
nand U13980 (N_13980,N_13751,N_13615);
xor U13981 (N_13981,N_13732,N_13711);
nor U13982 (N_13982,N_13793,N_13771);
nor U13983 (N_13983,N_13671,N_13765);
nand U13984 (N_13984,N_13628,N_13734);
and U13985 (N_13985,N_13610,N_13660);
and U13986 (N_13986,N_13693,N_13671);
nand U13987 (N_13987,N_13712,N_13741);
and U13988 (N_13988,N_13748,N_13678);
or U13989 (N_13989,N_13748,N_13745);
xnor U13990 (N_13990,N_13784,N_13678);
or U13991 (N_13991,N_13690,N_13645);
or U13992 (N_13992,N_13603,N_13633);
xor U13993 (N_13993,N_13653,N_13600);
and U13994 (N_13994,N_13645,N_13642);
or U13995 (N_13995,N_13719,N_13775);
nor U13996 (N_13996,N_13630,N_13651);
or U13997 (N_13997,N_13633,N_13757);
nor U13998 (N_13998,N_13660,N_13691);
xnor U13999 (N_13999,N_13724,N_13799);
or U14000 (N_14000,N_13953,N_13935);
nor U14001 (N_14001,N_13892,N_13917);
nor U14002 (N_14002,N_13849,N_13927);
nor U14003 (N_14003,N_13924,N_13966);
nor U14004 (N_14004,N_13813,N_13895);
nand U14005 (N_14005,N_13918,N_13990);
nand U14006 (N_14006,N_13902,N_13983);
and U14007 (N_14007,N_13908,N_13971);
and U14008 (N_14008,N_13838,N_13843);
nand U14009 (N_14009,N_13882,N_13993);
xnor U14010 (N_14010,N_13955,N_13840);
and U14011 (N_14011,N_13827,N_13820);
and U14012 (N_14012,N_13941,N_13867);
nand U14013 (N_14013,N_13981,N_13873);
or U14014 (N_14014,N_13959,N_13828);
and U14015 (N_14015,N_13804,N_13862);
or U14016 (N_14016,N_13894,N_13845);
xor U14017 (N_14017,N_13992,N_13961);
nor U14018 (N_14018,N_13920,N_13815);
xor U14019 (N_14019,N_13984,N_13914);
nand U14020 (N_14020,N_13853,N_13881);
and U14021 (N_14021,N_13883,N_13965);
nor U14022 (N_14022,N_13964,N_13814);
and U14023 (N_14023,N_13829,N_13926);
and U14024 (N_14024,N_13865,N_13887);
or U14025 (N_14025,N_13866,N_13831);
xnor U14026 (N_14026,N_13806,N_13989);
and U14027 (N_14027,N_13844,N_13839);
or U14028 (N_14028,N_13886,N_13995);
nor U14029 (N_14029,N_13904,N_13847);
nand U14030 (N_14030,N_13958,N_13808);
or U14031 (N_14031,N_13909,N_13852);
or U14032 (N_14032,N_13987,N_13925);
nand U14033 (N_14033,N_13817,N_13977);
xor U14034 (N_14034,N_13837,N_13871);
or U14035 (N_14035,N_13952,N_13994);
and U14036 (N_14036,N_13946,N_13930);
or U14037 (N_14037,N_13803,N_13949);
nor U14038 (N_14038,N_13963,N_13851);
nand U14039 (N_14039,N_13972,N_13985);
xnor U14040 (N_14040,N_13931,N_13915);
and U14041 (N_14041,N_13980,N_13822);
or U14042 (N_14042,N_13802,N_13923);
or U14043 (N_14043,N_13807,N_13929);
nand U14044 (N_14044,N_13970,N_13896);
nand U14045 (N_14045,N_13830,N_13968);
and U14046 (N_14046,N_13899,N_13922);
nand U14047 (N_14047,N_13835,N_13874);
and U14048 (N_14048,N_13864,N_13906);
nor U14049 (N_14049,N_13893,N_13880);
and U14050 (N_14050,N_13901,N_13816);
xor U14051 (N_14051,N_13832,N_13969);
nand U14052 (N_14052,N_13956,N_13942);
xor U14053 (N_14053,N_13868,N_13975);
xor U14054 (N_14054,N_13860,N_13944);
xnor U14055 (N_14055,N_13898,N_13863);
nor U14056 (N_14056,N_13848,N_13951);
nor U14057 (N_14057,N_13912,N_13945);
and U14058 (N_14058,N_13858,N_13879);
nor U14059 (N_14059,N_13876,N_13928);
and U14060 (N_14060,N_13823,N_13903);
xnor U14061 (N_14061,N_13910,N_13982);
nand U14062 (N_14062,N_13937,N_13996);
xor U14063 (N_14063,N_13861,N_13991);
and U14064 (N_14064,N_13940,N_13885);
nor U14065 (N_14065,N_13978,N_13809);
nor U14066 (N_14066,N_13960,N_13855);
nand U14067 (N_14067,N_13997,N_13810);
or U14068 (N_14068,N_13821,N_13934);
or U14069 (N_14069,N_13933,N_13811);
and U14070 (N_14070,N_13905,N_13936);
nor U14071 (N_14071,N_13998,N_13939);
and U14072 (N_14072,N_13836,N_13818);
nor U14073 (N_14073,N_13907,N_13801);
nand U14074 (N_14074,N_13800,N_13919);
or U14075 (N_14075,N_13859,N_13850);
xor U14076 (N_14076,N_13913,N_13842);
and U14077 (N_14077,N_13957,N_13884);
and U14078 (N_14078,N_13825,N_13878);
or U14079 (N_14079,N_13948,N_13979);
nand U14080 (N_14080,N_13834,N_13856);
nor U14081 (N_14081,N_13986,N_13889);
xor U14082 (N_14082,N_13897,N_13999);
nor U14083 (N_14083,N_13932,N_13872);
xnor U14084 (N_14084,N_13819,N_13841);
nand U14085 (N_14085,N_13805,N_13921);
nand U14086 (N_14086,N_13812,N_13833);
nand U14087 (N_14087,N_13890,N_13943);
nor U14088 (N_14088,N_13954,N_13857);
or U14089 (N_14089,N_13967,N_13891);
and U14090 (N_14090,N_13950,N_13938);
or U14091 (N_14091,N_13870,N_13869);
and U14092 (N_14092,N_13976,N_13875);
or U14093 (N_14093,N_13826,N_13962);
nand U14094 (N_14094,N_13947,N_13916);
and U14095 (N_14095,N_13854,N_13824);
and U14096 (N_14096,N_13988,N_13888);
or U14097 (N_14097,N_13911,N_13900);
nor U14098 (N_14098,N_13846,N_13877);
and U14099 (N_14099,N_13973,N_13974);
or U14100 (N_14100,N_13847,N_13915);
nor U14101 (N_14101,N_13915,N_13859);
nand U14102 (N_14102,N_13831,N_13963);
xnor U14103 (N_14103,N_13858,N_13920);
or U14104 (N_14104,N_13941,N_13861);
xnor U14105 (N_14105,N_13970,N_13881);
nand U14106 (N_14106,N_13991,N_13877);
or U14107 (N_14107,N_13897,N_13887);
nor U14108 (N_14108,N_13993,N_13856);
and U14109 (N_14109,N_13929,N_13983);
nor U14110 (N_14110,N_13864,N_13949);
and U14111 (N_14111,N_13808,N_13946);
nand U14112 (N_14112,N_13892,N_13886);
nor U14113 (N_14113,N_13936,N_13849);
nor U14114 (N_14114,N_13948,N_13967);
and U14115 (N_14115,N_13869,N_13899);
nand U14116 (N_14116,N_13830,N_13918);
and U14117 (N_14117,N_13913,N_13946);
and U14118 (N_14118,N_13967,N_13864);
nand U14119 (N_14119,N_13805,N_13925);
or U14120 (N_14120,N_13840,N_13931);
nor U14121 (N_14121,N_13838,N_13834);
and U14122 (N_14122,N_13862,N_13994);
xor U14123 (N_14123,N_13983,N_13868);
and U14124 (N_14124,N_13938,N_13906);
and U14125 (N_14125,N_13904,N_13935);
and U14126 (N_14126,N_13855,N_13928);
nor U14127 (N_14127,N_13981,N_13957);
and U14128 (N_14128,N_13881,N_13816);
nand U14129 (N_14129,N_13866,N_13965);
or U14130 (N_14130,N_13870,N_13913);
nand U14131 (N_14131,N_13910,N_13892);
and U14132 (N_14132,N_13851,N_13889);
nor U14133 (N_14133,N_13842,N_13845);
and U14134 (N_14134,N_13833,N_13895);
and U14135 (N_14135,N_13821,N_13980);
nand U14136 (N_14136,N_13876,N_13816);
nand U14137 (N_14137,N_13855,N_13847);
and U14138 (N_14138,N_13968,N_13859);
and U14139 (N_14139,N_13983,N_13947);
or U14140 (N_14140,N_13947,N_13995);
xor U14141 (N_14141,N_13867,N_13975);
nor U14142 (N_14142,N_13929,N_13896);
nand U14143 (N_14143,N_13935,N_13825);
and U14144 (N_14144,N_13885,N_13974);
and U14145 (N_14145,N_13977,N_13925);
and U14146 (N_14146,N_13936,N_13993);
or U14147 (N_14147,N_13908,N_13836);
nor U14148 (N_14148,N_13824,N_13925);
xnor U14149 (N_14149,N_13947,N_13893);
nor U14150 (N_14150,N_13885,N_13918);
or U14151 (N_14151,N_13877,N_13800);
and U14152 (N_14152,N_13804,N_13890);
xor U14153 (N_14153,N_13885,N_13842);
and U14154 (N_14154,N_13988,N_13952);
xnor U14155 (N_14155,N_13936,N_13940);
xor U14156 (N_14156,N_13924,N_13864);
and U14157 (N_14157,N_13853,N_13858);
nand U14158 (N_14158,N_13967,N_13957);
xnor U14159 (N_14159,N_13945,N_13891);
nor U14160 (N_14160,N_13825,N_13872);
and U14161 (N_14161,N_13993,N_13959);
xor U14162 (N_14162,N_13806,N_13819);
and U14163 (N_14163,N_13803,N_13875);
xnor U14164 (N_14164,N_13945,N_13866);
nand U14165 (N_14165,N_13888,N_13980);
nor U14166 (N_14166,N_13911,N_13955);
xor U14167 (N_14167,N_13890,N_13987);
nor U14168 (N_14168,N_13967,N_13998);
or U14169 (N_14169,N_13941,N_13852);
xor U14170 (N_14170,N_13892,N_13965);
nor U14171 (N_14171,N_13880,N_13974);
and U14172 (N_14172,N_13826,N_13998);
xnor U14173 (N_14173,N_13976,N_13983);
xor U14174 (N_14174,N_13992,N_13904);
nor U14175 (N_14175,N_13801,N_13864);
or U14176 (N_14176,N_13869,N_13817);
xnor U14177 (N_14177,N_13862,N_13964);
and U14178 (N_14178,N_13919,N_13987);
or U14179 (N_14179,N_13812,N_13973);
and U14180 (N_14180,N_13905,N_13942);
nand U14181 (N_14181,N_13870,N_13804);
nor U14182 (N_14182,N_13848,N_13985);
nor U14183 (N_14183,N_13973,N_13922);
xor U14184 (N_14184,N_13906,N_13896);
nor U14185 (N_14185,N_13885,N_13912);
xnor U14186 (N_14186,N_13812,N_13903);
nor U14187 (N_14187,N_13943,N_13953);
and U14188 (N_14188,N_13865,N_13827);
or U14189 (N_14189,N_13824,N_13879);
nor U14190 (N_14190,N_13826,N_13987);
nand U14191 (N_14191,N_13934,N_13901);
and U14192 (N_14192,N_13858,N_13921);
nand U14193 (N_14193,N_13973,N_13972);
nor U14194 (N_14194,N_13914,N_13994);
or U14195 (N_14195,N_13859,N_13905);
nor U14196 (N_14196,N_13842,N_13868);
and U14197 (N_14197,N_13835,N_13960);
or U14198 (N_14198,N_13901,N_13930);
xnor U14199 (N_14199,N_13941,N_13831);
xor U14200 (N_14200,N_14197,N_14004);
nor U14201 (N_14201,N_14021,N_14107);
or U14202 (N_14202,N_14164,N_14122);
xnor U14203 (N_14203,N_14047,N_14028);
or U14204 (N_14204,N_14114,N_14163);
and U14205 (N_14205,N_14043,N_14084);
or U14206 (N_14206,N_14187,N_14041);
or U14207 (N_14207,N_14133,N_14030);
nand U14208 (N_14208,N_14037,N_14170);
and U14209 (N_14209,N_14058,N_14108);
and U14210 (N_14210,N_14153,N_14008);
nor U14211 (N_14211,N_14131,N_14144);
nand U14212 (N_14212,N_14101,N_14134);
and U14213 (N_14213,N_14152,N_14066);
xnor U14214 (N_14214,N_14075,N_14129);
and U14215 (N_14215,N_14027,N_14160);
nor U14216 (N_14216,N_14154,N_14177);
nor U14217 (N_14217,N_14173,N_14125);
xnor U14218 (N_14218,N_14033,N_14046);
nor U14219 (N_14219,N_14087,N_14146);
nor U14220 (N_14220,N_14169,N_14198);
nor U14221 (N_14221,N_14090,N_14062);
xnor U14222 (N_14222,N_14113,N_14005);
or U14223 (N_14223,N_14091,N_14199);
nand U14224 (N_14224,N_14011,N_14151);
nor U14225 (N_14225,N_14132,N_14002);
and U14226 (N_14226,N_14168,N_14106);
nor U14227 (N_14227,N_14159,N_14086);
or U14228 (N_14228,N_14092,N_14055);
nand U14229 (N_14229,N_14098,N_14083);
nor U14230 (N_14230,N_14025,N_14023);
xnor U14231 (N_14231,N_14180,N_14149);
and U14232 (N_14232,N_14095,N_14182);
and U14233 (N_14233,N_14038,N_14079);
nor U14234 (N_14234,N_14121,N_14157);
or U14235 (N_14235,N_14116,N_14059);
or U14236 (N_14236,N_14103,N_14105);
nor U14237 (N_14237,N_14167,N_14060);
xor U14238 (N_14238,N_14150,N_14172);
nor U14239 (N_14239,N_14010,N_14053);
or U14240 (N_14240,N_14142,N_14089);
nor U14241 (N_14241,N_14094,N_14052);
xor U14242 (N_14242,N_14138,N_14127);
xor U14243 (N_14243,N_14147,N_14069);
nand U14244 (N_14244,N_14049,N_14067);
and U14245 (N_14245,N_14063,N_14034);
and U14246 (N_14246,N_14189,N_14136);
nand U14247 (N_14247,N_14191,N_14056);
nor U14248 (N_14248,N_14076,N_14186);
xnor U14249 (N_14249,N_14093,N_14143);
and U14250 (N_14250,N_14057,N_14019);
nand U14251 (N_14251,N_14035,N_14013);
or U14252 (N_14252,N_14074,N_14012);
nor U14253 (N_14253,N_14123,N_14139);
or U14254 (N_14254,N_14188,N_14158);
or U14255 (N_14255,N_14007,N_14088);
nor U14256 (N_14256,N_14175,N_14071);
or U14257 (N_14257,N_14064,N_14140);
nand U14258 (N_14258,N_14014,N_14009);
or U14259 (N_14259,N_14096,N_14048);
nand U14260 (N_14260,N_14085,N_14104);
and U14261 (N_14261,N_14174,N_14045);
and U14262 (N_14262,N_14166,N_14016);
and U14263 (N_14263,N_14073,N_14119);
or U14264 (N_14264,N_14161,N_14165);
nor U14265 (N_14265,N_14050,N_14178);
or U14266 (N_14266,N_14130,N_14137);
xor U14267 (N_14267,N_14051,N_14003);
or U14268 (N_14268,N_14078,N_14190);
xor U14269 (N_14269,N_14195,N_14109);
or U14270 (N_14270,N_14039,N_14081);
and U14271 (N_14271,N_14112,N_14036);
nor U14272 (N_14272,N_14061,N_14171);
and U14273 (N_14273,N_14141,N_14006);
nor U14274 (N_14274,N_14044,N_14031);
or U14275 (N_14275,N_14192,N_14026);
nand U14276 (N_14276,N_14184,N_14126);
or U14277 (N_14277,N_14054,N_14042);
xor U14278 (N_14278,N_14001,N_14162);
or U14279 (N_14279,N_14024,N_14100);
xor U14280 (N_14280,N_14135,N_14145);
nor U14281 (N_14281,N_14022,N_14097);
xnor U14282 (N_14282,N_14117,N_14179);
nor U14283 (N_14283,N_14102,N_14029);
xnor U14284 (N_14284,N_14082,N_14128);
nor U14285 (N_14285,N_14185,N_14111);
nor U14286 (N_14286,N_14077,N_14099);
and U14287 (N_14287,N_14018,N_14148);
or U14288 (N_14288,N_14080,N_14193);
xor U14289 (N_14289,N_14196,N_14124);
nor U14290 (N_14290,N_14176,N_14072);
xor U14291 (N_14291,N_14194,N_14065);
nor U14292 (N_14292,N_14017,N_14155);
nand U14293 (N_14293,N_14000,N_14156);
nand U14294 (N_14294,N_14118,N_14070);
nor U14295 (N_14295,N_14015,N_14120);
xnor U14296 (N_14296,N_14115,N_14181);
nand U14297 (N_14297,N_14032,N_14040);
xnor U14298 (N_14298,N_14110,N_14020);
or U14299 (N_14299,N_14183,N_14068);
xor U14300 (N_14300,N_14036,N_14004);
xnor U14301 (N_14301,N_14020,N_14027);
and U14302 (N_14302,N_14149,N_14195);
nand U14303 (N_14303,N_14160,N_14041);
and U14304 (N_14304,N_14045,N_14143);
nand U14305 (N_14305,N_14006,N_14116);
and U14306 (N_14306,N_14181,N_14174);
or U14307 (N_14307,N_14067,N_14057);
nor U14308 (N_14308,N_14168,N_14005);
nand U14309 (N_14309,N_14172,N_14142);
nand U14310 (N_14310,N_14166,N_14157);
nand U14311 (N_14311,N_14135,N_14095);
xnor U14312 (N_14312,N_14181,N_14187);
and U14313 (N_14313,N_14034,N_14148);
nand U14314 (N_14314,N_14169,N_14138);
xnor U14315 (N_14315,N_14028,N_14111);
nor U14316 (N_14316,N_14174,N_14012);
xnor U14317 (N_14317,N_14012,N_14063);
xnor U14318 (N_14318,N_14115,N_14100);
xor U14319 (N_14319,N_14030,N_14027);
or U14320 (N_14320,N_14124,N_14102);
xnor U14321 (N_14321,N_14038,N_14066);
or U14322 (N_14322,N_14181,N_14126);
nand U14323 (N_14323,N_14110,N_14060);
xor U14324 (N_14324,N_14171,N_14127);
nand U14325 (N_14325,N_14128,N_14112);
xor U14326 (N_14326,N_14107,N_14197);
nor U14327 (N_14327,N_14169,N_14099);
nand U14328 (N_14328,N_14141,N_14043);
and U14329 (N_14329,N_14144,N_14180);
or U14330 (N_14330,N_14190,N_14067);
and U14331 (N_14331,N_14004,N_14035);
and U14332 (N_14332,N_14062,N_14033);
and U14333 (N_14333,N_14101,N_14017);
or U14334 (N_14334,N_14003,N_14159);
xnor U14335 (N_14335,N_14111,N_14170);
or U14336 (N_14336,N_14051,N_14059);
xnor U14337 (N_14337,N_14087,N_14021);
nor U14338 (N_14338,N_14175,N_14065);
and U14339 (N_14339,N_14122,N_14027);
xor U14340 (N_14340,N_14171,N_14036);
or U14341 (N_14341,N_14129,N_14181);
nor U14342 (N_14342,N_14055,N_14014);
xnor U14343 (N_14343,N_14163,N_14109);
or U14344 (N_14344,N_14161,N_14120);
xnor U14345 (N_14345,N_14065,N_14142);
nand U14346 (N_14346,N_14155,N_14191);
xor U14347 (N_14347,N_14097,N_14092);
nand U14348 (N_14348,N_14134,N_14043);
and U14349 (N_14349,N_14091,N_14096);
and U14350 (N_14350,N_14026,N_14169);
or U14351 (N_14351,N_14013,N_14178);
nor U14352 (N_14352,N_14151,N_14114);
and U14353 (N_14353,N_14030,N_14116);
or U14354 (N_14354,N_14123,N_14000);
nand U14355 (N_14355,N_14107,N_14032);
xor U14356 (N_14356,N_14004,N_14178);
nand U14357 (N_14357,N_14154,N_14169);
nand U14358 (N_14358,N_14093,N_14114);
and U14359 (N_14359,N_14027,N_14061);
and U14360 (N_14360,N_14050,N_14006);
nand U14361 (N_14361,N_14024,N_14101);
and U14362 (N_14362,N_14103,N_14159);
xor U14363 (N_14363,N_14142,N_14014);
nand U14364 (N_14364,N_14095,N_14042);
or U14365 (N_14365,N_14006,N_14102);
nor U14366 (N_14366,N_14141,N_14070);
and U14367 (N_14367,N_14078,N_14025);
and U14368 (N_14368,N_14070,N_14162);
and U14369 (N_14369,N_14185,N_14015);
and U14370 (N_14370,N_14134,N_14198);
xnor U14371 (N_14371,N_14112,N_14164);
nor U14372 (N_14372,N_14147,N_14187);
nand U14373 (N_14373,N_14110,N_14133);
or U14374 (N_14374,N_14152,N_14115);
xnor U14375 (N_14375,N_14046,N_14127);
nand U14376 (N_14376,N_14175,N_14121);
nand U14377 (N_14377,N_14113,N_14102);
and U14378 (N_14378,N_14035,N_14031);
nand U14379 (N_14379,N_14167,N_14125);
nand U14380 (N_14380,N_14085,N_14149);
and U14381 (N_14381,N_14097,N_14031);
nand U14382 (N_14382,N_14176,N_14079);
and U14383 (N_14383,N_14064,N_14028);
nand U14384 (N_14384,N_14051,N_14114);
nand U14385 (N_14385,N_14116,N_14001);
xnor U14386 (N_14386,N_14161,N_14071);
xor U14387 (N_14387,N_14169,N_14061);
and U14388 (N_14388,N_14063,N_14177);
xor U14389 (N_14389,N_14026,N_14093);
nor U14390 (N_14390,N_14049,N_14193);
nor U14391 (N_14391,N_14165,N_14194);
and U14392 (N_14392,N_14010,N_14184);
nor U14393 (N_14393,N_14150,N_14034);
nor U14394 (N_14394,N_14063,N_14021);
or U14395 (N_14395,N_14010,N_14073);
or U14396 (N_14396,N_14151,N_14104);
or U14397 (N_14397,N_14187,N_14039);
nor U14398 (N_14398,N_14126,N_14190);
or U14399 (N_14399,N_14041,N_14199);
and U14400 (N_14400,N_14324,N_14227);
nand U14401 (N_14401,N_14240,N_14237);
nand U14402 (N_14402,N_14326,N_14226);
and U14403 (N_14403,N_14362,N_14220);
and U14404 (N_14404,N_14385,N_14327);
nor U14405 (N_14405,N_14278,N_14300);
nor U14406 (N_14406,N_14358,N_14242);
nor U14407 (N_14407,N_14205,N_14332);
xnor U14408 (N_14408,N_14233,N_14393);
nand U14409 (N_14409,N_14276,N_14222);
nor U14410 (N_14410,N_14335,N_14284);
nand U14411 (N_14411,N_14361,N_14244);
or U14412 (N_14412,N_14387,N_14263);
and U14413 (N_14413,N_14316,N_14225);
xnor U14414 (N_14414,N_14368,N_14345);
and U14415 (N_14415,N_14396,N_14304);
nand U14416 (N_14416,N_14252,N_14312);
or U14417 (N_14417,N_14323,N_14265);
nand U14418 (N_14418,N_14365,N_14218);
nand U14419 (N_14419,N_14319,N_14201);
xor U14420 (N_14420,N_14260,N_14357);
and U14421 (N_14421,N_14350,N_14337);
xor U14422 (N_14422,N_14334,N_14229);
or U14423 (N_14423,N_14208,N_14318);
nor U14424 (N_14424,N_14303,N_14230);
nor U14425 (N_14425,N_14247,N_14207);
xor U14426 (N_14426,N_14214,N_14235);
nor U14427 (N_14427,N_14363,N_14259);
and U14428 (N_14428,N_14277,N_14353);
nor U14429 (N_14429,N_14287,N_14272);
nor U14430 (N_14430,N_14397,N_14296);
and U14431 (N_14431,N_14254,N_14266);
and U14432 (N_14432,N_14267,N_14338);
or U14433 (N_14433,N_14269,N_14355);
xnor U14434 (N_14434,N_14360,N_14389);
xor U14435 (N_14435,N_14271,N_14394);
or U14436 (N_14436,N_14383,N_14221);
or U14437 (N_14437,N_14313,N_14307);
nand U14438 (N_14438,N_14314,N_14322);
and U14439 (N_14439,N_14372,N_14224);
and U14440 (N_14440,N_14380,N_14391);
xor U14441 (N_14441,N_14234,N_14399);
and U14442 (N_14442,N_14274,N_14333);
nor U14443 (N_14443,N_14211,N_14329);
nor U14444 (N_14444,N_14348,N_14310);
or U14445 (N_14445,N_14289,N_14308);
or U14446 (N_14446,N_14305,N_14299);
and U14447 (N_14447,N_14342,N_14306);
xor U14448 (N_14448,N_14210,N_14309);
and U14449 (N_14449,N_14204,N_14253);
nand U14450 (N_14450,N_14258,N_14216);
nor U14451 (N_14451,N_14370,N_14341);
and U14452 (N_14452,N_14371,N_14275);
xor U14453 (N_14453,N_14291,N_14261);
nand U14454 (N_14454,N_14364,N_14320);
nand U14455 (N_14455,N_14283,N_14301);
xor U14456 (N_14456,N_14395,N_14328);
and U14457 (N_14457,N_14325,N_14336);
nand U14458 (N_14458,N_14213,N_14366);
or U14459 (N_14459,N_14228,N_14206);
or U14460 (N_14460,N_14398,N_14349);
nor U14461 (N_14461,N_14251,N_14264);
nor U14462 (N_14462,N_14273,N_14203);
or U14463 (N_14463,N_14331,N_14217);
nor U14464 (N_14464,N_14382,N_14285);
xor U14465 (N_14465,N_14256,N_14293);
nor U14466 (N_14466,N_14209,N_14347);
and U14467 (N_14467,N_14317,N_14352);
xnor U14468 (N_14468,N_14238,N_14250);
xor U14469 (N_14469,N_14354,N_14290);
and U14470 (N_14470,N_14231,N_14257);
or U14471 (N_14471,N_14281,N_14268);
nand U14472 (N_14472,N_14315,N_14239);
and U14473 (N_14473,N_14330,N_14374);
nand U14474 (N_14474,N_14241,N_14367);
nand U14475 (N_14475,N_14294,N_14249);
nand U14476 (N_14476,N_14245,N_14339);
nand U14477 (N_14477,N_14248,N_14270);
xor U14478 (N_14478,N_14351,N_14298);
nand U14479 (N_14479,N_14375,N_14340);
or U14480 (N_14480,N_14288,N_14386);
and U14481 (N_14481,N_14388,N_14302);
nor U14482 (N_14482,N_14356,N_14279);
xnor U14483 (N_14483,N_14311,N_14215);
and U14484 (N_14484,N_14286,N_14202);
nor U14485 (N_14485,N_14381,N_14292);
and U14486 (N_14486,N_14390,N_14321);
xnor U14487 (N_14487,N_14384,N_14243);
xnor U14488 (N_14488,N_14236,N_14212);
and U14489 (N_14489,N_14378,N_14376);
or U14490 (N_14490,N_14379,N_14200);
xnor U14491 (N_14491,N_14359,N_14343);
xnor U14492 (N_14492,N_14346,N_14377);
nor U14493 (N_14493,N_14369,N_14392);
or U14494 (N_14494,N_14344,N_14219);
nand U14495 (N_14495,N_14255,N_14295);
nand U14496 (N_14496,N_14280,N_14282);
xnor U14497 (N_14497,N_14373,N_14246);
or U14498 (N_14498,N_14297,N_14262);
nand U14499 (N_14499,N_14232,N_14223);
nand U14500 (N_14500,N_14330,N_14267);
or U14501 (N_14501,N_14389,N_14288);
xnor U14502 (N_14502,N_14376,N_14280);
xnor U14503 (N_14503,N_14282,N_14390);
nand U14504 (N_14504,N_14357,N_14362);
and U14505 (N_14505,N_14242,N_14394);
xnor U14506 (N_14506,N_14306,N_14244);
xnor U14507 (N_14507,N_14253,N_14332);
and U14508 (N_14508,N_14268,N_14363);
or U14509 (N_14509,N_14317,N_14344);
and U14510 (N_14510,N_14256,N_14236);
or U14511 (N_14511,N_14382,N_14286);
and U14512 (N_14512,N_14319,N_14274);
and U14513 (N_14513,N_14353,N_14268);
xnor U14514 (N_14514,N_14294,N_14271);
nor U14515 (N_14515,N_14397,N_14339);
xor U14516 (N_14516,N_14210,N_14367);
and U14517 (N_14517,N_14235,N_14376);
nor U14518 (N_14518,N_14253,N_14242);
or U14519 (N_14519,N_14218,N_14345);
nor U14520 (N_14520,N_14365,N_14214);
nor U14521 (N_14521,N_14260,N_14373);
and U14522 (N_14522,N_14336,N_14398);
xnor U14523 (N_14523,N_14297,N_14290);
nand U14524 (N_14524,N_14207,N_14278);
nor U14525 (N_14525,N_14276,N_14263);
xor U14526 (N_14526,N_14321,N_14209);
or U14527 (N_14527,N_14246,N_14371);
or U14528 (N_14528,N_14295,N_14297);
and U14529 (N_14529,N_14312,N_14355);
and U14530 (N_14530,N_14207,N_14385);
xnor U14531 (N_14531,N_14338,N_14248);
or U14532 (N_14532,N_14390,N_14337);
nor U14533 (N_14533,N_14376,N_14325);
nand U14534 (N_14534,N_14251,N_14281);
nand U14535 (N_14535,N_14377,N_14200);
nor U14536 (N_14536,N_14371,N_14216);
nor U14537 (N_14537,N_14288,N_14283);
or U14538 (N_14538,N_14206,N_14220);
and U14539 (N_14539,N_14279,N_14375);
xor U14540 (N_14540,N_14335,N_14361);
nand U14541 (N_14541,N_14380,N_14399);
xnor U14542 (N_14542,N_14231,N_14370);
nor U14543 (N_14543,N_14374,N_14301);
nand U14544 (N_14544,N_14386,N_14257);
or U14545 (N_14545,N_14274,N_14202);
or U14546 (N_14546,N_14346,N_14231);
nor U14547 (N_14547,N_14248,N_14233);
and U14548 (N_14548,N_14316,N_14383);
nand U14549 (N_14549,N_14352,N_14256);
nor U14550 (N_14550,N_14391,N_14363);
nand U14551 (N_14551,N_14270,N_14373);
xor U14552 (N_14552,N_14357,N_14274);
or U14553 (N_14553,N_14241,N_14394);
nand U14554 (N_14554,N_14202,N_14238);
nand U14555 (N_14555,N_14338,N_14306);
and U14556 (N_14556,N_14299,N_14374);
and U14557 (N_14557,N_14334,N_14304);
nand U14558 (N_14558,N_14219,N_14313);
nand U14559 (N_14559,N_14349,N_14378);
or U14560 (N_14560,N_14225,N_14350);
and U14561 (N_14561,N_14363,N_14300);
nor U14562 (N_14562,N_14213,N_14261);
nor U14563 (N_14563,N_14267,N_14318);
or U14564 (N_14564,N_14229,N_14296);
xor U14565 (N_14565,N_14397,N_14209);
and U14566 (N_14566,N_14247,N_14385);
or U14567 (N_14567,N_14332,N_14398);
or U14568 (N_14568,N_14372,N_14237);
xnor U14569 (N_14569,N_14334,N_14321);
xor U14570 (N_14570,N_14348,N_14261);
nor U14571 (N_14571,N_14395,N_14320);
or U14572 (N_14572,N_14336,N_14309);
xnor U14573 (N_14573,N_14250,N_14242);
nor U14574 (N_14574,N_14279,N_14350);
xor U14575 (N_14575,N_14243,N_14216);
or U14576 (N_14576,N_14341,N_14242);
nor U14577 (N_14577,N_14279,N_14336);
nand U14578 (N_14578,N_14293,N_14360);
nor U14579 (N_14579,N_14312,N_14399);
nand U14580 (N_14580,N_14338,N_14337);
or U14581 (N_14581,N_14354,N_14393);
xnor U14582 (N_14582,N_14326,N_14384);
and U14583 (N_14583,N_14319,N_14383);
nor U14584 (N_14584,N_14365,N_14307);
xor U14585 (N_14585,N_14248,N_14207);
and U14586 (N_14586,N_14321,N_14320);
xor U14587 (N_14587,N_14307,N_14236);
xnor U14588 (N_14588,N_14327,N_14384);
or U14589 (N_14589,N_14391,N_14378);
nand U14590 (N_14590,N_14239,N_14368);
and U14591 (N_14591,N_14365,N_14278);
nor U14592 (N_14592,N_14296,N_14228);
and U14593 (N_14593,N_14395,N_14383);
and U14594 (N_14594,N_14380,N_14245);
or U14595 (N_14595,N_14377,N_14270);
or U14596 (N_14596,N_14358,N_14331);
or U14597 (N_14597,N_14305,N_14332);
nor U14598 (N_14598,N_14310,N_14292);
and U14599 (N_14599,N_14378,N_14335);
xnor U14600 (N_14600,N_14496,N_14541);
nor U14601 (N_14601,N_14431,N_14586);
or U14602 (N_14602,N_14515,N_14444);
nor U14603 (N_14603,N_14504,N_14443);
and U14604 (N_14604,N_14570,N_14451);
nand U14605 (N_14605,N_14582,N_14421);
or U14606 (N_14606,N_14539,N_14538);
nand U14607 (N_14607,N_14433,N_14599);
nand U14608 (N_14608,N_14470,N_14412);
and U14609 (N_14609,N_14467,N_14502);
or U14610 (N_14610,N_14516,N_14523);
xor U14611 (N_14611,N_14559,N_14505);
nor U14612 (N_14612,N_14514,N_14474);
nor U14613 (N_14613,N_14580,N_14503);
nand U14614 (N_14614,N_14456,N_14486);
nand U14615 (N_14615,N_14400,N_14551);
xor U14616 (N_14616,N_14497,N_14445);
xor U14617 (N_14617,N_14557,N_14425);
nor U14618 (N_14618,N_14415,N_14552);
xnor U14619 (N_14619,N_14487,N_14490);
nor U14620 (N_14620,N_14481,N_14519);
nand U14621 (N_14621,N_14578,N_14404);
nand U14622 (N_14622,N_14528,N_14436);
xnor U14623 (N_14623,N_14597,N_14583);
xor U14624 (N_14624,N_14414,N_14563);
nor U14625 (N_14625,N_14418,N_14524);
or U14626 (N_14626,N_14475,N_14413);
and U14627 (N_14627,N_14430,N_14408);
xnor U14628 (N_14628,N_14464,N_14417);
and U14629 (N_14629,N_14527,N_14498);
xor U14630 (N_14630,N_14457,N_14401);
or U14631 (N_14631,N_14458,N_14427);
xor U14632 (N_14632,N_14405,N_14591);
nand U14633 (N_14633,N_14598,N_14542);
or U14634 (N_14634,N_14564,N_14419);
nor U14635 (N_14635,N_14403,N_14536);
or U14636 (N_14636,N_14495,N_14587);
or U14637 (N_14637,N_14543,N_14416);
nand U14638 (N_14638,N_14531,N_14589);
nand U14639 (N_14639,N_14499,N_14548);
xor U14640 (N_14640,N_14571,N_14535);
nand U14641 (N_14641,N_14555,N_14500);
nor U14642 (N_14642,N_14459,N_14522);
and U14643 (N_14643,N_14572,N_14466);
xor U14644 (N_14644,N_14521,N_14573);
nand U14645 (N_14645,N_14429,N_14480);
or U14646 (N_14646,N_14455,N_14406);
nand U14647 (N_14647,N_14491,N_14526);
nor U14648 (N_14648,N_14460,N_14529);
nor U14649 (N_14649,N_14593,N_14574);
nand U14650 (N_14650,N_14410,N_14549);
nor U14651 (N_14651,N_14492,N_14588);
and U14652 (N_14652,N_14442,N_14435);
nor U14653 (N_14653,N_14512,N_14510);
or U14654 (N_14654,N_14447,N_14450);
or U14655 (N_14655,N_14452,N_14440);
nand U14656 (N_14656,N_14411,N_14508);
nor U14657 (N_14657,N_14509,N_14546);
and U14658 (N_14658,N_14566,N_14553);
and U14659 (N_14659,N_14585,N_14517);
and U14660 (N_14660,N_14596,N_14463);
xnor U14661 (N_14661,N_14488,N_14465);
nor U14662 (N_14662,N_14544,N_14432);
xor U14663 (N_14663,N_14560,N_14507);
and U14664 (N_14664,N_14562,N_14550);
or U14665 (N_14665,N_14407,N_14484);
xor U14666 (N_14666,N_14477,N_14468);
and U14667 (N_14667,N_14511,N_14462);
and U14668 (N_14668,N_14489,N_14426);
nand U14669 (N_14669,N_14449,N_14434);
and U14670 (N_14670,N_14420,N_14556);
xor U14671 (N_14671,N_14590,N_14422);
xor U14672 (N_14672,N_14575,N_14479);
nor U14673 (N_14673,N_14584,N_14437);
and U14674 (N_14674,N_14554,N_14438);
nor U14675 (N_14675,N_14561,N_14469);
or U14676 (N_14676,N_14592,N_14506);
or U14677 (N_14677,N_14423,N_14446);
nor U14678 (N_14678,N_14476,N_14409);
and U14679 (N_14679,N_14494,N_14472);
nand U14680 (N_14680,N_14534,N_14565);
and U14681 (N_14681,N_14547,N_14473);
nand U14682 (N_14682,N_14483,N_14533);
xor U14683 (N_14683,N_14518,N_14558);
or U14684 (N_14684,N_14594,N_14577);
or U14685 (N_14685,N_14428,N_14540);
xor U14686 (N_14686,N_14485,N_14454);
nand U14687 (N_14687,N_14441,N_14501);
nor U14688 (N_14688,N_14579,N_14532);
xor U14689 (N_14689,N_14471,N_14520);
xor U14690 (N_14690,N_14424,N_14530);
nor U14691 (N_14691,N_14439,N_14537);
xor U14692 (N_14692,N_14576,N_14568);
nand U14693 (N_14693,N_14461,N_14595);
xor U14694 (N_14694,N_14581,N_14448);
nand U14695 (N_14695,N_14478,N_14569);
and U14696 (N_14696,N_14493,N_14402);
or U14697 (N_14697,N_14567,N_14482);
or U14698 (N_14698,N_14453,N_14513);
nand U14699 (N_14699,N_14545,N_14525);
or U14700 (N_14700,N_14471,N_14525);
nor U14701 (N_14701,N_14452,N_14516);
nor U14702 (N_14702,N_14512,N_14545);
and U14703 (N_14703,N_14470,N_14523);
or U14704 (N_14704,N_14404,N_14496);
and U14705 (N_14705,N_14463,N_14439);
nand U14706 (N_14706,N_14468,N_14416);
nand U14707 (N_14707,N_14525,N_14577);
xor U14708 (N_14708,N_14516,N_14419);
nand U14709 (N_14709,N_14559,N_14563);
xor U14710 (N_14710,N_14433,N_14414);
or U14711 (N_14711,N_14540,N_14400);
nand U14712 (N_14712,N_14560,N_14556);
nand U14713 (N_14713,N_14514,N_14449);
and U14714 (N_14714,N_14521,N_14485);
xor U14715 (N_14715,N_14539,N_14461);
and U14716 (N_14716,N_14564,N_14489);
nor U14717 (N_14717,N_14565,N_14556);
and U14718 (N_14718,N_14411,N_14526);
xor U14719 (N_14719,N_14507,N_14581);
or U14720 (N_14720,N_14496,N_14465);
or U14721 (N_14721,N_14424,N_14433);
nor U14722 (N_14722,N_14558,N_14483);
and U14723 (N_14723,N_14514,N_14454);
nand U14724 (N_14724,N_14530,N_14504);
nor U14725 (N_14725,N_14457,N_14555);
nor U14726 (N_14726,N_14460,N_14555);
and U14727 (N_14727,N_14584,N_14519);
and U14728 (N_14728,N_14415,N_14512);
nand U14729 (N_14729,N_14560,N_14449);
nor U14730 (N_14730,N_14524,N_14456);
xor U14731 (N_14731,N_14539,N_14449);
or U14732 (N_14732,N_14555,N_14502);
nor U14733 (N_14733,N_14483,N_14597);
xor U14734 (N_14734,N_14443,N_14561);
xor U14735 (N_14735,N_14427,N_14424);
and U14736 (N_14736,N_14539,N_14472);
and U14737 (N_14737,N_14475,N_14524);
nand U14738 (N_14738,N_14530,N_14532);
or U14739 (N_14739,N_14599,N_14569);
xnor U14740 (N_14740,N_14523,N_14522);
nor U14741 (N_14741,N_14556,N_14406);
nand U14742 (N_14742,N_14477,N_14473);
or U14743 (N_14743,N_14408,N_14567);
nor U14744 (N_14744,N_14422,N_14538);
and U14745 (N_14745,N_14560,N_14498);
or U14746 (N_14746,N_14418,N_14502);
xor U14747 (N_14747,N_14598,N_14514);
or U14748 (N_14748,N_14462,N_14441);
and U14749 (N_14749,N_14415,N_14409);
nor U14750 (N_14750,N_14447,N_14548);
xor U14751 (N_14751,N_14476,N_14515);
or U14752 (N_14752,N_14483,N_14466);
nand U14753 (N_14753,N_14447,N_14452);
xor U14754 (N_14754,N_14461,N_14436);
and U14755 (N_14755,N_14475,N_14462);
nor U14756 (N_14756,N_14569,N_14523);
nand U14757 (N_14757,N_14562,N_14563);
nand U14758 (N_14758,N_14498,N_14400);
and U14759 (N_14759,N_14421,N_14461);
nor U14760 (N_14760,N_14581,N_14565);
and U14761 (N_14761,N_14544,N_14448);
nand U14762 (N_14762,N_14465,N_14455);
xor U14763 (N_14763,N_14589,N_14480);
nor U14764 (N_14764,N_14540,N_14452);
or U14765 (N_14765,N_14497,N_14545);
or U14766 (N_14766,N_14529,N_14493);
and U14767 (N_14767,N_14518,N_14560);
and U14768 (N_14768,N_14410,N_14541);
and U14769 (N_14769,N_14563,N_14478);
nor U14770 (N_14770,N_14575,N_14570);
xor U14771 (N_14771,N_14531,N_14481);
nor U14772 (N_14772,N_14535,N_14475);
nand U14773 (N_14773,N_14485,N_14402);
and U14774 (N_14774,N_14404,N_14568);
or U14775 (N_14775,N_14468,N_14448);
nand U14776 (N_14776,N_14511,N_14555);
xor U14777 (N_14777,N_14464,N_14499);
or U14778 (N_14778,N_14557,N_14537);
and U14779 (N_14779,N_14585,N_14480);
and U14780 (N_14780,N_14402,N_14575);
xnor U14781 (N_14781,N_14527,N_14562);
and U14782 (N_14782,N_14465,N_14447);
nor U14783 (N_14783,N_14489,N_14562);
nor U14784 (N_14784,N_14454,N_14538);
nand U14785 (N_14785,N_14540,N_14414);
nand U14786 (N_14786,N_14486,N_14414);
nand U14787 (N_14787,N_14473,N_14478);
xnor U14788 (N_14788,N_14437,N_14451);
nor U14789 (N_14789,N_14424,N_14527);
xnor U14790 (N_14790,N_14564,N_14542);
and U14791 (N_14791,N_14575,N_14487);
or U14792 (N_14792,N_14516,N_14530);
nand U14793 (N_14793,N_14447,N_14466);
and U14794 (N_14794,N_14418,N_14578);
nand U14795 (N_14795,N_14484,N_14412);
and U14796 (N_14796,N_14510,N_14473);
nand U14797 (N_14797,N_14429,N_14477);
nor U14798 (N_14798,N_14476,N_14540);
or U14799 (N_14799,N_14489,N_14491);
nand U14800 (N_14800,N_14779,N_14692);
xor U14801 (N_14801,N_14631,N_14797);
and U14802 (N_14802,N_14737,N_14796);
and U14803 (N_14803,N_14775,N_14665);
nand U14804 (N_14804,N_14622,N_14697);
xor U14805 (N_14805,N_14751,N_14689);
xor U14806 (N_14806,N_14722,N_14619);
or U14807 (N_14807,N_14641,N_14792);
nand U14808 (N_14808,N_14788,N_14648);
or U14809 (N_14809,N_14761,N_14770);
nand U14810 (N_14810,N_14702,N_14752);
nand U14811 (N_14811,N_14618,N_14623);
nand U14812 (N_14812,N_14759,N_14744);
nor U14813 (N_14813,N_14704,N_14762);
nand U14814 (N_14814,N_14705,N_14671);
xnor U14815 (N_14815,N_14636,N_14670);
xor U14816 (N_14816,N_14763,N_14643);
nor U14817 (N_14817,N_14718,N_14611);
nand U14818 (N_14818,N_14633,N_14728);
xor U14819 (N_14819,N_14601,N_14615);
or U14820 (N_14820,N_14773,N_14652);
and U14821 (N_14821,N_14666,N_14676);
nand U14822 (N_14822,N_14659,N_14644);
and U14823 (N_14823,N_14774,N_14607);
nor U14824 (N_14824,N_14629,N_14683);
or U14825 (N_14825,N_14771,N_14677);
or U14826 (N_14826,N_14639,N_14700);
and U14827 (N_14827,N_14725,N_14767);
or U14828 (N_14828,N_14664,N_14793);
nand U14829 (N_14829,N_14707,N_14685);
xor U14830 (N_14830,N_14701,N_14711);
xnor U14831 (N_14831,N_14777,N_14749);
nand U14832 (N_14832,N_14794,N_14758);
and U14833 (N_14833,N_14731,N_14772);
nor U14834 (N_14834,N_14778,N_14694);
nand U14835 (N_14835,N_14742,N_14653);
nor U14836 (N_14836,N_14745,N_14613);
or U14837 (N_14837,N_14733,N_14717);
nor U14838 (N_14838,N_14612,N_14712);
or U14839 (N_14839,N_14790,N_14709);
nor U14840 (N_14840,N_14706,N_14624);
nor U14841 (N_14841,N_14651,N_14713);
and U14842 (N_14842,N_14635,N_14691);
xor U14843 (N_14843,N_14736,N_14739);
xnor U14844 (N_14844,N_14663,N_14650);
nor U14845 (N_14845,N_14721,N_14795);
xnor U14846 (N_14846,N_14687,N_14646);
nor U14847 (N_14847,N_14740,N_14634);
xnor U14848 (N_14848,N_14708,N_14724);
nand U14849 (N_14849,N_14656,N_14746);
xnor U14850 (N_14850,N_14757,N_14783);
and U14851 (N_14851,N_14764,N_14786);
xnor U14852 (N_14852,N_14630,N_14662);
and U14853 (N_14853,N_14696,N_14698);
or U14854 (N_14854,N_14603,N_14715);
nor U14855 (N_14855,N_14682,N_14628);
and U14856 (N_14856,N_14620,N_14750);
nor U14857 (N_14857,N_14781,N_14710);
nand U14858 (N_14858,N_14719,N_14765);
or U14859 (N_14859,N_14784,N_14753);
xor U14860 (N_14860,N_14610,N_14727);
nand U14861 (N_14861,N_14743,N_14649);
and U14862 (N_14862,N_14729,N_14734);
or U14863 (N_14863,N_14616,N_14681);
nor U14864 (N_14864,N_14787,N_14695);
and U14865 (N_14865,N_14632,N_14627);
or U14866 (N_14866,N_14686,N_14768);
or U14867 (N_14867,N_14769,N_14798);
and U14868 (N_14868,N_14614,N_14608);
or U14869 (N_14869,N_14720,N_14638);
xor U14870 (N_14870,N_14658,N_14688);
xor U14871 (N_14871,N_14675,N_14645);
xor U14872 (N_14872,N_14660,N_14657);
nand U14873 (N_14873,N_14637,N_14680);
nand U14874 (N_14874,N_14785,N_14791);
nor U14875 (N_14875,N_14716,N_14766);
nand U14876 (N_14876,N_14754,N_14723);
and U14877 (N_14877,N_14626,N_14735);
nand U14878 (N_14878,N_14789,N_14693);
and U14879 (N_14879,N_14782,N_14776);
nor U14880 (N_14880,N_14741,N_14655);
and U14881 (N_14881,N_14690,N_14609);
xnor U14882 (N_14882,N_14760,N_14604);
nand U14883 (N_14883,N_14780,N_14640);
or U14884 (N_14884,N_14654,N_14730);
or U14885 (N_14885,N_14748,N_14661);
nor U14886 (N_14886,N_14600,N_14747);
nand U14887 (N_14887,N_14647,N_14738);
and U14888 (N_14888,N_14642,N_14667);
xnor U14889 (N_14889,N_14621,N_14678);
nor U14890 (N_14890,N_14732,N_14625);
nand U14891 (N_14891,N_14799,N_14714);
xnor U14892 (N_14892,N_14602,N_14605);
nand U14893 (N_14893,N_14755,N_14617);
nor U14894 (N_14894,N_14756,N_14606);
xnor U14895 (N_14895,N_14669,N_14679);
nand U14896 (N_14896,N_14668,N_14672);
and U14897 (N_14897,N_14684,N_14703);
or U14898 (N_14898,N_14726,N_14674);
or U14899 (N_14899,N_14673,N_14699);
or U14900 (N_14900,N_14637,N_14634);
and U14901 (N_14901,N_14644,N_14791);
and U14902 (N_14902,N_14791,N_14717);
or U14903 (N_14903,N_14754,N_14788);
and U14904 (N_14904,N_14625,N_14698);
xnor U14905 (N_14905,N_14752,N_14718);
nor U14906 (N_14906,N_14694,N_14776);
and U14907 (N_14907,N_14712,N_14669);
xnor U14908 (N_14908,N_14753,N_14676);
nor U14909 (N_14909,N_14709,N_14714);
or U14910 (N_14910,N_14795,N_14708);
xnor U14911 (N_14911,N_14677,N_14712);
and U14912 (N_14912,N_14796,N_14732);
or U14913 (N_14913,N_14754,N_14643);
nand U14914 (N_14914,N_14634,N_14688);
nor U14915 (N_14915,N_14679,N_14626);
nor U14916 (N_14916,N_14792,N_14653);
nand U14917 (N_14917,N_14614,N_14747);
nand U14918 (N_14918,N_14610,N_14622);
xor U14919 (N_14919,N_14656,N_14676);
nand U14920 (N_14920,N_14737,N_14698);
nor U14921 (N_14921,N_14785,N_14762);
nor U14922 (N_14922,N_14634,N_14645);
nor U14923 (N_14923,N_14679,N_14768);
and U14924 (N_14924,N_14787,N_14762);
xor U14925 (N_14925,N_14745,N_14650);
xor U14926 (N_14926,N_14678,N_14653);
or U14927 (N_14927,N_14691,N_14619);
nor U14928 (N_14928,N_14782,N_14676);
and U14929 (N_14929,N_14772,N_14632);
xnor U14930 (N_14930,N_14658,N_14743);
or U14931 (N_14931,N_14641,N_14640);
nor U14932 (N_14932,N_14626,N_14607);
nor U14933 (N_14933,N_14680,N_14738);
or U14934 (N_14934,N_14650,N_14746);
nand U14935 (N_14935,N_14770,N_14723);
nand U14936 (N_14936,N_14724,N_14670);
nor U14937 (N_14937,N_14643,N_14740);
nand U14938 (N_14938,N_14678,N_14746);
nor U14939 (N_14939,N_14676,N_14683);
nand U14940 (N_14940,N_14667,N_14608);
nand U14941 (N_14941,N_14792,N_14654);
or U14942 (N_14942,N_14629,N_14625);
nor U14943 (N_14943,N_14662,N_14692);
nand U14944 (N_14944,N_14687,N_14641);
nand U14945 (N_14945,N_14722,N_14740);
xor U14946 (N_14946,N_14677,N_14706);
xor U14947 (N_14947,N_14611,N_14796);
xor U14948 (N_14948,N_14770,N_14710);
xor U14949 (N_14949,N_14600,N_14677);
xor U14950 (N_14950,N_14685,N_14700);
xor U14951 (N_14951,N_14717,N_14702);
or U14952 (N_14952,N_14667,N_14657);
or U14953 (N_14953,N_14621,N_14785);
nand U14954 (N_14954,N_14772,N_14622);
nor U14955 (N_14955,N_14697,N_14653);
xnor U14956 (N_14956,N_14789,N_14715);
or U14957 (N_14957,N_14601,N_14772);
or U14958 (N_14958,N_14669,N_14642);
nand U14959 (N_14959,N_14607,N_14754);
and U14960 (N_14960,N_14714,N_14613);
or U14961 (N_14961,N_14638,N_14660);
or U14962 (N_14962,N_14630,N_14691);
and U14963 (N_14963,N_14798,N_14647);
or U14964 (N_14964,N_14723,N_14771);
nor U14965 (N_14965,N_14698,N_14729);
or U14966 (N_14966,N_14744,N_14603);
or U14967 (N_14967,N_14715,N_14757);
and U14968 (N_14968,N_14764,N_14749);
and U14969 (N_14969,N_14634,N_14773);
or U14970 (N_14970,N_14685,N_14634);
xor U14971 (N_14971,N_14694,N_14749);
nand U14972 (N_14972,N_14739,N_14752);
xor U14973 (N_14973,N_14753,N_14757);
nor U14974 (N_14974,N_14626,N_14677);
nand U14975 (N_14975,N_14774,N_14766);
or U14976 (N_14976,N_14729,N_14696);
or U14977 (N_14977,N_14608,N_14660);
and U14978 (N_14978,N_14660,N_14793);
nor U14979 (N_14979,N_14712,N_14643);
nand U14980 (N_14980,N_14663,N_14708);
or U14981 (N_14981,N_14770,N_14736);
nor U14982 (N_14982,N_14624,N_14659);
and U14983 (N_14983,N_14655,N_14707);
and U14984 (N_14984,N_14764,N_14665);
xor U14985 (N_14985,N_14795,N_14738);
nand U14986 (N_14986,N_14774,N_14665);
or U14987 (N_14987,N_14700,N_14705);
and U14988 (N_14988,N_14705,N_14752);
and U14989 (N_14989,N_14673,N_14779);
nand U14990 (N_14990,N_14731,N_14740);
nor U14991 (N_14991,N_14702,N_14780);
and U14992 (N_14992,N_14684,N_14632);
nand U14993 (N_14993,N_14718,N_14663);
xor U14994 (N_14994,N_14649,N_14659);
xnor U14995 (N_14995,N_14726,N_14702);
or U14996 (N_14996,N_14790,N_14665);
and U14997 (N_14997,N_14602,N_14729);
xnor U14998 (N_14998,N_14689,N_14757);
xnor U14999 (N_14999,N_14625,N_14669);
nand UO_0 (O_0,N_14924,N_14826);
or UO_1 (O_1,N_14834,N_14897);
nand UO_2 (O_2,N_14856,N_14864);
nor UO_3 (O_3,N_14860,N_14938);
xnor UO_4 (O_4,N_14997,N_14937);
or UO_5 (O_5,N_14979,N_14889);
and UO_6 (O_6,N_14893,N_14849);
nor UO_7 (O_7,N_14885,N_14944);
nor UO_8 (O_8,N_14802,N_14887);
xor UO_9 (O_9,N_14961,N_14874);
nand UO_10 (O_10,N_14950,N_14854);
xor UO_11 (O_11,N_14814,N_14931);
xor UO_12 (O_12,N_14913,N_14884);
nor UO_13 (O_13,N_14907,N_14993);
nand UO_14 (O_14,N_14922,N_14832);
and UO_15 (O_15,N_14844,N_14925);
and UO_16 (O_16,N_14878,N_14911);
nand UO_17 (O_17,N_14951,N_14901);
nand UO_18 (O_18,N_14984,N_14862);
or UO_19 (O_19,N_14936,N_14857);
or UO_20 (O_20,N_14945,N_14977);
nand UO_21 (O_21,N_14859,N_14808);
nor UO_22 (O_22,N_14833,N_14890);
nor UO_23 (O_23,N_14960,N_14918);
or UO_24 (O_24,N_14914,N_14953);
nor UO_25 (O_25,N_14866,N_14847);
or UO_26 (O_26,N_14822,N_14837);
nand UO_27 (O_27,N_14989,N_14980);
xor UO_28 (O_28,N_14910,N_14900);
and UO_29 (O_29,N_14823,N_14962);
nand UO_30 (O_30,N_14933,N_14899);
and UO_31 (O_31,N_14916,N_14992);
nor UO_32 (O_32,N_14972,N_14829);
nor UO_33 (O_33,N_14948,N_14982);
nand UO_34 (O_34,N_14846,N_14927);
nand UO_35 (O_35,N_14963,N_14958);
nand UO_36 (O_36,N_14881,N_14836);
and UO_37 (O_37,N_14942,N_14816);
nand UO_38 (O_38,N_14895,N_14880);
xor UO_39 (O_39,N_14845,N_14800);
or UO_40 (O_40,N_14828,N_14805);
xnor UO_41 (O_41,N_14801,N_14988);
or UO_42 (O_42,N_14850,N_14956);
and UO_43 (O_43,N_14926,N_14838);
nand UO_44 (O_44,N_14912,N_14919);
nor UO_45 (O_45,N_14873,N_14966);
and UO_46 (O_46,N_14921,N_14842);
nand UO_47 (O_47,N_14812,N_14939);
nand UO_48 (O_48,N_14985,N_14915);
nor UO_49 (O_49,N_14908,N_14923);
and UO_50 (O_50,N_14870,N_14806);
and UO_51 (O_51,N_14820,N_14947);
or UO_52 (O_52,N_14848,N_14970);
and UO_53 (O_53,N_14883,N_14855);
xor UO_54 (O_54,N_14902,N_14903);
or UO_55 (O_55,N_14949,N_14898);
xor UO_56 (O_56,N_14957,N_14803);
or UO_57 (O_57,N_14818,N_14930);
or UO_58 (O_58,N_14819,N_14810);
xor UO_59 (O_59,N_14978,N_14981);
xor UO_60 (O_60,N_14813,N_14943);
or UO_61 (O_61,N_14817,N_14959);
and UO_62 (O_62,N_14941,N_14967);
nor UO_63 (O_63,N_14867,N_14995);
and UO_64 (O_64,N_14882,N_14971);
nor UO_65 (O_65,N_14886,N_14876);
and UO_66 (O_66,N_14888,N_14852);
xor UO_67 (O_67,N_14917,N_14894);
nand UO_68 (O_68,N_14969,N_14973);
or UO_69 (O_69,N_14875,N_14872);
or UO_70 (O_70,N_14983,N_14807);
nor UO_71 (O_71,N_14935,N_14928);
nand UO_72 (O_72,N_14974,N_14904);
nand UO_73 (O_73,N_14879,N_14934);
nand UO_74 (O_74,N_14965,N_14858);
xnor UO_75 (O_75,N_14835,N_14841);
and UO_76 (O_76,N_14861,N_14853);
nand UO_77 (O_77,N_14843,N_14809);
xnor UO_78 (O_78,N_14906,N_14955);
nor UO_79 (O_79,N_14804,N_14998);
xnor UO_80 (O_80,N_14987,N_14891);
nand UO_81 (O_81,N_14869,N_14840);
nand UO_82 (O_82,N_14964,N_14892);
nor UO_83 (O_83,N_14868,N_14896);
or UO_84 (O_84,N_14986,N_14920);
and UO_85 (O_85,N_14905,N_14940);
nor UO_86 (O_86,N_14811,N_14929);
and UO_87 (O_87,N_14825,N_14821);
nor UO_88 (O_88,N_14839,N_14827);
nor UO_89 (O_89,N_14996,N_14954);
nor UO_90 (O_90,N_14952,N_14909);
nand UO_91 (O_91,N_14865,N_14975);
xor UO_92 (O_92,N_14976,N_14863);
nand UO_93 (O_93,N_14871,N_14968);
nand UO_94 (O_94,N_14824,N_14990);
nor UO_95 (O_95,N_14999,N_14994);
nand UO_96 (O_96,N_14830,N_14877);
xnor UO_97 (O_97,N_14991,N_14815);
or UO_98 (O_98,N_14851,N_14946);
and UO_99 (O_99,N_14932,N_14831);
nor UO_100 (O_100,N_14960,N_14994);
and UO_101 (O_101,N_14948,N_14931);
nor UO_102 (O_102,N_14893,N_14838);
and UO_103 (O_103,N_14843,N_14859);
and UO_104 (O_104,N_14959,N_14861);
nand UO_105 (O_105,N_14864,N_14924);
nor UO_106 (O_106,N_14987,N_14932);
nor UO_107 (O_107,N_14802,N_14950);
or UO_108 (O_108,N_14942,N_14971);
or UO_109 (O_109,N_14911,N_14936);
nor UO_110 (O_110,N_14900,N_14928);
and UO_111 (O_111,N_14988,N_14994);
xor UO_112 (O_112,N_14850,N_14977);
and UO_113 (O_113,N_14861,N_14911);
xnor UO_114 (O_114,N_14972,N_14818);
and UO_115 (O_115,N_14805,N_14929);
or UO_116 (O_116,N_14943,N_14970);
nand UO_117 (O_117,N_14844,N_14854);
nor UO_118 (O_118,N_14956,N_14815);
nand UO_119 (O_119,N_14979,N_14893);
or UO_120 (O_120,N_14895,N_14859);
xor UO_121 (O_121,N_14953,N_14928);
and UO_122 (O_122,N_14976,N_14951);
or UO_123 (O_123,N_14887,N_14925);
nand UO_124 (O_124,N_14977,N_14872);
nor UO_125 (O_125,N_14870,N_14820);
nor UO_126 (O_126,N_14870,N_14831);
or UO_127 (O_127,N_14905,N_14915);
nand UO_128 (O_128,N_14838,N_14890);
or UO_129 (O_129,N_14986,N_14952);
or UO_130 (O_130,N_14801,N_14963);
xnor UO_131 (O_131,N_14856,N_14844);
xnor UO_132 (O_132,N_14819,N_14885);
nor UO_133 (O_133,N_14831,N_14894);
and UO_134 (O_134,N_14891,N_14839);
nand UO_135 (O_135,N_14922,N_14806);
nor UO_136 (O_136,N_14976,N_14891);
or UO_137 (O_137,N_14805,N_14959);
and UO_138 (O_138,N_14838,N_14964);
nor UO_139 (O_139,N_14941,N_14857);
nor UO_140 (O_140,N_14846,N_14897);
nand UO_141 (O_141,N_14976,N_14850);
nand UO_142 (O_142,N_14988,N_14810);
and UO_143 (O_143,N_14868,N_14941);
and UO_144 (O_144,N_14857,N_14914);
and UO_145 (O_145,N_14904,N_14936);
xnor UO_146 (O_146,N_14892,N_14994);
and UO_147 (O_147,N_14819,N_14802);
xnor UO_148 (O_148,N_14969,N_14872);
or UO_149 (O_149,N_14965,N_14842);
nor UO_150 (O_150,N_14823,N_14906);
nor UO_151 (O_151,N_14979,N_14915);
and UO_152 (O_152,N_14907,N_14804);
xnor UO_153 (O_153,N_14944,N_14992);
xor UO_154 (O_154,N_14818,N_14898);
or UO_155 (O_155,N_14979,N_14957);
nor UO_156 (O_156,N_14857,N_14934);
and UO_157 (O_157,N_14854,N_14908);
and UO_158 (O_158,N_14907,N_14910);
xor UO_159 (O_159,N_14865,N_14884);
nand UO_160 (O_160,N_14939,N_14976);
or UO_161 (O_161,N_14960,N_14843);
nor UO_162 (O_162,N_14864,N_14907);
xor UO_163 (O_163,N_14867,N_14922);
or UO_164 (O_164,N_14977,N_14880);
nand UO_165 (O_165,N_14874,N_14937);
nor UO_166 (O_166,N_14905,N_14816);
xor UO_167 (O_167,N_14825,N_14869);
or UO_168 (O_168,N_14899,N_14895);
and UO_169 (O_169,N_14861,N_14845);
and UO_170 (O_170,N_14952,N_14825);
xor UO_171 (O_171,N_14934,N_14829);
and UO_172 (O_172,N_14808,N_14851);
nand UO_173 (O_173,N_14824,N_14883);
or UO_174 (O_174,N_14936,N_14802);
or UO_175 (O_175,N_14883,N_14880);
nand UO_176 (O_176,N_14952,N_14969);
nand UO_177 (O_177,N_14875,N_14876);
xor UO_178 (O_178,N_14807,N_14808);
nand UO_179 (O_179,N_14889,N_14953);
nand UO_180 (O_180,N_14890,N_14938);
and UO_181 (O_181,N_14852,N_14955);
nor UO_182 (O_182,N_14901,N_14940);
or UO_183 (O_183,N_14814,N_14824);
nand UO_184 (O_184,N_14965,N_14816);
or UO_185 (O_185,N_14976,N_14859);
or UO_186 (O_186,N_14891,N_14928);
or UO_187 (O_187,N_14822,N_14977);
xnor UO_188 (O_188,N_14964,N_14894);
or UO_189 (O_189,N_14945,N_14819);
or UO_190 (O_190,N_14919,N_14801);
xor UO_191 (O_191,N_14921,N_14912);
and UO_192 (O_192,N_14975,N_14945);
xor UO_193 (O_193,N_14892,N_14807);
or UO_194 (O_194,N_14838,N_14933);
or UO_195 (O_195,N_14968,N_14937);
and UO_196 (O_196,N_14899,N_14854);
nand UO_197 (O_197,N_14918,N_14898);
nand UO_198 (O_198,N_14985,N_14859);
nor UO_199 (O_199,N_14852,N_14831);
xnor UO_200 (O_200,N_14977,N_14938);
or UO_201 (O_201,N_14824,N_14982);
and UO_202 (O_202,N_14997,N_14839);
nand UO_203 (O_203,N_14981,N_14949);
and UO_204 (O_204,N_14988,N_14975);
and UO_205 (O_205,N_14961,N_14946);
nor UO_206 (O_206,N_14896,N_14946);
xnor UO_207 (O_207,N_14977,N_14884);
or UO_208 (O_208,N_14826,N_14932);
nor UO_209 (O_209,N_14895,N_14867);
nor UO_210 (O_210,N_14987,N_14822);
and UO_211 (O_211,N_14863,N_14922);
or UO_212 (O_212,N_14962,N_14809);
nor UO_213 (O_213,N_14974,N_14836);
nand UO_214 (O_214,N_14904,N_14810);
or UO_215 (O_215,N_14830,N_14839);
or UO_216 (O_216,N_14976,N_14827);
nand UO_217 (O_217,N_14883,N_14864);
xor UO_218 (O_218,N_14880,N_14830);
xnor UO_219 (O_219,N_14884,N_14992);
nor UO_220 (O_220,N_14959,N_14833);
and UO_221 (O_221,N_14878,N_14819);
or UO_222 (O_222,N_14818,N_14829);
nor UO_223 (O_223,N_14813,N_14907);
or UO_224 (O_224,N_14980,N_14866);
xor UO_225 (O_225,N_14960,N_14873);
and UO_226 (O_226,N_14928,N_14854);
nor UO_227 (O_227,N_14813,N_14996);
nor UO_228 (O_228,N_14988,N_14972);
and UO_229 (O_229,N_14879,N_14940);
and UO_230 (O_230,N_14917,N_14934);
and UO_231 (O_231,N_14841,N_14886);
or UO_232 (O_232,N_14861,N_14949);
and UO_233 (O_233,N_14866,N_14859);
nor UO_234 (O_234,N_14970,N_14827);
nor UO_235 (O_235,N_14960,N_14879);
nand UO_236 (O_236,N_14845,N_14888);
nand UO_237 (O_237,N_14817,N_14883);
or UO_238 (O_238,N_14913,N_14970);
nand UO_239 (O_239,N_14901,N_14984);
nor UO_240 (O_240,N_14814,N_14987);
xor UO_241 (O_241,N_14888,N_14995);
nand UO_242 (O_242,N_14898,N_14911);
nor UO_243 (O_243,N_14926,N_14947);
and UO_244 (O_244,N_14847,N_14948);
xnor UO_245 (O_245,N_14874,N_14936);
and UO_246 (O_246,N_14912,N_14896);
nor UO_247 (O_247,N_14841,N_14833);
xnor UO_248 (O_248,N_14925,N_14812);
or UO_249 (O_249,N_14973,N_14954);
or UO_250 (O_250,N_14982,N_14836);
nor UO_251 (O_251,N_14843,N_14803);
and UO_252 (O_252,N_14872,N_14902);
xnor UO_253 (O_253,N_14971,N_14801);
nand UO_254 (O_254,N_14869,N_14983);
xnor UO_255 (O_255,N_14919,N_14847);
nand UO_256 (O_256,N_14826,N_14896);
nor UO_257 (O_257,N_14903,N_14906);
and UO_258 (O_258,N_14831,N_14845);
or UO_259 (O_259,N_14847,N_14930);
nand UO_260 (O_260,N_14800,N_14822);
nor UO_261 (O_261,N_14916,N_14962);
xnor UO_262 (O_262,N_14963,N_14899);
nand UO_263 (O_263,N_14965,N_14982);
and UO_264 (O_264,N_14926,N_14988);
xor UO_265 (O_265,N_14848,N_14908);
or UO_266 (O_266,N_14906,N_14866);
nor UO_267 (O_267,N_14933,N_14939);
nor UO_268 (O_268,N_14917,N_14911);
and UO_269 (O_269,N_14920,N_14872);
nor UO_270 (O_270,N_14914,N_14836);
and UO_271 (O_271,N_14878,N_14920);
nand UO_272 (O_272,N_14896,N_14936);
nor UO_273 (O_273,N_14889,N_14981);
and UO_274 (O_274,N_14976,N_14849);
or UO_275 (O_275,N_14829,N_14990);
nand UO_276 (O_276,N_14987,N_14819);
or UO_277 (O_277,N_14984,N_14864);
and UO_278 (O_278,N_14879,N_14875);
or UO_279 (O_279,N_14838,N_14804);
or UO_280 (O_280,N_14870,N_14889);
nand UO_281 (O_281,N_14971,N_14923);
nand UO_282 (O_282,N_14908,N_14911);
or UO_283 (O_283,N_14812,N_14978);
nand UO_284 (O_284,N_14868,N_14892);
xnor UO_285 (O_285,N_14984,N_14950);
nor UO_286 (O_286,N_14972,N_14932);
nor UO_287 (O_287,N_14948,N_14897);
nor UO_288 (O_288,N_14920,N_14804);
nand UO_289 (O_289,N_14906,N_14807);
xor UO_290 (O_290,N_14971,N_14931);
or UO_291 (O_291,N_14914,N_14964);
nand UO_292 (O_292,N_14903,N_14874);
xor UO_293 (O_293,N_14963,N_14973);
xnor UO_294 (O_294,N_14957,N_14910);
nor UO_295 (O_295,N_14902,N_14942);
xor UO_296 (O_296,N_14871,N_14889);
xor UO_297 (O_297,N_14970,N_14972);
nand UO_298 (O_298,N_14943,N_14994);
xnor UO_299 (O_299,N_14920,N_14861);
nand UO_300 (O_300,N_14988,N_14997);
nor UO_301 (O_301,N_14951,N_14943);
nor UO_302 (O_302,N_14900,N_14967);
and UO_303 (O_303,N_14912,N_14975);
xnor UO_304 (O_304,N_14996,N_14960);
or UO_305 (O_305,N_14877,N_14940);
nand UO_306 (O_306,N_14897,N_14974);
nor UO_307 (O_307,N_14989,N_14907);
nor UO_308 (O_308,N_14904,N_14868);
and UO_309 (O_309,N_14946,N_14921);
or UO_310 (O_310,N_14830,N_14906);
xor UO_311 (O_311,N_14935,N_14832);
nand UO_312 (O_312,N_14996,N_14808);
xor UO_313 (O_313,N_14998,N_14850);
and UO_314 (O_314,N_14828,N_14947);
nor UO_315 (O_315,N_14938,N_14971);
nand UO_316 (O_316,N_14933,N_14809);
xnor UO_317 (O_317,N_14830,N_14923);
or UO_318 (O_318,N_14815,N_14931);
or UO_319 (O_319,N_14969,N_14997);
nor UO_320 (O_320,N_14800,N_14967);
and UO_321 (O_321,N_14995,N_14880);
nor UO_322 (O_322,N_14800,N_14979);
and UO_323 (O_323,N_14925,N_14813);
or UO_324 (O_324,N_14850,N_14848);
nand UO_325 (O_325,N_14924,N_14856);
nor UO_326 (O_326,N_14830,N_14868);
nand UO_327 (O_327,N_14974,N_14919);
or UO_328 (O_328,N_14907,N_14860);
and UO_329 (O_329,N_14872,N_14873);
nor UO_330 (O_330,N_14875,N_14818);
and UO_331 (O_331,N_14962,N_14903);
and UO_332 (O_332,N_14817,N_14937);
or UO_333 (O_333,N_14905,N_14995);
and UO_334 (O_334,N_14951,N_14964);
nor UO_335 (O_335,N_14841,N_14845);
or UO_336 (O_336,N_14814,N_14845);
nand UO_337 (O_337,N_14877,N_14927);
or UO_338 (O_338,N_14807,N_14913);
xor UO_339 (O_339,N_14849,N_14857);
nor UO_340 (O_340,N_14915,N_14832);
nand UO_341 (O_341,N_14887,N_14926);
nand UO_342 (O_342,N_14849,N_14869);
xor UO_343 (O_343,N_14824,N_14817);
xnor UO_344 (O_344,N_14822,N_14884);
or UO_345 (O_345,N_14914,N_14881);
nor UO_346 (O_346,N_14918,N_14903);
xor UO_347 (O_347,N_14899,N_14993);
nand UO_348 (O_348,N_14996,N_14878);
nand UO_349 (O_349,N_14924,N_14861);
nand UO_350 (O_350,N_14874,N_14879);
nor UO_351 (O_351,N_14822,N_14867);
xor UO_352 (O_352,N_14959,N_14857);
nor UO_353 (O_353,N_14898,N_14871);
or UO_354 (O_354,N_14837,N_14888);
or UO_355 (O_355,N_14890,N_14882);
nand UO_356 (O_356,N_14913,N_14810);
nor UO_357 (O_357,N_14830,N_14801);
nand UO_358 (O_358,N_14985,N_14894);
or UO_359 (O_359,N_14843,N_14883);
xor UO_360 (O_360,N_14858,N_14831);
nor UO_361 (O_361,N_14983,N_14803);
and UO_362 (O_362,N_14995,N_14967);
xnor UO_363 (O_363,N_14967,N_14987);
and UO_364 (O_364,N_14875,N_14922);
and UO_365 (O_365,N_14811,N_14956);
and UO_366 (O_366,N_14938,N_14986);
or UO_367 (O_367,N_14841,N_14924);
and UO_368 (O_368,N_14914,N_14838);
or UO_369 (O_369,N_14954,N_14827);
xor UO_370 (O_370,N_14862,N_14939);
nor UO_371 (O_371,N_14830,N_14903);
and UO_372 (O_372,N_14804,N_14911);
or UO_373 (O_373,N_14910,N_14888);
or UO_374 (O_374,N_14978,N_14926);
nand UO_375 (O_375,N_14955,N_14854);
nand UO_376 (O_376,N_14815,N_14838);
xnor UO_377 (O_377,N_14836,N_14906);
nor UO_378 (O_378,N_14848,N_14826);
and UO_379 (O_379,N_14821,N_14932);
xor UO_380 (O_380,N_14950,N_14909);
nand UO_381 (O_381,N_14841,N_14934);
and UO_382 (O_382,N_14914,N_14850);
xor UO_383 (O_383,N_14871,N_14838);
xnor UO_384 (O_384,N_14954,N_14824);
or UO_385 (O_385,N_14922,N_14872);
and UO_386 (O_386,N_14804,N_14876);
xnor UO_387 (O_387,N_14934,N_14996);
or UO_388 (O_388,N_14973,N_14906);
nand UO_389 (O_389,N_14866,N_14830);
xnor UO_390 (O_390,N_14996,N_14981);
or UO_391 (O_391,N_14940,N_14903);
and UO_392 (O_392,N_14922,N_14902);
xnor UO_393 (O_393,N_14812,N_14897);
and UO_394 (O_394,N_14957,N_14810);
nand UO_395 (O_395,N_14800,N_14846);
or UO_396 (O_396,N_14804,N_14973);
and UO_397 (O_397,N_14820,N_14854);
nand UO_398 (O_398,N_14803,N_14880);
or UO_399 (O_399,N_14827,N_14887);
nor UO_400 (O_400,N_14826,N_14801);
nor UO_401 (O_401,N_14935,N_14895);
and UO_402 (O_402,N_14838,N_14978);
or UO_403 (O_403,N_14978,N_14820);
xnor UO_404 (O_404,N_14807,N_14850);
nand UO_405 (O_405,N_14895,N_14904);
nor UO_406 (O_406,N_14818,N_14857);
and UO_407 (O_407,N_14986,N_14977);
nand UO_408 (O_408,N_14814,N_14990);
xnor UO_409 (O_409,N_14969,N_14908);
nor UO_410 (O_410,N_14826,N_14921);
nand UO_411 (O_411,N_14850,N_14939);
or UO_412 (O_412,N_14866,N_14805);
xor UO_413 (O_413,N_14856,N_14934);
and UO_414 (O_414,N_14911,N_14899);
nand UO_415 (O_415,N_14969,N_14994);
xor UO_416 (O_416,N_14812,N_14913);
or UO_417 (O_417,N_14807,N_14895);
or UO_418 (O_418,N_14920,N_14949);
nor UO_419 (O_419,N_14968,N_14973);
nand UO_420 (O_420,N_14837,N_14844);
and UO_421 (O_421,N_14878,N_14839);
nand UO_422 (O_422,N_14873,N_14824);
xnor UO_423 (O_423,N_14890,N_14831);
or UO_424 (O_424,N_14839,N_14874);
xor UO_425 (O_425,N_14942,N_14953);
xnor UO_426 (O_426,N_14981,N_14914);
nor UO_427 (O_427,N_14987,N_14883);
and UO_428 (O_428,N_14867,N_14933);
or UO_429 (O_429,N_14891,N_14990);
nand UO_430 (O_430,N_14922,N_14996);
or UO_431 (O_431,N_14840,N_14946);
and UO_432 (O_432,N_14931,N_14904);
or UO_433 (O_433,N_14822,N_14938);
nor UO_434 (O_434,N_14886,N_14962);
xnor UO_435 (O_435,N_14815,N_14970);
and UO_436 (O_436,N_14872,N_14845);
nand UO_437 (O_437,N_14822,N_14937);
nand UO_438 (O_438,N_14926,N_14976);
or UO_439 (O_439,N_14873,N_14981);
nor UO_440 (O_440,N_14951,N_14829);
nand UO_441 (O_441,N_14809,N_14852);
or UO_442 (O_442,N_14979,N_14918);
nor UO_443 (O_443,N_14985,N_14944);
nor UO_444 (O_444,N_14882,N_14908);
nand UO_445 (O_445,N_14979,N_14995);
or UO_446 (O_446,N_14970,N_14901);
and UO_447 (O_447,N_14950,N_14813);
nor UO_448 (O_448,N_14894,N_14995);
nor UO_449 (O_449,N_14912,N_14998);
nor UO_450 (O_450,N_14823,N_14848);
and UO_451 (O_451,N_14870,N_14818);
nand UO_452 (O_452,N_14976,N_14896);
nand UO_453 (O_453,N_14959,N_14915);
and UO_454 (O_454,N_14817,N_14831);
nand UO_455 (O_455,N_14907,N_14835);
nor UO_456 (O_456,N_14903,N_14859);
nor UO_457 (O_457,N_14983,N_14982);
nand UO_458 (O_458,N_14815,N_14813);
xor UO_459 (O_459,N_14886,N_14951);
or UO_460 (O_460,N_14861,N_14903);
nor UO_461 (O_461,N_14909,N_14817);
xor UO_462 (O_462,N_14823,N_14918);
xor UO_463 (O_463,N_14830,N_14803);
xor UO_464 (O_464,N_14943,N_14844);
nand UO_465 (O_465,N_14826,N_14821);
and UO_466 (O_466,N_14987,N_14805);
xnor UO_467 (O_467,N_14830,N_14919);
xor UO_468 (O_468,N_14827,N_14946);
or UO_469 (O_469,N_14863,N_14884);
xor UO_470 (O_470,N_14811,N_14962);
nor UO_471 (O_471,N_14898,N_14844);
and UO_472 (O_472,N_14870,N_14968);
or UO_473 (O_473,N_14828,N_14900);
xnor UO_474 (O_474,N_14814,N_14879);
nor UO_475 (O_475,N_14979,N_14884);
and UO_476 (O_476,N_14932,N_14906);
nand UO_477 (O_477,N_14984,N_14811);
xnor UO_478 (O_478,N_14928,N_14905);
nand UO_479 (O_479,N_14876,N_14811);
nand UO_480 (O_480,N_14995,N_14949);
xor UO_481 (O_481,N_14843,N_14963);
and UO_482 (O_482,N_14849,N_14956);
and UO_483 (O_483,N_14992,N_14836);
or UO_484 (O_484,N_14842,N_14927);
xnor UO_485 (O_485,N_14842,N_14879);
nand UO_486 (O_486,N_14982,N_14977);
or UO_487 (O_487,N_14804,N_14959);
or UO_488 (O_488,N_14911,N_14968);
xor UO_489 (O_489,N_14880,N_14822);
and UO_490 (O_490,N_14956,N_14889);
nor UO_491 (O_491,N_14972,N_14838);
xor UO_492 (O_492,N_14984,N_14870);
or UO_493 (O_493,N_14874,N_14848);
and UO_494 (O_494,N_14979,N_14987);
xor UO_495 (O_495,N_14812,N_14837);
or UO_496 (O_496,N_14849,N_14837);
nor UO_497 (O_497,N_14830,N_14905);
nor UO_498 (O_498,N_14828,N_14990);
and UO_499 (O_499,N_14899,N_14977);
or UO_500 (O_500,N_14935,N_14892);
nand UO_501 (O_501,N_14890,N_14957);
nand UO_502 (O_502,N_14850,N_14875);
nand UO_503 (O_503,N_14935,N_14851);
nand UO_504 (O_504,N_14973,N_14809);
nor UO_505 (O_505,N_14949,N_14834);
and UO_506 (O_506,N_14896,N_14908);
nor UO_507 (O_507,N_14921,N_14894);
nor UO_508 (O_508,N_14958,N_14935);
nor UO_509 (O_509,N_14800,N_14924);
xnor UO_510 (O_510,N_14869,N_14932);
xnor UO_511 (O_511,N_14890,N_14917);
nor UO_512 (O_512,N_14828,N_14814);
nand UO_513 (O_513,N_14828,N_14916);
and UO_514 (O_514,N_14823,N_14812);
xor UO_515 (O_515,N_14844,N_14813);
nand UO_516 (O_516,N_14916,N_14952);
or UO_517 (O_517,N_14948,N_14899);
nor UO_518 (O_518,N_14848,N_14840);
and UO_519 (O_519,N_14978,N_14805);
or UO_520 (O_520,N_14978,N_14879);
nand UO_521 (O_521,N_14853,N_14993);
xnor UO_522 (O_522,N_14964,N_14908);
nand UO_523 (O_523,N_14857,N_14837);
nor UO_524 (O_524,N_14904,N_14942);
nand UO_525 (O_525,N_14812,N_14932);
xnor UO_526 (O_526,N_14947,N_14849);
nand UO_527 (O_527,N_14915,N_14864);
nand UO_528 (O_528,N_14997,N_14907);
nor UO_529 (O_529,N_14970,N_14979);
xnor UO_530 (O_530,N_14806,N_14887);
nand UO_531 (O_531,N_14864,N_14801);
xnor UO_532 (O_532,N_14896,N_14820);
nand UO_533 (O_533,N_14936,N_14879);
and UO_534 (O_534,N_14920,N_14930);
nand UO_535 (O_535,N_14997,N_14950);
and UO_536 (O_536,N_14813,N_14854);
or UO_537 (O_537,N_14843,N_14869);
and UO_538 (O_538,N_14881,N_14917);
xnor UO_539 (O_539,N_14827,N_14847);
and UO_540 (O_540,N_14999,N_14968);
or UO_541 (O_541,N_14989,N_14884);
and UO_542 (O_542,N_14849,N_14886);
and UO_543 (O_543,N_14947,N_14984);
xor UO_544 (O_544,N_14814,N_14907);
and UO_545 (O_545,N_14926,N_14800);
and UO_546 (O_546,N_14840,N_14805);
nand UO_547 (O_547,N_14960,N_14804);
nor UO_548 (O_548,N_14959,N_14922);
nand UO_549 (O_549,N_14890,N_14979);
xnor UO_550 (O_550,N_14839,N_14981);
nor UO_551 (O_551,N_14978,N_14950);
or UO_552 (O_552,N_14989,N_14891);
and UO_553 (O_553,N_14844,N_14803);
or UO_554 (O_554,N_14813,N_14809);
nand UO_555 (O_555,N_14908,N_14819);
nand UO_556 (O_556,N_14957,N_14842);
or UO_557 (O_557,N_14937,N_14867);
nor UO_558 (O_558,N_14961,N_14996);
xor UO_559 (O_559,N_14814,N_14922);
and UO_560 (O_560,N_14968,N_14833);
and UO_561 (O_561,N_14856,N_14896);
or UO_562 (O_562,N_14850,N_14852);
nand UO_563 (O_563,N_14999,N_14901);
or UO_564 (O_564,N_14842,N_14952);
xnor UO_565 (O_565,N_14862,N_14856);
nor UO_566 (O_566,N_14871,N_14878);
nor UO_567 (O_567,N_14900,N_14971);
nand UO_568 (O_568,N_14851,N_14845);
or UO_569 (O_569,N_14952,N_14857);
and UO_570 (O_570,N_14945,N_14909);
nor UO_571 (O_571,N_14884,N_14839);
xor UO_572 (O_572,N_14990,N_14924);
nor UO_573 (O_573,N_14857,N_14807);
or UO_574 (O_574,N_14993,N_14891);
nor UO_575 (O_575,N_14818,N_14891);
and UO_576 (O_576,N_14999,N_14890);
or UO_577 (O_577,N_14843,N_14985);
and UO_578 (O_578,N_14971,N_14819);
xor UO_579 (O_579,N_14896,N_14840);
xor UO_580 (O_580,N_14844,N_14847);
nor UO_581 (O_581,N_14841,N_14868);
or UO_582 (O_582,N_14846,N_14970);
or UO_583 (O_583,N_14921,N_14976);
and UO_584 (O_584,N_14912,N_14990);
nand UO_585 (O_585,N_14832,N_14919);
xnor UO_586 (O_586,N_14945,N_14967);
and UO_587 (O_587,N_14843,N_14874);
xnor UO_588 (O_588,N_14843,N_14839);
or UO_589 (O_589,N_14852,N_14913);
and UO_590 (O_590,N_14998,N_14949);
nor UO_591 (O_591,N_14823,N_14972);
and UO_592 (O_592,N_14833,N_14830);
and UO_593 (O_593,N_14903,N_14845);
and UO_594 (O_594,N_14974,N_14931);
nand UO_595 (O_595,N_14805,N_14975);
nand UO_596 (O_596,N_14928,N_14922);
nor UO_597 (O_597,N_14966,N_14950);
nand UO_598 (O_598,N_14948,N_14988);
or UO_599 (O_599,N_14980,N_14931);
nand UO_600 (O_600,N_14846,N_14992);
xor UO_601 (O_601,N_14845,N_14895);
xnor UO_602 (O_602,N_14866,N_14880);
and UO_603 (O_603,N_14889,N_14942);
xor UO_604 (O_604,N_14879,N_14839);
and UO_605 (O_605,N_14821,N_14860);
nand UO_606 (O_606,N_14963,N_14811);
and UO_607 (O_607,N_14875,N_14885);
xor UO_608 (O_608,N_14967,N_14948);
nor UO_609 (O_609,N_14838,N_14984);
xor UO_610 (O_610,N_14866,N_14911);
nor UO_611 (O_611,N_14877,N_14829);
nor UO_612 (O_612,N_14864,N_14836);
xor UO_613 (O_613,N_14893,N_14847);
nor UO_614 (O_614,N_14954,N_14933);
nand UO_615 (O_615,N_14937,N_14991);
xnor UO_616 (O_616,N_14912,N_14954);
and UO_617 (O_617,N_14828,N_14942);
or UO_618 (O_618,N_14905,N_14874);
nor UO_619 (O_619,N_14939,N_14815);
and UO_620 (O_620,N_14904,N_14804);
xnor UO_621 (O_621,N_14913,N_14961);
nor UO_622 (O_622,N_14861,N_14973);
and UO_623 (O_623,N_14939,N_14810);
nand UO_624 (O_624,N_14929,N_14931);
and UO_625 (O_625,N_14872,N_14865);
nand UO_626 (O_626,N_14848,N_14967);
xor UO_627 (O_627,N_14836,N_14858);
nand UO_628 (O_628,N_14850,N_14973);
or UO_629 (O_629,N_14908,N_14974);
xnor UO_630 (O_630,N_14813,N_14994);
nand UO_631 (O_631,N_14805,N_14816);
nand UO_632 (O_632,N_14894,N_14878);
or UO_633 (O_633,N_14819,N_14960);
and UO_634 (O_634,N_14929,N_14867);
xor UO_635 (O_635,N_14915,N_14865);
nor UO_636 (O_636,N_14899,N_14966);
or UO_637 (O_637,N_14964,N_14830);
nand UO_638 (O_638,N_14962,N_14968);
xnor UO_639 (O_639,N_14882,N_14959);
and UO_640 (O_640,N_14865,N_14985);
xor UO_641 (O_641,N_14946,N_14854);
or UO_642 (O_642,N_14883,N_14926);
and UO_643 (O_643,N_14961,N_14865);
and UO_644 (O_644,N_14834,N_14945);
nor UO_645 (O_645,N_14842,N_14986);
xnor UO_646 (O_646,N_14974,N_14989);
nor UO_647 (O_647,N_14927,N_14838);
and UO_648 (O_648,N_14809,N_14896);
or UO_649 (O_649,N_14939,N_14981);
xor UO_650 (O_650,N_14945,N_14801);
nor UO_651 (O_651,N_14910,N_14905);
or UO_652 (O_652,N_14832,N_14999);
or UO_653 (O_653,N_14910,N_14840);
nand UO_654 (O_654,N_14960,N_14898);
nand UO_655 (O_655,N_14893,N_14868);
and UO_656 (O_656,N_14890,N_14857);
nand UO_657 (O_657,N_14964,N_14895);
nand UO_658 (O_658,N_14895,N_14958);
nor UO_659 (O_659,N_14863,N_14833);
and UO_660 (O_660,N_14919,N_14961);
and UO_661 (O_661,N_14863,N_14844);
xnor UO_662 (O_662,N_14903,N_14846);
nor UO_663 (O_663,N_14960,N_14941);
and UO_664 (O_664,N_14931,N_14939);
nor UO_665 (O_665,N_14838,N_14861);
nor UO_666 (O_666,N_14869,N_14961);
nor UO_667 (O_667,N_14933,N_14889);
or UO_668 (O_668,N_14869,N_14809);
or UO_669 (O_669,N_14842,N_14951);
nor UO_670 (O_670,N_14902,N_14938);
nor UO_671 (O_671,N_14963,N_14887);
or UO_672 (O_672,N_14801,N_14827);
nor UO_673 (O_673,N_14999,N_14872);
or UO_674 (O_674,N_14888,N_14911);
nand UO_675 (O_675,N_14935,N_14894);
xor UO_676 (O_676,N_14865,N_14814);
nand UO_677 (O_677,N_14884,N_14981);
nand UO_678 (O_678,N_14880,N_14818);
xor UO_679 (O_679,N_14960,N_14862);
or UO_680 (O_680,N_14987,N_14974);
and UO_681 (O_681,N_14814,N_14943);
xor UO_682 (O_682,N_14905,N_14867);
and UO_683 (O_683,N_14934,N_14992);
and UO_684 (O_684,N_14941,N_14970);
xor UO_685 (O_685,N_14950,N_14960);
nand UO_686 (O_686,N_14910,N_14838);
and UO_687 (O_687,N_14901,N_14986);
and UO_688 (O_688,N_14973,N_14880);
nor UO_689 (O_689,N_14842,N_14935);
and UO_690 (O_690,N_14871,N_14943);
and UO_691 (O_691,N_14869,N_14900);
nand UO_692 (O_692,N_14917,N_14965);
and UO_693 (O_693,N_14974,N_14992);
and UO_694 (O_694,N_14903,N_14969);
and UO_695 (O_695,N_14889,N_14911);
or UO_696 (O_696,N_14852,N_14875);
xor UO_697 (O_697,N_14954,N_14889);
and UO_698 (O_698,N_14963,N_14802);
nor UO_699 (O_699,N_14860,N_14829);
nand UO_700 (O_700,N_14964,N_14952);
or UO_701 (O_701,N_14964,N_14875);
and UO_702 (O_702,N_14863,N_14993);
or UO_703 (O_703,N_14948,N_14952);
nor UO_704 (O_704,N_14954,N_14994);
xor UO_705 (O_705,N_14856,N_14946);
xnor UO_706 (O_706,N_14909,N_14861);
and UO_707 (O_707,N_14857,N_14933);
or UO_708 (O_708,N_14964,N_14911);
and UO_709 (O_709,N_14915,N_14909);
nand UO_710 (O_710,N_14949,N_14853);
xnor UO_711 (O_711,N_14951,N_14862);
xnor UO_712 (O_712,N_14979,N_14828);
or UO_713 (O_713,N_14931,N_14874);
nand UO_714 (O_714,N_14876,N_14908);
or UO_715 (O_715,N_14893,N_14818);
nor UO_716 (O_716,N_14804,N_14984);
or UO_717 (O_717,N_14941,N_14887);
or UO_718 (O_718,N_14927,N_14912);
and UO_719 (O_719,N_14802,N_14909);
nor UO_720 (O_720,N_14904,N_14934);
or UO_721 (O_721,N_14914,N_14933);
and UO_722 (O_722,N_14907,N_14912);
xnor UO_723 (O_723,N_14903,N_14892);
nor UO_724 (O_724,N_14877,N_14957);
nor UO_725 (O_725,N_14899,N_14828);
and UO_726 (O_726,N_14814,N_14887);
xor UO_727 (O_727,N_14964,N_14831);
nor UO_728 (O_728,N_14932,N_14960);
or UO_729 (O_729,N_14874,N_14944);
nor UO_730 (O_730,N_14810,N_14809);
or UO_731 (O_731,N_14934,N_14982);
xnor UO_732 (O_732,N_14800,N_14920);
and UO_733 (O_733,N_14806,N_14937);
nand UO_734 (O_734,N_14807,N_14854);
or UO_735 (O_735,N_14984,N_14921);
xor UO_736 (O_736,N_14966,N_14973);
or UO_737 (O_737,N_14991,N_14996);
and UO_738 (O_738,N_14870,N_14962);
or UO_739 (O_739,N_14842,N_14898);
and UO_740 (O_740,N_14965,N_14814);
xor UO_741 (O_741,N_14810,N_14952);
nand UO_742 (O_742,N_14973,N_14812);
and UO_743 (O_743,N_14888,N_14913);
nand UO_744 (O_744,N_14887,N_14971);
xnor UO_745 (O_745,N_14873,N_14837);
or UO_746 (O_746,N_14972,N_14975);
nand UO_747 (O_747,N_14944,N_14857);
or UO_748 (O_748,N_14994,N_14913);
and UO_749 (O_749,N_14909,N_14948);
nand UO_750 (O_750,N_14954,N_14960);
nor UO_751 (O_751,N_14931,N_14803);
nor UO_752 (O_752,N_14877,N_14922);
nor UO_753 (O_753,N_14892,N_14942);
nor UO_754 (O_754,N_14886,N_14972);
or UO_755 (O_755,N_14895,N_14866);
or UO_756 (O_756,N_14813,N_14910);
nor UO_757 (O_757,N_14916,N_14978);
and UO_758 (O_758,N_14932,N_14895);
nand UO_759 (O_759,N_14983,N_14847);
xnor UO_760 (O_760,N_14867,N_14967);
xnor UO_761 (O_761,N_14867,N_14847);
nand UO_762 (O_762,N_14891,N_14851);
and UO_763 (O_763,N_14847,N_14965);
and UO_764 (O_764,N_14968,N_14861);
xnor UO_765 (O_765,N_14905,N_14861);
nand UO_766 (O_766,N_14813,N_14906);
and UO_767 (O_767,N_14824,N_14827);
xnor UO_768 (O_768,N_14892,N_14836);
and UO_769 (O_769,N_14881,N_14869);
or UO_770 (O_770,N_14941,N_14993);
nand UO_771 (O_771,N_14837,N_14806);
xor UO_772 (O_772,N_14880,N_14896);
nor UO_773 (O_773,N_14808,N_14802);
or UO_774 (O_774,N_14995,N_14957);
nand UO_775 (O_775,N_14800,N_14813);
or UO_776 (O_776,N_14862,N_14883);
nand UO_777 (O_777,N_14966,N_14853);
or UO_778 (O_778,N_14894,N_14930);
or UO_779 (O_779,N_14959,N_14835);
xor UO_780 (O_780,N_14844,N_14855);
nor UO_781 (O_781,N_14952,N_14906);
nor UO_782 (O_782,N_14927,N_14907);
nand UO_783 (O_783,N_14883,N_14831);
xor UO_784 (O_784,N_14813,N_14857);
xnor UO_785 (O_785,N_14826,N_14907);
nand UO_786 (O_786,N_14974,N_14876);
nor UO_787 (O_787,N_14916,N_14959);
xnor UO_788 (O_788,N_14925,N_14917);
xor UO_789 (O_789,N_14890,N_14928);
xnor UO_790 (O_790,N_14826,N_14995);
nor UO_791 (O_791,N_14959,N_14809);
nor UO_792 (O_792,N_14872,N_14810);
or UO_793 (O_793,N_14894,N_14994);
xnor UO_794 (O_794,N_14843,N_14903);
and UO_795 (O_795,N_14962,N_14872);
and UO_796 (O_796,N_14849,N_14883);
nand UO_797 (O_797,N_14835,N_14986);
or UO_798 (O_798,N_14837,N_14861);
nor UO_799 (O_799,N_14929,N_14812);
nor UO_800 (O_800,N_14968,N_14872);
or UO_801 (O_801,N_14875,N_14934);
xnor UO_802 (O_802,N_14984,N_14988);
or UO_803 (O_803,N_14917,N_14853);
nor UO_804 (O_804,N_14845,N_14965);
or UO_805 (O_805,N_14950,N_14943);
and UO_806 (O_806,N_14879,N_14979);
and UO_807 (O_807,N_14919,N_14837);
nand UO_808 (O_808,N_14952,N_14937);
nand UO_809 (O_809,N_14829,N_14969);
xor UO_810 (O_810,N_14932,N_14928);
and UO_811 (O_811,N_14845,N_14983);
xnor UO_812 (O_812,N_14805,N_14940);
nand UO_813 (O_813,N_14893,N_14973);
nand UO_814 (O_814,N_14892,N_14933);
nand UO_815 (O_815,N_14963,N_14828);
and UO_816 (O_816,N_14908,N_14956);
or UO_817 (O_817,N_14989,N_14841);
nor UO_818 (O_818,N_14806,N_14824);
nand UO_819 (O_819,N_14801,N_14901);
or UO_820 (O_820,N_14965,N_14835);
xnor UO_821 (O_821,N_14868,N_14943);
or UO_822 (O_822,N_14894,N_14857);
xor UO_823 (O_823,N_14837,N_14938);
nand UO_824 (O_824,N_14828,N_14832);
xor UO_825 (O_825,N_14968,N_14913);
nand UO_826 (O_826,N_14995,N_14922);
xor UO_827 (O_827,N_14883,N_14873);
or UO_828 (O_828,N_14802,N_14823);
nand UO_829 (O_829,N_14914,N_14934);
nor UO_830 (O_830,N_14984,N_14999);
nor UO_831 (O_831,N_14880,N_14949);
xnor UO_832 (O_832,N_14957,N_14930);
and UO_833 (O_833,N_14979,N_14932);
nor UO_834 (O_834,N_14807,N_14860);
nand UO_835 (O_835,N_14946,N_14990);
or UO_836 (O_836,N_14950,N_14857);
nor UO_837 (O_837,N_14818,N_14825);
nand UO_838 (O_838,N_14851,N_14860);
or UO_839 (O_839,N_14943,N_14815);
nand UO_840 (O_840,N_14844,N_14816);
xnor UO_841 (O_841,N_14813,N_14990);
nand UO_842 (O_842,N_14898,N_14919);
xnor UO_843 (O_843,N_14977,N_14925);
or UO_844 (O_844,N_14892,N_14872);
and UO_845 (O_845,N_14917,N_14828);
xnor UO_846 (O_846,N_14996,N_14939);
nand UO_847 (O_847,N_14832,N_14888);
and UO_848 (O_848,N_14949,N_14801);
xnor UO_849 (O_849,N_14937,N_14953);
xor UO_850 (O_850,N_14990,N_14801);
nor UO_851 (O_851,N_14913,N_14925);
xnor UO_852 (O_852,N_14923,N_14863);
or UO_853 (O_853,N_14811,N_14883);
nor UO_854 (O_854,N_14866,N_14901);
xor UO_855 (O_855,N_14844,N_14949);
and UO_856 (O_856,N_14891,N_14881);
xnor UO_857 (O_857,N_14880,N_14936);
and UO_858 (O_858,N_14951,N_14848);
or UO_859 (O_859,N_14878,N_14950);
and UO_860 (O_860,N_14951,N_14885);
nand UO_861 (O_861,N_14952,N_14987);
xor UO_862 (O_862,N_14949,N_14814);
nor UO_863 (O_863,N_14881,N_14832);
or UO_864 (O_864,N_14873,N_14907);
and UO_865 (O_865,N_14937,N_14951);
nor UO_866 (O_866,N_14821,N_14851);
or UO_867 (O_867,N_14920,N_14884);
xor UO_868 (O_868,N_14932,N_14943);
xor UO_869 (O_869,N_14908,N_14803);
or UO_870 (O_870,N_14972,N_14937);
and UO_871 (O_871,N_14817,N_14880);
and UO_872 (O_872,N_14824,N_14907);
nand UO_873 (O_873,N_14899,N_14909);
and UO_874 (O_874,N_14981,N_14941);
and UO_875 (O_875,N_14888,N_14915);
xor UO_876 (O_876,N_14860,N_14827);
nand UO_877 (O_877,N_14871,N_14905);
and UO_878 (O_878,N_14823,N_14819);
nor UO_879 (O_879,N_14837,N_14900);
nand UO_880 (O_880,N_14987,N_14829);
nor UO_881 (O_881,N_14942,N_14931);
nand UO_882 (O_882,N_14919,N_14930);
nor UO_883 (O_883,N_14962,N_14964);
or UO_884 (O_884,N_14923,N_14912);
xnor UO_885 (O_885,N_14849,N_14894);
xor UO_886 (O_886,N_14960,N_14871);
and UO_887 (O_887,N_14932,N_14982);
or UO_888 (O_888,N_14951,N_14866);
nand UO_889 (O_889,N_14895,N_14898);
nand UO_890 (O_890,N_14844,N_14916);
xnor UO_891 (O_891,N_14896,N_14853);
nor UO_892 (O_892,N_14856,N_14836);
or UO_893 (O_893,N_14850,N_14927);
or UO_894 (O_894,N_14861,N_14841);
xor UO_895 (O_895,N_14950,N_14889);
nor UO_896 (O_896,N_14838,N_14943);
or UO_897 (O_897,N_14979,N_14994);
and UO_898 (O_898,N_14965,N_14808);
and UO_899 (O_899,N_14926,N_14985);
or UO_900 (O_900,N_14842,N_14968);
nor UO_901 (O_901,N_14909,N_14800);
nor UO_902 (O_902,N_14986,N_14863);
or UO_903 (O_903,N_14981,N_14845);
nor UO_904 (O_904,N_14833,N_14847);
nand UO_905 (O_905,N_14977,N_14836);
nand UO_906 (O_906,N_14993,N_14918);
or UO_907 (O_907,N_14976,N_14958);
and UO_908 (O_908,N_14879,N_14896);
nand UO_909 (O_909,N_14914,N_14811);
xor UO_910 (O_910,N_14838,N_14982);
or UO_911 (O_911,N_14970,N_14849);
or UO_912 (O_912,N_14943,N_14909);
and UO_913 (O_913,N_14902,N_14891);
nand UO_914 (O_914,N_14944,N_14870);
or UO_915 (O_915,N_14904,N_14979);
or UO_916 (O_916,N_14998,N_14963);
nand UO_917 (O_917,N_14924,N_14957);
and UO_918 (O_918,N_14939,N_14924);
xnor UO_919 (O_919,N_14837,N_14815);
or UO_920 (O_920,N_14861,N_14875);
and UO_921 (O_921,N_14833,N_14999);
or UO_922 (O_922,N_14908,N_14808);
or UO_923 (O_923,N_14896,N_14982);
xnor UO_924 (O_924,N_14915,N_14951);
or UO_925 (O_925,N_14806,N_14879);
xnor UO_926 (O_926,N_14880,N_14863);
nor UO_927 (O_927,N_14963,N_14842);
nor UO_928 (O_928,N_14954,N_14831);
or UO_929 (O_929,N_14838,N_14903);
nor UO_930 (O_930,N_14839,N_14873);
nor UO_931 (O_931,N_14948,N_14956);
or UO_932 (O_932,N_14897,N_14873);
nor UO_933 (O_933,N_14936,N_14985);
nor UO_934 (O_934,N_14991,N_14874);
or UO_935 (O_935,N_14835,N_14852);
or UO_936 (O_936,N_14949,N_14944);
nand UO_937 (O_937,N_14932,N_14996);
nor UO_938 (O_938,N_14835,N_14952);
nand UO_939 (O_939,N_14934,N_14861);
and UO_940 (O_940,N_14965,N_14923);
and UO_941 (O_941,N_14826,N_14941);
and UO_942 (O_942,N_14864,N_14872);
and UO_943 (O_943,N_14855,N_14957);
or UO_944 (O_944,N_14803,N_14938);
nand UO_945 (O_945,N_14882,N_14861);
nor UO_946 (O_946,N_14922,N_14982);
nor UO_947 (O_947,N_14930,N_14892);
nand UO_948 (O_948,N_14976,N_14819);
xor UO_949 (O_949,N_14815,N_14872);
or UO_950 (O_950,N_14900,N_14858);
nand UO_951 (O_951,N_14829,N_14816);
xnor UO_952 (O_952,N_14941,N_14923);
or UO_953 (O_953,N_14906,N_14979);
or UO_954 (O_954,N_14866,N_14966);
nor UO_955 (O_955,N_14966,N_14895);
nor UO_956 (O_956,N_14941,N_14838);
and UO_957 (O_957,N_14973,N_14837);
nand UO_958 (O_958,N_14874,N_14886);
xnor UO_959 (O_959,N_14926,N_14879);
and UO_960 (O_960,N_14941,N_14871);
or UO_961 (O_961,N_14947,N_14862);
and UO_962 (O_962,N_14998,N_14875);
nor UO_963 (O_963,N_14893,N_14934);
xor UO_964 (O_964,N_14911,N_14923);
xnor UO_965 (O_965,N_14921,N_14804);
nand UO_966 (O_966,N_14901,N_14961);
nor UO_967 (O_967,N_14878,N_14955);
nor UO_968 (O_968,N_14968,N_14955);
xnor UO_969 (O_969,N_14997,N_14825);
or UO_970 (O_970,N_14853,N_14841);
nor UO_971 (O_971,N_14935,N_14924);
nand UO_972 (O_972,N_14832,N_14990);
nor UO_973 (O_973,N_14955,N_14979);
nor UO_974 (O_974,N_14883,N_14891);
xnor UO_975 (O_975,N_14999,N_14870);
nor UO_976 (O_976,N_14866,N_14997);
nand UO_977 (O_977,N_14931,N_14849);
or UO_978 (O_978,N_14835,N_14803);
and UO_979 (O_979,N_14967,N_14927);
nor UO_980 (O_980,N_14852,N_14810);
nand UO_981 (O_981,N_14859,N_14956);
or UO_982 (O_982,N_14919,N_14869);
nand UO_983 (O_983,N_14830,N_14958);
and UO_984 (O_984,N_14804,N_14974);
nor UO_985 (O_985,N_14938,N_14974);
nand UO_986 (O_986,N_14868,N_14847);
nor UO_987 (O_987,N_14906,N_14847);
or UO_988 (O_988,N_14888,N_14841);
nor UO_989 (O_989,N_14939,N_14954);
or UO_990 (O_990,N_14981,N_14842);
or UO_991 (O_991,N_14912,N_14894);
or UO_992 (O_992,N_14888,N_14881);
nand UO_993 (O_993,N_14953,N_14927);
nand UO_994 (O_994,N_14898,N_14902);
nor UO_995 (O_995,N_14926,N_14892);
or UO_996 (O_996,N_14949,N_14922);
or UO_997 (O_997,N_14853,N_14843);
and UO_998 (O_998,N_14958,N_14960);
or UO_999 (O_999,N_14847,N_14939);
nor UO_1000 (O_1000,N_14903,N_14932);
or UO_1001 (O_1001,N_14938,N_14806);
xor UO_1002 (O_1002,N_14928,N_14959);
or UO_1003 (O_1003,N_14992,N_14941);
nand UO_1004 (O_1004,N_14983,N_14829);
and UO_1005 (O_1005,N_14983,N_14850);
nor UO_1006 (O_1006,N_14961,N_14856);
or UO_1007 (O_1007,N_14810,N_14847);
or UO_1008 (O_1008,N_14842,N_14860);
xnor UO_1009 (O_1009,N_14924,N_14871);
nor UO_1010 (O_1010,N_14868,N_14971);
nor UO_1011 (O_1011,N_14833,N_14878);
xnor UO_1012 (O_1012,N_14906,N_14890);
nand UO_1013 (O_1013,N_14972,N_14997);
nand UO_1014 (O_1014,N_14985,N_14895);
and UO_1015 (O_1015,N_14920,N_14900);
or UO_1016 (O_1016,N_14986,N_14838);
or UO_1017 (O_1017,N_14885,N_14931);
or UO_1018 (O_1018,N_14859,N_14966);
xnor UO_1019 (O_1019,N_14817,N_14985);
or UO_1020 (O_1020,N_14998,N_14956);
xnor UO_1021 (O_1021,N_14821,N_14841);
nor UO_1022 (O_1022,N_14980,N_14844);
xor UO_1023 (O_1023,N_14917,N_14998);
and UO_1024 (O_1024,N_14937,N_14882);
nand UO_1025 (O_1025,N_14877,N_14812);
xor UO_1026 (O_1026,N_14960,N_14852);
nor UO_1027 (O_1027,N_14925,N_14996);
nand UO_1028 (O_1028,N_14863,N_14985);
nand UO_1029 (O_1029,N_14981,N_14980);
nand UO_1030 (O_1030,N_14988,N_14946);
or UO_1031 (O_1031,N_14987,N_14898);
or UO_1032 (O_1032,N_14931,N_14958);
nand UO_1033 (O_1033,N_14906,N_14883);
nand UO_1034 (O_1034,N_14846,N_14980);
or UO_1035 (O_1035,N_14957,N_14999);
or UO_1036 (O_1036,N_14933,N_14982);
nor UO_1037 (O_1037,N_14879,N_14927);
nand UO_1038 (O_1038,N_14809,N_14929);
nand UO_1039 (O_1039,N_14941,N_14852);
nor UO_1040 (O_1040,N_14864,N_14921);
nor UO_1041 (O_1041,N_14951,N_14807);
nand UO_1042 (O_1042,N_14931,N_14878);
or UO_1043 (O_1043,N_14941,N_14905);
nand UO_1044 (O_1044,N_14935,N_14850);
xor UO_1045 (O_1045,N_14998,N_14948);
or UO_1046 (O_1046,N_14947,N_14939);
or UO_1047 (O_1047,N_14879,N_14845);
nand UO_1048 (O_1048,N_14961,N_14986);
nand UO_1049 (O_1049,N_14801,N_14819);
or UO_1050 (O_1050,N_14937,N_14985);
nor UO_1051 (O_1051,N_14837,N_14817);
or UO_1052 (O_1052,N_14986,N_14820);
nor UO_1053 (O_1053,N_14902,N_14977);
nand UO_1054 (O_1054,N_14813,N_14802);
xnor UO_1055 (O_1055,N_14866,N_14996);
or UO_1056 (O_1056,N_14910,N_14997);
or UO_1057 (O_1057,N_14907,N_14806);
or UO_1058 (O_1058,N_14916,N_14862);
nand UO_1059 (O_1059,N_14897,N_14898);
nand UO_1060 (O_1060,N_14858,N_14968);
xnor UO_1061 (O_1061,N_14822,N_14962);
xor UO_1062 (O_1062,N_14900,N_14863);
xor UO_1063 (O_1063,N_14828,N_14978);
nor UO_1064 (O_1064,N_14922,N_14965);
nor UO_1065 (O_1065,N_14859,N_14831);
nor UO_1066 (O_1066,N_14868,N_14831);
nor UO_1067 (O_1067,N_14888,N_14981);
nand UO_1068 (O_1068,N_14962,N_14925);
or UO_1069 (O_1069,N_14907,N_14933);
or UO_1070 (O_1070,N_14987,N_14917);
xor UO_1071 (O_1071,N_14845,N_14890);
or UO_1072 (O_1072,N_14868,N_14806);
or UO_1073 (O_1073,N_14892,N_14838);
and UO_1074 (O_1074,N_14812,N_14910);
nor UO_1075 (O_1075,N_14909,N_14905);
and UO_1076 (O_1076,N_14967,N_14956);
nand UO_1077 (O_1077,N_14936,N_14947);
nor UO_1078 (O_1078,N_14810,N_14946);
xnor UO_1079 (O_1079,N_14973,N_14962);
nor UO_1080 (O_1080,N_14977,N_14921);
xor UO_1081 (O_1081,N_14988,N_14938);
nand UO_1082 (O_1082,N_14939,N_14987);
nor UO_1083 (O_1083,N_14842,N_14967);
or UO_1084 (O_1084,N_14946,N_14958);
xnor UO_1085 (O_1085,N_14834,N_14913);
and UO_1086 (O_1086,N_14884,N_14994);
or UO_1087 (O_1087,N_14970,N_14985);
xor UO_1088 (O_1088,N_14814,N_14979);
nand UO_1089 (O_1089,N_14983,N_14826);
nand UO_1090 (O_1090,N_14808,N_14854);
nand UO_1091 (O_1091,N_14946,N_14905);
nor UO_1092 (O_1092,N_14809,N_14953);
nand UO_1093 (O_1093,N_14886,N_14804);
nand UO_1094 (O_1094,N_14919,N_14957);
xnor UO_1095 (O_1095,N_14817,N_14861);
and UO_1096 (O_1096,N_14852,N_14948);
nand UO_1097 (O_1097,N_14980,N_14869);
nand UO_1098 (O_1098,N_14917,N_14844);
nor UO_1099 (O_1099,N_14946,N_14995);
or UO_1100 (O_1100,N_14901,N_14813);
or UO_1101 (O_1101,N_14800,N_14855);
nand UO_1102 (O_1102,N_14800,N_14932);
nor UO_1103 (O_1103,N_14950,N_14833);
nor UO_1104 (O_1104,N_14938,N_14853);
and UO_1105 (O_1105,N_14858,N_14873);
and UO_1106 (O_1106,N_14890,N_14815);
nand UO_1107 (O_1107,N_14975,N_14860);
or UO_1108 (O_1108,N_14840,N_14991);
and UO_1109 (O_1109,N_14889,N_14834);
xor UO_1110 (O_1110,N_14910,N_14803);
nand UO_1111 (O_1111,N_14801,N_14915);
xor UO_1112 (O_1112,N_14854,N_14921);
or UO_1113 (O_1113,N_14983,N_14870);
or UO_1114 (O_1114,N_14914,N_14939);
xnor UO_1115 (O_1115,N_14993,N_14971);
or UO_1116 (O_1116,N_14867,N_14859);
nand UO_1117 (O_1117,N_14893,N_14826);
xnor UO_1118 (O_1118,N_14818,N_14879);
nor UO_1119 (O_1119,N_14845,N_14843);
nor UO_1120 (O_1120,N_14826,N_14887);
or UO_1121 (O_1121,N_14910,N_14930);
nor UO_1122 (O_1122,N_14894,N_14876);
and UO_1123 (O_1123,N_14843,N_14888);
nor UO_1124 (O_1124,N_14838,N_14987);
nand UO_1125 (O_1125,N_14934,N_14997);
nand UO_1126 (O_1126,N_14881,N_14984);
and UO_1127 (O_1127,N_14986,N_14845);
xnor UO_1128 (O_1128,N_14925,N_14847);
and UO_1129 (O_1129,N_14974,N_14901);
nand UO_1130 (O_1130,N_14888,N_14939);
xor UO_1131 (O_1131,N_14965,N_14877);
or UO_1132 (O_1132,N_14852,N_14881);
nor UO_1133 (O_1133,N_14821,N_14955);
nor UO_1134 (O_1134,N_14843,N_14825);
nor UO_1135 (O_1135,N_14812,N_14966);
nand UO_1136 (O_1136,N_14947,N_14880);
xnor UO_1137 (O_1137,N_14844,N_14882);
nor UO_1138 (O_1138,N_14903,N_14890);
nor UO_1139 (O_1139,N_14833,N_14898);
nand UO_1140 (O_1140,N_14889,N_14908);
or UO_1141 (O_1141,N_14909,N_14960);
nand UO_1142 (O_1142,N_14948,N_14939);
xnor UO_1143 (O_1143,N_14807,N_14987);
nor UO_1144 (O_1144,N_14923,N_14838);
nor UO_1145 (O_1145,N_14856,N_14926);
or UO_1146 (O_1146,N_14885,N_14901);
or UO_1147 (O_1147,N_14800,N_14848);
xnor UO_1148 (O_1148,N_14804,N_14954);
nor UO_1149 (O_1149,N_14918,N_14926);
nor UO_1150 (O_1150,N_14808,N_14877);
or UO_1151 (O_1151,N_14853,N_14901);
nor UO_1152 (O_1152,N_14811,N_14995);
nor UO_1153 (O_1153,N_14853,N_14963);
nor UO_1154 (O_1154,N_14985,N_14921);
or UO_1155 (O_1155,N_14847,N_14916);
nor UO_1156 (O_1156,N_14895,N_14952);
nand UO_1157 (O_1157,N_14854,N_14931);
xnor UO_1158 (O_1158,N_14911,N_14920);
or UO_1159 (O_1159,N_14892,N_14825);
nor UO_1160 (O_1160,N_14890,N_14837);
and UO_1161 (O_1161,N_14972,N_14888);
and UO_1162 (O_1162,N_14952,N_14989);
or UO_1163 (O_1163,N_14841,N_14898);
nor UO_1164 (O_1164,N_14852,N_14860);
nand UO_1165 (O_1165,N_14892,N_14931);
and UO_1166 (O_1166,N_14906,N_14995);
nor UO_1167 (O_1167,N_14865,N_14982);
xnor UO_1168 (O_1168,N_14881,N_14886);
nand UO_1169 (O_1169,N_14967,N_14909);
nor UO_1170 (O_1170,N_14975,N_14837);
or UO_1171 (O_1171,N_14959,N_14973);
xor UO_1172 (O_1172,N_14988,N_14884);
and UO_1173 (O_1173,N_14999,N_14921);
or UO_1174 (O_1174,N_14823,N_14923);
nor UO_1175 (O_1175,N_14989,N_14963);
and UO_1176 (O_1176,N_14804,N_14926);
and UO_1177 (O_1177,N_14843,N_14844);
and UO_1178 (O_1178,N_14952,N_14900);
nor UO_1179 (O_1179,N_14955,N_14826);
nand UO_1180 (O_1180,N_14840,N_14965);
nor UO_1181 (O_1181,N_14947,N_14992);
xor UO_1182 (O_1182,N_14885,N_14933);
xor UO_1183 (O_1183,N_14890,N_14865);
nor UO_1184 (O_1184,N_14869,N_14824);
nor UO_1185 (O_1185,N_14966,N_14916);
nor UO_1186 (O_1186,N_14881,N_14950);
or UO_1187 (O_1187,N_14954,N_14987);
or UO_1188 (O_1188,N_14875,N_14924);
or UO_1189 (O_1189,N_14829,N_14819);
and UO_1190 (O_1190,N_14878,N_14824);
nand UO_1191 (O_1191,N_14848,N_14935);
and UO_1192 (O_1192,N_14831,N_14984);
xnor UO_1193 (O_1193,N_14935,N_14827);
xnor UO_1194 (O_1194,N_14971,N_14873);
xnor UO_1195 (O_1195,N_14820,N_14806);
nand UO_1196 (O_1196,N_14943,N_14864);
nand UO_1197 (O_1197,N_14842,N_14978);
and UO_1198 (O_1198,N_14987,N_14941);
or UO_1199 (O_1199,N_14983,N_14808);
xnor UO_1200 (O_1200,N_14920,N_14998);
nor UO_1201 (O_1201,N_14958,N_14873);
nand UO_1202 (O_1202,N_14881,N_14944);
or UO_1203 (O_1203,N_14822,N_14804);
xor UO_1204 (O_1204,N_14924,N_14943);
xnor UO_1205 (O_1205,N_14971,N_14875);
or UO_1206 (O_1206,N_14848,N_14906);
or UO_1207 (O_1207,N_14996,N_14926);
or UO_1208 (O_1208,N_14926,N_14817);
xor UO_1209 (O_1209,N_14933,N_14974);
or UO_1210 (O_1210,N_14876,N_14866);
nor UO_1211 (O_1211,N_14827,N_14812);
nand UO_1212 (O_1212,N_14891,N_14926);
nand UO_1213 (O_1213,N_14805,N_14906);
xnor UO_1214 (O_1214,N_14836,N_14886);
nand UO_1215 (O_1215,N_14989,N_14924);
and UO_1216 (O_1216,N_14910,N_14848);
nor UO_1217 (O_1217,N_14832,N_14890);
nor UO_1218 (O_1218,N_14887,N_14978);
xnor UO_1219 (O_1219,N_14945,N_14816);
or UO_1220 (O_1220,N_14921,N_14974);
xnor UO_1221 (O_1221,N_14975,N_14843);
xnor UO_1222 (O_1222,N_14865,N_14976);
nor UO_1223 (O_1223,N_14934,N_14909);
nand UO_1224 (O_1224,N_14900,N_14834);
nor UO_1225 (O_1225,N_14829,N_14924);
nand UO_1226 (O_1226,N_14871,N_14921);
xor UO_1227 (O_1227,N_14992,N_14904);
nand UO_1228 (O_1228,N_14844,N_14877);
and UO_1229 (O_1229,N_14969,N_14998);
xnor UO_1230 (O_1230,N_14977,N_14981);
and UO_1231 (O_1231,N_14990,N_14931);
nand UO_1232 (O_1232,N_14943,N_14961);
or UO_1233 (O_1233,N_14908,N_14805);
nand UO_1234 (O_1234,N_14882,N_14922);
or UO_1235 (O_1235,N_14856,N_14925);
or UO_1236 (O_1236,N_14857,N_14910);
xor UO_1237 (O_1237,N_14810,N_14856);
xor UO_1238 (O_1238,N_14958,N_14902);
xnor UO_1239 (O_1239,N_14858,N_14990);
nor UO_1240 (O_1240,N_14855,N_14887);
xor UO_1241 (O_1241,N_14936,N_14807);
xor UO_1242 (O_1242,N_14907,N_14988);
nor UO_1243 (O_1243,N_14806,N_14972);
or UO_1244 (O_1244,N_14814,N_14840);
or UO_1245 (O_1245,N_14888,N_14912);
or UO_1246 (O_1246,N_14897,N_14832);
nor UO_1247 (O_1247,N_14955,N_14827);
and UO_1248 (O_1248,N_14861,N_14969);
nand UO_1249 (O_1249,N_14818,N_14840);
and UO_1250 (O_1250,N_14925,N_14954);
nand UO_1251 (O_1251,N_14813,N_14871);
xor UO_1252 (O_1252,N_14923,N_14973);
and UO_1253 (O_1253,N_14900,N_14825);
nand UO_1254 (O_1254,N_14920,N_14992);
xor UO_1255 (O_1255,N_14860,N_14932);
nand UO_1256 (O_1256,N_14879,N_14817);
nand UO_1257 (O_1257,N_14872,N_14981);
or UO_1258 (O_1258,N_14991,N_14862);
and UO_1259 (O_1259,N_14968,N_14918);
and UO_1260 (O_1260,N_14856,N_14995);
or UO_1261 (O_1261,N_14818,N_14871);
nor UO_1262 (O_1262,N_14807,N_14842);
and UO_1263 (O_1263,N_14934,N_14998);
nor UO_1264 (O_1264,N_14977,N_14989);
nor UO_1265 (O_1265,N_14844,N_14828);
nor UO_1266 (O_1266,N_14934,N_14811);
nor UO_1267 (O_1267,N_14976,N_14842);
nand UO_1268 (O_1268,N_14819,N_14934);
xnor UO_1269 (O_1269,N_14837,N_14988);
nor UO_1270 (O_1270,N_14801,N_14829);
xnor UO_1271 (O_1271,N_14950,N_14921);
nor UO_1272 (O_1272,N_14819,N_14917);
and UO_1273 (O_1273,N_14847,N_14991);
nand UO_1274 (O_1274,N_14909,N_14941);
and UO_1275 (O_1275,N_14864,N_14938);
or UO_1276 (O_1276,N_14965,N_14926);
and UO_1277 (O_1277,N_14946,N_14809);
nand UO_1278 (O_1278,N_14805,N_14845);
nand UO_1279 (O_1279,N_14889,N_14874);
nand UO_1280 (O_1280,N_14811,N_14950);
xor UO_1281 (O_1281,N_14881,N_14996);
or UO_1282 (O_1282,N_14866,N_14806);
and UO_1283 (O_1283,N_14859,N_14829);
xnor UO_1284 (O_1284,N_14847,N_14839);
xor UO_1285 (O_1285,N_14828,N_14866);
nor UO_1286 (O_1286,N_14946,N_14819);
nand UO_1287 (O_1287,N_14907,N_14970);
and UO_1288 (O_1288,N_14947,N_14999);
nand UO_1289 (O_1289,N_14830,N_14897);
xor UO_1290 (O_1290,N_14973,N_14961);
nor UO_1291 (O_1291,N_14864,N_14820);
nand UO_1292 (O_1292,N_14839,N_14829);
nor UO_1293 (O_1293,N_14909,N_14824);
and UO_1294 (O_1294,N_14886,N_14816);
nor UO_1295 (O_1295,N_14816,N_14849);
or UO_1296 (O_1296,N_14902,N_14987);
nor UO_1297 (O_1297,N_14824,N_14981);
xnor UO_1298 (O_1298,N_14810,N_14909);
and UO_1299 (O_1299,N_14950,N_14911);
xor UO_1300 (O_1300,N_14895,N_14846);
xor UO_1301 (O_1301,N_14834,N_14835);
and UO_1302 (O_1302,N_14991,N_14997);
nor UO_1303 (O_1303,N_14828,N_14980);
and UO_1304 (O_1304,N_14826,N_14897);
nor UO_1305 (O_1305,N_14819,N_14813);
nor UO_1306 (O_1306,N_14887,N_14985);
xor UO_1307 (O_1307,N_14902,N_14814);
or UO_1308 (O_1308,N_14844,N_14879);
nand UO_1309 (O_1309,N_14966,N_14839);
xor UO_1310 (O_1310,N_14978,N_14929);
nand UO_1311 (O_1311,N_14893,N_14841);
xnor UO_1312 (O_1312,N_14969,N_14840);
nand UO_1313 (O_1313,N_14918,N_14956);
xnor UO_1314 (O_1314,N_14874,N_14861);
and UO_1315 (O_1315,N_14869,N_14870);
nor UO_1316 (O_1316,N_14863,N_14811);
or UO_1317 (O_1317,N_14811,N_14904);
or UO_1318 (O_1318,N_14819,N_14921);
nand UO_1319 (O_1319,N_14802,N_14838);
xor UO_1320 (O_1320,N_14927,N_14801);
and UO_1321 (O_1321,N_14810,N_14920);
nand UO_1322 (O_1322,N_14965,N_14914);
nor UO_1323 (O_1323,N_14857,N_14861);
or UO_1324 (O_1324,N_14889,N_14946);
nand UO_1325 (O_1325,N_14907,N_14802);
xnor UO_1326 (O_1326,N_14970,N_14867);
xor UO_1327 (O_1327,N_14801,N_14934);
xnor UO_1328 (O_1328,N_14979,N_14833);
and UO_1329 (O_1329,N_14804,N_14983);
xor UO_1330 (O_1330,N_14974,N_14927);
nand UO_1331 (O_1331,N_14807,N_14933);
nand UO_1332 (O_1332,N_14960,N_14955);
and UO_1333 (O_1333,N_14931,N_14801);
and UO_1334 (O_1334,N_14967,N_14861);
or UO_1335 (O_1335,N_14816,N_14904);
and UO_1336 (O_1336,N_14800,N_14826);
nand UO_1337 (O_1337,N_14936,N_14915);
and UO_1338 (O_1338,N_14973,N_14974);
xor UO_1339 (O_1339,N_14933,N_14826);
nor UO_1340 (O_1340,N_14890,N_14810);
xor UO_1341 (O_1341,N_14866,N_14894);
or UO_1342 (O_1342,N_14834,N_14856);
xnor UO_1343 (O_1343,N_14886,N_14979);
and UO_1344 (O_1344,N_14968,N_14873);
nor UO_1345 (O_1345,N_14914,N_14904);
xor UO_1346 (O_1346,N_14987,N_14887);
xnor UO_1347 (O_1347,N_14849,N_14888);
or UO_1348 (O_1348,N_14879,N_14928);
nor UO_1349 (O_1349,N_14975,N_14897);
nand UO_1350 (O_1350,N_14970,N_14814);
and UO_1351 (O_1351,N_14820,N_14800);
and UO_1352 (O_1352,N_14878,N_14919);
and UO_1353 (O_1353,N_14941,N_14922);
nand UO_1354 (O_1354,N_14877,N_14888);
and UO_1355 (O_1355,N_14880,N_14910);
and UO_1356 (O_1356,N_14928,N_14944);
nor UO_1357 (O_1357,N_14962,N_14839);
or UO_1358 (O_1358,N_14801,N_14947);
nor UO_1359 (O_1359,N_14906,N_14901);
nand UO_1360 (O_1360,N_14939,N_14963);
or UO_1361 (O_1361,N_14811,N_14823);
or UO_1362 (O_1362,N_14836,N_14808);
or UO_1363 (O_1363,N_14996,N_14896);
or UO_1364 (O_1364,N_14861,N_14961);
xor UO_1365 (O_1365,N_14978,N_14934);
xnor UO_1366 (O_1366,N_14937,N_14837);
nand UO_1367 (O_1367,N_14845,N_14885);
and UO_1368 (O_1368,N_14917,N_14900);
nand UO_1369 (O_1369,N_14902,N_14826);
xnor UO_1370 (O_1370,N_14979,N_14899);
nand UO_1371 (O_1371,N_14886,N_14830);
and UO_1372 (O_1372,N_14823,N_14875);
and UO_1373 (O_1373,N_14870,N_14996);
or UO_1374 (O_1374,N_14850,N_14918);
or UO_1375 (O_1375,N_14867,N_14979);
nand UO_1376 (O_1376,N_14941,N_14818);
nand UO_1377 (O_1377,N_14929,N_14885);
or UO_1378 (O_1378,N_14990,N_14903);
or UO_1379 (O_1379,N_14976,N_14945);
or UO_1380 (O_1380,N_14909,N_14937);
or UO_1381 (O_1381,N_14838,N_14872);
and UO_1382 (O_1382,N_14878,N_14863);
and UO_1383 (O_1383,N_14812,N_14944);
nor UO_1384 (O_1384,N_14999,N_14938);
or UO_1385 (O_1385,N_14889,N_14924);
and UO_1386 (O_1386,N_14825,N_14899);
and UO_1387 (O_1387,N_14813,N_14853);
nor UO_1388 (O_1388,N_14938,N_14995);
or UO_1389 (O_1389,N_14968,N_14905);
and UO_1390 (O_1390,N_14832,N_14842);
or UO_1391 (O_1391,N_14982,N_14959);
or UO_1392 (O_1392,N_14827,N_14828);
nand UO_1393 (O_1393,N_14833,N_14944);
or UO_1394 (O_1394,N_14886,N_14834);
xor UO_1395 (O_1395,N_14892,N_14843);
or UO_1396 (O_1396,N_14821,N_14961);
nand UO_1397 (O_1397,N_14827,N_14858);
nand UO_1398 (O_1398,N_14855,N_14905);
xnor UO_1399 (O_1399,N_14956,N_14812);
and UO_1400 (O_1400,N_14800,N_14995);
nand UO_1401 (O_1401,N_14883,N_14845);
xor UO_1402 (O_1402,N_14842,N_14954);
nand UO_1403 (O_1403,N_14954,N_14923);
or UO_1404 (O_1404,N_14931,N_14816);
nor UO_1405 (O_1405,N_14946,N_14959);
nand UO_1406 (O_1406,N_14861,N_14809);
nor UO_1407 (O_1407,N_14960,N_14976);
nand UO_1408 (O_1408,N_14910,N_14911);
nand UO_1409 (O_1409,N_14951,N_14830);
or UO_1410 (O_1410,N_14871,N_14808);
and UO_1411 (O_1411,N_14926,N_14805);
nor UO_1412 (O_1412,N_14944,N_14964);
and UO_1413 (O_1413,N_14995,N_14829);
and UO_1414 (O_1414,N_14906,N_14981);
xor UO_1415 (O_1415,N_14962,N_14891);
nor UO_1416 (O_1416,N_14902,N_14962);
xnor UO_1417 (O_1417,N_14854,N_14963);
or UO_1418 (O_1418,N_14954,N_14929);
or UO_1419 (O_1419,N_14868,N_14844);
xnor UO_1420 (O_1420,N_14876,N_14996);
nor UO_1421 (O_1421,N_14814,N_14957);
or UO_1422 (O_1422,N_14965,N_14956);
nor UO_1423 (O_1423,N_14997,N_14940);
or UO_1424 (O_1424,N_14842,N_14819);
xnor UO_1425 (O_1425,N_14917,N_14824);
or UO_1426 (O_1426,N_14978,N_14966);
and UO_1427 (O_1427,N_14915,N_14950);
nand UO_1428 (O_1428,N_14808,N_14827);
nand UO_1429 (O_1429,N_14896,N_14927);
and UO_1430 (O_1430,N_14899,N_14936);
nor UO_1431 (O_1431,N_14935,N_14805);
nor UO_1432 (O_1432,N_14810,N_14849);
nand UO_1433 (O_1433,N_14890,N_14824);
nand UO_1434 (O_1434,N_14838,N_14912);
and UO_1435 (O_1435,N_14942,N_14833);
and UO_1436 (O_1436,N_14939,N_14876);
or UO_1437 (O_1437,N_14921,N_14838);
or UO_1438 (O_1438,N_14940,N_14969);
nor UO_1439 (O_1439,N_14976,N_14925);
nand UO_1440 (O_1440,N_14850,N_14951);
nand UO_1441 (O_1441,N_14877,N_14980);
and UO_1442 (O_1442,N_14919,N_14996);
or UO_1443 (O_1443,N_14845,N_14969);
nor UO_1444 (O_1444,N_14823,N_14873);
nand UO_1445 (O_1445,N_14972,N_14843);
nor UO_1446 (O_1446,N_14835,N_14858);
or UO_1447 (O_1447,N_14856,N_14865);
nor UO_1448 (O_1448,N_14913,N_14840);
or UO_1449 (O_1449,N_14844,N_14912);
xnor UO_1450 (O_1450,N_14852,N_14845);
nor UO_1451 (O_1451,N_14823,N_14991);
nor UO_1452 (O_1452,N_14823,N_14938);
xnor UO_1453 (O_1453,N_14958,N_14886);
and UO_1454 (O_1454,N_14909,N_14964);
nand UO_1455 (O_1455,N_14876,N_14867);
nor UO_1456 (O_1456,N_14837,N_14909);
xor UO_1457 (O_1457,N_14863,N_14846);
nor UO_1458 (O_1458,N_14807,N_14901);
nor UO_1459 (O_1459,N_14890,N_14994);
and UO_1460 (O_1460,N_14981,N_14836);
nand UO_1461 (O_1461,N_14816,N_14939);
nor UO_1462 (O_1462,N_14996,N_14807);
or UO_1463 (O_1463,N_14923,N_14887);
xnor UO_1464 (O_1464,N_14825,N_14993);
or UO_1465 (O_1465,N_14848,N_14923);
or UO_1466 (O_1466,N_14996,N_14851);
nor UO_1467 (O_1467,N_14839,N_14958);
xor UO_1468 (O_1468,N_14962,N_14982);
nand UO_1469 (O_1469,N_14822,N_14854);
and UO_1470 (O_1470,N_14835,N_14981);
and UO_1471 (O_1471,N_14828,N_14993);
and UO_1472 (O_1472,N_14867,N_14960);
nand UO_1473 (O_1473,N_14860,N_14988);
xnor UO_1474 (O_1474,N_14929,N_14886);
nand UO_1475 (O_1475,N_14927,N_14820);
or UO_1476 (O_1476,N_14875,N_14960);
nor UO_1477 (O_1477,N_14978,N_14843);
nor UO_1478 (O_1478,N_14993,N_14826);
nor UO_1479 (O_1479,N_14998,N_14894);
xnor UO_1480 (O_1480,N_14962,N_14911);
and UO_1481 (O_1481,N_14834,N_14978);
xor UO_1482 (O_1482,N_14825,N_14976);
nand UO_1483 (O_1483,N_14852,N_14987);
xor UO_1484 (O_1484,N_14887,N_14830);
and UO_1485 (O_1485,N_14805,N_14909);
nand UO_1486 (O_1486,N_14944,N_14889);
or UO_1487 (O_1487,N_14818,N_14826);
or UO_1488 (O_1488,N_14960,N_14820);
nand UO_1489 (O_1489,N_14985,N_14971);
or UO_1490 (O_1490,N_14990,N_14846);
nand UO_1491 (O_1491,N_14816,N_14937);
xor UO_1492 (O_1492,N_14854,N_14997);
xnor UO_1493 (O_1493,N_14815,N_14897);
xor UO_1494 (O_1494,N_14991,N_14941);
xnor UO_1495 (O_1495,N_14988,N_14878);
or UO_1496 (O_1496,N_14881,N_14861);
and UO_1497 (O_1497,N_14951,N_14995);
or UO_1498 (O_1498,N_14900,N_14816);
nand UO_1499 (O_1499,N_14846,N_14975);
xnor UO_1500 (O_1500,N_14964,N_14934);
or UO_1501 (O_1501,N_14831,N_14810);
nand UO_1502 (O_1502,N_14987,N_14880);
nor UO_1503 (O_1503,N_14936,N_14828);
xor UO_1504 (O_1504,N_14810,N_14893);
nand UO_1505 (O_1505,N_14919,N_14887);
or UO_1506 (O_1506,N_14867,N_14915);
nand UO_1507 (O_1507,N_14928,N_14997);
nand UO_1508 (O_1508,N_14970,N_14874);
xnor UO_1509 (O_1509,N_14850,N_14898);
and UO_1510 (O_1510,N_14877,N_14880);
xnor UO_1511 (O_1511,N_14945,N_14841);
nand UO_1512 (O_1512,N_14900,N_14925);
nor UO_1513 (O_1513,N_14972,N_14801);
nand UO_1514 (O_1514,N_14881,N_14943);
and UO_1515 (O_1515,N_14863,N_14935);
and UO_1516 (O_1516,N_14845,N_14899);
nor UO_1517 (O_1517,N_14836,N_14922);
nand UO_1518 (O_1518,N_14901,N_14861);
or UO_1519 (O_1519,N_14806,N_14828);
or UO_1520 (O_1520,N_14810,N_14936);
and UO_1521 (O_1521,N_14870,N_14855);
xnor UO_1522 (O_1522,N_14971,N_14957);
xnor UO_1523 (O_1523,N_14951,N_14834);
xnor UO_1524 (O_1524,N_14848,N_14885);
nand UO_1525 (O_1525,N_14881,N_14981);
nand UO_1526 (O_1526,N_14819,N_14978);
xor UO_1527 (O_1527,N_14986,N_14871);
nand UO_1528 (O_1528,N_14958,N_14975);
or UO_1529 (O_1529,N_14829,N_14933);
nand UO_1530 (O_1530,N_14953,N_14903);
nor UO_1531 (O_1531,N_14838,N_14878);
nand UO_1532 (O_1532,N_14922,N_14850);
nor UO_1533 (O_1533,N_14857,N_14954);
and UO_1534 (O_1534,N_14819,N_14965);
nand UO_1535 (O_1535,N_14903,N_14868);
xnor UO_1536 (O_1536,N_14967,N_14838);
xor UO_1537 (O_1537,N_14921,N_14899);
and UO_1538 (O_1538,N_14865,N_14881);
xor UO_1539 (O_1539,N_14845,N_14826);
or UO_1540 (O_1540,N_14951,N_14892);
nor UO_1541 (O_1541,N_14835,N_14895);
nand UO_1542 (O_1542,N_14956,N_14999);
nand UO_1543 (O_1543,N_14909,N_14977);
nor UO_1544 (O_1544,N_14886,N_14818);
xnor UO_1545 (O_1545,N_14891,N_14979);
or UO_1546 (O_1546,N_14939,N_14821);
or UO_1547 (O_1547,N_14899,N_14864);
and UO_1548 (O_1548,N_14902,N_14851);
nand UO_1549 (O_1549,N_14888,N_14938);
nor UO_1550 (O_1550,N_14845,N_14947);
nand UO_1551 (O_1551,N_14923,N_14802);
or UO_1552 (O_1552,N_14908,N_14806);
and UO_1553 (O_1553,N_14824,N_14898);
nor UO_1554 (O_1554,N_14800,N_14988);
or UO_1555 (O_1555,N_14989,N_14824);
and UO_1556 (O_1556,N_14829,N_14981);
and UO_1557 (O_1557,N_14937,N_14917);
and UO_1558 (O_1558,N_14831,N_14933);
or UO_1559 (O_1559,N_14992,N_14964);
or UO_1560 (O_1560,N_14904,N_14828);
or UO_1561 (O_1561,N_14843,N_14926);
nor UO_1562 (O_1562,N_14960,N_14868);
nand UO_1563 (O_1563,N_14881,N_14814);
nand UO_1564 (O_1564,N_14975,N_14946);
nand UO_1565 (O_1565,N_14865,N_14953);
xnor UO_1566 (O_1566,N_14976,N_14841);
and UO_1567 (O_1567,N_14831,N_14835);
or UO_1568 (O_1568,N_14871,N_14915);
and UO_1569 (O_1569,N_14988,N_14802);
nand UO_1570 (O_1570,N_14849,N_14834);
and UO_1571 (O_1571,N_14915,N_14831);
and UO_1572 (O_1572,N_14912,N_14801);
xor UO_1573 (O_1573,N_14959,N_14977);
and UO_1574 (O_1574,N_14930,N_14912);
nor UO_1575 (O_1575,N_14961,N_14811);
or UO_1576 (O_1576,N_14980,N_14863);
nor UO_1577 (O_1577,N_14831,N_14861);
xor UO_1578 (O_1578,N_14869,N_14969);
nand UO_1579 (O_1579,N_14847,N_14860);
or UO_1580 (O_1580,N_14801,N_14884);
nor UO_1581 (O_1581,N_14993,N_14830);
nor UO_1582 (O_1582,N_14851,N_14966);
nor UO_1583 (O_1583,N_14951,N_14827);
xor UO_1584 (O_1584,N_14822,N_14972);
or UO_1585 (O_1585,N_14950,N_14870);
and UO_1586 (O_1586,N_14835,N_14997);
nand UO_1587 (O_1587,N_14992,N_14994);
or UO_1588 (O_1588,N_14812,N_14804);
nand UO_1589 (O_1589,N_14951,N_14970);
nand UO_1590 (O_1590,N_14818,N_14922);
nor UO_1591 (O_1591,N_14816,N_14988);
xnor UO_1592 (O_1592,N_14972,N_14841);
or UO_1593 (O_1593,N_14829,N_14832);
or UO_1594 (O_1594,N_14983,N_14955);
and UO_1595 (O_1595,N_14975,N_14880);
nand UO_1596 (O_1596,N_14852,N_14946);
or UO_1597 (O_1597,N_14885,N_14925);
and UO_1598 (O_1598,N_14996,N_14814);
or UO_1599 (O_1599,N_14845,N_14846);
xnor UO_1600 (O_1600,N_14933,N_14887);
xnor UO_1601 (O_1601,N_14856,N_14996);
or UO_1602 (O_1602,N_14898,N_14887);
or UO_1603 (O_1603,N_14805,N_14886);
nor UO_1604 (O_1604,N_14910,N_14994);
nor UO_1605 (O_1605,N_14898,N_14878);
and UO_1606 (O_1606,N_14808,N_14932);
nor UO_1607 (O_1607,N_14965,N_14809);
nor UO_1608 (O_1608,N_14951,N_14993);
and UO_1609 (O_1609,N_14857,N_14961);
nor UO_1610 (O_1610,N_14907,N_14847);
or UO_1611 (O_1611,N_14946,N_14877);
and UO_1612 (O_1612,N_14821,N_14895);
and UO_1613 (O_1613,N_14953,N_14820);
nand UO_1614 (O_1614,N_14886,N_14964);
and UO_1615 (O_1615,N_14973,N_14948);
nand UO_1616 (O_1616,N_14888,N_14899);
xnor UO_1617 (O_1617,N_14872,N_14914);
or UO_1618 (O_1618,N_14874,N_14996);
xor UO_1619 (O_1619,N_14815,N_14997);
nor UO_1620 (O_1620,N_14945,N_14811);
nand UO_1621 (O_1621,N_14961,N_14966);
and UO_1622 (O_1622,N_14904,N_14906);
nor UO_1623 (O_1623,N_14948,N_14810);
xor UO_1624 (O_1624,N_14963,N_14882);
xor UO_1625 (O_1625,N_14984,N_14887);
xor UO_1626 (O_1626,N_14997,N_14860);
xnor UO_1627 (O_1627,N_14906,N_14846);
or UO_1628 (O_1628,N_14924,N_14865);
nand UO_1629 (O_1629,N_14953,N_14924);
and UO_1630 (O_1630,N_14850,N_14985);
and UO_1631 (O_1631,N_14980,N_14996);
or UO_1632 (O_1632,N_14871,N_14972);
nor UO_1633 (O_1633,N_14824,N_14960);
xor UO_1634 (O_1634,N_14986,N_14826);
and UO_1635 (O_1635,N_14955,N_14897);
or UO_1636 (O_1636,N_14855,N_14937);
xor UO_1637 (O_1637,N_14856,N_14815);
and UO_1638 (O_1638,N_14804,N_14800);
nand UO_1639 (O_1639,N_14959,N_14934);
nor UO_1640 (O_1640,N_14900,N_14826);
nor UO_1641 (O_1641,N_14823,N_14810);
xnor UO_1642 (O_1642,N_14875,N_14871);
or UO_1643 (O_1643,N_14844,N_14819);
nor UO_1644 (O_1644,N_14958,N_14906);
xor UO_1645 (O_1645,N_14977,N_14806);
xor UO_1646 (O_1646,N_14903,N_14952);
and UO_1647 (O_1647,N_14915,N_14800);
and UO_1648 (O_1648,N_14962,N_14963);
xor UO_1649 (O_1649,N_14868,N_14864);
or UO_1650 (O_1650,N_14903,N_14997);
or UO_1651 (O_1651,N_14975,N_14829);
and UO_1652 (O_1652,N_14974,N_14961);
nand UO_1653 (O_1653,N_14995,N_14931);
or UO_1654 (O_1654,N_14960,N_14947);
or UO_1655 (O_1655,N_14830,N_14939);
nor UO_1656 (O_1656,N_14979,N_14986);
and UO_1657 (O_1657,N_14896,N_14850);
and UO_1658 (O_1658,N_14848,N_14957);
and UO_1659 (O_1659,N_14988,N_14819);
or UO_1660 (O_1660,N_14999,N_14880);
nand UO_1661 (O_1661,N_14836,N_14810);
nand UO_1662 (O_1662,N_14911,N_14894);
nand UO_1663 (O_1663,N_14871,N_14910);
nand UO_1664 (O_1664,N_14802,N_14878);
nor UO_1665 (O_1665,N_14818,N_14939);
nand UO_1666 (O_1666,N_14917,N_14959);
xnor UO_1667 (O_1667,N_14954,N_14975);
or UO_1668 (O_1668,N_14958,N_14889);
or UO_1669 (O_1669,N_14868,N_14815);
xor UO_1670 (O_1670,N_14810,N_14896);
xnor UO_1671 (O_1671,N_14935,N_14804);
and UO_1672 (O_1672,N_14863,N_14862);
or UO_1673 (O_1673,N_14985,N_14812);
and UO_1674 (O_1674,N_14920,N_14801);
nand UO_1675 (O_1675,N_14877,N_14866);
nor UO_1676 (O_1676,N_14860,N_14987);
nor UO_1677 (O_1677,N_14924,N_14852);
nor UO_1678 (O_1678,N_14899,N_14905);
nor UO_1679 (O_1679,N_14985,N_14800);
or UO_1680 (O_1680,N_14945,N_14857);
nor UO_1681 (O_1681,N_14915,N_14880);
and UO_1682 (O_1682,N_14881,N_14925);
nand UO_1683 (O_1683,N_14959,N_14810);
nand UO_1684 (O_1684,N_14933,N_14965);
xnor UO_1685 (O_1685,N_14983,N_14999);
or UO_1686 (O_1686,N_14812,N_14883);
and UO_1687 (O_1687,N_14868,N_14921);
and UO_1688 (O_1688,N_14981,N_14962);
xnor UO_1689 (O_1689,N_14847,N_14938);
nand UO_1690 (O_1690,N_14940,N_14899);
and UO_1691 (O_1691,N_14903,N_14910);
nand UO_1692 (O_1692,N_14988,N_14910);
nand UO_1693 (O_1693,N_14950,N_14936);
nor UO_1694 (O_1694,N_14838,N_14889);
or UO_1695 (O_1695,N_14839,N_14906);
and UO_1696 (O_1696,N_14864,N_14977);
xor UO_1697 (O_1697,N_14924,N_14984);
nand UO_1698 (O_1698,N_14928,N_14925);
nand UO_1699 (O_1699,N_14914,N_14871);
nor UO_1700 (O_1700,N_14962,N_14865);
nor UO_1701 (O_1701,N_14919,N_14817);
xnor UO_1702 (O_1702,N_14917,N_14845);
nor UO_1703 (O_1703,N_14876,N_14934);
xnor UO_1704 (O_1704,N_14991,N_14819);
nand UO_1705 (O_1705,N_14863,N_14879);
and UO_1706 (O_1706,N_14988,N_14826);
or UO_1707 (O_1707,N_14985,N_14993);
xnor UO_1708 (O_1708,N_14879,N_14847);
and UO_1709 (O_1709,N_14810,N_14880);
or UO_1710 (O_1710,N_14858,N_14898);
or UO_1711 (O_1711,N_14825,N_14816);
xnor UO_1712 (O_1712,N_14990,N_14879);
or UO_1713 (O_1713,N_14988,N_14871);
xor UO_1714 (O_1714,N_14970,N_14833);
xor UO_1715 (O_1715,N_14913,N_14866);
or UO_1716 (O_1716,N_14907,N_14871);
or UO_1717 (O_1717,N_14994,N_14822);
and UO_1718 (O_1718,N_14862,N_14814);
and UO_1719 (O_1719,N_14981,N_14974);
xnor UO_1720 (O_1720,N_14908,N_14999);
nand UO_1721 (O_1721,N_14902,N_14971);
and UO_1722 (O_1722,N_14900,N_14847);
and UO_1723 (O_1723,N_14931,N_14911);
xnor UO_1724 (O_1724,N_14917,N_14995);
or UO_1725 (O_1725,N_14872,N_14863);
xor UO_1726 (O_1726,N_14925,N_14815);
nand UO_1727 (O_1727,N_14890,N_14836);
nor UO_1728 (O_1728,N_14838,N_14832);
or UO_1729 (O_1729,N_14843,N_14894);
or UO_1730 (O_1730,N_14866,N_14857);
nand UO_1731 (O_1731,N_14997,N_14915);
xor UO_1732 (O_1732,N_14965,N_14852);
or UO_1733 (O_1733,N_14956,N_14876);
and UO_1734 (O_1734,N_14849,N_14841);
or UO_1735 (O_1735,N_14879,N_14991);
nor UO_1736 (O_1736,N_14880,N_14893);
nor UO_1737 (O_1737,N_14832,N_14809);
or UO_1738 (O_1738,N_14848,N_14866);
and UO_1739 (O_1739,N_14927,N_14883);
xor UO_1740 (O_1740,N_14823,N_14985);
nand UO_1741 (O_1741,N_14974,N_14819);
or UO_1742 (O_1742,N_14918,N_14907);
nand UO_1743 (O_1743,N_14856,N_14892);
nand UO_1744 (O_1744,N_14893,N_14902);
nor UO_1745 (O_1745,N_14949,N_14848);
nand UO_1746 (O_1746,N_14885,N_14887);
nor UO_1747 (O_1747,N_14807,N_14903);
and UO_1748 (O_1748,N_14890,N_14841);
or UO_1749 (O_1749,N_14843,N_14849);
xnor UO_1750 (O_1750,N_14877,N_14841);
or UO_1751 (O_1751,N_14906,N_14930);
or UO_1752 (O_1752,N_14978,N_14921);
nor UO_1753 (O_1753,N_14913,N_14869);
xnor UO_1754 (O_1754,N_14878,N_14941);
or UO_1755 (O_1755,N_14927,N_14854);
and UO_1756 (O_1756,N_14943,N_14857);
nor UO_1757 (O_1757,N_14851,N_14978);
nand UO_1758 (O_1758,N_14985,N_14988);
and UO_1759 (O_1759,N_14960,N_14966);
and UO_1760 (O_1760,N_14863,N_14920);
xor UO_1761 (O_1761,N_14811,N_14948);
xor UO_1762 (O_1762,N_14894,N_14855);
nand UO_1763 (O_1763,N_14944,N_14982);
nand UO_1764 (O_1764,N_14972,N_14812);
xor UO_1765 (O_1765,N_14931,N_14945);
or UO_1766 (O_1766,N_14982,N_14918);
nor UO_1767 (O_1767,N_14874,N_14833);
or UO_1768 (O_1768,N_14980,N_14928);
nand UO_1769 (O_1769,N_14976,N_14922);
xnor UO_1770 (O_1770,N_14820,N_14818);
xnor UO_1771 (O_1771,N_14856,N_14895);
and UO_1772 (O_1772,N_14864,N_14968);
or UO_1773 (O_1773,N_14906,N_14886);
xnor UO_1774 (O_1774,N_14945,N_14885);
and UO_1775 (O_1775,N_14893,N_14887);
nor UO_1776 (O_1776,N_14947,N_14895);
xor UO_1777 (O_1777,N_14979,N_14830);
or UO_1778 (O_1778,N_14923,N_14804);
and UO_1779 (O_1779,N_14981,N_14924);
nand UO_1780 (O_1780,N_14961,N_14831);
and UO_1781 (O_1781,N_14994,N_14951);
nor UO_1782 (O_1782,N_14894,N_14958);
and UO_1783 (O_1783,N_14996,N_14917);
nor UO_1784 (O_1784,N_14934,N_14890);
nor UO_1785 (O_1785,N_14954,N_14829);
and UO_1786 (O_1786,N_14855,N_14976);
nand UO_1787 (O_1787,N_14986,N_14874);
or UO_1788 (O_1788,N_14983,N_14975);
xor UO_1789 (O_1789,N_14881,N_14835);
nor UO_1790 (O_1790,N_14807,N_14977);
xor UO_1791 (O_1791,N_14962,N_14802);
and UO_1792 (O_1792,N_14932,N_14926);
xnor UO_1793 (O_1793,N_14981,N_14807);
nor UO_1794 (O_1794,N_14921,N_14816);
or UO_1795 (O_1795,N_14958,N_14984);
or UO_1796 (O_1796,N_14890,N_14866);
nor UO_1797 (O_1797,N_14932,N_14847);
and UO_1798 (O_1798,N_14802,N_14997);
and UO_1799 (O_1799,N_14821,N_14902);
nand UO_1800 (O_1800,N_14808,N_14985);
xnor UO_1801 (O_1801,N_14972,N_14996);
nor UO_1802 (O_1802,N_14918,N_14835);
and UO_1803 (O_1803,N_14954,N_14914);
and UO_1804 (O_1804,N_14927,N_14891);
nand UO_1805 (O_1805,N_14958,N_14867);
and UO_1806 (O_1806,N_14841,N_14974);
and UO_1807 (O_1807,N_14846,N_14983);
and UO_1808 (O_1808,N_14810,N_14848);
nand UO_1809 (O_1809,N_14861,N_14997);
and UO_1810 (O_1810,N_14969,N_14943);
nand UO_1811 (O_1811,N_14840,N_14977);
and UO_1812 (O_1812,N_14934,N_14967);
nand UO_1813 (O_1813,N_14877,N_14859);
or UO_1814 (O_1814,N_14808,N_14958);
and UO_1815 (O_1815,N_14951,N_14957);
and UO_1816 (O_1816,N_14976,N_14995);
nor UO_1817 (O_1817,N_14840,N_14851);
nor UO_1818 (O_1818,N_14996,N_14941);
nor UO_1819 (O_1819,N_14968,N_14800);
or UO_1820 (O_1820,N_14959,N_14897);
nand UO_1821 (O_1821,N_14965,N_14881);
xor UO_1822 (O_1822,N_14980,N_14890);
and UO_1823 (O_1823,N_14855,N_14941);
or UO_1824 (O_1824,N_14834,N_14894);
xnor UO_1825 (O_1825,N_14915,N_14942);
and UO_1826 (O_1826,N_14958,N_14924);
or UO_1827 (O_1827,N_14950,N_14919);
and UO_1828 (O_1828,N_14881,N_14975);
and UO_1829 (O_1829,N_14863,N_14967);
or UO_1830 (O_1830,N_14888,N_14860);
nor UO_1831 (O_1831,N_14895,N_14854);
and UO_1832 (O_1832,N_14964,N_14967);
nor UO_1833 (O_1833,N_14825,N_14897);
nand UO_1834 (O_1834,N_14837,N_14964);
nand UO_1835 (O_1835,N_14803,N_14812);
or UO_1836 (O_1836,N_14933,N_14855);
xor UO_1837 (O_1837,N_14950,N_14928);
xnor UO_1838 (O_1838,N_14996,N_14946);
nor UO_1839 (O_1839,N_14964,N_14863);
or UO_1840 (O_1840,N_14878,N_14949);
nand UO_1841 (O_1841,N_14892,N_14846);
nor UO_1842 (O_1842,N_14907,N_14831);
and UO_1843 (O_1843,N_14851,N_14812);
or UO_1844 (O_1844,N_14906,N_14931);
or UO_1845 (O_1845,N_14963,N_14888);
or UO_1846 (O_1846,N_14891,N_14924);
or UO_1847 (O_1847,N_14896,N_14910);
nor UO_1848 (O_1848,N_14967,N_14958);
and UO_1849 (O_1849,N_14935,N_14920);
xnor UO_1850 (O_1850,N_14921,N_14821);
or UO_1851 (O_1851,N_14912,N_14981);
nor UO_1852 (O_1852,N_14982,N_14961);
xor UO_1853 (O_1853,N_14959,N_14953);
and UO_1854 (O_1854,N_14857,N_14868);
or UO_1855 (O_1855,N_14907,N_14851);
and UO_1856 (O_1856,N_14811,N_14878);
and UO_1857 (O_1857,N_14962,N_14960);
nand UO_1858 (O_1858,N_14966,N_14920);
or UO_1859 (O_1859,N_14975,N_14929);
and UO_1860 (O_1860,N_14921,N_14802);
and UO_1861 (O_1861,N_14935,N_14962);
nand UO_1862 (O_1862,N_14970,N_14937);
nand UO_1863 (O_1863,N_14929,N_14990);
and UO_1864 (O_1864,N_14829,N_14901);
and UO_1865 (O_1865,N_14983,N_14957);
xor UO_1866 (O_1866,N_14984,N_14821);
or UO_1867 (O_1867,N_14890,N_14835);
xnor UO_1868 (O_1868,N_14854,N_14977);
xor UO_1869 (O_1869,N_14878,N_14806);
xor UO_1870 (O_1870,N_14987,N_14933);
nor UO_1871 (O_1871,N_14814,N_14807);
xor UO_1872 (O_1872,N_14839,N_14844);
nor UO_1873 (O_1873,N_14873,N_14979);
nor UO_1874 (O_1874,N_14812,N_14918);
nor UO_1875 (O_1875,N_14998,N_14853);
or UO_1876 (O_1876,N_14958,N_14802);
nor UO_1877 (O_1877,N_14965,N_14817);
nand UO_1878 (O_1878,N_14913,N_14875);
nor UO_1879 (O_1879,N_14910,N_14909);
xor UO_1880 (O_1880,N_14865,N_14896);
or UO_1881 (O_1881,N_14993,N_14964);
nor UO_1882 (O_1882,N_14931,N_14941);
nand UO_1883 (O_1883,N_14891,N_14859);
xor UO_1884 (O_1884,N_14810,N_14912);
nor UO_1885 (O_1885,N_14960,N_14815);
nand UO_1886 (O_1886,N_14914,N_14984);
xnor UO_1887 (O_1887,N_14812,N_14904);
or UO_1888 (O_1888,N_14860,N_14940);
xnor UO_1889 (O_1889,N_14825,N_14906);
xor UO_1890 (O_1890,N_14901,N_14812);
nor UO_1891 (O_1891,N_14803,N_14827);
xnor UO_1892 (O_1892,N_14986,N_14890);
nand UO_1893 (O_1893,N_14940,N_14914);
nor UO_1894 (O_1894,N_14804,N_14934);
nand UO_1895 (O_1895,N_14977,N_14912);
nand UO_1896 (O_1896,N_14949,N_14804);
nand UO_1897 (O_1897,N_14804,N_14993);
nor UO_1898 (O_1898,N_14954,N_14977);
or UO_1899 (O_1899,N_14994,N_14824);
or UO_1900 (O_1900,N_14834,N_14924);
or UO_1901 (O_1901,N_14821,N_14905);
nor UO_1902 (O_1902,N_14963,N_14895);
xor UO_1903 (O_1903,N_14992,N_14852);
xor UO_1904 (O_1904,N_14953,N_14816);
xor UO_1905 (O_1905,N_14859,N_14812);
xnor UO_1906 (O_1906,N_14877,N_14886);
and UO_1907 (O_1907,N_14867,N_14914);
nand UO_1908 (O_1908,N_14848,N_14847);
nor UO_1909 (O_1909,N_14922,N_14979);
nor UO_1910 (O_1910,N_14870,N_14875);
and UO_1911 (O_1911,N_14919,N_14901);
nor UO_1912 (O_1912,N_14974,N_14951);
nand UO_1913 (O_1913,N_14825,N_14894);
nor UO_1914 (O_1914,N_14956,N_14924);
nand UO_1915 (O_1915,N_14899,N_14914);
nor UO_1916 (O_1916,N_14883,N_14982);
nand UO_1917 (O_1917,N_14955,N_14964);
nand UO_1918 (O_1918,N_14822,N_14969);
or UO_1919 (O_1919,N_14812,N_14893);
xor UO_1920 (O_1920,N_14809,N_14902);
nor UO_1921 (O_1921,N_14994,N_14915);
nor UO_1922 (O_1922,N_14990,N_14881);
xor UO_1923 (O_1923,N_14923,N_14890);
and UO_1924 (O_1924,N_14985,N_14836);
or UO_1925 (O_1925,N_14943,N_14847);
or UO_1926 (O_1926,N_14852,N_14808);
and UO_1927 (O_1927,N_14911,N_14890);
nand UO_1928 (O_1928,N_14802,N_14800);
and UO_1929 (O_1929,N_14939,N_14895);
and UO_1930 (O_1930,N_14949,N_14900);
xnor UO_1931 (O_1931,N_14990,N_14812);
nor UO_1932 (O_1932,N_14908,N_14931);
nand UO_1933 (O_1933,N_14819,N_14931);
and UO_1934 (O_1934,N_14844,N_14812);
and UO_1935 (O_1935,N_14864,N_14922);
xnor UO_1936 (O_1936,N_14829,N_14914);
or UO_1937 (O_1937,N_14959,N_14863);
and UO_1938 (O_1938,N_14936,N_14962);
nor UO_1939 (O_1939,N_14899,N_14885);
nor UO_1940 (O_1940,N_14893,N_14981);
xnor UO_1941 (O_1941,N_14826,N_14996);
nor UO_1942 (O_1942,N_14912,N_14916);
xnor UO_1943 (O_1943,N_14830,N_14893);
or UO_1944 (O_1944,N_14981,N_14817);
xnor UO_1945 (O_1945,N_14959,N_14840);
xnor UO_1946 (O_1946,N_14810,N_14887);
and UO_1947 (O_1947,N_14967,N_14923);
and UO_1948 (O_1948,N_14974,N_14962);
and UO_1949 (O_1949,N_14870,N_14852);
nor UO_1950 (O_1950,N_14814,N_14803);
and UO_1951 (O_1951,N_14940,N_14978);
and UO_1952 (O_1952,N_14955,N_14957);
and UO_1953 (O_1953,N_14877,N_14976);
or UO_1954 (O_1954,N_14900,N_14897);
or UO_1955 (O_1955,N_14880,N_14887);
and UO_1956 (O_1956,N_14853,N_14831);
or UO_1957 (O_1957,N_14859,N_14935);
and UO_1958 (O_1958,N_14950,N_14988);
and UO_1959 (O_1959,N_14971,N_14983);
and UO_1960 (O_1960,N_14865,N_14870);
or UO_1961 (O_1961,N_14981,N_14832);
xor UO_1962 (O_1962,N_14933,N_14995);
or UO_1963 (O_1963,N_14955,N_14831);
nor UO_1964 (O_1964,N_14924,N_14857);
or UO_1965 (O_1965,N_14934,N_14901);
and UO_1966 (O_1966,N_14960,N_14924);
and UO_1967 (O_1967,N_14813,N_14924);
nor UO_1968 (O_1968,N_14926,N_14877);
xor UO_1969 (O_1969,N_14827,N_14907);
nand UO_1970 (O_1970,N_14905,N_14893);
or UO_1971 (O_1971,N_14927,N_14844);
xor UO_1972 (O_1972,N_14982,N_14818);
nor UO_1973 (O_1973,N_14864,N_14817);
and UO_1974 (O_1974,N_14857,N_14801);
nand UO_1975 (O_1975,N_14951,N_14802);
or UO_1976 (O_1976,N_14858,N_14933);
or UO_1977 (O_1977,N_14990,N_14966);
nor UO_1978 (O_1978,N_14833,N_14965);
xnor UO_1979 (O_1979,N_14827,N_14948);
and UO_1980 (O_1980,N_14884,N_14856);
xor UO_1981 (O_1981,N_14806,N_14874);
nand UO_1982 (O_1982,N_14850,N_14806);
nor UO_1983 (O_1983,N_14926,N_14900);
and UO_1984 (O_1984,N_14870,N_14933);
nor UO_1985 (O_1985,N_14918,N_14816);
or UO_1986 (O_1986,N_14939,N_14917);
or UO_1987 (O_1987,N_14819,N_14875);
and UO_1988 (O_1988,N_14964,N_14985);
and UO_1989 (O_1989,N_14810,N_14995);
nor UO_1990 (O_1990,N_14821,N_14944);
nand UO_1991 (O_1991,N_14951,N_14921);
nor UO_1992 (O_1992,N_14952,N_14954);
nor UO_1993 (O_1993,N_14915,N_14968);
or UO_1994 (O_1994,N_14894,N_14821);
or UO_1995 (O_1995,N_14830,N_14807);
or UO_1996 (O_1996,N_14803,N_14882);
or UO_1997 (O_1997,N_14906,N_14929);
xnor UO_1998 (O_1998,N_14834,N_14911);
nand UO_1999 (O_1999,N_14834,N_14877);
endmodule