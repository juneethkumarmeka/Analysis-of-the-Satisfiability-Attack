module basic_2000_20000_2500_4_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nor U0 (N_0,In_1289,In_226);
or U1 (N_1,In_411,In_1528);
and U2 (N_2,In_1630,In_1539);
nor U3 (N_3,In_720,In_298);
nor U4 (N_4,In_144,In_866);
or U5 (N_5,In_0,In_206);
and U6 (N_6,In_817,In_1298);
and U7 (N_7,In_1665,In_924);
and U8 (N_8,In_1522,In_1674);
xnor U9 (N_9,In_791,In_1594);
nor U10 (N_10,In_138,In_476);
xnor U11 (N_11,In_1913,In_1566);
or U12 (N_12,In_444,In_857);
xnor U13 (N_13,In_344,In_1580);
nor U14 (N_14,In_1670,In_1853);
nor U15 (N_15,In_67,In_1720);
and U16 (N_16,In_1965,In_1146);
nor U17 (N_17,In_1345,In_157);
xnor U18 (N_18,In_12,In_856);
nor U19 (N_19,In_1959,In_820);
nor U20 (N_20,In_1668,In_231);
nor U21 (N_21,In_597,In_164);
nor U22 (N_22,In_1824,In_1827);
nor U23 (N_23,In_1834,In_1467);
and U24 (N_24,In_1004,In_527);
or U25 (N_25,In_20,In_694);
xor U26 (N_26,In_1865,In_1535);
xnor U27 (N_27,In_1469,In_1125);
and U28 (N_28,In_1199,In_1214);
xnor U29 (N_29,In_279,In_288);
nand U30 (N_30,In_1031,In_1182);
xnor U31 (N_31,In_1129,In_859);
xor U32 (N_32,In_440,In_1860);
or U33 (N_33,In_1849,In_1902);
xor U34 (N_34,In_368,In_1758);
and U35 (N_35,In_1527,In_80);
xor U36 (N_36,In_271,In_1676);
or U37 (N_37,In_1634,In_168);
nand U38 (N_38,In_603,In_1615);
nand U39 (N_39,In_1940,In_1749);
nand U40 (N_40,In_618,In_1963);
xor U41 (N_41,In_1041,In_1568);
or U42 (N_42,In_256,In_222);
and U43 (N_43,In_1762,In_390);
xnor U44 (N_44,In_1974,In_1262);
xor U45 (N_45,In_1817,In_213);
nand U46 (N_46,In_1016,In_1867);
nand U47 (N_47,In_877,In_119);
nand U48 (N_48,In_1435,In_1459);
nor U49 (N_49,In_1699,In_1591);
or U50 (N_50,In_1662,In_1404);
and U51 (N_51,In_595,In_1037);
or U52 (N_52,In_1462,In_1126);
nand U53 (N_53,In_1000,In_1583);
or U54 (N_54,In_1702,In_1989);
nand U55 (N_55,In_386,In_742);
xor U56 (N_56,In_335,In_238);
xor U57 (N_57,In_683,In_1724);
and U58 (N_58,In_1056,In_1347);
nor U59 (N_59,In_1976,In_434);
nor U60 (N_60,In_1570,In_285);
nand U61 (N_61,In_1957,In_483);
or U62 (N_62,In_427,In_982);
xnor U63 (N_63,In_1838,In_1389);
nor U64 (N_64,In_1955,In_1585);
nand U65 (N_65,In_1365,In_718);
nor U66 (N_66,In_873,In_327);
xor U67 (N_67,In_248,In_738);
nor U68 (N_68,In_804,In_172);
and U69 (N_69,In_919,In_757);
and U70 (N_70,In_1076,In_1984);
and U71 (N_71,In_1780,In_1565);
xor U72 (N_72,In_1969,In_983);
or U73 (N_73,In_1240,In_489);
and U74 (N_74,In_428,In_659);
xnor U75 (N_75,In_346,In_1577);
nand U76 (N_76,In_140,In_38);
xor U77 (N_77,In_835,In_910);
nand U78 (N_78,In_1960,In_83);
nor U79 (N_79,In_1782,In_1966);
xor U80 (N_80,In_699,In_1332);
and U81 (N_81,In_837,In_648);
nor U82 (N_82,In_258,In_1313);
xnor U83 (N_83,In_1154,In_182);
nand U84 (N_84,In_980,In_14);
and U85 (N_85,In_568,In_1143);
nand U86 (N_86,In_1525,In_1465);
nand U87 (N_87,In_246,In_558);
and U88 (N_88,In_1318,In_51);
and U89 (N_89,In_1775,In_1480);
xor U90 (N_90,In_78,In_1430);
and U91 (N_91,In_240,In_1647);
or U92 (N_92,In_809,In_888);
nand U93 (N_93,In_446,In_740);
or U94 (N_94,In_633,In_1742);
and U95 (N_95,In_1048,In_579);
nor U96 (N_96,In_946,In_1491);
and U97 (N_97,In_548,In_1434);
or U98 (N_98,In_779,In_65);
xnor U99 (N_99,In_1152,In_1945);
or U100 (N_100,In_626,In_395);
and U101 (N_101,In_98,In_1600);
nor U102 (N_102,In_430,In_30);
nand U103 (N_103,In_281,In_725);
xnor U104 (N_104,In_1081,In_1850);
or U105 (N_105,In_829,In_135);
nor U106 (N_106,In_1296,In_1714);
and U107 (N_107,In_115,In_496);
nor U108 (N_108,In_825,In_1378);
nor U109 (N_109,In_1343,In_1516);
xnor U110 (N_110,In_1659,In_1169);
xnor U111 (N_111,In_33,In_559);
nor U112 (N_112,In_56,In_744);
or U113 (N_113,In_1291,In_7);
xor U114 (N_114,In_8,In_75);
or U115 (N_115,In_625,In_123);
or U116 (N_116,In_1401,In_1490);
xnor U117 (N_117,In_1983,In_761);
or U118 (N_118,In_1440,In_1320);
xor U119 (N_119,In_556,In_1202);
nand U120 (N_120,In_221,In_824);
and U121 (N_121,In_655,In_621);
nand U122 (N_122,In_19,In_1357);
and U123 (N_123,In_858,In_1299);
xnor U124 (N_124,In_1543,In_173);
nand U125 (N_125,In_1250,In_1903);
nand U126 (N_126,In_750,In_239);
xnor U127 (N_127,In_43,In_1086);
nor U128 (N_128,In_1641,In_1875);
nor U129 (N_129,In_1894,In_1830);
or U130 (N_130,In_861,In_723);
or U131 (N_131,In_1322,In_1718);
and U132 (N_132,In_1645,In_972);
xor U133 (N_133,In_1221,In_1682);
and U134 (N_134,In_1526,In_1941);
and U135 (N_135,In_1010,In_11);
or U136 (N_136,In_116,In_313);
nor U137 (N_137,In_1658,In_1093);
xnor U138 (N_138,In_21,In_810);
and U139 (N_139,In_249,In_117);
or U140 (N_140,In_87,In_1886);
xnor U141 (N_141,In_678,In_1579);
and U142 (N_142,In_1045,In_389);
and U143 (N_143,In_1334,In_673);
nand U144 (N_144,In_409,In_1964);
xor U145 (N_145,In_437,In_1495);
or U146 (N_146,In_1427,In_441);
nor U147 (N_147,In_355,In_1608);
xor U148 (N_148,In_1938,In_508);
and U149 (N_149,In_1800,In_1405);
and U150 (N_150,In_851,In_1596);
and U151 (N_151,In_730,In_696);
and U152 (N_152,In_475,In_1117);
or U153 (N_153,In_1962,In_1194);
and U154 (N_154,In_1071,In_1507);
xnor U155 (N_155,In_1703,In_1300);
nor U156 (N_156,In_964,In_406);
nor U157 (N_157,In_973,In_864);
xnor U158 (N_158,In_922,In_1090);
and U159 (N_159,In_917,In_1653);
nand U160 (N_160,In_846,In_867);
nand U161 (N_161,In_751,In_1277);
and U162 (N_162,In_1610,In_578);
or U163 (N_163,In_1673,In_1917);
nor U164 (N_164,In_665,In_773);
or U165 (N_165,In_736,In_1948);
and U166 (N_166,In_166,In_630);
nand U167 (N_167,In_515,In_1898);
or U168 (N_168,In_1359,In_216);
and U169 (N_169,In_177,In_789);
nand U170 (N_170,In_254,In_1926);
nor U171 (N_171,In_1951,In_1756);
nand U172 (N_172,In_686,In_628);
nand U173 (N_173,In_1191,In_901);
nor U174 (N_174,In_1342,In_848);
nand U175 (N_175,In_733,In_1141);
xnor U176 (N_176,In_379,In_1521);
xor U177 (N_177,In_1457,In_1773);
or U178 (N_178,In_1939,In_1801);
and U179 (N_179,In_860,In_844);
and U180 (N_180,In_1140,In_1746);
or U181 (N_181,In_1447,In_92);
nand U182 (N_182,In_1881,In_1196);
xnor U183 (N_183,In_1774,In_1757);
nand U184 (N_184,In_623,In_580);
nor U185 (N_185,In_1617,In_906);
and U186 (N_186,In_706,In_326);
xnor U187 (N_187,In_1413,In_612);
and U188 (N_188,In_1790,In_995);
nand U189 (N_189,In_1825,In_1449);
or U190 (N_190,In_654,In_698);
and U191 (N_191,In_870,In_1683);
xnor U192 (N_192,In_1590,In_933);
nor U193 (N_193,In_1063,In_1012);
nor U194 (N_194,In_1618,In_267);
nor U195 (N_195,In_1122,In_1421);
and U196 (N_196,In_494,In_1032);
or U197 (N_197,In_1576,In_1249);
and U198 (N_198,In_519,In_457);
or U199 (N_199,In_1377,In_885);
and U200 (N_200,In_1044,In_1123);
or U201 (N_201,In_445,In_1312);
xnor U202 (N_202,In_1292,In_1011);
or U203 (N_203,In_456,In_1935);
or U204 (N_204,In_1506,In_951);
and U205 (N_205,In_125,In_16);
and U206 (N_206,In_743,In_905);
xnor U207 (N_207,In_199,In_1017);
and U208 (N_208,In_598,In_1639);
nand U209 (N_209,In_265,In_1691);
and U210 (N_210,In_350,In_1943);
nor U211 (N_211,In_645,In_148);
and U212 (N_212,In_1584,In_304);
nand U213 (N_213,In_1247,In_937);
nand U214 (N_214,In_567,In_525);
and U215 (N_215,In_1918,In_377);
nand U216 (N_216,In_685,In_582);
nor U217 (N_217,In_721,In_1425);
and U218 (N_218,In_193,In_340);
nand U219 (N_219,In_63,In_419);
and U220 (N_220,In_55,In_1085);
xnor U221 (N_221,In_1680,In_22);
or U222 (N_222,In_1294,In_180);
nor U223 (N_223,In_1859,In_495);
or U224 (N_224,In_1787,In_1412);
nor U225 (N_225,In_322,In_1227);
and U226 (N_226,In_1233,In_1235);
xnor U227 (N_227,In_1632,In_328);
or U228 (N_228,In_1304,In_1986);
xor U229 (N_229,In_900,In_1253);
xnor U230 (N_230,In_42,In_786);
nor U231 (N_231,In_103,In_1609);
xor U232 (N_232,In_1133,In_975);
and U233 (N_233,In_40,In_1952);
or U234 (N_234,In_526,In_118);
nor U235 (N_235,In_590,In_1350);
or U236 (N_236,In_1733,In_1504);
nor U237 (N_237,In_94,In_473);
nor U238 (N_238,In_1878,In_514);
or U239 (N_239,In_478,In_537);
xor U240 (N_240,In_657,In_998);
xor U241 (N_241,In_1236,In_1667);
nand U242 (N_242,In_383,In_758);
and U243 (N_243,In_1264,In_1422);
nand U244 (N_244,In_879,In_1283);
or U245 (N_245,In_1772,In_703);
nand U246 (N_246,In_1643,In_155);
nand U247 (N_247,In_999,In_843);
xor U248 (N_248,In_1075,In_1372);
xnor U249 (N_249,In_588,In_1180);
xor U250 (N_250,In_1614,In_1338);
xnor U251 (N_251,In_324,In_1767);
or U252 (N_252,In_1319,In_968);
nor U253 (N_253,In_894,In_1700);
xor U254 (N_254,In_1669,In_109);
or U255 (N_255,In_245,In_1497);
xor U256 (N_256,In_1423,In_466);
nor U257 (N_257,In_503,In_1512);
and U258 (N_258,In_255,In_1722);
nand U259 (N_259,In_290,In_1464);
xnor U260 (N_260,In_1271,In_1181);
and U261 (N_261,In_192,In_1530);
and U262 (N_262,In_1324,In_981);
xor U263 (N_263,In_1567,In_566);
nand U264 (N_264,In_460,In_1050);
or U265 (N_265,In_1217,In_1198);
or U266 (N_266,In_1498,In_1764);
nor U267 (N_267,In_1042,In_371);
nor U268 (N_268,In_1348,In_287);
nor U269 (N_269,In_17,In_153);
or U270 (N_270,In_449,In_1248);
and U271 (N_271,In_1625,In_1686);
nor U272 (N_272,In_90,In_161);
nor U273 (N_273,In_638,In_957);
nand U274 (N_274,In_836,In_1145);
xor U275 (N_275,In_1376,In_302);
nor U276 (N_276,In_1893,In_1254);
and U277 (N_277,In_1173,In_1679);
xor U278 (N_278,In_1672,In_1390);
or U279 (N_279,In_251,In_1328);
and U280 (N_280,In_801,In_1367);
nand U281 (N_281,In_1361,In_1589);
xor U282 (N_282,In_1201,In_362);
or U283 (N_283,In_480,In_1139);
xnor U284 (N_284,In_978,In_1994);
and U285 (N_285,In_726,In_979);
nand U286 (N_286,In_930,In_993);
and U287 (N_287,In_450,In_112);
xor U288 (N_288,In_915,In_44);
nor U289 (N_289,In_1096,In_942);
or U290 (N_290,In_299,In_1315);
nand U291 (N_291,In_1097,In_724);
or U292 (N_292,In_1588,In_481);
nor U293 (N_293,In_1837,In_571);
and U294 (N_294,In_954,In_1057);
nor U295 (N_295,In_1207,In_1225);
xnor U296 (N_296,In_1744,In_1896);
or U297 (N_297,In_1545,In_1039);
or U298 (N_298,In_613,In_531);
and U299 (N_299,In_1740,In_1842);
nand U300 (N_300,In_1297,In_1794);
nand U301 (N_301,In_27,In_666);
or U302 (N_302,In_463,In_615);
and U303 (N_303,In_142,In_1078);
xor U304 (N_304,In_1985,In_762);
or U305 (N_305,In_1329,In_576);
nand U306 (N_306,In_1793,In_811);
nand U307 (N_307,In_1603,In_364);
nand U308 (N_308,In_1186,In_1748);
xnor U309 (N_309,In_339,In_1255);
nand U310 (N_310,In_622,In_181);
or U311 (N_311,In_1697,In_139);
nand U312 (N_312,In_1452,In_882);
xnor U313 (N_313,In_617,In_1677);
and U314 (N_314,In_1061,In_1923);
xor U315 (N_315,In_198,In_788);
nor U316 (N_316,In_1205,In_1038);
nor U317 (N_317,In_1455,In_374);
and U318 (N_318,In_1341,In_575);
nor U319 (N_319,In_640,In_672);
nand U320 (N_320,In_331,In_1754);
xnor U321 (N_321,In_93,In_1385);
and U322 (N_322,In_236,In_260);
and U323 (N_323,In_1408,In_1503);
nand U324 (N_324,In_1238,In_1845);
xor U325 (N_325,In_317,In_646);
nor U326 (N_326,In_1397,In_616);
nor U327 (N_327,In_701,In_841);
or U328 (N_328,In_544,In_128);
nor U329 (N_329,In_392,In_432);
xnor U330 (N_330,In_821,In_194);
or U331 (N_331,In_1765,In_822);
nor U332 (N_332,In_1021,In_491);
or U333 (N_333,In_1070,In_538);
or U334 (N_334,In_865,In_854);
and U335 (N_335,In_204,In_1534);
and U336 (N_336,In_32,In_1947);
or U337 (N_337,In_1106,In_1074);
xor U338 (N_338,In_547,In_1279);
and U339 (N_339,In_952,In_1396);
or U340 (N_340,In_420,In_1967);
nand U341 (N_341,In_436,In_1688);
nand U342 (N_342,In_372,In_1611);
xor U343 (N_343,In_827,In_1351);
nand U344 (N_344,In_1803,In_272);
and U345 (N_345,In_215,In_1177);
and U346 (N_346,In_1310,In_632);
nand U347 (N_347,In_29,In_1621);
or U348 (N_348,In_352,In_1587);
xor U349 (N_349,In_564,In_1442);
and U350 (N_350,In_295,In_716);
nor U351 (N_351,In_471,In_1922);
nand U352 (N_352,In_1147,In_1392);
xnor U353 (N_353,In_1415,In_874);
nand U354 (N_354,In_1899,In_818);
xor U355 (N_355,In_1987,In_1407);
and U356 (N_356,In_1119,In_1712);
nor U357 (N_357,In_405,In_1424);
nand U358 (N_358,In_1613,In_828);
and U359 (N_359,In_1114,In_1384);
xor U360 (N_360,In_1007,In_814);
nand U361 (N_361,In_513,In_1884);
nor U362 (N_362,In_777,In_842);
or U363 (N_363,In_1759,In_1747);
nand U364 (N_364,In_639,In_1906);
nand U365 (N_365,In_57,In_533);
or U366 (N_366,In_1436,In_1912);
xor U367 (N_367,In_675,In_967);
nand U368 (N_368,In_1655,In_1832);
xnor U369 (N_369,In_461,In_934);
or U370 (N_370,In_1726,In_212);
nand U371 (N_371,In_218,In_976);
nor U372 (N_372,In_1080,In_1159);
and U373 (N_373,In_1561,In_1520);
nand U374 (N_374,In_4,In_1373);
nor U375 (N_375,In_381,In_956);
and U376 (N_376,In_1308,In_1441);
or U377 (N_377,In_872,In_863);
and U378 (N_378,In_1946,In_1445);
xor U379 (N_379,In_1079,In_1598);
nand U380 (N_380,In_393,In_1992);
nor U381 (N_381,In_611,In_175);
and U382 (N_382,In_1224,In_1979);
xor U383 (N_383,In_689,In_482);
or U384 (N_384,In_1197,In_1393);
xor U385 (N_385,In_532,In_1137);
nor U386 (N_386,In_1226,In_439);
nor U387 (N_387,In_1750,In_1928);
or U388 (N_388,In_1820,In_1091);
nand U389 (N_389,In_219,In_1242);
xor U390 (N_390,In_1484,In_1326);
and U391 (N_391,In_282,In_969);
xor U392 (N_392,In_759,In_722);
xor U393 (N_393,In_876,In_1036);
or U394 (N_394,In_984,In_1810);
and U395 (N_395,In_1453,In_356);
xnor U396 (N_396,In_303,In_813);
xnor U397 (N_397,In_1931,In_1027);
nand U398 (N_398,In_243,In_1729);
or U399 (N_399,In_162,In_165);
or U400 (N_400,In_938,In_927);
nand U401 (N_401,In_768,In_120);
or U402 (N_402,In_708,In_262);
xnor U403 (N_403,In_1301,In_552);
and U404 (N_404,In_3,In_1921);
or U405 (N_405,In_1844,In_1494);
xor U406 (N_406,In_1822,In_619);
and U407 (N_407,In_1606,In_1175);
and U408 (N_408,In_1786,In_163);
and U409 (N_409,In_868,In_1161);
xor U410 (N_410,In_1371,In_1721);
and U411 (N_411,In_1446,In_755);
nand U412 (N_412,In_883,In_316);
and U413 (N_413,In_1745,In_634);
or U414 (N_414,In_1120,In_1950);
nor U415 (N_415,In_604,In_596);
nand U416 (N_416,In_96,In_1826);
and U417 (N_417,In_1261,In_1105);
xnor U418 (N_418,In_793,In_709);
nor U419 (N_419,In_375,In_932);
xor U420 (N_420,In_1666,In_1267);
nor U421 (N_421,In_1927,In_1956);
and U422 (N_422,In_944,In_1811);
and U423 (N_423,In_451,In_1164);
nor U424 (N_424,In_647,In_365);
xor U425 (N_425,In_985,In_940);
xnor U426 (N_426,In_502,In_18);
or U427 (N_427,In_929,In_1486);
or U428 (N_428,In_73,In_1211);
xnor U429 (N_429,In_1008,In_501);
nor U430 (N_430,In_1336,In_1709);
or U431 (N_431,In_1369,In_210);
nand U432 (N_432,In_230,In_1331);
or U433 (N_433,In_1508,In_792);
xor U434 (N_434,In_237,In_1458);
xor U435 (N_435,In_557,In_988);
nand U436 (N_436,In_417,In_1355);
nor U437 (N_437,In_1284,In_26);
xor U438 (N_438,In_1514,In_1174);
xnor U439 (N_439,In_1470,In_235);
nand U440 (N_440,In_289,In_284);
xor U441 (N_441,In_1185,In_1317);
nand U442 (N_442,In_908,In_643);
nor U443 (N_443,In_711,In_700);
xnor U444 (N_444,In_367,In_1382);
xnor U445 (N_445,In_1067,In_609);
nand U446 (N_446,In_1732,In_668);
and U447 (N_447,In_875,In_889);
xor U448 (N_448,In_1846,In_680);
nand U449 (N_449,In_1847,In_540);
or U450 (N_450,In_1633,In_431);
nand U451 (N_451,In_530,In_1409);
and U452 (N_452,In_1110,In_663);
and U453 (N_453,In_1562,In_1149);
or U454 (N_454,In_1478,In_1717);
xnor U455 (N_455,In_629,In_1907);
nand U456 (N_456,In_833,In_802);
nand U457 (N_457,In_948,In_1840);
nor U458 (N_458,In_61,In_1776);
xnor U459 (N_459,In_1339,In_1505);
nor U460 (N_460,In_1092,In_1560);
or U461 (N_461,In_1605,In_454);
nand U462 (N_462,In_1475,In_1874);
xor U463 (N_463,In_1542,In_130);
or U464 (N_464,In_562,In_418);
or U465 (N_465,In_220,In_1601);
nor U466 (N_466,In_1410,In_134);
xnor U467 (N_467,In_1022,In_987);
nand U468 (N_468,In_732,In_1306);
nor U469 (N_469,In_1961,In_1876);
xnor U470 (N_470,In_1942,In_704);
and U471 (N_471,In_1558,In_1072);
xor U472 (N_472,In_1635,In_516);
or U473 (N_473,In_196,In_297);
and U474 (N_474,In_806,In_382);
nor U475 (N_475,In_1996,In_1627);
xor U476 (N_476,In_1065,In_45);
nor U477 (N_477,In_1473,In_424);
nor U478 (N_478,In_34,In_563);
or U479 (N_479,In_561,In_171);
or U480 (N_480,In_426,In_1537);
and U481 (N_481,In_702,In_1132);
or U482 (N_482,In_1909,In_10);
nand U483 (N_483,In_385,In_1209);
and U484 (N_484,In_1461,In_150);
or U485 (N_485,In_1222,In_728);
xor U486 (N_486,In_765,In_1555);
and U487 (N_487,In_671,In_376);
xor U488 (N_488,In_1165,In_179);
xnor U489 (N_489,In_398,In_321);
and U490 (N_490,In_1841,In_485);
nand U491 (N_491,In_1115,In_1468);
and U492 (N_492,In_1930,In_1905);
nor U493 (N_493,In_69,In_234);
or U494 (N_494,In_545,In_1675);
xnor U495 (N_495,In_1089,In_1836);
or U496 (N_496,In_676,In_1231);
or U497 (N_497,In_209,In_136);
xnor U498 (N_498,In_25,In_1265);
nor U499 (N_499,In_1040,In_753);
or U500 (N_500,In_1855,In_624);
and U501 (N_501,In_1888,In_1064);
nor U502 (N_502,In_1519,In_1513);
nand U503 (N_503,In_347,In_1502);
xnor U504 (N_504,In_669,In_918);
and U505 (N_505,In_113,In_320);
and U506 (N_506,In_435,In_1919);
or U507 (N_507,In_453,In_366);
xnor U508 (N_508,In_584,In_1184);
nand U509 (N_509,In_1256,In_1171);
xor U510 (N_510,In_1597,In_357);
nor U511 (N_511,In_41,In_1575);
or U512 (N_512,In_23,In_1864);
xnor U513 (N_513,In_39,In_1274);
and U514 (N_514,In_183,In_1646);
or U515 (N_515,In_849,In_1599);
nor U516 (N_516,In_1536,In_920);
xor U517 (N_517,In_472,In_1971);
nor U518 (N_518,In_442,In_769);
nand U519 (N_519,In_715,In_276);
xnor U520 (N_520,In_1612,In_223);
xnor U521 (N_521,In_1901,In_586);
xnor U522 (N_522,In_1216,In_1548);
nand U523 (N_523,In_361,In_1541);
and U524 (N_524,In_400,In_707);
nand U525 (N_525,In_1783,In_528);
or U526 (N_526,In_1346,In_1770);
nor U527 (N_527,In_1309,In_1073);
and U528 (N_528,In_897,In_247);
and U529 (N_529,In_1472,In_1015);
nor U530 (N_530,In_553,In_1356);
nand U531 (N_531,In_1999,In_35);
nand U532 (N_532,In_1684,In_1135);
nor U533 (N_533,In_487,In_1370);
xnor U534 (N_534,In_631,In_845);
nand U535 (N_535,In_1915,In_132);
nor U536 (N_536,In_891,In_1381);
or U537 (N_537,In_794,In_1657);
nor U538 (N_538,In_1087,In_1690);
nand U539 (N_539,In_652,In_534);
nor U540 (N_540,In_1843,In_176);
nor U541 (N_541,In_644,In_959);
and U542 (N_542,In_767,In_1887);
xor U543 (N_543,In_1559,In_1725);
nor U544 (N_544,In_790,In_1908);
and U545 (N_545,In_1595,In_1788);
and U546 (N_546,In_1051,In_396);
and U547 (N_547,In_263,In_1344);
and U548 (N_548,In_577,In_1157);
and U549 (N_549,In_1949,In_1028);
nand U550 (N_550,In_587,In_1980);
xor U551 (N_551,In_600,In_971);
nand U552 (N_552,In_923,In_1387);
xor U553 (N_553,In_925,In_474);
nor U554 (N_554,In_1349,In_1431);
nand U555 (N_555,In_1880,In_48);
xor U556 (N_556,In_653,In_756);
nor U557 (N_557,In_1270,In_1795);
or U558 (N_558,In_1020,In_1807);
and U559 (N_559,In_966,In_1619);
nand U560 (N_560,In_661,In_1571);
nand U561 (N_561,In_1977,In_1815);
and U562 (N_562,In_913,In_1364);
nor U563 (N_563,In_111,In_1395);
and U564 (N_564,In_369,In_5);
xor U565 (N_565,In_286,In_641);
nand U566 (N_566,In_49,In_1206);
and U567 (N_567,In_573,In_550);
nand U568 (N_568,In_974,In_1998);
nand U569 (N_569,In_729,In_1698);
xnor U570 (N_570,In_31,In_1804);
and U571 (N_571,In_931,In_614);
xor U572 (N_572,In_1869,In_1035);
or U573 (N_573,In_1866,In_855);
xor U574 (N_574,In_1816,In_151);
xor U575 (N_575,In_105,In_705);
or U576 (N_576,In_748,In_1652);
nand U577 (N_577,In_852,In_250);
nand U578 (N_578,In_1550,In_735);
xnor U579 (N_579,In_1856,In_554);
nor U580 (N_580,In_1778,In_211);
and U581 (N_581,In_928,In_1481);
and U582 (N_582,In_1398,In_413);
and U583 (N_583,In_1258,In_752);
and U584 (N_584,In_710,In_1200);
nand U585 (N_585,In_1650,In_121);
and U586 (N_586,In_330,In_225);
xnor U587 (N_587,In_1743,In_1162);
nor U588 (N_588,In_1779,In_1572);
nor U589 (N_589,In_656,In_1981);
and U590 (N_590,In_1252,In_1671);
or U591 (N_591,In_884,In_325);
and U592 (N_592,In_1303,In_1552);
and U593 (N_593,In_880,In_1730);
nor U594 (N_594,In_1829,In_59);
nand U595 (N_595,In_737,In_1708);
nand U596 (N_596,In_493,In_781);
xnor U597 (N_597,In_1229,In_1379);
xnor U598 (N_598,In_1889,In_504);
xnor U599 (N_599,In_1190,In_1799);
nand U600 (N_600,In_1958,In_1230);
and U601 (N_601,In_1103,In_1433);
nor U602 (N_602,In_1604,In_687);
and U603 (N_603,In_1482,In_1187);
and U604 (N_604,In_1366,In_338);
xor U605 (N_605,In_315,In_214);
or U606 (N_606,In_1269,In_862);
and U607 (N_607,In_1544,In_149);
and U608 (N_608,In_823,In_1863);
nand U609 (N_609,In_359,In_143);
nor U610 (N_610,In_1978,In_1418);
nand U611 (N_611,In_1890,In_803);
xor U612 (N_612,In_1879,In_731);
xnor U613 (N_613,In_660,In_1789);
xnor U614 (N_614,In_84,In_1403);
or U615 (N_615,In_1664,In_1134);
or U616 (N_616,In_784,In_1399);
or U617 (N_617,In_1069,In_602);
xor U618 (N_618,In_1813,In_1131);
and U619 (N_619,In_749,In_1629);
nand U620 (N_620,In_1529,In_1100);
or U621 (N_621,In_1488,In_484);
nand U622 (N_622,In_1259,In_1239);
nor U623 (N_623,In_1553,In_348);
nand U624 (N_624,In_1066,In_943);
xnor U625 (N_625,In_1660,In_569);
xor U626 (N_626,In_1861,In_1932);
xnor U627 (N_627,In_912,In_847);
nand U628 (N_628,In_252,In_1654);
nor U629 (N_629,In_64,In_363);
and U630 (N_630,In_447,In_787);
nand U631 (N_631,In_1054,In_1777);
xor U632 (N_632,In_941,In_593);
nand U633 (N_633,In_1101,In_1735);
and U634 (N_634,In_591,In_543);
or U635 (N_635,In_1275,In_308);
and U636 (N_636,In_1213,In_950);
nand U637 (N_637,In_1972,In_1648);
or U638 (N_638,In_838,In_408);
xor U639 (N_639,In_620,In_1130);
and U640 (N_640,In_808,In_1644);
and U641 (N_641,In_273,In_1220);
or U642 (N_642,In_895,In_570);
or U643 (N_643,In_682,In_510);
nand U644 (N_644,In_869,In_1474);
and U645 (N_645,In_1479,In_300);
and U646 (N_646,In_423,In_1466);
nor U647 (N_647,In_380,In_1203);
and U648 (N_648,In_77,In_780);
nor U649 (N_649,In_904,In_1797);
nand U650 (N_650,In_1163,In_1781);
xnor U651 (N_651,In_1068,In_1593);
or U652 (N_652,In_154,In_191);
and U653 (N_653,In_775,In_1053);
or U654 (N_654,In_71,In_24);
and U655 (N_655,In_850,In_524);
nand U656 (N_656,In_1689,In_853);
or U657 (N_657,In_1538,In_970);
xnor U658 (N_658,In_1936,In_926);
xor U659 (N_659,In_1188,In_1739);
or U660 (N_660,In_1574,In_1483);
and U661 (N_661,In_1937,In_1707);
nor U662 (N_662,In_360,In_1245);
and U663 (N_663,In_195,In_812);
nand U664 (N_664,In_1681,In_1082);
nand U665 (N_665,In_1150,In_1183);
xor U666 (N_666,In_152,In_1193);
nand U667 (N_667,In_1819,In_517);
xnor U668 (N_668,In_1752,In_72);
nand U669 (N_669,In_1102,In_2);
xor U670 (N_670,In_443,In_91);
xnor U671 (N_671,In_697,In_1362);
xnor U672 (N_672,In_1451,In_291);
and U673 (N_673,In_253,In_1138);
xor U674 (N_674,In_1586,In_692);
nand U675 (N_675,In_1426,In_429);
xnor U676 (N_676,In_1892,In_54);
nor U677 (N_677,In_1713,In_1852);
xor U678 (N_678,In_1107,In_52);
nor U679 (N_679,In_81,In_890);
and U680 (N_680,In_921,In_1380);
and U681 (N_681,In_292,In_452);
nor U682 (N_682,In_1170,In_261);
nand U683 (N_683,In_1975,In_1034);
nor U684 (N_684,In_684,In_1112);
xnor U685 (N_685,In_1151,In_1511);
or U686 (N_686,In_1900,In_1215);
nand U687 (N_687,In_605,In_1833);
nand U688 (N_688,In_607,In_1168);
nor U689 (N_689,In_1563,In_310);
xor U690 (N_690,In_1127,In_1564);
nor U691 (N_691,In_509,In_965);
or U692 (N_692,In_264,In_1616);
or U693 (N_693,In_1523,In_1854);
xnor U694 (N_694,In_1710,In_770);
or U695 (N_695,In_469,In_782);
or U696 (N_696,In_283,In_1891);
nor U697 (N_697,In_785,In_512);
and U698 (N_698,In_124,In_244);
nor U699 (N_699,In_1995,In_1406);
nor U700 (N_700,In_881,In_500);
xnor U701 (N_701,In_1158,In_62);
nand U702 (N_702,In_1160,In_1116);
nand U703 (N_703,In_189,In_1546);
and U704 (N_704,In_312,In_1386);
or U705 (N_705,In_939,In_228);
or U706 (N_706,In_714,In_693);
or U707 (N_707,In_960,In_1383);
nand U708 (N_708,In_1701,In_462);
or U709 (N_709,In_896,In_394);
xor U710 (N_710,In_1013,In_333);
nor U711 (N_711,In_402,In_1047);
and U712 (N_712,In_9,In_1391);
and U713 (N_713,In_110,In_506);
or U714 (N_714,In_1411,In_898);
and U715 (N_715,In_1755,In_1327);
nor U716 (N_716,In_1305,In_601);
nand U717 (N_717,In_1153,In_100);
nand U718 (N_718,In_949,In_1109);
or U719 (N_719,In_1244,In_1280);
or U720 (N_720,In_412,In_1924);
or U721 (N_721,In_1,In_670);
nor U722 (N_722,In_1492,In_1084);
and U723 (N_723,In_1897,In_1736);
nor U724 (N_724,In_589,In_892);
xor U725 (N_725,In_871,In_1785);
or U726 (N_726,In_1933,In_1642);
or U727 (N_727,In_996,In_1263);
xor U728 (N_728,In_85,In_796);
xnor U729 (N_729,In_1241,In_296);
nand U730 (N_730,In_1678,In_169);
xor U731 (N_731,In_1095,In_127);
or U732 (N_732,In_774,In_47);
xnor U733 (N_733,In_1792,In_1210);
nand U734 (N_734,In_1791,In_1910);
or U735 (N_735,In_1456,In_958);
xnor U736 (N_736,In_373,In_1569);
and U737 (N_737,In_1839,In_1685);
nor U738 (N_738,In_1374,In_637);
nand U739 (N_739,In_266,In_887);
xor U740 (N_740,In_1195,In_1706);
and U741 (N_741,In_1970,In_1731);
or U742 (N_742,In_314,In_1622);
or U743 (N_743,In_1172,In_1204);
xor U744 (N_744,In_991,In_1805);
and U745 (N_745,In_1156,In_141);
nand U746 (N_746,In_1573,In_754);
and U747 (N_747,In_1741,In_1432);
nand U748 (N_748,In_1113,In_1273);
nand U749 (N_749,In_679,In_378);
nand U750 (N_750,In_1607,In_658);
nand U751 (N_751,In_1402,In_305);
nand U752 (N_752,In_1232,In_610);
xor U753 (N_753,In_1873,In_122);
or U754 (N_754,In_549,In_170);
or U755 (N_755,In_86,In_1499);
xor U756 (N_756,In_592,In_907);
nand U757 (N_757,In_911,In_13);
nor U758 (N_758,In_555,In_772);
and U759 (N_759,In_1394,In_798);
nand U760 (N_760,In_800,In_1476);
nand U761 (N_761,In_1851,In_1695);
nor U762 (N_762,In_492,In_370);
and U763 (N_763,In_1055,In_1796);
xor U764 (N_764,In_1419,In_74);
or U765 (N_765,In_1014,In_1524);
nand U766 (N_766,In_1868,In_1531);
and U767 (N_767,In_997,In_207);
nor U768 (N_768,In_421,In_1895);
xor U769 (N_769,In_1532,In_158);
xor U770 (N_770,In_520,In_1148);
or U771 (N_771,In_583,In_536);
nor U772 (N_772,In_15,In_323);
and U773 (N_773,In_886,In_511);
or U774 (N_774,In_1623,In_1862);
xnor U775 (N_775,In_1489,In_1753);
or U776 (N_776,In_203,In_760);
nor U777 (N_777,In_1460,In_1260);
nand U778 (N_778,In_415,In_899);
and U779 (N_779,In_187,In_1354);
nand U780 (N_780,In_1018,In_1223);
or U781 (N_781,In_1340,In_989);
or U782 (N_782,In_1993,In_1973);
xor U783 (N_783,In_159,In_224);
nor U784 (N_784,In_1167,In_903);
or U785 (N_785,In_1477,In_416);
and U786 (N_786,In_916,In_521);
or U787 (N_787,In_1118,In_307);
or U788 (N_788,In_1715,In_1052);
xor U789 (N_789,In_1437,In_763);
or U790 (N_790,In_28,In_594);
nor U791 (N_791,In_1321,In_1046);
nor U792 (N_792,In_1814,In_1293);
or U793 (N_793,In_349,In_425);
nor U794 (N_794,In_1696,In_1029);
and U795 (N_795,In_114,In_1771);
nor U796 (N_796,In_565,In_1818);
nor U797 (N_797,In_1798,In_499);
xor U798 (N_798,In_455,In_351);
nor U799 (N_799,In_145,In_1111);
and U800 (N_800,In_1178,In_274);
nand U801 (N_801,In_1953,In_994);
or U802 (N_802,In_961,In_397);
and U803 (N_803,In_1885,In_318);
nor U804 (N_804,In_257,In_1218);
nor U805 (N_805,In_53,In_1155);
and U806 (N_806,In_99,In_1212);
xor U807 (N_807,In_1192,In_358);
nand U808 (N_808,In_58,In_1719);
and U809 (N_809,In_160,In_830);
xnor U810 (N_810,In_1582,In_1023);
xor U811 (N_811,In_747,In_1448);
and U812 (N_812,In_797,In_1858);
xnor U813 (N_813,In_688,In_522);
or U814 (N_814,In_1638,In_200);
or U815 (N_815,In_97,In_1444);
nor U816 (N_816,In_497,In_336);
nand U817 (N_817,In_717,In_1663);
and U818 (N_818,In_197,In_1062);
nor U819 (N_819,In_1316,In_1551);
and U820 (N_820,In_201,In_1251);
or U821 (N_821,In_102,In_217);
nor U822 (N_822,In_1692,In_1266);
nand U823 (N_823,In_832,In_1420);
or U824 (N_824,In_1228,In_1030);
nor U825 (N_825,In_560,In_129);
or U826 (N_826,In_1920,In_1982);
nand U827 (N_827,In_1325,In_1661);
and U828 (N_828,In_178,In_1121);
nor U829 (N_829,In_690,In_1626);
nand U830 (N_830,In_909,In_208);
nand U831 (N_831,In_1761,In_1831);
and U832 (N_832,In_1485,In_1509);
nor U833 (N_833,In_147,In_1059);
xor U834 (N_834,In_795,In_1925);
xnor U835 (N_835,In_523,In_1904);
or U836 (N_836,In_1179,In_636);
xor U837 (N_837,In_1246,In_343);
xnor U838 (N_838,In_963,In_746);
or U839 (N_839,In_764,In_319);
nor U840 (N_840,In_190,In_778);
nand U841 (N_841,In_1694,In_667);
nand U842 (N_842,In_1911,In_1517);
xnor U843 (N_843,In_1003,In_280);
or U844 (N_844,In_345,In_1043);
nor U845 (N_845,In_1549,In_1916);
or U846 (N_846,In_414,In_1094);
and U847 (N_847,In_1823,In_1991);
xor U848 (N_848,In_1337,In_1723);
or U849 (N_849,In_805,In_677);
or U850 (N_850,In_1104,In_488);
and U851 (N_851,In_635,In_1234);
nand U852 (N_852,In_232,In_1352);
nor U853 (N_853,In_293,In_1002);
xnor U854 (N_854,In_1968,In_242);
and U855 (N_855,In_807,In_1438);
nand U856 (N_856,In_353,In_1636);
nand U857 (N_857,In_403,In_1997);
nand U858 (N_858,In_1006,In_301);
or U859 (N_859,In_1219,In_1734);
or U860 (N_860,In_95,In_771);
xor U861 (N_861,In_388,In_1278);
or U862 (N_862,In_188,In_106);
xnor U863 (N_863,In_1108,In_1768);
nand U864 (N_864,In_205,In_1716);
and U865 (N_865,In_404,In_518);
xnor U866 (N_866,In_337,In_88);
and U867 (N_867,In_834,In_1828);
and U868 (N_868,In_1687,In_185);
xnor U869 (N_869,In_1624,In_167);
or U870 (N_870,In_186,In_1314);
xor U871 (N_871,In_1540,In_229);
nand U872 (N_872,In_1019,In_1307);
xor U873 (N_873,In_1914,In_1812);
xor U874 (N_874,In_893,In_137);
or U875 (N_875,In_1295,In_1501);
nand U876 (N_876,In_1784,In_1281);
and U877 (N_877,In_642,In_464);
nor U878 (N_878,In_306,In_107);
and U879 (N_879,In_1429,In_986);
and U880 (N_880,In_1417,In_783);
nor U881 (N_881,In_1286,In_1060);
xor U882 (N_882,In_1290,In_1033);
and U883 (N_883,In_878,In_902);
xnor U884 (N_884,In_691,In_36);
and U885 (N_885,In_674,In_608);
nor U886 (N_886,In_840,In_1882);
or U887 (N_887,In_477,In_1360);
and U888 (N_888,In_1237,In_606);
and U889 (N_889,In_1176,In_574);
nand U890 (N_890,In_990,In_1848);
xnor U891 (N_891,In_50,In_1870);
or U892 (N_892,In_407,In_1288);
xor U893 (N_893,In_1124,In_1189);
or U894 (N_894,In_387,In_1450);
nor U895 (N_895,In_627,In_1809);
nand U896 (N_896,In_1988,In_936);
or U897 (N_897,In_233,In_410);
or U898 (N_898,In_294,In_278);
nor U899 (N_899,In_1443,In_1821);
nor U900 (N_900,In_37,In_551);
nand U901 (N_901,In_1705,In_66);
or U902 (N_902,In_341,In_1649);
nand U903 (N_903,In_1471,In_712);
and U904 (N_904,In_599,In_1428);
nor U905 (N_905,In_1704,In_1333);
xor U906 (N_906,In_1871,In_831);
nand U907 (N_907,In_1323,In_68);
xor U908 (N_908,In_1136,In_82);
and U909 (N_909,In_1276,In_719);
or U910 (N_910,In_467,In_1728);
and U911 (N_911,In_745,In_1857);
xor U912 (N_912,In_1557,In_1578);
or U913 (N_913,In_1077,In_354);
xor U914 (N_914,In_713,In_46);
or U915 (N_915,In_1416,In_1808);
nand U916 (N_916,In_1547,In_819);
and U917 (N_917,In_1208,In_1375);
and U918 (N_918,In_1620,In_776);
nand U919 (N_919,In_131,In_1368);
and U920 (N_920,In_174,In_1400);
or U921 (N_921,In_1058,In_1944);
nor U922 (N_922,In_1806,In_311);
nand U923 (N_923,In_935,In_479);
and U924 (N_924,In_1166,In_468);
nand U925 (N_925,In_1282,In_535);
nor U926 (N_926,In_1769,In_1802);
and U927 (N_927,In_1049,In_1496);
and U928 (N_928,In_1024,In_945);
xor U929 (N_929,In_727,In_470);
nor U930 (N_930,In_1088,In_465);
nand U931 (N_931,In_839,In_664);
nand U932 (N_932,In_1602,In_1388);
nor U933 (N_933,In_1099,In_104);
nor U934 (N_934,In_1353,In_1272);
or U935 (N_935,In_1243,In_184);
nor U936 (N_936,In_490,In_108);
nand U937 (N_937,In_259,In_650);
and U938 (N_938,In_1487,In_1518);
or U939 (N_939,In_741,In_539);
xor U940 (N_940,In_585,In_541);
and U941 (N_941,In_1500,In_422);
nor U942 (N_942,In_1711,In_6);
or U943 (N_943,In_651,In_241);
and U944 (N_944,In_1311,In_1656);
nand U945 (N_945,In_401,In_992);
nand U946 (N_946,In_1144,In_433);
and U947 (N_947,In_79,In_1693);
or U948 (N_948,In_695,In_1651);
nor U949 (N_949,In_268,In_438);
nor U950 (N_950,In_202,In_1727);
nand U951 (N_951,In_816,In_1737);
and U952 (N_952,In_1883,In_227);
nor U953 (N_953,In_156,In_384);
nand U954 (N_954,In_546,In_766);
nand U955 (N_955,In_815,In_1877);
nand U956 (N_956,In_572,In_1454);
nand U957 (N_957,In_1026,In_1358);
xor U958 (N_958,In_1142,In_1005);
nand U959 (N_959,In_101,In_1493);
or U960 (N_960,In_269,In_1009);
or U961 (N_961,In_1766,In_146);
xor U962 (N_962,In_458,In_1631);
nand U963 (N_963,In_89,In_1001);
and U964 (N_964,In_962,In_1025);
nor U965 (N_965,In_399,In_799);
or U966 (N_966,In_1533,In_1285);
nand U967 (N_967,In_1581,In_953);
or U968 (N_968,In_1098,In_332);
or U969 (N_969,In_739,In_681);
nand U970 (N_970,In_126,In_275);
nor U971 (N_971,In_529,In_826);
xor U972 (N_972,In_486,In_60);
or U973 (N_973,In_391,In_1929);
or U974 (N_974,In_1515,In_1556);
and U975 (N_975,In_734,In_1083);
xor U976 (N_976,In_1439,In_1738);
and U977 (N_977,In_1363,In_1510);
or U978 (N_978,In_581,In_498);
xnor U979 (N_979,In_329,In_1835);
nand U980 (N_980,In_505,In_914);
or U981 (N_981,In_309,In_1637);
nand U982 (N_982,In_1463,In_507);
nand U983 (N_983,In_1760,In_1414);
nand U984 (N_984,In_1302,In_277);
xnor U985 (N_985,In_662,In_1954);
nand U986 (N_986,In_977,In_70);
xor U987 (N_987,In_1268,In_1640);
or U988 (N_988,In_448,In_334);
nand U989 (N_989,In_459,In_1554);
xor U990 (N_990,In_76,In_1763);
and U991 (N_991,In_1628,In_1335);
xnor U992 (N_992,In_1934,In_133);
and U993 (N_993,In_1257,In_1330);
and U994 (N_994,In_542,In_955);
and U995 (N_995,In_342,In_1592);
or U996 (N_996,In_1872,In_1287);
nor U997 (N_997,In_947,In_270);
xnor U998 (N_998,In_649,In_1128);
xnor U999 (N_999,In_1990,In_1751);
nor U1000 (N_1000,In_1800,In_1434);
nor U1001 (N_1001,In_1015,In_226);
or U1002 (N_1002,In_563,In_1693);
or U1003 (N_1003,In_1739,In_1876);
nand U1004 (N_1004,In_1516,In_1159);
xnor U1005 (N_1005,In_1895,In_552);
xor U1006 (N_1006,In_597,In_1368);
and U1007 (N_1007,In_118,In_807);
nand U1008 (N_1008,In_787,In_1850);
nand U1009 (N_1009,In_1721,In_938);
and U1010 (N_1010,In_1766,In_1627);
nor U1011 (N_1011,In_1730,In_578);
and U1012 (N_1012,In_1797,In_781);
xor U1013 (N_1013,In_1102,In_58);
xnor U1014 (N_1014,In_1919,In_289);
and U1015 (N_1015,In_520,In_620);
nand U1016 (N_1016,In_393,In_1298);
nand U1017 (N_1017,In_715,In_317);
nand U1018 (N_1018,In_1058,In_1091);
and U1019 (N_1019,In_245,In_1505);
and U1020 (N_1020,In_1259,In_1310);
nand U1021 (N_1021,In_877,In_1542);
nand U1022 (N_1022,In_632,In_1595);
and U1023 (N_1023,In_1209,In_1754);
or U1024 (N_1024,In_542,In_49);
and U1025 (N_1025,In_298,In_178);
xnor U1026 (N_1026,In_7,In_434);
or U1027 (N_1027,In_214,In_703);
or U1028 (N_1028,In_1530,In_119);
nor U1029 (N_1029,In_539,In_1849);
xor U1030 (N_1030,In_276,In_1247);
and U1031 (N_1031,In_1853,In_17);
nand U1032 (N_1032,In_143,In_418);
nand U1033 (N_1033,In_185,In_578);
nand U1034 (N_1034,In_1819,In_1238);
or U1035 (N_1035,In_924,In_621);
xor U1036 (N_1036,In_77,In_392);
and U1037 (N_1037,In_1075,In_721);
or U1038 (N_1038,In_16,In_872);
or U1039 (N_1039,In_1204,In_1733);
or U1040 (N_1040,In_764,In_756);
nor U1041 (N_1041,In_728,In_659);
or U1042 (N_1042,In_485,In_503);
or U1043 (N_1043,In_1760,In_364);
and U1044 (N_1044,In_1264,In_978);
or U1045 (N_1045,In_524,In_887);
nand U1046 (N_1046,In_1807,In_9);
xnor U1047 (N_1047,In_1396,In_1345);
and U1048 (N_1048,In_246,In_946);
or U1049 (N_1049,In_152,In_1194);
xnor U1050 (N_1050,In_1362,In_466);
xor U1051 (N_1051,In_96,In_62);
and U1052 (N_1052,In_463,In_952);
or U1053 (N_1053,In_597,In_531);
and U1054 (N_1054,In_1829,In_849);
nor U1055 (N_1055,In_1020,In_1968);
xnor U1056 (N_1056,In_770,In_1809);
nand U1057 (N_1057,In_1015,In_643);
nand U1058 (N_1058,In_1139,In_1976);
nand U1059 (N_1059,In_580,In_275);
or U1060 (N_1060,In_415,In_361);
or U1061 (N_1061,In_1625,In_1137);
and U1062 (N_1062,In_775,In_1277);
nand U1063 (N_1063,In_167,In_761);
nand U1064 (N_1064,In_1518,In_1676);
or U1065 (N_1065,In_1824,In_145);
nand U1066 (N_1066,In_1867,In_1752);
xor U1067 (N_1067,In_693,In_1094);
nor U1068 (N_1068,In_585,In_362);
nor U1069 (N_1069,In_820,In_663);
xor U1070 (N_1070,In_1457,In_162);
nor U1071 (N_1071,In_1341,In_1256);
and U1072 (N_1072,In_469,In_1830);
nor U1073 (N_1073,In_234,In_463);
xnor U1074 (N_1074,In_1095,In_320);
or U1075 (N_1075,In_762,In_1005);
xor U1076 (N_1076,In_311,In_410);
nor U1077 (N_1077,In_627,In_1259);
nand U1078 (N_1078,In_1499,In_1765);
and U1079 (N_1079,In_572,In_598);
nor U1080 (N_1080,In_825,In_1628);
xnor U1081 (N_1081,In_1778,In_1873);
nor U1082 (N_1082,In_4,In_1925);
and U1083 (N_1083,In_1177,In_1362);
nor U1084 (N_1084,In_1882,In_1228);
and U1085 (N_1085,In_1488,In_1050);
xor U1086 (N_1086,In_1774,In_70);
or U1087 (N_1087,In_269,In_905);
and U1088 (N_1088,In_1362,In_292);
nor U1089 (N_1089,In_903,In_650);
nand U1090 (N_1090,In_164,In_337);
or U1091 (N_1091,In_1844,In_97);
and U1092 (N_1092,In_391,In_1870);
nor U1093 (N_1093,In_937,In_1266);
nor U1094 (N_1094,In_1471,In_1684);
nor U1095 (N_1095,In_1272,In_405);
or U1096 (N_1096,In_261,In_34);
or U1097 (N_1097,In_1438,In_1966);
nand U1098 (N_1098,In_949,In_500);
xnor U1099 (N_1099,In_538,In_1798);
and U1100 (N_1100,In_1058,In_1513);
and U1101 (N_1101,In_1365,In_1081);
and U1102 (N_1102,In_242,In_969);
nor U1103 (N_1103,In_1328,In_1285);
or U1104 (N_1104,In_1840,In_1260);
nand U1105 (N_1105,In_1698,In_255);
xnor U1106 (N_1106,In_536,In_710);
xor U1107 (N_1107,In_1043,In_498);
and U1108 (N_1108,In_176,In_1821);
nand U1109 (N_1109,In_584,In_1233);
and U1110 (N_1110,In_902,In_35);
nand U1111 (N_1111,In_450,In_429);
nor U1112 (N_1112,In_325,In_1490);
or U1113 (N_1113,In_262,In_498);
or U1114 (N_1114,In_1677,In_1273);
xor U1115 (N_1115,In_939,In_399);
nor U1116 (N_1116,In_699,In_1155);
nand U1117 (N_1117,In_355,In_1670);
nor U1118 (N_1118,In_301,In_899);
nor U1119 (N_1119,In_1796,In_443);
nor U1120 (N_1120,In_1342,In_1327);
nor U1121 (N_1121,In_1312,In_202);
xor U1122 (N_1122,In_31,In_1764);
or U1123 (N_1123,In_1652,In_982);
and U1124 (N_1124,In_842,In_341);
nor U1125 (N_1125,In_466,In_856);
and U1126 (N_1126,In_325,In_1929);
or U1127 (N_1127,In_1639,In_18);
xnor U1128 (N_1128,In_1444,In_1559);
nor U1129 (N_1129,In_736,In_805);
xnor U1130 (N_1130,In_1113,In_1542);
or U1131 (N_1131,In_1271,In_1086);
nand U1132 (N_1132,In_1671,In_1121);
nor U1133 (N_1133,In_167,In_911);
nand U1134 (N_1134,In_896,In_751);
xnor U1135 (N_1135,In_1046,In_1387);
nand U1136 (N_1136,In_1025,In_1382);
nor U1137 (N_1137,In_74,In_1409);
nand U1138 (N_1138,In_1220,In_195);
nand U1139 (N_1139,In_17,In_457);
and U1140 (N_1140,In_738,In_515);
nor U1141 (N_1141,In_126,In_1675);
nand U1142 (N_1142,In_1823,In_1812);
xor U1143 (N_1143,In_1907,In_76);
and U1144 (N_1144,In_1220,In_1896);
and U1145 (N_1145,In_1383,In_1703);
xnor U1146 (N_1146,In_1605,In_1494);
or U1147 (N_1147,In_1136,In_1119);
or U1148 (N_1148,In_1071,In_127);
nand U1149 (N_1149,In_59,In_1413);
and U1150 (N_1150,In_746,In_38);
nand U1151 (N_1151,In_566,In_1068);
xnor U1152 (N_1152,In_1740,In_1405);
nor U1153 (N_1153,In_853,In_1875);
nor U1154 (N_1154,In_637,In_1801);
or U1155 (N_1155,In_1632,In_217);
nand U1156 (N_1156,In_149,In_275);
nand U1157 (N_1157,In_313,In_888);
or U1158 (N_1158,In_982,In_149);
xnor U1159 (N_1159,In_3,In_510);
nor U1160 (N_1160,In_989,In_712);
and U1161 (N_1161,In_453,In_438);
and U1162 (N_1162,In_1015,In_1177);
and U1163 (N_1163,In_1639,In_1216);
and U1164 (N_1164,In_878,In_111);
nor U1165 (N_1165,In_558,In_1114);
xor U1166 (N_1166,In_664,In_1665);
nor U1167 (N_1167,In_1307,In_1556);
nand U1168 (N_1168,In_538,In_1491);
nand U1169 (N_1169,In_1250,In_640);
and U1170 (N_1170,In_498,In_767);
or U1171 (N_1171,In_1749,In_401);
nor U1172 (N_1172,In_1172,In_79);
or U1173 (N_1173,In_1342,In_920);
or U1174 (N_1174,In_681,In_466);
xor U1175 (N_1175,In_1317,In_1488);
xnor U1176 (N_1176,In_594,In_534);
and U1177 (N_1177,In_1812,In_546);
and U1178 (N_1178,In_809,In_1683);
and U1179 (N_1179,In_124,In_656);
xor U1180 (N_1180,In_621,In_723);
or U1181 (N_1181,In_1419,In_1788);
nand U1182 (N_1182,In_1512,In_751);
xnor U1183 (N_1183,In_1117,In_1787);
nand U1184 (N_1184,In_438,In_1767);
or U1185 (N_1185,In_1028,In_1761);
nand U1186 (N_1186,In_365,In_881);
or U1187 (N_1187,In_1129,In_1074);
xnor U1188 (N_1188,In_1465,In_1225);
xnor U1189 (N_1189,In_1328,In_1127);
nand U1190 (N_1190,In_1329,In_200);
nor U1191 (N_1191,In_1722,In_315);
nand U1192 (N_1192,In_299,In_1448);
or U1193 (N_1193,In_1789,In_51);
nand U1194 (N_1194,In_1848,In_823);
xor U1195 (N_1195,In_10,In_777);
or U1196 (N_1196,In_1313,In_685);
and U1197 (N_1197,In_1816,In_317);
or U1198 (N_1198,In_1339,In_955);
nor U1199 (N_1199,In_1616,In_1960);
or U1200 (N_1200,In_1960,In_61);
or U1201 (N_1201,In_1247,In_1814);
or U1202 (N_1202,In_1137,In_17);
and U1203 (N_1203,In_1428,In_35);
xnor U1204 (N_1204,In_1367,In_631);
or U1205 (N_1205,In_467,In_1025);
nor U1206 (N_1206,In_71,In_1311);
nand U1207 (N_1207,In_1587,In_793);
xor U1208 (N_1208,In_1155,In_1266);
xor U1209 (N_1209,In_1629,In_830);
and U1210 (N_1210,In_897,In_452);
or U1211 (N_1211,In_1490,In_566);
nand U1212 (N_1212,In_890,In_808);
or U1213 (N_1213,In_629,In_929);
and U1214 (N_1214,In_789,In_1706);
and U1215 (N_1215,In_1570,In_1581);
nand U1216 (N_1216,In_1020,In_530);
xnor U1217 (N_1217,In_1405,In_1052);
xnor U1218 (N_1218,In_1732,In_1596);
or U1219 (N_1219,In_1752,In_1983);
nand U1220 (N_1220,In_248,In_1990);
nand U1221 (N_1221,In_188,In_164);
xor U1222 (N_1222,In_1681,In_583);
nor U1223 (N_1223,In_1654,In_1666);
nor U1224 (N_1224,In_1524,In_424);
xor U1225 (N_1225,In_607,In_84);
or U1226 (N_1226,In_1304,In_331);
or U1227 (N_1227,In_1000,In_1832);
nor U1228 (N_1228,In_1161,In_1155);
nor U1229 (N_1229,In_412,In_275);
or U1230 (N_1230,In_1271,In_886);
or U1231 (N_1231,In_1144,In_494);
and U1232 (N_1232,In_123,In_442);
or U1233 (N_1233,In_1683,In_947);
xor U1234 (N_1234,In_1555,In_1241);
nor U1235 (N_1235,In_1348,In_401);
xnor U1236 (N_1236,In_906,In_1900);
xor U1237 (N_1237,In_1928,In_169);
xor U1238 (N_1238,In_927,In_261);
nor U1239 (N_1239,In_1660,In_307);
xnor U1240 (N_1240,In_1357,In_1369);
xnor U1241 (N_1241,In_1110,In_1151);
and U1242 (N_1242,In_326,In_43);
or U1243 (N_1243,In_783,In_1907);
xnor U1244 (N_1244,In_1203,In_813);
nor U1245 (N_1245,In_527,In_1069);
and U1246 (N_1246,In_315,In_492);
xor U1247 (N_1247,In_477,In_537);
or U1248 (N_1248,In_1175,In_1170);
xnor U1249 (N_1249,In_1267,In_1599);
xor U1250 (N_1250,In_932,In_1633);
or U1251 (N_1251,In_287,In_658);
or U1252 (N_1252,In_991,In_1132);
xnor U1253 (N_1253,In_935,In_1216);
and U1254 (N_1254,In_106,In_973);
or U1255 (N_1255,In_1957,In_1477);
nand U1256 (N_1256,In_152,In_262);
xor U1257 (N_1257,In_61,In_1310);
nand U1258 (N_1258,In_1411,In_1708);
nand U1259 (N_1259,In_579,In_1457);
nor U1260 (N_1260,In_332,In_1705);
nand U1261 (N_1261,In_1587,In_117);
nor U1262 (N_1262,In_1003,In_1386);
xnor U1263 (N_1263,In_1418,In_73);
nor U1264 (N_1264,In_1960,In_1819);
and U1265 (N_1265,In_423,In_224);
xnor U1266 (N_1266,In_1716,In_369);
and U1267 (N_1267,In_438,In_1209);
or U1268 (N_1268,In_1830,In_1757);
and U1269 (N_1269,In_1162,In_1494);
nor U1270 (N_1270,In_343,In_1020);
nor U1271 (N_1271,In_1157,In_235);
nand U1272 (N_1272,In_1313,In_1218);
and U1273 (N_1273,In_185,In_520);
nor U1274 (N_1274,In_1403,In_1136);
and U1275 (N_1275,In_1681,In_1099);
nand U1276 (N_1276,In_1526,In_564);
nand U1277 (N_1277,In_698,In_1508);
nor U1278 (N_1278,In_63,In_560);
xnor U1279 (N_1279,In_1125,In_633);
or U1280 (N_1280,In_1233,In_467);
xor U1281 (N_1281,In_1736,In_1561);
nor U1282 (N_1282,In_857,In_1920);
nand U1283 (N_1283,In_1669,In_1318);
nand U1284 (N_1284,In_933,In_1938);
or U1285 (N_1285,In_1047,In_1827);
xor U1286 (N_1286,In_750,In_307);
or U1287 (N_1287,In_1882,In_97);
nand U1288 (N_1288,In_1627,In_634);
and U1289 (N_1289,In_211,In_1221);
and U1290 (N_1290,In_266,In_212);
xnor U1291 (N_1291,In_174,In_1835);
nand U1292 (N_1292,In_853,In_1199);
nand U1293 (N_1293,In_504,In_561);
nand U1294 (N_1294,In_1421,In_1881);
or U1295 (N_1295,In_1222,In_422);
and U1296 (N_1296,In_377,In_1572);
nor U1297 (N_1297,In_1733,In_308);
nor U1298 (N_1298,In_1814,In_599);
nor U1299 (N_1299,In_1939,In_905);
or U1300 (N_1300,In_1383,In_585);
xnor U1301 (N_1301,In_509,In_1112);
nor U1302 (N_1302,In_14,In_1211);
nor U1303 (N_1303,In_745,In_716);
or U1304 (N_1304,In_1371,In_1628);
or U1305 (N_1305,In_1502,In_237);
or U1306 (N_1306,In_582,In_349);
nand U1307 (N_1307,In_1378,In_522);
nor U1308 (N_1308,In_1448,In_1282);
or U1309 (N_1309,In_986,In_1616);
or U1310 (N_1310,In_28,In_450);
xor U1311 (N_1311,In_1799,In_170);
nand U1312 (N_1312,In_295,In_462);
nand U1313 (N_1313,In_222,In_1219);
or U1314 (N_1314,In_506,In_1011);
nor U1315 (N_1315,In_850,In_1499);
and U1316 (N_1316,In_303,In_1960);
xor U1317 (N_1317,In_258,In_517);
xor U1318 (N_1318,In_684,In_542);
or U1319 (N_1319,In_424,In_1692);
nand U1320 (N_1320,In_919,In_1964);
and U1321 (N_1321,In_475,In_1018);
and U1322 (N_1322,In_1332,In_380);
xor U1323 (N_1323,In_1561,In_750);
xnor U1324 (N_1324,In_544,In_193);
nand U1325 (N_1325,In_844,In_1381);
nor U1326 (N_1326,In_574,In_359);
nand U1327 (N_1327,In_1560,In_1018);
nand U1328 (N_1328,In_1365,In_1854);
nand U1329 (N_1329,In_1618,In_1661);
or U1330 (N_1330,In_624,In_1421);
and U1331 (N_1331,In_1971,In_1397);
and U1332 (N_1332,In_601,In_1324);
or U1333 (N_1333,In_1025,In_1437);
nand U1334 (N_1334,In_1835,In_1205);
xnor U1335 (N_1335,In_645,In_1293);
nand U1336 (N_1336,In_597,In_1742);
nor U1337 (N_1337,In_158,In_959);
and U1338 (N_1338,In_1001,In_1557);
nand U1339 (N_1339,In_439,In_337);
or U1340 (N_1340,In_1086,In_1741);
nor U1341 (N_1341,In_1410,In_1351);
nor U1342 (N_1342,In_1171,In_1838);
or U1343 (N_1343,In_1529,In_1199);
and U1344 (N_1344,In_1386,In_544);
and U1345 (N_1345,In_1409,In_135);
xnor U1346 (N_1346,In_1696,In_1170);
xnor U1347 (N_1347,In_1587,In_1240);
and U1348 (N_1348,In_677,In_834);
nand U1349 (N_1349,In_881,In_1560);
nor U1350 (N_1350,In_288,In_421);
nand U1351 (N_1351,In_1616,In_646);
and U1352 (N_1352,In_362,In_1910);
nand U1353 (N_1353,In_430,In_848);
xnor U1354 (N_1354,In_1086,In_525);
and U1355 (N_1355,In_1145,In_697);
nor U1356 (N_1356,In_492,In_1487);
nor U1357 (N_1357,In_1112,In_1144);
nor U1358 (N_1358,In_163,In_445);
or U1359 (N_1359,In_1106,In_1000);
nor U1360 (N_1360,In_1548,In_649);
nand U1361 (N_1361,In_85,In_467);
xnor U1362 (N_1362,In_1692,In_1930);
xnor U1363 (N_1363,In_472,In_1514);
and U1364 (N_1364,In_1132,In_1305);
xnor U1365 (N_1365,In_1448,In_1477);
and U1366 (N_1366,In_675,In_1533);
nand U1367 (N_1367,In_1004,In_1492);
or U1368 (N_1368,In_1857,In_407);
nand U1369 (N_1369,In_354,In_43);
nand U1370 (N_1370,In_923,In_1088);
nand U1371 (N_1371,In_918,In_383);
xor U1372 (N_1372,In_597,In_889);
and U1373 (N_1373,In_901,In_1451);
nand U1374 (N_1374,In_246,In_949);
and U1375 (N_1375,In_1366,In_414);
and U1376 (N_1376,In_812,In_694);
xnor U1377 (N_1377,In_1372,In_1901);
and U1378 (N_1378,In_507,In_714);
or U1379 (N_1379,In_1161,In_1194);
xnor U1380 (N_1380,In_3,In_694);
nor U1381 (N_1381,In_1274,In_831);
and U1382 (N_1382,In_556,In_1771);
nor U1383 (N_1383,In_858,In_1573);
nand U1384 (N_1384,In_444,In_1834);
nand U1385 (N_1385,In_1073,In_1308);
and U1386 (N_1386,In_517,In_1064);
xor U1387 (N_1387,In_1417,In_1282);
or U1388 (N_1388,In_1828,In_853);
xor U1389 (N_1389,In_1316,In_23);
nand U1390 (N_1390,In_1725,In_1967);
nand U1391 (N_1391,In_259,In_1487);
nand U1392 (N_1392,In_1085,In_250);
or U1393 (N_1393,In_1958,In_168);
nor U1394 (N_1394,In_1883,In_946);
nand U1395 (N_1395,In_1629,In_1519);
nor U1396 (N_1396,In_549,In_1279);
or U1397 (N_1397,In_1539,In_872);
nor U1398 (N_1398,In_1984,In_100);
and U1399 (N_1399,In_1583,In_1285);
nor U1400 (N_1400,In_1240,In_377);
xnor U1401 (N_1401,In_1367,In_334);
and U1402 (N_1402,In_1642,In_651);
or U1403 (N_1403,In_1331,In_1503);
nand U1404 (N_1404,In_1363,In_353);
or U1405 (N_1405,In_1107,In_687);
and U1406 (N_1406,In_485,In_1896);
or U1407 (N_1407,In_440,In_1418);
or U1408 (N_1408,In_403,In_1299);
nor U1409 (N_1409,In_1694,In_1936);
nand U1410 (N_1410,In_1256,In_103);
xnor U1411 (N_1411,In_881,In_134);
nor U1412 (N_1412,In_161,In_1346);
nor U1413 (N_1413,In_415,In_1121);
xor U1414 (N_1414,In_487,In_784);
nor U1415 (N_1415,In_355,In_1079);
or U1416 (N_1416,In_173,In_227);
nand U1417 (N_1417,In_1133,In_1880);
nor U1418 (N_1418,In_195,In_1954);
xnor U1419 (N_1419,In_1603,In_822);
xnor U1420 (N_1420,In_907,In_416);
and U1421 (N_1421,In_1340,In_1070);
and U1422 (N_1422,In_49,In_955);
nand U1423 (N_1423,In_874,In_1553);
nand U1424 (N_1424,In_87,In_1314);
and U1425 (N_1425,In_113,In_208);
nand U1426 (N_1426,In_1611,In_578);
and U1427 (N_1427,In_525,In_551);
nand U1428 (N_1428,In_0,In_1217);
or U1429 (N_1429,In_576,In_1070);
or U1430 (N_1430,In_1341,In_90);
and U1431 (N_1431,In_61,In_653);
nor U1432 (N_1432,In_1374,In_997);
or U1433 (N_1433,In_650,In_1562);
nand U1434 (N_1434,In_538,In_1080);
nor U1435 (N_1435,In_1405,In_595);
nand U1436 (N_1436,In_1172,In_666);
or U1437 (N_1437,In_818,In_833);
xnor U1438 (N_1438,In_1593,In_945);
and U1439 (N_1439,In_1924,In_931);
nand U1440 (N_1440,In_1650,In_582);
or U1441 (N_1441,In_1873,In_1082);
nor U1442 (N_1442,In_141,In_1410);
nand U1443 (N_1443,In_238,In_1464);
and U1444 (N_1444,In_78,In_1152);
nor U1445 (N_1445,In_1973,In_1752);
nor U1446 (N_1446,In_1189,In_1243);
and U1447 (N_1447,In_1050,In_1595);
or U1448 (N_1448,In_862,In_1761);
and U1449 (N_1449,In_557,In_1033);
nor U1450 (N_1450,In_1824,In_1515);
nand U1451 (N_1451,In_521,In_1674);
and U1452 (N_1452,In_1852,In_127);
xnor U1453 (N_1453,In_816,In_1205);
nand U1454 (N_1454,In_1358,In_875);
or U1455 (N_1455,In_1452,In_599);
nor U1456 (N_1456,In_934,In_1594);
or U1457 (N_1457,In_1327,In_300);
xnor U1458 (N_1458,In_66,In_53);
nor U1459 (N_1459,In_1634,In_449);
xnor U1460 (N_1460,In_1803,In_812);
xor U1461 (N_1461,In_245,In_1971);
and U1462 (N_1462,In_210,In_183);
or U1463 (N_1463,In_991,In_632);
xnor U1464 (N_1464,In_241,In_1046);
nor U1465 (N_1465,In_1880,In_1174);
nor U1466 (N_1466,In_808,In_1283);
or U1467 (N_1467,In_1154,In_1951);
xnor U1468 (N_1468,In_1112,In_2);
and U1469 (N_1469,In_700,In_1933);
nor U1470 (N_1470,In_1853,In_1647);
nand U1471 (N_1471,In_652,In_1216);
or U1472 (N_1472,In_1375,In_1800);
nand U1473 (N_1473,In_745,In_1899);
nor U1474 (N_1474,In_956,In_978);
nor U1475 (N_1475,In_1858,In_323);
nor U1476 (N_1476,In_887,In_114);
nor U1477 (N_1477,In_1655,In_541);
or U1478 (N_1478,In_1700,In_769);
nand U1479 (N_1479,In_892,In_1214);
nand U1480 (N_1480,In_1402,In_1627);
nand U1481 (N_1481,In_1504,In_42);
nor U1482 (N_1482,In_1032,In_748);
xor U1483 (N_1483,In_1001,In_72);
xor U1484 (N_1484,In_1889,In_490);
xor U1485 (N_1485,In_875,In_1425);
nand U1486 (N_1486,In_136,In_1733);
or U1487 (N_1487,In_902,In_793);
or U1488 (N_1488,In_1307,In_588);
and U1489 (N_1489,In_1825,In_1913);
and U1490 (N_1490,In_1443,In_1765);
nand U1491 (N_1491,In_1855,In_1327);
nor U1492 (N_1492,In_1549,In_288);
nor U1493 (N_1493,In_1327,In_1144);
or U1494 (N_1494,In_1198,In_1730);
nor U1495 (N_1495,In_439,In_1849);
nand U1496 (N_1496,In_1855,In_1372);
nor U1497 (N_1497,In_1745,In_1482);
or U1498 (N_1498,In_409,In_1639);
xor U1499 (N_1499,In_217,In_889);
nand U1500 (N_1500,In_1832,In_145);
or U1501 (N_1501,In_1435,In_1767);
xor U1502 (N_1502,In_286,In_281);
xor U1503 (N_1503,In_54,In_5);
nor U1504 (N_1504,In_1677,In_449);
or U1505 (N_1505,In_1748,In_1841);
nand U1506 (N_1506,In_15,In_1140);
or U1507 (N_1507,In_1337,In_838);
and U1508 (N_1508,In_1732,In_1117);
and U1509 (N_1509,In_495,In_382);
xor U1510 (N_1510,In_315,In_1302);
xor U1511 (N_1511,In_935,In_1607);
and U1512 (N_1512,In_875,In_1157);
nor U1513 (N_1513,In_1609,In_1024);
or U1514 (N_1514,In_344,In_1638);
xnor U1515 (N_1515,In_281,In_1132);
and U1516 (N_1516,In_1805,In_1208);
and U1517 (N_1517,In_1357,In_677);
nand U1518 (N_1518,In_567,In_1768);
or U1519 (N_1519,In_1800,In_1998);
and U1520 (N_1520,In_91,In_1831);
xnor U1521 (N_1521,In_1874,In_1157);
xnor U1522 (N_1522,In_1601,In_1127);
or U1523 (N_1523,In_506,In_896);
nor U1524 (N_1524,In_185,In_312);
and U1525 (N_1525,In_868,In_1127);
nor U1526 (N_1526,In_1142,In_709);
and U1527 (N_1527,In_1528,In_193);
or U1528 (N_1528,In_1495,In_854);
or U1529 (N_1529,In_868,In_1290);
xor U1530 (N_1530,In_300,In_555);
nor U1531 (N_1531,In_1828,In_870);
and U1532 (N_1532,In_2,In_437);
nor U1533 (N_1533,In_1686,In_309);
nor U1534 (N_1534,In_276,In_1204);
or U1535 (N_1535,In_758,In_1878);
nand U1536 (N_1536,In_1776,In_943);
xnor U1537 (N_1537,In_1628,In_229);
nand U1538 (N_1538,In_358,In_779);
and U1539 (N_1539,In_427,In_1863);
nand U1540 (N_1540,In_122,In_1778);
and U1541 (N_1541,In_79,In_17);
or U1542 (N_1542,In_542,In_1129);
and U1543 (N_1543,In_63,In_1047);
or U1544 (N_1544,In_1506,In_828);
and U1545 (N_1545,In_1250,In_1682);
and U1546 (N_1546,In_350,In_1313);
nand U1547 (N_1547,In_1525,In_112);
and U1548 (N_1548,In_1668,In_1823);
and U1549 (N_1549,In_247,In_119);
and U1550 (N_1550,In_751,In_365);
and U1551 (N_1551,In_1848,In_954);
or U1552 (N_1552,In_974,In_1957);
or U1553 (N_1553,In_524,In_1707);
nand U1554 (N_1554,In_325,In_608);
and U1555 (N_1555,In_577,In_1175);
nor U1556 (N_1556,In_44,In_1179);
and U1557 (N_1557,In_1073,In_179);
nor U1558 (N_1558,In_1879,In_489);
xnor U1559 (N_1559,In_343,In_1543);
nand U1560 (N_1560,In_1120,In_1731);
nor U1561 (N_1561,In_1363,In_1805);
or U1562 (N_1562,In_94,In_648);
or U1563 (N_1563,In_1217,In_528);
or U1564 (N_1564,In_422,In_1527);
or U1565 (N_1565,In_712,In_140);
nor U1566 (N_1566,In_945,In_715);
xor U1567 (N_1567,In_344,In_635);
or U1568 (N_1568,In_1617,In_1506);
xnor U1569 (N_1569,In_802,In_389);
xnor U1570 (N_1570,In_852,In_1951);
nor U1571 (N_1571,In_663,In_69);
and U1572 (N_1572,In_1674,In_1055);
nand U1573 (N_1573,In_1241,In_1589);
or U1574 (N_1574,In_818,In_1345);
or U1575 (N_1575,In_952,In_70);
xor U1576 (N_1576,In_325,In_191);
nor U1577 (N_1577,In_1048,In_190);
or U1578 (N_1578,In_1438,In_41);
nor U1579 (N_1579,In_409,In_911);
nand U1580 (N_1580,In_331,In_1229);
and U1581 (N_1581,In_318,In_1014);
nor U1582 (N_1582,In_1527,In_325);
nand U1583 (N_1583,In_1541,In_691);
xor U1584 (N_1584,In_159,In_960);
and U1585 (N_1585,In_782,In_276);
nor U1586 (N_1586,In_857,In_1045);
and U1587 (N_1587,In_772,In_345);
nand U1588 (N_1588,In_1643,In_607);
or U1589 (N_1589,In_892,In_1747);
xnor U1590 (N_1590,In_810,In_1007);
nand U1591 (N_1591,In_1614,In_271);
and U1592 (N_1592,In_825,In_563);
xor U1593 (N_1593,In_11,In_1080);
nand U1594 (N_1594,In_1510,In_756);
nand U1595 (N_1595,In_1714,In_862);
nand U1596 (N_1596,In_46,In_516);
or U1597 (N_1597,In_1562,In_103);
nor U1598 (N_1598,In_90,In_252);
nand U1599 (N_1599,In_754,In_227);
nand U1600 (N_1600,In_945,In_787);
xnor U1601 (N_1601,In_29,In_655);
or U1602 (N_1602,In_1439,In_1662);
xnor U1603 (N_1603,In_447,In_1949);
and U1604 (N_1604,In_1045,In_701);
and U1605 (N_1605,In_1359,In_1631);
or U1606 (N_1606,In_1506,In_1985);
or U1607 (N_1607,In_1625,In_1715);
and U1608 (N_1608,In_732,In_1302);
or U1609 (N_1609,In_1359,In_1507);
nand U1610 (N_1610,In_1794,In_1356);
and U1611 (N_1611,In_547,In_1560);
or U1612 (N_1612,In_289,In_1879);
nand U1613 (N_1613,In_964,In_19);
or U1614 (N_1614,In_1185,In_1154);
or U1615 (N_1615,In_1532,In_1234);
nor U1616 (N_1616,In_90,In_1292);
nor U1617 (N_1617,In_1125,In_122);
xnor U1618 (N_1618,In_1067,In_1640);
or U1619 (N_1619,In_1795,In_1614);
nand U1620 (N_1620,In_260,In_187);
xor U1621 (N_1621,In_1673,In_530);
and U1622 (N_1622,In_244,In_1654);
nand U1623 (N_1623,In_1677,In_182);
nand U1624 (N_1624,In_1734,In_1098);
nand U1625 (N_1625,In_1715,In_295);
nand U1626 (N_1626,In_1315,In_1130);
nor U1627 (N_1627,In_934,In_504);
nor U1628 (N_1628,In_496,In_1751);
xnor U1629 (N_1629,In_1962,In_1928);
xnor U1630 (N_1630,In_1010,In_421);
nand U1631 (N_1631,In_1941,In_1635);
nor U1632 (N_1632,In_978,In_938);
nor U1633 (N_1633,In_262,In_1201);
nand U1634 (N_1634,In_754,In_1232);
or U1635 (N_1635,In_527,In_1348);
xor U1636 (N_1636,In_886,In_1757);
or U1637 (N_1637,In_1688,In_693);
xor U1638 (N_1638,In_1013,In_1036);
or U1639 (N_1639,In_84,In_351);
or U1640 (N_1640,In_1786,In_1893);
xor U1641 (N_1641,In_429,In_198);
xnor U1642 (N_1642,In_1977,In_86);
and U1643 (N_1643,In_1957,In_1334);
xor U1644 (N_1644,In_58,In_551);
xnor U1645 (N_1645,In_430,In_302);
and U1646 (N_1646,In_597,In_957);
xnor U1647 (N_1647,In_1843,In_1058);
nor U1648 (N_1648,In_511,In_898);
or U1649 (N_1649,In_1105,In_168);
nor U1650 (N_1650,In_692,In_754);
or U1651 (N_1651,In_352,In_1522);
and U1652 (N_1652,In_1567,In_1453);
xor U1653 (N_1653,In_350,In_520);
xnor U1654 (N_1654,In_1789,In_1510);
nor U1655 (N_1655,In_1614,In_1315);
xnor U1656 (N_1656,In_442,In_1017);
xor U1657 (N_1657,In_71,In_255);
nand U1658 (N_1658,In_335,In_664);
or U1659 (N_1659,In_736,In_434);
nor U1660 (N_1660,In_1344,In_584);
nor U1661 (N_1661,In_74,In_970);
nor U1662 (N_1662,In_1717,In_660);
xnor U1663 (N_1663,In_258,In_853);
or U1664 (N_1664,In_969,In_221);
xnor U1665 (N_1665,In_1661,In_1212);
nand U1666 (N_1666,In_1813,In_596);
xor U1667 (N_1667,In_171,In_1713);
nor U1668 (N_1668,In_208,In_1525);
nand U1669 (N_1669,In_160,In_1823);
or U1670 (N_1670,In_443,In_1619);
and U1671 (N_1671,In_764,In_489);
nor U1672 (N_1672,In_1751,In_1580);
or U1673 (N_1673,In_757,In_1231);
or U1674 (N_1674,In_309,In_186);
and U1675 (N_1675,In_1758,In_1965);
nor U1676 (N_1676,In_891,In_1220);
and U1677 (N_1677,In_962,In_1578);
nand U1678 (N_1678,In_321,In_1606);
nor U1679 (N_1679,In_1340,In_1832);
and U1680 (N_1680,In_1469,In_32);
nand U1681 (N_1681,In_1992,In_375);
and U1682 (N_1682,In_714,In_208);
or U1683 (N_1683,In_495,In_1782);
xor U1684 (N_1684,In_1817,In_157);
nor U1685 (N_1685,In_1667,In_464);
xnor U1686 (N_1686,In_341,In_1205);
nand U1687 (N_1687,In_703,In_876);
nor U1688 (N_1688,In_920,In_766);
nand U1689 (N_1689,In_32,In_515);
or U1690 (N_1690,In_1070,In_943);
or U1691 (N_1691,In_1364,In_1923);
nor U1692 (N_1692,In_1081,In_280);
nand U1693 (N_1693,In_362,In_1443);
xor U1694 (N_1694,In_1716,In_971);
and U1695 (N_1695,In_1263,In_573);
or U1696 (N_1696,In_1393,In_732);
nor U1697 (N_1697,In_226,In_529);
or U1698 (N_1698,In_798,In_318);
and U1699 (N_1699,In_15,In_1069);
xor U1700 (N_1700,In_811,In_607);
or U1701 (N_1701,In_1728,In_380);
and U1702 (N_1702,In_225,In_910);
or U1703 (N_1703,In_1837,In_1020);
and U1704 (N_1704,In_1123,In_1461);
or U1705 (N_1705,In_1054,In_693);
or U1706 (N_1706,In_1122,In_367);
or U1707 (N_1707,In_1411,In_402);
or U1708 (N_1708,In_543,In_1426);
nand U1709 (N_1709,In_362,In_95);
xor U1710 (N_1710,In_1162,In_42);
nand U1711 (N_1711,In_1434,In_1326);
nor U1712 (N_1712,In_1908,In_531);
xor U1713 (N_1713,In_166,In_873);
nor U1714 (N_1714,In_726,In_264);
or U1715 (N_1715,In_1162,In_1271);
or U1716 (N_1716,In_428,In_1782);
and U1717 (N_1717,In_449,In_651);
nor U1718 (N_1718,In_872,In_1321);
xnor U1719 (N_1719,In_814,In_1294);
xor U1720 (N_1720,In_1502,In_1741);
xor U1721 (N_1721,In_1457,In_320);
and U1722 (N_1722,In_1772,In_1878);
nor U1723 (N_1723,In_121,In_325);
nand U1724 (N_1724,In_1554,In_1599);
nor U1725 (N_1725,In_1902,In_1948);
xor U1726 (N_1726,In_1295,In_282);
or U1727 (N_1727,In_1054,In_631);
and U1728 (N_1728,In_412,In_143);
xor U1729 (N_1729,In_482,In_1742);
nor U1730 (N_1730,In_51,In_1604);
and U1731 (N_1731,In_1971,In_102);
nand U1732 (N_1732,In_1170,In_1737);
and U1733 (N_1733,In_253,In_1629);
and U1734 (N_1734,In_1242,In_978);
xor U1735 (N_1735,In_1686,In_1822);
xnor U1736 (N_1736,In_900,In_586);
or U1737 (N_1737,In_1909,In_716);
nor U1738 (N_1738,In_420,In_1039);
or U1739 (N_1739,In_1375,In_187);
nand U1740 (N_1740,In_631,In_1620);
nor U1741 (N_1741,In_1686,In_320);
nand U1742 (N_1742,In_720,In_616);
nor U1743 (N_1743,In_1320,In_1297);
and U1744 (N_1744,In_994,In_221);
or U1745 (N_1745,In_1640,In_1009);
xnor U1746 (N_1746,In_525,In_397);
nand U1747 (N_1747,In_404,In_242);
nor U1748 (N_1748,In_926,In_1745);
or U1749 (N_1749,In_510,In_192);
xnor U1750 (N_1750,In_1440,In_140);
or U1751 (N_1751,In_958,In_689);
nand U1752 (N_1752,In_1624,In_1703);
xnor U1753 (N_1753,In_410,In_313);
nor U1754 (N_1754,In_1657,In_1241);
or U1755 (N_1755,In_1268,In_130);
nand U1756 (N_1756,In_665,In_335);
and U1757 (N_1757,In_1891,In_1567);
nor U1758 (N_1758,In_1271,In_489);
xnor U1759 (N_1759,In_578,In_371);
nand U1760 (N_1760,In_803,In_557);
or U1761 (N_1761,In_1197,In_1275);
nor U1762 (N_1762,In_1949,In_1897);
xor U1763 (N_1763,In_475,In_718);
or U1764 (N_1764,In_1132,In_1150);
or U1765 (N_1765,In_695,In_1878);
nand U1766 (N_1766,In_613,In_1119);
nor U1767 (N_1767,In_1569,In_714);
and U1768 (N_1768,In_1603,In_1589);
nand U1769 (N_1769,In_202,In_1202);
xnor U1770 (N_1770,In_762,In_982);
and U1771 (N_1771,In_193,In_661);
nand U1772 (N_1772,In_1014,In_1432);
xor U1773 (N_1773,In_1731,In_1989);
xor U1774 (N_1774,In_468,In_759);
nand U1775 (N_1775,In_914,In_1441);
nor U1776 (N_1776,In_1146,In_1894);
nand U1777 (N_1777,In_121,In_1014);
nor U1778 (N_1778,In_106,In_1281);
nor U1779 (N_1779,In_1135,In_962);
xor U1780 (N_1780,In_1659,In_835);
or U1781 (N_1781,In_916,In_297);
or U1782 (N_1782,In_1764,In_228);
nand U1783 (N_1783,In_1242,In_1124);
and U1784 (N_1784,In_450,In_802);
nand U1785 (N_1785,In_1103,In_1148);
or U1786 (N_1786,In_710,In_197);
or U1787 (N_1787,In_596,In_755);
nand U1788 (N_1788,In_1952,In_1954);
nor U1789 (N_1789,In_1254,In_1923);
or U1790 (N_1790,In_224,In_757);
xor U1791 (N_1791,In_1891,In_335);
and U1792 (N_1792,In_53,In_262);
nor U1793 (N_1793,In_1161,In_1005);
xor U1794 (N_1794,In_790,In_679);
nor U1795 (N_1795,In_1753,In_350);
xor U1796 (N_1796,In_356,In_1562);
nand U1797 (N_1797,In_468,In_1581);
xnor U1798 (N_1798,In_652,In_290);
nor U1799 (N_1799,In_1901,In_1177);
nand U1800 (N_1800,In_1008,In_735);
and U1801 (N_1801,In_1995,In_1264);
nor U1802 (N_1802,In_1632,In_570);
nand U1803 (N_1803,In_1883,In_1914);
and U1804 (N_1804,In_1785,In_1375);
nor U1805 (N_1805,In_1112,In_1014);
and U1806 (N_1806,In_171,In_345);
nand U1807 (N_1807,In_125,In_1541);
and U1808 (N_1808,In_371,In_174);
nor U1809 (N_1809,In_591,In_1722);
and U1810 (N_1810,In_672,In_183);
and U1811 (N_1811,In_297,In_961);
nand U1812 (N_1812,In_1246,In_1433);
nor U1813 (N_1813,In_1663,In_1331);
nand U1814 (N_1814,In_664,In_1488);
nand U1815 (N_1815,In_371,In_1919);
xnor U1816 (N_1816,In_505,In_867);
xnor U1817 (N_1817,In_155,In_1520);
nor U1818 (N_1818,In_1333,In_1306);
nand U1819 (N_1819,In_268,In_589);
and U1820 (N_1820,In_1674,In_594);
and U1821 (N_1821,In_676,In_1142);
or U1822 (N_1822,In_1159,In_1620);
nor U1823 (N_1823,In_671,In_303);
nor U1824 (N_1824,In_559,In_27);
nand U1825 (N_1825,In_252,In_1700);
nand U1826 (N_1826,In_1114,In_908);
nand U1827 (N_1827,In_1699,In_560);
nand U1828 (N_1828,In_1452,In_550);
and U1829 (N_1829,In_972,In_1659);
nor U1830 (N_1830,In_256,In_1515);
or U1831 (N_1831,In_1542,In_1439);
nor U1832 (N_1832,In_1841,In_1313);
nor U1833 (N_1833,In_1091,In_1453);
or U1834 (N_1834,In_1294,In_440);
xor U1835 (N_1835,In_854,In_1930);
or U1836 (N_1836,In_1439,In_11);
nor U1837 (N_1837,In_1208,In_906);
or U1838 (N_1838,In_1768,In_1174);
or U1839 (N_1839,In_1515,In_397);
xnor U1840 (N_1840,In_305,In_745);
and U1841 (N_1841,In_1777,In_679);
nand U1842 (N_1842,In_607,In_1768);
or U1843 (N_1843,In_242,In_985);
xor U1844 (N_1844,In_1049,In_680);
nor U1845 (N_1845,In_334,In_1285);
xnor U1846 (N_1846,In_505,In_1714);
and U1847 (N_1847,In_1039,In_715);
and U1848 (N_1848,In_968,In_131);
nor U1849 (N_1849,In_1057,In_1442);
nor U1850 (N_1850,In_401,In_1645);
or U1851 (N_1851,In_102,In_1462);
nand U1852 (N_1852,In_801,In_1135);
nor U1853 (N_1853,In_1460,In_934);
xor U1854 (N_1854,In_1479,In_331);
nand U1855 (N_1855,In_239,In_1153);
and U1856 (N_1856,In_1744,In_256);
or U1857 (N_1857,In_1008,In_314);
xnor U1858 (N_1858,In_1964,In_1419);
nor U1859 (N_1859,In_1928,In_1872);
nor U1860 (N_1860,In_523,In_573);
xor U1861 (N_1861,In_1844,In_340);
nand U1862 (N_1862,In_1356,In_1706);
xor U1863 (N_1863,In_93,In_391);
or U1864 (N_1864,In_255,In_419);
nor U1865 (N_1865,In_1470,In_976);
or U1866 (N_1866,In_911,In_1303);
or U1867 (N_1867,In_1887,In_1290);
and U1868 (N_1868,In_1432,In_477);
or U1869 (N_1869,In_1995,In_1558);
and U1870 (N_1870,In_929,In_769);
nand U1871 (N_1871,In_1479,In_1048);
nand U1872 (N_1872,In_1766,In_1645);
nor U1873 (N_1873,In_1793,In_1104);
and U1874 (N_1874,In_1814,In_1385);
nand U1875 (N_1875,In_1691,In_564);
xor U1876 (N_1876,In_1469,In_1728);
nor U1877 (N_1877,In_871,In_1226);
nand U1878 (N_1878,In_1916,In_580);
nor U1879 (N_1879,In_1296,In_20);
and U1880 (N_1880,In_1215,In_1060);
or U1881 (N_1881,In_1999,In_772);
xor U1882 (N_1882,In_1431,In_50);
nor U1883 (N_1883,In_1544,In_1173);
nor U1884 (N_1884,In_399,In_157);
and U1885 (N_1885,In_354,In_1027);
and U1886 (N_1886,In_6,In_790);
or U1887 (N_1887,In_723,In_354);
xnor U1888 (N_1888,In_380,In_49);
or U1889 (N_1889,In_549,In_1449);
nor U1890 (N_1890,In_915,In_1456);
nand U1891 (N_1891,In_1043,In_303);
nor U1892 (N_1892,In_941,In_1880);
and U1893 (N_1893,In_593,In_970);
xor U1894 (N_1894,In_329,In_832);
nand U1895 (N_1895,In_1252,In_1830);
xor U1896 (N_1896,In_1110,In_1582);
or U1897 (N_1897,In_299,In_1262);
nor U1898 (N_1898,In_939,In_924);
and U1899 (N_1899,In_262,In_490);
nand U1900 (N_1900,In_476,In_1776);
or U1901 (N_1901,In_996,In_499);
or U1902 (N_1902,In_1437,In_709);
xnor U1903 (N_1903,In_677,In_803);
nand U1904 (N_1904,In_553,In_810);
nor U1905 (N_1905,In_1224,In_1450);
nor U1906 (N_1906,In_702,In_1798);
or U1907 (N_1907,In_1128,In_65);
nor U1908 (N_1908,In_444,In_832);
nor U1909 (N_1909,In_1361,In_117);
or U1910 (N_1910,In_323,In_1770);
xor U1911 (N_1911,In_1313,In_1170);
nor U1912 (N_1912,In_1370,In_1341);
and U1913 (N_1913,In_718,In_647);
or U1914 (N_1914,In_1508,In_1441);
and U1915 (N_1915,In_286,In_90);
nor U1916 (N_1916,In_1716,In_1394);
or U1917 (N_1917,In_1086,In_11);
xnor U1918 (N_1918,In_1318,In_303);
nand U1919 (N_1919,In_1855,In_1906);
nor U1920 (N_1920,In_300,In_902);
and U1921 (N_1921,In_1776,In_1117);
xor U1922 (N_1922,In_1349,In_1699);
xnor U1923 (N_1923,In_1960,In_1881);
and U1924 (N_1924,In_1482,In_1276);
nor U1925 (N_1925,In_666,In_557);
nor U1926 (N_1926,In_1656,In_1045);
xor U1927 (N_1927,In_1482,In_1173);
xor U1928 (N_1928,In_197,In_1935);
or U1929 (N_1929,In_1507,In_484);
nand U1930 (N_1930,In_576,In_746);
nor U1931 (N_1931,In_1838,In_1524);
or U1932 (N_1932,In_1590,In_462);
or U1933 (N_1933,In_533,In_801);
and U1934 (N_1934,In_743,In_1178);
nor U1935 (N_1935,In_249,In_1108);
and U1936 (N_1936,In_461,In_1019);
and U1937 (N_1937,In_995,In_1306);
nor U1938 (N_1938,In_620,In_869);
nand U1939 (N_1939,In_1824,In_636);
nor U1940 (N_1940,In_1099,In_1821);
and U1941 (N_1941,In_1695,In_1281);
nand U1942 (N_1942,In_1704,In_1808);
xnor U1943 (N_1943,In_551,In_244);
nor U1944 (N_1944,In_79,In_169);
nor U1945 (N_1945,In_1738,In_738);
nand U1946 (N_1946,In_542,In_1593);
xnor U1947 (N_1947,In_421,In_204);
nand U1948 (N_1948,In_831,In_173);
or U1949 (N_1949,In_1318,In_1094);
nor U1950 (N_1950,In_1845,In_746);
nor U1951 (N_1951,In_1683,In_638);
and U1952 (N_1952,In_563,In_1854);
xor U1953 (N_1953,In_612,In_1072);
or U1954 (N_1954,In_896,In_725);
xor U1955 (N_1955,In_227,In_300);
nand U1956 (N_1956,In_1063,In_1086);
xor U1957 (N_1957,In_1145,In_1111);
and U1958 (N_1958,In_823,In_1768);
xnor U1959 (N_1959,In_12,In_492);
nor U1960 (N_1960,In_658,In_1435);
nor U1961 (N_1961,In_12,In_1050);
nor U1962 (N_1962,In_713,In_1769);
and U1963 (N_1963,In_1934,In_1784);
nand U1964 (N_1964,In_1152,In_329);
xnor U1965 (N_1965,In_1220,In_825);
nand U1966 (N_1966,In_987,In_836);
xnor U1967 (N_1967,In_1927,In_392);
nand U1968 (N_1968,In_250,In_568);
or U1969 (N_1969,In_1159,In_1775);
xnor U1970 (N_1970,In_928,In_1239);
or U1971 (N_1971,In_1846,In_1961);
nand U1972 (N_1972,In_195,In_363);
or U1973 (N_1973,In_583,In_251);
nor U1974 (N_1974,In_128,In_732);
or U1975 (N_1975,In_1764,In_599);
and U1976 (N_1976,In_1306,In_1041);
or U1977 (N_1977,In_929,In_1698);
nor U1978 (N_1978,In_1991,In_638);
nor U1979 (N_1979,In_1726,In_1179);
xnor U1980 (N_1980,In_655,In_325);
xnor U1981 (N_1981,In_1738,In_769);
nand U1982 (N_1982,In_1425,In_1573);
or U1983 (N_1983,In_1640,In_600);
or U1984 (N_1984,In_397,In_1960);
xor U1985 (N_1985,In_690,In_295);
nand U1986 (N_1986,In_1249,In_324);
or U1987 (N_1987,In_133,In_1123);
nor U1988 (N_1988,In_1574,In_1216);
nand U1989 (N_1989,In_634,In_1995);
nand U1990 (N_1990,In_1288,In_1095);
nor U1991 (N_1991,In_985,In_565);
or U1992 (N_1992,In_411,In_1473);
and U1993 (N_1993,In_998,In_1410);
or U1994 (N_1994,In_1277,In_1180);
or U1995 (N_1995,In_339,In_818);
and U1996 (N_1996,In_19,In_1718);
and U1997 (N_1997,In_989,In_635);
nor U1998 (N_1998,In_80,In_1774);
xor U1999 (N_1999,In_1296,In_297);
or U2000 (N_2000,In_818,In_1048);
nor U2001 (N_2001,In_1840,In_1053);
and U2002 (N_2002,In_1099,In_661);
nand U2003 (N_2003,In_1967,In_161);
or U2004 (N_2004,In_361,In_1172);
nand U2005 (N_2005,In_420,In_1937);
and U2006 (N_2006,In_560,In_1055);
nor U2007 (N_2007,In_1566,In_1894);
nand U2008 (N_2008,In_389,In_1308);
or U2009 (N_2009,In_1479,In_512);
or U2010 (N_2010,In_604,In_757);
and U2011 (N_2011,In_1509,In_1995);
nor U2012 (N_2012,In_1754,In_278);
and U2013 (N_2013,In_1589,In_1050);
nor U2014 (N_2014,In_95,In_1423);
nor U2015 (N_2015,In_396,In_1866);
nand U2016 (N_2016,In_1551,In_469);
and U2017 (N_2017,In_1816,In_1270);
xnor U2018 (N_2018,In_420,In_867);
nor U2019 (N_2019,In_1407,In_253);
nor U2020 (N_2020,In_1237,In_1670);
nand U2021 (N_2021,In_4,In_339);
nor U2022 (N_2022,In_501,In_11);
and U2023 (N_2023,In_1069,In_1762);
nor U2024 (N_2024,In_1530,In_1273);
xnor U2025 (N_2025,In_1680,In_1345);
nand U2026 (N_2026,In_291,In_780);
nor U2027 (N_2027,In_1616,In_1814);
nand U2028 (N_2028,In_1354,In_820);
nor U2029 (N_2029,In_206,In_1026);
xnor U2030 (N_2030,In_1127,In_1523);
nor U2031 (N_2031,In_1512,In_37);
or U2032 (N_2032,In_311,In_1790);
nand U2033 (N_2033,In_259,In_1141);
xor U2034 (N_2034,In_1197,In_1883);
nand U2035 (N_2035,In_1137,In_1660);
or U2036 (N_2036,In_1149,In_1893);
xor U2037 (N_2037,In_1301,In_868);
or U2038 (N_2038,In_1267,In_1082);
xor U2039 (N_2039,In_804,In_1994);
nand U2040 (N_2040,In_1151,In_1438);
and U2041 (N_2041,In_1619,In_1471);
or U2042 (N_2042,In_1088,In_1193);
nor U2043 (N_2043,In_1073,In_806);
nor U2044 (N_2044,In_1327,In_1739);
or U2045 (N_2045,In_891,In_1403);
nand U2046 (N_2046,In_1616,In_1139);
and U2047 (N_2047,In_1383,In_1042);
or U2048 (N_2048,In_293,In_1779);
and U2049 (N_2049,In_1908,In_1708);
and U2050 (N_2050,In_245,In_1208);
nor U2051 (N_2051,In_1792,In_1147);
xor U2052 (N_2052,In_1250,In_86);
and U2053 (N_2053,In_1161,In_1427);
xor U2054 (N_2054,In_206,In_15);
and U2055 (N_2055,In_620,In_934);
nor U2056 (N_2056,In_1165,In_932);
or U2057 (N_2057,In_673,In_1391);
and U2058 (N_2058,In_663,In_1473);
nand U2059 (N_2059,In_1858,In_1475);
nor U2060 (N_2060,In_917,In_34);
and U2061 (N_2061,In_1755,In_67);
and U2062 (N_2062,In_1604,In_1414);
and U2063 (N_2063,In_1031,In_684);
nor U2064 (N_2064,In_698,In_469);
and U2065 (N_2065,In_1258,In_719);
nand U2066 (N_2066,In_1806,In_1969);
or U2067 (N_2067,In_437,In_319);
and U2068 (N_2068,In_1662,In_1447);
and U2069 (N_2069,In_867,In_1652);
or U2070 (N_2070,In_309,In_1346);
and U2071 (N_2071,In_174,In_1739);
nor U2072 (N_2072,In_1248,In_1915);
nand U2073 (N_2073,In_1425,In_545);
or U2074 (N_2074,In_490,In_1231);
and U2075 (N_2075,In_156,In_1494);
xor U2076 (N_2076,In_821,In_1457);
nand U2077 (N_2077,In_1449,In_1207);
and U2078 (N_2078,In_1289,In_1545);
xor U2079 (N_2079,In_1229,In_738);
and U2080 (N_2080,In_537,In_227);
xnor U2081 (N_2081,In_883,In_345);
and U2082 (N_2082,In_1104,In_1258);
nand U2083 (N_2083,In_760,In_422);
or U2084 (N_2084,In_116,In_1455);
nand U2085 (N_2085,In_108,In_107);
xor U2086 (N_2086,In_1750,In_1516);
and U2087 (N_2087,In_1547,In_2);
xor U2088 (N_2088,In_58,In_638);
and U2089 (N_2089,In_872,In_256);
and U2090 (N_2090,In_1929,In_943);
xnor U2091 (N_2091,In_1237,In_1663);
nand U2092 (N_2092,In_1768,In_1112);
nor U2093 (N_2093,In_380,In_1979);
or U2094 (N_2094,In_1990,In_215);
or U2095 (N_2095,In_1383,In_1140);
nand U2096 (N_2096,In_1641,In_914);
or U2097 (N_2097,In_405,In_567);
nand U2098 (N_2098,In_300,In_1657);
nand U2099 (N_2099,In_674,In_909);
nor U2100 (N_2100,In_802,In_1213);
xor U2101 (N_2101,In_166,In_1761);
xnor U2102 (N_2102,In_1777,In_25);
nor U2103 (N_2103,In_138,In_353);
xnor U2104 (N_2104,In_1501,In_359);
nor U2105 (N_2105,In_501,In_1555);
xnor U2106 (N_2106,In_1983,In_788);
xor U2107 (N_2107,In_953,In_1961);
and U2108 (N_2108,In_1800,In_549);
nor U2109 (N_2109,In_1598,In_84);
or U2110 (N_2110,In_905,In_1048);
nand U2111 (N_2111,In_1258,In_292);
xor U2112 (N_2112,In_291,In_179);
xor U2113 (N_2113,In_878,In_1302);
or U2114 (N_2114,In_532,In_1858);
nand U2115 (N_2115,In_398,In_834);
nor U2116 (N_2116,In_971,In_1835);
xor U2117 (N_2117,In_1586,In_339);
nor U2118 (N_2118,In_1446,In_1517);
xnor U2119 (N_2119,In_1493,In_769);
xor U2120 (N_2120,In_1028,In_621);
nand U2121 (N_2121,In_106,In_57);
nor U2122 (N_2122,In_1488,In_726);
or U2123 (N_2123,In_1791,In_549);
nand U2124 (N_2124,In_692,In_607);
and U2125 (N_2125,In_1456,In_714);
and U2126 (N_2126,In_125,In_1207);
and U2127 (N_2127,In_682,In_38);
xnor U2128 (N_2128,In_504,In_228);
or U2129 (N_2129,In_409,In_379);
nor U2130 (N_2130,In_1276,In_1635);
xnor U2131 (N_2131,In_1972,In_659);
and U2132 (N_2132,In_1620,In_1718);
nor U2133 (N_2133,In_891,In_425);
and U2134 (N_2134,In_938,In_945);
nor U2135 (N_2135,In_1248,In_1326);
and U2136 (N_2136,In_454,In_561);
xor U2137 (N_2137,In_377,In_1641);
or U2138 (N_2138,In_1456,In_514);
and U2139 (N_2139,In_479,In_1123);
nand U2140 (N_2140,In_1633,In_302);
nor U2141 (N_2141,In_1702,In_1621);
nor U2142 (N_2142,In_1058,In_843);
xor U2143 (N_2143,In_926,In_585);
and U2144 (N_2144,In_468,In_89);
and U2145 (N_2145,In_195,In_1747);
nor U2146 (N_2146,In_1246,In_1449);
nor U2147 (N_2147,In_1545,In_686);
and U2148 (N_2148,In_1473,In_526);
or U2149 (N_2149,In_494,In_1899);
nor U2150 (N_2150,In_1885,In_234);
nor U2151 (N_2151,In_1018,In_1443);
and U2152 (N_2152,In_656,In_422);
nor U2153 (N_2153,In_822,In_1025);
nand U2154 (N_2154,In_884,In_1884);
and U2155 (N_2155,In_904,In_1840);
nor U2156 (N_2156,In_241,In_414);
and U2157 (N_2157,In_660,In_1265);
and U2158 (N_2158,In_1728,In_868);
nand U2159 (N_2159,In_613,In_1148);
and U2160 (N_2160,In_1477,In_346);
and U2161 (N_2161,In_278,In_306);
nand U2162 (N_2162,In_1086,In_1130);
nand U2163 (N_2163,In_450,In_599);
nor U2164 (N_2164,In_193,In_354);
xor U2165 (N_2165,In_104,In_718);
and U2166 (N_2166,In_702,In_688);
nor U2167 (N_2167,In_502,In_1009);
xnor U2168 (N_2168,In_1464,In_1584);
xnor U2169 (N_2169,In_414,In_1070);
nand U2170 (N_2170,In_291,In_192);
xor U2171 (N_2171,In_1268,In_1333);
xor U2172 (N_2172,In_284,In_462);
nor U2173 (N_2173,In_1543,In_1128);
nand U2174 (N_2174,In_946,In_939);
nand U2175 (N_2175,In_1653,In_795);
xnor U2176 (N_2176,In_1696,In_857);
or U2177 (N_2177,In_1941,In_991);
or U2178 (N_2178,In_378,In_1500);
nand U2179 (N_2179,In_1248,In_676);
xor U2180 (N_2180,In_1146,In_423);
nand U2181 (N_2181,In_1402,In_1883);
xor U2182 (N_2182,In_9,In_937);
nand U2183 (N_2183,In_786,In_317);
nor U2184 (N_2184,In_685,In_1037);
nor U2185 (N_2185,In_1293,In_145);
and U2186 (N_2186,In_1930,In_78);
nand U2187 (N_2187,In_1444,In_1350);
nor U2188 (N_2188,In_1144,In_975);
and U2189 (N_2189,In_1095,In_703);
nor U2190 (N_2190,In_1681,In_1570);
xnor U2191 (N_2191,In_1836,In_1490);
nor U2192 (N_2192,In_1326,In_158);
and U2193 (N_2193,In_966,In_1417);
or U2194 (N_2194,In_1055,In_1839);
xnor U2195 (N_2195,In_577,In_187);
xnor U2196 (N_2196,In_608,In_502);
nor U2197 (N_2197,In_1394,In_1693);
or U2198 (N_2198,In_387,In_819);
nor U2199 (N_2199,In_22,In_1707);
nor U2200 (N_2200,In_634,In_440);
and U2201 (N_2201,In_809,In_1105);
xor U2202 (N_2202,In_1960,In_1157);
nand U2203 (N_2203,In_1141,In_420);
or U2204 (N_2204,In_1959,In_1934);
nor U2205 (N_2205,In_1047,In_1);
nand U2206 (N_2206,In_1862,In_1822);
or U2207 (N_2207,In_1302,In_742);
or U2208 (N_2208,In_713,In_882);
or U2209 (N_2209,In_1446,In_1209);
xor U2210 (N_2210,In_1642,In_854);
and U2211 (N_2211,In_405,In_407);
or U2212 (N_2212,In_1048,In_1693);
and U2213 (N_2213,In_488,In_936);
xor U2214 (N_2214,In_183,In_1433);
and U2215 (N_2215,In_949,In_1473);
and U2216 (N_2216,In_301,In_758);
xor U2217 (N_2217,In_271,In_1567);
and U2218 (N_2218,In_701,In_782);
or U2219 (N_2219,In_1936,In_980);
nor U2220 (N_2220,In_1288,In_1449);
nand U2221 (N_2221,In_1041,In_1242);
and U2222 (N_2222,In_1060,In_278);
and U2223 (N_2223,In_1887,In_1992);
and U2224 (N_2224,In_1697,In_1661);
nand U2225 (N_2225,In_1372,In_153);
nor U2226 (N_2226,In_1827,In_1576);
nand U2227 (N_2227,In_1875,In_103);
or U2228 (N_2228,In_1453,In_1804);
xor U2229 (N_2229,In_355,In_193);
nor U2230 (N_2230,In_324,In_1896);
nor U2231 (N_2231,In_1749,In_1787);
or U2232 (N_2232,In_1240,In_629);
nor U2233 (N_2233,In_547,In_684);
xor U2234 (N_2234,In_798,In_1472);
nand U2235 (N_2235,In_1416,In_1810);
xnor U2236 (N_2236,In_1999,In_779);
or U2237 (N_2237,In_1330,In_1426);
and U2238 (N_2238,In_871,In_1025);
and U2239 (N_2239,In_905,In_1439);
xnor U2240 (N_2240,In_1292,In_1688);
nor U2241 (N_2241,In_1502,In_809);
or U2242 (N_2242,In_1513,In_462);
nand U2243 (N_2243,In_770,In_1128);
nor U2244 (N_2244,In_694,In_469);
and U2245 (N_2245,In_1734,In_79);
and U2246 (N_2246,In_183,In_0);
nor U2247 (N_2247,In_691,In_1847);
and U2248 (N_2248,In_165,In_339);
xor U2249 (N_2249,In_1294,In_269);
and U2250 (N_2250,In_1085,In_674);
and U2251 (N_2251,In_1208,In_666);
or U2252 (N_2252,In_383,In_558);
nand U2253 (N_2253,In_1754,In_595);
or U2254 (N_2254,In_231,In_764);
nand U2255 (N_2255,In_148,In_1959);
nand U2256 (N_2256,In_1611,In_276);
xnor U2257 (N_2257,In_325,In_782);
nor U2258 (N_2258,In_36,In_1002);
and U2259 (N_2259,In_772,In_528);
and U2260 (N_2260,In_570,In_1802);
nor U2261 (N_2261,In_1822,In_355);
or U2262 (N_2262,In_1862,In_950);
nor U2263 (N_2263,In_1170,In_462);
or U2264 (N_2264,In_1341,In_844);
and U2265 (N_2265,In_1217,In_1949);
and U2266 (N_2266,In_1095,In_218);
or U2267 (N_2267,In_1398,In_1204);
or U2268 (N_2268,In_877,In_1725);
or U2269 (N_2269,In_1853,In_849);
and U2270 (N_2270,In_1694,In_1244);
or U2271 (N_2271,In_476,In_1561);
nand U2272 (N_2272,In_21,In_203);
nor U2273 (N_2273,In_1734,In_1021);
nor U2274 (N_2274,In_768,In_154);
and U2275 (N_2275,In_787,In_1159);
or U2276 (N_2276,In_628,In_1544);
nor U2277 (N_2277,In_1030,In_251);
nand U2278 (N_2278,In_1209,In_5);
nor U2279 (N_2279,In_791,In_1357);
and U2280 (N_2280,In_1684,In_1500);
nand U2281 (N_2281,In_730,In_735);
nor U2282 (N_2282,In_1515,In_58);
xor U2283 (N_2283,In_1094,In_277);
nand U2284 (N_2284,In_1688,In_119);
and U2285 (N_2285,In_379,In_1491);
and U2286 (N_2286,In_196,In_61);
and U2287 (N_2287,In_1935,In_519);
nor U2288 (N_2288,In_1627,In_1456);
xor U2289 (N_2289,In_1129,In_975);
xnor U2290 (N_2290,In_826,In_655);
or U2291 (N_2291,In_1453,In_379);
xor U2292 (N_2292,In_83,In_832);
nand U2293 (N_2293,In_1546,In_1213);
or U2294 (N_2294,In_1875,In_1939);
and U2295 (N_2295,In_557,In_1421);
or U2296 (N_2296,In_1617,In_1343);
or U2297 (N_2297,In_1664,In_1630);
xnor U2298 (N_2298,In_1191,In_212);
nor U2299 (N_2299,In_81,In_1074);
nor U2300 (N_2300,In_20,In_1277);
nand U2301 (N_2301,In_587,In_299);
or U2302 (N_2302,In_818,In_765);
xor U2303 (N_2303,In_1049,In_1174);
nand U2304 (N_2304,In_578,In_1591);
or U2305 (N_2305,In_1055,In_116);
and U2306 (N_2306,In_541,In_487);
nor U2307 (N_2307,In_754,In_279);
nor U2308 (N_2308,In_1962,In_639);
nor U2309 (N_2309,In_1962,In_1884);
nor U2310 (N_2310,In_1342,In_1985);
nand U2311 (N_2311,In_1003,In_1835);
and U2312 (N_2312,In_239,In_721);
or U2313 (N_2313,In_614,In_1377);
nor U2314 (N_2314,In_1669,In_1227);
or U2315 (N_2315,In_1379,In_873);
or U2316 (N_2316,In_95,In_1926);
nor U2317 (N_2317,In_1983,In_216);
nand U2318 (N_2318,In_1038,In_1079);
or U2319 (N_2319,In_799,In_1822);
xnor U2320 (N_2320,In_724,In_124);
xor U2321 (N_2321,In_1761,In_1916);
or U2322 (N_2322,In_417,In_737);
xor U2323 (N_2323,In_1366,In_1901);
nor U2324 (N_2324,In_748,In_629);
nor U2325 (N_2325,In_995,In_1805);
nand U2326 (N_2326,In_1587,In_1814);
nand U2327 (N_2327,In_639,In_649);
and U2328 (N_2328,In_826,In_955);
nor U2329 (N_2329,In_1256,In_1143);
xor U2330 (N_2330,In_405,In_1103);
or U2331 (N_2331,In_615,In_14);
and U2332 (N_2332,In_596,In_581);
xnor U2333 (N_2333,In_208,In_1521);
nand U2334 (N_2334,In_750,In_701);
xnor U2335 (N_2335,In_65,In_1470);
and U2336 (N_2336,In_1941,In_780);
xor U2337 (N_2337,In_662,In_1312);
and U2338 (N_2338,In_1410,In_757);
and U2339 (N_2339,In_1203,In_104);
nand U2340 (N_2340,In_1334,In_182);
nor U2341 (N_2341,In_602,In_1989);
nand U2342 (N_2342,In_1721,In_970);
or U2343 (N_2343,In_1837,In_911);
and U2344 (N_2344,In_377,In_19);
nor U2345 (N_2345,In_19,In_1251);
nor U2346 (N_2346,In_1808,In_424);
nor U2347 (N_2347,In_781,In_599);
or U2348 (N_2348,In_1705,In_70);
xnor U2349 (N_2349,In_932,In_1572);
xor U2350 (N_2350,In_588,In_1757);
nor U2351 (N_2351,In_1050,In_1992);
nand U2352 (N_2352,In_1887,In_1014);
xnor U2353 (N_2353,In_449,In_481);
xnor U2354 (N_2354,In_389,In_1143);
nor U2355 (N_2355,In_617,In_824);
or U2356 (N_2356,In_626,In_1101);
or U2357 (N_2357,In_824,In_1474);
and U2358 (N_2358,In_444,In_1978);
nand U2359 (N_2359,In_1128,In_1782);
or U2360 (N_2360,In_1879,In_1801);
and U2361 (N_2361,In_1204,In_760);
xor U2362 (N_2362,In_13,In_1482);
nand U2363 (N_2363,In_867,In_1454);
and U2364 (N_2364,In_582,In_1187);
and U2365 (N_2365,In_3,In_1491);
and U2366 (N_2366,In_163,In_1944);
and U2367 (N_2367,In_1230,In_1804);
nand U2368 (N_2368,In_1344,In_241);
xnor U2369 (N_2369,In_98,In_844);
xor U2370 (N_2370,In_1317,In_1839);
and U2371 (N_2371,In_943,In_1239);
nand U2372 (N_2372,In_1186,In_1360);
and U2373 (N_2373,In_1495,In_1581);
nor U2374 (N_2374,In_317,In_1661);
nand U2375 (N_2375,In_825,In_836);
or U2376 (N_2376,In_1797,In_880);
and U2377 (N_2377,In_1740,In_590);
and U2378 (N_2378,In_1551,In_146);
nand U2379 (N_2379,In_584,In_987);
or U2380 (N_2380,In_1481,In_1559);
nor U2381 (N_2381,In_571,In_65);
nor U2382 (N_2382,In_1647,In_389);
or U2383 (N_2383,In_1718,In_314);
xnor U2384 (N_2384,In_657,In_1662);
and U2385 (N_2385,In_1656,In_1528);
xnor U2386 (N_2386,In_891,In_440);
and U2387 (N_2387,In_1165,In_1913);
nand U2388 (N_2388,In_1908,In_1005);
nor U2389 (N_2389,In_573,In_742);
xor U2390 (N_2390,In_89,In_1380);
nor U2391 (N_2391,In_573,In_1427);
nand U2392 (N_2392,In_122,In_1480);
or U2393 (N_2393,In_1890,In_1519);
and U2394 (N_2394,In_770,In_50);
xor U2395 (N_2395,In_22,In_865);
and U2396 (N_2396,In_1692,In_1009);
nor U2397 (N_2397,In_99,In_1462);
nand U2398 (N_2398,In_1886,In_1078);
or U2399 (N_2399,In_1759,In_1988);
xnor U2400 (N_2400,In_200,In_1909);
xor U2401 (N_2401,In_205,In_217);
nand U2402 (N_2402,In_1751,In_222);
nor U2403 (N_2403,In_370,In_1685);
nor U2404 (N_2404,In_1842,In_1758);
and U2405 (N_2405,In_839,In_585);
and U2406 (N_2406,In_1187,In_1262);
nor U2407 (N_2407,In_1736,In_1240);
and U2408 (N_2408,In_1239,In_897);
nand U2409 (N_2409,In_852,In_1978);
xor U2410 (N_2410,In_357,In_979);
or U2411 (N_2411,In_1211,In_1186);
nor U2412 (N_2412,In_1198,In_697);
xnor U2413 (N_2413,In_1866,In_7);
and U2414 (N_2414,In_1390,In_666);
nor U2415 (N_2415,In_621,In_754);
xnor U2416 (N_2416,In_313,In_573);
or U2417 (N_2417,In_1758,In_1906);
xnor U2418 (N_2418,In_284,In_1267);
and U2419 (N_2419,In_1976,In_944);
or U2420 (N_2420,In_191,In_853);
nor U2421 (N_2421,In_23,In_1874);
nand U2422 (N_2422,In_1637,In_1536);
nand U2423 (N_2423,In_1880,In_352);
nor U2424 (N_2424,In_510,In_1368);
or U2425 (N_2425,In_1887,In_831);
and U2426 (N_2426,In_891,In_1584);
and U2427 (N_2427,In_1429,In_1659);
nand U2428 (N_2428,In_1325,In_613);
and U2429 (N_2429,In_1196,In_899);
xnor U2430 (N_2430,In_1719,In_1849);
nor U2431 (N_2431,In_335,In_1988);
nor U2432 (N_2432,In_745,In_1717);
and U2433 (N_2433,In_1331,In_783);
xnor U2434 (N_2434,In_973,In_554);
or U2435 (N_2435,In_910,In_938);
xnor U2436 (N_2436,In_755,In_1632);
nor U2437 (N_2437,In_66,In_1565);
nand U2438 (N_2438,In_545,In_1883);
and U2439 (N_2439,In_1751,In_1121);
nor U2440 (N_2440,In_1618,In_1619);
and U2441 (N_2441,In_1401,In_1258);
and U2442 (N_2442,In_1001,In_1254);
nor U2443 (N_2443,In_102,In_1172);
and U2444 (N_2444,In_780,In_1349);
or U2445 (N_2445,In_1402,In_1024);
nor U2446 (N_2446,In_1046,In_1043);
and U2447 (N_2447,In_1763,In_1701);
nand U2448 (N_2448,In_1790,In_1436);
nor U2449 (N_2449,In_1895,In_292);
nor U2450 (N_2450,In_1317,In_1650);
nand U2451 (N_2451,In_892,In_524);
nor U2452 (N_2452,In_1403,In_455);
or U2453 (N_2453,In_1037,In_44);
or U2454 (N_2454,In_526,In_1456);
nand U2455 (N_2455,In_936,In_287);
or U2456 (N_2456,In_823,In_992);
nor U2457 (N_2457,In_31,In_273);
or U2458 (N_2458,In_445,In_1277);
and U2459 (N_2459,In_1707,In_294);
nand U2460 (N_2460,In_1443,In_222);
or U2461 (N_2461,In_1235,In_1888);
and U2462 (N_2462,In_1879,In_1585);
nand U2463 (N_2463,In_351,In_438);
or U2464 (N_2464,In_159,In_1826);
nor U2465 (N_2465,In_1622,In_1333);
and U2466 (N_2466,In_1918,In_1971);
nor U2467 (N_2467,In_609,In_1899);
or U2468 (N_2468,In_1529,In_1494);
or U2469 (N_2469,In_668,In_10);
and U2470 (N_2470,In_664,In_787);
or U2471 (N_2471,In_22,In_117);
and U2472 (N_2472,In_640,In_1440);
or U2473 (N_2473,In_1609,In_852);
xnor U2474 (N_2474,In_1280,In_412);
and U2475 (N_2475,In_186,In_218);
and U2476 (N_2476,In_1140,In_1669);
and U2477 (N_2477,In_1764,In_789);
xor U2478 (N_2478,In_471,In_1146);
or U2479 (N_2479,In_1833,In_2);
and U2480 (N_2480,In_1924,In_31);
xor U2481 (N_2481,In_1777,In_1202);
nor U2482 (N_2482,In_1506,In_899);
nor U2483 (N_2483,In_681,In_1428);
nand U2484 (N_2484,In_1094,In_847);
nor U2485 (N_2485,In_844,In_1649);
nor U2486 (N_2486,In_305,In_1874);
and U2487 (N_2487,In_309,In_1762);
xor U2488 (N_2488,In_1967,In_1934);
nand U2489 (N_2489,In_352,In_1810);
and U2490 (N_2490,In_2,In_648);
and U2491 (N_2491,In_1510,In_320);
nor U2492 (N_2492,In_1788,In_1328);
nand U2493 (N_2493,In_1561,In_956);
nand U2494 (N_2494,In_1909,In_1329);
nand U2495 (N_2495,In_1007,In_1544);
and U2496 (N_2496,In_226,In_1930);
nor U2497 (N_2497,In_415,In_719);
nor U2498 (N_2498,In_331,In_1326);
xor U2499 (N_2499,In_391,In_374);
and U2500 (N_2500,In_322,In_1010);
or U2501 (N_2501,In_1576,In_1729);
nor U2502 (N_2502,In_976,In_1230);
and U2503 (N_2503,In_638,In_1324);
or U2504 (N_2504,In_1651,In_665);
or U2505 (N_2505,In_1643,In_1421);
xor U2506 (N_2506,In_916,In_1397);
xnor U2507 (N_2507,In_385,In_1532);
or U2508 (N_2508,In_1652,In_1779);
nor U2509 (N_2509,In_793,In_1810);
xnor U2510 (N_2510,In_1020,In_818);
or U2511 (N_2511,In_488,In_1459);
or U2512 (N_2512,In_1659,In_1282);
and U2513 (N_2513,In_431,In_143);
and U2514 (N_2514,In_143,In_205);
xnor U2515 (N_2515,In_1364,In_1195);
or U2516 (N_2516,In_1330,In_1639);
xnor U2517 (N_2517,In_1508,In_324);
nor U2518 (N_2518,In_953,In_1003);
xnor U2519 (N_2519,In_1684,In_1989);
nand U2520 (N_2520,In_673,In_1628);
xnor U2521 (N_2521,In_586,In_582);
and U2522 (N_2522,In_1335,In_106);
nor U2523 (N_2523,In_727,In_494);
nand U2524 (N_2524,In_1014,In_1025);
nand U2525 (N_2525,In_1343,In_1822);
and U2526 (N_2526,In_579,In_1392);
and U2527 (N_2527,In_1138,In_1665);
nand U2528 (N_2528,In_161,In_496);
or U2529 (N_2529,In_8,In_67);
xnor U2530 (N_2530,In_1659,In_220);
or U2531 (N_2531,In_1639,In_328);
or U2532 (N_2532,In_344,In_1172);
and U2533 (N_2533,In_90,In_1218);
xor U2534 (N_2534,In_1261,In_1591);
xnor U2535 (N_2535,In_230,In_1740);
nor U2536 (N_2536,In_1782,In_1624);
and U2537 (N_2537,In_673,In_1480);
and U2538 (N_2538,In_474,In_1936);
nand U2539 (N_2539,In_356,In_476);
xnor U2540 (N_2540,In_1546,In_900);
and U2541 (N_2541,In_1762,In_128);
xor U2542 (N_2542,In_1367,In_1178);
or U2543 (N_2543,In_783,In_825);
xor U2544 (N_2544,In_993,In_1493);
or U2545 (N_2545,In_547,In_454);
or U2546 (N_2546,In_1273,In_6);
nor U2547 (N_2547,In_1071,In_54);
nand U2548 (N_2548,In_89,In_1480);
and U2549 (N_2549,In_1120,In_1797);
or U2550 (N_2550,In_326,In_933);
or U2551 (N_2551,In_448,In_918);
xnor U2552 (N_2552,In_1830,In_1176);
nand U2553 (N_2553,In_155,In_1815);
nor U2554 (N_2554,In_793,In_1461);
or U2555 (N_2555,In_1185,In_296);
and U2556 (N_2556,In_1789,In_573);
nand U2557 (N_2557,In_1665,In_1022);
nand U2558 (N_2558,In_1640,In_335);
nand U2559 (N_2559,In_416,In_430);
xnor U2560 (N_2560,In_107,In_56);
nand U2561 (N_2561,In_1895,In_243);
xor U2562 (N_2562,In_720,In_1661);
or U2563 (N_2563,In_163,In_1205);
and U2564 (N_2564,In_1803,In_1935);
or U2565 (N_2565,In_1690,In_1231);
or U2566 (N_2566,In_1564,In_1873);
and U2567 (N_2567,In_1235,In_869);
and U2568 (N_2568,In_1488,In_1071);
and U2569 (N_2569,In_461,In_1808);
nor U2570 (N_2570,In_650,In_1020);
xnor U2571 (N_2571,In_1273,In_1025);
xor U2572 (N_2572,In_1936,In_1940);
xor U2573 (N_2573,In_1578,In_1822);
xor U2574 (N_2574,In_547,In_1838);
nand U2575 (N_2575,In_1618,In_784);
nand U2576 (N_2576,In_1722,In_1841);
and U2577 (N_2577,In_1314,In_133);
xor U2578 (N_2578,In_818,In_1133);
nor U2579 (N_2579,In_1999,In_1580);
nor U2580 (N_2580,In_550,In_1911);
and U2581 (N_2581,In_833,In_539);
xor U2582 (N_2582,In_1612,In_1337);
xnor U2583 (N_2583,In_829,In_1885);
or U2584 (N_2584,In_1959,In_1313);
xor U2585 (N_2585,In_339,In_365);
nor U2586 (N_2586,In_219,In_940);
and U2587 (N_2587,In_1282,In_6);
xnor U2588 (N_2588,In_1785,In_432);
and U2589 (N_2589,In_961,In_181);
nand U2590 (N_2590,In_1732,In_346);
xor U2591 (N_2591,In_1409,In_1323);
or U2592 (N_2592,In_366,In_70);
and U2593 (N_2593,In_1010,In_1116);
xor U2594 (N_2594,In_347,In_662);
nor U2595 (N_2595,In_71,In_1623);
xor U2596 (N_2596,In_983,In_1099);
and U2597 (N_2597,In_345,In_1010);
or U2598 (N_2598,In_1019,In_313);
nor U2599 (N_2599,In_1625,In_135);
and U2600 (N_2600,In_170,In_346);
and U2601 (N_2601,In_1184,In_1604);
nor U2602 (N_2602,In_387,In_1342);
xor U2603 (N_2603,In_406,In_13);
nor U2604 (N_2604,In_1246,In_1478);
and U2605 (N_2605,In_726,In_1998);
nand U2606 (N_2606,In_1751,In_1818);
xnor U2607 (N_2607,In_73,In_936);
or U2608 (N_2608,In_1959,In_1474);
nand U2609 (N_2609,In_576,In_1411);
xor U2610 (N_2610,In_1137,In_419);
nor U2611 (N_2611,In_1607,In_1909);
nor U2612 (N_2612,In_165,In_1063);
xnor U2613 (N_2613,In_1644,In_510);
or U2614 (N_2614,In_1840,In_1546);
or U2615 (N_2615,In_1777,In_267);
or U2616 (N_2616,In_142,In_394);
or U2617 (N_2617,In_1554,In_1279);
or U2618 (N_2618,In_1484,In_69);
nor U2619 (N_2619,In_511,In_1179);
or U2620 (N_2620,In_485,In_1811);
xnor U2621 (N_2621,In_1415,In_850);
or U2622 (N_2622,In_425,In_833);
nor U2623 (N_2623,In_1457,In_1708);
or U2624 (N_2624,In_1996,In_165);
nor U2625 (N_2625,In_709,In_1430);
and U2626 (N_2626,In_1154,In_410);
or U2627 (N_2627,In_1147,In_598);
nor U2628 (N_2628,In_257,In_1071);
nor U2629 (N_2629,In_1564,In_706);
or U2630 (N_2630,In_1416,In_1883);
xnor U2631 (N_2631,In_1335,In_1341);
xor U2632 (N_2632,In_132,In_1767);
xnor U2633 (N_2633,In_70,In_290);
nand U2634 (N_2634,In_1085,In_1940);
nor U2635 (N_2635,In_909,In_1077);
or U2636 (N_2636,In_1455,In_1531);
xor U2637 (N_2637,In_1155,In_751);
and U2638 (N_2638,In_1270,In_196);
or U2639 (N_2639,In_1797,In_477);
nor U2640 (N_2640,In_1561,In_1848);
nor U2641 (N_2641,In_204,In_45);
and U2642 (N_2642,In_116,In_217);
xnor U2643 (N_2643,In_766,In_440);
nand U2644 (N_2644,In_681,In_1890);
or U2645 (N_2645,In_251,In_1419);
nor U2646 (N_2646,In_325,In_221);
or U2647 (N_2647,In_861,In_1198);
and U2648 (N_2648,In_1969,In_1176);
nand U2649 (N_2649,In_688,In_329);
or U2650 (N_2650,In_82,In_1585);
nor U2651 (N_2651,In_354,In_52);
or U2652 (N_2652,In_312,In_1245);
nor U2653 (N_2653,In_935,In_214);
nand U2654 (N_2654,In_651,In_52);
xnor U2655 (N_2655,In_222,In_580);
xor U2656 (N_2656,In_1796,In_1568);
or U2657 (N_2657,In_1749,In_935);
or U2658 (N_2658,In_574,In_1553);
xor U2659 (N_2659,In_799,In_604);
nor U2660 (N_2660,In_169,In_20);
xor U2661 (N_2661,In_740,In_250);
or U2662 (N_2662,In_918,In_365);
xor U2663 (N_2663,In_1186,In_1288);
xor U2664 (N_2664,In_695,In_1018);
or U2665 (N_2665,In_530,In_962);
and U2666 (N_2666,In_1408,In_102);
and U2667 (N_2667,In_1513,In_1813);
nand U2668 (N_2668,In_636,In_1152);
or U2669 (N_2669,In_94,In_162);
xor U2670 (N_2670,In_977,In_1945);
or U2671 (N_2671,In_1839,In_1432);
or U2672 (N_2672,In_1497,In_125);
nor U2673 (N_2673,In_635,In_687);
nand U2674 (N_2674,In_1190,In_777);
or U2675 (N_2675,In_34,In_506);
nand U2676 (N_2676,In_1093,In_212);
xor U2677 (N_2677,In_1292,In_1076);
nor U2678 (N_2678,In_756,In_559);
xor U2679 (N_2679,In_912,In_515);
nand U2680 (N_2680,In_1264,In_750);
xnor U2681 (N_2681,In_1157,In_1943);
and U2682 (N_2682,In_858,In_202);
or U2683 (N_2683,In_1966,In_474);
and U2684 (N_2684,In_1671,In_1484);
or U2685 (N_2685,In_366,In_1582);
or U2686 (N_2686,In_1041,In_1975);
or U2687 (N_2687,In_696,In_1133);
nor U2688 (N_2688,In_96,In_416);
or U2689 (N_2689,In_1153,In_774);
xnor U2690 (N_2690,In_1685,In_1348);
nor U2691 (N_2691,In_180,In_1730);
nor U2692 (N_2692,In_355,In_396);
and U2693 (N_2693,In_1722,In_823);
or U2694 (N_2694,In_1968,In_868);
or U2695 (N_2695,In_252,In_722);
nor U2696 (N_2696,In_1952,In_1105);
nor U2697 (N_2697,In_1149,In_1519);
xnor U2698 (N_2698,In_546,In_154);
nor U2699 (N_2699,In_1468,In_350);
xnor U2700 (N_2700,In_1046,In_632);
nand U2701 (N_2701,In_857,In_769);
nand U2702 (N_2702,In_1806,In_19);
xor U2703 (N_2703,In_1836,In_901);
xnor U2704 (N_2704,In_249,In_1023);
and U2705 (N_2705,In_283,In_1658);
or U2706 (N_2706,In_1814,In_20);
or U2707 (N_2707,In_411,In_1194);
and U2708 (N_2708,In_1076,In_1700);
or U2709 (N_2709,In_771,In_1522);
or U2710 (N_2710,In_1366,In_1342);
nand U2711 (N_2711,In_1858,In_413);
nand U2712 (N_2712,In_1032,In_305);
nand U2713 (N_2713,In_1376,In_1448);
or U2714 (N_2714,In_334,In_1038);
xor U2715 (N_2715,In_1196,In_840);
nand U2716 (N_2716,In_1212,In_217);
nand U2717 (N_2717,In_1159,In_915);
and U2718 (N_2718,In_1574,In_356);
xnor U2719 (N_2719,In_595,In_779);
and U2720 (N_2720,In_1078,In_1725);
or U2721 (N_2721,In_1129,In_583);
or U2722 (N_2722,In_1883,In_1082);
or U2723 (N_2723,In_1409,In_249);
and U2724 (N_2724,In_1562,In_1483);
or U2725 (N_2725,In_144,In_550);
and U2726 (N_2726,In_360,In_828);
xnor U2727 (N_2727,In_1182,In_404);
and U2728 (N_2728,In_337,In_121);
and U2729 (N_2729,In_1773,In_1173);
nor U2730 (N_2730,In_253,In_164);
xnor U2731 (N_2731,In_1844,In_329);
nand U2732 (N_2732,In_1237,In_1154);
xnor U2733 (N_2733,In_721,In_766);
nand U2734 (N_2734,In_684,In_1127);
nand U2735 (N_2735,In_1873,In_1915);
or U2736 (N_2736,In_1803,In_1868);
nand U2737 (N_2737,In_1601,In_1015);
nand U2738 (N_2738,In_1552,In_1928);
xor U2739 (N_2739,In_290,In_1322);
nor U2740 (N_2740,In_1278,In_1179);
nor U2741 (N_2741,In_1181,In_1948);
nor U2742 (N_2742,In_324,In_687);
or U2743 (N_2743,In_1769,In_1935);
xnor U2744 (N_2744,In_933,In_227);
and U2745 (N_2745,In_1200,In_1257);
nor U2746 (N_2746,In_1415,In_1546);
nand U2747 (N_2747,In_1008,In_327);
xor U2748 (N_2748,In_1632,In_1463);
nor U2749 (N_2749,In_1288,In_1873);
nor U2750 (N_2750,In_94,In_1042);
xor U2751 (N_2751,In_831,In_70);
and U2752 (N_2752,In_805,In_888);
nand U2753 (N_2753,In_1936,In_1283);
nor U2754 (N_2754,In_1203,In_560);
or U2755 (N_2755,In_375,In_1163);
nor U2756 (N_2756,In_389,In_464);
nand U2757 (N_2757,In_1570,In_1034);
or U2758 (N_2758,In_471,In_255);
nand U2759 (N_2759,In_1025,In_1738);
xor U2760 (N_2760,In_270,In_1148);
nand U2761 (N_2761,In_259,In_1784);
or U2762 (N_2762,In_1424,In_1135);
and U2763 (N_2763,In_943,In_1556);
xor U2764 (N_2764,In_1300,In_400);
nand U2765 (N_2765,In_1450,In_62);
nand U2766 (N_2766,In_1251,In_232);
or U2767 (N_2767,In_1973,In_1764);
nor U2768 (N_2768,In_112,In_1111);
nor U2769 (N_2769,In_370,In_1128);
nor U2770 (N_2770,In_1416,In_586);
nor U2771 (N_2771,In_1178,In_1782);
xor U2772 (N_2772,In_193,In_242);
nand U2773 (N_2773,In_1812,In_1979);
or U2774 (N_2774,In_260,In_971);
nor U2775 (N_2775,In_810,In_789);
nor U2776 (N_2776,In_545,In_4);
nand U2777 (N_2777,In_205,In_1739);
nand U2778 (N_2778,In_1301,In_150);
nand U2779 (N_2779,In_748,In_1687);
or U2780 (N_2780,In_97,In_990);
or U2781 (N_2781,In_1867,In_1099);
or U2782 (N_2782,In_820,In_576);
or U2783 (N_2783,In_1585,In_1511);
or U2784 (N_2784,In_322,In_1185);
nor U2785 (N_2785,In_1924,In_1058);
xor U2786 (N_2786,In_520,In_1748);
nand U2787 (N_2787,In_1011,In_420);
nand U2788 (N_2788,In_1125,In_1180);
nor U2789 (N_2789,In_8,In_361);
xor U2790 (N_2790,In_343,In_480);
nor U2791 (N_2791,In_53,In_752);
xnor U2792 (N_2792,In_752,In_1935);
and U2793 (N_2793,In_1459,In_108);
nor U2794 (N_2794,In_1602,In_550);
nor U2795 (N_2795,In_460,In_1707);
or U2796 (N_2796,In_839,In_1785);
nand U2797 (N_2797,In_1293,In_823);
xnor U2798 (N_2798,In_1815,In_1334);
and U2799 (N_2799,In_934,In_1075);
nand U2800 (N_2800,In_1241,In_617);
nand U2801 (N_2801,In_1613,In_211);
nor U2802 (N_2802,In_271,In_968);
or U2803 (N_2803,In_1994,In_1121);
xnor U2804 (N_2804,In_1158,In_1333);
nor U2805 (N_2805,In_920,In_1510);
nand U2806 (N_2806,In_1819,In_1597);
or U2807 (N_2807,In_588,In_738);
nor U2808 (N_2808,In_1527,In_511);
or U2809 (N_2809,In_31,In_1104);
and U2810 (N_2810,In_226,In_565);
or U2811 (N_2811,In_356,In_519);
xnor U2812 (N_2812,In_1832,In_1715);
and U2813 (N_2813,In_1985,In_1167);
nand U2814 (N_2814,In_559,In_134);
nand U2815 (N_2815,In_276,In_1375);
nand U2816 (N_2816,In_770,In_765);
nor U2817 (N_2817,In_1872,In_601);
or U2818 (N_2818,In_172,In_1278);
nand U2819 (N_2819,In_713,In_221);
nand U2820 (N_2820,In_1437,In_1417);
or U2821 (N_2821,In_1575,In_1366);
or U2822 (N_2822,In_1694,In_161);
xnor U2823 (N_2823,In_1118,In_871);
nand U2824 (N_2824,In_1278,In_501);
xnor U2825 (N_2825,In_1879,In_1937);
xor U2826 (N_2826,In_1805,In_1836);
and U2827 (N_2827,In_1118,In_626);
and U2828 (N_2828,In_1508,In_23);
and U2829 (N_2829,In_666,In_1534);
or U2830 (N_2830,In_40,In_1865);
or U2831 (N_2831,In_245,In_1360);
nand U2832 (N_2832,In_327,In_1257);
and U2833 (N_2833,In_209,In_594);
or U2834 (N_2834,In_653,In_1355);
nand U2835 (N_2835,In_108,In_1752);
and U2836 (N_2836,In_1330,In_133);
and U2837 (N_2837,In_940,In_475);
nor U2838 (N_2838,In_190,In_1671);
or U2839 (N_2839,In_216,In_803);
xor U2840 (N_2840,In_1351,In_302);
xnor U2841 (N_2841,In_1344,In_291);
nor U2842 (N_2842,In_1141,In_1457);
nor U2843 (N_2843,In_1534,In_1470);
xnor U2844 (N_2844,In_1598,In_1695);
xor U2845 (N_2845,In_1931,In_1357);
nand U2846 (N_2846,In_385,In_1921);
nor U2847 (N_2847,In_1181,In_916);
nor U2848 (N_2848,In_885,In_1719);
xor U2849 (N_2849,In_433,In_224);
and U2850 (N_2850,In_557,In_133);
and U2851 (N_2851,In_1304,In_1129);
or U2852 (N_2852,In_322,In_268);
xor U2853 (N_2853,In_1463,In_137);
or U2854 (N_2854,In_462,In_1650);
nor U2855 (N_2855,In_1077,In_685);
and U2856 (N_2856,In_1468,In_499);
or U2857 (N_2857,In_1445,In_544);
xor U2858 (N_2858,In_1744,In_1632);
xnor U2859 (N_2859,In_1756,In_1363);
nor U2860 (N_2860,In_1477,In_1171);
nor U2861 (N_2861,In_1877,In_1658);
xor U2862 (N_2862,In_1559,In_268);
nand U2863 (N_2863,In_923,In_94);
nor U2864 (N_2864,In_1797,In_1898);
nand U2865 (N_2865,In_1081,In_734);
nor U2866 (N_2866,In_770,In_1725);
nor U2867 (N_2867,In_481,In_691);
or U2868 (N_2868,In_1636,In_621);
nor U2869 (N_2869,In_391,In_723);
and U2870 (N_2870,In_1257,In_1157);
nand U2871 (N_2871,In_61,In_1039);
nor U2872 (N_2872,In_532,In_1627);
and U2873 (N_2873,In_1705,In_1382);
or U2874 (N_2874,In_1004,In_1878);
nor U2875 (N_2875,In_1765,In_1078);
or U2876 (N_2876,In_1665,In_1991);
xor U2877 (N_2877,In_1244,In_620);
or U2878 (N_2878,In_1458,In_222);
nand U2879 (N_2879,In_1393,In_185);
nor U2880 (N_2880,In_1912,In_1831);
nand U2881 (N_2881,In_915,In_816);
nand U2882 (N_2882,In_1967,In_879);
or U2883 (N_2883,In_1423,In_488);
nor U2884 (N_2884,In_1527,In_940);
and U2885 (N_2885,In_251,In_619);
nand U2886 (N_2886,In_435,In_991);
xnor U2887 (N_2887,In_1295,In_265);
nand U2888 (N_2888,In_1115,In_841);
nor U2889 (N_2889,In_139,In_301);
or U2890 (N_2890,In_1128,In_204);
nand U2891 (N_2891,In_720,In_1193);
and U2892 (N_2892,In_1761,In_844);
nor U2893 (N_2893,In_684,In_1747);
nor U2894 (N_2894,In_533,In_1059);
or U2895 (N_2895,In_798,In_1949);
and U2896 (N_2896,In_1471,In_1434);
nor U2897 (N_2897,In_1390,In_661);
xor U2898 (N_2898,In_1908,In_1586);
nand U2899 (N_2899,In_90,In_865);
and U2900 (N_2900,In_1475,In_1202);
nand U2901 (N_2901,In_1405,In_1888);
nor U2902 (N_2902,In_10,In_1984);
and U2903 (N_2903,In_1589,In_1000);
nor U2904 (N_2904,In_520,In_1067);
or U2905 (N_2905,In_464,In_46);
and U2906 (N_2906,In_1075,In_1601);
or U2907 (N_2907,In_78,In_608);
xnor U2908 (N_2908,In_1459,In_73);
nand U2909 (N_2909,In_434,In_1554);
and U2910 (N_2910,In_1344,In_1829);
or U2911 (N_2911,In_1370,In_1711);
or U2912 (N_2912,In_1778,In_1860);
nand U2913 (N_2913,In_664,In_417);
xor U2914 (N_2914,In_1384,In_1161);
and U2915 (N_2915,In_1118,In_17);
nand U2916 (N_2916,In_1790,In_850);
nand U2917 (N_2917,In_1726,In_164);
nor U2918 (N_2918,In_789,In_111);
or U2919 (N_2919,In_1423,In_1323);
nand U2920 (N_2920,In_803,In_1604);
nor U2921 (N_2921,In_1545,In_1439);
or U2922 (N_2922,In_744,In_1822);
nand U2923 (N_2923,In_292,In_1304);
nor U2924 (N_2924,In_147,In_1757);
or U2925 (N_2925,In_1715,In_1478);
or U2926 (N_2926,In_948,In_1001);
nor U2927 (N_2927,In_417,In_1364);
and U2928 (N_2928,In_365,In_568);
and U2929 (N_2929,In_1434,In_732);
or U2930 (N_2930,In_1108,In_1373);
and U2931 (N_2931,In_672,In_572);
or U2932 (N_2932,In_304,In_1021);
xor U2933 (N_2933,In_1881,In_219);
nand U2934 (N_2934,In_24,In_1897);
or U2935 (N_2935,In_1476,In_1489);
or U2936 (N_2936,In_1464,In_833);
nand U2937 (N_2937,In_68,In_262);
and U2938 (N_2938,In_28,In_224);
or U2939 (N_2939,In_56,In_1603);
nand U2940 (N_2940,In_1279,In_936);
xnor U2941 (N_2941,In_1746,In_875);
nor U2942 (N_2942,In_246,In_1093);
nand U2943 (N_2943,In_719,In_883);
or U2944 (N_2944,In_1806,In_1671);
or U2945 (N_2945,In_1150,In_1679);
and U2946 (N_2946,In_1429,In_703);
xnor U2947 (N_2947,In_822,In_1663);
xnor U2948 (N_2948,In_490,In_375);
and U2949 (N_2949,In_511,In_1890);
xnor U2950 (N_2950,In_1239,In_1574);
and U2951 (N_2951,In_1303,In_126);
or U2952 (N_2952,In_1859,In_961);
or U2953 (N_2953,In_559,In_2);
xnor U2954 (N_2954,In_1507,In_250);
xnor U2955 (N_2955,In_1912,In_1541);
nor U2956 (N_2956,In_865,In_1924);
and U2957 (N_2957,In_277,In_1996);
xnor U2958 (N_2958,In_213,In_1660);
or U2959 (N_2959,In_1976,In_1832);
or U2960 (N_2960,In_1287,In_908);
or U2961 (N_2961,In_2,In_1010);
or U2962 (N_2962,In_1342,In_294);
and U2963 (N_2963,In_1217,In_952);
or U2964 (N_2964,In_1546,In_1981);
or U2965 (N_2965,In_274,In_262);
xor U2966 (N_2966,In_229,In_122);
nand U2967 (N_2967,In_1002,In_1160);
xnor U2968 (N_2968,In_847,In_1052);
and U2969 (N_2969,In_951,In_794);
nor U2970 (N_2970,In_1231,In_201);
nand U2971 (N_2971,In_1457,In_1978);
xor U2972 (N_2972,In_1489,In_874);
or U2973 (N_2973,In_1654,In_76);
xor U2974 (N_2974,In_1006,In_566);
and U2975 (N_2975,In_1432,In_156);
xnor U2976 (N_2976,In_1593,In_1177);
or U2977 (N_2977,In_711,In_290);
nor U2978 (N_2978,In_142,In_1847);
or U2979 (N_2979,In_11,In_1219);
or U2980 (N_2980,In_1735,In_373);
xnor U2981 (N_2981,In_1408,In_950);
and U2982 (N_2982,In_259,In_545);
and U2983 (N_2983,In_1477,In_1724);
and U2984 (N_2984,In_1347,In_393);
nor U2985 (N_2985,In_290,In_1069);
or U2986 (N_2986,In_1856,In_273);
nand U2987 (N_2987,In_137,In_1177);
xor U2988 (N_2988,In_1262,In_905);
nand U2989 (N_2989,In_1854,In_729);
and U2990 (N_2990,In_876,In_410);
nand U2991 (N_2991,In_268,In_1441);
and U2992 (N_2992,In_1764,In_908);
xnor U2993 (N_2993,In_1987,In_335);
nand U2994 (N_2994,In_1040,In_1730);
or U2995 (N_2995,In_1259,In_601);
xnor U2996 (N_2996,In_1582,In_1338);
and U2997 (N_2997,In_915,In_195);
or U2998 (N_2998,In_1163,In_68);
nand U2999 (N_2999,In_1954,In_1706);
xor U3000 (N_3000,In_164,In_776);
nor U3001 (N_3001,In_1942,In_1808);
or U3002 (N_3002,In_1734,In_872);
and U3003 (N_3003,In_52,In_1311);
or U3004 (N_3004,In_1041,In_58);
and U3005 (N_3005,In_1089,In_1767);
or U3006 (N_3006,In_766,In_317);
xor U3007 (N_3007,In_716,In_53);
nor U3008 (N_3008,In_349,In_167);
nand U3009 (N_3009,In_1309,In_1058);
xor U3010 (N_3010,In_1571,In_1374);
nor U3011 (N_3011,In_1959,In_1184);
or U3012 (N_3012,In_1794,In_1110);
xnor U3013 (N_3013,In_1547,In_309);
and U3014 (N_3014,In_819,In_304);
nor U3015 (N_3015,In_1513,In_688);
xor U3016 (N_3016,In_1501,In_171);
or U3017 (N_3017,In_1231,In_1011);
nor U3018 (N_3018,In_1567,In_199);
and U3019 (N_3019,In_775,In_265);
and U3020 (N_3020,In_1671,In_521);
and U3021 (N_3021,In_1290,In_112);
nand U3022 (N_3022,In_1285,In_53);
nand U3023 (N_3023,In_150,In_900);
nor U3024 (N_3024,In_98,In_1740);
nand U3025 (N_3025,In_212,In_1064);
and U3026 (N_3026,In_1227,In_1368);
xnor U3027 (N_3027,In_1037,In_566);
xnor U3028 (N_3028,In_1649,In_638);
or U3029 (N_3029,In_611,In_417);
nand U3030 (N_3030,In_1574,In_1751);
or U3031 (N_3031,In_575,In_287);
or U3032 (N_3032,In_824,In_1675);
and U3033 (N_3033,In_1216,In_1715);
and U3034 (N_3034,In_960,In_605);
xnor U3035 (N_3035,In_1349,In_64);
or U3036 (N_3036,In_498,In_1144);
nor U3037 (N_3037,In_660,In_1484);
xnor U3038 (N_3038,In_200,In_1947);
nor U3039 (N_3039,In_1395,In_1344);
nand U3040 (N_3040,In_508,In_1413);
and U3041 (N_3041,In_520,In_652);
and U3042 (N_3042,In_222,In_90);
xnor U3043 (N_3043,In_1171,In_702);
nand U3044 (N_3044,In_139,In_1611);
nand U3045 (N_3045,In_413,In_1044);
or U3046 (N_3046,In_1175,In_1051);
xnor U3047 (N_3047,In_1690,In_763);
nand U3048 (N_3048,In_856,In_383);
or U3049 (N_3049,In_1851,In_1872);
and U3050 (N_3050,In_809,In_331);
xnor U3051 (N_3051,In_935,In_290);
or U3052 (N_3052,In_507,In_1089);
nand U3053 (N_3053,In_434,In_1744);
xnor U3054 (N_3054,In_741,In_1536);
xor U3055 (N_3055,In_123,In_892);
xnor U3056 (N_3056,In_1552,In_561);
xnor U3057 (N_3057,In_364,In_204);
nand U3058 (N_3058,In_93,In_1380);
xor U3059 (N_3059,In_1123,In_620);
and U3060 (N_3060,In_1045,In_1352);
xor U3061 (N_3061,In_444,In_240);
nand U3062 (N_3062,In_1016,In_1959);
or U3063 (N_3063,In_1556,In_90);
nor U3064 (N_3064,In_1640,In_1226);
nor U3065 (N_3065,In_478,In_50);
or U3066 (N_3066,In_1468,In_1509);
and U3067 (N_3067,In_1080,In_692);
xnor U3068 (N_3068,In_1522,In_580);
nand U3069 (N_3069,In_1960,In_80);
or U3070 (N_3070,In_1252,In_610);
xnor U3071 (N_3071,In_785,In_818);
xnor U3072 (N_3072,In_1282,In_296);
or U3073 (N_3073,In_1260,In_658);
xor U3074 (N_3074,In_1605,In_700);
xor U3075 (N_3075,In_508,In_1288);
or U3076 (N_3076,In_1729,In_1511);
or U3077 (N_3077,In_1215,In_1458);
and U3078 (N_3078,In_946,In_1631);
and U3079 (N_3079,In_1083,In_305);
and U3080 (N_3080,In_1528,In_279);
or U3081 (N_3081,In_1336,In_1332);
xnor U3082 (N_3082,In_150,In_1785);
or U3083 (N_3083,In_1620,In_1962);
xnor U3084 (N_3084,In_1465,In_1497);
xor U3085 (N_3085,In_358,In_1774);
nor U3086 (N_3086,In_1064,In_1247);
and U3087 (N_3087,In_103,In_1261);
or U3088 (N_3088,In_1358,In_571);
or U3089 (N_3089,In_27,In_374);
and U3090 (N_3090,In_1794,In_871);
or U3091 (N_3091,In_1057,In_536);
nand U3092 (N_3092,In_172,In_1555);
xnor U3093 (N_3093,In_1389,In_1915);
nand U3094 (N_3094,In_1065,In_1624);
nor U3095 (N_3095,In_189,In_1744);
nand U3096 (N_3096,In_458,In_1108);
nand U3097 (N_3097,In_623,In_1551);
and U3098 (N_3098,In_722,In_1397);
and U3099 (N_3099,In_425,In_167);
and U3100 (N_3100,In_374,In_262);
and U3101 (N_3101,In_851,In_1523);
and U3102 (N_3102,In_337,In_61);
nor U3103 (N_3103,In_1290,In_348);
nor U3104 (N_3104,In_824,In_1148);
xnor U3105 (N_3105,In_1142,In_54);
nor U3106 (N_3106,In_991,In_1651);
xnor U3107 (N_3107,In_1839,In_698);
nor U3108 (N_3108,In_981,In_1892);
xnor U3109 (N_3109,In_1884,In_1679);
xor U3110 (N_3110,In_1095,In_767);
nor U3111 (N_3111,In_586,In_1686);
or U3112 (N_3112,In_742,In_237);
xor U3113 (N_3113,In_711,In_32);
nor U3114 (N_3114,In_1766,In_114);
nand U3115 (N_3115,In_747,In_1140);
nor U3116 (N_3116,In_1335,In_776);
and U3117 (N_3117,In_856,In_585);
nand U3118 (N_3118,In_1813,In_392);
nor U3119 (N_3119,In_1799,In_1750);
and U3120 (N_3120,In_946,In_1269);
nand U3121 (N_3121,In_705,In_1076);
nand U3122 (N_3122,In_852,In_1519);
or U3123 (N_3123,In_735,In_915);
nor U3124 (N_3124,In_1001,In_1911);
xor U3125 (N_3125,In_414,In_1132);
and U3126 (N_3126,In_1346,In_601);
xnor U3127 (N_3127,In_230,In_6);
xnor U3128 (N_3128,In_1729,In_1997);
nor U3129 (N_3129,In_1534,In_281);
and U3130 (N_3130,In_595,In_1706);
nand U3131 (N_3131,In_597,In_997);
or U3132 (N_3132,In_585,In_1217);
and U3133 (N_3133,In_1049,In_1846);
or U3134 (N_3134,In_603,In_178);
or U3135 (N_3135,In_1353,In_921);
nand U3136 (N_3136,In_688,In_1267);
xnor U3137 (N_3137,In_504,In_1001);
or U3138 (N_3138,In_666,In_1074);
or U3139 (N_3139,In_32,In_1087);
nand U3140 (N_3140,In_214,In_1534);
xnor U3141 (N_3141,In_1960,In_1734);
nand U3142 (N_3142,In_1127,In_644);
xor U3143 (N_3143,In_1255,In_1024);
and U3144 (N_3144,In_1116,In_1274);
nand U3145 (N_3145,In_355,In_1410);
nand U3146 (N_3146,In_816,In_181);
nor U3147 (N_3147,In_612,In_1825);
or U3148 (N_3148,In_1306,In_1957);
and U3149 (N_3149,In_548,In_879);
nand U3150 (N_3150,In_1323,In_691);
and U3151 (N_3151,In_1100,In_630);
or U3152 (N_3152,In_1028,In_638);
or U3153 (N_3153,In_1377,In_1657);
nor U3154 (N_3154,In_1112,In_906);
and U3155 (N_3155,In_1633,In_1832);
nor U3156 (N_3156,In_538,In_1784);
nor U3157 (N_3157,In_559,In_1119);
or U3158 (N_3158,In_1013,In_849);
xor U3159 (N_3159,In_430,In_1698);
xor U3160 (N_3160,In_546,In_507);
and U3161 (N_3161,In_967,In_1775);
xor U3162 (N_3162,In_265,In_723);
nor U3163 (N_3163,In_643,In_101);
and U3164 (N_3164,In_651,In_767);
xor U3165 (N_3165,In_927,In_1383);
xnor U3166 (N_3166,In_1657,In_1373);
xor U3167 (N_3167,In_1231,In_646);
and U3168 (N_3168,In_41,In_1135);
xor U3169 (N_3169,In_1418,In_1882);
nor U3170 (N_3170,In_1833,In_965);
and U3171 (N_3171,In_1367,In_435);
nor U3172 (N_3172,In_1669,In_1477);
and U3173 (N_3173,In_710,In_951);
or U3174 (N_3174,In_1875,In_192);
nand U3175 (N_3175,In_587,In_74);
and U3176 (N_3176,In_889,In_236);
or U3177 (N_3177,In_664,In_185);
and U3178 (N_3178,In_281,In_850);
nor U3179 (N_3179,In_1726,In_1142);
xor U3180 (N_3180,In_1700,In_1783);
nor U3181 (N_3181,In_1727,In_201);
nand U3182 (N_3182,In_1063,In_575);
nor U3183 (N_3183,In_936,In_1928);
nor U3184 (N_3184,In_1128,In_1876);
xor U3185 (N_3185,In_1968,In_645);
nand U3186 (N_3186,In_222,In_586);
and U3187 (N_3187,In_101,In_128);
and U3188 (N_3188,In_247,In_1835);
nand U3189 (N_3189,In_662,In_893);
or U3190 (N_3190,In_1706,In_1157);
nor U3191 (N_3191,In_559,In_384);
or U3192 (N_3192,In_562,In_389);
or U3193 (N_3193,In_19,In_898);
and U3194 (N_3194,In_411,In_1386);
nor U3195 (N_3195,In_34,In_1915);
or U3196 (N_3196,In_1330,In_1873);
and U3197 (N_3197,In_831,In_957);
xnor U3198 (N_3198,In_1852,In_1718);
or U3199 (N_3199,In_562,In_475);
xnor U3200 (N_3200,In_1356,In_53);
and U3201 (N_3201,In_216,In_1071);
xor U3202 (N_3202,In_1868,In_1408);
and U3203 (N_3203,In_391,In_90);
and U3204 (N_3204,In_1777,In_731);
and U3205 (N_3205,In_981,In_1479);
and U3206 (N_3206,In_626,In_199);
nand U3207 (N_3207,In_683,In_1261);
nand U3208 (N_3208,In_69,In_289);
nand U3209 (N_3209,In_435,In_1947);
nor U3210 (N_3210,In_209,In_1048);
xnor U3211 (N_3211,In_1958,In_1279);
nor U3212 (N_3212,In_462,In_282);
and U3213 (N_3213,In_366,In_113);
and U3214 (N_3214,In_1694,In_511);
nand U3215 (N_3215,In_1044,In_1306);
xor U3216 (N_3216,In_1489,In_1134);
nor U3217 (N_3217,In_1332,In_1501);
nand U3218 (N_3218,In_173,In_739);
or U3219 (N_3219,In_1318,In_516);
and U3220 (N_3220,In_681,In_1699);
nand U3221 (N_3221,In_1179,In_902);
nand U3222 (N_3222,In_1058,In_197);
nand U3223 (N_3223,In_1477,In_1612);
or U3224 (N_3224,In_368,In_1607);
nand U3225 (N_3225,In_45,In_793);
nand U3226 (N_3226,In_581,In_1896);
or U3227 (N_3227,In_1034,In_665);
nand U3228 (N_3228,In_569,In_1267);
xnor U3229 (N_3229,In_1113,In_751);
xor U3230 (N_3230,In_1755,In_806);
or U3231 (N_3231,In_58,In_1753);
and U3232 (N_3232,In_1448,In_1752);
xnor U3233 (N_3233,In_442,In_454);
nand U3234 (N_3234,In_478,In_1847);
or U3235 (N_3235,In_1846,In_807);
nor U3236 (N_3236,In_846,In_567);
or U3237 (N_3237,In_1002,In_1332);
nand U3238 (N_3238,In_934,In_1969);
and U3239 (N_3239,In_1673,In_1296);
xnor U3240 (N_3240,In_746,In_1644);
nand U3241 (N_3241,In_669,In_436);
and U3242 (N_3242,In_150,In_561);
or U3243 (N_3243,In_1740,In_1745);
nand U3244 (N_3244,In_875,In_732);
and U3245 (N_3245,In_864,In_58);
nor U3246 (N_3246,In_563,In_1846);
xor U3247 (N_3247,In_1037,In_1714);
nor U3248 (N_3248,In_376,In_1741);
nand U3249 (N_3249,In_18,In_144);
and U3250 (N_3250,In_676,In_986);
nor U3251 (N_3251,In_640,In_894);
nand U3252 (N_3252,In_455,In_350);
nor U3253 (N_3253,In_33,In_1615);
nand U3254 (N_3254,In_1899,In_1802);
xnor U3255 (N_3255,In_185,In_1418);
nand U3256 (N_3256,In_114,In_166);
xor U3257 (N_3257,In_1143,In_1504);
xor U3258 (N_3258,In_1732,In_732);
xor U3259 (N_3259,In_624,In_1344);
and U3260 (N_3260,In_931,In_919);
xor U3261 (N_3261,In_1392,In_1826);
nand U3262 (N_3262,In_1094,In_1225);
or U3263 (N_3263,In_1053,In_64);
nor U3264 (N_3264,In_590,In_1961);
and U3265 (N_3265,In_1533,In_1724);
or U3266 (N_3266,In_1270,In_746);
nor U3267 (N_3267,In_1813,In_891);
nand U3268 (N_3268,In_666,In_234);
nand U3269 (N_3269,In_882,In_1887);
xnor U3270 (N_3270,In_293,In_715);
nor U3271 (N_3271,In_456,In_1291);
or U3272 (N_3272,In_1484,In_1331);
xnor U3273 (N_3273,In_557,In_1806);
and U3274 (N_3274,In_1134,In_1224);
and U3275 (N_3275,In_1468,In_1352);
nand U3276 (N_3276,In_902,In_879);
or U3277 (N_3277,In_966,In_760);
xnor U3278 (N_3278,In_7,In_572);
xnor U3279 (N_3279,In_1132,In_1900);
xor U3280 (N_3280,In_470,In_116);
xor U3281 (N_3281,In_812,In_1323);
nand U3282 (N_3282,In_1418,In_248);
nand U3283 (N_3283,In_489,In_412);
and U3284 (N_3284,In_1836,In_1832);
or U3285 (N_3285,In_128,In_1531);
or U3286 (N_3286,In_993,In_541);
nor U3287 (N_3287,In_820,In_1172);
and U3288 (N_3288,In_1153,In_377);
or U3289 (N_3289,In_989,In_1687);
nand U3290 (N_3290,In_1374,In_623);
or U3291 (N_3291,In_1638,In_1285);
nand U3292 (N_3292,In_569,In_950);
or U3293 (N_3293,In_948,In_56);
nand U3294 (N_3294,In_902,In_1897);
or U3295 (N_3295,In_305,In_402);
xor U3296 (N_3296,In_1816,In_926);
nand U3297 (N_3297,In_812,In_1282);
nand U3298 (N_3298,In_217,In_1897);
and U3299 (N_3299,In_1983,In_829);
xnor U3300 (N_3300,In_1718,In_186);
and U3301 (N_3301,In_990,In_1565);
nor U3302 (N_3302,In_1309,In_1645);
and U3303 (N_3303,In_1585,In_1258);
nand U3304 (N_3304,In_1641,In_1107);
and U3305 (N_3305,In_101,In_1806);
nand U3306 (N_3306,In_995,In_812);
nor U3307 (N_3307,In_869,In_1013);
and U3308 (N_3308,In_1063,In_1825);
or U3309 (N_3309,In_1408,In_6);
and U3310 (N_3310,In_708,In_1922);
and U3311 (N_3311,In_1814,In_1682);
xnor U3312 (N_3312,In_219,In_1876);
nor U3313 (N_3313,In_981,In_1104);
or U3314 (N_3314,In_1042,In_1827);
and U3315 (N_3315,In_1772,In_131);
and U3316 (N_3316,In_709,In_1040);
nor U3317 (N_3317,In_190,In_1267);
nand U3318 (N_3318,In_1744,In_1302);
nand U3319 (N_3319,In_1338,In_899);
or U3320 (N_3320,In_492,In_365);
nor U3321 (N_3321,In_137,In_123);
xnor U3322 (N_3322,In_634,In_1683);
xor U3323 (N_3323,In_809,In_271);
xor U3324 (N_3324,In_739,In_1835);
xor U3325 (N_3325,In_379,In_1558);
nand U3326 (N_3326,In_425,In_1111);
or U3327 (N_3327,In_1027,In_1129);
xor U3328 (N_3328,In_778,In_818);
nor U3329 (N_3329,In_1234,In_1034);
nand U3330 (N_3330,In_957,In_1551);
nand U3331 (N_3331,In_1900,In_1901);
and U3332 (N_3332,In_348,In_834);
nand U3333 (N_3333,In_50,In_923);
xor U3334 (N_3334,In_66,In_614);
and U3335 (N_3335,In_323,In_403);
nand U3336 (N_3336,In_1333,In_410);
nand U3337 (N_3337,In_1281,In_983);
nand U3338 (N_3338,In_1294,In_1318);
and U3339 (N_3339,In_48,In_1708);
or U3340 (N_3340,In_1701,In_1410);
xnor U3341 (N_3341,In_1626,In_890);
nor U3342 (N_3342,In_1372,In_1516);
or U3343 (N_3343,In_1963,In_1254);
and U3344 (N_3344,In_1983,In_723);
xor U3345 (N_3345,In_90,In_157);
nand U3346 (N_3346,In_47,In_1702);
and U3347 (N_3347,In_893,In_181);
nor U3348 (N_3348,In_564,In_222);
or U3349 (N_3349,In_685,In_1124);
and U3350 (N_3350,In_609,In_897);
or U3351 (N_3351,In_180,In_1734);
and U3352 (N_3352,In_1641,In_102);
and U3353 (N_3353,In_573,In_1337);
nor U3354 (N_3354,In_1336,In_1865);
and U3355 (N_3355,In_1122,In_688);
xnor U3356 (N_3356,In_1403,In_1617);
xor U3357 (N_3357,In_1541,In_1102);
nand U3358 (N_3358,In_1418,In_418);
or U3359 (N_3359,In_1471,In_759);
nand U3360 (N_3360,In_481,In_773);
nor U3361 (N_3361,In_989,In_592);
xor U3362 (N_3362,In_1386,In_620);
xor U3363 (N_3363,In_165,In_1259);
nand U3364 (N_3364,In_1071,In_325);
and U3365 (N_3365,In_1750,In_783);
nand U3366 (N_3366,In_493,In_664);
nand U3367 (N_3367,In_885,In_1442);
nor U3368 (N_3368,In_685,In_1325);
and U3369 (N_3369,In_1266,In_367);
nor U3370 (N_3370,In_1579,In_1213);
xnor U3371 (N_3371,In_722,In_1941);
nor U3372 (N_3372,In_601,In_252);
or U3373 (N_3373,In_1179,In_1632);
xnor U3374 (N_3374,In_1050,In_1197);
nor U3375 (N_3375,In_312,In_1657);
and U3376 (N_3376,In_925,In_1224);
nand U3377 (N_3377,In_390,In_1478);
or U3378 (N_3378,In_815,In_1384);
and U3379 (N_3379,In_1007,In_1661);
nand U3380 (N_3380,In_232,In_641);
xor U3381 (N_3381,In_531,In_1592);
nor U3382 (N_3382,In_1858,In_817);
nand U3383 (N_3383,In_1528,In_269);
nor U3384 (N_3384,In_1878,In_32);
nand U3385 (N_3385,In_54,In_899);
nand U3386 (N_3386,In_174,In_870);
nor U3387 (N_3387,In_1421,In_90);
nor U3388 (N_3388,In_981,In_1449);
and U3389 (N_3389,In_173,In_1772);
or U3390 (N_3390,In_1458,In_794);
nand U3391 (N_3391,In_963,In_799);
or U3392 (N_3392,In_1349,In_607);
nand U3393 (N_3393,In_1564,In_1284);
xnor U3394 (N_3394,In_418,In_1121);
and U3395 (N_3395,In_1464,In_7);
and U3396 (N_3396,In_972,In_1459);
and U3397 (N_3397,In_678,In_1306);
xor U3398 (N_3398,In_502,In_627);
and U3399 (N_3399,In_1404,In_121);
or U3400 (N_3400,In_892,In_1989);
nor U3401 (N_3401,In_1539,In_417);
or U3402 (N_3402,In_1653,In_92);
nand U3403 (N_3403,In_1962,In_193);
xnor U3404 (N_3404,In_1138,In_918);
nand U3405 (N_3405,In_1687,In_15);
nor U3406 (N_3406,In_1646,In_1630);
nor U3407 (N_3407,In_1197,In_1225);
nor U3408 (N_3408,In_163,In_580);
xor U3409 (N_3409,In_1577,In_826);
or U3410 (N_3410,In_1540,In_1020);
or U3411 (N_3411,In_1614,In_503);
xnor U3412 (N_3412,In_1234,In_1600);
xnor U3413 (N_3413,In_1945,In_1238);
xnor U3414 (N_3414,In_247,In_659);
nand U3415 (N_3415,In_1971,In_288);
xor U3416 (N_3416,In_312,In_436);
xor U3417 (N_3417,In_317,In_1000);
xor U3418 (N_3418,In_1907,In_786);
nor U3419 (N_3419,In_1834,In_579);
xnor U3420 (N_3420,In_65,In_1);
nand U3421 (N_3421,In_1726,In_371);
and U3422 (N_3422,In_1790,In_1453);
nand U3423 (N_3423,In_569,In_1672);
or U3424 (N_3424,In_1825,In_1584);
nand U3425 (N_3425,In_1825,In_1034);
or U3426 (N_3426,In_1432,In_375);
or U3427 (N_3427,In_1698,In_456);
nor U3428 (N_3428,In_210,In_1345);
nand U3429 (N_3429,In_1306,In_1357);
nor U3430 (N_3430,In_647,In_1052);
nand U3431 (N_3431,In_1121,In_663);
nor U3432 (N_3432,In_1205,In_491);
and U3433 (N_3433,In_1632,In_1228);
nor U3434 (N_3434,In_1058,In_600);
xor U3435 (N_3435,In_714,In_116);
or U3436 (N_3436,In_898,In_1166);
and U3437 (N_3437,In_1724,In_751);
nand U3438 (N_3438,In_374,In_1695);
nor U3439 (N_3439,In_1264,In_1250);
or U3440 (N_3440,In_611,In_734);
xor U3441 (N_3441,In_1271,In_271);
nand U3442 (N_3442,In_839,In_1494);
nand U3443 (N_3443,In_54,In_586);
or U3444 (N_3444,In_1374,In_536);
and U3445 (N_3445,In_1125,In_833);
xor U3446 (N_3446,In_1621,In_1596);
and U3447 (N_3447,In_373,In_408);
and U3448 (N_3448,In_610,In_1566);
nand U3449 (N_3449,In_1861,In_1081);
and U3450 (N_3450,In_1493,In_1085);
nand U3451 (N_3451,In_1646,In_962);
xor U3452 (N_3452,In_1065,In_1658);
nor U3453 (N_3453,In_1916,In_225);
xor U3454 (N_3454,In_967,In_1);
and U3455 (N_3455,In_1486,In_1435);
xor U3456 (N_3456,In_1950,In_128);
and U3457 (N_3457,In_405,In_471);
and U3458 (N_3458,In_1127,In_1655);
nor U3459 (N_3459,In_483,In_1584);
and U3460 (N_3460,In_1709,In_1572);
nand U3461 (N_3461,In_891,In_493);
nor U3462 (N_3462,In_267,In_1532);
nand U3463 (N_3463,In_498,In_143);
nand U3464 (N_3464,In_1662,In_1388);
nor U3465 (N_3465,In_1415,In_466);
nand U3466 (N_3466,In_562,In_252);
and U3467 (N_3467,In_501,In_631);
and U3468 (N_3468,In_597,In_871);
nor U3469 (N_3469,In_1067,In_784);
nor U3470 (N_3470,In_1464,In_109);
nand U3471 (N_3471,In_666,In_1374);
or U3472 (N_3472,In_96,In_1264);
and U3473 (N_3473,In_135,In_602);
nor U3474 (N_3474,In_1492,In_1480);
and U3475 (N_3475,In_1358,In_439);
or U3476 (N_3476,In_296,In_1011);
or U3477 (N_3477,In_1093,In_1899);
xnor U3478 (N_3478,In_279,In_1911);
nand U3479 (N_3479,In_297,In_1665);
nor U3480 (N_3480,In_1481,In_797);
nand U3481 (N_3481,In_1653,In_897);
nand U3482 (N_3482,In_1167,In_1596);
or U3483 (N_3483,In_560,In_936);
nor U3484 (N_3484,In_199,In_3);
nor U3485 (N_3485,In_1088,In_1727);
and U3486 (N_3486,In_1755,In_650);
xor U3487 (N_3487,In_1172,In_7);
nor U3488 (N_3488,In_403,In_220);
or U3489 (N_3489,In_1290,In_614);
nand U3490 (N_3490,In_901,In_1037);
and U3491 (N_3491,In_652,In_1125);
or U3492 (N_3492,In_1937,In_381);
and U3493 (N_3493,In_1300,In_742);
and U3494 (N_3494,In_1533,In_175);
or U3495 (N_3495,In_251,In_921);
xnor U3496 (N_3496,In_1008,In_638);
nand U3497 (N_3497,In_1678,In_511);
nor U3498 (N_3498,In_1812,In_1946);
nand U3499 (N_3499,In_630,In_1745);
or U3500 (N_3500,In_1255,In_206);
nand U3501 (N_3501,In_1651,In_571);
nor U3502 (N_3502,In_1404,In_1143);
or U3503 (N_3503,In_1033,In_1541);
xnor U3504 (N_3504,In_776,In_275);
and U3505 (N_3505,In_506,In_1146);
xnor U3506 (N_3506,In_514,In_21);
nor U3507 (N_3507,In_0,In_596);
nor U3508 (N_3508,In_72,In_600);
or U3509 (N_3509,In_1172,In_971);
xor U3510 (N_3510,In_1520,In_93);
nand U3511 (N_3511,In_136,In_729);
or U3512 (N_3512,In_591,In_220);
nand U3513 (N_3513,In_857,In_838);
nor U3514 (N_3514,In_1927,In_1378);
xor U3515 (N_3515,In_1093,In_294);
nand U3516 (N_3516,In_64,In_1006);
or U3517 (N_3517,In_933,In_381);
or U3518 (N_3518,In_366,In_1044);
nor U3519 (N_3519,In_1102,In_1743);
nand U3520 (N_3520,In_1827,In_841);
xor U3521 (N_3521,In_1348,In_1644);
nand U3522 (N_3522,In_1747,In_937);
xor U3523 (N_3523,In_1879,In_1966);
or U3524 (N_3524,In_1913,In_1612);
or U3525 (N_3525,In_1854,In_1166);
and U3526 (N_3526,In_679,In_1220);
and U3527 (N_3527,In_977,In_1228);
nor U3528 (N_3528,In_1319,In_301);
or U3529 (N_3529,In_980,In_419);
nand U3530 (N_3530,In_579,In_1402);
or U3531 (N_3531,In_1852,In_833);
xor U3532 (N_3532,In_1844,In_662);
nor U3533 (N_3533,In_773,In_1314);
nand U3534 (N_3534,In_1905,In_1214);
xor U3535 (N_3535,In_1261,In_1624);
xnor U3536 (N_3536,In_1219,In_452);
nand U3537 (N_3537,In_1109,In_611);
and U3538 (N_3538,In_1564,In_564);
and U3539 (N_3539,In_767,In_1271);
or U3540 (N_3540,In_693,In_1879);
xnor U3541 (N_3541,In_1165,In_1671);
and U3542 (N_3542,In_647,In_777);
nor U3543 (N_3543,In_253,In_1805);
and U3544 (N_3544,In_1141,In_571);
and U3545 (N_3545,In_62,In_1900);
xor U3546 (N_3546,In_1756,In_552);
or U3547 (N_3547,In_1377,In_245);
and U3548 (N_3548,In_694,In_653);
nor U3549 (N_3549,In_537,In_1935);
and U3550 (N_3550,In_441,In_590);
nand U3551 (N_3551,In_1866,In_617);
nor U3552 (N_3552,In_1025,In_1544);
xnor U3553 (N_3553,In_273,In_1242);
xor U3554 (N_3554,In_979,In_1728);
xor U3555 (N_3555,In_637,In_1106);
nand U3556 (N_3556,In_1594,In_1203);
or U3557 (N_3557,In_1313,In_1586);
xnor U3558 (N_3558,In_1219,In_1700);
xnor U3559 (N_3559,In_1053,In_355);
xor U3560 (N_3560,In_790,In_681);
and U3561 (N_3561,In_926,In_883);
and U3562 (N_3562,In_1601,In_411);
nand U3563 (N_3563,In_1164,In_1523);
xor U3564 (N_3564,In_1660,In_1428);
or U3565 (N_3565,In_279,In_1829);
nor U3566 (N_3566,In_1381,In_1331);
nor U3567 (N_3567,In_69,In_367);
or U3568 (N_3568,In_1123,In_743);
and U3569 (N_3569,In_1702,In_938);
nor U3570 (N_3570,In_216,In_1053);
nor U3571 (N_3571,In_1409,In_1601);
and U3572 (N_3572,In_856,In_360);
xor U3573 (N_3573,In_727,In_544);
nor U3574 (N_3574,In_1849,In_1048);
xnor U3575 (N_3575,In_680,In_1551);
nand U3576 (N_3576,In_1636,In_286);
xor U3577 (N_3577,In_1405,In_1751);
and U3578 (N_3578,In_1604,In_1139);
nor U3579 (N_3579,In_478,In_1022);
xnor U3580 (N_3580,In_800,In_1452);
or U3581 (N_3581,In_374,In_62);
nand U3582 (N_3582,In_1804,In_106);
xor U3583 (N_3583,In_1708,In_1505);
nand U3584 (N_3584,In_1619,In_1070);
or U3585 (N_3585,In_1595,In_1170);
nor U3586 (N_3586,In_1916,In_937);
nand U3587 (N_3587,In_1305,In_253);
nand U3588 (N_3588,In_417,In_1975);
nand U3589 (N_3589,In_1609,In_984);
nand U3590 (N_3590,In_1243,In_1321);
or U3591 (N_3591,In_644,In_1955);
or U3592 (N_3592,In_1684,In_805);
and U3593 (N_3593,In_1384,In_180);
nor U3594 (N_3594,In_641,In_768);
nor U3595 (N_3595,In_99,In_1028);
nand U3596 (N_3596,In_1913,In_977);
xor U3597 (N_3597,In_1672,In_1960);
and U3598 (N_3598,In_45,In_1341);
or U3599 (N_3599,In_1618,In_186);
and U3600 (N_3600,In_715,In_708);
xor U3601 (N_3601,In_1396,In_1277);
and U3602 (N_3602,In_1177,In_418);
xor U3603 (N_3603,In_761,In_838);
xor U3604 (N_3604,In_796,In_1484);
nor U3605 (N_3605,In_1422,In_467);
xor U3606 (N_3606,In_1357,In_284);
and U3607 (N_3607,In_733,In_1304);
or U3608 (N_3608,In_898,In_910);
xor U3609 (N_3609,In_772,In_475);
and U3610 (N_3610,In_1741,In_629);
nor U3611 (N_3611,In_393,In_845);
nand U3612 (N_3612,In_444,In_1403);
nand U3613 (N_3613,In_1217,In_11);
or U3614 (N_3614,In_1775,In_1926);
xor U3615 (N_3615,In_1458,In_10);
and U3616 (N_3616,In_1025,In_69);
or U3617 (N_3617,In_41,In_694);
and U3618 (N_3618,In_1848,In_1894);
nor U3619 (N_3619,In_569,In_196);
xnor U3620 (N_3620,In_253,In_1067);
nand U3621 (N_3621,In_635,In_709);
xor U3622 (N_3622,In_1126,In_345);
and U3623 (N_3623,In_671,In_378);
nor U3624 (N_3624,In_1745,In_389);
xnor U3625 (N_3625,In_621,In_1664);
xnor U3626 (N_3626,In_853,In_1190);
xor U3627 (N_3627,In_955,In_1167);
or U3628 (N_3628,In_1968,In_343);
nand U3629 (N_3629,In_25,In_1590);
nor U3630 (N_3630,In_1803,In_1464);
and U3631 (N_3631,In_126,In_564);
nor U3632 (N_3632,In_1692,In_1071);
or U3633 (N_3633,In_487,In_1055);
nor U3634 (N_3634,In_1837,In_1691);
and U3635 (N_3635,In_1235,In_700);
or U3636 (N_3636,In_1416,In_937);
xor U3637 (N_3637,In_1045,In_1820);
and U3638 (N_3638,In_1023,In_1652);
or U3639 (N_3639,In_759,In_463);
nor U3640 (N_3640,In_1261,In_478);
and U3641 (N_3641,In_1854,In_1436);
or U3642 (N_3642,In_1412,In_129);
or U3643 (N_3643,In_566,In_1010);
or U3644 (N_3644,In_344,In_181);
and U3645 (N_3645,In_959,In_222);
nor U3646 (N_3646,In_1957,In_197);
and U3647 (N_3647,In_277,In_91);
and U3648 (N_3648,In_1169,In_444);
nor U3649 (N_3649,In_1620,In_293);
nand U3650 (N_3650,In_1516,In_1758);
xor U3651 (N_3651,In_1490,In_1807);
and U3652 (N_3652,In_867,In_589);
or U3653 (N_3653,In_1320,In_364);
nor U3654 (N_3654,In_1002,In_902);
nor U3655 (N_3655,In_427,In_1145);
and U3656 (N_3656,In_1491,In_1969);
nand U3657 (N_3657,In_859,In_1373);
or U3658 (N_3658,In_1275,In_1969);
nor U3659 (N_3659,In_36,In_1685);
nor U3660 (N_3660,In_637,In_1723);
nor U3661 (N_3661,In_510,In_232);
and U3662 (N_3662,In_655,In_139);
xor U3663 (N_3663,In_486,In_149);
nand U3664 (N_3664,In_495,In_1252);
or U3665 (N_3665,In_960,In_1381);
xnor U3666 (N_3666,In_583,In_1518);
or U3667 (N_3667,In_621,In_1837);
or U3668 (N_3668,In_1104,In_251);
nand U3669 (N_3669,In_973,In_800);
nor U3670 (N_3670,In_329,In_379);
nand U3671 (N_3671,In_1657,In_1554);
nand U3672 (N_3672,In_1311,In_976);
xor U3673 (N_3673,In_950,In_369);
nand U3674 (N_3674,In_1642,In_1636);
xor U3675 (N_3675,In_1750,In_160);
xor U3676 (N_3676,In_1404,In_1035);
xor U3677 (N_3677,In_928,In_684);
nor U3678 (N_3678,In_1310,In_236);
or U3679 (N_3679,In_1939,In_309);
xor U3680 (N_3680,In_498,In_977);
nand U3681 (N_3681,In_1863,In_1175);
and U3682 (N_3682,In_1969,In_358);
and U3683 (N_3683,In_1425,In_565);
and U3684 (N_3684,In_1339,In_500);
nor U3685 (N_3685,In_426,In_1348);
xor U3686 (N_3686,In_904,In_176);
nor U3687 (N_3687,In_1491,In_1106);
or U3688 (N_3688,In_1419,In_1329);
or U3689 (N_3689,In_1431,In_1886);
nor U3690 (N_3690,In_1241,In_82);
and U3691 (N_3691,In_285,In_1422);
or U3692 (N_3692,In_262,In_1194);
or U3693 (N_3693,In_627,In_1198);
nor U3694 (N_3694,In_568,In_1850);
nand U3695 (N_3695,In_1956,In_1181);
nor U3696 (N_3696,In_1100,In_1233);
xnor U3697 (N_3697,In_1653,In_1352);
nand U3698 (N_3698,In_1434,In_1409);
nand U3699 (N_3699,In_1745,In_1058);
nor U3700 (N_3700,In_1389,In_1337);
and U3701 (N_3701,In_1703,In_1627);
or U3702 (N_3702,In_1988,In_45);
or U3703 (N_3703,In_559,In_1634);
xor U3704 (N_3704,In_1113,In_702);
nor U3705 (N_3705,In_1854,In_1986);
nor U3706 (N_3706,In_1111,In_99);
nor U3707 (N_3707,In_546,In_745);
or U3708 (N_3708,In_195,In_1440);
or U3709 (N_3709,In_287,In_1041);
xnor U3710 (N_3710,In_1181,In_1721);
xnor U3711 (N_3711,In_1033,In_57);
and U3712 (N_3712,In_1446,In_1641);
nand U3713 (N_3713,In_1096,In_1067);
or U3714 (N_3714,In_471,In_834);
nor U3715 (N_3715,In_1610,In_17);
nor U3716 (N_3716,In_1777,In_921);
xnor U3717 (N_3717,In_756,In_95);
and U3718 (N_3718,In_838,In_20);
nand U3719 (N_3719,In_606,In_1318);
nor U3720 (N_3720,In_1142,In_1221);
nand U3721 (N_3721,In_1826,In_792);
xor U3722 (N_3722,In_1826,In_391);
xor U3723 (N_3723,In_251,In_230);
nand U3724 (N_3724,In_1312,In_1110);
xnor U3725 (N_3725,In_77,In_1799);
nand U3726 (N_3726,In_741,In_677);
nand U3727 (N_3727,In_1036,In_850);
nand U3728 (N_3728,In_143,In_80);
nand U3729 (N_3729,In_1747,In_1676);
nand U3730 (N_3730,In_1159,In_924);
xnor U3731 (N_3731,In_1338,In_809);
and U3732 (N_3732,In_307,In_827);
or U3733 (N_3733,In_419,In_1325);
nand U3734 (N_3734,In_1495,In_23);
nor U3735 (N_3735,In_542,In_1243);
or U3736 (N_3736,In_1951,In_345);
nor U3737 (N_3737,In_1526,In_1845);
and U3738 (N_3738,In_1117,In_612);
or U3739 (N_3739,In_1352,In_1886);
nor U3740 (N_3740,In_1989,In_395);
xnor U3741 (N_3741,In_1292,In_513);
and U3742 (N_3742,In_1361,In_725);
or U3743 (N_3743,In_1494,In_1010);
and U3744 (N_3744,In_118,In_621);
nand U3745 (N_3745,In_981,In_315);
xnor U3746 (N_3746,In_1102,In_897);
or U3747 (N_3747,In_1554,In_1391);
xor U3748 (N_3748,In_1811,In_1177);
or U3749 (N_3749,In_1002,In_1317);
nand U3750 (N_3750,In_95,In_985);
and U3751 (N_3751,In_160,In_51);
and U3752 (N_3752,In_1214,In_1067);
nor U3753 (N_3753,In_1609,In_412);
nor U3754 (N_3754,In_239,In_858);
and U3755 (N_3755,In_1985,In_1215);
nor U3756 (N_3756,In_1886,In_1961);
nand U3757 (N_3757,In_579,In_847);
xor U3758 (N_3758,In_886,In_1454);
or U3759 (N_3759,In_1451,In_747);
xor U3760 (N_3760,In_1338,In_1659);
nand U3761 (N_3761,In_1308,In_983);
xnor U3762 (N_3762,In_230,In_680);
or U3763 (N_3763,In_1288,In_1430);
nor U3764 (N_3764,In_1645,In_1723);
or U3765 (N_3765,In_808,In_772);
xnor U3766 (N_3766,In_1756,In_262);
or U3767 (N_3767,In_1706,In_132);
and U3768 (N_3768,In_931,In_808);
or U3769 (N_3769,In_867,In_1489);
or U3770 (N_3770,In_464,In_163);
or U3771 (N_3771,In_828,In_219);
or U3772 (N_3772,In_1511,In_1842);
nand U3773 (N_3773,In_1705,In_647);
xnor U3774 (N_3774,In_1902,In_153);
nand U3775 (N_3775,In_1723,In_852);
xor U3776 (N_3776,In_1989,In_1294);
xnor U3777 (N_3777,In_565,In_277);
xnor U3778 (N_3778,In_1711,In_860);
nor U3779 (N_3779,In_288,In_1099);
nand U3780 (N_3780,In_90,In_1790);
nor U3781 (N_3781,In_1521,In_1634);
nand U3782 (N_3782,In_1883,In_838);
or U3783 (N_3783,In_1277,In_719);
xor U3784 (N_3784,In_460,In_1724);
or U3785 (N_3785,In_833,In_691);
nand U3786 (N_3786,In_456,In_1405);
nand U3787 (N_3787,In_698,In_260);
nor U3788 (N_3788,In_1130,In_1368);
nor U3789 (N_3789,In_1947,In_1326);
nor U3790 (N_3790,In_965,In_1114);
nor U3791 (N_3791,In_1319,In_1976);
or U3792 (N_3792,In_307,In_655);
nor U3793 (N_3793,In_1041,In_1414);
nor U3794 (N_3794,In_1207,In_1245);
nand U3795 (N_3795,In_1135,In_1744);
nand U3796 (N_3796,In_1696,In_596);
and U3797 (N_3797,In_140,In_371);
nor U3798 (N_3798,In_748,In_1208);
nand U3799 (N_3799,In_414,In_714);
nor U3800 (N_3800,In_1045,In_900);
nor U3801 (N_3801,In_1780,In_333);
nor U3802 (N_3802,In_1860,In_1463);
nand U3803 (N_3803,In_1233,In_42);
nor U3804 (N_3804,In_1451,In_1244);
nand U3805 (N_3805,In_398,In_553);
or U3806 (N_3806,In_1413,In_1158);
or U3807 (N_3807,In_1396,In_1993);
xor U3808 (N_3808,In_1327,In_839);
xor U3809 (N_3809,In_1121,In_475);
or U3810 (N_3810,In_189,In_1183);
nor U3811 (N_3811,In_1348,In_111);
nor U3812 (N_3812,In_1892,In_627);
xor U3813 (N_3813,In_361,In_686);
or U3814 (N_3814,In_553,In_937);
and U3815 (N_3815,In_336,In_1575);
nand U3816 (N_3816,In_929,In_998);
nor U3817 (N_3817,In_1348,In_1905);
and U3818 (N_3818,In_956,In_848);
nor U3819 (N_3819,In_1682,In_201);
or U3820 (N_3820,In_329,In_224);
and U3821 (N_3821,In_343,In_981);
nor U3822 (N_3822,In_442,In_492);
nor U3823 (N_3823,In_1182,In_1211);
nor U3824 (N_3824,In_1391,In_1355);
nor U3825 (N_3825,In_924,In_1433);
nand U3826 (N_3826,In_1166,In_1289);
and U3827 (N_3827,In_1707,In_1452);
xnor U3828 (N_3828,In_1780,In_632);
and U3829 (N_3829,In_861,In_78);
and U3830 (N_3830,In_817,In_1297);
nand U3831 (N_3831,In_1887,In_763);
nor U3832 (N_3832,In_442,In_1019);
nor U3833 (N_3833,In_1552,In_136);
nand U3834 (N_3834,In_595,In_323);
or U3835 (N_3835,In_835,In_1664);
nor U3836 (N_3836,In_1412,In_313);
or U3837 (N_3837,In_683,In_1448);
or U3838 (N_3838,In_1283,In_1102);
nor U3839 (N_3839,In_810,In_1562);
or U3840 (N_3840,In_1128,In_687);
nand U3841 (N_3841,In_510,In_1711);
nor U3842 (N_3842,In_319,In_439);
and U3843 (N_3843,In_730,In_1635);
and U3844 (N_3844,In_536,In_854);
nand U3845 (N_3845,In_24,In_1324);
or U3846 (N_3846,In_1720,In_386);
xor U3847 (N_3847,In_368,In_41);
or U3848 (N_3848,In_1398,In_216);
xor U3849 (N_3849,In_1803,In_619);
nand U3850 (N_3850,In_347,In_1239);
nor U3851 (N_3851,In_512,In_514);
nand U3852 (N_3852,In_1498,In_1823);
nor U3853 (N_3853,In_1836,In_239);
and U3854 (N_3854,In_1351,In_620);
or U3855 (N_3855,In_1363,In_1270);
nand U3856 (N_3856,In_1408,In_525);
nor U3857 (N_3857,In_61,In_37);
nor U3858 (N_3858,In_434,In_404);
and U3859 (N_3859,In_1464,In_368);
or U3860 (N_3860,In_137,In_1473);
and U3861 (N_3861,In_155,In_1465);
xnor U3862 (N_3862,In_845,In_1928);
nor U3863 (N_3863,In_293,In_1070);
and U3864 (N_3864,In_1923,In_395);
nor U3865 (N_3865,In_1562,In_1402);
or U3866 (N_3866,In_1863,In_708);
nand U3867 (N_3867,In_1720,In_54);
or U3868 (N_3868,In_1693,In_1766);
nand U3869 (N_3869,In_1881,In_1351);
xor U3870 (N_3870,In_1775,In_1413);
xor U3871 (N_3871,In_370,In_238);
nor U3872 (N_3872,In_1791,In_115);
and U3873 (N_3873,In_452,In_488);
and U3874 (N_3874,In_1701,In_1800);
or U3875 (N_3875,In_1735,In_706);
xnor U3876 (N_3876,In_1651,In_709);
or U3877 (N_3877,In_1960,In_973);
and U3878 (N_3878,In_598,In_57);
xor U3879 (N_3879,In_159,In_582);
nand U3880 (N_3880,In_636,In_553);
or U3881 (N_3881,In_158,In_854);
or U3882 (N_3882,In_137,In_1294);
xnor U3883 (N_3883,In_1597,In_1162);
nor U3884 (N_3884,In_1895,In_1230);
or U3885 (N_3885,In_459,In_781);
nor U3886 (N_3886,In_674,In_435);
nand U3887 (N_3887,In_280,In_135);
xor U3888 (N_3888,In_408,In_1973);
xor U3889 (N_3889,In_1816,In_711);
nand U3890 (N_3890,In_1103,In_1765);
xor U3891 (N_3891,In_933,In_691);
and U3892 (N_3892,In_3,In_884);
nand U3893 (N_3893,In_397,In_285);
xor U3894 (N_3894,In_1598,In_1746);
or U3895 (N_3895,In_1366,In_505);
or U3896 (N_3896,In_1,In_2);
or U3897 (N_3897,In_4,In_1384);
and U3898 (N_3898,In_1687,In_321);
nand U3899 (N_3899,In_142,In_476);
nor U3900 (N_3900,In_584,In_1872);
nor U3901 (N_3901,In_1884,In_572);
and U3902 (N_3902,In_427,In_208);
xnor U3903 (N_3903,In_429,In_1758);
nand U3904 (N_3904,In_1224,In_1663);
or U3905 (N_3905,In_1692,In_366);
and U3906 (N_3906,In_1401,In_1636);
or U3907 (N_3907,In_1572,In_1215);
or U3908 (N_3908,In_148,In_1920);
or U3909 (N_3909,In_842,In_220);
or U3910 (N_3910,In_1414,In_1308);
xor U3911 (N_3911,In_683,In_1108);
xor U3912 (N_3912,In_1374,In_1289);
and U3913 (N_3913,In_995,In_1616);
nand U3914 (N_3914,In_1191,In_1608);
xnor U3915 (N_3915,In_406,In_25);
xnor U3916 (N_3916,In_302,In_851);
and U3917 (N_3917,In_926,In_889);
xnor U3918 (N_3918,In_1609,In_71);
xnor U3919 (N_3919,In_1812,In_357);
and U3920 (N_3920,In_1706,In_671);
nor U3921 (N_3921,In_330,In_835);
or U3922 (N_3922,In_1567,In_781);
nand U3923 (N_3923,In_488,In_986);
and U3924 (N_3924,In_1758,In_1360);
nor U3925 (N_3925,In_623,In_1027);
nand U3926 (N_3926,In_814,In_1467);
and U3927 (N_3927,In_1968,In_1184);
and U3928 (N_3928,In_466,In_716);
nand U3929 (N_3929,In_1378,In_321);
or U3930 (N_3930,In_1133,In_730);
nor U3931 (N_3931,In_1924,In_603);
or U3932 (N_3932,In_499,In_886);
nand U3933 (N_3933,In_1513,In_889);
and U3934 (N_3934,In_990,In_33);
nand U3935 (N_3935,In_1167,In_613);
or U3936 (N_3936,In_1294,In_1442);
nand U3937 (N_3937,In_249,In_1686);
xnor U3938 (N_3938,In_831,In_588);
xor U3939 (N_3939,In_457,In_577);
nor U3940 (N_3940,In_763,In_178);
and U3941 (N_3941,In_1778,In_731);
nand U3942 (N_3942,In_480,In_637);
nor U3943 (N_3943,In_471,In_1428);
and U3944 (N_3944,In_579,In_954);
xor U3945 (N_3945,In_638,In_1768);
nor U3946 (N_3946,In_62,In_1354);
xor U3947 (N_3947,In_1374,In_1552);
nand U3948 (N_3948,In_563,In_990);
nor U3949 (N_3949,In_1154,In_1942);
nand U3950 (N_3950,In_515,In_238);
nand U3951 (N_3951,In_1948,In_1021);
nor U3952 (N_3952,In_1714,In_740);
xor U3953 (N_3953,In_1265,In_1468);
and U3954 (N_3954,In_150,In_420);
nor U3955 (N_3955,In_593,In_445);
xor U3956 (N_3956,In_1481,In_1291);
xor U3957 (N_3957,In_169,In_1419);
xnor U3958 (N_3958,In_1264,In_1538);
and U3959 (N_3959,In_425,In_1391);
xor U3960 (N_3960,In_1776,In_215);
or U3961 (N_3961,In_171,In_1663);
or U3962 (N_3962,In_197,In_310);
nand U3963 (N_3963,In_996,In_1904);
nand U3964 (N_3964,In_704,In_1015);
and U3965 (N_3965,In_1400,In_589);
or U3966 (N_3966,In_572,In_1241);
and U3967 (N_3967,In_89,In_157);
nor U3968 (N_3968,In_1160,In_1453);
and U3969 (N_3969,In_1993,In_1073);
and U3970 (N_3970,In_229,In_552);
and U3971 (N_3971,In_1226,In_570);
xnor U3972 (N_3972,In_1023,In_668);
or U3973 (N_3973,In_1662,In_912);
nand U3974 (N_3974,In_1886,In_1371);
and U3975 (N_3975,In_179,In_429);
or U3976 (N_3976,In_982,In_121);
and U3977 (N_3977,In_879,In_1075);
xor U3978 (N_3978,In_178,In_1712);
or U3979 (N_3979,In_30,In_1070);
nand U3980 (N_3980,In_1600,In_1408);
nand U3981 (N_3981,In_1458,In_890);
xnor U3982 (N_3982,In_1750,In_440);
nor U3983 (N_3983,In_793,In_1606);
and U3984 (N_3984,In_457,In_1898);
and U3985 (N_3985,In_402,In_464);
and U3986 (N_3986,In_1131,In_57);
xor U3987 (N_3987,In_798,In_1647);
or U3988 (N_3988,In_995,In_277);
and U3989 (N_3989,In_105,In_3);
or U3990 (N_3990,In_123,In_1575);
or U3991 (N_3991,In_1536,In_1445);
or U3992 (N_3992,In_1816,In_1725);
and U3993 (N_3993,In_1225,In_1902);
and U3994 (N_3994,In_3,In_1054);
nor U3995 (N_3995,In_1758,In_727);
xnor U3996 (N_3996,In_1872,In_1017);
and U3997 (N_3997,In_643,In_1906);
or U3998 (N_3998,In_220,In_1693);
or U3999 (N_3999,In_1272,In_47);
and U4000 (N_4000,In_89,In_1352);
or U4001 (N_4001,In_1424,In_1395);
and U4002 (N_4002,In_1202,In_1091);
nor U4003 (N_4003,In_253,In_1766);
or U4004 (N_4004,In_697,In_521);
xor U4005 (N_4005,In_486,In_1824);
nand U4006 (N_4006,In_596,In_1532);
xor U4007 (N_4007,In_467,In_1505);
nor U4008 (N_4008,In_151,In_1814);
or U4009 (N_4009,In_1606,In_350);
xnor U4010 (N_4010,In_1858,In_1224);
and U4011 (N_4011,In_1131,In_1525);
nand U4012 (N_4012,In_736,In_1998);
xnor U4013 (N_4013,In_1304,In_20);
xnor U4014 (N_4014,In_721,In_447);
and U4015 (N_4015,In_767,In_1318);
nor U4016 (N_4016,In_1673,In_640);
and U4017 (N_4017,In_1967,In_504);
xnor U4018 (N_4018,In_1323,In_1500);
nand U4019 (N_4019,In_102,In_1701);
nor U4020 (N_4020,In_47,In_1194);
nor U4021 (N_4021,In_37,In_1754);
nand U4022 (N_4022,In_1984,In_1694);
and U4023 (N_4023,In_179,In_607);
or U4024 (N_4024,In_5,In_345);
nor U4025 (N_4025,In_1258,In_1404);
and U4026 (N_4026,In_790,In_538);
nand U4027 (N_4027,In_1177,In_656);
xnor U4028 (N_4028,In_309,In_1277);
or U4029 (N_4029,In_1734,In_1264);
xnor U4030 (N_4030,In_1475,In_1434);
and U4031 (N_4031,In_781,In_1178);
nor U4032 (N_4032,In_1387,In_554);
xor U4033 (N_4033,In_1120,In_360);
or U4034 (N_4034,In_1353,In_1568);
and U4035 (N_4035,In_73,In_903);
xnor U4036 (N_4036,In_978,In_585);
xor U4037 (N_4037,In_1353,In_816);
nor U4038 (N_4038,In_66,In_344);
nor U4039 (N_4039,In_1074,In_1050);
xnor U4040 (N_4040,In_255,In_308);
and U4041 (N_4041,In_236,In_512);
xnor U4042 (N_4042,In_1043,In_1011);
and U4043 (N_4043,In_1691,In_1330);
xor U4044 (N_4044,In_283,In_89);
xor U4045 (N_4045,In_1237,In_1411);
nand U4046 (N_4046,In_1855,In_716);
nand U4047 (N_4047,In_746,In_345);
and U4048 (N_4048,In_622,In_1076);
and U4049 (N_4049,In_580,In_227);
nand U4050 (N_4050,In_1920,In_745);
and U4051 (N_4051,In_624,In_279);
xnor U4052 (N_4052,In_1912,In_86);
xor U4053 (N_4053,In_1930,In_1044);
nor U4054 (N_4054,In_445,In_1336);
xnor U4055 (N_4055,In_1512,In_747);
xor U4056 (N_4056,In_829,In_194);
nor U4057 (N_4057,In_647,In_1419);
or U4058 (N_4058,In_1535,In_452);
nor U4059 (N_4059,In_1313,In_803);
nand U4060 (N_4060,In_1017,In_1914);
or U4061 (N_4061,In_1121,In_1470);
nor U4062 (N_4062,In_309,In_1031);
or U4063 (N_4063,In_114,In_343);
nor U4064 (N_4064,In_809,In_758);
xnor U4065 (N_4065,In_1113,In_1031);
nor U4066 (N_4066,In_167,In_367);
nand U4067 (N_4067,In_1935,In_1816);
xnor U4068 (N_4068,In_1216,In_1449);
nand U4069 (N_4069,In_1853,In_1919);
nand U4070 (N_4070,In_216,In_105);
or U4071 (N_4071,In_1822,In_777);
nor U4072 (N_4072,In_292,In_298);
nand U4073 (N_4073,In_1129,In_269);
nor U4074 (N_4074,In_927,In_1208);
nor U4075 (N_4075,In_1154,In_368);
and U4076 (N_4076,In_1873,In_306);
or U4077 (N_4077,In_1801,In_982);
nor U4078 (N_4078,In_516,In_534);
nor U4079 (N_4079,In_145,In_398);
nand U4080 (N_4080,In_1446,In_870);
nand U4081 (N_4081,In_1707,In_1405);
nor U4082 (N_4082,In_648,In_1884);
and U4083 (N_4083,In_1030,In_55);
or U4084 (N_4084,In_1537,In_314);
nor U4085 (N_4085,In_1885,In_300);
nand U4086 (N_4086,In_1543,In_1662);
or U4087 (N_4087,In_1673,In_644);
nor U4088 (N_4088,In_563,In_1721);
nor U4089 (N_4089,In_907,In_289);
nor U4090 (N_4090,In_1041,In_669);
nand U4091 (N_4091,In_1965,In_856);
or U4092 (N_4092,In_1508,In_1743);
nor U4093 (N_4093,In_429,In_1877);
and U4094 (N_4094,In_1230,In_1581);
nor U4095 (N_4095,In_1058,In_721);
nand U4096 (N_4096,In_1228,In_341);
nand U4097 (N_4097,In_1141,In_130);
nor U4098 (N_4098,In_587,In_519);
and U4099 (N_4099,In_1847,In_1704);
or U4100 (N_4100,In_1034,In_648);
or U4101 (N_4101,In_1357,In_1826);
xor U4102 (N_4102,In_1887,In_52);
nand U4103 (N_4103,In_38,In_1303);
or U4104 (N_4104,In_1776,In_1832);
xor U4105 (N_4105,In_165,In_1503);
and U4106 (N_4106,In_101,In_1143);
nor U4107 (N_4107,In_466,In_318);
nor U4108 (N_4108,In_39,In_266);
xor U4109 (N_4109,In_86,In_1493);
nand U4110 (N_4110,In_1408,In_921);
nor U4111 (N_4111,In_1869,In_499);
nor U4112 (N_4112,In_1681,In_689);
nand U4113 (N_4113,In_601,In_909);
xor U4114 (N_4114,In_664,In_1708);
xnor U4115 (N_4115,In_1753,In_303);
xnor U4116 (N_4116,In_521,In_1133);
xor U4117 (N_4117,In_476,In_1711);
or U4118 (N_4118,In_529,In_1938);
nor U4119 (N_4119,In_1866,In_18);
xnor U4120 (N_4120,In_818,In_189);
and U4121 (N_4121,In_1175,In_1870);
or U4122 (N_4122,In_745,In_1493);
nand U4123 (N_4123,In_1015,In_1909);
nor U4124 (N_4124,In_680,In_563);
xnor U4125 (N_4125,In_1319,In_1683);
and U4126 (N_4126,In_1772,In_1714);
nor U4127 (N_4127,In_1223,In_1123);
nand U4128 (N_4128,In_284,In_367);
or U4129 (N_4129,In_912,In_1625);
nor U4130 (N_4130,In_1024,In_372);
nor U4131 (N_4131,In_1215,In_1958);
nand U4132 (N_4132,In_507,In_816);
and U4133 (N_4133,In_1601,In_865);
nor U4134 (N_4134,In_1832,In_444);
or U4135 (N_4135,In_135,In_6);
and U4136 (N_4136,In_839,In_719);
xnor U4137 (N_4137,In_1583,In_176);
xor U4138 (N_4138,In_1416,In_1585);
nor U4139 (N_4139,In_724,In_285);
and U4140 (N_4140,In_1005,In_1718);
or U4141 (N_4141,In_540,In_2);
and U4142 (N_4142,In_212,In_13);
nand U4143 (N_4143,In_179,In_67);
or U4144 (N_4144,In_1603,In_1158);
nor U4145 (N_4145,In_153,In_1563);
xor U4146 (N_4146,In_983,In_1212);
nor U4147 (N_4147,In_375,In_598);
xnor U4148 (N_4148,In_690,In_136);
nand U4149 (N_4149,In_605,In_728);
nand U4150 (N_4150,In_99,In_1842);
or U4151 (N_4151,In_1894,In_1120);
xnor U4152 (N_4152,In_1081,In_1565);
nor U4153 (N_4153,In_659,In_1752);
and U4154 (N_4154,In_769,In_1024);
and U4155 (N_4155,In_1592,In_1992);
nor U4156 (N_4156,In_466,In_172);
and U4157 (N_4157,In_1665,In_1547);
nand U4158 (N_4158,In_1417,In_1012);
nand U4159 (N_4159,In_1773,In_1406);
or U4160 (N_4160,In_6,In_870);
or U4161 (N_4161,In_1921,In_315);
and U4162 (N_4162,In_740,In_814);
and U4163 (N_4163,In_1528,In_1377);
xor U4164 (N_4164,In_366,In_1549);
nor U4165 (N_4165,In_160,In_197);
nor U4166 (N_4166,In_772,In_924);
or U4167 (N_4167,In_1614,In_1684);
and U4168 (N_4168,In_1517,In_1656);
nor U4169 (N_4169,In_1270,In_1247);
xor U4170 (N_4170,In_997,In_225);
xor U4171 (N_4171,In_1128,In_1334);
xnor U4172 (N_4172,In_156,In_501);
or U4173 (N_4173,In_1493,In_947);
nand U4174 (N_4174,In_1917,In_974);
nor U4175 (N_4175,In_1378,In_1533);
xnor U4176 (N_4176,In_744,In_1836);
and U4177 (N_4177,In_709,In_1563);
nor U4178 (N_4178,In_1014,In_1204);
and U4179 (N_4179,In_1073,In_1814);
xor U4180 (N_4180,In_1306,In_349);
xnor U4181 (N_4181,In_1197,In_1971);
nand U4182 (N_4182,In_1701,In_713);
and U4183 (N_4183,In_1058,In_436);
and U4184 (N_4184,In_331,In_1024);
nand U4185 (N_4185,In_1507,In_850);
nor U4186 (N_4186,In_868,In_333);
xor U4187 (N_4187,In_1520,In_1181);
and U4188 (N_4188,In_63,In_1319);
and U4189 (N_4189,In_252,In_666);
or U4190 (N_4190,In_545,In_831);
xor U4191 (N_4191,In_711,In_1961);
and U4192 (N_4192,In_74,In_1240);
or U4193 (N_4193,In_1674,In_1208);
xor U4194 (N_4194,In_1291,In_208);
nor U4195 (N_4195,In_79,In_1419);
xnor U4196 (N_4196,In_1706,In_52);
or U4197 (N_4197,In_1273,In_406);
or U4198 (N_4198,In_427,In_1489);
or U4199 (N_4199,In_1475,In_1284);
nand U4200 (N_4200,In_753,In_51);
or U4201 (N_4201,In_1326,In_249);
or U4202 (N_4202,In_349,In_1989);
xnor U4203 (N_4203,In_1598,In_1594);
and U4204 (N_4204,In_639,In_1584);
nand U4205 (N_4205,In_873,In_514);
xor U4206 (N_4206,In_672,In_635);
xnor U4207 (N_4207,In_1861,In_1259);
nand U4208 (N_4208,In_4,In_1321);
nand U4209 (N_4209,In_1994,In_1147);
xor U4210 (N_4210,In_322,In_353);
nand U4211 (N_4211,In_287,In_998);
nor U4212 (N_4212,In_1026,In_417);
nor U4213 (N_4213,In_915,In_767);
nand U4214 (N_4214,In_1811,In_249);
nor U4215 (N_4215,In_1557,In_996);
and U4216 (N_4216,In_815,In_232);
nor U4217 (N_4217,In_1017,In_510);
xnor U4218 (N_4218,In_1530,In_1332);
nand U4219 (N_4219,In_1864,In_1077);
xor U4220 (N_4220,In_911,In_1322);
and U4221 (N_4221,In_214,In_780);
and U4222 (N_4222,In_226,In_1316);
nor U4223 (N_4223,In_1347,In_1244);
nand U4224 (N_4224,In_1977,In_48);
or U4225 (N_4225,In_906,In_918);
xnor U4226 (N_4226,In_1815,In_1937);
or U4227 (N_4227,In_1705,In_358);
nand U4228 (N_4228,In_666,In_1002);
nor U4229 (N_4229,In_1341,In_1220);
nor U4230 (N_4230,In_964,In_1904);
nor U4231 (N_4231,In_1374,In_307);
nand U4232 (N_4232,In_1966,In_1937);
or U4233 (N_4233,In_1882,In_1701);
nor U4234 (N_4234,In_320,In_1652);
nand U4235 (N_4235,In_986,In_878);
nand U4236 (N_4236,In_746,In_416);
nor U4237 (N_4237,In_1066,In_1679);
nand U4238 (N_4238,In_975,In_684);
nand U4239 (N_4239,In_822,In_834);
or U4240 (N_4240,In_1391,In_17);
or U4241 (N_4241,In_13,In_1630);
nand U4242 (N_4242,In_588,In_684);
nor U4243 (N_4243,In_1060,In_33);
nand U4244 (N_4244,In_1932,In_971);
or U4245 (N_4245,In_1512,In_1161);
and U4246 (N_4246,In_202,In_1530);
and U4247 (N_4247,In_1472,In_290);
xnor U4248 (N_4248,In_181,In_1161);
or U4249 (N_4249,In_1418,In_572);
and U4250 (N_4250,In_184,In_1290);
nand U4251 (N_4251,In_911,In_1101);
or U4252 (N_4252,In_134,In_275);
xnor U4253 (N_4253,In_1405,In_1219);
nor U4254 (N_4254,In_1149,In_688);
and U4255 (N_4255,In_1343,In_1909);
nor U4256 (N_4256,In_1753,In_1135);
and U4257 (N_4257,In_591,In_613);
xor U4258 (N_4258,In_1323,In_1036);
and U4259 (N_4259,In_1025,In_1774);
and U4260 (N_4260,In_396,In_836);
nor U4261 (N_4261,In_272,In_1211);
and U4262 (N_4262,In_855,In_419);
or U4263 (N_4263,In_552,In_1761);
or U4264 (N_4264,In_1884,In_1595);
or U4265 (N_4265,In_688,In_1515);
nand U4266 (N_4266,In_1347,In_300);
or U4267 (N_4267,In_1727,In_801);
nor U4268 (N_4268,In_1664,In_690);
xnor U4269 (N_4269,In_147,In_1401);
and U4270 (N_4270,In_57,In_526);
and U4271 (N_4271,In_1532,In_1585);
xor U4272 (N_4272,In_1137,In_52);
and U4273 (N_4273,In_432,In_1695);
nand U4274 (N_4274,In_417,In_258);
nand U4275 (N_4275,In_173,In_781);
and U4276 (N_4276,In_1938,In_586);
nand U4277 (N_4277,In_1387,In_831);
and U4278 (N_4278,In_1984,In_951);
or U4279 (N_4279,In_624,In_775);
or U4280 (N_4280,In_1340,In_690);
nand U4281 (N_4281,In_406,In_1026);
and U4282 (N_4282,In_1439,In_698);
nor U4283 (N_4283,In_1593,In_983);
nor U4284 (N_4284,In_1908,In_636);
xnor U4285 (N_4285,In_1497,In_1705);
and U4286 (N_4286,In_1604,In_785);
and U4287 (N_4287,In_1335,In_1636);
nand U4288 (N_4288,In_892,In_497);
or U4289 (N_4289,In_882,In_1035);
xor U4290 (N_4290,In_119,In_1323);
xnor U4291 (N_4291,In_800,In_1214);
and U4292 (N_4292,In_1309,In_20);
xnor U4293 (N_4293,In_101,In_568);
and U4294 (N_4294,In_951,In_1761);
nor U4295 (N_4295,In_74,In_897);
or U4296 (N_4296,In_480,In_108);
nor U4297 (N_4297,In_1415,In_1328);
xnor U4298 (N_4298,In_446,In_101);
or U4299 (N_4299,In_1195,In_1595);
and U4300 (N_4300,In_1676,In_1645);
nor U4301 (N_4301,In_1246,In_36);
and U4302 (N_4302,In_936,In_812);
or U4303 (N_4303,In_1031,In_573);
nand U4304 (N_4304,In_50,In_14);
xor U4305 (N_4305,In_422,In_959);
nor U4306 (N_4306,In_1125,In_1847);
nor U4307 (N_4307,In_103,In_1336);
xor U4308 (N_4308,In_904,In_787);
xnor U4309 (N_4309,In_1469,In_605);
nand U4310 (N_4310,In_497,In_1669);
nor U4311 (N_4311,In_991,In_1546);
or U4312 (N_4312,In_38,In_501);
or U4313 (N_4313,In_1573,In_656);
nand U4314 (N_4314,In_818,In_773);
nand U4315 (N_4315,In_1638,In_1500);
xnor U4316 (N_4316,In_1659,In_1432);
nand U4317 (N_4317,In_153,In_1306);
or U4318 (N_4318,In_1079,In_504);
nand U4319 (N_4319,In_1811,In_1798);
nand U4320 (N_4320,In_701,In_890);
xnor U4321 (N_4321,In_424,In_362);
xnor U4322 (N_4322,In_1845,In_253);
nand U4323 (N_4323,In_1927,In_900);
nor U4324 (N_4324,In_631,In_1641);
or U4325 (N_4325,In_1357,In_876);
nor U4326 (N_4326,In_1219,In_1039);
nand U4327 (N_4327,In_43,In_1396);
or U4328 (N_4328,In_965,In_1066);
xnor U4329 (N_4329,In_1104,In_732);
nor U4330 (N_4330,In_194,In_1536);
or U4331 (N_4331,In_631,In_35);
nand U4332 (N_4332,In_1478,In_872);
xnor U4333 (N_4333,In_772,In_697);
or U4334 (N_4334,In_1612,In_1481);
nor U4335 (N_4335,In_1687,In_798);
and U4336 (N_4336,In_1430,In_1450);
or U4337 (N_4337,In_1574,In_1103);
nand U4338 (N_4338,In_1401,In_1894);
or U4339 (N_4339,In_38,In_704);
nor U4340 (N_4340,In_235,In_807);
nor U4341 (N_4341,In_663,In_540);
or U4342 (N_4342,In_1773,In_821);
or U4343 (N_4343,In_606,In_632);
nor U4344 (N_4344,In_1293,In_848);
and U4345 (N_4345,In_1754,In_1355);
or U4346 (N_4346,In_1625,In_994);
or U4347 (N_4347,In_1601,In_1268);
xor U4348 (N_4348,In_812,In_1991);
nand U4349 (N_4349,In_2,In_1996);
nand U4350 (N_4350,In_1873,In_1493);
xor U4351 (N_4351,In_624,In_423);
xnor U4352 (N_4352,In_1595,In_1063);
and U4353 (N_4353,In_1825,In_822);
or U4354 (N_4354,In_502,In_871);
xnor U4355 (N_4355,In_1470,In_302);
and U4356 (N_4356,In_1910,In_1051);
xnor U4357 (N_4357,In_221,In_966);
or U4358 (N_4358,In_632,In_1253);
nand U4359 (N_4359,In_161,In_1246);
nor U4360 (N_4360,In_236,In_297);
and U4361 (N_4361,In_1466,In_797);
nor U4362 (N_4362,In_1990,In_1000);
xor U4363 (N_4363,In_1339,In_1209);
nand U4364 (N_4364,In_1247,In_907);
and U4365 (N_4365,In_1890,In_1244);
or U4366 (N_4366,In_1559,In_107);
and U4367 (N_4367,In_1778,In_1660);
and U4368 (N_4368,In_1664,In_1256);
or U4369 (N_4369,In_1194,In_1152);
nand U4370 (N_4370,In_1086,In_100);
nor U4371 (N_4371,In_1007,In_109);
or U4372 (N_4372,In_381,In_1804);
or U4373 (N_4373,In_160,In_1237);
xnor U4374 (N_4374,In_994,In_1122);
nor U4375 (N_4375,In_966,In_385);
and U4376 (N_4376,In_192,In_477);
xor U4377 (N_4377,In_1044,In_741);
nand U4378 (N_4378,In_374,In_1012);
and U4379 (N_4379,In_1515,In_1863);
nor U4380 (N_4380,In_1998,In_675);
nor U4381 (N_4381,In_1288,In_1509);
and U4382 (N_4382,In_128,In_390);
nor U4383 (N_4383,In_1742,In_1828);
or U4384 (N_4384,In_81,In_1279);
nor U4385 (N_4385,In_382,In_1859);
nand U4386 (N_4386,In_1078,In_649);
or U4387 (N_4387,In_1216,In_814);
or U4388 (N_4388,In_1934,In_742);
nor U4389 (N_4389,In_649,In_588);
and U4390 (N_4390,In_1913,In_1129);
and U4391 (N_4391,In_450,In_1114);
nor U4392 (N_4392,In_818,In_1378);
and U4393 (N_4393,In_1276,In_770);
nor U4394 (N_4394,In_607,In_757);
or U4395 (N_4395,In_1425,In_1074);
or U4396 (N_4396,In_1329,In_1756);
or U4397 (N_4397,In_87,In_747);
xnor U4398 (N_4398,In_1017,In_458);
nand U4399 (N_4399,In_408,In_179);
or U4400 (N_4400,In_1755,In_453);
xnor U4401 (N_4401,In_10,In_1031);
nor U4402 (N_4402,In_1556,In_171);
nand U4403 (N_4403,In_1267,In_1331);
xnor U4404 (N_4404,In_46,In_1567);
nor U4405 (N_4405,In_1429,In_1038);
xor U4406 (N_4406,In_1613,In_96);
or U4407 (N_4407,In_1078,In_1690);
nand U4408 (N_4408,In_1109,In_1517);
and U4409 (N_4409,In_1300,In_43);
nor U4410 (N_4410,In_1179,In_200);
nand U4411 (N_4411,In_653,In_139);
and U4412 (N_4412,In_1676,In_1013);
and U4413 (N_4413,In_1113,In_1277);
nor U4414 (N_4414,In_219,In_1437);
or U4415 (N_4415,In_514,In_547);
xnor U4416 (N_4416,In_1477,In_1221);
or U4417 (N_4417,In_78,In_1367);
or U4418 (N_4418,In_1131,In_1832);
or U4419 (N_4419,In_1408,In_238);
or U4420 (N_4420,In_339,In_1216);
nor U4421 (N_4421,In_1812,In_316);
nor U4422 (N_4422,In_1952,In_428);
and U4423 (N_4423,In_1472,In_871);
and U4424 (N_4424,In_1429,In_39);
xnor U4425 (N_4425,In_1315,In_37);
and U4426 (N_4426,In_813,In_461);
and U4427 (N_4427,In_538,In_220);
xor U4428 (N_4428,In_824,In_451);
nor U4429 (N_4429,In_369,In_1146);
nor U4430 (N_4430,In_204,In_1541);
xnor U4431 (N_4431,In_1218,In_1562);
and U4432 (N_4432,In_1788,In_1773);
nand U4433 (N_4433,In_1508,In_1309);
nor U4434 (N_4434,In_1268,In_1463);
nor U4435 (N_4435,In_664,In_230);
and U4436 (N_4436,In_1942,In_1805);
or U4437 (N_4437,In_773,In_653);
xnor U4438 (N_4438,In_1680,In_1622);
nand U4439 (N_4439,In_347,In_1675);
or U4440 (N_4440,In_466,In_1641);
and U4441 (N_4441,In_156,In_1750);
and U4442 (N_4442,In_34,In_1510);
nand U4443 (N_4443,In_139,In_997);
nand U4444 (N_4444,In_685,In_1596);
or U4445 (N_4445,In_1193,In_1840);
xnor U4446 (N_4446,In_1999,In_1520);
nor U4447 (N_4447,In_208,In_736);
and U4448 (N_4448,In_1296,In_927);
nand U4449 (N_4449,In_902,In_1042);
nand U4450 (N_4450,In_1251,In_1128);
nand U4451 (N_4451,In_1487,In_196);
nor U4452 (N_4452,In_1955,In_558);
nor U4453 (N_4453,In_1884,In_943);
or U4454 (N_4454,In_1870,In_78);
xor U4455 (N_4455,In_1574,In_1711);
nand U4456 (N_4456,In_495,In_319);
nor U4457 (N_4457,In_571,In_1057);
nand U4458 (N_4458,In_1270,In_601);
and U4459 (N_4459,In_1131,In_1201);
and U4460 (N_4460,In_386,In_347);
and U4461 (N_4461,In_1139,In_1529);
and U4462 (N_4462,In_547,In_1422);
xor U4463 (N_4463,In_867,In_584);
and U4464 (N_4464,In_186,In_1024);
or U4465 (N_4465,In_1365,In_250);
xor U4466 (N_4466,In_1531,In_346);
nand U4467 (N_4467,In_574,In_1973);
or U4468 (N_4468,In_1280,In_672);
or U4469 (N_4469,In_496,In_288);
xor U4470 (N_4470,In_1014,In_3);
xor U4471 (N_4471,In_1668,In_1435);
or U4472 (N_4472,In_462,In_51);
xor U4473 (N_4473,In_1741,In_55);
or U4474 (N_4474,In_1240,In_523);
or U4475 (N_4475,In_399,In_917);
and U4476 (N_4476,In_1219,In_1938);
nor U4477 (N_4477,In_1526,In_1301);
or U4478 (N_4478,In_1136,In_36);
or U4479 (N_4479,In_1523,In_1373);
nand U4480 (N_4480,In_1049,In_127);
nor U4481 (N_4481,In_1490,In_480);
or U4482 (N_4482,In_1068,In_185);
xor U4483 (N_4483,In_1671,In_847);
or U4484 (N_4484,In_180,In_1757);
nor U4485 (N_4485,In_589,In_1446);
or U4486 (N_4486,In_787,In_1264);
nand U4487 (N_4487,In_542,In_1444);
nand U4488 (N_4488,In_1231,In_1833);
and U4489 (N_4489,In_582,In_1983);
or U4490 (N_4490,In_1034,In_1380);
or U4491 (N_4491,In_109,In_504);
or U4492 (N_4492,In_1092,In_1378);
nand U4493 (N_4493,In_1336,In_1691);
nand U4494 (N_4494,In_708,In_785);
xnor U4495 (N_4495,In_1241,In_1354);
xor U4496 (N_4496,In_97,In_720);
xor U4497 (N_4497,In_1827,In_1343);
nor U4498 (N_4498,In_733,In_546);
nor U4499 (N_4499,In_266,In_1475);
or U4500 (N_4500,In_652,In_988);
nor U4501 (N_4501,In_281,In_1895);
and U4502 (N_4502,In_1195,In_1399);
or U4503 (N_4503,In_429,In_65);
xnor U4504 (N_4504,In_1392,In_1802);
or U4505 (N_4505,In_926,In_428);
nand U4506 (N_4506,In_911,In_528);
or U4507 (N_4507,In_575,In_645);
and U4508 (N_4508,In_1689,In_206);
xnor U4509 (N_4509,In_1869,In_385);
nand U4510 (N_4510,In_690,In_1218);
nand U4511 (N_4511,In_937,In_1853);
nand U4512 (N_4512,In_792,In_952);
nor U4513 (N_4513,In_976,In_1799);
and U4514 (N_4514,In_449,In_641);
or U4515 (N_4515,In_1445,In_1379);
or U4516 (N_4516,In_1484,In_1681);
nor U4517 (N_4517,In_1946,In_1801);
or U4518 (N_4518,In_1697,In_662);
and U4519 (N_4519,In_1489,In_835);
or U4520 (N_4520,In_432,In_903);
nor U4521 (N_4521,In_369,In_974);
and U4522 (N_4522,In_1388,In_479);
xor U4523 (N_4523,In_488,In_468);
or U4524 (N_4524,In_115,In_1476);
or U4525 (N_4525,In_1794,In_122);
nor U4526 (N_4526,In_239,In_1314);
and U4527 (N_4527,In_1652,In_1071);
nand U4528 (N_4528,In_1693,In_893);
xnor U4529 (N_4529,In_22,In_23);
and U4530 (N_4530,In_624,In_1197);
nand U4531 (N_4531,In_152,In_227);
nand U4532 (N_4532,In_358,In_1521);
or U4533 (N_4533,In_650,In_794);
xnor U4534 (N_4534,In_1158,In_1874);
nand U4535 (N_4535,In_832,In_111);
or U4536 (N_4536,In_1905,In_1997);
or U4537 (N_4537,In_613,In_952);
nand U4538 (N_4538,In_1541,In_1992);
and U4539 (N_4539,In_161,In_1432);
or U4540 (N_4540,In_871,In_225);
and U4541 (N_4541,In_877,In_719);
and U4542 (N_4542,In_1765,In_565);
nor U4543 (N_4543,In_356,In_83);
and U4544 (N_4544,In_1718,In_1770);
xor U4545 (N_4545,In_1901,In_1051);
and U4546 (N_4546,In_679,In_1174);
nand U4547 (N_4547,In_1589,In_126);
or U4548 (N_4548,In_1219,In_1201);
nor U4549 (N_4549,In_829,In_878);
xor U4550 (N_4550,In_1112,In_1306);
or U4551 (N_4551,In_1161,In_176);
nor U4552 (N_4552,In_1421,In_1476);
nor U4553 (N_4553,In_1863,In_287);
or U4554 (N_4554,In_143,In_1365);
xnor U4555 (N_4555,In_1666,In_536);
nand U4556 (N_4556,In_1321,In_693);
nand U4557 (N_4557,In_560,In_779);
and U4558 (N_4558,In_674,In_1757);
xnor U4559 (N_4559,In_1490,In_61);
or U4560 (N_4560,In_245,In_1009);
nand U4561 (N_4561,In_1207,In_558);
or U4562 (N_4562,In_226,In_26);
nand U4563 (N_4563,In_1483,In_430);
or U4564 (N_4564,In_159,In_130);
xnor U4565 (N_4565,In_1570,In_357);
nand U4566 (N_4566,In_1417,In_230);
nand U4567 (N_4567,In_98,In_680);
nor U4568 (N_4568,In_1910,In_1975);
xor U4569 (N_4569,In_1095,In_276);
nor U4570 (N_4570,In_1303,In_65);
or U4571 (N_4571,In_131,In_793);
nor U4572 (N_4572,In_1067,In_208);
and U4573 (N_4573,In_1246,In_433);
nand U4574 (N_4574,In_1382,In_468);
and U4575 (N_4575,In_994,In_76);
or U4576 (N_4576,In_1346,In_1465);
nor U4577 (N_4577,In_881,In_1125);
or U4578 (N_4578,In_1788,In_1868);
xor U4579 (N_4579,In_376,In_1234);
or U4580 (N_4580,In_602,In_1824);
or U4581 (N_4581,In_842,In_1879);
xnor U4582 (N_4582,In_1707,In_1783);
nand U4583 (N_4583,In_1381,In_1225);
nor U4584 (N_4584,In_857,In_1609);
and U4585 (N_4585,In_802,In_237);
nor U4586 (N_4586,In_821,In_1013);
or U4587 (N_4587,In_94,In_563);
nor U4588 (N_4588,In_325,In_251);
xor U4589 (N_4589,In_1004,In_559);
nand U4590 (N_4590,In_216,In_1159);
and U4591 (N_4591,In_1776,In_650);
and U4592 (N_4592,In_1658,In_710);
nand U4593 (N_4593,In_1089,In_557);
nand U4594 (N_4594,In_302,In_889);
xnor U4595 (N_4595,In_1884,In_1521);
nor U4596 (N_4596,In_782,In_1273);
or U4597 (N_4597,In_213,In_1486);
and U4598 (N_4598,In_1072,In_323);
or U4599 (N_4599,In_15,In_941);
nor U4600 (N_4600,In_1930,In_1490);
and U4601 (N_4601,In_1173,In_681);
nand U4602 (N_4602,In_150,In_438);
or U4603 (N_4603,In_1945,In_116);
nor U4604 (N_4604,In_1376,In_760);
or U4605 (N_4605,In_713,In_1465);
nand U4606 (N_4606,In_1855,In_307);
and U4607 (N_4607,In_1954,In_1090);
xnor U4608 (N_4608,In_600,In_91);
or U4609 (N_4609,In_141,In_1734);
and U4610 (N_4610,In_826,In_1389);
nor U4611 (N_4611,In_1817,In_1822);
nor U4612 (N_4612,In_1384,In_272);
nand U4613 (N_4613,In_1121,In_43);
nand U4614 (N_4614,In_314,In_1381);
or U4615 (N_4615,In_1701,In_684);
xnor U4616 (N_4616,In_576,In_1011);
xnor U4617 (N_4617,In_1891,In_894);
nor U4618 (N_4618,In_1271,In_265);
nand U4619 (N_4619,In_924,In_1430);
and U4620 (N_4620,In_1980,In_1694);
and U4621 (N_4621,In_754,In_804);
xor U4622 (N_4622,In_399,In_818);
and U4623 (N_4623,In_1331,In_1288);
nor U4624 (N_4624,In_1129,In_1153);
or U4625 (N_4625,In_276,In_901);
and U4626 (N_4626,In_1008,In_1633);
and U4627 (N_4627,In_454,In_721);
or U4628 (N_4628,In_895,In_606);
nand U4629 (N_4629,In_1916,In_1636);
or U4630 (N_4630,In_995,In_675);
or U4631 (N_4631,In_1441,In_813);
nor U4632 (N_4632,In_756,In_298);
xnor U4633 (N_4633,In_1150,In_334);
xnor U4634 (N_4634,In_1427,In_393);
and U4635 (N_4635,In_695,In_1075);
xnor U4636 (N_4636,In_1523,In_682);
nor U4637 (N_4637,In_756,In_146);
and U4638 (N_4638,In_1481,In_1690);
nand U4639 (N_4639,In_40,In_486);
and U4640 (N_4640,In_840,In_440);
nor U4641 (N_4641,In_604,In_620);
nor U4642 (N_4642,In_729,In_899);
or U4643 (N_4643,In_51,In_311);
nor U4644 (N_4644,In_221,In_1244);
nand U4645 (N_4645,In_1019,In_534);
or U4646 (N_4646,In_1683,In_901);
and U4647 (N_4647,In_74,In_317);
or U4648 (N_4648,In_1930,In_1120);
nor U4649 (N_4649,In_40,In_1130);
nor U4650 (N_4650,In_1883,In_1096);
nor U4651 (N_4651,In_1286,In_52);
or U4652 (N_4652,In_922,In_206);
xnor U4653 (N_4653,In_575,In_1167);
nor U4654 (N_4654,In_1379,In_1138);
and U4655 (N_4655,In_1143,In_1837);
nor U4656 (N_4656,In_782,In_1920);
xor U4657 (N_4657,In_1351,In_1834);
xnor U4658 (N_4658,In_1887,In_698);
xor U4659 (N_4659,In_452,In_856);
xor U4660 (N_4660,In_1876,In_29);
and U4661 (N_4661,In_1655,In_1918);
or U4662 (N_4662,In_1001,In_1867);
nor U4663 (N_4663,In_854,In_1752);
and U4664 (N_4664,In_1796,In_117);
nor U4665 (N_4665,In_12,In_879);
nor U4666 (N_4666,In_1812,In_1008);
or U4667 (N_4667,In_231,In_1600);
nand U4668 (N_4668,In_532,In_1025);
and U4669 (N_4669,In_717,In_352);
or U4670 (N_4670,In_824,In_1278);
nor U4671 (N_4671,In_202,In_1895);
xnor U4672 (N_4672,In_1447,In_822);
and U4673 (N_4673,In_1288,In_174);
xnor U4674 (N_4674,In_1750,In_378);
nand U4675 (N_4675,In_1989,In_79);
or U4676 (N_4676,In_1238,In_741);
xnor U4677 (N_4677,In_1929,In_1980);
and U4678 (N_4678,In_175,In_1377);
nand U4679 (N_4679,In_910,In_1225);
xnor U4680 (N_4680,In_1805,In_1357);
or U4681 (N_4681,In_1526,In_1355);
or U4682 (N_4682,In_1290,In_615);
xor U4683 (N_4683,In_1066,In_1493);
nand U4684 (N_4684,In_1274,In_1996);
nand U4685 (N_4685,In_1886,In_1761);
nand U4686 (N_4686,In_736,In_1078);
nand U4687 (N_4687,In_1143,In_1696);
nor U4688 (N_4688,In_1334,In_1747);
or U4689 (N_4689,In_1984,In_1987);
nand U4690 (N_4690,In_1808,In_1832);
nand U4691 (N_4691,In_618,In_450);
xor U4692 (N_4692,In_55,In_1367);
and U4693 (N_4693,In_226,In_1142);
and U4694 (N_4694,In_431,In_1137);
xnor U4695 (N_4695,In_1060,In_1583);
xnor U4696 (N_4696,In_1319,In_611);
or U4697 (N_4697,In_511,In_1109);
nor U4698 (N_4698,In_798,In_1230);
xnor U4699 (N_4699,In_1035,In_129);
xnor U4700 (N_4700,In_1952,In_575);
nand U4701 (N_4701,In_712,In_1952);
nand U4702 (N_4702,In_1196,In_1527);
xor U4703 (N_4703,In_896,In_1954);
xnor U4704 (N_4704,In_568,In_949);
or U4705 (N_4705,In_123,In_702);
or U4706 (N_4706,In_1554,In_317);
nand U4707 (N_4707,In_1262,In_1869);
nand U4708 (N_4708,In_292,In_1620);
or U4709 (N_4709,In_1183,In_1848);
or U4710 (N_4710,In_1439,In_1786);
or U4711 (N_4711,In_1079,In_498);
nand U4712 (N_4712,In_1561,In_64);
nor U4713 (N_4713,In_697,In_1747);
nor U4714 (N_4714,In_1271,In_660);
xor U4715 (N_4715,In_1510,In_938);
or U4716 (N_4716,In_1272,In_362);
and U4717 (N_4717,In_997,In_975);
and U4718 (N_4718,In_722,In_1008);
nand U4719 (N_4719,In_270,In_1846);
or U4720 (N_4720,In_135,In_568);
nand U4721 (N_4721,In_1079,In_291);
or U4722 (N_4722,In_228,In_34);
xnor U4723 (N_4723,In_27,In_1488);
or U4724 (N_4724,In_204,In_1892);
xor U4725 (N_4725,In_219,In_997);
or U4726 (N_4726,In_1607,In_1032);
or U4727 (N_4727,In_1404,In_1951);
xor U4728 (N_4728,In_1470,In_1491);
xnor U4729 (N_4729,In_1809,In_803);
nor U4730 (N_4730,In_898,In_647);
nand U4731 (N_4731,In_1631,In_1909);
nand U4732 (N_4732,In_1328,In_1329);
and U4733 (N_4733,In_1824,In_363);
nor U4734 (N_4734,In_972,In_1262);
and U4735 (N_4735,In_988,In_1890);
nor U4736 (N_4736,In_1287,In_197);
or U4737 (N_4737,In_1747,In_876);
and U4738 (N_4738,In_275,In_270);
or U4739 (N_4739,In_62,In_1909);
or U4740 (N_4740,In_1547,In_1424);
and U4741 (N_4741,In_93,In_936);
xnor U4742 (N_4742,In_1819,In_1292);
nor U4743 (N_4743,In_242,In_143);
or U4744 (N_4744,In_673,In_77);
nor U4745 (N_4745,In_92,In_1371);
nor U4746 (N_4746,In_287,In_211);
nor U4747 (N_4747,In_1049,In_656);
or U4748 (N_4748,In_666,In_1884);
xor U4749 (N_4749,In_1040,In_1538);
and U4750 (N_4750,In_1120,In_1910);
nor U4751 (N_4751,In_756,In_1134);
nand U4752 (N_4752,In_668,In_1154);
nor U4753 (N_4753,In_1084,In_1897);
nor U4754 (N_4754,In_1799,In_935);
nand U4755 (N_4755,In_957,In_977);
xor U4756 (N_4756,In_125,In_1392);
nor U4757 (N_4757,In_984,In_1485);
xor U4758 (N_4758,In_1872,In_1364);
nand U4759 (N_4759,In_1484,In_41);
xnor U4760 (N_4760,In_1670,In_1657);
and U4761 (N_4761,In_1942,In_458);
nand U4762 (N_4762,In_415,In_1967);
or U4763 (N_4763,In_774,In_659);
and U4764 (N_4764,In_221,In_1806);
nor U4765 (N_4765,In_1089,In_712);
nor U4766 (N_4766,In_1800,In_388);
or U4767 (N_4767,In_621,In_318);
or U4768 (N_4768,In_1634,In_1942);
or U4769 (N_4769,In_943,In_58);
and U4770 (N_4770,In_195,In_1933);
nor U4771 (N_4771,In_1555,In_748);
xnor U4772 (N_4772,In_1303,In_297);
or U4773 (N_4773,In_1988,In_96);
and U4774 (N_4774,In_1702,In_1321);
xor U4775 (N_4775,In_1623,In_1359);
nand U4776 (N_4776,In_1123,In_1579);
and U4777 (N_4777,In_500,In_1438);
nand U4778 (N_4778,In_518,In_1609);
or U4779 (N_4779,In_374,In_394);
nor U4780 (N_4780,In_1881,In_761);
or U4781 (N_4781,In_471,In_283);
or U4782 (N_4782,In_944,In_991);
xnor U4783 (N_4783,In_487,In_608);
or U4784 (N_4784,In_602,In_664);
xnor U4785 (N_4785,In_45,In_486);
xnor U4786 (N_4786,In_497,In_1191);
nand U4787 (N_4787,In_1362,In_1216);
nand U4788 (N_4788,In_265,In_288);
xnor U4789 (N_4789,In_909,In_361);
nand U4790 (N_4790,In_1010,In_24);
xnor U4791 (N_4791,In_1874,In_164);
and U4792 (N_4792,In_661,In_754);
nor U4793 (N_4793,In_1069,In_88);
or U4794 (N_4794,In_1018,In_1821);
or U4795 (N_4795,In_718,In_1858);
xnor U4796 (N_4796,In_1399,In_1687);
and U4797 (N_4797,In_1034,In_1328);
and U4798 (N_4798,In_230,In_470);
nor U4799 (N_4799,In_444,In_1074);
nor U4800 (N_4800,In_592,In_570);
nor U4801 (N_4801,In_1913,In_393);
nor U4802 (N_4802,In_77,In_427);
and U4803 (N_4803,In_859,In_1242);
and U4804 (N_4804,In_630,In_290);
or U4805 (N_4805,In_1772,In_211);
nor U4806 (N_4806,In_1479,In_1358);
nor U4807 (N_4807,In_635,In_1874);
nor U4808 (N_4808,In_727,In_577);
xnor U4809 (N_4809,In_1997,In_723);
xnor U4810 (N_4810,In_258,In_970);
or U4811 (N_4811,In_1902,In_1361);
or U4812 (N_4812,In_1661,In_1276);
nand U4813 (N_4813,In_1914,In_1978);
nor U4814 (N_4814,In_1104,In_1427);
and U4815 (N_4815,In_1628,In_1006);
nand U4816 (N_4816,In_1348,In_564);
nor U4817 (N_4817,In_244,In_893);
or U4818 (N_4818,In_1748,In_725);
nand U4819 (N_4819,In_1365,In_1493);
nand U4820 (N_4820,In_1334,In_1589);
xnor U4821 (N_4821,In_38,In_875);
and U4822 (N_4822,In_1945,In_1397);
nor U4823 (N_4823,In_260,In_660);
or U4824 (N_4824,In_98,In_1302);
nand U4825 (N_4825,In_182,In_1467);
xnor U4826 (N_4826,In_1678,In_777);
nor U4827 (N_4827,In_572,In_868);
nor U4828 (N_4828,In_967,In_376);
nor U4829 (N_4829,In_903,In_310);
or U4830 (N_4830,In_745,In_928);
nand U4831 (N_4831,In_304,In_1499);
nor U4832 (N_4832,In_1309,In_1480);
and U4833 (N_4833,In_1737,In_805);
and U4834 (N_4834,In_1606,In_841);
nand U4835 (N_4835,In_1373,In_571);
nand U4836 (N_4836,In_893,In_1900);
nand U4837 (N_4837,In_1743,In_1718);
nand U4838 (N_4838,In_685,In_1041);
nor U4839 (N_4839,In_1480,In_226);
and U4840 (N_4840,In_558,In_1579);
xor U4841 (N_4841,In_5,In_1160);
xor U4842 (N_4842,In_290,In_1724);
nand U4843 (N_4843,In_1415,In_14);
and U4844 (N_4844,In_970,In_554);
nand U4845 (N_4845,In_1020,In_692);
xor U4846 (N_4846,In_1797,In_1163);
or U4847 (N_4847,In_1142,In_57);
nor U4848 (N_4848,In_533,In_596);
and U4849 (N_4849,In_1743,In_1998);
xnor U4850 (N_4850,In_1343,In_20);
xnor U4851 (N_4851,In_1317,In_1162);
nand U4852 (N_4852,In_1483,In_1493);
nor U4853 (N_4853,In_1098,In_497);
nor U4854 (N_4854,In_1928,In_1256);
nor U4855 (N_4855,In_411,In_355);
and U4856 (N_4856,In_501,In_843);
nor U4857 (N_4857,In_1642,In_1629);
or U4858 (N_4858,In_265,In_763);
or U4859 (N_4859,In_1586,In_1952);
and U4860 (N_4860,In_92,In_1760);
or U4861 (N_4861,In_56,In_1836);
nor U4862 (N_4862,In_202,In_968);
or U4863 (N_4863,In_884,In_19);
nor U4864 (N_4864,In_1264,In_1270);
and U4865 (N_4865,In_666,In_977);
and U4866 (N_4866,In_375,In_1069);
xnor U4867 (N_4867,In_463,In_392);
or U4868 (N_4868,In_627,In_1529);
xor U4869 (N_4869,In_207,In_1838);
and U4870 (N_4870,In_58,In_1847);
or U4871 (N_4871,In_910,In_1607);
or U4872 (N_4872,In_1080,In_67);
and U4873 (N_4873,In_837,In_1425);
and U4874 (N_4874,In_902,In_467);
or U4875 (N_4875,In_1539,In_450);
and U4876 (N_4876,In_267,In_1699);
nand U4877 (N_4877,In_1756,In_1897);
and U4878 (N_4878,In_1806,In_1799);
and U4879 (N_4879,In_1072,In_879);
or U4880 (N_4880,In_778,In_30);
xnor U4881 (N_4881,In_998,In_1831);
nor U4882 (N_4882,In_1853,In_1222);
xnor U4883 (N_4883,In_1632,In_331);
xor U4884 (N_4884,In_1928,In_1855);
nand U4885 (N_4885,In_1555,In_680);
nand U4886 (N_4886,In_1421,In_1945);
nor U4887 (N_4887,In_125,In_469);
nand U4888 (N_4888,In_1877,In_1521);
nand U4889 (N_4889,In_1718,In_1285);
or U4890 (N_4890,In_1295,In_1020);
nor U4891 (N_4891,In_551,In_1337);
and U4892 (N_4892,In_1508,In_791);
or U4893 (N_4893,In_788,In_1048);
nand U4894 (N_4894,In_1962,In_412);
or U4895 (N_4895,In_1953,In_306);
xnor U4896 (N_4896,In_815,In_175);
nand U4897 (N_4897,In_223,In_1940);
and U4898 (N_4898,In_273,In_575);
or U4899 (N_4899,In_1680,In_1056);
nand U4900 (N_4900,In_73,In_1398);
nor U4901 (N_4901,In_276,In_1040);
and U4902 (N_4902,In_1280,In_1879);
nand U4903 (N_4903,In_100,In_1237);
nor U4904 (N_4904,In_1045,In_1576);
nand U4905 (N_4905,In_1822,In_78);
or U4906 (N_4906,In_1668,In_1009);
nor U4907 (N_4907,In_1160,In_1102);
nand U4908 (N_4908,In_832,In_296);
nor U4909 (N_4909,In_409,In_1200);
xor U4910 (N_4910,In_1121,In_1231);
or U4911 (N_4911,In_240,In_1449);
and U4912 (N_4912,In_1264,In_413);
or U4913 (N_4913,In_79,In_1703);
nor U4914 (N_4914,In_1136,In_1259);
or U4915 (N_4915,In_1437,In_1781);
nor U4916 (N_4916,In_1538,In_677);
or U4917 (N_4917,In_123,In_292);
xnor U4918 (N_4918,In_1655,In_356);
nand U4919 (N_4919,In_9,In_1911);
xnor U4920 (N_4920,In_567,In_897);
xor U4921 (N_4921,In_607,In_1457);
nand U4922 (N_4922,In_901,In_1527);
or U4923 (N_4923,In_181,In_96);
nand U4924 (N_4924,In_1967,In_441);
xor U4925 (N_4925,In_1086,In_1749);
nor U4926 (N_4926,In_1798,In_240);
nor U4927 (N_4927,In_1417,In_964);
xnor U4928 (N_4928,In_765,In_158);
nor U4929 (N_4929,In_1567,In_951);
nand U4930 (N_4930,In_660,In_795);
xnor U4931 (N_4931,In_742,In_466);
or U4932 (N_4932,In_944,In_549);
and U4933 (N_4933,In_1281,In_506);
nand U4934 (N_4934,In_26,In_1622);
nand U4935 (N_4935,In_1392,In_1298);
nor U4936 (N_4936,In_386,In_1132);
xnor U4937 (N_4937,In_1416,In_1865);
or U4938 (N_4938,In_31,In_1932);
nand U4939 (N_4939,In_1926,In_1725);
and U4940 (N_4940,In_254,In_704);
or U4941 (N_4941,In_592,In_457);
nand U4942 (N_4942,In_295,In_864);
nor U4943 (N_4943,In_954,In_747);
nor U4944 (N_4944,In_338,In_1756);
nor U4945 (N_4945,In_846,In_1857);
xnor U4946 (N_4946,In_1320,In_1993);
or U4947 (N_4947,In_899,In_511);
nor U4948 (N_4948,In_490,In_604);
and U4949 (N_4949,In_698,In_1074);
and U4950 (N_4950,In_1117,In_1421);
nor U4951 (N_4951,In_1390,In_1152);
or U4952 (N_4952,In_99,In_775);
nand U4953 (N_4953,In_233,In_1761);
nand U4954 (N_4954,In_1465,In_706);
or U4955 (N_4955,In_513,In_285);
nand U4956 (N_4956,In_683,In_1476);
nand U4957 (N_4957,In_1587,In_34);
nand U4958 (N_4958,In_1098,In_640);
nand U4959 (N_4959,In_1462,In_1049);
and U4960 (N_4960,In_170,In_227);
nand U4961 (N_4961,In_1373,In_1489);
and U4962 (N_4962,In_393,In_1133);
or U4963 (N_4963,In_1849,In_96);
xor U4964 (N_4964,In_811,In_1466);
nor U4965 (N_4965,In_884,In_1686);
nand U4966 (N_4966,In_1644,In_777);
xnor U4967 (N_4967,In_239,In_897);
and U4968 (N_4968,In_1527,In_1267);
nand U4969 (N_4969,In_413,In_972);
or U4970 (N_4970,In_476,In_542);
nand U4971 (N_4971,In_1811,In_1297);
xnor U4972 (N_4972,In_1063,In_1105);
or U4973 (N_4973,In_846,In_203);
nor U4974 (N_4974,In_1104,In_1629);
nor U4975 (N_4975,In_426,In_1256);
nand U4976 (N_4976,In_857,In_53);
xor U4977 (N_4977,In_1943,In_1628);
and U4978 (N_4978,In_39,In_386);
or U4979 (N_4979,In_1871,In_906);
and U4980 (N_4980,In_992,In_20);
and U4981 (N_4981,In_1882,In_667);
xor U4982 (N_4982,In_515,In_812);
nand U4983 (N_4983,In_291,In_665);
nor U4984 (N_4984,In_126,In_1843);
and U4985 (N_4985,In_1010,In_1953);
or U4986 (N_4986,In_177,In_1621);
or U4987 (N_4987,In_1755,In_52);
or U4988 (N_4988,In_1929,In_628);
and U4989 (N_4989,In_1986,In_336);
and U4990 (N_4990,In_199,In_1140);
and U4991 (N_4991,In_951,In_964);
nor U4992 (N_4992,In_1154,In_864);
nand U4993 (N_4993,In_359,In_1132);
xnor U4994 (N_4994,In_347,In_1720);
xor U4995 (N_4995,In_772,In_20);
and U4996 (N_4996,In_1312,In_919);
or U4997 (N_4997,In_1000,In_1896);
and U4998 (N_4998,In_1331,In_276);
nand U4999 (N_4999,In_1614,In_1064);
xor U5000 (N_5000,N_44,N_2909);
xor U5001 (N_5001,N_2699,N_1615);
nand U5002 (N_5002,N_4863,N_1691);
nor U5003 (N_5003,N_1,N_1189);
nand U5004 (N_5004,N_2392,N_2937);
nor U5005 (N_5005,N_146,N_2565);
xor U5006 (N_5006,N_2185,N_1588);
nand U5007 (N_5007,N_3344,N_1136);
or U5008 (N_5008,N_3210,N_1815);
and U5009 (N_5009,N_3161,N_4677);
and U5010 (N_5010,N_2441,N_3758);
and U5011 (N_5011,N_2611,N_1260);
nand U5012 (N_5012,N_2356,N_699);
and U5013 (N_5013,N_4419,N_4026);
xnor U5014 (N_5014,N_1750,N_2207);
xnor U5015 (N_5015,N_2638,N_2732);
nand U5016 (N_5016,N_887,N_1419);
nor U5017 (N_5017,N_539,N_3932);
xor U5018 (N_5018,N_90,N_3386);
nand U5019 (N_5019,N_2537,N_617);
nor U5020 (N_5020,N_4631,N_4766);
xnor U5021 (N_5021,N_930,N_1655);
or U5022 (N_5022,N_3508,N_1491);
nand U5023 (N_5023,N_4099,N_911);
xor U5024 (N_5024,N_2456,N_2758);
xnor U5025 (N_5025,N_2958,N_2544);
xor U5026 (N_5026,N_673,N_1767);
and U5027 (N_5027,N_2385,N_3786);
nand U5028 (N_5028,N_3804,N_4415);
or U5029 (N_5029,N_3167,N_23);
nor U5030 (N_5030,N_4877,N_949);
or U5031 (N_5031,N_2703,N_3733);
nand U5032 (N_5032,N_4842,N_1503);
or U5033 (N_5033,N_1965,N_4034);
xnor U5034 (N_5034,N_1004,N_2679);
nor U5035 (N_5035,N_2196,N_4079);
or U5036 (N_5036,N_4919,N_450);
and U5037 (N_5037,N_2495,N_1169);
nand U5038 (N_5038,N_4222,N_3059);
nand U5039 (N_5039,N_3005,N_414);
xor U5040 (N_5040,N_2457,N_2307);
or U5041 (N_5041,N_3654,N_1879);
nand U5042 (N_5042,N_2038,N_106);
or U5043 (N_5043,N_4769,N_4319);
nand U5044 (N_5044,N_1974,N_3954);
or U5045 (N_5045,N_1353,N_2523);
nand U5046 (N_5046,N_2923,N_3855);
xnor U5047 (N_5047,N_536,N_1309);
nor U5048 (N_5048,N_3384,N_884);
nor U5049 (N_5049,N_260,N_3044);
nor U5050 (N_5050,N_4829,N_2686);
nand U5051 (N_5051,N_1976,N_920);
nand U5052 (N_5052,N_3459,N_2625);
nor U5053 (N_5053,N_2733,N_1720);
nand U5054 (N_5054,N_712,N_3807);
or U5055 (N_5055,N_2498,N_2464);
nand U5056 (N_5056,N_2828,N_2993);
nand U5057 (N_5057,N_4851,N_1159);
nor U5058 (N_5058,N_2979,N_4111);
nor U5059 (N_5059,N_4186,N_679);
nand U5060 (N_5060,N_3628,N_3477);
xnor U5061 (N_5061,N_126,N_1301);
or U5062 (N_5062,N_1031,N_772);
or U5063 (N_5063,N_1852,N_3076);
and U5064 (N_5064,N_3526,N_4812);
xnor U5065 (N_5065,N_2566,N_1039);
nand U5066 (N_5066,N_2424,N_2559);
and U5067 (N_5067,N_2587,N_1064);
xor U5068 (N_5068,N_705,N_4762);
or U5069 (N_5069,N_1683,N_4834);
and U5070 (N_5070,N_893,N_2721);
or U5071 (N_5071,N_4441,N_1649);
and U5072 (N_5072,N_4515,N_1404);
or U5073 (N_5073,N_1798,N_2235);
xor U5074 (N_5074,N_1687,N_812);
xor U5075 (N_5075,N_1198,N_833);
xor U5076 (N_5076,N_1607,N_4809);
or U5077 (N_5077,N_4593,N_2402);
and U5078 (N_5078,N_4131,N_3458);
and U5079 (N_5079,N_141,N_1343);
nor U5080 (N_5080,N_4152,N_1475);
or U5081 (N_5081,N_1785,N_3613);
xor U5082 (N_5082,N_1188,N_4890);
xnor U5083 (N_5083,N_490,N_4835);
xnor U5084 (N_5084,N_3764,N_4101);
and U5085 (N_5085,N_4523,N_296);
nand U5086 (N_5086,N_4015,N_4090);
or U5087 (N_5087,N_3684,N_2555);
nand U5088 (N_5088,N_4698,N_2560);
nor U5089 (N_5089,N_1375,N_26);
or U5090 (N_5090,N_3399,N_825);
nor U5091 (N_5091,N_7,N_1949);
or U5092 (N_5092,N_3826,N_4761);
nand U5093 (N_5093,N_2126,N_4917);
nand U5094 (N_5094,N_4732,N_2972);
or U5095 (N_5095,N_602,N_159);
or U5096 (N_5096,N_694,N_1313);
nor U5097 (N_5097,N_4146,N_666);
and U5098 (N_5098,N_4003,N_1902);
xnor U5099 (N_5099,N_3061,N_1308);
and U5100 (N_5100,N_2195,N_3986);
and U5101 (N_5101,N_4781,N_1211);
or U5102 (N_5102,N_3974,N_3506);
xnor U5103 (N_5103,N_1812,N_3294);
and U5104 (N_5104,N_3325,N_1730);
nand U5105 (N_5105,N_1816,N_950);
nor U5106 (N_5106,N_678,N_243);
or U5107 (N_5107,N_3748,N_4516);
or U5108 (N_5108,N_3484,N_4109);
and U5109 (N_5109,N_3619,N_83);
nand U5110 (N_5110,N_2744,N_4774);
and U5111 (N_5111,N_4342,N_4243);
nand U5112 (N_5112,N_81,N_1387);
xor U5113 (N_5113,N_4276,N_780);
and U5114 (N_5114,N_1851,N_1326);
or U5115 (N_5115,N_760,N_10);
nor U5116 (N_5116,N_3078,N_4576);
or U5117 (N_5117,N_4310,N_1899);
or U5118 (N_5118,N_276,N_316);
or U5119 (N_5119,N_227,N_1924);
nor U5120 (N_5120,N_4849,N_2573);
or U5121 (N_5121,N_2206,N_2757);
and U5122 (N_5122,N_4929,N_2709);
nand U5123 (N_5123,N_733,N_171);
nand U5124 (N_5124,N_3162,N_4689);
and U5125 (N_5125,N_2528,N_1487);
and U5126 (N_5126,N_1534,N_2026);
or U5127 (N_5127,N_909,N_4081);
and U5128 (N_5128,N_2877,N_2610);
xnor U5129 (N_5129,N_2605,N_3412);
and U5130 (N_5130,N_2364,N_706);
or U5131 (N_5131,N_2443,N_1719);
or U5132 (N_5132,N_2811,N_3434);
nand U5133 (N_5133,N_2924,N_293);
or U5134 (N_5134,N_357,N_4258);
or U5135 (N_5135,N_4174,N_1954);
nand U5136 (N_5136,N_2349,N_3001);
and U5137 (N_5137,N_116,N_4251);
xor U5138 (N_5138,N_716,N_3272);
and U5139 (N_5139,N_4316,N_3569);
or U5140 (N_5140,N_4436,N_324);
nor U5141 (N_5141,N_1286,N_3347);
and U5142 (N_5142,N_1060,N_3949);
xor U5143 (N_5143,N_703,N_3847);
and U5144 (N_5144,N_2850,N_790);
xor U5145 (N_5145,N_1782,N_3732);
nor U5146 (N_5146,N_1645,N_3035);
and U5147 (N_5147,N_2664,N_1075);
nor U5148 (N_5148,N_1323,N_2191);
or U5149 (N_5149,N_1870,N_522);
nand U5150 (N_5150,N_1805,N_933);
or U5151 (N_5151,N_5,N_1803);
nand U5152 (N_5152,N_3086,N_2120);
and U5153 (N_5153,N_4971,N_4730);
and U5154 (N_5154,N_4140,N_3580);
and U5155 (N_5155,N_1081,N_3181);
nand U5156 (N_5156,N_4786,N_3878);
and U5157 (N_5157,N_3025,N_624);
xor U5158 (N_5158,N_601,N_4855);
and U5159 (N_5159,N_4748,N_1756);
or U5160 (N_5160,N_4616,N_1408);
and U5161 (N_5161,N_3124,N_1495);
and U5162 (N_5162,N_4254,N_2722);
or U5163 (N_5163,N_2561,N_4473);
xnor U5164 (N_5164,N_2070,N_1436);
nand U5165 (N_5165,N_1276,N_4826);
xor U5166 (N_5166,N_2752,N_2230);
or U5167 (N_5167,N_85,N_12);
nor U5168 (N_5168,N_3268,N_4053);
and U5169 (N_5169,N_2779,N_439);
and U5170 (N_5170,N_2332,N_3743);
xor U5171 (N_5171,N_4154,N_1700);
nor U5172 (N_5172,N_3907,N_4901);
nand U5173 (N_5173,N_3132,N_2751);
or U5174 (N_5174,N_365,N_3447);
xor U5175 (N_5175,N_1836,N_2174);
and U5176 (N_5176,N_438,N_2730);
and U5177 (N_5177,N_3564,N_550);
nand U5178 (N_5178,N_1073,N_3455);
or U5179 (N_5179,N_2306,N_613);
nand U5180 (N_5180,N_585,N_4136);
nor U5181 (N_5181,N_1917,N_1510);
or U5182 (N_5182,N_1233,N_3203);
xor U5183 (N_5183,N_4626,N_4644);
nand U5184 (N_5184,N_3623,N_2028);
or U5185 (N_5185,N_738,N_724);
and U5186 (N_5186,N_1479,N_1009);
or U5187 (N_5187,N_4670,N_2795);
and U5188 (N_5188,N_1012,N_1653);
and U5189 (N_5189,N_1628,N_735);
nand U5190 (N_5190,N_4183,N_1279);
nand U5191 (N_5191,N_4997,N_2266);
xor U5192 (N_5192,N_2759,N_3287);
nand U5193 (N_5193,N_2525,N_824);
xnor U5194 (N_5194,N_3728,N_4611);
nor U5195 (N_5195,N_938,N_4429);
xor U5196 (N_5196,N_3921,N_2139);
nor U5197 (N_5197,N_702,N_4780);
nor U5198 (N_5198,N_1593,N_2150);
or U5199 (N_5199,N_2548,N_1726);
and U5200 (N_5200,N_300,N_2347);
nand U5201 (N_5201,N_4510,N_2395);
nand U5202 (N_5202,N_4042,N_3840);
nand U5203 (N_5203,N_320,N_2475);
xnor U5204 (N_5204,N_4420,N_4668);
xnor U5205 (N_5205,N_3343,N_2900);
xor U5206 (N_5206,N_4142,N_3130);
or U5207 (N_5207,N_4925,N_4295);
nor U5208 (N_5208,N_3095,N_4367);
and U5209 (N_5209,N_3571,N_247);
nand U5210 (N_5210,N_1239,N_3525);
nand U5211 (N_5211,N_294,N_1786);
nor U5212 (N_5212,N_2868,N_395);
nand U5213 (N_5213,N_202,N_762);
and U5214 (N_5214,N_2472,N_2245);
nand U5215 (N_5215,N_4160,N_4023);
xor U5216 (N_5216,N_562,N_421);
nand U5217 (N_5217,N_2595,N_1922);
nand U5218 (N_5218,N_2662,N_3869);
or U5219 (N_5219,N_3256,N_526);
and U5220 (N_5220,N_1265,N_3875);
nand U5221 (N_5221,N_1509,N_1227);
xor U5222 (N_5222,N_1877,N_3607);
or U5223 (N_5223,N_1472,N_1523);
and U5224 (N_5224,N_4701,N_637);
and U5225 (N_5225,N_4041,N_4578);
nor U5226 (N_5226,N_3006,N_866);
xor U5227 (N_5227,N_1961,N_2378);
nand U5228 (N_5228,N_4092,N_3717);
xnor U5229 (N_5229,N_3558,N_351);
or U5230 (N_5230,N_3754,N_4487);
xnor U5231 (N_5231,N_928,N_3596);
or U5232 (N_5232,N_3839,N_1888);
or U5233 (N_5233,N_1111,N_2036);
nand U5234 (N_5234,N_2153,N_318);
nand U5235 (N_5235,N_1040,N_1838);
and U5236 (N_5236,N_4802,N_1406);
or U5237 (N_5237,N_3296,N_1102);
or U5238 (N_5238,N_4195,N_1195);
xor U5239 (N_5239,N_400,N_4902);
or U5240 (N_5240,N_3277,N_3850);
or U5241 (N_5241,N_184,N_249);
xnor U5242 (N_5242,N_902,N_3300);
or U5243 (N_5243,N_4903,N_212);
and U5244 (N_5244,N_2350,N_4170);
nor U5245 (N_5245,N_393,N_587);
xnor U5246 (N_5246,N_1988,N_3150);
nand U5247 (N_5247,N_1642,N_2483);
nor U5248 (N_5248,N_3977,N_3282);
xor U5249 (N_5249,N_549,N_51);
nand U5250 (N_5250,N_2321,N_1396);
nand U5251 (N_5251,N_1698,N_4642);
and U5252 (N_5252,N_4466,N_2453);
nand U5253 (N_5253,N_3135,N_3438);
nor U5254 (N_5254,N_1861,N_4763);
or U5255 (N_5255,N_389,N_4662);
and U5256 (N_5256,N_2033,N_1977);
nand U5257 (N_5257,N_1018,N_3170);
nor U5258 (N_5258,N_4098,N_4134);
nor U5259 (N_5259,N_3196,N_2115);
nor U5260 (N_5260,N_3252,N_2113);
or U5261 (N_5261,N_3278,N_4318);
or U5262 (N_5262,N_4753,N_2249);
nand U5263 (N_5263,N_2550,N_2878);
and U5264 (N_5264,N_1054,N_599);
or U5265 (N_5265,N_286,N_1675);
and U5266 (N_5266,N_388,N_3998);
xor U5267 (N_5267,N_4444,N_1104);
nor U5268 (N_5268,N_4707,N_2545);
or U5269 (N_5269,N_2193,N_2578);
xor U5270 (N_5270,N_3114,N_4872);
or U5271 (N_5271,N_2939,N_3534);
and U5272 (N_5272,N_4681,N_3916);
or U5273 (N_5273,N_2770,N_3267);
nand U5274 (N_5274,N_2990,N_2767);
or U5275 (N_5275,N_2058,N_3109);
xnor U5276 (N_5276,N_3538,N_245);
nand U5277 (N_5277,N_3612,N_4029);
nor U5278 (N_5278,N_1654,N_2604);
and U5279 (N_5279,N_885,N_1445);
nor U5280 (N_5280,N_2098,N_3696);
nand U5281 (N_5281,N_3679,N_3497);
nand U5282 (N_5282,N_3244,N_1332);
and U5283 (N_5283,N_818,N_1597);
nand U5284 (N_5284,N_4619,N_3249);
xor U5285 (N_5285,N_2375,N_1783);
and U5286 (N_5286,N_1604,N_4756);
nor U5287 (N_5287,N_1422,N_157);
xnor U5288 (N_5288,N_3159,N_1605);
nand U5289 (N_5289,N_4953,N_3302);
xor U5290 (N_5290,N_1666,N_572);
or U5291 (N_5291,N_3835,N_3482);
and U5292 (N_5292,N_2184,N_2745);
nand U5293 (N_5293,N_3094,N_840);
nand U5294 (N_5294,N_2064,N_1894);
xnor U5295 (N_5295,N_4566,N_682);
and U5296 (N_5296,N_4063,N_1292);
or U5297 (N_5297,N_259,N_3065);
nand U5298 (N_5298,N_2187,N_2589);
nor U5299 (N_5299,N_476,N_3970);
and U5300 (N_5300,N_1179,N_2959);
and U5301 (N_5301,N_648,N_2598);
xnor U5302 (N_5302,N_397,N_2642);
nand U5303 (N_5303,N_3652,N_3121);
nor U5304 (N_5304,N_3367,N_4502);
or U5305 (N_5305,N_2030,N_4333);
nand U5306 (N_5306,N_1724,N_4285);
or U5307 (N_5307,N_4513,N_177);
xnor U5308 (N_5308,N_495,N_1950);
or U5309 (N_5309,N_3326,N_656);
or U5310 (N_5310,N_1860,N_4723);
or U5311 (N_5311,N_4227,N_3259);
nor U5312 (N_5312,N_698,N_4361);
xor U5313 (N_5313,N_3923,N_24);
and U5314 (N_5314,N_3332,N_3904);
xor U5315 (N_5315,N_2482,N_263);
nand U5316 (N_5316,N_2613,N_3700);
or U5317 (N_5317,N_4692,N_2237);
xor U5318 (N_5318,N_588,N_4097);
or U5319 (N_5319,N_2117,N_1152);
xor U5320 (N_5320,N_367,N_2403);
or U5321 (N_5321,N_3541,N_4171);
or U5322 (N_5322,N_798,N_3688);
or U5323 (N_5323,N_845,N_621);
or U5324 (N_5324,N_1055,N_221);
nand U5325 (N_5325,N_3408,N_4458);
nand U5326 (N_5326,N_4749,N_3649);
xor U5327 (N_5327,N_2931,N_3957);
nand U5328 (N_5328,N_4291,N_4622);
xor U5329 (N_5329,N_3711,N_2712);
xnor U5330 (N_5330,N_558,N_929);
nor U5331 (N_5331,N_3663,N_3392);
nor U5332 (N_5332,N_3015,N_3156);
and U5333 (N_5333,N_4998,N_4703);
nor U5334 (N_5334,N_2217,N_1516);
nand U5335 (N_5335,N_862,N_848);
nor U5336 (N_5336,N_2966,N_4175);
or U5337 (N_5337,N_3264,N_2971);
nor U5338 (N_5338,N_2810,N_4271);
xor U5339 (N_5339,N_2913,N_1017);
xnor U5340 (N_5340,N_3544,N_3504);
or U5341 (N_5341,N_1809,N_3183);
nor U5342 (N_5342,N_3036,N_2691);
and U5343 (N_5343,N_3788,N_939);
and U5344 (N_5344,N_748,N_4082);
or U5345 (N_5345,N_4655,N_3604);
xor U5346 (N_5346,N_275,N_160);
nor U5347 (N_5347,N_1267,N_3131);
nor U5348 (N_5348,N_2491,N_690);
or U5349 (N_5349,N_3549,N_4169);
xnor U5350 (N_5350,N_886,N_3755);
and U5351 (N_5351,N_3242,N_291);
or U5352 (N_5352,N_4193,N_2128);
nand U5353 (N_5353,N_2081,N_3677);
or U5354 (N_5354,N_248,N_3443);
nor U5355 (N_5355,N_2327,N_219);
nor U5356 (N_5356,N_1513,N_2200);
and U5357 (N_5357,N_806,N_2474);
xnor U5358 (N_5358,N_543,N_3540);
or U5359 (N_5359,N_1699,N_3342);
and U5360 (N_5360,N_4714,N_2859);
xnor U5361 (N_5361,N_4439,N_2362);
and U5362 (N_5362,N_4044,N_3553);
xor U5363 (N_5363,N_3351,N_4830);
and U5364 (N_5364,N_125,N_209);
and U5365 (N_5365,N_1268,N_1757);
and U5366 (N_5366,N_3080,N_1282);
and U5367 (N_5367,N_57,N_1667);
nor U5368 (N_5368,N_3092,N_246);
nand U5369 (N_5369,N_3423,N_3585);
xor U5370 (N_5370,N_2738,N_3225);
xnor U5371 (N_5371,N_4575,N_238);
nand U5372 (N_5372,N_4261,N_2114);
nor U5373 (N_5373,N_4218,N_3417);
nand U5374 (N_5374,N_4446,N_2146);
and U5375 (N_5375,N_577,N_3703);
nand U5376 (N_5376,N_1840,N_4399);
nor U5377 (N_5377,N_354,N_657);
and U5378 (N_5378,N_4443,N_4697);
or U5379 (N_5379,N_4246,N_3985);
xnor U5380 (N_5380,N_4646,N_1049);
xor U5381 (N_5381,N_4100,N_321);
nor U5382 (N_5382,N_1237,N_3993);
and U5383 (N_5383,N_1606,N_3435);
nor U5384 (N_5384,N_4226,N_3237);
and U5385 (N_5385,N_1148,N_2546);
and U5386 (N_5386,N_3168,N_908);
xnor U5387 (N_5387,N_1201,N_3727);
xnor U5388 (N_5388,N_2369,N_1705);
and U5389 (N_5389,N_3273,N_4283);
nand U5390 (N_5390,N_2821,N_1945);
or U5391 (N_5391,N_2264,N_2554);
xnor U5392 (N_5392,N_1372,N_1355);
nor U5393 (N_5393,N_100,N_4584);
nor U5394 (N_5394,N_4754,N_528);
nor U5395 (N_5395,N_3782,N_2156);
xnor U5396 (N_5396,N_692,N_306);
nand U5397 (N_5397,N_1310,N_3429);
xor U5398 (N_5398,N_3556,N_3683);
xnor U5399 (N_5399,N_59,N_4352);
nor U5400 (N_5400,N_1426,N_461);
nor U5401 (N_5401,N_1327,N_854);
nand U5402 (N_5402,N_2422,N_611);
or U5403 (N_5403,N_2,N_2967);
nand U5404 (N_5404,N_3873,N_4077);
nand U5405 (N_5405,N_1057,N_1361);
nand U5406 (N_5406,N_2932,N_372);
and U5407 (N_5407,N_1067,N_1957);
nor U5408 (N_5408,N_3651,N_3773);
nand U5409 (N_5409,N_3557,N_802);
nand U5410 (N_5410,N_4667,N_1576);
nand U5411 (N_5411,N_4017,N_4602);
and U5412 (N_5412,N_853,N_746);
nor U5413 (N_5413,N_2848,N_4485);
xnor U5414 (N_5414,N_2594,N_2681);
and U5415 (N_5415,N_4543,N_1328);
nor U5416 (N_5416,N_3362,N_1377);
nand U5417 (N_5417,N_3298,N_831);
nand U5418 (N_5418,N_88,N_2487);
or U5419 (N_5419,N_1741,N_2085);
or U5420 (N_5420,N_3039,N_565);
nor U5421 (N_5421,N_4435,N_517);
or U5422 (N_5422,N_2011,N_1787);
nand U5423 (N_5423,N_1373,N_3999);
and U5424 (N_5424,N_3934,N_1482);
nor U5425 (N_5425,N_4883,N_4268);
and U5426 (N_5426,N_688,N_4617);
and U5427 (N_5427,N_548,N_2326);
or U5428 (N_5428,N_3348,N_3009);
xnor U5429 (N_5429,N_3910,N_1156);
nor U5430 (N_5430,N_4528,N_361);
xnor U5431 (N_5431,N_3153,N_2445);
xnor U5432 (N_5432,N_1418,N_162);
or U5433 (N_5433,N_4634,N_4201);
or U5434 (N_5434,N_4897,N_3802);
nand U5435 (N_5435,N_3308,N_4560);
and U5436 (N_5436,N_3263,N_4460);
xnor U5437 (N_5437,N_1680,N_3337);
nor U5438 (N_5438,N_1740,N_1481);
nor U5439 (N_5439,N_1972,N_2763);
and U5440 (N_5440,N_2399,N_2965);
nor U5441 (N_5441,N_1229,N_1703);
nand U5442 (N_5442,N_1315,N_3618);
or U5443 (N_5443,N_619,N_152);
nand U5444 (N_5444,N_1682,N_1764);
or U5445 (N_5445,N_3591,N_272);
and U5446 (N_5446,N_4165,N_477);
and U5447 (N_5447,N_2895,N_169);
nor U5448 (N_5448,N_3646,N_3548);
nand U5449 (N_5449,N_1424,N_2090);
and U5450 (N_5450,N_3994,N_2363);
xor U5451 (N_5451,N_3695,N_4741);
nand U5452 (N_5452,N_2209,N_491);
and U5453 (N_5453,N_2769,N_4067);
nand U5454 (N_5454,N_424,N_4032);
xor U5455 (N_5455,N_4228,N_750);
and U5456 (N_5456,N_683,N_914);
nand U5457 (N_5457,N_2372,N_118);
nor U5458 (N_5458,N_3295,N_3730);
nor U5459 (N_5459,N_1697,N_4069);
and U5460 (N_5460,N_3621,N_3990);
nor U5461 (N_5461,N_1739,N_2096);
nand U5462 (N_5462,N_2896,N_1349);
nor U5463 (N_5463,N_1540,N_1685);
nand U5464 (N_5464,N_1997,N_3146);
nand U5465 (N_5465,N_3486,N_113);
nand U5466 (N_5466,N_1927,N_4290);
and U5467 (N_5467,N_2439,N_4370);
nand U5468 (N_5468,N_3499,N_799);
xor U5469 (N_5469,N_4686,N_3178);
and U5470 (N_5470,N_4810,N_1109);
xor U5471 (N_5471,N_1579,N_176);
nor U5472 (N_5472,N_4920,N_817);
or U5473 (N_5473,N_4733,N_4861);
xor U5474 (N_5474,N_2083,N_258);
or U5475 (N_5475,N_2067,N_3317);
xnor U5476 (N_5476,N_2341,N_1598);
nand U5477 (N_5477,N_1347,N_3493);
and U5478 (N_5478,N_2801,N_2713);
nand U5479 (N_5479,N_131,N_1470);
and U5480 (N_5480,N_164,N_3336);
nand U5481 (N_5481,N_955,N_1723);
and U5482 (N_5482,N_2138,N_2783);
and U5483 (N_5483,N_2890,N_4350);
xnor U5484 (N_5484,N_3631,N_4968);
nand U5485 (N_5485,N_4132,N_1993);
or U5486 (N_5486,N_3953,N_801);
and U5487 (N_5487,N_1320,N_774);
and U5488 (N_5488,N_4220,N_3547);
or U5489 (N_5489,N_161,N_1302);
xnor U5490 (N_5490,N_4095,N_2458);
nor U5491 (N_5491,N_2335,N_1446);
and U5492 (N_5492,N_4540,N_4671);
or U5493 (N_5493,N_114,N_2619);
nand U5494 (N_5494,N_1543,N_2022);
nor U5495 (N_5495,N_2715,N_4314);
nand U5496 (N_5496,N_4094,N_2558);
and U5497 (N_5497,N_2618,N_485);
nor U5498 (N_5498,N_256,N_3202);
nand U5499 (N_5499,N_4815,N_3038);
and U5500 (N_5500,N_4060,N_4530);
and U5501 (N_5501,N_2084,N_4269);
xnor U5502 (N_5502,N_1880,N_1601);
nand U5503 (N_5503,N_4740,N_2933);
and U5504 (N_5504,N_1566,N_4989);
or U5505 (N_5505,N_2202,N_4596);
and U5506 (N_5506,N_255,N_3812);
xnor U5507 (N_5507,N_1360,N_129);
xnor U5508 (N_5508,N_2060,N_1011);
xor U5509 (N_5509,N_3007,N_3357);
or U5510 (N_5510,N_1351,N_534);
nand U5511 (N_5511,N_2236,N_4612);
xor U5512 (N_5512,N_3860,N_1317);
and U5513 (N_5513,N_3245,N_1219);
and U5514 (N_5514,N_1641,N_3657);
nand U5515 (N_5515,N_2218,N_3893);
or U5516 (N_5516,N_1975,N_768);
xnor U5517 (N_5517,N_4311,N_2072);
or U5518 (N_5518,N_2917,N_2701);
xnor U5519 (N_5519,N_1007,N_1839);
nor U5520 (N_5520,N_2749,N_2088);
or U5521 (N_5521,N_2864,N_575);
or U5522 (N_5522,N_1795,N_3089);
and U5523 (N_5523,N_4280,N_2969);
nand U5524 (N_5524,N_3761,N_4093);
nor U5525 (N_5525,N_4259,N_891);
xor U5526 (N_5526,N_1664,N_360);
xnor U5527 (N_5527,N_3961,N_1564);
or U5528 (N_5528,N_3037,N_18);
and U5529 (N_5529,N_2617,N_1557);
nand U5530 (N_5530,N_2826,N_881);
xor U5531 (N_5531,N_993,N_1693);
xnor U5532 (N_5532,N_1886,N_154);
or U5533 (N_5533,N_2814,N_218);
or U5534 (N_5534,N_379,N_4382);
and U5535 (N_5535,N_2232,N_2567);
xor U5536 (N_5536,N_1635,N_4991);
and U5537 (N_5537,N_4488,N_3609);
nor U5538 (N_5538,N_2127,N_576);
nor U5539 (N_5539,N_283,N_1097);
nor U5540 (N_5540,N_994,N_4351);
nand U5541 (N_5541,N_266,N_271);
and U5542 (N_5542,N_187,N_4794);
xnor U5543 (N_5543,N_1574,N_667);
xnor U5544 (N_5544,N_1618,N_155);
or U5545 (N_5545,N_2037,N_1497);
nand U5546 (N_5546,N_307,N_3718);
or U5547 (N_5547,N_2585,N_3948);
nand U5548 (N_5548,N_2302,N_1908);
xnor U5549 (N_5549,N_3891,N_4256);
xor U5550 (N_5550,N_2951,N_2380);
nor U5551 (N_5551,N_3390,N_3331);
and U5552 (N_5552,N_3741,N_163);
nor U5553 (N_5553,N_3480,N_972);
xnor U5554 (N_5554,N_4267,N_3783);
or U5555 (N_5555,N_1953,N_2787);
xor U5556 (N_5556,N_4221,N_3502);
xor U5557 (N_5557,N_3822,N_4993);
or U5558 (N_5558,N_4345,N_2695);
or U5559 (N_5559,N_3361,N_2112);
or U5560 (N_5560,N_231,N_377);
xnor U5561 (N_5561,N_1966,N_96);
and U5562 (N_5562,N_4640,N_1112);
nor U5563 (N_5563,N_3456,N_3026);
nand U5564 (N_5564,N_230,N_2666);
or U5565 (N_5565,N_1340,N_3537);
nor U5566 (N_5566,N_2056,N_3615);
xnor U5567 (N_5567,N_3262,N_1874);
nand U5568 (N_5568,N_1827,N_3966);
and U5569 (N_5569,N_1433,N_868);
xor U5570 (N_5570,N_658,N_211);
nand U5571 (N_5571,N_1824,N_1727);
and U5572 (N_5572,N_3592,N_1603);
and U5573 (N_5573,N_4820,N_2173);
nor U5574 (N_5574,N_3081,N_3177);
nor U5575 (N_5575,N_4659,N_573);
xnor U5576 (N_5576,N_3586,N_1989);
or U5577 (N_5577,N_2032,N_2446);
and U5578 (N_5578,N_4790,N_3391);
xnor U5579 (N_5579,N_3909,N_2998);
xor U5580 (N_5580,N_3285,N_3884);
or U5581 (N_5581,N_3368,N_650);
nor U5582 (N_5582,N_4529,N_2693);
and U5583 (N_5583,N_4661,N_1001);
xor U5584 (N_5584,N_139,N_4182);
xnor U5585 (N_5585,N_2734,N_2303);
nor U5586 (N_5586,N_1884,N_3676);
xor U5587 (N_5587,N_282,N_1170);
nand U5588 (N_5588,N_91,N_757);
nand U5589 (N_5589,N_4875,N_2886);
and U5590 (N_5590,N_4507,N_3712);
and U5591 (N_5591,N_1376,N_686);
nor U5592 (N_5592,N_4847,N_4406);
nand U5593 (N_5593,N_2640,N_2016);
or U5594 (N_5594,N_46,N_2093);
nor U5595 (N_5595,N_441,N_3945);
xor U5596 (N_5596,N_4112,N_2031);
or U5597 (N_5597,N_2576,N_4304);
or U5598 (N_5598,N_2556,N_4054);
nand U5599 (N_5599,N_2569,N_1923);
xnor U5600 (N_5600,N_375,N_1386);
xor U5601 (N_5601,N_1336,N_4893);
nor U5602 (N_5602,N_1688,N_4873);
or U5603 (N_5603,N_2387,N_1184);
nor U5604 (N_5604,N_3091,N_3494);
and U5605 (N_5605,N_4949,N_1910);
nor U5606 (N_5606,N_1980,N_1458);
and U5607 (N_5607,N_4755,N_1554);
xnor U5608 (N_5608,N_844,N_867);
xor U5609 (N_5609,N_334,N_2052);
nor U5610 (N_5610,N_4138,N_4139);
nand U5611 (N_5611,N_567,N_3902);
or U5612 (N_5612,N_226,N_4106);
and U5613 (N_5613,N_3995,N_257);
or U5614 (N_5614,N_4585,N_1059);
xnor U5615 (N_5615,N_1477,N_186);
nand U5616 (N_5616,N_530,N_3842);
nor U5617 (N_5617,N_4669,N_3501);
nand U5618 (N_5618,N_2935,N_4009);
or U5619 (N_5619,N_208,N_4947);
xnor U5620 (N_5620,N_1629,N_2504);
or U5621 (N_5621,N_841,N_4789);
and U5622 (N_5622,N_4103,N_4497);
xor U5623 (N_5623,N_4430,N_4784);
xnor U5624 (N_5624,N_2359,N_743);
nand U5625 (N_5625,N_728,N_244);
and U5626 (N_5626,N_3462,N_4180);
nor U5627 (N_5627,N_3349,N_2466);
nand U5628 (N_5628,N_1000,N_4932);
nand U5629 (N_5629,N_4804,N_4305);
nand U5630 (N_5630,N_2463,N_538);
nor U5631 (N_5631,N_4008,N_773);
nand U5632 (N_5632,N_4581,N_975);
or U5633 (N_5633,N_4588,N_720);
xor U5634 (N_5634,N_3376,N_789);
nor U5635 (N_5635,N_4595,N_1494);
and U5636 (N_5636,N_204,N_4533);
nand U5637 (N_5637,N_3846,N_1389);
xor U5638 (N_5638,N_1398,N_4571);
or U5639 (N_5639,N_416,N_2835);
xnor U5640 (N_5640,N_2515,N_2132);
and U5641 (N_5641,N_2885,N_1480);
nor U5642 (N_5642,N_4004,N_4484);
and U5643 (N_5643,N_1183,N_2631);
xnor U5644 (N_5644,N_4062,N_995);
xor U5645 (N_5645,N_2590,N_121);
and U5646 (N_5646,N_4599,N_1126);
xnor U5647 (N_5647,N_2658,N_3067);
and U5648 (N_5648,N_1425,N_697);
nor U5649 (N_5649,N_3485,N_4738);
or U5650 (N_5650,N_1412,N_4931);
or U5651 (N_5651,N_915,N_3396);
or U5652 (N_5652,N_409,N_4468);
nand U5653 (N_5653,N_3213,N_764);
nand U5654 (N_5654,N_2047,N_2852);
xor U5655 (N_5655,N_519,N_2526);
and U5656 (N_5656,N_425,N_1460);
nand U5657 (N_5657,N_4687,N_4313);
or U5658 (N_5658,N_4546,N_4411);
or U5659 (N_5659,N_1285,N_2930);
and U5660 (N_5660,N_1702,N_1679);
xor U5661 (N_5661,N_2710,N_2557);
and U5662 (N_5662,N_362,N_3536);
nor U5663 (N_5663,N_3102,N_3303);
nor U5664 (N_5664,N_2421,N_1171);
xor U5665 (N_5665,N_4570,N_4113);
nor U5666 (N_5666,N_2639,N_1578);
xnor U5667 (N_5667,N_726,N_3630);
or U5668 (N_5668,N_2632,N_1103);
nand U5669 (N_5669,N_4159,N_4278);
xor U5670 (N_5670,N_4391,N_2471);
nor U5671 (N_5671,N_1359,N_2145);
nor U5672 (N_5672,N_3468,N_2339);
xor U5673 (N_5673,N_2148,N_1047);
nor U5674 (N_5674,N_2807,N_3513);
and U5675 (N_5675,N_2988,N_786);
or U5676 (N_5676,N_2348,N_1665);
xnor U5677 (N_5677,N_4393,N_3057);
nand U5678 (N_5678,N_4120,N_2333);
nand U5679 (N_5679,N_1637,N_4561);
and U5680 (N_5680,N_2428,N_3316);
and U5681 (N_5681,N_4061,N_1083);
and U5682 (N_5682,N_1599,N_1094);
and U5683 (N_5683,N_115,N_1199);
nor U5684 (N_5684,N_822,N_3862);
nor U5685 (N_5685,N_297,N_312);
xor U5686 (N_5686,N_4957,N_668);
nand U5687 (N_5687,N_1455,N_2278);
xnor U5688 (N_5688,N_3100,N_2340);
nor U5689 (N_5689,N_1643,N_3885);
nor U5690 (N_5690,N_75,N_2162);
or U5691 (N_5691,N_77,N_1021);
and U5692 (N_5692,N_3704,N_4057);
xnor U5693 (N_5693,N_4675,N_2221);
or U5694 (N_5694,N_1488,N_4867);
or U5695 (N_5695,N_3883,N_4002);
nor U5696 (N_5696,N_4204,N_3925);
xnor U5697 (N_5697,N_3013,N_4556);
or U5698 (N_5698,N_3906,N_2660);
xor U5699 (N_5699,N_4459,N_4203);
or U5700 (N_5700,N_1182,N_4822);
nand U5701 (N_5701,N_1848,N_4544);
and U5702 (N_5702,N_14,N_2694);
and U5703 (N_5703,N_3290,N_268);
nand U5704 (N_5704,N_3474,N_1165);
xnor U5705 (N_5705,N_687,N_628);
or U5706 (N_5706,N_4292,N_1442);
nor U5707 (N_5707,N_4388,N_4735);
and U5708 (N_5708,N_4477,N_2989);
and U5709 (N_5709,N_3967,N_471);
nor U5710 (N_5710,N_205,N_4527);
nor U5711 (N_5711,N_3662,N_4791);
and U5712 (N_5712,N_857,N_1690);
or U5713 (N_5713,N_47,N_3120);
nand U5714 (N_5714,N_518,N_3247);
and U5715 (N_5715,N_1796,N_524);
nand U5716 (N_5716,N_3601,N_4200);
nand U5717 (N_5717,N_3859,N_4463);
xnor U5718 (N_5718,N_3573,N_240);
nand U5719 (N_5719,N_2130,N_2199);
nand U5720 (N_5720,N_3824,N_3466);
xor U5721 (N_5721,N_2802,N_384);
nand U5722 (N_5722,N_4688,N_3831);
nor U5723 (N_5723,N_796,N_4632);
or U5724 (N_5724,N_1454,N_251);
xnor U5725 (N_5725,N_4255,N_3236);
nor U5726 (N_5726,N_3112,N_4322);
nand U5727 (N_5727,N_4068,N_1329);
or U5728 (N_5728,N_3724,N_3809);
or U5729 (N_5729,N_3425,N_3313);
or U5730 (N_5730,N_3255,N_1232);
xor U5731 (N_5731,N_4482,N_3473);
or U5732 (N_5732,N_3402,N_951);
nor U5733 (N_5733,N_4603,N_107);
or U5734 (N_5734,N_420,N_4505);
and U5735 (N_5735,N_3753,N_3944);
or U5736 (N_5736,N_4337,N_4064);
nor U5737 (N_5737,N_1147,N_3275);
or U5738 (N_5738,N_2034,N_2762);
nor U5739 (N_5739,N_3561,N_1528);
and U5740 (N_5740,N_3694,N_1909);
nor U5741 (N_5741,N_2980,N_1397);
nor U5742 (N_5742,N_4736,N_2823);
xor U5743 (N_5743,N_2599,N_529);
xnor U5744 (N_5744,N_509,N_475);
nor U5745 (N_5745,N_4143,N_4058);
nor U5746 (N_5746,N_148,N_1843);
or U5747 (N_5747,N_3224,N_561);
and U5748 (N_5748,N_681,N_1420);
nor U5749 (N_5749,N_2874,N_3629);
or U5750 (N_5750,N_2602,N_1985);
nand U5751 (N_5751,N_1911,N_2087);
nand U5752 (N_5752,N_3658,N_3137);
nor U5753 (N_5753,N_4975,N_4911);
nor U5754 (N_5754,N_339,N_1781);
nor U5755 (N_5755,N_4704,N_3426);
nand U5756 (N_5756,N_2419,N_3004);
xor U5757 (N_5757,N_3416,N_858);
and U5758 (N_5758,N_1345,N_4018);
xnor U5759 (N_5759,N_1525,N_287);
xnor U5760 (N_5760,N_3072,N_3174);
and U5761 (N_5761,N_912,N_1873);
xor U5762 (N_5762,N_3739,N_390);
or U5763 (N_5763,N_3433,N_3445);
nor U5764 (N_5764,N_4198,N_3241);
xnor U5765 (N_5765,N_3903,N_328);
nor U5766 (N_5766,N_1969,N_2853);
nor U5767 (N_5767,N_1612,N_3584);
xor U5768 (N_5768,N_3415,N_4951);
nor U5769 (N_5769,N_713,N_2503);
nand U5770 (N_5770,N_2568,N_2608);
nor U5771 (N_5771,N_1378,N_2519);
nand U5772 (N_5772,N_4312,N_1501);
and U5773 (N_5773,N_2597,N_4624);
xnor U5774 (N_5774,N_2337,N_2812);
nand U5775 (N_5775,N_4765,N_777);
or U5776 (N_5776,N_2296,N_3436);
nor U5777 (N_5777,N_153,N_4614);
or U5778 (N_5778,N_1444,N_3803);
nand U5779 (N_5779,N_1485,N_1529);
nand U5780 (N_5780,N_4874,N_4078);
or U5781 (N_5781,N_1451,N_4938);
nor U5782 (N_5782,N_4958,N_2746);
xor U5783 (N_5783,N_4685,N_2953);
nand U5784 (N_5784,N_2893,N_2477);
xor U5785 (N_5785,N_4731,N_1714);
and U5786 (N_5786,N_4977,N_3371);
or U5787 (N_5787,N_2371,N_4114);
and U5788 (N_5788,N_143,N_1167);
nand U5789 (N_5789,N_3246,N_3470);
or U5790 (N_5790,N_3689,N_415);
nor U5791 (N_5791,N_4623,N_1240);
nand U5792 (N_5792,N_1381,N_4070);
xor U5793 (N_5793,N_2178,N_2100);
and U5794 (N_5794,N_4964,N_4177);
or U5795 (N_5795,N_863,N_3933);
or U5796 (N_5796,N_1234,N_2524);
and U5797 (N_5797,N_445,N_1251);
and U5798 (N_5798,N_4242,N_2905);
and U5799 (N_5799,N_4462,N_3108);
xnor U5800 (N_5800,N_4678,N_3791);
xor U5801 (N_5801,N_1651,N_4628);
nand U5802 (N_5802,N_2797,N_2884);
nor U5803 (N_5803,N_2542,N_1298);
nor U5804 (N_5804,N_3817,N_1335);
nand U5805 (N_5805,N_1294,N_4557);
xnor U5806 (N_5806,N_4757,N_1410);
nor U5807 (N_5807,N_569,N_4816);
xnor U5808 (N_5808,N_783,N_52);
xnor U5809 (N_5809,N_3077,N_4751);
nor U5810 (N_5810,N_498,N_2772);
xor U5811 (N_5811,N_3233,N_337);
or U5812 (N_5812,N_1062,N_3397);
or U5813 (N_5813,N_4438,N_4192);
nor U5814 (N_5814,N_3806,N_4641);
nand U5815 (N_5815,N_2451,N_1568);
xor U5816 (N_5816,N_4479,N_984);
nor U5817 (N_5817,N_2004,N_763);
nand U5818 (N_5818,N_2241,N_363);
or U5819 (N_5819,N_3971,N_2079);
nand U5820 (N_5820,N_791,N_3119);
and U5821 (N_5821,N_731,N_804);
or U5822 (N_5822,N_4110,N_604);
nor U5823 (N_5823,N_4574,N_941);
nor U5824 (N_5824,N_4467,N_1711);
nor U5825 (N_5825,N_766,N_4338);
xor U5826 (N_5826,N_2771,N_3031);
or U5827 (N_5827,N_566,N_3048);
or U5828 (N_5828,N_4185,N_1948);
or U5829 (N_5829,N_1552,N_4604);
xnor U5830 (N_5830,N_3771,N_3284);
or U5831 (N_5831,N_3968,N_4715);
nand U5832 (N_5832,N_1402,N_166);
or U5833 (N_5833,N_1042,N_2764);
xor U5834 (N_5834,N_4620,N_1290);
and U5835 (N_5835,N_4744,N_3071);
and U5836 (N_5836,N_1504,N_4207);
nand U5837 (N_5837,N_4856,N_2902);
nor U5838 (N_5838,N_1287,N_2508);
xor U5839 (N_5839,N_4364,N_3605);
or U5840 (N_5840,N_4349,N_358);
or U5841 (N_5841,N_3587,N_4580);
and U5842 (N_5842,N_170,N_4638);
or U5843 (N_5843,N_290,N_3437);
or U5844 (N_5844,N_1357,N_469);
or U5845 (N_5845,N_4888,N_856);
xnor U5846 (N_5846,N_2962,N_537);
or U5847 (N_5847,N_649,N_2338);
and U5848 (N_5848,N_664,N_1056);
xnor U5849 (N_5849,N_1849,N_2683);
nor U5850 (N_5850,N_4955,N_3424);
or U5851 (N_5851,N_4627,N_1196);
nand U5852 (N_5852,N_191,N_373);
and U5853 (N_5853,N_1684,N_4592);
or U5854 (N_5854,N_2668,N_4840);
xnor U5855 (N_5855,N_3309,N_2538);
nor U5856 (N_5856,N_3010,N_795);
xor U5857 (N_5857,N_736,N_4555);
and U5858 (N_5858,N_4357,N_4144);
nand U5859 (N_5859,N_3315,N_1943);
nand U5860 (N_5860,N_4190,N_4248);
or U5861 (N_5861,N_4408,N_3230);
nor U5862 (N_5862,N_4022,N_4265);
or U5863 (N_5863,N_1982,N_622);
or U5864 (N_5864,N_4649,N_535);
and U5865 (N_5865,N_1044,N_216);
and U5866 (N_5866,N_4086,N_4954);
or U5867 (N_5867,N_4445,N_1575);
xor U5868 (N_5868,N_4868,N_563);
xor U5869 (N_5869,N_1155,N_3567);
and U5870 (N_5870,N_2078,N_429);
nand U5871 (N_5871,N_3341,N_1393);
nor U5872 (N_5872,N_1800,N_4301);
nand U5873 (N_5873,N_4848,N_1617);
nand U5874 (N_5874,N_2459,N_4838);
nand U5875 (N_5875,N_1258,N_2514);
nor U5876 (N_5876,N_4940,N_1569);
and U5877 (N_5877,N_2761,N_1058);
nor U5878 (N_5878,N_4859,N_842);
and U5879 (N_5879,N_1938,N_4263);
or U5880 (N_5880,N_1533,N_4776);
nand U5881 (N_5881,N_2448,N_3643);
nor U5882 (N_5882,N_484,N_3531);
xnor U5883 (N_5883,N_3642,N_3637);
xor U5884 (N_5884,N_2914,N_1819);
nor U5885 (N_5885,N_1123,N_2300);
nand U5886 (N_5886,N_1421,N_3257);
and U5887 (N_5887,N_4341,N_4962);
nand U5888 (N_5888,N_3191,N_4233);
nor U5889 (N_5889,N_4724,N_1158);
or U5890 (N_5890,N_508,N_1520);
nor U5891 (N_5891,N_4066,N_2727);
xnor U5892 (N_5892,N_482,N_1273);
or U5893 (N_5893,N_3404,N_3118);
nor U5894 (N_5894,N_274,N_1272);
nand U5895 (N_5895,N_369,N_3281);
nand U5896 (N_5896,N_4785,N_4084);
nor U5897 (N_5897,N_3490,N_1356);
and U5898 (N_5898,N_627,N_138);
xor U5899 (N_5899,N_86,N_3350);
nor U5900 (N_5900,N_3590,N_344);
nand U5901 (N_5901,N_413,N_48);
and U5902 (N_5902,N_2984,N_1429);
nand U5903 (N_5903,N_1986,N_4939);
and U5904 (N_5904,N_4385,N_2943);
xor U5905 (N_5905,N_544,N_899);
and U5906 (N_5906,N_189,N_3411);
or U5907 (N_5907,N_3723,N_876);
nor U5908 (N_5908,N_1363,N_3726);
nand U5909 (N_5909,N_1416,N_2588);
nand U5910 (N_5910,N_923,N_2136);
nor U5911 (N_5911,N_2455,N_2685);
nand U5912 (N_5912,N_194,N_182);
nand U5913 (N_5913,N_600,N_2600);
xor U5914 (N_5914,N_1792,N_501);
or U5915 (N_5915,N_2839,N_3395);
nor U5916 (N_5916,N_2134,N_2481);
and U5917 (N_5917,N_3511,N_874);
and U5918 (N_5918,N_4682,N_2665);
xor U5919 (N_5919,N_872,N_1745);
xnor U5920 (N_5920,N_4329,N_2726);
and U5921 (N_5921,N_3896,N_584);
nor U5922 (N_5922,N_1625,N_870);
nand U5923 (N_5923,N_3503,N_1857);
and U5924 (N_5924,N_2396,N_3154);
xnor U5925 (N_5925,N_1297,N_496);
and U5926 (N_5926,N_4717,N_8);
or U5927 (N_5927,N_1992,N_4384);
nand U5928 (N_5928,N_2898,N_2478);
nand U5929 (N_5929,N_1197,N_3519);
xnor U5930 (N_5930,N_285,N_4270);
xor U5931 (N_5931,N_3705,N_4206);
nor U5932 (N_5932,N_4922,N_3670);
or U5933 (N_5933,N_2142,N_1715);
and U5934 (N_5934,N_1291,N_3597);
xnor U5935 (N_5935,N_1657,N_2706);
nor U5936 (N_5936,N_2756,N_578);
xnor U5937 (N_5937,N_2025,N_4734);
and U5938 (N_5938,N_606,N_4421);
and U5939 (N_5939,N_1262,N_1817);
xor U5940 (N_5940,N_1423,N_983);
nor U5941 (N_5941,N_2551,N_1385);
nand U5942 (N_5942,N_175,N_3410);
or U5943 (N_5943,N_428,N_4817);
nand U5944 (N_5944,N_3595,N_3975);
xnor U5945 (N_5945,N_2440,N_849);
xnor U5946 (N_5946,N_758,N_986);
xnor U5947 (N_5947,N_634,N_4133);
or U5948 (N_5948,N_403,N_3314);
and U5949 (N_5949,N_3889,N_1374);
nand U5950 (N_5950,N_1008,N_2728);
nor U5951 (N_5951,N_3144,N_1511);
and U5952 (N_5952,N_2690,N_2825);
and U5953 (N_5953,N_3028,N_1143);
and U5954 (N_5954,N_4605,N_2506);
or U5955 (N_5955,N_2915,N_2647);
nor U5956 (N_5956,N_2938,N_3211);
nor U5957 (N_5957,N_2111,N_1793);
and U5958 (N_5958,N_3058,N_3805);
xnor U5959 (N_5959,N_1616,N_540);
or U5960 (N_5960,N_1085,N_4716);
nand U5961 (N_5961,N_2256,N_4331);
xnor U5962 (N_5962,N_3890,N_1725);
xnor U5963 (N_5963,N_2377,N_3340);
or U5964 (N_5964,N_3509,N_3867);
nor U5965 (N_5965,N_3145,N_3450);
xor U5966 (N_5966,N_4808,N_3943);
xor U5967 (N_5967,N_56,N_1048);
or U5968 (N_5968,N_1539,N_3858);
nand U5969 (N_5969,N_4645,N_2881);
and U5970 (N_5970,N_3227,N_4725);
nor U5971 (N_5971,N_3815,N_4205);
nor U5972 (N_5972,N_3528,N_2204);
nand U5973 (N_5973,N_1934,N_4011);
nand U5974 (N_5974,N_4935,N_3864);
and U5975 (N_5975,N_2423,N_2454);
or U5976 (N_5976,N_3749,N_797);
and U5977 (N_5977,N_2029,N_2684);
nand U5978 (N_5978,N_1489,N_3354);
or U5979 (N_5979,N_2616,N_2406);
nor U5980 (N_5980,N_2541,N_739);
nor U5981 (N_5981,N_1146,N_3087);
or U5982 (N_5982,N_1766,N_4400);
and U5983 (N_5983,N_3234,N_940);
nor U5984 (N_5984,N_1210,N_1092);
or U5985 (N_5985,N_593,N_3160);
nor U5986 (N_5986,N_2871,N_1522);
or U5987 (N_5987,N_765,N_1695);
nor U5988 (N_5988,N_3175,N_1981);
xnor U5989 (N_5989,N_3543,N_2832);
and U5990 (N_5990,N_3816,N_1086);
nor U5991 (N_5991,N_2437,N_761);
xnor U5992 (N_5992,N_1333,N_214);
xnor U5993 (N_5993,N_4650,N_4801);
xnor U5994 (N_5994,N_4517,N_2614);
nand U5995 (N_5995,N_1390,N_1771);
nand U5996 (N_5996,N_3576,N_2901);
nand U5997 (N_5997,N_3271,N_239);
and U5998 (N_5998,N_1288,N_3451);
nor U5999 (N_5999,N_2766,N_3489);
and U6000 (N_6000,N_2982,N_1648);
xor U6001 (N_6001,N_1431,N_1850);
nand U6002 (N_6002,N_1813,N_4690);
or U6003 (N_6003,N_1537,N_3002);
nor U6004 (N_6004,N_1250,N_2974);
nand U6005 (N_6005,N_2531,N_2842);
nor U6006 (N_6006,N_322,N_4891);
xor U6007 (N_6007,N_1707,N_4038);
xnor U6008 (N_6008,N_4519,N_788);
nor U6009 (N_6009,N_2325,N_1428);
or U6010 (N_6010,N_4179,N_2792);
and U6011 (N_6011,N_4470,N_2648);
nor U6012 (N_6012,N_3589,N_1069);
or U6013 (N_6013,N_2334,N_3373);
xor U6014 (N_6014,N_94,N_3882);
xor U6015 (N_6015,N_4,N_55);
and U6016 (N_6016,N_2747,N_3322);
and U6017 (N_6017,N_2841,N_1776);
and U6018 (N_6018,N_4176,N_228);
or U6019 (N_6019,N_1474,N_3760);
and U6020 (N_6020,N_359,N_4966);
or U6021 (N_6021,N_2818,N_734);
nand U6022 (N_6022,N_1713,N_3871);
nor U6023 (N_6023,N_2601,N_1777);
or U6024 (N_6024,N_3034,N_3675);
nand U6025 (N_6025,N_3363,N_442);
or U6026 (N_6026,N_3301,N_996);
or U6027 (N_6027,N_2803,N_579);
and U6028 (N_6028,N_456,N_1563);
and U6029 (N_6029,N_1636,N_4324);
or U6030 (N_6030,N_4796,N_1391);
or U6031 (N_6031,N_2285,N_3625);
nor U6032 (N_6032,N_4141,N_3063);
nor U6033 (N_6033,N_444,N_532);
nand U6034 (N_6034,N_759,N_564);
or U6035 (N_6035,N_2782,N_3421);
or U6036 (N_6036,N_1627,N_3111);
or U6037 (N_6037,N_4450,N_449);
nor U6038 (N_6038,N_3866,N_4520);
nor U6039 (N_6039,N_3166,N_1941);
nor U6040 (N_6040,N_2829,N_4216);
xnor U6041 (N_6041,N_3691,N_3116);
and U6042 (N_6042,N_2680,N_4075);
nand U6043 (N_6043,N_2316,N_3706);
or U6044 (N_6044,N_3060,N_3616);
or U6045 (N_6045,N_2789,N_2622);
or U6046 (N_6046,N_3205,N_1280);
nor U6047 (N_6047,N_2008,N_1077);
or U6048 (N_6048,N_3787,N_976);
and U6049 (N_6049,N_4249,N_835);
or U6050 (N_6050,N_4824,N_3664);
or U6051 (N_6051,N_3918,N_3976);
nor U6052 (N_6052,N_1769,N_2833);
or U6053 (N_6053,N_4178,N_4047);
nand U6054 (N_6054,N_823,N_4672);
and U6055 (N_6055,N_1125,N_2345);
nor U6056 (N_6056,N_4635,N_971);
or U6057 (N_6057,N_1999,N_1116);
nor U6058 (N_6058,N_2404,N_1177);
xor U6059 (N_6059,N_352,N_2317);
xor U6060 (N_6060,N_2432,N_236);
or U6061 (N_6061,N_1205,N_4210);
or U6062 (N_6062,N_1066,N_2354);
or U6063 (N_6063,N_631,N_1252);
xor U6064 (N_6064,N_4866,N_225);
nor U6065 (N_6065,N_610,N_6);
nand U6066 (N_6066,N_4684,N_298);
or U6067 (N_6067,N_3699,N_3280);
nand U6068 (N_6068,N_3857,N_1990);
or U6069 (N_6069,N_839,N_3555);
and U6070 (N_6070,N_1744,N_3745);
nand U6071 (N_6071,N_3856,N_253);
xnor U6072 (N_6072,N_3000,N_2261);
nor U6073 (N_6073,N_2987,N_151);
nand U6074 (N_6074,N_4912,N_3678);
nor U6075 (N_6075,N_92,N_2426);
nor U6076 (N_6076,N_1050,N_838);
nand U6077 (N_6077,N_1362,N_3453);
nand U6078 (N_6078,N_580,N_478);
or U6079 (N_6079,N_1716,N_4434);
nand U6080 (N_6080,N_516,N_2040);
and U6081 (N_6081,N_2645,N_4793);
and U6082 (N_6082,N_4432,N_4116);
nor U6083 (N_6083,N_1865,N_3659);
and U6084 (N_6084,N_655,N_4996);
or U6085 (N_6085,N_4918,N_1099);
and U6086 (N_6086,N_1319,N_3622);
xor U6087 (N_6087,N_1249,N_3345);
nand U6088 (N_6088,N_913,N_2313);
nand U6089 (N_6089,N_1942,N_1122);
and U6090 (N_6090,N_1266,N_2006);
xnor U6091 (N_6091,N_2160,N_4960);
nand U6092 (N_6092,N_1241,N_3110);
or U6093 (N_6093,N_591,N_2141);
and U6094 (N_6094,N_2869,N_1916);
and U6095 (N_6095,N_730,N_1514);
nand U6096 (N_6096,N_1672,N_4980);
and U6097 (N_6097,N_4262,N_521);
and U6098 (N_6098,N_4309,N_3358);
xor U6099 (N_6099,N_685,N_4403);
or U6100 (N_6100,N_3082,N_2502);
or U6101 (N_6101,N_2671,N_1919);
or U6102 (N_6102,N_4320,N_3818);
or U6103 (N_6103,N_1869,N_2652);
or U6104 (N_6104,N_1996,N_34);
and U6105 (N_6105,N_326,N_3766);
or U6106 (N_6106,N_3199,N_371);
and U6107 (N_6107,N_4712,N_583);
nor U6108 (N_6108,N_1737,N_3492);
nand U6109 (N_6109,N_4260,N_948);
and U6110 (N_6110,N_1202,N_4188);
and U6111 (N_6111,N_4708,N_4274);
or U6112 (N_6112,N_4702,N_1300);
xor U6113 (N_6113,N_1935,N_4914);
nor U6114 (N_6114,N_2675,N_2046);
nand U6115 (N_6115,N_2867,N_590);
nor U6116 (N_6116,N_546,N_1778);
or U6117 (N_6117,N_4151,N_2678);
xor U6118 (N_6118,N_65,N_4639);
and U6119 (N_6119,N_3073,N_1548);
and U6120 (N_6120,N_458,N_1613);
or U6121 (N_6121,N_4071,N_102);
nand U6122 (N_6122,N_3989,N_2768);
or U6123 (N_6123,N_2368,N_4244);
or U6124 (N_6124,N_1663,N_1382);
xnor U6125 (N_6125,N_2168,N_423);
nand U6126 (N_6126,N_1022,N_2563);
nor U6127 (N_6127,N_3047,N_4489);
nand U6128 (N_6128,N_3216,N_2172);
nor U6129 (N_6129,N_4166,N_1076);
nand U6130 (N_6130,N_850,N_2863);
or U6131 (N_6131,N_1765,N_54);
xnor U6132 (N_6132,N_1400,N_3562);
nor U6133 (N_6133,N_4948,N_241);
or U6134 (N_6134,N_4355,N_4928);
nand U6135 (N_6135,N_4279,N_4001);
or U6136 (N_6136,N_3033,N_1499);
or U6137 (N_6137,N_327,N_1856);
xnor U6138 (N_6138,N_553,N_3475);
and U6139 (N_6139,N_2125,N_4821);
nor U6140 (N_6140,N_4509,N_3248);
or U6141 (N_6141,N_917,N_1991);
nor U6142 (N_6142,N_999,N_3339);
and U6143 (N_6143,N_4535,N_527);
and U6144 (N_6144,N_488,N_2672);
xnor U6145 (N_6145,N_4783,N_2583);
and U6146 (N_6146,N_3905,N_727);
or U6147 (N_6147,N_1091,N_1678);
nor U6148 (N_6148,N_1107,N_3133);
nor U6149 (N_6149,N_4904,N_4155);
and U6150 (N_6150,N_1016,N_4721);
and U6151 (N_6151,N_1570,N_217);
nor U6152 (N_6152,N_3046,N_1435);
nand U6153 (N_6153,N_2397,N_2805);
xor U6154 (N_6154,N_3554,N_4496);
and U6155 (N_6155,N_742,N_3461);
and U6156 (N_6156,N_3365,N_2057);
nand U6157 (N_6157,N_3229,N_3956);
xnor U6158 (N_6158,N_3129,N_708);
or U6159 (N_6159,N_1939,N_1452);
xnor U6160 (N_6160,N_2941,N_1209);
nor U6161 (N_6161,N_2225,N_2208);
or U6162 (N_6162,N_109,N_1689);
nand U6163 (N_6163,N_4750,N_2283);
and U6164 (N_6164,N_1732,N_1788);
or U6165 (N_6165,N_1565,N_1964);
xnor U6166 (N_6166,N_2641,N_836);
xor U6167 (N_6167,N_1166,N_1163);
xor U6168 (N_6168,N_4569,N_2161);
nand U6169 (N_6169,N_4157,N_2053);
or U6170 (N_6170,N_4910,N_122);
and U6171 (N_6171,N_4764,N_4414);
or U6172 (N_6172,N_1581,N_4946);
or U6173 (N_6173,N_3157,N_407);
nand U6174 (N_6174,N_436,N_452);
or U6175 (N_6175,N_3915,N_2827);
and U6176 (N_6176,N_3644,N_4287);
nor U6177 (N_6177,N_144,N_828);
or U6178 (N_6178,N_2919,N_4225);
xnor U6179 (N_6179,N_3193,N_2534);
xnor U6180 (N_6180,N_4108,N_4035);
or U6181 (N_6181,N_3722,N_2222);
xor U6182 (N_6182,N_4590,N_2310);
or U6183 (N_6183,N_3834,N_2244);
nor U6184 (N_6184,N_1255,N_53);
nand U6185 (N_6185,N_196,N_4158);
xnor U6186 (N_6186,N_3522,N_3735);
nand U6187 (N_6187,N_1223,N_1150);
or U6188 (N_6188,N_665,N_4526);
xor U6189 (N_6189,N_2465,N_4722);
xnor U6190 (N_6190,N_1231,N_1465);
and U6191 (N_6191,N_1380,N_4237);
nor U6192 (N_6192,N_3958,N_1638);
nor U6193 (N_6193,N_3865,N_3184);
nand U6194 (N_6194,N_700,N_3223);
and U6195 (N_6195,N_1906,N_4524);
and U6196 (N_6196,N_3018,N_531);
or U6197 (N_6197,N_2412,N_651);
xor U6198 (N_6198,N_2572,N_935);
and U6199 (N_6199,N_4039,N_1119);
nand U6200 (N_6200,N_2501,N_1096);
xnor U6201 (N_6201,N_135,N_2092);
or U6202 (N_6202,N_1023,N_878);
xnor U6203 (N_6203,N_4896,N_2781);
nand U6204 (N_6204,N_2386,N_4440);
or U6205 (N_6205,N_3085,N_4819);
xnor U6206 (N_6206,N_4969,N_473);
xor U6207 (N_6207,N_2636,N_2985);
or U6208 (N_6208,N_3532,N_769);
or U6209 (N_6209,N_988,N_1928);
xor U6210 (N_6210,N_3942,N_1005);
xor U6211 (N_6211,N_618,N_4074);
nand U6212 (N_6212,N_4814,N_1006);
xnor U6213 (N_6213,N_4583,N_3292);
nor U6214 (N_6214,N_2182,N_966);
and U6215 (N_6215,N_3320,N_1028);
xnor U6216 (N_6216,N_2013,N_1440);
nand U6217 (N_6217,N_1128,N_4806);
nand U6218 (N_6218,N_3746,N_4354);
nor U6219 (N_6219,N_133,N_1591);
or U6220 (N_6220,N_2840,N_3539);
and U6221 (N_6221,N_1395,N_200);
or U6222 (N_6222,N_3003,N_2963);
and U6223 (N_6223,N_4398,N_4149);
and U6224 (N_6224,N_4286,N_2044);
and U6225 (N_6225,N_2942,N_4876);
nor U6226 (N_6226,N_2082,N_670);
nor U6227 (N_6227,N_615,N_1113);
or U6228 (N_6228,N_4552,N_1464);
or U6229 (N_6229,N_3982,N_826);
and U6230 (N_6230,N_2231,N_2536);
nand U6231 (N_6231,N_3495,N_2836);
nand U6232 (N_6232,N_689,N_2643);
and U6233 (N_6233,N_136,N_4030);
nand U6234 (N_6234,N_1517,N_1161);
and U6235 (N_6235,N_1098,N_954);
and U6236 (N_6236,N_4547,N_1221);
and U6237 (N_6237,N_4402,N_4972);
nor U6238 (N_6238,N_992,N_3877);
and U6239 (N_6239,N_1493,N_3062);
xor U6240 (N_6240,N_1518,N_1900);
xor U6241 (N_6241,N_910,N_3617);
nor U6242 (N_6242,N_376,N_4202);
xnor U6243 (N_6243,N_2255,N_2108);
nor U6244 (N_6244,N_3825,N_693);
and U6245 (N_6245,N_3950,N_2151);
and U6246 (N_6246,N_4012,N_3093);
xnor U6247 (N_6247,N_3800,N_1145);
or U6248 (N_6248,N_924,N_943);
or U6249 (N_6249,N_2581,N_3693);
and U6250 (N_6250,N_2394,N_4568);
nand U6251 (N_6251,N_847,N_3117);
and U6252 (N_6252,N_725,N_234);
or U6253 (N_6253,N_2997,N_402);
or U6254 (N_6254,N_3901,N_178);
xor U6255 (N_6255,N_2293,N_3790);
xnor U6256 (N_6256,N_292,N_470);
and U6257 (N_6257,N_2644,N_2281);
xor U6258 (N_6258,N_4752,N_4913);
xor U6259 (N_6259,N_1106,N_792);
nand U6260 (N_6260,N_1872,N_2784);
or U6261 (N_6261,N_3823,N_466);
and U6262 (N_6262,N_1248,N_270);
xnor U6263 (N_6263,N_3991,N_2177);
nand U6264 (N_6264,N_181,N_560);
and U6265 (N_6265,N_2328,N_629);
or U6266 (N_6266,N_1556,N_982);
or U6267 (N_6267,N_1828,N_1450);
nor U6268 (N_6268,N_1437,N_350);
and U6269 (N_6269,N_341,N_4926);
nand U6270 (N_6270,N_4831,N_4636);
nor U6271 (N_6271,N_3192,N_3550);
nand U6272 (N_6272,N_103,N_2346);
or U6273 (N_6273,N_4857,N_4240);
or U6274 (N_6274,N_3400,N_504);
or U6275 (N_6275,N_2407,N_3731);
nor U6276 (N_6276,N_4072,N_752);
nand U6277 (N_6277,N_2398,N_3572);
nor U6278 (N_6278,N_793,N_4521);
nand U6279 (N_6279,N_3066,N_2849);
and U6280 (N_6280,N_1095,N_3533);
nand U6281 (N_6281,N_3327,N_880);
xor U6282 (N_6282,N_3140,N_2263);
xor U6283 (N_6283,N_1341,N_3757);
nor U6284 (N_6284,N_3032,N_3829);
nand U6285 (N_6285,N_1032,N_3720);
nor U6286 (N_6286,N_41,N_4453);
nor U6287 (N_6287,N_1101,N_4378);
xor U6288 (N_6288,N_633,N_1129);
and U6289 (N_6289,N_3147,N_2741);
nand U6290 (N_6290,N_2343,N_4990);
or U6291 (N_6291,N_1138,N_596);
nor U6292 (N_6292,N_947,N_1907);
nand U6293 (N_6293,N_3775,N_4597);
xnor U6294 (N_6294,N_669,N_3512);
nor U6295 (N_6295,N_571,N_4630);
or U6296 (N_6296,N_93,N_4936);
nor U6297 (N_6297,N_38,N_3020);
or U6298 (N_6298,N_4330,N_2314);
nor U6299 (N_6299,N_964,N_2299);
or U6300 (N_6300,N_1185,N_2374);
nor U6301 (N_6301,N_1010,N_1862);
nor U6302 (N_6302,N_2571,N_2215);
nor U6303 (N_6303,N_4247,N_4359);
nor U6304 (N_6304,N_4377,N_4371);
or U6305 (N_6305,N_4492,N_718);
or U6306 (N_6306,N_4409,N_1920);
xnor U6307 (N_6307,N_2564,N_3215);
nand U6308 (N_6308,N_1936,N_4860);
or U6309 (N_6309,N_2301,N_696);
nand U6310 (N_6310,N_1696,N_2268);
or U6311 (N_6311,N_4898,N_4709);
or U6312 (N_6312,N_1330,N_2068);
and U6313 (N_6313,N_3090,N_4746);
nand U6314 (N_6314,N_3,N_1259);
nor U6315 (N_6315,N_2800,N_3105);
nand U6316 (N_6316,N_2183,N_998);
xor U6317 (N_6317,N_4959,N_366);
nor U6318 (N_6318,N_4973,N_815);
xor U6319 (N_6319,N_3454,N_2494);
or U6320 (N_6320,N_4389,N_779);
and U6321 (N_6321,N_3624,N_4043);
xor U6322 (N_6322,N_4737,N_4909);
nor U6323 (N_6323,N_4726,N_1090);
nand U6324 (N_6324,N_3797,N_2687);
xnor U6325 (N_6325,N_2365,N_2861);
xor U6326 (N_6326,N_2039,N_2846);
nor U6327 (N_6327,N_2948,N_542);
or U6328 (N_6328,N_3796,N_3476);
and U6329 (N_6329,N_412,N_2819);
nor U6330 (N_6330,N_1293,N_4115);
nor U6331 (N_6331,N_489,N_785);
or U6332 (N_6332,N_4615,N_2270);
nor U6333 (N_6333,N_3813,N_1020);
or U6334 (N_6334,N_1334,N_1947);
and U6335 (N_6335,N_2157,N_620);
or U6336 (N_6336,N_1045,N_3774);
or U6337 (N_6337,N_1003,N_199);
nor U6338 (N_6338,N_1274,N_480);
nor U6339 (N_6339,N_2186,N_4777);
or U6340 (N_6340,N_2080,N_500);
xnor U6341 (N_6341,N_1434,N_502);
nand U6342 (N_6342,N_2649,N_2674);
or U6343 (N_6343,N_457,N_3660);
xnor U6344 (N_6344,N_2580,N_4383);
nand U6345 (N_6345,N_2430,N_864);
xor U6346 (N_6346,N_873,N_1608);
or U6347 (N_6347,N_4564,N_4000);
nand U6348 (N_6348,N_3721,N_4652);
nor U6349 (N_6349,N_3979,N_2045);
nor U6350 (N_6350,N_2102,N_3919);
and U6351 (N_6351,N_1206,N_1668);
nor U6352 (N_6352,N_4881,N_4213);
nand U6353 (N_6353,N_4772,N_3401);
nor U6354 (N_6354,N_4549,N_3872);
or U6355 (N_6355,N_1984,N_3311);
and U6356 (N_6356,N_1853,N_2949);
nand U6357 (N_6357,N_1868,N_3419);
nand U6358 (N_6358,N_1652,N_3254);
nor U6359 (N_6359,N_2719,N_3984);
and U6360 (N_6360,N_901,N_1366);
nor U6361 (N_6361,N_4423,N_3852);
xnor U6362 (N_6362,N_2621,N_1312);
and U6363 (N_6363,N_751,N_2308);
or U6364 (N_6364,N_1701,N_4558);
nor U6365 (N_6365,N_4076,N_3164);
nor U6366 (N_6366,N_3243,N_3830);
or U6367 (N_6367,N_3770,N_4005);
and U6368 (N_6368,N_1718,N_1542);
nor U6369 (N_6369,N_640,N_2352);
or U6370 (N_6370,N_3667,N_989);
xor U6371 (N_6371,N_2725,N_808);
nor U6372 (N_6372,N_1162,N_3442);
nand U6373 (N_6373,N_4307,N_3138);
and U6374 (N_6374,N_2851,N_3844);
and U6375 (N_6375,N_2522,N_3707);
or U6376 (N_6376,N_3261,N_2765);
nor U6377 (N_6377,N_4811,N_2952);
xnor U6378 (N_6378,N_4196,N_396);
xor U6379 (N_6379,N_3172,N_2543);
xnor U6380 (N_6380,N_1457,N_3431);
nor U6381 (N_6381,N_1794,N_313);
and U6382 (N_6382,N_4522,N_1038);
or U6383 (N_6383,N_1743,N_4944);
nand U6384 (N_6384,N_1921,N_4865);
nor U6385 (N_6385,N_4275,N_4895);
and U6386 (N_6386,N_2925,N_1784);
and U6387 (N_6387,N_180,N_4608);
or U6388 (N_6388,N_2091,N_837);
or U6389 (N_6389,N_3751,N_1746);
xnor U6390 (N_6390,N_3385,N_4425);
or U6391 (N_6391,N_2627,N_2484);
and U6392 (N_6392,N_3578,N_4373);
xor U6393 (N_6393,N_1407,N_220);
xnor U6394 (N_6394,N_1801,N_2488);
xor U6395 (N_6395,N_1979,N_4422);
xor U6396 (N_6396,N_2469,N_1555);
or U6397 (N_6397,N_3819,N_2535);
nor U6398 (N_6398,N_4577,N_3635);
and U6399 (N_6399,N_1443,N_215);
nand U6400 (N_6400,N_4366,N_435);
nand U6401 (N_6401,N_250,N_448);
nor U6402 (N_6402,N_3821,N_2530);
nor U6403 (N_6403,N_3113,N_3931);
nor U6404 (N_6404,N_784,N_2707);
xor U6405 (N_6405,N_2612,N_3898);
and U6406 (N_6406,N_3148,N_525);
and U6407 (N_6407,N_3524,N_2630);
nor U6408 (N_6408,N_2499,N_3598);
and U6409 (N_6409,N_2968,N_4923);
nor U6410 (N_6410,N_1187,N_4532);
nand U6411 (N_6411,N_3552,N_1583);
nand U6412 (N_6412,N_4413,N_4410);
nor U6413 (N_6413,N_4358,N_3165);
nand U6414 (N_6414,N_1925,N_781);
nand U6415 (N_6415,N_2048,N_2780);
and U6416 (N_6416,N_1467,N_3049);
nand U6417 (N_6417,N_1194,N_936);
nor U6418 (N_6418,N_4353,N_1632);
or U6419 (N_6419,N_3516,N_1114);
and U6420 (N_6420,N_4567,N_882);
nand U6421 (N_6421,N_329,N_2131);
and U6422 (N_6422,N_3043,N_1203);
nor U6423 (N_6423,N_2704,N_4693);
and U6424 (N_6424,N_3692,N_4130);
xnor U6425 (N_6425,N_860,N_4273);
nand U6426 (N_6426,N_31,N_1580);
and U6427 (N_6427,N_3881,N_2169);
xnor U6428 (N_6428,N_468,N_4189);
xor U6429 (N_6429,N_1447,N_1432);
xor U6430 (N_6430,N_942,N_3965);
or U6431 (N_6431,N_568,N_1305);
nand U6432 (N_6432,N_1736,N_4871);
nor U6433 (N_6433,N_437,N_3523);
or U6434 (N_6434,N_4347,N_2411);
nand U6435 (N_6435,N_168,N_3312);
nand U6436 (N_6436,N_2517,N_2233);
nand U6437 (N_6437,N_1905,N_1821);
nor U6438 (N_6438,N_3012,N_4021);
nor U6439 (N_6439,N_2246,N_1897);
nand U6440 (N_6440,N_4869,N_431);
or U6441 (N_6441,N_3265,N_625);
nor U6442 (N_6442,N_406,N_3288);
nor U6443 (N_6443,N_967,N_301);
nor U6444 (N_6444,N_195,N_2049);
nand U6445 (N_6445,N_684,N_3518);
xor U6446 (N_6446,N_1710,N_1864);
nand U6447 (N_6447,N_4083,N_4498);
xnor U6448 (N_6448,N_3973,N_4332);
nand U6449 (N_6449,N_101,N_557);
and U6450 (N_6450,N_2908,N_2073);
or U6451 (N_6451,N_4148,N_284);
or U6452 (N_6452,N_4289,N_3892);
xnor U6453 (N_6453,N_4073,N_4317);
nor U6454 (N_6454,N_1832,N_2750);
and U6455 (N_6455,N_2830,N_4334);
nor U6456 (N_6456,N_3457,N_3152);
and U6457 (N_6457,N_1411,N_4551);
or U6458 (N_6458,N_890,N_2158);
and U6459 (N_6459,N_201,N_4238);
nand U6460 (N_6460,N_2020,N_385);
and U6461 (N_6461,N_2214,N_2205);
or U6462 (N_6462,N_919,N_4710);
nor U6463 (N_6463,N_69,N_411);
xor U6464 (N_6464,N_3258,N_608);
and U6465 (N_6465,N_3270,N_340);
or U6466 (N_6466,N_843,N_4031);
nor U6467 (N_6467,N_2427,N_3449);
nor U6468 (N_6468,N_2540,N_630);
nor U6469 (N_6469,N_4945,N_4978);
xor U6470 (N_6470,N_433,N_3383);
xnor U6471 (N_6471,N_381,N_1963);
and U6472 (N_6472,N_1932,N_3937);
nor U6473 (N_6473,N_3432,N_483);
nor U6474 (N_6474,N_3551,N_2910);
and U6475 (N_6475,N_3381,N_117);
and U6476 (N_6476,N_2311,N_1807);
and U6477 (N_6477,N_1164,N_2986);
or U6478 (N_6478,N_811,N_2574);
and U6479 (N_6479,N_2210,N_4173);
and U6480 (N_6480,N_1956,N_430);
and U6481 (N_6481,N_1070,N_446);
or U6482 (N_6482,N_2170,N_3920);
nor U6483 (N_6483,N_4380,N_3139);
or U6484 (N_6484,N_554,N_2773);
or U6485 (N_6485,N_505,N_3964);
xnor U6486 (N_6486,N_2716,N_3022);
nand U6487 (N_6487,N_308,N_2003);
and U6488 (N_6488,N_2063,N_3068);
nand U6489 (N_6489,N_506,N_3680);
or U6490 (N_6490,N_1735,N_4374);
nand U6491 (N_6491,N_1670,N_4481);
xor U6492 (N_6492,N_2994,N_2107);
or U6493 (N_6493,N_1370,N_545);
xor U6494 (N_6494,N_2620,N_1134);
and U6495 (N_6495,N_4699,N_511);
and U6496 (N_6496,N_1072,N_2014);
and U6497 (N_6497,N_443,N_1438);
and U6498 (N_6498,N_1441,N_1881);
nor U6499 (N_6499,N_1149,N_1958);
and U6500 (N_6500,N_1245,N_3665);
xnor U6501 (N_6501,N_2711,N_2742);
nand U6502 (N_6502,N_2262,N_1913);
or U6503 (N_6503,N_1151,N_2737);
xnor U6504 (N_6504,N_2870,N_2353);
xor U6505 (N_6505,N_4089,N_2021);
or U6506 (N_6506,N_2410,N_1562);
xor U6507 (N_6507,N_1034,N_3483);
nor U6508 (N_6508,N_3123,N_2000);
or U6509 (N_6509,N_871,N_3330);
nand U6510 (N_6510,N_1855,N_1449);
nand U6511 (N_6511,N_1078,N_4493);
nand U6512 (N_6512,N_3194,N_3570);
nand U6513 (N_6513,N_1439,N_3639);
xor U6514 (N_6514,N_3136,N_2956);
and U6515 (N_6515,N_3023,N_61);
nand U6516 (N_6516,N_4982,N_70);
nand U6517 (N_6517,N_2920,N_2140);
or U6518 (N_6518,N_4607,N_4016);
nor U6519 (N_6519,N_4163,N_800);
nor U6520 (N_6520,N_4407,N_2061);
nand U6521 (N_6521,N_4921,N_1405);
or U6522 (N_6522,N_4451,N_3335);
xor U6523 (N_6523,N_4298,N_295);
and U6524 (N_6524,N_875,N_805);
xor U6525 (N_6525,N_3360,N_4554);
xnor U6526 (N_6526,N_1692,N_2179);
nor U6527 (N_6527,N_2857,N_965);
nand U6528 (N_6528,N_127,N_4601);
nand U6529 (N_6529,N_78,N_4153);
and U6530 (N_6530,N_3768,N_2393);
and U6531 (N_6531,N_1087,N_1338);
nand U6532 (N_6532,N_4792,N_3702);
or U6533 (N_6533,N_2181,N_4051);
xor U6534 (N_6534,N_3413,N_4253);
xnor U6535 (N_6535,N_934,N_331);
and U6536 (N_6536,N_3924,N_2790);
or U6537 (N_6537,N_662,N_3155);
xnor U6538 (N_6538,N_832,N_1208);
xnor U6539 (N_6539,N_3602,N_900);
nor U6540 (N_6540,N_2042,N_3440);
xnor U6541 (N_6541,N_3633,N_3297);
nand U6542 (N_6542,N_957,N_156);
nand U6543 (N_6543,N_4629,N_3430);
xnor U6544 (N_6544,N_3103,N_4934);
or U6545 (N_6545,N_3214,N_638);
nand U6546 (N_6546,N_1365,N_4424);
and U6547 (N_6547,N_1448,N_4818);
nand U6548 (N_6548,N_2220,N_1532);
xor U6549 (N_6549,N_2101,N_2813);
nand U6550 (N_6550,N_2243,N_2981);
xor U6551 (N_6551,N_4899,N_2273);
nand U6552 (N_6552,N_1354,N_2461);
or U6553 (N_6553,N_84,N_4223);
or U6554 (N_6554,N_4858,N_1244);
xor U6555 (N_6555,N_1955,N_128);
xnor U6556 (N_6556,N_1180,N_4483);
or U6557 (N_6557,N_626,N_4209);
nand U6558 (N_6558,N_956,N_213);
nor U6559 (N_6559,N_3611,N_3414);
nand U6560 (N_6560,N_3126,N_4296);
or U6561 (N_6561,N_1289,N_2373);
and U6562 (N_6562,N_451,N_816);
and U6563 (N_6563,N_3820,N_408);
nand U6564 (N_6564,N_4052,N_4531);
nor U6565 (N_6565,N_603,N_852);
nand U6566 (N_6566,N_132,N_2533);
nand U6567 (N_6567,N_4091,N_3719);
xnor U6568 (N_6568,N_2297,N_3498);
xor U6569 (N_6569,N_1584,N_2122);
xor U6570 (N_6570,N_1002,N_865);
and U6571 (N_6571,N_921,N_4600);
nand U6572 (N_6572,N_2109,N_3650);
xor U6573 (N_6573,N_4125,N_4887);
nand U6574 (N_6574,N_2654,N_4308);
or U6575 (N_6575,N_1502,N_2735);
nor U6576 (N_6576,N_3291,N_2344);
and U6577 (N_6577,N_4536,N_744);
or U6578 (N_6578,N_598,N_2320);
and U6579 (N_6579,N_2094,N_1536);
nor U6580 (N_6580,N_4181,N_1903);
xor U6581 (N_6581,N_4379,N_4499);
nor U6582 (N_6582,N_1774,N_813);
and U6583 (N_6583,N_2520,N_2579);
nand U6584 (N_6584,N_3319,N_4431);
xor U6585 (N_6585,N_4007,N_859);
and U6586 (N_6586,N_3799,N_3465);
or U6587 (N_6587,N_3690,N_3014);
nand U6588 (N_6588,N_3403,N_1561);
xnor U6589 (N_6589,N_325,N_1620);
and U6590 (N_6590,N_4534,N_1524);
nor U6591 (N_6591,N_2635,N_1131);
nor U6592 (N_6592,N_1137,N_4386);
or U6593 (N_6593,N_1133,N_1473);
and U6594 (N_6594,N_981,N_514);
or U6595 (N_6595,N_3777,N_861);
nand U6596 (N_6596,N_2673,N_1978);
nand U6597 (N_6597,N_455,N_1243);
and U6598 (N_6598,N_2820,N_4119);
xor U6599 (N_6599,N_4779,N_4886);
nor U6600 (N_6600,N_3088,N_4992);
and U6601 (N_6601,N_2089,N_4348);
and U6602 (N_6602,N_4055,N_4199);
and U6603 (N_6603,N_4768,N_1242);
or U6604 (N_6604,N_4428,N_2940);
xor U6605 (N_6605,N_4589,N_1417);
nand U6606 (N_6606,N_335,N_4916);
nand U6607 (N_6607,N_2754,N_332);
or U6608 (N_6608,N_1806,N_1751);
nand U6609 (N_6609,N_888,N_4618);
nand U6610 (N_6610,N_652,N_2010);
nor U6611 (N_6611,N_2165,N_3106);
xnor U6612 (N_6612,N_3446,N_4412);
and U6613 (N_6613,N_1117,N_37);
xor U6614 (N_6614,N_4024,N_1469);
or U6615 (N_6615,N_3527,N_661);
or U6616 (N_6616,N_1930,N_3064);
and U6617 (N_6617,N_1515,N_4718);
and U6618 (N_6618,N_2250,N_4889);
or U6619 (N_6619,N_2785,N_315);
nor U6620 (N_6620,N_4020,N_1053);
and U6621 (N_6621,N_1721,N_2239);
or U6622 (N_6622,N_1246,N_4862);
and U6623 (N_6623,N_1079,N_2190);
xnor U6624 (N_6624,N_3514,N_1644);
xnor U6625 (N_6625,N_3814,N_1669);
and U6626 (N_6626,N_265,N_2212);
and U6627 (N_6627,N_2817,N_269);
xor U6628 (N_6628,N_2050,N_317);
nor U6629 (N_6629,N_1626,N_2357);
nand U6630 (N_6630,N_2906,N_2019);
nor U6631 (N_6631,N_2603,N_4771);
or U6632 (N_6632,N_4381,N_1842);
nor U6633 (N_6633,N_2592,N_1773);
xor U6634 (N_6634,N_172,N_4832);
nand U6635 (N_6635,N_903,N_1176);
nor U6636 (N_6636,N_4999,N_4625);
xnor U6637 (N_6637,N_595,N_3359);
xor U6638 (N_6638,N_2577,N_980);
nand U6639 (N_6639,N_2381,N_422);
nand U6640 (N_6640,N_3978,N_2774);
xnor U6641 (N_6641,N_3142,N_304);
nor U6642 (N_6642,N_472,N_1959);
xor U6643 (N_6643,N_4184,N_1348);
or U6644 (N_6644,N_3672,N_2897);
nand U6645 (N_6645,N_2891,N_374);
and U6646 (N_6646,N_2547,N_3669);
and U6647 (N_6647,N_4850,N_1770);
or U6648 (N_6648,N_3266,N_3874);
or U6649 (N_6649,N_2383,N_3097);
nand U6650 (N_6650,N_4961,N_985);
or U6651 (N_6651,N_969,N_2121);
and U6652 (N_6652,N_4676,N_4613);
or U6653 (N_6653,N_3785,N_1413);
nand U6654 (N_6654,N_2714,N_1080);
xor U6655 (N_6655,N_4518,N_4606);
nor U6656 (N_6656,N_1403,N_3913);
and U6657 (N_6657,N_2288,N_2606);
nor U6658 (N_6658,N_1496,N_3407);
or U6659 (N_6659,N_67,N_3228);
or U6660 (N_6660,N_2650,N_3306);
nor U6661 (N_6661,N_1369,N_4368);
and U6662 (N_6662,N_302,N_747);
and U6663 (N_6663,N_4994,N_4299);
or U6664 (N_6664,N_1762,N_1519);
xor U6665 (N_6665,N_2051,N_3052);
nand U6666 (N_6666,N_1306,N_4162);
nand U6667 (N_6667,N_4503,N_1582);
or U6668 (N_6668,N_3778,N_11);
and U6669 (N_6669,N_4027,N_2305);
nor U6670 (N_6670,N_3056,N_4050);
nor U6671 (N_6671,N_574,N_2309);
or U6672 (N_6672,N_2485,N_916);
and U6673 (N_6673,N_3190,N_2934);
nor U6674 (N_6674,N_1712,N_1027);
xnor U6675 (N_6675,N_3756,N_3382);
xor U6676 (N_6676,N_3127,N_932);
xor U6677 (N_6677,N_50,N_1594);
xnor U6678 (N_6678,N_3084,N_2831);
xor U6679 (N_6679,N_927,N_3276);
or U6680 (N_6680,N_3444,N_1535);
or U6681 (N_6681,N_3708,N_2809);
or U6682 (N_6682,N_1733,N_197);
nor U6683 (N_6683,N_4648,N_2361);
and U6684 (N_6684,N_2242,N_130);
and U6685 (N_6685,N_3239,N_1673);
or U6686 (N_6686,N_72,N_3428);
and U6687 (N_6687,N_1898,N_338);
xnor U6688 (N_6688,N_3505,N_1296);
and U6689 (N_6689,N_1749,N_3930);
xnor U6690 (N_6690,N_4454,N_3083);
or U6691 (N_6691,N_3232,N_4970);
nand U6692 (N_6692,N_1780,N_3379);
or U6693 (N_6693,N_4541,N_1019);
or U6694 (N_6694,N_3394,N_2175);
xor U6695 (N_6695,N_1717,N_4511);
xnor U6696 (N_6696,N_2152,N_1573);
xnor U6697 (N_6697,N_32,N_1476);
or U6698 (N_6698,N_261,N_4833);
or U6699 (N_6699,N_4778,N_2099);
xnor U6700 (N_6700,N_3151,N_922);
nand U6701 (N_6701,N_3212,N_27);
nor U6702 (N_6702,N_2197,N_1358);
nor U6703 (N_6703,N_4813,N_1456);
and U6704 (N_6704,N_745,N_2360);
xor U6705 (N_6705,N_1311,N_399);
xor U6706 (N_6706,N_310,N_1646);
and U6707 (N_6707,N_3638,N_2401);
nand U6708 (N_6708,N_4336,N_770);
xnor U6709 (N_6709,N_2420,N_3565);
or U6710 (N_6710,N_2950,N_404);
and U6711 (N_6711,N_834,N_3251);
or U6712 (N_6712,N_1339,N_520);
xnor U6713 (N_6713,N_1589,N_4742);
and U6714 (N_6714,N_2663,N_2159);
nand U6715 (N_6715,N_1388,N_3599);
or U6716 (N_6716,N_4565,N_3546);
xor U6717 (N_6717,N_1686,N_3713);
nand U6718 (N_6718,N_2876,N_89);
or U6719 (N_6719,N_1940,N_454);
nand U6720 (N_6720,N_4327,N_1430);
or U6721 (N_6721,N_3648,N_281);
nor U6722 (N_6722,N_232,N_3581);
nand U6723 (N_6723,N_2415,N_4653);
nand U6724 (N_6724,N_4525,N_1036);
xor U6725 (N_6725,N_1168,N_3217);
nor U6726 (N_6726,N_541,N_674);
or U6727 (N_6727,N_1858,N_4514);
xor U6728 (N_6728,N_2961,N_2103);
xor U6729 (N_6729,N_556,N_2389);
nand U6730 (N_6730,N_952,N_4979);
and U6731 (N_6731,N_3960,N_2634);
nor U6732 (N_6732,N_3559,N_2976);
xnor U6733 (N_6733,N_2806,N_1761);
xor U6734 (N_6734,N_2277,N_2945);
nand U6735 (N_6735,N_2775,N_1768);
or U6736 (N_6736,N_2509,N_2743);
or U6737 (N_6737,N_2434,N_1994);
and U6738 (N_6738,N_134,N_1658);
xor U6739 (N_6739,N_3521,N_4974);
nand U6740 (N_6740,N_1871,N_2269);
nand U6741 (N_6741,N_3848,N_4880);
xnor U6742 (N_6742,N_1530,N_3008);
and U6743 (N_6743,N_906,N_1043);
xnor U6744 (N_6744,N_2219,N_1130);
nand U6745 (N_6745,N_343,N_3583);
xnor U6746 (N_6746,N_2024,N_2899);
and U6747 (N_6747,N_1674,N_2095);
nor U6748 (N_6748,N_2384,N_740);
xor U6749 (N_6749,N_4773,N_2808);
nand U6750 (N_6750,N_3173,N_1527);
and U6751 (N_6751,N_4767,N_2267);
or U6752 (N_6752,N_493,N_609);
xnor U6753 (N_6753,N_2163,N_1885);
xor U6754 (N_6754,N_1791,N_2688);
or U6755 (N_6755,N_95,N_2460);
nand U6756 (N_6756,N_60,N_3762);
nand U6757 (N_6757,N_2379,N_978);
xor U6758 (N_6758,N_2724,N_383);
xor U6759 (N_6759,N_252,N_4933);
or U6760 (N_6760,N_2017,N_3329);
nor U6761 (N_6761,N_2844,N_19);
xnor U6762 (N_6762,N_3169,N_4995);
nor U6763 (N_6763,N_4344,N_3837);
nand U6764 (N_6764,N_150,N_4729);
and U6765 (N_6765,N_4365,N_4449);
nand U6766 (N_6766,N_45,N_410);
nor U6767 (N_6767,N_3698,N_1318);
or U6768 (N_6768,N_2435,N_3479);
nor U6769 (N_6769,N_4651,N_1281);
or U6770 (N_6770,N_3380,N_4105);
xor U6771 (N_6771,N_2607,N_2880);
and U6772 (N_6772,N_4448,N_3496);
or U6773 (N_6773,N_3911,N_2164);
xor U6774 (N_6774,N_1526,N_2238);
nor U6775 (N_6775,N_242,N_2135);
nor U6776 (N_6776,N_4654,N_3914);
nand U6777 (N_6777,N_1215,N_2858);
xnor U6778 (N_6778,N_3021,N_671);
or U6779 (N_6779,N_869,N_1779);
or U6780 (N_6780,N_2521,N_2149);
nand U6781 (N_6781,N_4147,N_3969);
nand U6782 (N_6782,N_3464,N_2669);
nand U6783 (N_6783,N_1204,N_3886);
and U6784 (N_6784,N_3115,N_346);
and U6785 (N_6785,N_1200,N_3908);
nor U6786 (N_6786,N_2907,N_1033);
and U6787 (N_6787,N_3141,N_2390);
nand U6788 (N_6788,N_4924,N_2862);
nand U6789 (N_6789,N_2322,N_4293);
or U6790 (N_6790,N_1316,N_1461);
nand U6791 (N_6791,N_1968,N_4825);
nor U6792 (N_6792,N_4325,N_636);
xnor U6793 (N_6793,N_4343,N_380);
nand U6794 (N_6794,N_2553,N_1577);
or U6795 (N_6795,N_2229,N_3134);
xor U6796 (N_6796,N_2718,N_2879);
and U6797 (N_6797,N_1704,N_4306);
nor U6798 (N_6798,N_401,N_2926);
or U6799 (N_6799,N_3355,N_1708);
xnor U6800 (N_6800,N_3740,N_3610);
xor U6801 (N_6801,N_3593,N_66);
nand U6802 (N_6802,N_2319,N_3854);
nor U6803 (N_6803,N_4167,N_1545);
or U6804 (N_6804,N_723,N_3369);
and U6805 (N_6805,N_1154,N_1823);
and U6806 (N_6806,N_3460,N_1427);
nor U6807 (N_6807,N_2001,N_4985);
and U6808 (N_6808,N_1661,N_2947);
and U6809 (N_6809,N_3653,N_552);
nand U6810 (N_6810,N_4770,N_3370);
xor U6811 (N_6811,N_2106,N_2633);
and U6812 (N_6812,N_663,N_4037);
nand U6813 (N_6813,N_4745,N_1270);
or U6814 (N_6814,N_4085,N_2702);
xor U6815 (N_6815,N_1676,N_2272);
and U6816 (N_6816,N_1547,N_1483);
nand U6817 (N_6817,N_711,N_3051);
xnor U6818 (N_6818,N_3472,N_926);
and U6819 (N_6819,N_3838,N_1760);
and U6820 (N_6820,N_4025,N_1846);
or U6821 (N_6821,N_9,N_1191);
and U6822 (N_6822,N_3752,N_581);
nor U6823 (N_6823,N_819,N_4894);
or U6824 (N_6824,N_3510,N_188);
nor U6825 (N_6825,N_179,N_2450);
nor U6826 (N_6826,N_2425,N_4674);
nor U6827 (N_6827,N_4288,N_223);
nand U6828 (N_6828,N_3289,N_418);
and U6829 (N_6829,N_2562,N_3364);
and U6830 (N_6830,N_3575,N_2189);
xnor U6831 (N_6831,N_3880,N_2480);
nor U6832 (N_6832,N_2376,N_4828);
xnor U6833 (N_6833,N_4019,N_2518);
nor U6834 (N_6834,N_4490,N_4096);
and U6835 (N_6835,N_2194,N_737);
or U6836 (N_6836,N_1946,N_3016);
xnor U6837 (N_6837,N_3996,N_3149);
xnor U6838 (N_6838,N_794,N_2076);
xnor U6839 (N_6839,N_4234,N_1295);
xor U6840 (N_6840,N_4404,N_3180);
and U6841 (N_6841,N_3321,N_2110);
xor U6842 (N_6842,N_405,N_3759);
or U6843 (N_6843,N_2955,N_4621);
xor U6844 (N_6844,N_2697,N_112);
nand U6845 (N_6845,N_1647,N_370);
nand U6846 (N_6846,N_1763,N_4390);
and U6847 (N_6847,N_2667,N_4129);
nand U6848 (N_6848,N_1889,N_3253);
or U6849 (N_6849,N_547,N_3158);
and U6850 (N_6850,N_1995,N_1207);
or U6851 (N_6851,N_717,N_222);
nor U6852 (N_6852,N_3912,N_492);
nand U6853 (N_6853,N_3283,N_2918);
nand U6854 (N_6854,N_4376,N_2291);
nand U6855 (N_6855,N_4845,N_345);
xor U6856 (N_6856,N_305,N_2843);
or U6857 (N_6857,N_2240,N_4803);
and U6858 (N_6858,N_3346,N_643);
nor U6859 (N_6859,N_2292,N_4937);
and U6860 (N_6860,N_597,N_460);
or U6861 (N_6861,N_474,N_4706);
nand U6862 (N_6862,N_2490,N_775);
xor U6863 (N_6863,N_756,N_3737);
and U6864 (N_6864,N_1567,N_1383);
and U6865 (N_6865,N_1225,N_1854);
xnor U6866 (N_6866,N_2282,N_1623);
nor U6867 (N_6867,N_3389,N_3793);
nor U6868 (N_6868,N_570,N_1415);
or U6869 (N_6869,N_314,N_4372);
nand U6870 (N_6870,N_953,N_2928);
or U6871 (N_6871,N_973,N_680);
xor U6872 (N_6872,N_4465,N_2452);
or U6873 (N_6873,N_1278,N_137);
and U6874 (N_6874,N_821,N_937);
and U6875 (N_6875,N_2936,N_3011);
nand U6876 (N_6876,N_123,N_4469);
nor U6877 (N_6877,N_3079,N_1830);
nand U6878 (N_6878,N_4550,N_3030);
and U6879 (N_6879,N_787,N_2066);
or U6880 (N_6880,N_3393,N_4495);
and U6881 (N_6881,N_279,N_2248);
and U6882 (N_6882,N_3710,N_3197);
or U6883 (N_6883,N_2251,N_2431);
or U6884 (N_6884,N_4356,N_3794);
nor U6885 (N_6885,N_4795,N_499);
nor U6886 (N_6886,N_3027,N_3687);
or U6887 (N_6887,N_1706,N_3200);
and U6888 (N_6888,N_3926,N_704);
and U6889 (N_6889,N_607,N_1867);
nor U6890 (N_6890,N_4211,N_3515);
xor U6891 (N_6891,N_3941,N_1213);
nand U6892 (N_6892,N_4405,N_391);
and U6893 (N_6893,N_2470,N_2847);
and U6894 (N_6894,N_192,N_2796);
xnor U6895 (N_6895,N_962,N_2062);
or U6896 (N_6896,N_3917,N_3674);
nand U6897 (N_6897,N_4539,N_3963);
or U6898 (N_6898,N_4943,N_1218);
xnor U6899 (N_6899,N_4427,N_3530);
and U6900 (N_6900,N_4447,N_2059);
or U6901 (N_6901,N_2400,N_2865);
nor U6902 (N_6902,N_3636,N_4562);
nor U6903 (N_6903,N_2593,N_3828);
xor U6904 (N_6904,N_1303,N_2854);
or U6905 (N_6905,N_1325,N_1121);
and U6906 (N_6906,N_434,N_4172);
or U6907 (N_6907,N_392,N_1074);
nor U6908 (N_6908,N_3409,N_2417);
nor U6909 (N_6909,N_1738,N_1471);
and U6910 (N_6910,N_1967,N_2247);
or U6911 (N_6911,N_3220,N_1160);
nand U6912 (N_6912,N_3849,N_1926);
and U6913 (N_6913,N_3988,N_1035);
or U6914 (N_6914,N_110,N_1951);
xor U6915 (N_6915,N_3305,N_3250);
nand U6916 (N_6916,N_1190,N_1531);
xor U6917 (N_6917,N_4500,N_1694);
and U6918 (N_6918,N_3274,N_3709);
and U6919 (N_6919,N_336,N_1214);
and U6920 (N_6920,N_16,N_190);
or U6921 (N_6921,N_3853,N_2873);
and U6922 (N_6922,N_3069,N_4965);
nor U6923 (N_6923,N_1896,N_2005);
nor U6924 (N_6924,N_2954,N_4582);
or U6925 (N_6925,N_918,N_97);
nor U6926 (N_6926,N_3208,N_1409);
xor U6927 (N_6927,N_4747,N_4232);
nor U6928 (N_6928,N_3627,N_1790);
and U6929 (N_6929,N_4598,N_4486);
or U6930 (N_6930,N_2659,N_3656);
xnor U6931 (N_6931,N_3040,N_1379);
or U6932 (N_6932,N_1492,N_3673);
and U6933 (N_6933,N_2887,N_1275);
xnor U6934 (N_6934,N_4839,N_3938);
nor U6935 (N_6935,N_616,N_2329);
nand U6936 (N_6936,N_87,N_2041);
or U6937 (N_6937,N_1216,N_1814);
or U6938 (N_6938,N_1173,N_2075);
nor U6939 (N_6939,N_4494,N_3104);
nand U6940 (N_6940,N_3972,N_3772);
nand U6941 (N_6941,N_987,N_2147);
or U6942 (N_6942,N_264,N_4215);
and U6943 (N_6943,N_2992,N_659);
and U6944 (N_6944,N_2226,N_2275);
and U6945 (N_6945,N_3318,N_1677);
xnor U6946 (N_6946,N_4028,N_1283);
nor U6947 (N_6947,N_277,N_1468);
xor U6948 (N_6948,N_1228,N_76);
and U6949 (N_6949,N_677,N_1226);
xnor U6950 (N_6950,N_2065,N_3620);
xnor U6951 (N_6951,N_3427,N_1631);
nor U6952 (N_6952,N_3795,N_1175);
nor U6953 (N_6953,N_4145,N_3041);
nand U6954 (N_6954,N_639,N_2866);
nand U6955 (N_6955,N_1271,N_4118);
xnor U6956 (N_6956,N_2529,N_4369);
nand U6957 (N_6957,N_3176,N_1742);
nand U6958 (N_6958,N_173,N_3600);
nor U6959 (N_6959,N_2786,N_185);
nand U6960 (N_6960,N_3307,N_1722);
xnor U6961 (N_6961,N_4700,N_1141);
xor U6962 (N_6962,N_3647,N_3668);
xor U6963 (N_6963,N_2418,N_3776);
and U6964 (N_6964,N_2331,N_2171);
xnor U6965 (N_6965,N_1015,N_1753);
or U6966 (N_6966,N_3843,N_2815);
nor U6967 (N_6967,N_2351,N_2286);
and U6968 (N_6968,N_2035,N_3377);
and U6969 (N_6969,N_1299,N_4048);
and U6970 (N_6970,N_1181,N_3734);
and U6971 (N_6971,N_4036,N_2656);
or U6972 (N_6972,N_660,N_4508);
nand U6973 (N_6973,N_2500,N_4905);
xor U6974 (N_6974,N_356,N_4837);
or U6975 (N_6975,N_3238,N_3922);
and U6976 (N_6976,N_2720,N_1609);
and U6977 (N_6977,N_1041,N_3681);
and U6978 (N_6978,N_4457,N_2015);
nor U6979 (N_6979,N_4461,N_1314);
and U6980 (N_6980,N_1998,N_1610);
xnor U6981 (N_6981,N_695,N_1459);
nand U6982 (N_6982,N_2007,N_1859);
or U6983 (N_6983,N_4720,N_2892);
and U6984 (N_6984,N_1611,N_614);
and U6985 (N_6985,N_3520,N_2944);
nor U6986 (N_6986,N_3469,N_4387);
xor U6987 (N_6987,N_1254,N_2027);
nand U6988 (N_6988,N_2216,N_647);
and U6989 (N_6989,N_1962,N_3832);
or U6990 (N_6990,N_1284,N_2476);
xnor U6991 (N_6991,N_3042,N_1024);
xnor U6992 (N_6992,N_2740,N_4252);
xnor U6993 (N_6993,N_4976,N_2167);
or U6994 (N_6994,N_3640,N_3811);
or U6995 (N_6995,N_4241,N_4045);
or U6996 (N_6996,N_3222,N_2922);
nand U6997 (N_6997,N_4480,N_74);
nand U6998 (N_6998,N_4587,N_3588);
or U6999 (N_6999,N_2549,N_4277);
and U7000 (N_7000,N_207,N_3188);
nand U7001 (N_7001,N_394,N_1882);
or U7002 (N_7002,N_1394,N_463);
nor U7003 (N_7003,N_3500,N_4956);
xnor U7004 (N_7004,N_4161,N_3189);
nor U7005 (N_7005,N_2921,N_4853);
and U7006 (N_7006,N_1025,N_3900);
and U7007 (N_7007,N_147,N_4864);
and U7008 (N_7008,N_3810,N_2856);
nand U7009 (N_7009,N_675,N_3582);
and U7010 (N_7010,N_2318,N_4827);
nand U7011 (N_7011,N_3185,N_895);
xor U7012 (N_7012,N_4799,N_3626);
and U7013 (N_7013,N_4217,N_2192);
nor U7014 (N_7014,N_4264,N_3997);
xnor U7015 (N_7015,N_33,N_104);
xor U7016 (N_7016,N_977,N_497);
nand U7017 (N_7017,N_398,N_3195);
and U7018 (N_7018,N_3545,N_4121);
and U7019 (N_7019,N_1633,N_2736);
nand U7020 (N_7020,N_142,N_2433);
xor U7021 (N_7021,N_1660,N_4573);
nand U7022 (N_7022,N_510,N_22);
nor U7023 (N_7023,N_1639,N_1512);
xnor U7024 (N_7024,N_465,N_3328);
and U7025 (N_7025,N_4537,N_2582);
and U7026 (N_7026,N_3655,N_1269);
or U7027 (N_7027,N_1371,N_3899);
nor U7028 (N_7028,N_2129,N_4476);
nor U7029 (N_7029,N_2584,N_3645);
or U7030 (N_7030,N_2074,N_4156);
nand U7031 (N_7031,N_1478,N_782);
and U7032 (N_7032,N_3983,N_1970);
or U7033 (N_7033,N_105,N_1466);
xnor U7034 (N_7034,N_2904,N_4229);
nor U7035 (N_7035,N_1825,N_1342);
or U7036 (N_7036,N_2143,N_1912);
xor U7037 (N_7037,N_1634,N_2358);
and U7038 (N_7038,N_4908,N_3293);
nor U7039 (N_7039,N_386,N_2513);
nand U7040 (N_7040,N_1212,N_4637);
nand U7041 (N_7041,N_1490,N_4401);
or U7042 (N_7042,N_646,N_2492);
or U7043 (N_7043,N_2086,N_1346);
and U7044 (N_7044,N_4455,N_82);
and U7045 (N_7045,N_1324,N_1217);
nor U7046 (N_7046,N_3260,N_4231);
nor U7047 (N_7047,N_3074,N_1322);
or U7048 (N_7048,N_3323,N_3861);
xnor U7049 (N_7049,N_4797,N_2234);
or U7050 (N_7050,N_4579,N_4046);
xnor U7051 (N_7051,N_2700,N_4014);
xnor U7052 (N_7052,N_1538,N_970);
xor U7053 (N_7053,N_2279,N_4798);
nand U7054 (N_7054,N_1709,N_3939);
nand U7055 (N_7055,N_2855,N_3186);
nand U7056 (N_7056,N_776,N_1728);
or U7057 (N_7057,N_319,N_2336);
xnor U7058 (N_7058,N_1144,N_997);
xnor U7059 (N_7059,N_364,N_3936);
and U7060 (N_7060,N_1650,N_108);
or U7061 (N_7061,N_459,N_1915);
or U7062 (N_7062,N_894,N_2442);
and U7063 (N_7063,N_273,N_98);
nor U7064 (N_7064,N_3143,N_1754);
nor U7065 (N_7065,N_2002,N_2983);
xor U7066 (N_7066,N_4474,N_1051);
or U7067 (N_7067,N_4963,N_925);
or U7068 (N_7068,N_4679,N_4553);
or U7069 (N_7069,N_2409,N_4633);
and U7070 (N_7070,N_1904,N_1747);
xor U7071 (N_7071,N_1892,N_4464);
xnor U7072 (N_7072,N_2253,N_944);
or U7073 (N_7073,N_2105,N_1368);
nor U7074 (N_7074,N_2228,N_4548);
xnor U7075 (N_7075,N_3017,N_3304);
nor U7076 (N_7076,N_632,N_1140);
nand U7077 (N_7077,N_3946,N_4647);
nor U7078 (N_7078,N_206,N_2539);
nand U7079 (N_7079,N_347,N_3632);
nor U7080 (N_7080,N_4294,N_2698);
or U7081 (N_7081,N_820,N_2355);
or U7082 (N_7082,N_4841,N_4987);
nand U7083 (N_7083,N_741,N_1453);
xor U7084 (N_7084,N_4281,N_4656);
nand U7085 (N_7085,N_3608,N_1037);
nand U7086 (N_7086,N_2860,N_2257);
nor U7087 (N_7087,N_467,N_3697);
nor U7088 (N_7088,N_2486,N_810);
xnor U7089 (N_7089,N_2298,N_3418);
nand U7090 (N_7090,N_2798,N_267);
nor U7091 (N_7091,N_945,N_507);
nor U7092 (N_7092,N_1186,N_2696);
or U7093 (N_7093,N_2912,N_487);
xnor U7094 (N_7094,N_715,N_2653);
or U7095 (N_7095,N_3686,N_755);
nand U7096 (N_7096,N_15,N_4418);
nor U7097 (N_7097,N_814,N_224);
nor U7098 (N_7098,N_387,N_771);
or U7099 (N_7099,N_426,N_4870);
nor U7100 (N_7100,N_605,N_2677);
and U7101 (N_7101,N_4665,N_803);
or U7102 (N_7102,N_3935,N_2609);
nand U7103 (N_7103,N_2223,N_3845);
nor U7104 (N_7104,N_4456,N_710);
nor U7105 (N_7105,N_4950,N_4506);
or U7106 (N_7106,N_1833,N_4080);
and U7107 (N_7107,N_672,N_851);
xor U7108 (N_7108,N_1068,N_149);
nor U7109 (N_7109,N_3594,N_4360);
xor U7110 (N_7110,N_513,N_2999);
nand U7111 (N_7111,N_1681,N_299);
nor U7112 (N_7112,N_4663,N_4339);
nand U7113 (N_7113,N_2324,N_2570);
nand U7114 (N_7114,N_1505,N_3163);
xor U7115 (N_7115,N_4224,N_2799);
nand U7116 (N_7116,N_417,N_1987);
and U7117 (N_7117,N_1550,N_1622);
nor U7118 (N_7118,N_1498,N_4941);
or U7119 (N_7119,N_3452,N_1808);
or U7120 (N_7120,N_4878,N_4884);
nor U7121 (N_7121,N_378,N_3928);
nand U7122 (N_7122,N_2144,N_4394);
nor U7123 (N_7123,N_4302,N_1384);
xnor U7124 (N_7124,N_494,N_4128);
and U7125 (N_7125,N_719,N_1931);
and U7126 (N_7126,N_2315,N_1193);
nor U7127 (N_7127,N_3682,N_4695);
nor U7128 (N_7128,N_1063,N_42);
xnor U7129 (N_7129,N_2405,N_4879);
nand U7130 (N_7130,N_1261,N_4433);
nor U7131 (N_7131,N_4475,N_3701);
or U7132 (N_7132,N_4983,N_2753);
nor U7133 (N_7133,N_39,N_1105);
and U7134 (N_7134,N_210,N_1558);
xor U7135 (N_7135,N_3388,N_183);
or U7136 (N_7136,N_586,N_3870);
nor U7137 (N_7137,N_2227,N_4194);
or U7138 (N_7138,N_62,N_1971);
or U7139 (N_7139,N_4230,N_3744);
or U7140 (N_7140,N_235,N_4542);
or U7141 (N_7141,N_4854,N_3980);
nand U7142 (N_7142,N_4087,N_2155);
xor U7143 (N_7143,N_3863,N_4437);
nor U7144 (N_7144,N_229,N_4563);
and U7145 (N_7145,N_1659,N_2438);
and U7146 (N_7146,N_1100,N_2188);
xnor U7147 (N_7147,N_4807,N_140);
xor U7148 (N_7148,N_1973,N_1013);
or U7149 (N_7149,N_1835,N_1937);
xor U7150 (N_7150,N_2493,N_2077);
nand U7151 (N_7151,N_3356,N_17);
or U7152 (N_7152,N_691,N_4907);
and U7153 (N_7153,N_1331,N_3448);
xor U7154 (N_7154,N_1876,N_2532);
nor U7155 (N_7155,N_846,N_4124);
and U7156 (N_7156,N_1257,N_4942);
nand U7157 (N_7157,N_4297,N_2180);
nor U7158 (N_7158,N_2655,N_635);
nor U7159 (N_7159,N_1752,N_2875);
or U7160 (N_7160,N_3478,N_3366);
or U7161 (N_7161,N_2755,N_4117);
nand U7162 (N_7162,N_2123,N_2408);
nand U7163 (N_7163,N_645,N_2646);
and U7164 (N_7164,N_754,N_1587);
nor U7165 (N_7165,N_3231,N_1484);
or U7166 (N_7166,N_3517,N_2295);
and U7167 (N_7167,N_462,N_2883);
and U7168 (N_7168,N_233,N_3353);
and U7169 (N_7169,N_2201,N_749);
and U7170 (N_7170,N_2777,N_1127);
or U7171 (N_7171,N_3574,N_2964);
or U7172 (N_7172,N_3888,N_1401);
xor U7173 (N_7173,N_368,N_2788);
or U7174 (N_7174,N_1541,N_960);
nand U7175 (N_7175,N_1546,N_73);
or U7176 (N_7176,N_4660,N_3324);
nand U7177 (N_7177,N_21,N_280);
and U7178 (N_7178,N_2054,N_4609);
xnor U7179 (N_7179,N_453,N_427);
and U7180 (N_7180,N_898,N_3981);
nor U7181 (N_7181,N_99,N_1729);
xor U7182 (N_7182,N_1820,N_4375);
or U7183 (N_7183,N_4882,N_4788);
nor U7184 (N_7184,N_4572,N_4049);
nor U7185 (N_7185,N_2211,N_1944);
and U7186 (N_7186,N_3334,N_3579);
xnor U7187 (N_7187,N_2198,N_1236);
and U7188 (N_7188,N_3729,N_968);
nand U7189 (N_7189,N_4326,N_3398);
or U7190 (N_7190,N_49,N_2290);
xnor U7191 (N_7191,N_278,N_2176);
nor U7192 (N_7192,N_1224,N_3463);
and U7193 (N_7193,N_555,N_1463);
or U7194 (N_7194,N_3279,N_2804);
nor U7195 (N_7195,N_1264,N_3055);
nand U7196 (N_7196,N_3738,N_1222);
and U7197 (N_7197,N_1108,N_2689);
xnor U7198 (N_7198,N_1822,N_3269);
nand U7199 (N_7199,N_4728,N_4743);
nor U7200 (N_7200,N_1506,N_1084);
and U7201 (N_7201,N_4758,N_4315);
and U7202 (N_7202,N_348,N_1799);
nor U7203 (N_7203,N_2872,N_2637);
and U7204 (N_7204,N_1878,N_4984);
nand U7205 (N_7205,N_2575,N_2729);
nor U7206 (N_7206,N_3187,N_714);
nand U7207 (N_7207,N_64,N_1253);
or U7208 (N_7208,N_3050,N_3833);
xor U7209 (N_7209,N_2927,N_654);
xor U7210 (N_7210,N_4491,N_1486);
nor U7211 (N_7211,N_1621,N_503);
xnor U7212 (N_7212,N_623,N_2723);
nand U7213 (N_7213,N_1364,N_3836);
nand U7214 (N_7214,N_3927,N_2739);
nor U7215 (N_7215,N_3075,N_3439);
nand U7216 (N_7216,N_4321,N_1235);
nand U7217 (N_7217,N_111,N_3019);
xnor U7218 (N_7218,N_4478,N_3789);
and U7219 (N_7219,N_3240,N_174);
and U7220 (N_7220,N_3481,N_4823);
and U7221 (N_7221,N_1592,N_79);
or U7222 (N_7222,N_3529,N_3209);
and U7223 (N_7223,N_355,N_701);
and U7224 (N_7224,N_3661,N_2748);
or U7225 (N_7225,N_4930,N_30);
xnor U7226 (N_7226,N_1065,N_4239);
xnor U7227 (N_7227,N_3742,N_897);
nor U7228 (N_7228,N_2367,N_4782);
and U7229 (N_7229,N_4673,N_3716);
or U7230 (N_7230,N_1549,N_3897);
nand U7231 (N_7231,N_2903,N_809);
or U7232 (N_7232,N_1500,N_2330);
nor U7233 (N_7233,N_3375,N_2254);
nor U7234 (N_7234,N_3685,N_2416);
nand U7235 (N_7235,N_2166,N_4846);
nor U7236 (N_7236,N_1414,N_3876);
nor U7237 (N_7237,N_4168,N_4362);
nor U7238 (N_7238,N_2137,N_594);
and U7239 (N_7239,N_2265,N_1139);
nand U7240 (N_7240,N_2778,N_1551);
nand U7241 (N_7241,N_1572,N_2946);
xor U7242 (N_7242,N_2252,N_1952);
xor U7243 (N_7243,N_3868,N_3488);
nand U7244 (N_7244,N_961,N_1157);
or U7245 (N_7245,N_1153,N_2342);
or U7246 (N_7246,N_807,N_1758);
or U7247 (N_7247,N_829,N_512);
and U7248 (N_7248,N_4538,N_4122);
or U7249 (N_7249,N_4208,N_2717);
or U7250 (N_7250,N_1337,N_1192);
or U7251 (N_7251,N_2388,N_80);
or U7252 (N_7252,N_1811,N_1656);
nor U7253 (N_7253,N_4392,N_2507);
and U7254 (N_7254,N_883,N_4844);
nor U7255 (N_7255,N_4927,N_1734);
nand U7256 (N_7256,N_1029,N_333);
and U7257 (N_7257,N_1797,N_1731);
xor U7258 (N_7258,N_2276,N_2259);
or U7259 (N_7259,N_551,N_1026);
nor U7260 (N_7260,N_1887,N_1630);
xor U7261 (N_7261,N_2629,N_4727);
nor U7262 (N_7262,N_2496,N_4127);
xnor U7263 (N_7263,N_3182,N_3352);
nor U7264 (N_7264,N_2628,N_3947);
nand U7265 (N_7265,N_3827,N_879);
xor U7266 (N_7266,N_3715,N_4102);
nand U7267 (N_7267,N_479,N_991);
and U7268 (N_7268,N_2889,N_1918);
and U7269 (N_7269,N_1030,N_515);
xnor U7270 (N_7270,N_2596,N_330);
xor U7271 (N_7271,N_3333,N_1759);
or U7272 (N_7272,N_3542,N_1914);
and U7273 (N_7273,N_2527,N_2097);
xnor U7274 (N_7274,N_4805,N_3765);
nand U7275 (N_7275,N_1619,N_3299);
nor U7276 (N_7276,N_653,N_1172);
nand U7277 (N_7277,N_40,N_4013);
nor U7278 (N_7278,N_2069,N_1590);
nand U7279 (N_7279,N_1544,N_198);
or U7280 (N_7280,N_1247,N_3218);
nand U7281 (N_7281,N_1230,N_582);
nand U7282 (N_7282,N_1120,N_165);
and U7283 (N_7283,N_1115,N_3226);
or U7284 (N_7284,N_4266,N_2447);
nor U7285 (N_7285,N_3024,N_2280);
or U7286 (N_7286,N_2294,N_3422);
and U7287 (N_7287,N_1124,N_2009);
xnor U7288 (N_7288,N_1845,N_4104);
and U7289 (N_7289,N_4236,N_2479);
xnor U7290 (N_7290,N_707,N_4760);
and U7291 (N_7291,N_2591,N_3566);
nor U7292 (N_7292,N_1321,N_3198);
nand U7293 (N_7293,N_3372,N_3441);
xnor U7294 (N_7294,N_3568,N_1118);
xnor U7295 (N_7295,N_2692,N_3798);
or U7296 (N_7296,N_2023,N_2467);
or U7297 (N_7297,N_3045,N_3808);
or U7298 (N_7298,N_892,N_4666);
xnor U7299 (N_7299,N_974,N_4335);
nand U7300 (N_7300,N_2258,N_4852);
and U7301 (N_7301,N_931,N_2304);
nor U7302 (N_7302,N_1893,N_905);
and U7303 (N_7303,N_979,N_778);
nand U7304 (N_7304,N_4775,N_3666);
nand U7305 (N_7305,N_68,N_2929);
nor U7306 (N_7306,N_29,N_2104);
nor U7307 (N_7307,N_3070,N_4800);
nor U7308 (N_7308,N_1367,N_1142);
nor U7309 (N_7309,N_3792,N_2670);
xor U7310 (N_7310,N_2776,N_2274);
or U7311 (N_7311,N_4643,N_2991);
and U7312 (N_7312,N_2043,N_533);
or U7313 (N_7313,N_3491,N_2473);
and U7314 (N_7314,N_289,N_3606);
nand U7315 (N_7315,N_2370,N_1595);
xor U7316 (N_7316,N_3992,N_4135);
and U7317 (N_7317,N_2055,N_4472);
nor U7318 (N_7318,N_896,N_3987);
xor U7319 (N_7319,N_3286,N_262);
or U7320 (N_7320,N_1399,N_4691);
nand U7321 (N_7321,N_1624,N_1352);
nand U7322 (N_7322,N_1834,N_1844);
and U7323 (N_7323,N_3959,N_323);
or U7324 (N_7324,N_4065,N_3725);
and U7325 (N_7325,N_3471,N_3955);
xor U7326 (N_7326,N_1089,N_1462);
nand U7327 (N_7327,N_4137,N_1929);
xor U7328 (N_7328,N_4836,N_1088);
and U7329 (N_7329,N_2510,N_2838);
and U7330 (N_7330,N_2957,N_2118);
and U7331 (N_7331,N_2682,N_2845);
and U7332 (N_7332,N_2793,N_1602);
nand U7333 (N_7333,N_4759,N_2615);
nand U7334 (N_7334,N_612,N_3614);
and U7335 (N_7335,N_2382,N_2449);
nor U7336 (N_7336,N_3763,N_1775);
and U7337 (N_7337,N_1829,N_1596);
nand U7338 (N_7338,N_3053,N_1521);
nor U7339 (N_7339,N_4610,N_4559);
xor U7340 (N_7340,N_3535,N_4501);
nand U7341 (N_7341,N_1810,N_3420);
and U7342 (N_7342,N_3603,N_237);
nand U7343 (N_7343,N_1178,N_4010);
nor U7344 (N_7344,N_4346,N_2366);
and U7345 (N_7345,N_4300,N_2911);
and U7346 (N_7346,N_1960,N_3671);
or U7347 (N_7347,N_4512,N_4323);
or U7348 (N_7348,N_4694,N_3714);
or U7349 (N_7349,N_1061,N_3784);
nor U7350 (N_7350,N_946,N_592);
xnor U7351 (N_7351,N_4426,N_1132);
and U7352 (N_7352,N_1600,N_1831);
xor U7353 (N_7353,N_2287,N_4900);
or U7354 (N_7354,N_4150,N_4303);
and U7355 (N_7355,N_721,N_2289);
nor U7356 (N_7356,N_3310,N_1883);
nand U7357 (N_7357,N_1586,N_1818);
or U7358 (N_7358,N_4033,N_1277);
nor U7359 (N_7359,N_2414,N_2429);
and U7360 (N_7360,N_2462,N_4219);
xor U7361 (N_7361,N_3634,N_3951);
nand U7362 (N_7362,N_1875,N_732);
nand U7363 (N_7363,N_4257,N_2973);
xor U7364 (N_7364,N_353,N_2323);
nand U7365 (N_7365,N_3487,N_2916);
and U7366 (N_7366,N_4123,N_2133);
nor U7367 (N_7367,N_2661,N_1755);
xor U7368 (N_7368,N_1826,N_3374);
nand U7369 (N_7369,N_4986,N_722);
xor U7370 (N_7370,N_855,N_1093);
nand U7371 (N_7371,N_3781,N_1662);
or U7372 (N_7372,N_4284,N_1508);
nand U7373 (N_7373,N_3128,N_4396);
xnor U7374 (N_7374,N_729,N_309);
nor U7375 (N_7375,N_1895,N_641);
and U7376 (N_7376,N_3940,N_2512);
nor U7377 (N_7377,N_35,N_3962);
and U7378 (N_7378,N_4843,N_2824);
or U7379 (N_7379,N_3378,N_3895);
or U7380 (N_7380,N_3750,N_4981);
xor U7381 (N_7381,N_2623,N_642);
xnor U7382 (N_7382,N_2018,N_3338);
xnor U7383 (N_7383,N_486,N_3894);
xnor U7384 (N_7384,N_3179,N_1983);
xnor U7385 (N_7385,N_753,N_3122);
nor U7386 (N_7386,N_1571,N_827);
xnor U7387 (N_7387,N_4191,N_1046);
nor U7388 (N_7388,N_990,N_3952);
xor U7389 (N_7389,N_958,N_889);
xor U7390 (N_7390,N_464,N_2960);
xor U7391 (N_7391,N_3563,N_3029);
or U7392 (N_7392,N_119,N_2626);
xnor U7393 (N_7393,N_3767,N_2224);
xor U7394 (N_7394,N_120,N_1804);
nand U7395 (N_7395,N_3507,N_1307);
and U7396 (N_7396,N_2888,N_830);
nand U7397 (N_7397,N_3099,N_767);
or U7398 (N_7398,N_3204,N_440);
xor U7399 (N_7399,N_3747,N_1901);
nand U7400 (N_7400,N_447,N_1772);
and U7401 (N_7401,N_4664,N_2894);
nand U7402 (N_7402,N_4040,N_1507);
nor U7403 (N_7403,N_1082,N_2505);
xor U7404 (N_7404,N_2676,N_2586);
and U7405 (N_7405,N_4952,N_432);
nand U7406 (N_7406,N_4235,N_4657);
xor U7407 (N_7407,N_1640,N_25);
nand U7408 (N_7408,N_4594,N_4272);
or U7409 (N_7409,N_877,N_4711);
nor U7410 (N_7410,N_145,N_167);
or U7411 (N_7411,N_419,N_2497);
nor U7412 (N_7412,N_1263,N_2705);
nor U7413 (N_7413,N_3171,N_3560);
nor U7414 (N_7414,N_63,N_2312);
xor U7415 (N_7415,N_3219,N_1866);
xor U7416 (N_7416,N_3207,N_4471);
xnor U7417 (N_7417,N_4967,N_3779);
nand U7418 (N_7418,N_1220,N_907);
and U7419 (N_7419,N_203,N_4187);
or U7420 (N_7420,N_4197,N_523);
xnor U7421 (N_7421,N_3769,N_3101);
nor U7422 (N_7422,N_13,N_58);
xor U7423 (N_7423,N_4417,N_4006);
xor U7424 (N_7424,N_4452,N_3054);
nor U7425 (N_7425,N_2260,N_1863);
nor U7426 (N_7426,N_3405,N_1052);
nor U7427 (N_7427,N_1553,N_4059);
and U7428 (N_7428,N_2436,N_4658);
xnor U7429 (N_7429,N_2996,N_3206);
nand U7430 (N_7430,N_2116,N_1789);
nand U7431 (N_7431,N_1841,N_3467);
nor U7432 (N_7432,N_1890,N_1802);
xor U7433 (N_7433,N_4282,N_3887);
and U7434 (N_7434,N_1344,N_1585);
nand U7435 (N_7435,N_4713,N_4397);
and U7436 (N_7436,N_589,N_3929);
nor U7437 (N_7437,N_1933,N_2012);
nand U7438 (N_7438,N_2794,N_2213);
xor U7439 (N_7439,N_559,N_4250);
nand U7440 (N_7440,N_28,N_2391);
xor U7441 (N_7441,N_4214,N_4340);
xnor U7442 (N_7442,N_2444,N_4591);
or U7443 (N_7443,N_2791,N_3736);
nand U7444 (N_7444,N_4680,N_2978);
or U7445 (N_7445,N_4088,N_2731);
or U7446 (N_7446,N_4885,N_158);
or U7447 (N_7447,N_3577,N_342);
or U7448 (N_7448,N_4056,N_2203);
nand U7449 (N_7449,N_4126,N_3406);
and U7450 (N_7450,N_3235,N_4892);
xor U7451 (N_7451,N_3801,N_3851);
and U7452 (N_7452,N_4395,N_1304);
and U7453 (N_7453,N_2413,N_2708);
and U7454 (N_7454,N_3125,N_1847);
nand U7455 (N_7455,N_382,N_1671);
nand U7456 (N_7456,N_43,N_3201);
nor U7457 (N_7457,N_2882,N_709);
xnor U7458 (N_7458,N_1110,N_2977);
nor U7459 (N_7459,N_3096,N_4416);
xnor U7460 (N_7460,N_2468,N_1256);
nand U7461 (N_7461,N_4328,N_1014);
and U7462 (N_7462,N_2651,N_1392);
or U7463 (N_7463,N_1559,N_959);
and U7464 (N_7464,N_2834,N_4705);
nor U7465 (N_7465,N_288,N_2489);
nand U7466 (N_7466,N_4245,N_4164);
nor U7467 (N_7467,N_2624,N_2071);
xnor U7468 (N_7468,N_3387,N_4906);
nand U7469 (N_7469,N_4683,N_963);
xnor U7470 (N_7470,N_0,N_1350);
or U7471 (N_7471,N_1071,N_124);
nand U7472 (N_7472,N_36,N_1837);
xnor U7473 (N_7473,N_2284,N_4988);
nand U7474 (N_7474,N_4363,N_4739);
nor U7475 (N_7475,N_4586,N_4719);
and U7476 (N_7476,N_349,N_1174);
nor U7477 (N_7477,N_2995,N_3107);
xor U7478 (N_7478,N_2657,N_2552);
nor U7479 (N_7479,N_2271,N_2970);
nand U7480 (N_7480,N_4212,N_4696);
nand U7481 (N_7481,N_3780,N_303);
nand U7482 (N_7482,N_4787,N_1748);
nor U7483 (N_7483,N_4442,N_2975);
nor U7484 (N_7484,N_1891,N_4915);
xnor U7485 (N_7485,N_1614,N_3098);
nand U7486 (N_7486,N_2516,N_311);
or U7487 (N_7487,N_1560,N_2760);
or U7488 (N_7488,N_193,N_2822);
and U7489 (N_7489,N_20,N_3641);
and U7490 (N_7490,N_904,N_481);
and U7491 (N_7491,N_254,N_1135);
or U7492 (N_7492,N_4545,N_4107);
nand U7493 (N_7493,N_2124,N_3221);
and U7494 (N_7494,N_644,N_2154);
nor U7495 (N_7495,N_4504,N_2119);
nor U7496 (N_7496,N_2511,N_676);
nand U7497 (N_7497,N_71,N_1238);
or U7498 (N_7498,N_2816,N_3841);
xor U7499 (N_7499,N_2837,N_3879);
and U7500 (N_7500,N_1107,N_4196);
or U7501 (N_7501,N_1551,N_4189);
nor U7502 (N_7502,N_2002,N_3085);
nor U7503 (N_7503,N_3977,N_154);
nor U7504 (N_7504,N_2794,N_959);
and U7505 (N_7505,N_3404,N_4435);
or U7506 (N_7506,N_824,N_3772);
nand U7507 (N_7507,N_3754,N_4412);
nor U7508 (N_7508,N_4544,N_1253);
nand U7509 (N_7509,N_1734,N_3089);
xor U7510 (N_7510,N_3214,N_1089);
nand U7511 (N_7511,N_54,N_3328);
nand U7512 (N_7512,N_4761,N_1523);
nor U7513 (N_7513,N_2393,N_4591);
xnor U7514 (N_7514,N_1228,N_2658);
xor U7515 (N_7515,N_3423,N_2566);
or U7516 (N_7516,N_2047,N_3465);
nand U7517 (N_7517,N_4448,N_2734);
and U7518 (N_7518,N_2731,N_233);
or U7519 (N_7519,N_3154,N_3050);
nand U7520 (N_7520,N_1185,N_1866);
nor U7521 (N_7521,N_4378,N_4150);
nand U7522 (N_7522,N_458,N_3697);
or U7523 (N_7523,N_4871,N_2017);
nand U7524 (N_7524,N_1814,N_4140);
and U7525 (N_7525,N_4637,N_1018);
and U7526 (N_7526,N_814,N_2767);
or U7527 (N_7527,N_370,N_2328);
and U7528 (N_7528,N_1327,N_3670);
xnor U7529 (N_7529,N_4913,N_4393);
or U7530 (N_7530,N_1427,N_3637);
xor U7531 (N_7531,N_270,N_1886);
nor U7532 (N_7532,N_1564,N_76);
xor U7533 (N_7533,N_3735,N_4138);
or U7534 (N_7534,N_4565,N_4018);
nor U7535 (N_7535,N_2015,N_3047);
xor U7536 (N_7536,N_3496,N_1246);
xor U7537 (N_7537,N_57,N_2917);
nor U7538 (N_7538,N_1661,N_1423);
or U7539 (N_7539,N_1704,N_1466);
nand U7540 (N_7540,N_4369,N_4631);
or U7541 (N_7541,N_821,N_1462);
and U7542 (N_7542,N_200,N_1561);
nand U7543 (N_7543,N_471,N_2282);
nand U7544 (N_7544,N_3552,N_3703);
or U7545 (N_7545,N_2827,N_1080);
and U7546 (N_7546,N_2457,N_4094);
nand U7547 (N_7547,N_4133,N_4933);
nor U7548 (N_7548,N_4060,N_4866);
xor U7549 (N_7549,N_3066,N_556);
xnor U7550 (N_7550,N_748,N_1323);
nor U7551 (N_7551,N_4733,N_3417);
xor U7552 (N_7552,N_2252,N_1284);
nor U7553 (N_7553,N_2206,N_4816);
and U7554 (N_7554,N_4573,N_2318);
and U7555 (N_7555,N_1515,N_3996);
or U7556 (N_7556,N_1436,N_4127);
and U7557 (N_7557,N_3802,N_1116);
xnor U7558 (N_7558,N_3396,N_2090);
and U7559 (N_7559,N_3600,N_4617);
and U7560 (N_7560,N_2335,N_940);
and U7561 (N_7561,N_1081,N_4098);
nor U7562 (N_7562,N_324,N_1355);
xor U7563 (N_7563,N_1712,N_2706);
xor U7564 (N_7564,N_794,N_983);
xnor U7565 (N_7565,N_3096,N_1357);
nor U7566 (N_7566,N_2927,N_4516);
nand U7567 (N_7567,N_4318,N_1430);
xor U7568 (N_7568,N_4873,N_1352);
and U7569 (N_7569,N_2455,N_889);
nand U7570 (N_7570,N_4006,N_253);
xor U7571 (N_7571,N_1991,N_400);
and U7572 (N_7572,N_2354,N_3149);
or U7573 (N_7573,N_198,N_3072);
nand U7574 (N_7574,N_3822,N_1003);
or U7575 (N_7575,N_3844,N_4522);
xnor U7576 (N_7576,N_2489,N_2862);
nor U7577 (N_7577,N_4122,N_3021);
or U7578 (N_7578,N_1002,N_1610);
nand U7579 (N_7579,N_4869,N_2588);
xnor U7580 (N_7580,N_3825,N_2086);
nor U7581 (N_7581,N_3657,N_354);
and U7582 (N_7582,N_2385,N_4012);
nand U7583 (N_7583,N_381,N_3314);
nand U7584 (N_7584,N_1097,N_2456);
or U7585 (N_7585,N_2304,N_4288);
nor U7586 (N_7586,N_4159,N_3442);
nand U7587 (N_7587,N_1651,N_939);
and U7588 (N_7588,N_44,N_4800);
xor U7589 (N_7589,N_2754,N_382);
xor U7590 (N_7590,N_2585,N_3452);
xor U7591 (N_7591,N_3504,N_4684);
nor U7592 (N_7592,N_2909,N_4183);
nor U7593 (N_7593,N_3439,N_3378);
and U7594 (N_7594,N_3927,N_4915);
nor U7595 (N_7595,N_2290,N_3163);
nor U7596 (N_7596,N_712,N_1326);
and U7597 (N_7597,N_1615,N_3004);
nor U7598 (N_7598,N_430,N_3525);
xnor U7599 (N_7599,N_1530,N_1415);
xor U7600 (N_7600,N_3884,N_295);
nand U7601 (N_7601,N_468,N_1771);
and U7602 (N_7602,N_3086,N_2454);
and U7603 (N_7603,N_3749,N_4487);
and U7604 (N_7604,N_1760,N_1736);
xor U7605 (N_7605,N_4957,N_1395);
nand U7606 (N_7606,N_2856,N_4168);
nor U7607 (N_7607,N_3991,N_2829);
or U7608 (N_7608,N_2546,N_1227);
and U7609 (N_7609,N_2603,N_513);
nor U7610 (N_7610,N_1132,N_1346);
and U7611 (N_7611,N_4069,N_3155);
or U7612 (N_7612,N_2633,N_4928);
nand U7613 (N_7613,N_3908,N_4214);
xnor U7614 (N_7614,N_933,N_3957);
and U7615 (N_7615,N_381,N_524);
or U7616 (N_7616,N_2679,N_123);
and U7617 (N_7617,N_3320,N_2640);
nor U7618 (N_7618,N_2689,N_2579);
nor U7619 (N_7619,N_2219,N_3910);
nor U7620 (N_7620,N_4682,N_1546);
and U7621 (N_7621,N_3980,N_4878);
nor U7622 (N_7622,N_750,N_1877);
nand U7623 (N_7623,N_3157,N_4118);
or U7624 (N_7624,N_4476,N_3119);
or U7625 (N_7625,N_4377,N_1549);
xnor U7626 (N_7626,N_609,N_4607);
xnor U7627 (N_7627,N_1799,N_2759);
nand U7628 (N_7628,N_2314,N_742);
and U7629 (N_7629,N_2887,N_2936);
and U7630 (N_7630,N_3511,N_1405);
nor U7631 (N_7631,N_1318,N_3391);
xnor U7632 (N_7632,N_3139,N_3314);
xor U7633 (N_7633,N_2814,N_4640);
or U7634 (N_7634,N_1005,N_388);
xor U7635 (N_7635,N_949,N_1421);
or U7636 (N_7636,N_3043,N_4167);
nor U7637 (N_7637,N_633,N_925);
nor U7638 (N_7638,N_2692,N_1705);
nor U7639 (N_7639,N_2736,N_2520);
xnor U7640 (N_7640,N_4004,N_3754);
and U7641 (N_7641,N_1615,N_3195);
nor U7642 (N_7642,N_1939,N_3447);
or U7643 (N_7643,N_1798,N_2661);
nand U7644 (N_7644,N_3852,N_1655);
or U7645 (N_7645,N_4065,N_4974);
nand U7646 (N_7646,N_3258,N_1945);
nand U7647 (N_7647,N_3620,N_3029);
nor U7648 (N_7648,N_4319,N_929);
nand U7649 (N_7649,N_3049,N_4441);
and U7650 (N_7650,N_1410,N_4620);
nand U7651 (N_7651,N_4668,N_603);
xnor U7652 (N_7652,N_1293,N_37);
or U7653 (N_7653,N_2619,N_2081);
nand U7654 (N_7654,N_1705,N_2238);
xnor U7655 (N_7655,N_1342,N_34);
nor U7656 (N_7656,N_1282,N_3494);
and U7657 (N_7657,N_3239,N_604);
or U7658 (N_7658,N_170,N_413);
or U7659 (N_7659,N_4633,N_4213);
nand U7660 (N_7660,N_4309,N_435);
xnor U7661 (N_7661,N_3369,N_3706);
nor U7662 (N_7662,N_2871,N_1607);
nand U7663 (N_7663,N_373,N_4260);
and U7664 (N_7664,N_3024,N_4557);
and U7665 (N_7665,N_1530,N_4202);
and U7666 (N_7666,N_3100,N_4540);
nand U7667 (N_7667,N_3807,N_2475);
nor U7668 (N_7668,N_2749,N_4401);
or U7669 (N_7669,N_2494,N_3432);
nand U7670 (N_7670,N_4043,N_1113);
or U7671 (N_7671,N_2347,N_2070);
or U7672 (N_7672,N_1597,N_96);
and U7673 (N_7673,N_4109,N_361);
xnor U7674 (N_7674,N_3912,N_884);
nand U7675 (N_7675,N_2950,N_3917);
or U7676 (N_7676,N_1755,N_3818);
or U7677 (N_7677,N_1026,N_867);
or U7678 (N_7678,N_3376,N_4923);
nor U7679 (N_7679,N_1604,N_2100);
xnor U7680 (N_7680,N_1824,N_2753);
xor U7681 (N_7681,N_3171,N_3034);
nand U7682 (N_7682,N_1532,N_176);
nand U7683 (N_7683,N_2460,N_1001);
or U7684 (N_7684,N_2635,N_207);
nand U7685 (N_7685,N_2701,N_1978);
or U7686 (N_7686,N_4066,N_902);
or U7687 (N_7687,N_1301,N_191);
xnor U7688 (N_7688,N_1925,N_3599);
xor U7689 (N_7689,N_3110,N_1253);
or U7690 (N_7690,N_4517,N_3016);
nand U7691 (N_7691,N_1535,N_339);
or U7692 (N_7692,N_3592,N_831);
nand U7693 (N_7693,N_1250,N_236);
xor U7694 (N_7694,N_3466,N_3037);
and U7695 (N_7695,N_3173,N_4739);
or U7696 (N_7696,N_1735,N_3526);
nand U7697 (N_7697,N_1344,N_3978);
nor U7698 (N_7698,N_159,N_3542);
and U7699 (N_7699,N_127,N_3258);
or U7700 (N_7700,N_4633,N_2385);
nor U7701 (N_7701,N_4987,N_2764);
or U7702 (N_7702,N_4596,N_395);
nor U7703 (N_7703,N_2424,N_4011);
nor U7704 (N_7704,N_1244,N_4379);
and U7705 (N_7705,N_247,N_2422);
xor U7706 (N_7706,N_684,N_2680);
nand U7707 (N_7707,N_1690,N_3749);
nor U7708 (N_7708,N_3326,N_4507);
and U7709 (N_7709,N_3377,N_4923);
or U7710 (N_7710,N_1494,N_1075);
xnor U7711 (N_7711,N_3030,N_3869);
and U7712 (N_7712,N_2660,N_259);
and U7713 (N_7713,N_1840,N_692);
nor U7714 (N_7714,N_4121,N_3915);
nand U7715 (N_7715,N_3449,N_3234);
or U7716 (N_7716,N_4794,N_4696);
and U7717 (N_7717,N_2653,N_1472);
xnor U7718 (N_7718,N_4837,N_2860);
or U7719 (N_7719,N_3575,N_947);
nand U7720 (N_7720,N_2585,N_1836);
and U7721 (N_7721,N_1739,N_4841);
nor U7722 (N_7722,N_2877,N_980);
nor U7723 (N_7723,N_854,N_2876);
nand U7724 (N_7724,N_340,N_3805);
nand U7725 (N_7725,N_1975,N_1896);
or U7726 (N_7726,N_3490,N_4222);
xnor U7727 (N_7727,N_3084,N_196);
xor U7728 (N_7728,N_2781,N_302);
xor U7729 (N_7729,N_1027,N_3895);
xor U7730 (N_7730,N_2332,N_3029);
nor U7731 (N_7731,N_4264,N_4356);
xor U7732 (N_7732,N_4017,N_1452);
or U7733 (N_7733,N_60,N_3747);
nor U7734 (N_7734,N_2322,N_365);
or U7735 (N_7735,N_341,N_1301);
and U7736 (N_7736,N_1509,N_2851);
nand U7737 (N_7737,N_3543,N_3596);
or U7738 (N_7738,N_4581,N_471);
xor U7739 (N_7739,N_373,N_1219);
nand U7740 (N_7740,N_1327,N_2745);
nand U7741 (N_7741,N_357,N_1536);
nor U7742 (N_7742,N_531,N_280);
xnor U7743 (N_7743,N_3946,N_1776);
xor U7744 (N_7744,N_3866,N_1167);
xor U7745 (N_7745,N_2024,N_2968);
nand U7746 (N_7746,N_1653,N_4087);
and U7747 (N_7747,N_4192,N_3393);
xnor U7748 (N_7748,N_439,N_4979);
or U7749 (N_7749,N_746,N_3775);
nand U7750 (N_7750,N_1627,N_95);
or U7751 (N_7751,N_2283,N_3246);
nand U7752 (N_7752,N_3170,N_2333);
xnor U7753 (N_7753,N_1291,N_466);
and U7754 (N_7754,N_1895,N_4447);
nand U7755 (N_7755,N_3032,N_131);
or U7756 (N_7756,N_212,N_3317);
nor U7757 (N_7757,N_1061,N_3292);
xnor U7758 (N_7758,N_2201,N_4734);
nand U7759 (N_7759,N_505,N_2231);
nor U7760 (N_7760,N_2842,N_4134);
and U7761 (N_7761,N_1474,N_3676);
xnor U7762 (N_7762,N_1560,N_3981);
and U7763 (N_7763,N_2770,N_1458);
xor U7764 (N_7764,N_3530,N_2401);
or U7765 (N_7765,N_4394,N_226);
and U7766 (N_7766,N_1589,N_3966);
xor U7767 (N_7767,N_126,N_4560);
xor U7768 (N_7768,N_1379,N_3506);
or U7769 (N_7769,N_3794,N_3225);
or U7770 (N_7770,N_4806,N_3458);
or U7771 (N_7771,N_1013,N_363);
nor U7772 (N_7772,N_549,N_4817);
xor U7773 (N_7773,N_3029,N_1837);
xnor U7774 (N_7774,N_3109,N_212);
and U7775 (N_7775,N_264,N_1181);
or U7776 (N_7776,N_2165,N_649);
or U7777 (N_7777,N_4289,N_2534);
or U7778 (N_7778,N_365,N_3354);
xnor U7779 (N_7779,N_254,N_1973);
or U7780 (N_7780,N_3298,N_2071);
xor U7781 (N_7781,N_2102,N_4737);
or U7782 (N_7782,N_1835,N_1274);
nor U7783 (N_7783,N_1789,N_2370);
nand U7784 (N_7784,N_2112,N_4198);
and U7785 (N_7785,N_685,N_3710);
and U7786 (N_7786,N_4632,N_3779);
xor U7787 (N_7787,N_3258,N_643);
nor U7788 (N_7788,N_70,N_3506);
or U7789 (N_7789,N_2157,N_512);
nor U7790 (N_7790,N_3451,N_919);
xor U7791 (N_7791,N_4933,N_4849);
and U7792 (N_7792,N_4519,N_4984);
or U7793 (N_7793,N_712,N_3386);
or U7794 (N_7794,N_3830,N_2184);
nand U7795 (N_7795,N_3751,N_2479);
and U7796 (N_7796,N_704,N_3732);
nand U7797 (N_7797,N_3048,N_4620);
nor U7798 (N_7798,N_3554,N_4724);
nor U7799 (N_7799,N_2166,N_3746);
xor U7800 (N_7800,N_3130,N_3752);
xor U7801 (N_7801,N_1270,N_2566);
nand U7802 (N_7802,N_930,N_2775);
xor U7803 (N_7803,N_1997,N_984);
nor U7804 (N_7804,N_2947,N_1758);
or U7805 (N_7805,N_193,N_4258);
or U7806 (N_7806,N_4510,N_4033);
or U7807 (N_7807,N_51,N_4117);
and U7808 (N_7808,N_3411,N_180);
and U7809 (N_7809,N_2348,N_1143);
or U7810 (N_7810,N_3967,N_231);
nor U7811 (N_7811,N_2779,N_3208);
nand U7812 (N_7812,N_2916,N_1779);
nor U7813 (N_7813,N_963,N_349);
xnor U7814 (N_7814,N_260,N_3103);
or U7815 (N_7815,N_1291,N_4751);
xnor U7816 (N_7816,N_4132,N_3908);
xor U7817 (N_7817,N_4364,N_884);
nor U7818 (N_7818,N_3943,N_1196);
xnor U7819 (N_7819,N_1330,N_2313);
xnor U7820 (N_7820,N_1345,N_3364);
or U7821 (N_7821,N_4574,N_3522);
or U7822 (N_7822,N_1051,N_1);
xor U7823 (N_7823,N_77,N_3478);
or U7824 (N_7824,N_783,N_3968);
nand U7825 (N_7825,N_1040,N_1128);
xor U7826 (N_7826,N_207,N_1468);
xnor U7827 (N_7827,N_3852,N_859);
nand U7828 (N_7828,N_1211,N_120);
or U7829 (N_7829,N_433,N_2533);
xor U7830 (N_7830,N_2958,N_1961);
and U7831 (N_7831,N_4910,N_3204);
xor U7832 (N_7832,N_25,N_2417);
xnor U7833 (N_7833,N_52,N_398);
and U7834 (N_7834,N_4759,N_819);
and U7835 (N_7835,N_3657,N_2800);
and U7836 (N_7836,N_3088,N_4626);
and U7837 (N_7837,N_2006,N_3684);
nor U7838 (N_7838,N_4787,N_893);
nand U7839 (N_7839,N_2133,N_2506);
and U7840 (N_7840,N_2157,N_772);
nor U7841 (N_7841,N_1701,N_1310);
nand U7842 (N_7842,N_305,N_4635);
nor U7843 (N_7843,N_3058,N_2787);
xnor U7844 (N_7844,N_2573,N_1403);
xor U7845 (N_7845,N_1359,N_784);
and U7846 (N_7846,N_3356,N_2505);
xor U7847 (N_7847,N_3426,N_4183);
or U7848 (N_7848,N_1626,N_3462);
xnor U7849 (N_7849,N_2888,N_600);
and U7850 (N_7850,N_1178,N_2684);
nand U7851 (N_7851,N_2363,N_637);
or U7852 (N_7852,N_3317,N_1840);
nand U7853 (N_7853,N_1223,N_455);
nand U7854 (N_7854,N_3658,N_3226);
or U7855 (N_7855,N_3735,N_2399);
or U7856 (N_7856,N_3284,N_1202);
or U7857 (N_7857,N_1424,N_2672);
and U7858 (N_7858,N_118,N_4456);
and U7859 (N_7859,N_4252,N_1195);
and U7860 (N_7860,N_4897,N_243);
and U7861 (N_7861,N_532,N_1600);
nand U7862 (N_7862,N_3271,N_2434);
xnor U7863 (N_7863,N_3832,N_2660);
xor U7864 (N_7864,N_747,N_903);
nand U7865 (N_7865,N_1081,N_2542);
nand U7866 (N_7866,N_853,N_4944);
xnor U7867 (N_7867,N_4514,N_4400);
or U7868 (N_7868,N_3033,N_1891);
or U7869 (N_7869,N_4369,N_1129);
and U7870 (N_7870,N_1400,N_1531);
xor U7871 (N_7871,N_1109,N_172);
nand U7872 (N_7872,N_308,N_1694);
nand U7873 (N_7873,N_453,N_117);
and U7874 (N_7874,N_3859,N_3300);
nor U7875 (N_7875,N_375,N_2424);
and U7876 (N_7876,N_1238,N_4744);
nor U7877 (N_7877,N_3232,N_4522);
or U7878 (N_7878,N_1058,N_4247);
nand U7879 (N_7879,N_590,N_850);
or U7880 (N_7880,N_3975,N_2714);
nor U7881 (N_7881,N_3776,N_4344);
and U7882 (N_7882,N_169,N_2955);
or U7883 (N_7883,N_2000,N_1885);
nor U7884 (N_7884,N_580,N_4308);
nand U7885 (N_7885,N_4228,N_2865);
or U7886 (N_7886,N_4846,N_51);
or U7887 (N_7887,N_1329,N_4927);
xnor U7888 (N_7888,N_27,N_4769);
nor U7889 (N_7889,N_1946,N_1709);
nand U7890 (N_7890,N_2219,N_4128);
nor U7891 (N_7891,N_2586,N_4941);
nand U7892 (N_7892,N_1901,N_1572);
xor U7893 (N_7893,N_3741,N_4412);
nand U7894 (N_7894,N_456,N_3061);
xnor U7895 (N_7895,N_3305,N_837);
and U7896 (N_7896,N_2615,N_349);
nor U7897 (N_7897,N_4456,N_4799);
and U7898 (N_7898,N_2539,N_1280);
nor U7899 (N_7899,N_4499,N_4660);
or U7900 (N_7900,N_3261,N_4443);
nand U7901 (N_7901,N_81,N_3369);
nand U7902 (N_7902,N_1558,N_3544);
and U7903 (N_7903,N_3367,N_1049);
xor U7904 (N_7904,N_1680,N_2818);
nor U7905 (N_7905,N_1035,N_1290);
and U7906 (N_7906,N_65,N_1847);
nand U7907 (N_7907,N_3307,N_4492);
or U7908 (N_7908,N_998,N_569);
or U7909 (N_7909,N_3694,N_4625);
nand U7910 (N_7910,N_4569,N_1107);
nor U7911 (N_7911,N_1412,N_4405);
or U7912 (N_7912,N_3929,N_710);
and U7913 (N_7913,N_1769,N_4644);
xor U7914 (N_7914,N_833,N_1509);
or U7915 (N_7915,N_1212,N_2604);
or U7916 (N_7916,N_1906,N_4037);
nor U7917 (N_7917,N_3578,N_711);
and U7918 (N_7918,N_2893,N_1879);
nor U7919 (N_7919,N_2753,N_2173);
nand U7920 (N_7920,N_1803,N_410);
nor U7921 (N_7921,N_2845,N_4349);
or U7922 (N_7922,N_1210,N_476);
or U7923 (N_7923,N_2185,N_1100);
and U7924 (N_7924,N_531,N_4220);
xnor U7925 (N_7925,N_2186,N_3901);
and U7926 (N_7926,N_1533,N_587);
nand U7927 (N_7927,N_1306,N_2207);
nand U7928 (N_7928,N_4933,N_4561);
or U7929 (N_7929,N_1328,N_2051);
nand U7930 (N_7930,N_3045,N_3078);
nor U7931 (N_7931,N_206,N_4558);
xor U7932 (N_7932,N_4552,N_3601);
and U7933 (N_7933,N_1615,N_1214);
nand U7934 (N_7934,N_2700,N_4463);
nand U7935 (N_7935,N_4277,N_2972);
nor U7936 (N_7936,N_3366,N_4807);
and U7937 (N_7937,N_1569,N_1616);
nor U7938 (N_7938,N_2383,N_3528);
nor U7939 (N_7939,N_4074,N_4130);
nand U7940 (N_7940,N_2638,N_630);
xnor U7941 (N_7941,N_785,N_1348);
xor U7942 (N_7942,N_4827,N_3579);
nor U7943 (N_7943,N_2220,N_3955);
xor U7944 (N_7944,N_4072,N_3069);
nor U7945 (N_7945,N_872,N_2338);
nand U7946 (N_7946,N_2927,N_334);
nand U7947 (N_7947,N_4977,N_2744);
nand U7948 (N_7948,N_2706,N_4319);
xnor U7949 (N_7949,N_2513,N_1441);
nand U7950 (N_7950,N_561,N_446);
nand U7951 (N_7951,N_146,N_1773);
xnor U7952 (N_7952,N_2515,N_4085);
or U7953 (N_7953,N_3095,N_2434);
or U7954 (N_7954,N_4810,N_2988);
and U7955 (N_7955,N_3991,N_1011);
xor U7956 (N_7956,N_3411,N_3620);
and U7957 (N_7957,N_2780,N_3913);
nor U7958 (N_7958,N_2003,N_1363);
nor U7959 (N_7959,N_1412,N_4779);
and U7960 (N_7960,N_1563,N_4802);
and U7961 (N_7961,N_1898,N_1303);
or U7962 (N_7962,N_1428,N_2329);
xnor U7963 (N_7963,N_3411,N_392);
nor U7964 (N_7964,N_2810,N_2646);
xnor U7965 (N_7965,N_2633,N_3459);
nor U7966 (N_7966,N_1000,N_194);
nand U7967 (N_7967,N_408,N_4620);
or U7968 (N_7968,N_3985,N_2407);
nand U7969 (N_7969,N_2132,N_2627);
and U7970 (N_7970,N_2445,N_4525);
nor U7971 (N_7971,N_3845,N_2507);
nor U7972 (N_7972,N_4295,N_1485);
xor U7973 (N_7973,N_4289,N_3700);
or U7974 (N_7974,N_3280,N_727);
nor U7975 (N_7975,N_2676,N_4568);
or U7976 (N_7976,N_945,N_386);
and U7977 (N_7977,N_3499,N_3104);
nand U7978 (N_7978,N_2328,N_4766);
nor U7979 (N_7979,N_4470,N_853);
or U7980 (N_7980,N_3052,N_1246);
xnor U7981 (N_7981,N_2135,N_3736);
and U7982 (N_7982,N_1634,N_1860);
and U7983 (N_7983,N_4345,N_1770);
or U7984 (N_7984,N_3680,N_2180);
or U7985 (N_7985,N_3916,N_2143);
xor U7986 (N_7986,N_1210,N_786);
xnor U7987 (N_7987,N_3476,N_2421);
and U7988 (N_7988,N_3738,N_3838);
xnor U7989 (N_7989,N_3647,N_768);
or U7990 (N_7990,N_2570,N_3453);
nand U7991 (N_7991,N_1394,N_2349);
nor U7992 (N_7992,N_2558,N_3489);
and U7993 (N_7993,N_1737,N_4228);
and U7994 (N_7994,N_2674,N_4628);
nand U7995 (N_7995,N_572,N_10);
xor U7996 (N_7996,N_253,N_3639);
nand U7997 (N_7997,N_1465,N_4348);
xor U7998 (N_7998,N_4394,N_4606);
or U7999 (N_7999,N_4255,N_2958);
nor U8000 (N_8000,N_4142,N_1526);
or U8001 (N_8001,N_4360,N_3602);
and U8002 (N_8002,N_4295,N_538);
and U8003 (N_8003,N_4240,N_1846);
nand U8004 (N_8004,N_607,N_3604);
and U8005 (N_8005,N_4119,N_4079);
xnor U8006 (N_8006,N_252,N_3178);
or U8007 (N_8007,N_2669,N_2487);
nand U8008 (N_8008,N_3534,N_1711);
or U8009 (N_8009,N_4597,N_3188);
nor U8010 (N_8010,N_4571,N_3933);
nand U8011 (N_8011,N_2295,N_3429);
and U8012 (N_8012,N_3380,N_2672);
and U8013 (N_8013,N_4738,N_1773);
nand U8014 (N_8014,N_4708,N_1914);
or U8015 (N_8015,N_1323,N_2407);
and U8016 (N_8016,N_282,N_2969);
nand U8017 (N_8017,N_3507,N_4996);
xor U8018 (N_8018,N_1366,N_2409);
or U8019 (N_8019,N_3177,N_3806);
and U8020 (N_8020,N_562,N_12);
nor U8021 (N_8021,N_2302,N_980);
nand U8022 (N_8022,N_4898,N_2759);
nor U8023 (N_8023,N_2309,N_2585);
or U8024 (N_8024,N_4710,N_3283);
nand U8025 (N_8025,N_2211,N_2669);
xor U8026 (N_8026,N_1297,N_2247);
or U8027 (N_8027,N_4290,N_343);
xnor U8028 (N_8028,N_1829,N_3679);
or U8029 (N_8029,N_2994,N_4870);
or U8030 (N_8030,N_28,N_3974);
nor U8031 (N_8031,N_3880,N_768);
or U8032 (N_8032,N_2020,N_410);
or U8033 (N_8033,N_3430,N_4714);
xnor U8034 (N_8034,N_2197,N_64);
xnor U8035 (N_8035,N_319,N_3180);
nor U8036 (N_8036,N_1793,N_4529);
or U8037 (N_8037,N_3111,N_219);
nand U8038 (N_8038,N_919,N_2364);
nor U8039 (N_8039,N_217,N_930);
nand U8040 (N_8040,N_1198,N_3806);
nor U8041 (N_8041,N_1960,N_743);
nor U8042 (N_8042,N_980,N_3642);
nor U8043 (N_8043,N_2951,N_4228);
nor U8044 (N_8044,N_2984,N_1906);
xor U8045 (N_8045,N_3782,N_1422);
and U8046 (N_8046,N_2621,N_1025);
nand U8047 (N_8047,N_2645,N_3353);
or U8048 (N_8048,N_983,N_2512);
xnor U8049 (N_8049,N_1120,N_1920);
nor U8050 (N_8050,N_305,N_13);
nor U8051 (N_8051,N_1360,N_3919);
nor U8052 (N_8052,N_3125,N_4417);
xor U8053 (N_8053,N_463,N_1891);
xor U8054 (N_8054,N_1109,N_924);
and U8055 (N_8055,N_4368,N_1263);
nor U8056 (N_8056,N_1537,N_1514);
and U8057 (N_8057,N_4477,N_3050);
or U8058 (N_8058,N_386,N_3076);
and U8059 (N_8059,N_2691,N_2048);
or U8060 (N_8060,N_4404,N_3363);
nand U8061 (N_8061,N_299,N_2240);
and U8062 (N_8062,N_3829,N_2239);
nand U8063 (N_8063,N_4399,N_3784);
nor U8064 (N_8064,N_2192,N_603);
nor U8065 (N_8065,N_3987,N_4090);
or U8066 (N_8066,N_2049,N_1690);
xnor U8067 (N_8067,N_420,N_7);
xnor U8068 (N_8068,N_1951,N_3227);
xnor U8069 (N_8069,N_4457,N_2761);
xnor U8070 (N_8070,N_4867,N_819);
nor U8071 (N_8071,N_3581,N_3866);
nand U8072 (N_8072,N_1600,N_3384);
and U8073 (N_8073,N_4076,N_337);
nand U8074 (N_8074,N_2933,N_4825);
nor U8075 (N_8075,N_2481,N_3353);
and U8076 (N_8076,N_1255,N_3921);
xor U8077 (N_8077,N_4593,N_2541);
nand U8078 (N_8078,N_2498,N_4968);
nand U8079 (N_8079,N_2602,N_3713);
xor U8080 (N_8080,N_237,N_3435);
nor U8081 (N_8081,N_282,N_3032);
nor U8082 (N_8082,N_1362,N_4582);
or U8083 (N_8083,N_1344,N_2212);
or U8084 (N_8084,N_2865,N_1882);
xor U8085 (N_8085,N_991,N_980);
xnor U8086 (N_8086,N_206,N_3585);
and U8087 (N_8087,N_2424,N_1834);
xor U8088 (N_8088,N_3192,N_4971);
and U8089 (N_8089,N_2402,N_3777);
and U8090 (N_8090,N_1996,N_1109);
and U8091 (N_8091,N_2816,N_3215);
nor U8092 (N_8092,N_4483,N_3867);
nand U8093 (N_8093,N_4993,N_286);
nand U8094 (N_8094,N_2029,N_70);
nand U8095 (N_8095,N_2474,N_183);
nand U8096 (N_8096,N_4284,N_4167);
or U8097 (N_8097,N_26,N_3613);
xnor U8098 (N_8098,N_4070,N_2559);
or U8099 (N_8099,N_2016,N_1863);
or U8100 (N_8100,N_4715,N_2755);
xnor U8101 (N_8101,N_866,N_4018);
and U8102 (N_8102,N_1445,N_3582);
nand U8103 (N_8103,N_3582,N_2651);
and U8104 (N_8104,N_4559,N_1060);
and U8105 (N_8105,N_2101,N_3849);
or U8106 (N_8106,N_1236,N_3623);
and U8107 (N_8107,N_1136,N_1502);
or U8108 (N_8108,N_4194,N_61);
and U8109 (N_8109,N_2270,N_4846);
xor U8110 (N_8110,N_4322,N_2920);
xor U8111 (N_8111,N_2153,N_3655);
or U8112 (N_8112,N_4659,N_2704);
or U8113 (N_8113,N_2353,N_4967);
and U8114 (N_8114,N_3498,N_1363);
or U8115 (N_8115,N_1970,N_2115);
and U8116 (N_8116,N_4426,N_1703);
nand U8117 (N_8117,N_101,N_1981);
or U8118 (N_8118,N_781,N_3982);
or U8119 (N_8119,N_1691,N_2104);
nand U8120 (N_8120,N_1506,N_1914);
xor U8121 (N_8121,N_2992,N_855);
nor U8122 (N_8122,N_465,N_3922);
nor U8123 (N_8123,N_95,N_503);
or U8124 (N_8124,N_2503,N_977);
and U8125 (N_8125,N_4484,N_592);
nand U8126 (N_8126,N_3315,N_2865);
or U8127 (N_8127,N_4508,N_4856);
nor U8128 (N_8128,N_1133,N_2755);
xnor U8129 (N_8129,N_2166,N_3966);
nor U8130 (N_8130,N_3801,N_2385);
or U8131 (N_8131,N_2861,N_926);
xor U8132 (N_8132,N_350,N_2992);
xor U8133 (N_8133,N_2422,N_355);
nor U8134 (N_8134,N_212,N_1903);
or U8135 (N_8135,N_944,N_3622);
nand U8136 (N_8136,N_3565,N_1126);
nor U8137 (N_8137,N_4782,N_3470);
and U8138 (N_8138,N_2267,N_3283);
and U8139 (N_8139,N_2737,N_1807);
nand U8140 (N_8140,N_2211,N_2499);
and U8141 (N_8141,N_4239,N_2665);
nand U8142 (N_8142,N_4173,N_2771);
xnor U8143 (N_8143,N_1651,N_3359);
or U8144 (N_8144,N_1994,N_2043);
nand U8145 (N_8145,N_2433,N_3357);
nor U8146 (N_8146,N_561,N_3833);
nand U8147 (N_8147,N_3615,N_352);
nand U8148 (N_8148,N_896,N_4126);
nand U8149 (N_8149,N_938,N_2046);
xor U8150 (N_8150,N_2578,N_3495);
nand U8151 (N_8151,N_704,N_4584);
nand U8152 (N_8152,N_1131,N_1364);
or U8153 (N_8153,N_425,N_3753);
nand U8154 (N_8154,N_2726,N_262);
nand U8155 (N_8155,N_2298,N_2868);
or U8156 (N_8156,N_1120,N_672);
and U8157 (N_8157,N_1259,N_1769);
or U8158 (N_8158,N_2486,N_1478);
nand U8159 (N_8159,N_552,N_985);
or U8160 (N_8160,N_889,N_4250);
nand U8161 (N_8161,N_19,N_2231);
xor U8162 (N_8162,N_1601,N_997);
xor U8163 (N_8163,N_3596,N_678);
nand U8164 (N_8164,N_935,N_4731);
xnor U8165 (N_8165,N_4882,N_4470);
or U8166 (N_8166,N_3143,N_2140);
nor U8167 (N_8167,N_3294,N_3240);
nor U8168 (N_8168,N_3092,N_2971);
nand U8169 (N_8169,N_4812,N_2747);
xnor U8170 (N_8170,N_3215,N_3070);
nand U8171 (N_8171,N_4737,N_4124);
nor U8172 (N_8172,N_2776,N_663);
and U8173 (N_8173,N_2567,N_4925);
xor U8174 (N_8174,N_3405,N_765);
or U8175 (N_8175,N_4184,N_111);
and U8176 (N_8176,N_4674,N_4935);
nand U8177 (N_8177,N_2815,N_2575);
nor U8178 (N_8178,N_927,N_1558);
or U8179 (N_8179,N_1165,N_2107);
nand U8180 (N_8180,N_508,N_1442);
nand U8181 (N_8181,N_1835,N_4319);
and U8182 (N_8182,N_2905,N_2935);
nand U8183 (N_8183,N_1053,N_3587);
nand U8184 (N_8184,N_1304,N_2692);
nor U8185 (N_8185,N_4424,N_3338);
and U8186 (N_8186,N_52,N_3671);
nor U8187 (N_8187,N_2848,N_268);
nand U8188 (N_8188,N_2410,N_2481);
nand U8189 (N_8189,N_2350,N_2942);
nor U8190 (N_8190,N_2515,N_1363);
nand U8191 (N_8191,N_1172,N_1398);
nand U8192 (N_8192,N_413,N_2641);
nand U8193 (N_8193,N_176,N_4406);
nor U8194 (N_8194,N_1202,N_15);
nor U8195 (N_8195,N_3007,N_2487);
nor U8196 (N_8196,N_1773,N_4953);
nor U8197 (N_8197,N_645,N_3299);
and U8198 (N_8198,N_2733,N_1070);
and U8199 (N_8199,N_2799,N_3047);
and U8200 (N_8200,N_4610,N_2804);
nand U8201 (N_8201,N_3047,N_2136);
xor U8202 (N_8202,N_2082,N_1596);
and U8203 (N_8203,N_3235,N_1102);
or U8204 (N_8204,N_2543,N_3093);
nand U8205 (N_8205,N_4114,N_2930);
and U8206 (N_8206,N_1783,N_1170);
xnor U8207 (N_8207,N_126,N_1761);
nand U8208 (N_8208,N_1732,N_2016);
and U8209 (N_8209,N_4378,N_73);
xor U8210 (N_8210,N_3,N_4796);
xnor U8211 (N_8211,N_3172,N_3855);
xor U8212 (N_8212,N_105,N_2794);
xnor U8213 (N_8213,N_2903,N_4225);
nand U8214 (N_8214,N_4780,N_318);
and U8215 (N_8215,N_3913,N_2404);
xnor U8216 (N_8216,N_2379,N_954);
nand U8217 (N_8217,N_541,N_1456);
nor U8218 (N_8218,N_2380,N_833);
xor U8219 (N_8219,N_4181,N_2462);
xnor U8220 (N_8220,N_2326,N_1958);
xnor U8221 (N_8221,N_2248,N_2898);
nand U8222 (N_8222,N_1809,N_1106);
nor U8223 (N_8223,N_4892,N_2457);
xor U8224 (N_8224,N_3578,N_2914);
and U8225 (N_8225,N_4652,N_3958);
or U8226 (N_8226,N_2207,N_4693);
xor U8227 (N_8227,N_2750,N_283);
nor U8228 (N_8228,N_4806,N_2272);
or U8229 (N_8229,N_1790,N_4503);
and U8230 (N_8230,N_1764,N_993);
and U8231 (N_8231,N_1936,N_2789);
and U8232 (N_8232,N_2441,N_746);
nor U8233 (N_8233,N_1924,N_2389);
and U8234 (N_8234,N_4996,N_4946);
xnor U8235 (N_8235,N_1847,N_710);
or U8236 (N_8236,N_1173,N_3366);
nand U8237 (N_8237,N_2361,N_4917);
and U8238 (N_8238,N_2505,N_1284);
and U8239 (N_8239,N_3248,N_393);
and U8240 (N_8240,N_2177,N_3303);
xnor U8241 (N_8241,N_1587,N_3374);
and U8242 (N_8242,N_3213,N_3875);
and U8243 (N_8243,N_2144,N_2104);
xor U8244 (N_8244,N_1365,N_4590);
xor U8245 (N_8245,N_3819,N_2161);
nand U8246 (N_8246,N_2659,N_889);
nand U8247 (N_8247,N_2054,N_4502);
or U8248 (N_8248,N_4178,N_4837);
or U8249 (N_8249,N_4657,N_3420);
nand U8250 (N_8250,N_4332,N_847);
and U8251 (N_8251,N_4813,N_1708);
nor U8252 (N_8252,N_4213,N_4889);
xnor U8253 (N_8253,N_4575,N_3461);
nand U8254 (N_8254,N_2519,N_4721);
xor U8255 (N_8255,N_4485,N_1907);
or U8256 (N_8256,N_4841,N_77);
nand U8257 (N_8257,N_568,N_683);
or U8258 (N_8258,N_1394,N_4701);
or U8259 (N_8259,N_1502,N_1551);
and U8260 (N_8260,N_3666,N_1653);
and U8261 (N_8261,N_4011,N_2974);
and U8262 (N_8262,N_1735,N_4104);
or U8263 (N_8263,N_743,N_1674);
or U8264 (N_8264,N_3687,N_2720);
nand U8265 (N_8265,N_2560,N_2126);
nor U8266 (N_8266,N_3997,N_769);
and U8267 (N_8267,N_305,N_3805);
nand U8268 (N_8268,N_982,N_2292);
xor U8269 (N_8269,N_2655,N_4968);
and U8270 (N_8270,N_267,N_1590);
nand U8271 (N_8271,N_3037,N_2445);
nor U8272 (N_8272,N_1861,N_489);
xnor U8273 (N_8273,N_1681,N_503);
and U8274 (N_8274,N_1104,N_1851);
and U8275 (N_8275,N_2021,N_613);
or U8276 (N_8276,N_776,N_1707);
nand U8277 (N_8277,N_2733,N_590);
or U8278 (N_8278,N_583,N_1242);
and U8279 (N_8279,N_1461,N_2114);
or U8280 (N_8280,N_3100,N_131);
or U8281 (N_8281,N_275,N_2537);
nor U8282 (N_8282,N_582,N_1515);
xor U8283 (N_8283,N_1313,N_3935);
and U8284 (N_8284,N_4151,N_3896);
nand U8285 (N_8285,N_4381,N_4023);
and U8286 (N_8286,N_1897,N_649);
or U8287 (N_8287,N_911,N_4254);
xor U8288 (N_8288,N_4421,N_4324);
xor U8289 (N_8289,N_1213,N_3275);
and U8290 (N_8290,N_4261,N_53);
nand U8291 (N_8291,N_3374,N_396);
or U8292 (N_8292,N_725,N_2096);
or U8293 (N_8293,N_1011,N_3471);
nor U8294 (N_8294,N_883,N_3125);
xnor U8295 (N_8295,N_251,N_273);
nand U8296 (N_8296,N_3915,N_2296);
or U8297 (N_8297,N_2154,N_567);
nand U8298 (N_8298,N_3098,N_3682);
or U8299 (N_8299,N_1168,N_2313);
nand U8300 (N_8300,N_4453,N_3584);
nand U8301 (N_8301,N_1624,N_2341);
xnor U8302 (N_8302,N_2487,N_2692);
nor U8303 (N_8303,N_455,N_2607);
nor U8304 (N_8304,N_1968,N_1807);
nand U8305 (N_8305,N_4108,N_2402);
nor U8306 (N_8306,N_769,N_2779);
nand U8307 (N_8307,N_2777,N_3243);
or U8308 (N_8308,N_467,N_2600);
nor U8309 (N_8309,N_1591,N_855);
nor U8310 (N_8310,N_2359,N_197);
or U8311 (N_8311,N_217,N_119);
xnor U8312 (N_8312,N_610,N_507);
xor U8313 (N_8313,N_3946,N_1044);
and U8314 (N_8314,N_2057,N_1090);
and U8315 (N_8315,N_717,N_95);
nand U8316 (N_8316,N_2684,N_1624);
and U8317 (N_8317,N_1027,N_42);
or U8318 (N_8318,N_4385,N_1587);
nor U8319 (N_8319,N_269,N_1951);
nand U8320 (N_8320,N_3670,N_4885);
and U8321 (N_8321,N_1117,N_4132);
or U8322 (N_8322,N_3771,N_4040);
and U8323 (N_8323,N_4839,N_1819);
xnor U8324 (N_8324,N_594,N_4311);
xor U8325 (N_8325,N_1447,N_1332);
and U8326 (N_8326,N_2594,N_4942);
or U8327 (N_8327,N_3563,N_3186);
and U8328 (N_8328,N_4116,N_3689);
nor U8329 (N_8329,N_484,N_4870);
and U8330 (N_8330,N_4642,N_172);
nand U8331 (N_8331,N_544,N_2715);
xnor U8332 (N_8332,N_4016,N_2578);
or U8333 (N_8333,N_3746,N_1431);
xnor U8334 (N_8334,N_3605,N_1620);
and U8335 (N_8335,N_3717,N_267);
or U8336 (N_8336,N_1732,N_260);
nand U8337 (N_8337,N_4157,N_4437);
or U8338 (N_8338,N_4684,N_3191);
and U8339 (N_8339,N_4198,N_753);
and U8340 (N_8340,N_2868,N_2662);
xnor U8341 (N_8341,N_1554,N_4093);
and U8342 (N_8342,N_1145,N_55);
or U8343 (N_8343,N_2573,N_1482);
and U8344 (N_8344,N_789,N_2751);
nand U8345 (N_8345,N_1064,N_2197);
and U8346 (N_8346,N_1398,N_2937);
and U8347 (N_8347,N_345,N_2930);
or U8348 (N_8348,N_4000,N_1778);
nor U8349 (N_8349,N_4521,N_690);
and U8350 (N_8350,N_1946,N_467);
and U8351 (N_8351,N_4836,N_1731);
nand U8352 (N_8352,N_3777,N_745);
or U8353 (N_8353,N_4349,N_3155);
and U8354 (N_8354,N_1786,N_4561);
or U8355 (N_8355,N_3888,N_587);
and U8356 (N_8356,N_1083,N_1009);
and U8357 (N_8357,N_3113,N_4971);
nand U8358 (N_8358,N_514,N_370);
or U8359 (N_8359,N_1648,N_3835);
xor U8360 (N_8360,N_343,N_875);
and U8361 (N_8361,N_2206,N_2634);
nor U8362 (N_8362,N_2858,N_3847);
or U8363 (N_8363,N_3197,N_2252);
nor U8364 (N_8364,N_1827,N_2150);
xor U8365 (N_8365,N_3880,N_4864);
nand U8366 (N_8366,N_3551,N_2781);
or U8367 (N_8367,N_507,N_2683);
nor U8368 (N_8368,N_1039,N_4881);
nor U8369 (N_8369,N_1910,N_2049);
and U8370 (N_8370,N_2394,N_2051);
or U8371 (N_8371,N_2952,N_4951);
and U8372 (N_8372,N_3113,N_3881);
or U8373 (N_8373,N_3037,N_3453);
nand U8374 (N_8374,N_1548,N_3480);
nor U8375 (N_8375,N_495,N_1657);
nand U8376 (N_8376,N_25,N_1183);
xor U8377 (N_8377,N_4396,N_3507);
nor U8378 (N_8378,N_4454,N_2071);
or U8379 (N_8379,N_491,N_2003);
nor U8380 (N_8380,N_3645,N_1522);
nand U8381 (N_8381,N_1533,N_2367);
or U8382 (N_8382,N_4001,N_1250);
nand U8383 (N_8383,N_863,N_1669);
nand U8384 (N_8384,N_305,N_1866);
and U8385 (N_8385,N_3281,N_4357);
nand U8386 (N_8386,N_2069,N_1080);
xnor U8387 (N_8387,N_3591,N_574);
and U8388 (N_8388,N_1349,N_1875);
nor U8389 (N_8389,N_2344,N_1008);
or U8390 (N_8390,N_533,N_1945);
and U8391 (N_8391,N_1843,N_202);
nand U8392 (N_8392,N_370,N_3823);
nand U8393 (N_8393,N_4847,N_1907);
or U8394 (N_8394,N_575,N_911);
or U8395 (N_8395,N_2945,N_4530);
nand U8396 (N_8396,N_3746,N_2229);
xor U8397 (N_8397,N_345,N_2418);
nor U8398 (N_8398,N_2074,N_262);
xor U8399 (N_8399,N_2752,N_4865);
and U8400 (N_8400,N_406,N_4970);
nand U8401 (N_8401,N_4879,N_3495);
or U8402 (N_8402,N_1845,N_494);
xor U8403 (N_8403,N_3864,N_2544);
nand U8404 (N_8404,N_2037,N_2032);
and U8405 (N_8405,N_147,N_4838);
nand U8406 (N_8406,N_1140,N_2298);
nor U8407 (N_8407,N_854,N_3689);
and U8408 (N_8408,N_4208,N_233);
nand U8409 (N_8409,N_3369,N_3132);
nor U8410 (N_8410,N_2867,N_4700);
xnor U8411 (N_8411,N_1908,N_3056);
nor U8412 (N_8412,N_3580,N_4933);
and U8413 (N_8413,N_598,N_1199);
or U8414 (N_8414,N_4697,N_2593);
nand U8415 (N_8415,N_893,N_2067);
xor U8416 (N_8416,N_1464,N_1935);
and U8417 (N_8417,N_3765,N_4102);
or U8418 (N_8418,N_1548,N_1779);
nor U8419 (N_8419,N_3992,N_858);
nor U8420 (N_8420,N_1598,N_19);
or U8421 (N_8421,N_2406,N_2273);
and U8422 (N_8422,N_486,N_4697);
or U8423 (N_8423,N_2823,N_1811);
and U8424 (N_8424,N_1899,N_399);
or U8425 (N_8425,N_866,N_1452);
xor U8426 (N_8426,N_2123,N_4568);
or U8427 (N_8427,N_387,N_4648);
xnor U8428 (N_8428,N_2430,N_4656);
xor U8429 (N_8429,N_368,N_1193);
xnor U8430 (N_8430,N_1103,N_1626);
nand U8431 (N_8431,N_1363,N_4319);
or U8432 (N_8432,N_3522,N_2528);
xor U8433 (N_8433,N_1520,N_2234);
nor U8434 (N_8434,N_4985,N_3359);
nand U8435 (N_8435,N_1230,N_2214);
nand U8436 (N_8436,N_2998,N_767);
nand U8437 (N_8437,N_3886,N_2166);
xnor U8438 (N_8438,N_541,N_4633);
and U8439 (N_8439,N_2525,N_3055);
or U8440 (N_8440,N_2864,N_2721);
and U8441 (N_8441,N_3632,N_339);
nor U8442 (N_8442,N_4843,N_1189);
nand U8443 (N_8443,N_4642,N_3586);
nand U8444 (N_8444,N_3406,N_4907);
nor U8445 (N_8445,N_1686,N_2868);
nor U8446 (N_8446,N_369,N_1940);
xnor U8447 (N_8447,N_196,N_2279);
and U8448 (N_8448,N_3713,N_2928);
or U8449 (N_8449,N_153,N_3606);
nand U8450 (N_8450,N_1007,N_2277);
nand U8451 (N_8451,N_2070,N_1401);
nand U8452 (N_8452,N_2076,N_1424);
and U8453 (N_8453,N_1554,N_309);
nor U8454 (N_8454,N_4969,N_4836);
or U8455 (N_8455,N_2298,N_3022);
nand U8456 (N_8456,N_4570,N_2892);
and U8457 (N_8457,N_2344,N_4461);
or U8458 (N_8458,N_4691,N_938);
nor U8459 (N_8459,N_2128,N_2522);
and U8460 (N_8460,N_4099,N_4240);
nor U8461 (N_8461,N_401,N_2404);
xnor U8462 (N_8462,N_4714,N_4421);
and U8463 (N_8463,N_688,N_4862);
xnor U8464 (N_8464,N_2540,N_475);
or U8465 (N_8465,N_2689,N_2067);
or U8466 (N_8466,N_1666,N_4953);
nand U8467 (N_8467,N_3399,N_225);
nand U8468 (N_8468,N_3203,N_2871);
nand U8469 (N_8469,N_1657,N_2924);
and U8470 (N_8470,N_2114,N_3357);
and U8471 (N_8471,N_992,N_4888);
nor U8472 (N_8472,N_421,N_532);
and U8473 (N_8473,N_914,N_1575);
xnor U8474 (N_8474,N_3514,N_2414);
xor U8475 (N_8475,N_1030,N_325);
xor U8476 (N_8476,N_1038,N_2590);
nand U8477 (N_8477,N_3613,N_2176);
and U8478 (N_8478,N_956,N_567);
and U8479 (N_8479,N_4118,N_234);
and U8480 (N_8480,N_3444,N_3991);
and U8481 (N_8481,N_4575,N_80);
nor U8482 (N_8482,N_4941,N_1552);
or U8483 (N_8483,N_1364,N_4958);
and U8484 (N_8484,N_2115,N_4236);
and U8485 (N_8485,N_3279,N_983);
and U8486 (N_8486,N_1260,N_1988);
nand U8487 (N_8487,N_363,N_4455);
nor U8488 (N_8488,N_3040,N_1908);
and U8489 (N_8489,N_2231,N_2043);
nor U8490 (N_8490,N_247,N_488);
or U8491 (N_8491,N_2618,N_3205);
nand U8492 (N_8492,N_2362,N_559);
xnor U8493 (N_8493,N_4133,N_3329);
xnor U8494 (N_8494,N_1838,N_2311);
nand U8495 (N_8495,N_607,N_4968);
nor U8496 (N_8496,N_2487,N_897);
nand U8497 (N_8497,N_2037,N_2920);
xor U8498 (N_8498,N_601,N_987);
nand U8499 (N_8499,N_4072,N_3735);
or U8500 (N_8500,N_3519,N_4221);
nor U8501 (N_8501,N_2196,N_1592);
nand U8502 (N_8502,N_582,N_1604);
nand U8503 (N_8503,N_910,N_3308);
nor U8504 (N_8504,N_2721,N_4107);
nor U8505 (N_8505,N_1699,N_1136);
xor U8506 (N_8506,N_2438,N_4365);
xnor U8507 (N_8507,N_2586,N_973);
xnor U8508 (N_8508,N_3449,N_1896);
xor U8509 (N_8509,N_4754,N_1504);
or U8510 (N_8510,N_1437,N_2513);
nand U8511 (N_8511,N_466,N_2148);
nor U8512 (N_8512,N_88,N_408);
or U8513 (N_8513,N_3499,N_1370);
nand U8514 (N_8514,N_3972,N_34);
or U8515 (N_8515,N_392,N_3097);
and U8516 (N_8516,N_284,N_3960);
and U8517 (N_8517,N_2624,N_2849);
nand U8518 (N_8518,N_3331,N_2049);
xor U8519 (N_8519,N_2332,N_3787);
xor U8520 (N_8520,N_1247,N_258);
nand U8521 (N_8521,N_4934,N_4638);
and U8522 (N_8522,N_1503,N_99);
nor U8523 (N_8523,N_2443,N_2070);
nor U8524 (N_8524,N_3535,N_4237);
or U8525 (N_8525,N_441,N_3648);
xor U8526 (N_8526,N_4506,N_197);
or U8527 (N_8527,N_3336,N_3382);
and U8528 (N_8528,N_1951,N_1166);
or U8529 (N_8529,N_1484,N_3371);
and U8530 (N_8530,N_750,N_433);
nor U8531 (N_8531,N_1706,N_9);
nor U8532 (N_8532,N_3506,N_4689);
and U8533 (N_8533,N_3642,N_20);
nand U8534 (N_8534,N_449,N_2340);
or U8535 (N_8535,N_3457,N_1134);
and U8536 (N_8536,N_309,N_2846);
xnor U8537 (N_8537,N_2385,N_4780);
xor U8538 (N_8538,N_655,N_4663);
or U8539 (N_8539,N_4281,N_1020);
nand U8540 (N_8540,N_1319,N_1148);
or U8541 (N_8541,N_1082,N_70);
xnor U8542 (N_8542,N_4513,N_2788);
nor U8543 (N_8543,N_882,N_2651);
or U8544 (N_8544,N_1579,N_800);
and U8545 (N_8545,N_2020,N_1935);
nor U8546 (N_8546,N_1412,N_3539);
nand U8547 (N_8547,N_1617,N_1110);
and U8548 (N_8548,N_1422,N_4845);
nand U8549 (N_8549,N_4956,N_962);
or U8550 (N_8550,N_2018,N_4121);
and U8551 (N_8551,N_1127,N_4291);
and U8552 (N_8552,N_1524,N_202);
nand U8553 (N_8553,N_4577,N_3893);
nand U8554 (N_8554,N_1022,N_2005);
or U8555 (N_8555,N_1454,N_2);
xnor U8556 (N_8556,N_509,N_3374);
nor U8557 (N_8557,N_4110,N_4645);
nand U8558 (N_8558,N_2722,N_1593);
and U8559 (N_8559,N_3435,N_4793);
nor U8560 (N_8560,N_4520,N_4869);
or U8561 (N_8561,N_3127,N_3892);
nor U8562 (N_8562,N_3371,N_1712);
nand U8563 (N_8563,N_2389,N_4613);
xnor U8564 (N_8564,N_3720,N_126);
nor U8565 (N_8565,N_3607,N_2680);
xnor U8566 (N_8566,N_4017,N_1555);
nor U8567 (N_8567,N_1292,N_2359);
xnor U8568 (N_8568,N_766,N_3610);
xor U8569 (N_8569,N_4688,N_4286);
xnor U8570 (N_8570,N_879,N_4702);
nand U8571 (N_8571,N_3449,N_1180);
or U8572 (N_8572,N_2065,N_4235);
nand U8573 (N_8573,N_2869,N_955);
xor U8574 (N_8574,N_1397,N_3765);
and U8575 (N_8575,N_2475,N_2497);
and U8576 (N_8576,N_2320,N_4210);
and U8577 (N_8577,N_3209,N_4228);
and U8578 (N_8578,N_774,N_2066);
and U8579 (N_8579,N_3275,N_1890);
and U8580 (N_8580,N_2086,N_4164);
or U8581 (N_8581,N_2006,N_4158);
nor U8582 (N_8582,N_355,N_2462);
and U8583 (N_8583,N_910,N_525);
and U8584 (N_8584,N_1428,N_429);
or U8585 (N_8585,N_2369,N_3007);
xor U8586 (N_8586,N_2296,N_3002);
or U8587 (N_8587,N_3048,N_1440);
nand U8588 (N_8588,N_826,N_2382);
nand U8589 (N_8589,N_2078,N_4393);
and U8590 (N_8590,N_70,N_2471);
xnor U8591 (N_8591,N_1690,N_1421);
nor U8592 (N_8592,N_4393,N_596);
or U8593 (N_8593,N_1805,N_3051);
nor U8594 (N_8594,N_3429,N_920);
xor U8595 (N_8595,N_1284,N_3513);
nand U8596 (N_8596,N_1964,N_3119);
or U8597 (N_8597,N_3362,N_404);
or U8598 (N_8598,N_3636,N_3011);
or U8599 (N_8599,N_136,N_781);
nand U8600 (N_8600,N_2318,N_4954);
or U8601 (N_8601,N_4445,N_289);
or U8602 (N_8602,N_1138,N_2433);
nor U8603 (N_8603,N_4492,N_2605);
xnor U8604 (N_8604,N_4412,N_622);
and U8605 (N_8605,N_1604,N_1348);
or U8606 (N_8606,N_1647,N_2067);
and U8607 (N_8607,N_3442,N_3242);
nand U8608 (N_8608,N_2860,N_4659);
xor U8609 (N_8609,N_1386,N_696);
nand U8610 (N_8610,N_751,N_643);
nor U8611 (N_8611,N_2046,N_3328);
nand U8612 (N_8612,N_1393,N_4566);
nand U8613 (N_8613,N_4053,N_2776);
xnor U8614 (N_8614,N_2545,N_942);
and U8615 (N_8615,N_2322,N_142);
nor U8616 (N_8616,N_4880,N_4833);
nor U8617 (N_8617,N_1666,N_3998);
nand U8618 (N_8618,N_453,N_1587);
nor U8619 (N_8619,N_2513,N_2273);
nor U8620 (N_8620,N_3815,N_4567);
nand U8621 (N_8621,N_1784,N_3612);
xnor U8622 (N_8622,N_672,N_267);
nand U8623 (N_8623,N_463,N_395);
and U8624 (N_8624,N_3524,N_1182);
or U8625 (N_8625,N_557,N_4685);
nor U8626 (N_8626,N_1469,N_1270);
or U8627 (N_8627,N_320,N_2866);
nand U8628 (N_8628,N_2467,N_3988);
xnor U8629 (N_8629,N_1244,N_2652);
nor U8630 (N_8630,N_1437,N_757);
nand U8631 (N_8631,N_2102,N_4480);
nor U8632 (N_8632,N_3388,N_2999);
xnor U8633 (N_8633,N_3438,N_365);
or U8634 (N_8634,N_2999,N_2098);
or U8635 (N_8635,N_3552,N_4669);
xor U8636 (N_8636,N_1787,N_1139);
and U8637 (N_8637,N_3799,N_1482);
nor U8638 (N_8638,N_1478,N_3852);
or U8639 (N_8639,N_2920,N_844);
nand U8640 (N_8640,N_2868,N_3740);
nand U8641 (N_8641,N_3546,N_4860);
or U8642 (N_8642,N_4022,N_4270);
xor U8643 (N_8643,N_3792,N_4430);
xnor U8644 (N_8644,N_1490,N_4242);
and U8645 (N_8645,N_3639,N_193);
nand U8646 (N_8646,N_3858,N_3538);
nor U8647 (N_8647,N_1977,N_13);
nand U8648 (N_8648,N_996,N_3788);
and U8649 (N_8649,N_668,N_2431);
and U8650 (N_8650,N_2273,N_43);
nand U8651 (N_8651,N_3033,N_400);
and U8652 (N_8652,N_2535,N_2385);
and U8653 (N_8653,N_1835,N_12);
nor U8654 (N_8654,N_2142,N_4543);
xnor U8655 (N_8655,N_2002,N_2431);
or U8656 (N_8656,N_2147,N_4253);
nand U8657 (N_8657,N_3297,N_2668);
nand U8658 (N_8658,N_2067,N_362);
xnor U8659 (N_8659,N_3330,N_324);
or U8660 (N_8660,N_4657,N_2743);
nand U8661 (N_8661,N_1983,N_1871);
and U8662 (N_8662,N_3605,N_3896);
nor U8663 (N_8663,N_2668,N_4607);
or U8664 (N_8664,N_2461,N_191);
and U8665 (N_8665,N_3185,N_1369);
nand U8666 (N_8666,N_4041,N_1172);
and U8667 (N_8667,N_3775,N_4159);
and U8668 (N_8668,N_1964,N_4141);
nand U8669 (N_8669,N_4055,N_3964);
nor U8670 (N_8670,N_4006,N_1785);
nand U8671 (N_8671,N_252,N_2985);
nand U8672 (N_8672,N_1671,N_2358);
or U8673 (N_8673,N_3429,N_3326);
nor U8674 (N_8674,N_3069,N_213);
and U8675 (N_8675,N_2533,N_3364);
xnor U8676 (N_8676,N_3269,N_4280);
nor U8677 (N_8677,N_4101,N_2869);
and U8678 (N_8678,N_1816,N_4491);
and U8679 (N_8679,N_4955,N_4443);
xor U8680 (N_8680,N_1015,N_1136);
nand U8681 (N_8681,N_807,N_3918);
nand U8682 (N_8682,N_3633,N_1536);
nand U8683 (N_8683,N_1269,N_3333);
xor U8684 (N_8684,N_3889,N_2981);
and U8685 (N_8685,N_416,N_2375);
and U8686 (N_8686,N_2294,N_1265);
nand U8687 (N_8687,N_2406,N_2721);
or U8688 (N_8688,N_4556,N_3348);
xnor U8689 (N_8689,N_3004,N_1073);
xnor U8690 (N_8690,N_4906,N_3210);
and U8691 (N_8691,N_1331,N_4651);
and U8692 (N_8692,N_3308,N_1615);
or U8693 (N_8693,N_1343,N_1501);
nor U8694 (N_8694,N_4825,N_3104);
or U8695 (N_8695,N_4460,N_4371);
nor U8696 (N_8696,N_328,N_2751);
xnor U8697 (N_8697,N_758,N_3511);
nor U8698 (N_8698,N_1886,N_360);
nor U8699 (N_8699,N_1777,N_629);
xor U8700 (N_8700,N_3423,N_1080);
nor U8701 (N_8701,N_4044,N_996);
xor U8702 (N_8702,N_2937,N_973);
nand U8703 (N_8703,N_2574,N_4036);
nand U8704 (N_8704,N_3236,N_4492);
xor U8705 (N_8705,N_1638,N_373);
nor U8706 (N_8706,N_4692,N_1683);
xnor U8707 (N_8707,N_1704,N_2801);
or U8708 (N_8708,N_4800,N_2707);
nor U8709 (N_8709,N_557,N_2612);
xnor U8710 (N_8710,N_1141,N_1723);
or U8711 (N_8711,N_327,N_1494);
or U8712 (N_8712,N_2193,N_909);
nand U8713 (N_8713,N_792,N_3185);
and U8714 (N_8714,N_3835,N_2776);
and U8715 (N_8715,N_4145,N_2556);
and U8716 (N_8716,N_2843,N_868);
or U8717 (N_8717,N_2878,N_3740);
or U8718 (N_8718,N_975,N_1182);
or U8719 (N_8719,N_3918,N_1438);
nor U8720 (N_8720,N_4371,N_2443);
nand U8721 (N_8721,N_1216,N_300);
nor U8722 (N_8722,N_469,N_3005);
and U8723 (N_8723,N_929,N_1604);
nor U8724 (N_8724,N_1685,N_3759);
xor U8725 (N_8725,N_2525,N_1079);
and U8726 (N_8726,N_898,N_2458);
nand U8727 (N_8727,N_3462,N_1509);
nand U8728 (N_8728,N_1221,N_1048);
or U8729 (N_8729,N_103,N_2318);
xnor U8730 (N_8730,N_3938,N_1371);
and U8731 (N_8731,N_1748,N_2042);
nor U8732 (N_8732,N_2618,N_1198);
nand U8733 (N_8733,N_1247,N_3117);
nand U8734 (N_8734,N_3870,N_3544);
or U8735 (N_8735,N_2735,N_2642);
and U8736 (N_8736,N_1062,N_1575);
nand U8737 (N_8737,N_2285,N_3181);
and U8738 (N_8738,N_2593,N_3729);
xnor U8739 (N_8739,N_4615,N_605);
and U8740 (N_8740,N_467,N_3595);
and U8741 (N_8741,N_1894,N_407);
xnor U8742 (N_8742,N_2241,N_1348);
or U8743 (N_8743,N_3146,N_3509);
nand U8744 (N_8744,N_2819,N_3805);
or U8745 (N_8745,N_2791,N_4961);
and U8746 (N_8746,N_3912,N_498);
nor U8747 (N_8747,N_2116,N_4924);
xor U8748 (N_8748,N_2676,N_3719);
and U8749 (N_8749,N_1811,N_45);
nor U8750 (N_8750,N_4024,N_4499);
or U8751 (N_8751,N_4452,N_4241);
or U8752 (N_8752,N_4609,N_2936);
or U8753 (N_8753,N_4794,N_2004);
and U8754 (N_8754,N_1423,N_4901);
nand U8755 (N_8755,N_4376,N_4149);
nor U8756 (N_8756,N_804,N_2406);
or U8757 (N_8757,N_1588,N_1492);
xor U8758 (N_8758,N_3278,N_3083);
nand U8759 (N_8759,N_3955,N_3085);
nor U8760 (N_8760,N_3474,N_2453);
nand U8761 (N_8761,N_2124,N_2036);
or U8762 (N_8762,N_4013,N_51);
and U8763 (N_8763,N_4436,N_2633);
xnor U8764 (N_8764,N_611,N_1616);
nor U8765 (N_8765,N_1678,N_4385);
or U8766 (N_8766,N_2438,N_2951);
and U8767 (N_8767,N_1687,N_1033);
or U8768 (N_8768,N_3266,N_3374);
and U8769 (N_8769,N_687,N_3549);
xnor U8770 (N_8770,N_2665,N_4934);
and U8771 (N_8771,N_3741,N_1413);
nor U8772 (N_8772,N_2435,N_775);
xor U8773 (N_8773,N_1534,N_3083);
or U8774 (N_8774,N_4351,N_2846);
or U8775 (N_8775,N_3425,N_637);
nor U8776 (N_8776,N_1356,N_111);
and U8777 (N_8777,N_1599,N_1903);
and U8778 (N_8778,N_484,N_1854);
xnor U8779 (N_8779,N_1691,N_2665);
and U8780 (N_8780,N_3384,N_524);
and U8781 (N_8781,N_1209,N_715);
and U8782 (N_8782,N_2485,N_1987);
nor U8783 (N_8783,N_2148,N_2451);
nand U8784 (N_8784,N_4896,N_2847);
and U8785 (N_8785,N_632,N_71);
nor U8786 (N_8786,N_2128,N_3573);
nand U8787 (N_8787,N_4215,N_3198);
xor U8788 (N_8788,N_2556,N_2226);
and U8789 (N_8789,N_3522,N_783);
or U8790 (N_8790,N_3422,N_4189);
nor U8791 (N_8791,N_1763,N_1918);
nand U8792 (N_8792,N_951,N_663);
nor U8793 (N_8793,N_112,N_175);
or U8794 (N_8794,N_4048,N_2600);
nand U8795 (N_8795,N_1587,N_1389);
xor U8796 (N_8796,N_1818,N_1747);
nor U8797 (N_8797,N_241,N_1231);
and U8798 (N_8798,N_1386,N_1681);
or U8799 (N_8799,N_1378,N_223);
nor U8800 (N_8800,N_2887,N_3623);
nor U8801 (N_8801,N_3900,N_2095);
xnor U8802 (N_8802,N_3016,N_2050);
nand U8803 (N_8803,N_4503,N_3267);
and U8804 (N_8804,N_3085,N_3848);
or U8805 (N_8805,N_2658,N_1166);
xor U8806 (N_8806,N_973,N_2005);
or U8807 (N_8807,N_148,N_3431);
and U8808 (N_8808,N_3379,N_2301);
nand U8809 (N_8809,N_3371,N_1804);
and U8810 (N_8810,N_3581,N_4664);
or U8811 (N_8811,N_2889,N_3318);
or U8812 (N_8812,N_2572,N_2655);
nor U8813 (N_8813,N_3903,N_4260);
nor U8814 (N_8814,N_463,N_1961);
nor U8815 (N_8815,N_1042,N_2106);
or U8816 (N_8816,N_1929,N_1922);
or U8817 (N_8817,N_1112,N_3538);
nand U8818 (N_8818,N_3949,N_4278);
or U8819 (N_8819,N_1995,N_1409);
and U8820 (N_8820,N_1608,N_2295);
or U8821 (N_8821,N_477,N_749);
xor U8822 (N_8822,N_1824,N_2484);
and U8823 (N_8823,N_271,N_291);
nand U8824 (N_8824,N_4479,N_4244);
nor U8825 (N_8825,N_2320,N_1973);
or U8826 (N_8826,N_2093,N_469);
nor U8827 (N_8827,N_2926,N_1772);
nand U8828 (N_8828,N_3051,N_2507);
or U8829 (N_8829,N_1376,N_4247);
nor U8830 (N_8830,N_3224,N_984);
and U8831 (N_8831,N_4501,N_853);
nor U8832 (N_8832,N_1430,N_3729);
or U8833 (N_8833,N_3382,N_1881);
nand U8834 (N_8834,N_4119,N_2830);
and U8835 (N_8835,N_1300,N_930);
nand U8836 (N_8836,N_2776,N_1649);
nor U8837 (N_8837,N_2149,N_3693);
xor U8838 (N_8838,N_736,N_1483);
nor U8839 (N_8839,N_4844,N_1825);
nor U8840 (N_8840,N_873,N_2535);
or U8841 (N_8841,N_2315,N_807);
nor U8842 (N_8842,N_552,N_2342);
nor U8843 (N_8843,N_3584,N_2313);
xor U8844 (N_8844,N_3404,N_95);
xnor U8845 (N_8845,N_1883,N_4724);
nand U8846 (N_8846,N_1840,N_1405);
nand U8847 (N_8847,N_921,N_3712);
or U8848 (N_8848,N_4575,N_3224);
xnor U8849 (N_8849,N_14,N_3799);
nor U8850 (N_8850,N_4985,N_4283);
and U8851 (N_8851,N_2210,N_3649);
and U8852 (N_8852,N_1538,N_3811);
or U8853 (N_8853,N_3467,N_832);
or U8854 (N_8854,N_4806,N_4131);
nand U8855 (N_8855,N_3017,N_2265);
or U8856 (N_8856,N_4620,N_3206);
or U8857 (N_8857,N_1818,N_4371);
xor U8858 (N_8858,N_3990,N_1007);
xor U8859 (N_8859,N_390,N_222);
and U8860 (N_8860,N_2204,N_3152);
xnor U8861 (N_8861,N_536,N_2832);
xor U8862 (N_8862,N_2299,N_4929);
and U8863 (N_8863,N_3816,N_4262);
or U8864 (N_8864,N_4985,N_3191);
nand U8865 (N_8865,N_4163,N_4997);
or U8866 (N_8866,N_3557,N_1961);
nor U8867 (N_8867,N_1245,N_1536);
xnor U8868 (N_8868,N_3792,N_3484);
xor U8869 (N_8869,N_1983,N_1454);
and U8870 (N_8870,N_1045,N_3978);
xnor U8871 (N_8871,N_2330,N_3465);
nor U8872 (N_8872,N_1611,N_336);
nand U8873 (N_8873,N_3504,N_4200);
nor U8874 (N_8874,N_2017,N_1767);
nand U8875 (N_8875,N_2145,N_2328);
nor U8876 (N_8876,N_3375,N_2890);
nor U8877 (N_8877,N_2956,N_3194);
or U8878 (N_8878,N_4171,N_1027);
xor U8879 (N_8879,N_3002,N_4464);
nand U8880 (N_8880,N_1263,N_2430);
xor U8881 (N_8881,N_2757,N_3807);
xnor U8882 (N_8882,N_2295,N_4731);
xor U8883 (N_8883,N_2609,N_4088);
or U8884 (N_8884,N_2469,N_4708);
nand U8885 (N_8885,N_4084,N_4587);
nor U8886 (N_8886,N_554,N_4559);
and U8887 (N_8887,N_4016,N_4108);
or U8888 (N_8888,N_1714,N_4690);
or U8889 (N_8889,N_1237,N_3037);
nor U8890 (N_8890,N_464,N_3121);
nor U8891 (N_8891,N_4466,N_3496);
and U8892 (N_8892,N_3913,N_4275);
and U8893 (N_8893,N_3780,N_428);
nand U8894 (N_8894,N_1024,N_1258);
and U8895 (N_8895,N_2750,N_4266);
and U8896 (N_8896,N_941,N_302);
and U8897 (N_8897,N_919,N_1235);
nor U8898 (N_8898,N_1444,N_743);
nor U8899 (N_8899,N_3891,N_3829);
and U8900 (N_8900,N_832,N_2067);
nand U8901 (N_8901,N_1337,N_2551);
nand U8902 (N_8902,N_1177,N_994);
or U8903 (N_8903,N_3130,N_4840);
xor U8904 (N_8904,N_1565,N_3472);
and U8905 (N_8905,N_4901,N_3754);
xor U8906 (N_8906,N_3140,N_1583);
and U8907 (N_8907,N_3107,N_1214);
xor U8908 (N_8908,N_3990,N_3089);
nand U8909 (N_8909,N_1806,N_4499);
xor U8910 (N_8910,N_3086,N_2725);
nand U8911 (N_8911,N_4291,N_2513);
and U8912 (N_8912,N_4176,N_1040);
xor U8913 (N_8913,N_1732,N_2256);
xnor U8914 (N_8914,N_491,N_2719);
nor U8915 (N_8915,N_504,N_3550);
nor U8916 (N_8916,N_2156,N_2843);
and U8917 (N_8917,N_1758,N_2001);
or U8918 (N_8918,N_1646,N_4495);
xor U8919 (N_8919,N_4265,N_1933);
xor U8920 (N_8920,N_3623,N_573);
nand U8921 (N_8921,N_2155,N_1024);
and U8922 (N_8922,N_3031,N_1576);
xor U8923 (N_8923,N_892,N_1027);
nand U8924 (N_8924,N_1169,N_1246);
and U8925 (N_8925,N_3005,N_4451);
and U8926 (N_8926,N_3350,N_4187);
xnor U8927 (N_8927,N_3838,N_2226);
nand U8928 (N_8928,N_3644,N_673);
and U8929 (N_8929,N_2583,N_989);
and U8930 (N_8930,N_2403,N_1670);
and U8931 (N_8931,N_2230,N_196);
and U8932 (N_8932,N_3309,N_2471);
and U8933 (N_8933,N_1751,N_3460);
nor U8934 (N_8934,N_1722,N_826);
or U8935 (N_8935,N_76,N_1678);
or U8936 (N_8936,N_529,N_1997);
nand U8937 (N_8937,N_1419,N_2180);
xnor U8938 (N_8938,N_1246,N_4437);
xnor U8939 (N_8939,N_2692,N_2520);
nand U8940 (N_8940,N_1455,N_1879);
nand U8941 (N_8941,N_3847,N_820);
nor U8942 (N_8942,N_3123,N_3073);
nor U8943 (N_8943,N_1006,N_1231);
or U8944 (N_8944,N_577,N_3335);
or U8945 (N_8945,N_2747,N_2829);
or U8946 (N_8946,N_820,N_4139);
nand U8947 (N_8947,N_3020,N_4894);
nand U8948 (N_8948,N_4293,N_3832);
xnor U8949 (N_8949,N_3840,N_205);
nand U8950 (N_8950,N_3663,N_867);
xor U8951 (N_8951,N_3612,N_3112);
nand U8952 (N_8952,N_640,N_3088);
or U8953 (N_8953,N_4402,N_4111);
or U8954 (N_8954,N_4559,N_4726);
and U8955 (N_8955,N_393,N_4311);
nor U8956 (N_8956,N_3993,N_32);
xor U8957 (N_8957,N_1802,N_764);
nor U8958 (N_8958,N_2896,N_4950);
and U8959 (N_8959,N_912,N_2814);
xor U8960 (N_8960,N_4899,N_208);
or U8961 (N_8961,N_3447,N_3728);
nand U8962 (N_8962,N_152,N_4559);
nand U8963 (N_8963,N_2242,N_1913);
xnor U8964 (N_8964,N_4519,N_3292);
or U8965 (N_8965,N_1001,N_3373);
and U8966 (N_8966,N_951,N_973);
xnor U8967 (N_8967,N_1117,N_3897);
nand U8968 (N_8968,N_3115,N_4507);
nand U8969 (N_8969,N_1628,N_2894);
nand U8970 (N_8970,N_4077,N_2282);
and U8971 (N_8971,N_1639,N_2757);
nor U8972 (N_8972,N_4673,N_4856);
or U8973 (N_8973,N_2713,N_4491);
xor U8974 (N_8974,N_1893,N_4048);
nor U8975 (N_8975,N_2494,N_1326);
and U8976 (N_8976,N_3817,N_2505);
nand U8977 (N_8977,N_4004,N_1846);
and U8978 (N_8978,N_4313,N_324);
nand U8979 (N_8979,N_1000,N_3023);
nand U8980 (N_8980,N_1709,N_1718);
and U8981 (N_8981,N_4314,N_3142);
nor U8982 (N_8982,N_3186,N_725);
and U8983 (N_8983,N_2927,N_152);
and U8984 (N_8984,N_1269,N_4321);
nor U8985 (N_8985,N_4229,N_4237);
xor U8986 (N_8986,N_4606,N_2449);
or U8987 (N_8987,N_4795,N_3506);
nor U8988 (N_8988,N_2902,N_3142);
xor U8989 (N_8989,N_4881,N_2195);
xor U8990 (N_8990,N_4675,N_3399);
and U8991 (N_8991,N_4481,N_3169);
nand U8992 (N_8992,N_118,N_326);
nor U8993 (N_8993,N_4331,N_2202);
and U8994 (N_8994,N_3035,N_3934);
nand U8995 (N_8995,N_1013,N_1059);
or U8996 (N_8996,N_482,N_2364);
or U8997 (N_8997,N_1405,N_4170);
nand U8998 (N_8998,N_3034,N_2782);
or U8999 (N_8999,N_1730,N_585);
nand U9000 (N_9000,N_3347,N_284);
nor U9001 (N_9001,N_4920,N_4862);
nor U9002 (N_9002,N_3783,N_2663);
nor U9003 (N_9003,N_3118,N_4082);
nor U9004 (N_9004,N_3317,N_3328);
nand U9005 (N_9005,N_3140,N_2693);
or U9006 (N_9006,N_3163,N_2042);
nand U9007 (N_9007,N_674,N_4388);
xor U9008 (N_9008,N_3872,N_4607);
nand U9009 (N_9009,N_3152,N_3273);
nor U9010 (N_9010,N_3037,N_2046);
nand U9011 (N_9011,N_4117,N_3806);
nand U9012 (N_9012,N_3032,N_965);
and U9013 (N_9013,N_4837,N_2904);
or U9014 (N_9014,N_4097,N_2947);
xor U9015 (N_9015,N_2104,N_3939);
nand U9016 (N_9016,N_1205,N_1863);
xnor U9017 (N_9017,N_4449,N_1539);
and U9018 (N_9018,N_2748,N_1034);
nand U9019 (N_9019,N_1940,N_582);
and U9020 (N_9020,N_2250,N_906);
or U9021 (N_9021,N_3023,N_2605);
nand U9022 (N_9022,N_4195,N_4211);
xnor U9023 (N_9023,N_3131,N_4177);
xnor U9024 (N_9024,N_4700,N_3780);
nor U9025 (N_9025,N_4465,N_3198);
nand U9026 (N_9026,N_1422,N_689);
or U9027 (N_9027,N_778,N_951);
nor U9028 (N_9028,N_1932,N_517);
nor U9029 (N_9029,N_963,N_2560);
xnor U9030 (N_9030,N_4636,N_3323);
nand U9031 (N_9031,N_4532,N_1745);
or U9032 (N_9032,N_4637,N_77);
or U9033 (N_9033,N_3945,N_3133);
and U9034 (N_9034,N_3385,N_4480);
and U9035 (N_9035,N_3317,N_277);
or U9036 (N_9036,N_789,N_4420);
xor U9037 (N_9037,N_3124,N_1398);
or U9038 (N_9038,N_4651,N_2066);
nand U9039 (N_9039,N_733,N_2548);
or U9040 (N_9040,N_3415,N_957);
and U9041 (N_9041,N_1671,N_1358);
or U9042 (N_9042,N_3181,N_2317);
or U9043 (N_9043,N_338,N_804);
nor U9044 (N_9044,N_142,N_48);
xor U9045 (N_9045,N_106,N_1540);
nor U9046 (N_9046,N_3231,N_528);
or U9047 (N_9047,N_2453,N_1795);
xor U9048 (N_9048,N_2302,N_800);
xor U9049 (N_9049,N_1985,N_3596);
and U9050 (N_9050,N_3181,N_2323);
nand U9051 (N_9051,N_1854,N_4226);
and U9052 (N_9052,N_1037,N_1666);
nor U9053 (N_9053,N_4155,N_2246);
and U9054 (N_9054,N_3290,N_4580);
and U9055 (N_9055,N_2410,N_2577);
and U9056 (N_9056,N_3325,N_2625);
nand U9057 (N_9057,N_4212,N_3244);
or U9058 (N_9058,N_4066,N_1381);
xor U9059 (N_9059,N_3939,N_3715);
or U9060 (N_9060,N_3985,N_2971);
xnor U9061 (N_9061,N_1017,N_3131);
nand U9062 (N_9062,N_1180,N_2619);
nor U9063 (N_9063,N_1069,N_2034);
xor U9064 (N_9064,N_4622,N_4453);
or U9065 (N_9065,N_4239,N_1642);
or U9066 (N_9066,N_1826,N_4706);
or U9067 (N_9067,N_394,N_533);
nor U9068 (N_9068,N_516,N_3895);
and U9069 (N_9069,N_504,N_4000);
and U9070 (N_9070,N_2388,N_3591);
xor U9071 (N_9071,N_2279,N_2375);
nand U9072 (N_9072,N_2328,N_3688);
xor U9073 (N_9073,N_3689,N_3299);
and U9074 (N_9074,N_2603,N_1346);
and U9075 (N_9075,N_4007,N_3164);
nor U9076 (N_9076,N_2918,N_4812);
nand U9077 (N_9077,N_3585,N_4897);
xnor U9078 (N_9078,N_427,N_2546);
nand U9079 (N_9079,N_2621,N_1673);
nor U9080 (N_9080,N_4860,N_4586);
nand U9081 (N_9081,N_2596,N_1391);
nor U9082 (N_9082,N_1839,N_131);
nand U9083 (N_9083,N_2748,N_731);
nand U9084 (N_9084,N_2504,N_108);
nor U9085 (N_9085,N_913,N_1018);
and U9086 (N_9086,N_4135,N_67);
nand U9087 (N_9087,N_1179,N_4376);
or U9088 (N_9088,N_1937,N_1701);
or U9089 (N_9089,N_3482,N_296);
nand U9090 (N_9090,N_4436,N_2261);
nand U9091 (N_9091,N_4801,N_4336);
xor U9092 (N_9092,N_4977,N_1910);
and U9093 (N_9093,N_2553,N_3037);
and U9094 (N_9094,N_3122,N_4431);
or U9095 (N_9095,N_1402,N_865);
nor U9096 (N_9096,N_2844,N_998);
or U9097 (N_9097,N_4382,N_2533);
xnor U9098 (N_9098,N_4596,N_1201);
xnor U9099 (N_9099,N_3864,N_511);
or U9100 (N_9100,N_4399,N_2490);
or U9101 (N_9101,N_646,N_573);
and U9102 (N_9102,N_1665,N_1847);
xnor U9103 (N_9103,N_816,N_2662);
or U9104 (N_9104,N_4874,N_4467);
or U9105 (N_9105,N_4557,N_4004);
and U9106 (N_9106,N_3061,N_2548);
nand U9107 (N_9107,N_2927,N_1097);
xor U9108 (N_9108,N_4702,N_4092);
xnor U9109 (N_9109,N_818,N_4220);
xnor U9110 (N_9110,N_3300,N_3936);
nor U9111 (N_9111,N_4032,N_1042);
nor U9112 (N_9112,N_1209,N_2532);
xor U9113 (N_9113,N_2358,N_1428);
or U9114 (N_9114,N_3534,N_294);
nor U9115 (N_9115,N_2624,N_3836);
nor U9116 (N_9116,N_2017,N_8);
nand U9117 (N_9117,N_2630,N_321);
nor U9118 (N_9118,N_1309,N_462);
xor U9119 (N_9119,N_3894,N_2622);
xnor U9120 (N_9120,N_2930,N_2383);
nor U9121 (N_9121,N_3150,N_1734);
nor U9122 (N_9122,N_2915,N_732);
nand U9123 (N_9123,N_2475,N_1501);
xor U9124 (N_9124,N_4400,N_3595);
or U9125 (N_9125,N_2493,N_2598);
nor U9126 (N_9126,N_598,N_4623);
nand U9127 (N_9127,N_3942,N_1806);
nand U9128 (N_9128,N_2858,N_4136);
and U9129 (N_9129,N_1428,N_3763);
or U9130 (N_9130,N_4341,N_1273);
or U9131 (N_9131,N_2426,N_3585);
nor U9132 (N_9132,N_824,N_1920);
or U9133 (N_9133,N_296,N_2436);
nor U9134 (N_9134,N_2271,N_1294);
or U9135 (N_9135,N_4439,N_1591);
nand U9136 (N_9136,N_2297,N_1159);
or U9137 (N_9137,N_3175,N_2269);
or U9138 (N_9138,N_2632,N_2355);
xor U9139 (N_9139,N_4081,N_3763);
nor U9140 (N_9140,N_2928,N_2181);
and U9141 (N_9141,N_2058,N_4756);
xor U9142 (N_9142,N_4290,N_2519);
xor U9143 (N_9143,N_2379,N_2325);
xor U9144 (N_9144,N_1384,N_2342);
and U9145 (N_9145,N_2876,N_4135);
and U9146 (N_9146,N_2584,N_1943);
and U9147 (N_9147,N_770,N_3361);
xnor U9148 (N_9148,N_4225,N_2931);
nor U9149 (N_9149,N_1409,N_569);
and U9150 (N_9150,N_168,N_2081);
xor U9151 (N_9151,N_1332,N_804);
xnor U9152 (N_9152,N_1491,N_3338);
and U9153 (N_9153,N_3533,N_4612);
and U9154 (N_9154,N_1167,N_459);
and U9155 (N_9155,N_2732,N_3211);
xor U9156 (N_9156,N_3654,N_1297);
and U9157 (N_9157,N_702,N_3874);
nor U9158 (N_9158,N_768,N_3300);
nand U9159 (N_9159,N_1209,N_4702);
nand U9160 (N_9160,N_1369,N_573);
or U9161 (N_9161,N_4493,N_829);
or U9162 (N_9162,N_1975,N_578);
nor U9163 (N_9163,N_1288,N_3134);
xnor U9164 (N_9164,N_729,N_4435);
xor U9165 (N_9165,N_1922,N_285);
nand U9166 (N_9166,N_1184,N_2728);
xor U9167 (N_9167,N_3441,N_653);
xnor U9168 (N_9168,N_4818,N_2556);
and U9169 (N_9169,N_3320,N_2618);
xnor U9170 (N_9170,N_3465,N_4150);
nand U9171 (N_9171,N_4033,N_224);
and U9172 (N_9172,N_1203,N_64);
nor U9173 (N_9173,N_643,N_2452);
nor U9174 (N_9174,N_4036,N_2309);
and U9175 (N_9175,N_1768,N_147);
and U9176 (N_9176,N_984,N_888);
nor U9177 (N_9177,N_4918,N_508);
and U9178 (N_9178,N_1613,N_3962);
or U9179 (N_9179,N_660,N_658);
xnor U9180 (N_9180,N_4374,N_4032);
nor U9181 (N_9181,N_1034,N_3854);
nor U9182 (N_9182,N_783,N_1243);
nand U9183 (N_9183,N_4019,N_4116);
and U9184 (N_9184,N_858,N_2704);
and U9185 (N_9185,N_3096,N_2445);
nor U9186 (N_9186,N_786,N_4749);
nand U9187 (N_9187,N_2096,N_1142);
xor U9188 (N_9188,N_2418,N_2151);
or U9189 (N_9189,N_4029,N_1343);
and U9190 (N_9190,N_881,N_1479);
nand U9191 (N_9191,N_1281,N_3458);
or U9192 (N_9192,N_2950,N_178);
and U9193 (N_9193,N_1381,N_4240);
nand U9194 (N_9194,N_916,N_4351);
xor U9195 (N_9195,N_3317,N_1187);
and U9196 (N_9196,N_3343,N_4975);
nor U9197 (N_9197,N_4023,N_3032);
or U9198 (N_9198,N_3031,N_946);
and U9199 (N_9199,N_1587,N_1515);
xnor U9200 (N_9200,N_628,N_1584);
nand U9201 (N_9201,N_638,N_2162);
or U9202 (N_9202,N_4061,N_1536);
or U9203 (N_9203,N_2927,N_318);
nor U9204 (N_9204,N_3012,N_3521);
xor U9205 (N_9205,N_3660,N_4838);
xnor U9206 (N_9206,N_4935,N_2582);
and U9207 (N_9207,N_958,N_3992);
nand U9208 (N_9208,N_2622,N_2968);
and U9209 (N_9209,N_2596,N_2057);
xor U9210 (N_9210,N_4818,N_3815);
xnor U9211 (N_9211,N_1126,N_1989);
or U9212 (N_9212,N_1413,N_2053);
nand U9213 (N_9213,N_728,N_3960);
and U9214 (N_9214,N_4463,N_3368);
xor U9215 (N_9215,N_1635,N_3610);
xor U9216 (N_9216,N_2098,N_762);
and U9217 (N_9217,N_2154,N_510);
and U9218 (N_9218,N_1693,N_3969);
or U9219 (N_9219,N_2598,N_753);
or U9220 (N_9220,N_4741,N_1847);
nor U9221 (N_9221,N_4136,N_967);
nor U9222 (N_9222,N_4454,N_21);
xor U9223 (N_9223,N_4347,N_536);
nand U9224 (N_9224,N_3277,N_3770);
or U9225 (N_9225,N_2382,N_2695);
xor U9226 (N_9226,N_312,N_4678);
and U9227 (N_9227,N_1663,N_487);
xnor U9228 (N_9228,N_3411,N_3185);
or U9229 (N_9229,N_4842,N_3641);
nor U9230 (N_9230,N_3622,N_4619);
nor U9231 (N_9231,N_696,N_2606);
nor U9232 (N_9232,N_1203,N_1286);
xor U9233 (N_9233,N_4391,N_1926);
and U9234 (N_9234,N_4481,N_2429);
xor U9235 (N_9235,N_3218,N_3495);
nand U9236 (N_9236,N_2108,N_2278);
or U9237 (N_9237,N_4040,N_1345);
and U9238 (N_9238,N_1961,N_4645);
and U9239 (N_9239,N_3234,N_1704);
and U9240 (N_9240,N_3401,N_3998);
nand U9241 (N_9241,N_1934,N_3261);
xnor U9242 (N_9242,N_517,N_520);
nor U9243 (N_9243,N_371,N_4911);
nand U9244 (N_9244,N_4657,N_3467);
nor U9245 (N_9245,N_3146,N_3378);
xnor U9246 (N_9246,N_4911,N_2259);
nand U9247 (N_9247,N_2465,N_575);
xor U9248 (N_9248,N_3105,N_2559);
or U9249 (N_9249,N_1787,N_4660);
nor U9250 (N_9250,N_4406,N_1109);
and U9251 (N_9251,N_278,N_2704);
nand U9252 (N_9252,N_176,N_4319);
nor U9253 (N_9253,N_1632,N_98);
nor U9254 (N_9254,N_4314,N_2741);
nand U9255 (N_9255,N_4406,N_1015);
and U9256 (N_9256,N_2989,N_4167);
nor U9257 (N_9257,N_1104,N_1414);
or U9258 (N_9258,N_3200,N_912);
nand U9259 (N_9259,N_2653,N_3566);
and U9260 (N_9260,N_1640,N_1076);
or U9261 (N_9261,N_3272,N_2773);
xnor U9262 (N_9262,N_1115,N_2962);
or U9263 (N_9263,N_4652,N_920);
nand U9264 (N_9264,N_2831,N_2081);
nand U9265 (N_9265,N_2052,N_986);
or U9266 (N_9266,N_365,N_214);
or U9267 (N_9267,N_3603,N_2511);
and U9268 (N_9268,N_130,N_4670);
nand U9269 (N_9269,N_1634,N_3169);
nor U9270 (N_9270,N_4696,N_3806);
nand U9271 (N_9271,N_1132,N_1584);
xor U9272 (N_9272,N_2729,N_3604);
or U9273 (N_9273,N_1409,N_2180);
xor U9274 (N_9274,N_4019,N_829);
nand U9275 (N_9275,N_4636,N_4675);
or U9276 (N_9276,N_4397,N_1980);
or U9277 (N_9277,N_3504,N_3705);
nor U9278 (N_9278,N_4356,N_3905);
or U9279 (N_9279,N_3758,N_4028);
or U9280 (N_9280,N_3480,N_3655);
nor U9281 (N_9281,N_828,N_3409);
xnor U9282 (N_9282,N_2928,N_1879);
nand U9283 (N_9283,N_506,N_3582);
and U9284 (N_9284,N_2155,N_3507);
and U9285 (N_9285,N_1933,N_4954);
xnor U9286 (N_9286,N_2646,N_4097);
nand U9287 (N_9287,N_3178,N_3661);
nor U9288 (N_9288,N_620,N_3573);
or U9289 (N_9289,N_3519,N_3555);
or U9290 (N_9290,N_4573,N_3526);
and U9291 (N_9291,N_2082,N_3015);
nand U9292 (N_9292,N_1080,N_4287);
or U9293 (N_9293,N_4768,N_1364);
or U9294 (N_9294,N_2623,N_4232);
xnor U9295 (N_9295,N_3370,N_2565);
nand U9296 (N_9296,N_3893,N_2678);
nor U9297 (N_9297,N_1427,N_1974);
and U9298 (N_9298,N_2277,N_3383);
nor U9299 (N_9299,N_4740,N_4630);
nor U9300 (N_9300,N_1069,N_588);
nand U9301 (N_9301,N_1043,N_2248);
nor U9302 (N_9302,N_2045,N_1088);
nor U9303 (N_9303,N_4476,N_1701);
or U9304 (N_9304,N_4282,N_343);
or U9305 (N_9305,N_2960,N_4041);
xnor U9306 (N_9306,N_4268,N_4127);
nand U9307 (N_9307,N_4509,N_2631);
or U9308 (N_9308,N_3336,N_1743);
and U9309 (N_9309,N_1053,N_3174);
xor U9310 (N_9310,N_1685,N_1743);
nor U9311 (N_9311,N_1184,N_933);
nor U9312 (N_9312,N_2688,N_2565);
and U9313 (N_9313,N_2896,N_2155);
or U9314 (N_9314,N_2150,N_2836);
xor U9315 (N_9315,N_1033,N_1153);
xor U9316 (N_9316,N_1563,N_567);
or U9317 (N_9317,N_465,N_3311);
nor U9318 (N_9318,N_2,N_912);
nand U9319 (N_9319,N_3135,N_2817);
and U9320 (N_9320,N_2537,N_209);
xor U9321 (N_9321,N_3387,N_684);
nand U9322 (N_9322,N_263,N_3024);
or U9323 (N_9323,N_24,N_2392);
nand U9324 (N_9324,N_259,N_2834);
and U9325 (N_9325,N_4937,N_3920);
or U9326 (N_9326,N_1981,N_4844);
xnor U9327 (N_9327,N_2132,N_2245);
or U9328 (N_9328,N_2973,N_4);
xor U9329 (N_9329,N_4894,N_2075);
xnor U9330 (N_9330,N_4166,N_2202);
nor U9331 (N_9331,N_3394,N_1716);
and U9332 (N_9332,N_2618,N_4786);
or U9333 (N_9333,N_2577,N_2826);
xor U9334 (N_9334,N_2869,N_956);
nor U9335 (N_9335,N_4062,N_1790);
and U9336 (N_9336,N_2073,N_2858);
and U9337 (N_9337,N_1556,N_4925);
xnor U9338 (N_9338,N_180,N_4235);
nand U9339 (N_9339,N_605,N_3318);
nor U9340 (N_9340,N_3330,N_351);
nor U9341 (N_9341,N_1119,N_4202);
and U9342 (N_9342,N_590,N_3040);
nand U9343 (N_9343,N_1396,N_3421);
xnor U9344 (N_9344,N_1451,N_2475);
xor U9345 (N_9345,N_3920,N_2652);
nand U9346 (N_9346,N_4387,N_273);
xnor U9347 (N_9347,N_4463,N_2331);
or U9348 (N_9348,N_3728,N_2052);
nor U9349 (N_9349,N_4691,N_4092);
nor U9350 (N_9350,N_4843,N_1827);
xnor U9351 (N_9351,N_422,N_3007);
nor U9352 (N_9352,N_920,N_4721);
nand U9353 (N_9353,N_4456,N_2038);
xor U9354 (N_9354,N_4183,N_2270);
nor U9355 (N_9355,N_2288,N_2610);
nor U9356 (N_9356,N_3787,N_1600);
nor U9357 (N_9357,N_1175,N_2584);
or U9358 (N_9358,N_2065,N_594);
nand U9359 (N_9359,N_4633,N_4091);
nand U9360 (N_9360,N_3790,N_1368);
nand U9361 (N_9361,N_2998,N_260);
nand U9362 (N_9362,N_896,N_4053);
nand U9363 (N_9363,N_1374,N_3342);
xor U9364 (N_9364,N_3340,N_2541);
nor U9365 (N_9365,N_870,N_1065);
or U9366 (N_9366,N_1849,N_2342);
and U9367 (N_9367,N_3177,N_1119);
nor U9368 (N_9368,N_2418,N_1821);
nand U9369 (N_9369,N_1210,N_4091);
and U9370 (N_9370,N_2502,N_545);
or U9371 (N_9371,N_738,N_1031);
nor U9372 (N_9372,N_1151,N_3782);
or U9373 (N_9373,N_774,N_1456);
nor U9374 (N_9374,N_1388,N_4145);
xor U9375 (N_9375,N_4610,N_3653);
xnor U9376 (N_9376,N_571,N_3153);
nand U9377 (N_9377,N_386,N_4726);
xor U9378 (N_9378,N_4563,N_1292);
and U9379 (N_9379,N_3671,N_2713);
nand U9380 (N_9380,N_4294,N_603);
nor U9381 (N_9381,N_557,N_2011);
or U9382 (N_9382,N_2869,N_2636);
nand U9383 (N_9383,N_2175,N_642);
nor U9384 (N_9384,N_683,N_776);
nand U9385 (N_9385,N_3793,N_795);
xnor U9386 (N_9386,N_3082,N_567);
and U9387 (N_9387,N_3767,N_3850);
nand U9388 (N_9388,N_4833,N_3220);
nor U9389 (N_9389,N_2811,N_3065);
and U9390 (N_9390,N_2503,N_710);
and U9391 (N_9391,N_1435,N_1143);
nand U9392 (N_9392,N_3152,N_4503);
xnor U9393 (N_9393,N_939,N_4573);
nor U9394 (N_9394,N_4878,N_2800);
xnor U9395 (N_9395,N_3035,N_698);
xor U9396 (N_9396,N_2744,N_3576);
xnor U9397 (N_9397,N_2798,N_184);
and U9398 (N_9398,N_2762,N_2729);
nor U9399 (N_9399,N_2964,N_2269);
nor U9400 (N_9400,N_3287,N_277);
nor U9401 (N_9401,N_2976,N_2225);
nand U9402 (N_9402,N_1493,N_2572);
or U9403 (N_9403,N_4281,N_2367);
or U9404 (N_9404,N_2498,N_1137);
xor U9405 (N_9405,N_1821,N_4855);
nand U9406 (N_9406,N_2876,N_1489);
or U9407 (N_9407,N_4062,N_3284);
nand U9408 (N_9408,N_1621,N_320);
nand U9409 (N_9409,N_3320,N_1967);
nand U9410 (N_9410,N_3525,N_602);
or U9411 (N_9411,N_3895,N_750);
or U9412 (N_9412,N_2773,N_378);
nand U9413 (N_9413,N_329,N_1402);
nand U9414 (N_9414,N_3716,N_2756);
nand U9415 (N_9415,N_2763,N_3028);
nand U9416 (N_9416,N_4714,N_4077);
or U9417 (N_9417,N_1204,N_4146);
xnor U9418 (N_9418,N_2082,N_3187);
and U9419 (N_9419,N_2136,N_4504);
nand U9420 (N_9420,N_4520,N_259);
and U9421 (N_9421,N_2371,N_462);
nor U9422 (N_9422,N_2808,N_1214);
nor U9423 (N_9423,N_2759,N_4981);
nand U9424 (N_9424,N_678,N_2945);
nand U9425 (N_9425,N_741,N_1883);
nor U9426 (N_9426,N_2693,N_2734);
or U9427 (N_9427,N_137,N_2068);
or U9428 (N_9428,N_836,N_1672);
or U9429 (N_9429,N_2555,N_389);
nor U9430 (N_9430,N_2725,N_4072);
nor U9431 (N_9431,N_2419,N_2841);
and U9432 (N_9432,N_3593,N_453);
nand U9433 (N_9433,N_4180,N_4594);
or U9434 (N_9434,N_3835,N_2063);
nand U9435 (N_9435,N_2118,N_970);
and U9436 (N_9436,N_1206,N_409);
nand U9437 (N_9437,N_2741,N_4356);
and U9438 (N_9438,N_4046,N_3963);
nor U9439 (N_9439,N_2130,N_629);
nand U9440 (N_9440,N_1644,N_2030);
nor U9441 (N_9441,N_4447,N_4911);
or U9442 (N_9442,N_4708,N_3970);
xor U9443 (N_9443,N_4294,N_2622);
xnor U9444 (N_9444,N_1378,N_1335);
and U9445 (N_9445,N_4551,N_4310);
nand U9446 (N_9446,N_1104,N_681);
nor U9447 (N_9447,N_949,N_103);
nor U9448 (N_9448,N_1437,N_1039);
nand U9449 (N_9449,N_243,N_113);
xor U9450 (N_9450,N_2140,N_50);
nand U9451 (N_9451,N_1369,N_2936);
nor U9452 (N_9452,N_1130,N_2136);
or U9453 (N_9453,N_4390,N_951);
and U9454 (N_9454,N_510,N_2412);
nand U9455 (N_9455,N_75,N_1239);
xor U9456 (N_9456,N_999,N_3396);
and U9457 (N_9457,N_4944,N_3165);
xor U9458 (N_9458,N_250,N_2884);
xor U9459 (N_9459,N_3189,N_4572);
and U9460 (N_9460,N_3138,N_3090);
or U9461 (N_9461,N_3533,N_2516);
or U9462 (N_9462,N_4213,N_3724);
or U9463 (N_9463,N_1900,N_4542);
nand U9464 (N_9464,N_1035,N_1482);
and U9465 (N_9465,N_512,N_2486);
xnor U9466 (N_9466,N_3914,N_132);
and U9467 (N_9467,N_3849,N_449);
xor U9468 (N_9468,N_4373,N_1759);
and U9469 (N_9469,N_2288,N_1141);
nand U9470 (N_9470,N_2774,N_2124);
and U9471 (N_9471,N_1098,N_3646);
and U9472 (N_9472,N_2835,N_3628);
nor U9473 (N_9473,N_1738,N_4280);
xor U9474 (N_9474,N_3648,N_124);
or U9475 (N_9475,N_716,N_1324);
nand U9476 (N_9476,N_861,N_3289);
nor U9477 (N_9477,N_4936,N_4325);
nor U9478 (N_9478,N_461,N_3560);
nor U9479 (N_9479,N_4919,N_2751);
or U9480 (N_9480,N_1469,N_2928);
nand U9481 (N_9481,N_1837,N_4735);
xnor U9482 (N_9482,N_4942,N_807);
nor U9483 (N_9483,N_3086,N_1135);
nand U9484 (N_9484,N_4233,N_2436);
xor U9485 (N_9485,N_4,N_1968);
or U9486 (N_9486,N_3082,N_3019);
nand U9487 (N_9487,N_1700,N_3801);
nor U9488 (N_9488,N_872,N_3323);
or U9489 (N_9489,N_193,N_2380);
xor U9490 (N_9490,N_818,N_3820);
nand U9491 (N_9491,N_2292,N_4585);
and U9492 (N_9492,N_2388,N_4492);
nor U9493 (N_9493,N_2216,N_4767);
and U9494 (N_9494,N_2704,N_2798);
or U9495 (N_9495,N_2836,N_1702);
nand U9496 (N_9496,N_3718,N_3365);
xnor U9497 (N_9497,N_3655,N_1651);
and U9498 (N_9498,N_1183,N_3469);
and U9499 (N_9499,N_3989,N_3185);
nand U9500 (N_9500,N_4697,N_3188);
nor U9501 (N_9501,N_2242,N_3511);
or U9502 (N_9502,N_3821,N_1500);
nor U9503 (N_9503,N_3478,N_2820);
nor U9504 (N_9504,N_667,N_1745);
xor U9505 (N_9505,N_882,N_4781);
nor U9506 (N_9506,N_8,N_3836);
xnor U9507 (N_9507,N_4730,N_4209);
and U9508 (N_9508,N_3659,N_4693);
and U9509 (N_9509,N_3457,N_401);
xnor U9510 (N_9510,N_2403,N_2185);
and U9511 (N_9511,N_631,N_3730);
nor U9512 (N_9512,N_2923,N_2201);
or U9513 (N_9513,N_1321,N_2285);
and U9514 (N_9514,N_169,N_4991);
nor U9515 (N_9515,N_4022,N_783);
nand U9516 (N_9516,N_1242,N_3371);
or U9517 (N_9517,N_252,N_4578);
and U9518 (N_9518,N_2257,N_3348);
nor U9519 (N_9519,N_109,N_4185);
nand U9520 (N_9520,N_2901,N_4104);
or U9521 (N_9521,N_4052,N_4995);
nor U9522 (N_9522,N_1949,N_4456);
nand U9523 (N_9523,N_2257,N_2207);
or U9524 (N_9524,N_1229,N_4850);
xnor U9525 (N_9525,N_510,N_3464);
or U9526 (N_9526,N_2698,N_4994);
and U9527 (N_9527,N_364,N_3302);
nand U9528 (N_9528,N_2263,N_3409);
or U9529 (N_9529,N_1254,N_563);
or U9530 (N_9530,N_3792,N_2526);
xnor U9531 (N_9531,N_4682,N_1239);
or U9532 (N_9532,N_481,N_4245);
and U9533 (N_9533,N_1790,N_2258);
or U9534 (N_9534,N_791,N_3947);
or U9535 (N_9535,N_808,N_83);
and U9536 (N_9536,N_913,N_3157);
or U9537 (N_9537,N_2696,N_1551);
nor U9538 (N_9538,N_3035,N_3468);
nor U9539 (N_9539,N_2345,N_573);
xor U9540 (N_9540,N_1865,N_1834);
or U9541 (N_9541,N_4545,N_3087);
nand U9542 (N_9542,N_67,N_1227);
xnor U9543 (N_9543,N_4842,N_3824);
nor U9544 (N_9544,N_3644,N_2997);
nand U9545 (N_9545,N_4169,N_4697);
nor U9546 (N_9546,N_4150,N_1393);
nand U9547 (N_9547,N_3952,N_4763);
and U9548 (N_9548,N_4367,N_4453);
nand U9549 (N_9549,N_2181,N_2463);
nor U9550 (N_9550,N_4938,N_2350);
or U9551 (N_9551,N_3123,N_1675);
nand U9552 (N_9552,N_2189,N_1296);
nor U9553 (N_9553,N_2375,N_4474);
nor U9554 (N_9554,N_3770,N_4112);
and U9555 (N_9555,N_606,N_4886);
nand U9556 (N_9556,N_1733,N_2621);
xor U9557 (N_9557,N_505,N_4283);
nor U9558 (N_9558,N_3095,N_3785);
nor U9559 (N_9559,N_4872,N_2035);
nor U9560 (N_9560,N_396,N_4316);
xor U9561 (N_9561,N_154,N_4900);
and U9562 (N_9562,N_1693,N_4559);
and U9563 (N_9563,N_4685,N_3395);
or U9564 (N_9564,N_3728,N_856);
and U9565 (N_9565,N_3433,N_4585);
xor U9566 (N_9566,N_3318,N_1787);
and U9567 (N_9567,N_1525,N_3591);
nor U9568 (N_9568,N_3090,N_1227);
xnor U9569 (N_9569,N_4216,N_4931);
nor U9570 (N_9570,N_499,N_2258);
and U9571 (N_9571,N_1874,N_2950);
nand U9572 (N_9572,N_2295,N_920);
or U9573 (N_9573,N_3225,N_3665);
xnor U9574 (N_9574,N_1139,N_117);
or U9575 (N_9575,N_3589,N_3817);
nand U9576 (N_9576,N_3920,N_137);
nand U9577 (N_9577,N_4062,N_319);
nor U9578 (N_9578,N_562,N_982);
or U9579 (N_9579,N_1994,N_4995);
or U9580 (N_9580,N_4231,N_1428);
xnor U9581 (N_9581,N_849,N_2163);
nor U9582 (N_9582,N_3329,N_3131);
or U9583 (N_9583,N_3651,N_3856);
nor U9584 (N_9584,N_4594,N_4094);
or U9585 (N_9585,N_3623,N_2181);
xnor U9586 (N_9586,N_4278,N_339);
and U9587 (N_9587,N_3719,N_4017);
nand U9588 (N_9588,N_3159,N_1837);
nand U9589 (N_9589,N_3881,N_3612);
xnor U9590 (N_9590,N_3517,N_2489);
or U9591 (N_9591,N_1108,N_1876);
nor U9592 (N_9592,N_3229,N_1267);
nand U9593 (N_9593,N_1941,N_3344);
and U9594 (N_9594,N_4403,N_4228);
or U9595 (N_9595,N_1392,N_3304);
nor U9596 (N_9596,N_1794,N_4835);
and U9597 (N_9597,N_4792,N_2216);
nor U9598 (N_9598,N_2938,N_629);
xnor U9599 (N_9599,N_3219,N_4595);
xor U9600 (N_9600,N_413,N_4634);
nand U9601 (N_9601,N_806,N_887);
nor U9602 (N_9602,N_3464,N_1156);
or U9603 (N_9603,N_2656,N_740);
and U9604 (N_9604,N_2771,N_2242);
nand U9605 (N_9605,N_2979,N_577);
nand U9606 (N_9606,N_9,N_238);
nor U9607 (N_9607,N_4477,N_4758);
nor U9608 (N_9608,N_1300,N_3921);
or U9609 (N_9609,N_507,N_2646);
nor U9610 (N_9610,N_4702,N_4065);
nand U9611 (N_9611,N_481,N_2099);
and U9612 (N_9612,N_2903,N_807);
or U9613 (N_9613,N_4972,N_3217);
or U9614 (N_9614,N_3912,N_4060);
and U9615 (N_9615,N_1565,N_4527);
nand U9616 (N_9616,N_2542,N_474);
and U9617 (N_9617,N_134,N_3285);
nand U9618 (N_9618,N_1200,N_1577);
and U9619 (N_9619,N_542,N_3549);
or U9620 (N_9620,N_897,N_2749);
nor U9621 (N_9621,N_2904,N_3772);
nor U9622 (N_9622,N_1455,N_518);
and U9623 (N_9623,N_3336,N_3365);
or U9624 (N_9624,N_3606,N_4532);
and U9625 (N_9625,N_1942,N_1613);
or U9626 (N_9626,N_926,N_4838);
and U9627 (N_9627,N_2569,N_838);
nor U9628 (N_9628,N_4830,N_1617);
and U9629 (N_9629,N_3288,N_2564);
nand U9630 (N_9630,N_152,N_1905);
and U9631 (N_9631,N_2086,N_831);
nor U9632 (N_9632,N_3676,N_2120);
xor U9633 (N_9633,N_3284,N_3373);
nor U9634 (N_9634,N_2927,N_3085);
xnor U9635 (N_9635,N_3772,N_3666);
and U9636 (N_9636,N_2578,N_3631);
nor U9637 (N_9637,N_3762,N_3838);
xnor U9638 (N_9638,N_3553,N_3699);
or U9639 (N_9639,N_1450,N_4912);
nor U9640 (N_9640,N_3717,N_3433);
and U9641 (N_9641,N_4362,N_3870);
and U9642 (N_9642,N_2924,N_1809);
nand U9643 (N_9643,N_1613,N_4029);
xor U9644 (N_9644,N_1149,N_63);
nand U9645 (N_9645,N_634,N_2740);
nand U9646 (N_9646,N_1946,N_2013);
nor U9647 (N_9647,N_394,N_3637);
nand U9648 (N_9648,N_634,N_4558);
xnor U9649 (N_9649,N_1910,N_1775);
nand U9650 (N_9650,N_2408,N_3339);
nand U9651 (N_9651,N_3138,N_3019);
and U9652 (N_9652,N_3342,N_2865);
and U9653 (N_9653,N_4825,N_3457);
nand U9654 (N_9654,N_4536,N_279);
nand U9655 (N_9655,N_4051,N_2252);
nor U9656 (N_9656,N_4474,N_187);
xor U9657 (N_9657,N_1432,N_2331);
nor U9658 (N_9658,N_2042,N_2527);
nand U9659 (N_9659,N_3032,N_4575);
or U9660 (N_9660,N_2768,N_2273);
nand U9661 (N_9661,N_4628,N_3764);
or U9662 (N_9662,N_1294,N_3990);
or U9663 (N_9663,N_352,N_1870);
xor U9664 (N_9664,N_3707,N_1693);
xor U9665 (N_9665,N_3404,N_4173);
and U9666 (N_9666,N_4566,N_3544);
xor U9667 (N_9667,N_3054,N_1165);
or U9668 (N_9668,N_4450,N_3445);
nand U9669 (N_9669,N_4791,N_210);
nor U9670 (N_9670,N_4661,N_2193);
or U9671 (N_9671,N_2052,N_2672);
xor U9672 (N_9672,N_4855,N_1309);
nor U9673 (N_9673,N_287,N_2678);
xnor U9674 (N_9674,N_1266,N_497);
and U9675 (N_9675,N_3149,N_3902);
or U9676 (N_9676,N_2079,N_4451);
or U9677 (N_9677,N_2706,N_3020);
nand U9678 (N_9678,N_2662,N_3138);
nand U9679 (N_9679,N_1689,N_3802);
nor U9680 (N_9680,N_4952,N_2093);
xor U9681 (N_9681,N_508,N_2134);
and U9682 (N_9682,N_3277,N_4239);
nand U9683 (N_9683,N_273,N_1654);
or U9684 (N_9684,N_1652,N_3896);
nor U9685 (N_9685,N_4551,N_3642);
and U9686 (N_9686,N_1431,N_966);
nor U9687 (N_9687,N_3887,N_3172);
nor U9688 (N_9688,N_584,N_4928);
or U9689 (N_9689,N_2293,N_101);
xnor U9690 (N_9690,N_4820,N_2045);
xnor U9691 (N_9691,N_3138,N_3330);
xnor U9692 (N_9692,N_4752,N_2994);
or U9693 (N_9693,N_1333,N_2575);
xor U9694 (N_9694,N_743,N_125);
xnor U9695 (N_9695,N_1219,N_4680);
xnor U9696 (N_9696,N_2296,N_1058);
nor U9697 (N_9697,N_74,N_3717);
nand U9698 (N_9698,N_3427,N_3835);
nand U9699 (N_9699,N_4771,N_4671);
and U9700 (N_9700,N_2817,N_368);
and U9701 (N_9701,N_1696,N_4109);
and U9702 (N_9702,N_3391,N_3093);
and U9703 (N_9703,N_3534,N_1197);
or U9704 (N_9704,N_1513,N_3756);
nand U9705 (N_9705,N_3403,N_4362);
nor U9706 (N_9706,N_807,N_1343);
nor U9707 (N_9707,N_4200,N_2283);
xnor U9708 (N_9708,N_170,N_3080);
xnor U9709 (N_9709,N_2601,N_2981);
nand U9710 (N_9710,N_1968,N_1346);
xnor U9711 (N_9711,N_3542,N_3295);
or U9712 (N_9712,N_1596,N_608);
xnor U9713 (N_9713,N_2947,N_1935);
or U9714 (N_9714,N_355,N_3328);
nand U9715 (N_9715,N_541,N_1872);
and U9716 (N_9716,N_2746,N_3321);
nor U9717 (N_9717,N_3428,N_1979);
xor U9718 (N_9718,N_2471,N_2034);
xor U9719 (N_9719,N_1669,N_4971);
or U9720 (N_9720,N_272,N_2042);
and U9721 (N_9721,N_2835,N_4749);
and U9722 (N_9722,N_4546,N_2367);
or U9723 (N_9723,N_2526,N_2047);
nor U9724 (N_9724,N_1195,N_198);
or U9725 (N_9725,N_894,N_2427);
or U9726 (N_9726,N_3089,N_4157);
or U9727 (N_9727,N_4642,N_4061);
or U9728 (N_9728,N_486,N_589);
nand U9729 (N_9729,N_1220,N_2501);
nor U9730 (N_9730,N_91,N_2977);
nor U9731 (N_9731,N_2267,N_928);
nand U9732 (N_9732,N_2386,N_30);
xor U9733 (N_9733,N_3360,N_3815);
nor U9734 (N_9734,N_844,N_2865);
nor U9735 (N_9735,N_2909,N_3344);
nand U9736 (N_9736,N_2444,N_1460);
xor U9737 (N_9737,N_3631,N_4733);
and U9738 (N_9738,N_2316,N_1574);
nand U9739 (N_9739,N_795,N_4003);
or U9740 (N_9740,N_3530,N_1746);
nor U9741 (N_9741,N_1382,N_619);
xnor U9742 (N_9742,N_2844,N_3395);
and U9743 (N_9743,N_4339,N_1429);
or U9744 (N_9744,N_4596,N_1115);
nand U9745 (N_9745,N_4879,N_1929);
nor U9746 (N_9746,N_1592,N_851);
nor U9747 (N_9747,N_3911,N_3330);
and U9748 (N_9748,N_1887,N_2118);
nor U9749 (N_9749,N_2131,N_449);
and U9750 (N_9750,N_1525,N_4435);
and U9751 (N_9751,N_3476,N_395);
nor U9752 (N_9752,N_3887,N_2074);
and U9753 (N_9753,N_4712,N_2735);
nand U9754 (N_9754,N_4713,N_4585);
nor U9755 (N_9755,N_945,N_206);
or U9756 (N_9756,N_2849,N_141);
nand U9757 (N_9757,N_1641,N_1635);
xor U9758 (N_9758,N_942,N_615);
nor U9759 (N_9759,N_3728,N_2088);
nor U9760 (N_9760,N_3449,N_1943);
nor U9761 (N_9761,N_858,N_1589);
nand U9762 (N_9762,N_1391,N_2178);
nor U9763 (N_9763,N_2015,N_1029);
nor U9764 (N_9764,N_579,N_4176);
or U9765 (N_9765,N_242,N_3246);
xnor U9766 (N_9766,N_2054,N_1457);
or U9767 (N_9767,N_2991,N_1875);
nor U9768 (N_9768,N_2916,N_4777);
or U9769 (N_9769,N_132,N_1955);
nand U9770 (N_9770,N_1067,N_3059);
nor U9771 (N_9771,N_4173,N_4968);
xnor U9772 (N_9772,N_426,N_4305);
or U9773 (N_9773,N_94,N_1902);
xnor U9774 (N_9774,N_4154,N_1233);
nor U9775 (N_9775,N_986,N_4634);
nand U9776 (N_9776,N_2422,N_3240);
nand U9777 (N_9777,N_4695,N_1605);
or U9778 (N_9778,N_4441,N_4091);
and U9779 (N_9779,N_4406,N_703);
nor U9780 (N_9780,N_3330,N_318);
nor U9781 (N_9781,N_2435,N_3534);
nand U9782 (N_9782,N_1283,N_117);
nor U9783 (N_9783,N_4436,N_1305);
or U9784 (N_9784,N_1179,N_2329);
and U9785 (N_9785,N_2025,N_3977);
nor U9786 (N_9786,N_4362,N_1581);
nor U9787 (N_9787,N_4157,N_3460);
xnor U9788 (N_9788,N_11,N_2142);
and U9789 (N_9789,N_2427,N_952);
and U9790 (N_9790,N_2548,N_4594);
and U9791 (N_9791,N_2131,N_3413);
nor U9792 (N_9792,N_4566,N_4347);
nor U9793 (N_9793,N_3502,N_4197);
xor U9794 (N_9794,N_1973,N_3864);
nand U9795 (N_9795,N_3116,N_4346);
nor U9796 (N_9796,N_2406,N_2607);
nor U9797 (N_9797,N_2327,N_949);
nor U9798 (N_9798,N_4421,N_1630);
nor U9799 (N_9799,N_846,N_4049);
nor U9800 (N_9800,N_4990,N_3038);
xor U9801 (N_9801,N_925,N_956);
or U9802 (N_9802,N_730,N_2668);
nand U9803 (N_9803,N_3678,N_4415);
nor U9804 (N_9804,N_2394,N_3086);
or U9805 (N_9805,N_2864,N_4449);
xor U9806 (N_9806,N_962,N_4100);
nand U9807 (N_9807,N_1927,N_292);
and U9808 (N_9808,N_1303,N_2163);
nand U9809 (N_9809,N_560,N_2662);
and U9810 (N_9810,N_2659,N_2942);
or U9811 (N_9811,N_3308,N_3394);
nor U9812 (N_9812,N_4388,N_1612);
and U9813 (N_9813,N_4075,N_187);
or U9814 (N_9814,N_3410,N_4664);
nor U9815 (N_9815,N_4870,N_229);
or U9816 (N_9816,N_4604,N_459);
xnor U9817 (N_9817,N_1624,N_591);
nor U9818 (N_9818,N_180,N_2712);
and U9819 (N_9819,N_986,N_14);
nand U9820 (N_9820,N_818,N_2949);
and U9821 (N_9821,N_2881,N_897);
nor U9822 (N_9822,N_2405,N_3188);
xnor U9823 (N_9823,N_779,N_233);
and U9824 (N_9824,N_1606,N_3683);
or U9825 (N_9825,N_4843,N_77);
xnor U9826 (N_9826,N_4510,N_965);
or U9827 (N_9827,N_1771,N_364);
nand U9828 (N_9828,N_1983,N_1661);
nand U9829 (N_9829,N_2564,N_2430);
xor U9830 (N_9830,N_1720,N_2402);
nand U9831 (N_9831,N_2193,N_1199);
nand U9832 (N_9832,N_4258,N_3903);
or U9833 (N_9833,N_2898,N_841);
or U9834 (N_9834,N_520,N_130);
and U9835 (N_9835,N_2073,N_2783);
nand U9836 (N_9836,N_491,N_4329);
nor U9837 (N_9837,N_1849,N_937);
nor U9838 (N_9838,N_1297,N_1081);
xor U9839 (N_9839,N_625,N_1531);
nand U9840 (N_9840,N_2247,N_2867);
and U9841 (N_9841,N_647,N_4297);
nor U9842 (N_9842,N_3544,N_983);
and U9843 (N_9843,N_236,N_2009);
nand U9844 (N_9844,N_3314,N_2008);
nand U9845 (N_9845,N_4207,N_2604);
xor U9846 (N_9846,N_3511,N_2184);
or U9847 (N_9847,N_417,N_1213);
xnor U9848 (N_9848,N_4517,N_2793);
xor U9849 (N_9849,N_1234,N_513);
or U9850 (N_9850,N_4047,N_3660);
nor U9851 (N_9851,N_134,N_1566);
or U9852 (N_9852,N_1908,N_873);
nand U9853 (N_9853,N_1740,N_355);
nor U9854 (N_9854,N_2935,N_3246);
xnor U9855 (N_9855,N_3152,N_148);
and U9856 (N_9856,N_4677,N_1877);
and U9857 (N_9857,N_4037,N_4342);
nand U9858 (N_9858,N_74,N_2947);
and U9859 (N_9859,N_3554,N_1087);
xnor U9860 (N_9860,N_2978,N_4400);
xnor U9861 (N_9861,N_4920,N_1162);
xor U9862 (N_9862,N_1659,N_2060);
nor U9863 (N_9863,N_1692,N_4874);
or U9864 (N_9864,N_4316,N_3494);
or U9865 (N_9865,N_2012,N_1316);
xor U9866 (N_9866,N_4999,N_5);
nand U9867 (N_9867,N_2074,N_864);
or U9868 (N_9868,N_3301,N_3732);
nand U9869 (N_9869,N_2386,N_2575);
nor U9870 (N_9870,N_4575,N_1288);
or U9871 (N_9871,N_1520,N_4221);
xnor U9872 (N_9872,N_2575,N_481);
or U9873 (N_9873,N_2565,N_885);
nand U9874 (N_9874,N_2092,N_4886);
nor U9875 (N_9875,N_2495,N_2477);
xor U9876 (N_9876,N_711,N_2795);
xnor U9877 (N_9877,N_4686,N_1837);
or U9878 (N_9878,N_8,N_569);
nor U9879 (N_9879,N_2927,N_4025);
nand U9880 (N_9880,N_2416,N_3126);
nor U9881 (N_9881,N_4121,N_2215);
or U9882 (N_9882,N_3153,N_1617);
and U9883 (N_9883,N_2666,N_2091);
xnor U9884 (N_9884,N_3070,N_4801);
xor U9885 (N_9885,N_3533,N_1453);
or U9886 (N_9886,N_4817,N_3280);
xnor U9887 (N_9887,N_268,N_158);
and U9888 (N_9888,N_4831,N_3643);
or U9889 (N_9889,N_1624,N_321);
xnor U9890 (N_9890,N_695,N_4995);
and U9891 (N_9891,N_1040,N_3565);
and U9892 (N_9892,N_3192,N_4075);
xnor U9893 (N_9893,N_3284,N_3515);
nand U9894 (N_9894,N_334,N_2683);
xor U9895 (N_9895,N_629,N_3700);
nor U9896 (N_9896,N_2219,N_4476);
nor U9897 (N_9897,N_367,N_4506);
nor U9898 (N_9898,N_3297,N_2722);
or U9899 (N_9899,N_4825,N_4368);
and U9900 (N_9900,N_1531,N_2269);
nor U9901 (N_9901,N_269,N_1997);
nor U9902 (N_9902,N_3245,N_1614);
xor U9903 (N_9903,N_1896,N_4282);
and U9904 (N_9904,N_4320,N_4570);
nand U9905 (N_9905,N_1933,N_528);
and U9906 (N_9906,N_2300,N_3362);
nand U9907 (N_9907,N_3551,N_1316);
xnor U9908 (N_9908,N_4242,N_2030);
and U9909 (N_9909,N_4718,N_4734);
nand U9910 (N_9910,N_196,N_2122);
nor U9911 (N_9911,N_940,N_573);
or U9912 (N_9912,N_1970,N_1058);
and U9913 (N_9913,N_4678,N_3743);
nand U9914 (N_9914,N_4457,N_471);
nand U9915 (N_9915,N_281,N_1045);
and U9916 (N_9916,N_2881,N_3997);
nand U9917 (N_9917,N_978,N_4424);
nor U9918 (N_9918,N_4644,N_1327);
nand U9919 (N_9919,N_2174,N_4223);
xor U9920 (N_9920,N_2549,N_2858);
nor U9921 (N_9921,N_1513,N_4664);
and U9922 (N_9922,N_3371,N_4539);
or U9923 (N_9923,N_4096,N_3067);
xor U9924 (N_9924,N_603,N_4627);
nand U9925 (N_9925,N_376,N_1494);
nor U9926 (N_9926,N_4169,N_4800);
xnor U9927 (N_9927,N_1640,N_3181);
nand U9928 (N_9928,N_2886,N_4099);
nand U9929 (N_9929,N_1254,N_783);
nor U9930 (N_9930,N_4524,N_4648);
xor U9931 (N_9931,N_4421,N_2385);
nor U9932 (N_9932,N_4075,N_4497);
xnor U9933 (N_9933,N_1061,N_4696);
and U9934 (N_9934,N_602,N_1022);
nor U9935 (N_9935,N_288,N_4259);
nand U9936 (N_9936,N_536,N_178);
nor U9937 (N_9937,N_1008,N_3531);
xor U9938 (N_9938,N_692,N_1143);
nand U9939 (N_9939,N_2369,N_4612);
or U9940 (N_9940,N_3882,N_4983);
or U9941 (N_9941,N_2515,N_760);
or U9942 (N_9942,N_2803,N_4696);
nor U9943 (N_9943,N_1620,N_1226);
and U9944 (N_9944,N_1467,N_2606);
xnor U9945 (N_9945,N_2772,N_3073);
xor U9946 (N_9946,N_1221,N_2827);
nor U9947 (N_9947,N_1255,N_341);
xnor U9948 (N_9948,N_1457,N_1298);
nor U9949 (N_9949,N_1660,N_2709);
nand U9950 (N_9950,N_3018,N_2879);
nor U9951 (N_9951,N_3050,N_1558);
xor U9952 (N_9952,N_1584,N_4023);
and U9953 (N_9953,N_763,N_4539);
and U9954 (N_9954,N_4016,N_633);
and U9955 (N_9955,N_638,N_932);
and U9956 (N_9956,N_1817,N_2221);
xor U9957 (N_9957,N_347,N_3904);
nor U9958 (N_9958,N_2672,N_3201);
nor U9959 (N_9959,N_4555,N_4481);
xnor U9960 (N_9960,N_1128,N_3593);
and U9961 (N_9961,N_2805,N_2828);
and U9962 (N_9962,N_3475,N_1523);
xnor U9963 (N_9963,N_3045,N_336);
nor U9964 (N_9964,N_2292,N_3327);
xnor U9965 (N_9965,N_1382,N_427);
and U9966 (N_9966,N_1919,N_2551);
or U9967 (N_9967,N_1253,N_3231);
nand U9968 (N_9968,N_525,N_3932);
nand U9969 (N_9969,N_885,N_2291);
nand U9970 (N_9970,N_986,N_3637);
xor U9971 (N_9971,N_1306,N_4926);
nand U9972 (N_9972,N_2801,N_1210);
or U9973 (N_9973,N_4553,N_4155);
or U9974 (N_9974,N_2962,N_2883);
nand U9975 (N_9975,N_3362,N_3991);
xnor U9976 (N_9976,N_2925,N_1130);
nor U9977 (N_9977,N_1273,N_1246);
and U9978 (N_9978,N_1197,N_3457);
xnor U9979 (N_9979,N_2801,N_1516);
xnor U9980 (N_9980,N_1386,N_1660);
and U9981 (N_9981,N_731,N_4204);
and U9982 (N_9982,N_3165,N_4301);
and U9983 (N_9983,N_1869,N_1745);
nor U9984 (N_9984,N_2026,N_4364);
xor U9985 (N_9985,N_2965,N_3856);
or U9986 (N_9986,N_566,N_1100);
nand U9987 (N_9987,N_871,N_1080);
nand U9988 (N_9988,N_618,N_1893);
and U9989 (N_9989,N_4560,N_3586);
nand U9990 (N_9990,N_4205,N_4834);
and U9991 (N_9991,N_1760,N_740);
nor U9992 (N_9992,N_1014,N_3607);
or U9993 (N_9993,N_613,N_1164);
nor U9994 (N_9994,N_4322,N_3884);
and U9995 (N_9995,N_3633,N_2965);
or U9996 (N_9996,N_3932,N_2650);
or U9997 (N_9997,N_2970,N_2314);
and U9998 (N_9998,N_1143,N_4945);
or U9999 (N_9999,N_4595,N_2525);
nor U10000 (N_10000,N_5339,N_6893);
and U10001 (N_10001,N_5448,N_7796);
xor U10002 (N_10002,N_9261,N_9019);
or U10003 (N_10003,N_7914,N_9571);
and U10004 (N_10004,N_7049,N_7157);
and U10005 (N_10005,N_6082,N_8389);
or U10006 (N_10006,N_9493,N_5771);
or U10007 (N_10007,N_8541,N_7865);
xnor U10008 (N_10008,N_9271,N_6738);
nor U10009 (N_10009,N_8551,N_6721);
or U10010 (N_10010,N_6276,N_5981);
and U10011 (N_10011,N_5127,N_8979);
nor U10012 (N_10012,N_7687,N_6417);
or U10013 (N_10013,N_7283,N_8303);
nand U10014 (N_10014,N_5973,N_9276);
nand U10015 (N_10015,N_6023,N_6752);
and U10016 (N_10016,N_7192,N_8639);
or U10017 (N_10017,N_9086,N_7316);
xor U10018 (N_10018,N_6411,N_8894);
nor U10019 (N_10019,N_9504,N_8549);
and U10020 (N_10020,N_6537,N_9673);
nor U10021 (N_10021,N_9329,N_8466);
and U10022 (N_10022,N_6008,N_8161);
and U10023 (N_10023,N_8497,N_9353);
and U10024 (N_10024,N_7949,N_9847);
xnor U10025 (N_10025,N_6891,N_5547);
and U10026 (N_10026,N_9422,N_6274);
xnor U10027 (N_10027,N_8873,N_5883);
nor U10028 (N_10028,N_9802,N_6763);
or U10029 (N_10029,N_9318,N_9440);
nor U10030 (N_10030,N_5685,N_9899);
and U10031 (N_10031,N_9039,N_7263);
nor U10032 (N_10032,N_5637,N_8495);
nor U10033 (N_10033,N_8626,N_7787);
and U10034 (N_10034,N_7030,N_7414);
nand U10035 (N_10035,N_6283,N_8859);
nor U10036 (N_10036,N_9354,N_9822);
and U10037 (N_10037,N_5316,N_7760);
and U10038 (N_10038,N_9020,N_9588);
nor U10039 (N_10039,N_9550,N_5922);
and U10040 (N_10040,N_6733,N_9264);
nor U10041 (N_10041,N_5134,N_9911);
and U10042 (N_10042,N_5331,N_6527);
nand U10043 (N_10043,N_8785,N_6977);
or U10044 (N_10044,N_7714,N_5359);
nor U10045 (N_10045,N_8328,N_9249);
and U10046 (N_10046,N_8183,N_6967);
xor U10047 (N_10047,N_5944,N_6884);
or U10048 (N_10048,N_5354,N_6689);
or U10049 (N_10049,N_6823,N_7958);
and U10050 (N_10050,N_5274,N_6771);
nor U10051 (N_10051,N_6372,N_6592);
nand U10052 (N_10052,N_8063,N_5932);
nor U10053 (N_10053,N_9838,N_6926);
nor U10054 (N_10054,N_6369,N_5878);
xnor U10055 (N_10055,N_6818,N_7487);
and U10056 (N_10056,N_8510,N_9175);
xnor U10057 (N_10057,N_5465,N_8274);
nand U10058 (N_10058,N_5728,N_8489);
or U10059 (N_10059,N_6001,N_6457);
nor U10060 (N_10060,N_5721,N_9235);
xor U10061 (N_10061,N_8338,N_7609);
or U10062 (N_10062,N_7089,N_8532);
or U10063 (N_10063,N_7538,N_9827);
nor U10064 (N_10064,N_5398,N_5201);
nand U10065 (N_10065,N_5928,N_6599);
xor U10066 (N_10066,N_5399,N_6514);
xnor U10067 (N_10067,N_8622,N_9172);
or U10068 (N_10068,N_9918,N_5697);
and U10069 (N_10069,N_7684,N_7943);
nor U10070 (N_10070,N_9589,N_5933);
xor U10071 (N_10071,N_5596,N_6261);
and U10072 (N_10072,N_8576,N_7925);
nor U10073 (N_10073,N_5449,N_9715);
nor U10074 (N_10074,N_6556,N_9404);
nand U10075 (N_10075,N_8716,N_8924);
nor U10076 (N_10076,N_7685,N_7850);
xor U10077 (N_10077,N_5905,N_7152);
xnor U10078 (N_10078,N_5683,N_6557);
xnor U10079 (N_10079,N_7540,N_8147);
xor U10080 (N_10080,N_8269,N_9923);
nand U10081 (N_10081,N_5349,N_7178);
nand U10082 (N_10082,N_6743,N_9635);
xor U10083 (N_10083,N_8281,N_8855);
xnor U10084 (N_10084,N_9122,N_5435);
nand U10085 (N_10085,N_7432,N_8007);
or U10086 (N_10086,N_9164,N_8872);
or U10087 (N_10087,N_7401,N_6503);
nor U10088 (N_10088,N_7219,N_8131);
nor U10089 (N_10089,N_8585,N_9717);
nand U10090 (N_10090,N_7273,N_5816);
and U10091 (N_10091,N_6118,N_8414);
nor U10092 (N_10092,N_7123,N_6177);
xor U10093 (N_10093,N_6227,N_5256);
nand U10094 (N_10094,N_9869,N_5780);
and U10095 (N_10095,N_6157,N_8702);
and U10096 (N_10096,N_7183,N_7149);
or U10097 (N_10097,N_9628,N_7305);
xor U10098 (N_10098,N_9285,N_5891);
or U10099 (N_10099,N_6642,N_9182);
or U10100 (N_10100,N_9372,N_5236);
or U10101 (N_10101,N_6998,N_9791);
nor U10102 (N_10102,N_9035,N_6346);
xnor U10103 (N_10103,N_8448,N_5084);
nor U10104 (N_10104,N_5415,N_7058);
nand U10105 (N_10105,N_6751,N_7362);
xnor U10106 (N_10106,N_8179,N_8341);
nand U10107 (N_10107,N_9104,N_6479);
nand U10108 (N_10108,N_6236,N_5145);
and U10109 (N_10109,N_5047,N_7902);
or U10110 (N_10110,N_6344,N_7349);
or U10111 (N_10111,N_7783,N_9545);
xor U10112 (N_10112,N_5551,N_6467);
nand U10113 (N_10113,N_7103,N_5174);
or U10114 (N_10114,N_8444,N_7972);
and U10115 (N_10115,N_7872,N_5381);
or U10116 (N_10116,N_5811,N_8198);
and U10117 (N_10117,N_5620,N_8140);
and U10118 (N_10118,N_7016,N_7809);
xor U10119 (N_10119,N_5074,N_8429);
nor U10120 (N_10120,N_7476,N_5890);
or U10121 (N_10121,N_9700,N_5095);
nor U10122 (N_10122,N_6682,N_9755);
and U10123 (N_10123,N_5288,N_7614);
and U10124 (N_10124,N_7951,N_8579);
or U10125 (N_10125,N_8111,N_6913);
xnor U10126 (N_10126,N_6130,N_5871);
and U10127 (N_10127,N_5327,N_9524);
nor U10128 (N_10128,N_5247,N_9084);
nand U10129 (N_10129,N_7091,N_9358);
xnor U10130 (N_10130,N_6927,N_8825);
and U10131 (N_10131,N_9582,N_8482);
nor U10132 (N_10132,N_5525,N_9389);
nand U10133 (N_10133,N_6137,N_8415);
or U10134 (N_10134,N_9239,N_8788);
and U10135 (N_10135,N_6535,N_7489);
nand U10136 (N_10136,N_7915,N_8737);
xnor U10137 (N_10137,N_8762,N_8770);
and U10138 (N_10138,N_5439,N_7334);
xnor U10139 (N_10139,N_8801,N_9113);
and U10140 (N_10140,N_7288,N_9114);
nand U10141 (N_10141,N_9789,N_6154);
nand U10142 (N_10142,N_8453,N_9679);
nor U10143 (N_10143,N_9048,N_5323);
and U10144 (N_10144,N_7140,N_8763);
and U10145 (N_10145,N_5284,N_8214);
or U10146 (N_10146,N_6859,N_9117);
xor U10147 (N_10147,N_9941,N_5726);
or U10148 (N_10148,N_9989,N_7791);
xnor U10149 (N_10149,N_9740,N_5320);
xor U10150 (N_10150,N_6560,N_9417);
nor U10151 (N_10151,N_6074,N_8952);
nand U10152 (N_10152,N_7019,N_5834);
xor U10153 (N_10153,N_5817,N_7442);
nand U10154 (N_10154,N_7920,N_6269);
nand U10155 (N_10155,N_5627,N_7254);
or U10156 (N_10156,N_6002,N_5797);
and U10157 (N_10157,N_6633,N_5594);
nor U10158 (N_10158,N_7342,N_8534);
and U10159 (N_10159,N_9624,N_6934);
or U10160 (N_10160,N_9696,N_9505);
nor U10161 (N_10161,N_8750,N_9368);
or U10162 (N_10162,N_9139,N_7388);
nor U10163 (N_10163,N_5750,N_9845);
nand U10164 (N_10164,N_8597,N_9999);
xnor U10165 (N_10165,N_7161,N_6219);
xor U10166 (N_10166,N_8700,N_5286);
xnor U10167 (N_10167,N_5993,N_6401);
or U10168 (N_10168,N_7446,N_7968);
and U10169 (N_10169,N_5505,N_9096);
nand U10170 (N_10170,N_9608,N_9163);
or U10171 (N_10171,N_9920,N_9129);
nor U10172 (N_10172,N_5629,N_8629);
nor U10173 (N_10173,N_9597,N_9111);
nor U10174 (N_10174,N_6121,N_8745);
xnor U10175 (N_10175,N_6617,N_9592);
nor U10176 (N_10176,N_8790,N_5920);
and U10177 (N_10177,N_5033,N_5161);
and U10178 (N_10178,N_6309,N_6942);
xor U10179 (N_10179,N_6516,N_8166);
nand U10180 (N_10180,N_7232,N_6968);
or U10181 (N_10181,N_7500,N_7758);
xor U10182 (N_10182,N_8216,N_8255);
and U10183 (N_10183,N_5004,N_5874);
nand U10184 (N_10184,N_8436,N_6638);
or U10185 (N_10185,N_6984,N_7395);
xnor U10186 (N_10186,N_7078,N_6160);
or U10187 (N_10187,N_6523,N_5077);
or U10188 (N_10188,N_9880,N_5096);
or U10189 (N_10189,N_7536,N_6107);
xor U10190 (N_10190,N_9294,N_9398);
and U10191 (N_10191,N_8187,N_7450);
nand U10192 (N_10192,N_8324,N_6452);
nand U10193 (N_10193,N_6209,N_7096);
nor U10194 (N_10194,N_9565,N_5020);
nor U10195 (N_10195,N_8595,N_8402);
nand U10196 (N_10196,N_6899,N_5178);
nor U10197 (N_10197,N_7742,N_9409);
xnor U10198 (N_10198,N_7418,N_5378);
xnor U10199 (N_10199,N_7174,N_5831);
nand U10200 (N_10200,N_6900,N_9030);
or U10201 (N_10201,N_8256,N_5242);
nand U10202 (N_10202,N_9652,N_7693);
xnor U10203 (N_10203,N_8781,N_9718);
nor U10204 (N_10204,N_7033,N_5254);
or U10205 (N_10205,N_7979,N_6122);
nor U10206 (N_10206,N_7804,N_6675);
and U10207 (N_10207,N_7132,N_6273);
nor U10208 (N_10208,N_8713,N_8386);
nor U10209 (N_10209,N_7842,N_9851);
xor U10210 (N_10210,N_6777,N_9537);
and U10211 (N_10211,N_6448,N_9638);
or U10212 (N_10212,N_6760,N_7937);
nor U10213 (N_10213,N_8587,N_6242);
nor U10214 (N_10214,N_9522,N_6920);
or U10215 (N_10215,N_9749,N_8773);
nor U10216 (N_10216,N_6325,N_7838);
or U10217 (N_10217,N_5836,N_5187);
nor U10218 (N_10218,N_7271,N_9681);
nor U10219 (N_10219,N_5042,N_9091);
and U10220 (N_10220,N_8461,N_5692);
and U10221 (N_10221,N_6343,N_7831);
nand U10222 (N_10222,N_8698,N_6607);
and U10223 (N_10223,N_8620,N_5467);
xnor U10224 (N_10224,N_5510,N_8027);
nand U10225 (N_10225,N_8196,N_9022);
or U10226 (N_10226,N_7942,N_8372);
or U10227 (N_10227,N_5367,N_8542);
nor U10228 (N_10228,N_5607,N_5877);
nand U10229 (N_10229,N_8206,N_8837);
or U10230 (N_10230,N_8031,N_7986);
or U10231 (N_10231,N_5233,N_7667);
or U10232 (N_10232,N_5305,N_7989);
or U10233 (N_10233,N_8765,N_8623);
or U10234 (N_10234,N_8876,N_9152);
nor U10235 (N_10235,N_6761,N_6814);
or U10236 (N_10236,N_5490,N_9757);
or U10237 (N_10237,N_7572,N_6996);
and U10238 (N_10238,N_7191,N_9983);
nor U10239 (N_10239,N_7618,N_5794);
or U10240 (N_10240,N_9561,N_9702);
and U10241 (N_10241,N_7812,N_9997);
and U10242 (N_10242,N_7464,N_8057);
xnor U10243 (N_10243,N_9664,N_6707);
or U10244 (N_10244,N_7596,N_6508);
nand U10245 (N_10245,N_9461,N_5545);
nor U10246 (N_10246,N_5132,N_5902);
and U10247 (N_10247,N_7364,N_8574);
and U10248 (N_10248,N_9917,N_7526);
and U10249 (N_10249,N_5508,N_8138);
and U10250 (N_10250,N_9429,N_6288);
nand U10251 (N_10251,N_6474,N_5803);
or U10252 (N_10252,N_7524,N_7390);
or U10253 (N_10253,N_6300,N_5763);
xor U10254 (N_10254,N_7413,N_7659);
nor U10255 (N_10255,N_6446,N_7563);
or U10256 (N_10256,N_9270,N_7604);
or U10257 (N_10257,N_9839,N_7138);
xor U10258 (N_10258,N_9761,N_5036);
nand U10259 (N_10259,N_6709,N_6433);
nor U10260 (N_10260,N_5110,N_6562);
nand U10261 (N_10261,N_5542,N_8567);
or U10262 (N_10262,N_6941,N_7820);
xor U10263 (N_10263,N_7880,N_7059);
nand U10264 (N_10264,N_8478,N_8520);
xnor U10265 (N_10265,N_7289,N_5614);
nor U10266 (N_10266,N_8679,N_7185);
nand U10267 (N_10267,N_7286,N_5023);
and U10268 (N_10268,N_7293,N_6625);
xor U10269 (N_10269,N_8706,N_8973);
xor U10270 (N_10270,N_9556,N_6588);
xor U10271 (N_10271,N_8565,N_7176);
nand U10272 (N_10272,N_7180,N_6917);
or U10273 (N_10273,N_8897,N_9347);
and U10274 (N_10274,N_8182,N_7483);
or U10275 (N_10275,N_6631,N_9290);
and U10276 (N_10276,N_6870,N_6032);
or U10277 (N_10277,N_5353,N_6907);
xor U10278 (N_10278,N_8868,N_9259);
nor U10279 (N_10279,N_9547,N_6955);
xor U10280 (N_10280,N_8778,N_5571);
nor U10281 (N_10281,N_6442,N_5300);
nor U10282 (N_10282,N_9765,N_5277);
nand U10283 (N_10283,N_6059,N_6040);
or U10284 (N_10284,N_6525,N_6971);
nand U10285 (N_10285,N_6394,N_8406);
nand U10286 (N_10286,N_8445,N_7456);
and U10287 (N_10287,N_7862,N_5793);
nand U10288 (N_10288,N_5203,N_5946);
nor U10289 (N_10289,N_5584,N_8991);
nand U10290 (N_10290,N_5494,N_5104);
xor U10291 (N_10291,N_9726,N_9289);
nor U10292 (N_10292,N_7681,N_7086);
and U10293 (N_10293,N_6197,N_7368);
or U10294 (N_10294,N_5740,N_7508);
nor U10295 (N_10295,N_8601,N_8385);
nand U10296 (N_10296,N_8544,N_7075);
nor U10297 (N_10297,N_7210,N_5258);
or U10298 (N_10298,N_8840,N_8939);
xor U10299 (N_10299,N_6914,N_8374);
nand U10300 (N_10300,N_5009,N_5580);
xor U10301 (N_10301,N_7042,N_5606);
nor U10302 (N_10302,N_5833,N_9732);
and U10303 (N_10303,N_7668,N_5264);
nor U10304 (N_10304,N_9188,N_6250);
and U10305 (N_10305,N_7061,N_8383);
or U10306 (N_10306,N_6991,N_5462);
and U10307 (N_10307,N_6702,N_8285);
nand U10308 (N_10308,N_6813,N_8531);
and U10309 (N_10309,N_5079,N_6392);
nand U10310 (N_10310,N_7891,N_8686);
nor U10311 (N_10311,N_8076,N_6362);
nand U10312 (N_10312,N_9458,N_6788);
xor U10313 (N_10313,N_9144,N_8172);
nand U10314 (N_10314,N_9350,N_9621);
or U10315 (N_10315,N_5950,N_8848);
and U10316 (N_10316,N_9884,N_7122);
and U10317 (N_10317,N_6165,N_5361);
nand U10318 (N_10318,N_9173,N_9669);
nor U10319 (N_10319,N_7557,N_9243);
nor U10320 (N_10320,N_9600,N_8624);
and U10321 (N_10321,N_9455,N_8224);
nor U10322 (N_10322,N_9841,N_9663);
xnor U10323 (N_10323,N_8230,N_9946);
nand U10324 (N_10324,N_5860,N_8866);
or U10325 (N_10325,N_6710,N_6769);
or U10326 (N_10326,N_5452,N_9451);
nor U10327 (N_10327,N_6257,N_6854);
and U10328 (N_10328,N_5842,N_6935);
and U10329 (N_10329,N_6726,N_9287);
and U10330 (N_10330,N_7012,N_8008);
and U10331 (N_10331,N_8356,N_6051);
or U10332 (N_10332,N_6974,N_8263);
xnor U10333 (N_10333,N_9288,N_7298);
and U10334 (N_10334,N_9089,N_6739);
nand U10335 (N_10335,N_5645,N_7339);
xnor U10336 (N_10336,N_7265,N_6522);
and U10337 (N_10337,N_6153,N_6932);
nand U10338 (N_10338,N_6725,N_5484);
nor U10339 (N_10339,N_9305,N_8692);
or U10340 (N_10340,N_5898,N_8169);
or U10341 (N_10341,N_9636,N_7907);
nand U10342 (N_10342,N_5152,N_9058);
nand U10343 (N_10343,N_8509,N_7076);
nor U10344 (N_10344,N_6778,N_6445);
xor U10345 (N_10345,N_5705,N_8833);
or U10346 (N_10346,N_7922,N_5347);
or U10347 (N_10347,N_7374,N_7018);
or U10348 (N_10348,N_7744,N_6294);
nor U10349 (N_10349,N_9646,N_7953);
or U10350 (N_10350,N_5723,N_7532);
or U10351 (N_10351,N_6663,N_6683);
or U10352 (N_10352,N_7869,N_8552);
xnor U10353 (N_10353,N_9128,N_8742);
or U10354 (N_10354,N_5759,N_8287);
and U10355 (N_10355,N_5273,N_8307);
and U10356 (N_10356,N_9734,N_6119);
nand U10357 (N_10357,N_7249,N_9009);
nand U10358 (N_10358,N_6524,N_5285);
and U10359 (N_10359,N_6179,N_6238);
or U10360 (N_10360,N_6217,N_6779);
or U10361 (N_10361,N_9703,N_6380);
xor U10362 (N_10362,N_8295,N_8993);
or U10363 (N_10363,N_7348,N_6794);
nor U10364 (N_10364,N_9780,N_6058);
xor U10365 (N_10365,N_6052,N_6285);
xnor U10366 (N_10366,N_6124,N_9807);
xor U10367 (N_10367,N_9436,N_9119);
or U10368 (N_10368,N_7810,N_6469);
or U10369 (N_10369,N_9192,N_8102);
or U10370 (N_10370,N_5919,N_5301);
and U10371 (N_10371,N_8245,N_8756);
nor U10372 (N_10372,N_9252,N_9612);
xnor U10373 (N_10373,N_9410,N_5578);
nor U10374 (N_10374,N_6612,N_6155);
xor U10375 (N_10375,N_9064,N_6246);
nor U10376 (N_10376,N_5954,N_5234);
or U10377 (N_10377,N_8375,N_8896);
or U10378 (N_10378,N_8598,N_8013);
nor U10379 (N_10379,N_7044,N_7438);
or U10380 (N_10380,N_5395,N_8504);
and U10381 (N_10381,N_7694,N_8923);
nor U10382 (N_10382,N_9639,N_6020);
and U10383 (N_10383,N_7468,N_7246);
and U10384 (N_10384,N_8612,N_8451);
nand U10385 (N_10385,N_9370,N_6026);
nand U10386 (N_10386,N_7155,N_9102);
and U10387 (N_10387,N_8194,N_8809);
and U10388 (N_10388,N_9959,N_6376);
xor U10389 (N_10389,N_7427,N_9557);
nand U10390 (N_10390,N_6200,N_5798);
nand U10391 (N_10391,N_6151,N_5191);
and U10392 (N_10392,N_8288,N_6969);
nand U10393 (N_10393,N_6549,N_7741);
and U10394 (N_10394,N_9306,N_7952);
nand U10395 (N_10395,N_9897,N_5088);
or U10396 (N_10396,N_7743,N_7491);
xor U10397 (N_10397,N_8603,N_6742);
or U10398 (N_10398,N_6125,N_5795);
nor U10399 (N_10399,N_7244,N_8911);
and U10400 (N_10400,N_7097,N_5529);
and U10401 (N_10401,N_9196,N_5263);
or U10402 (N_10402,N_5107,N_9668);
nor U10403 (N_10403,N_5425,N_7890);
nor U10404 (N_10404,N_9683,N_6251);
or U10405 (N_10405,N_7679,N_7597);
and U10406 (N_10406,N_9453,N_5155);
xnor U10407 (N_10407,N_6199,N_8367);
nand U10408 (N_10408,N_5764,N_8468);
nand U10409 (N_10409,N_5619,N_9883);
nor U10410 (N_10410,N_7875,N_9691);
nand U10411 (N_10411,N_8380,N_7518);
or U10412 (N_10412,N_6308,N_5847);
and U10413 (N_10413,N_6053,N_7696);
nor U10414 (N_10414,N_8831,N_9319);
and U10415 (N_10415,N_8953,N_5369);
and U10416 (N_10416,N_8523,N_5472);
xor U10417 (N_10417,N_9836,N_5884);
and U10418 (N_10418,N_9631,N_9189);
xnor U10419 (N_10419,N_9846,N_9707);
nor U10420 (N_10420,N_7522,N_8673);
or U10421 (N_10421,N_5496,N_6229);
and U10422 (N_10422,N_9245,N_7347);
or U10423 (N_10423,N_8658,N_5731);
and U10424 (N_10424,N_7656,N_5761);
xor U10425 (N_10425,N_9230,N_8180);
or U10426 (N_10426,N_5734,N_5024);
or U10427 (N_10427,N_6443,N_6212);
nor U10428 (N_10428,N_5965,N_8339);
nand U10429 (N_10429,N_6608,N_9242);
nand U10430 (N_10430,N_9955,N_7165);
nor U10431 (N_10431,N_7380,N_6962);
nor U10432 (N_10432,N_8961,N_9088);
or U10433 (N_10433,N_5060,N_8120);
nor U10434 (N_10434,N_7213,N_7372);
xnor U10435 (N_10435,N_9938,N_6911);
or U10436 (N_10436,N_9994,N_5968);
or U10437 (N_10437,N_5593,N_9303);
xor U10438 (N_10438,N_8486,N_5502);
xor U10439 (N_10439,N_9892,N_8471);
nor U10440 (N_10440,N_9336,N_9298);
xor U10441 (N_10441,N_9864,N_8930);
and U10442 (N_10442,N_6353,N_7315);
and U10443 (N_10443,N_9540,N_9081);
xnor U10444 (N_10444,N_9337,N_6845);
xnor U10445 (N_10445,N_9282,N_8695);
nand U10446 (N_10446,N_5120,N_7803);
nor U10447 (N_10447,N_8087,N_9507);
xor U10448 (N_10448,N_5570,N_8362);
xor U10449 (N_10449,N_5405,N_5861);
and U10450 (N_10450,N_7221,N_8846);
nand U10451 (N_10451,N_6732,N_6100);
or U10452 (N_10452,N_7546,N_8197);
nand U10453 (N_10453,N_7017,N_8656);
or U10454 (N_10454,N_6168,N_5086);
nor U10455 (N_10455,N_7556,N_7959);
and U10456 (N_10456,N_5586,N_5599);
nor U10457 (N_10457,N_9183,N_6025);
or U10458 (N_10458,N_6510,N_9485);
nor U10459 (N_10459,N_9891,N_5711);
nand U10460 (N_10460,N_8633,N_8919);
nor U10461 (N_10461,N_5377,N_7026);
and U10462 (N_10462,N_5411,N_8559);
and U10463 (N_10463,N_6647,N_9871);
nand U10464 (N_10464,N_6450,N_9903);
or U10465 (N_10465,N_8439,N_9302);
xnor U10466 (N_10466,N_5640,N_6885);
nor U10467 (N_10467,N_6918,N_5862);
or U10468 (N_10468,N_5111,N_5999);
nor U10469 (N_10469,N_7345,N_7674);
xor U10470 (N_10470,N_5699,N_8358);
and U10471 (N_10471,N_6488,N_5719);
and U10472 (N_10472,N_6489,N_5625);
nor U10473 (N_10473,N_5013,N_5059);
nor U10474 (N_10474,N_5207,N_5141);
nor U10475 (N_10475,N_6018,N_9415);
and U10476 (N_10476,N_6678,N_5035);
nor U10477 (N_10477,N_6708,N_9850);
xnor U10478 (N_10478,N_8830,N_7663);
or U10479 (N_10479,N_5000,N_8980);
nor U10480 (N_10480,N_7829,N_5848);
xnor U10481 (N_10481,N_6048,N_7921);
and U10482 (N_10482,N_9324,N_9616);
xor U10483 (N_10483,N_7874,N_6005);
or U10484 (N_10484,N_5148,N_9974);
nor U10485 (N_10485,N_9200,N_6143);
nor U10486 (N_10486,N_5295,N_5183);
or U10487 (N_10487,N_8240,N_9414);
nand U10488 (N_10488,N_7023,N_8655);
xnor U10489 (N_10489,N_5666,N_8975);
or U10490 (N_10490,N_7126,N_9169);
and U10491 (N_10491,N_8515,N_6776);
xor U10492 (N_10492,N_9979,N_8677);
and U10493 (N_10493,N_6712,N_6298);
nor U10494 (N_10494,N_9885,N_9161);
or U10495 (N_10495,N_6277,N_5012);
xor U10496 (N_10496,N_9790,N_7041);
or U10497 (N_10497,N_9286,N_8122);
nand U10498 (N_10498,N_5324,N_9135);
or U10499 (N_10499,N_9047,N_5595);
or U10500 (N_10500,N_5559,N_8412);
nor U10501 (N_10501,N_5403,N_5591);
or U10502 (N_10502,N_5958,N_7690);
or U10503 (N_10503,N_8755,N_7085);
and U10504 (N_10504,N_6014,N_6483);
and U10505 (N_10505,N_6495,N_8313);
nand U10506 (N_10506,N_8420,N_6613);
xnor U10507 (N_10507,N_8646,N_5030);
nor U10508 (N_10508,N_6736,N_9021);
nand U10509 (N_10509,N_5298,N_7750);
or U10510 (N_10510,N_5015,N_5010);
xor U10511 (N_10511,N_5802,N_8165);
and U10512 (N_10512,N_7194,N_6011);
nand U10513 (N_10513,N_7243,N_5669);
nor U10514 (N_10514,N_9082,N_9629);
or U10515 (N_10515,N_9462,N_7726);
xnor U10516 (N_10516,N_6582,N_7034);
or U10517 (N_10517,N_5352,N_8901);
nor U10518 (N_10518,N_5427,N_5548);
xnor U10519 (N_10519,N_7773,N_9926);
nand U10520 (N_10520,N_9400,N_8107);
nor U10521 (N_10521,N_6349,N_6939);
xnor U10522 (N_10522,N_7153,N_6314);
nand U10523 (N_10523,N_7504,N_8964);
xnor U10524 (N_10524,N_8934,N_9538);
nand U10525 (N_10525,N_7731,N_7386);
or U10526 (N_10526,N_8738,N_7987);
nor U10527 (N_10527,N_5772,N_7159);
and U10528 (N_10528,N_9000,N_5908);
xor U10529 (N_10529,N_6545,N_7899);
or U10530 (N_10530,N_6825,N_6339);
or U10531 (N_10531,N_9008,N_8446);
or U10532 (N_10532,N_5546,N_9684);
and U10533 (N_10533,N_6080,N_5479);
nor U10534 (N_10534,N_7167,N_7431);
nor U10535 (N_10535,N_6869,N_6649);
or U10536 (N_10536,N_5910,N_7736);
nand U10537 (N_10537,N_6873,N_8508);
or U10538 (N_10538,N_7599,N_7624);
or U10539 (N_10539,N_7746,N_8527);
or U10540 (N_10540,N_5445,N_9025);
nor U10541 (N_10541,N_8135,N_8889);
and U10542 (N_10542,N_6838,N_6464);
and U10543 (N_10543,N_5604,N_6359);
or U10544 (N_10544,N_6850,N_5690);
and U10545 (N_10545,N_5678,N_7939);
and U10546 (N_10546,N_8047,N_8936);
nor U10547 (N_10547,N_6952,N_5424);
or U10548 (N_10548,N_5947,N_6054);
nand U10549 (N_10549,N_5837,N_5262);
xor U10550 (N_10550,N_5539,N_5296);
nand U10551 (N_10551,N_6785,N_9413);
nand U10552 (N_10552,N_7932,N_9360);
and U10553 (N_10553,N_5839,N_5245);
or U10554 (N_10554,N_7686,N_7666);
nand U10555 (N_10555,N_7886,N_7634);
or U10556 (N_10556,N_9446,N_9226);
nand U10557 (N_10557,N_9502,N_5556);
or U10558 (N_10558,N_5210,N_8862);
nor U10559 (N_10559,N_8805,N_6305);
or U10560 (N_10560,N_7762,N_5554);
nand U10561 (N_10561,N_9486,N_9204);
nand U10562 (N_10562,N_6138,N_8546);
nand U10563 (N_10563,N_9345,N_8289);
or U10564 (N_10564,N_9518,N_5280);
nand U10565 (N_10565,N_5090,N_7037);
and U10566 (N_10566,N_8450,N_8690);
xor U10567 (N_10567,N_6248,N_6271);
nor U10568 (N_10568,N_7848,N_8296);
nor U10569 (N_10569,N_8176,N_5918);
and U10570 (N_10570,N_5497,N_7145);
and U10571 (N_10571,N_8032,N_8564);
xor U10572 (N_10572,N_8721,N_7955);
xnor U10573 (N_10573,N_8957,N_6088);
or U10574 (N_10574,N_9754,N_6186);
nand U10575 (N_10575,N_8665,N_5007);
or U10576 (N_10576,N_5949,N_6834);
or U10577 (N_10577,N_8346,N_9411);
nor U10578 (N_10578,N_5799,N_5072);
or U10579 (N_10579,N_5975,N_6644);
or U10580 (N_10580,N_5366,N_7625);
nand U10581 (N_10581,N_9216,N_7099);
nor U10582 (N_10582,N_8152,N_7574);
and U10583 (N_10583,N_7992,N_6264);
or U10584 (N_10584,N_9211,N_6010);
or U10585 (N_10585,N_8938,N_5239);
xnor U10586 (N_10586,N_6497,N_5776);
or U10587 (N_10587,N_7575,N_7358);
and U10588 (N_10588,N_8012,N_7929);
and U10589 (N_10589,N_9007,N_6097);
or U10590 (N_10590,N_9623,N_6912);
and U10591 (N_10591,N_5376,N_8315);
and U10592 (N_10592,N_7445,N_9861);
nand U10593 (N_10593,N_6843,N_9103);
or U10594 (N_10594,N_6840,N_6141);
nor U10595 (N_10595,N_5257,N_8349);
nand U10596 (N_10596,N_8611,N_5244);
nand U10597 (N_10597,N_9056,N_9002);
xor U10598 (N_10598,N_9428,N_6995);
or U10599 (N_10599,N_9107,N_8393);
xor U10600 (N_10600,N_7201,N_5184);
nor U10601 (N_10601,N_7507,N_8469);
and U10602 (N_10602,N_5456,N_8246);
xnor U10603 (N_10603,N_6440,N_8079);
or U10604 (N_10604,N_6116,N_8674);
xor U10605 (N_10605,N_6256,N_7467);
xnor U10606 (N_10606,N_8907,N_6016);
or U10607 (N_10607,N_8282,N_5078);
nand U10608 (N_10608,N_9546,N_7028);
nand U10609 (N_10609,N_8299,N_8253);
nand U10610 (N_10610,N_8184,N_5641);
nor U10611 (N_10611,N_5226,N_9153);
nand U10612 (N_10612,N_8318,N_5017);
or U10613 (N_10613,N_5282,N_9363);
xnor U10614 (N_10614,N_9803,N_9065);
nand U10615 (N_10615,N_6847,N_5784);
and U10616 (N_10616,N_8098,N_7941);
nor U10617 (N_10617,N_6473,N_6808);
and U10618 (N_10618,N_6335,N_7903);
or U10619 (N_10619,N_5680,N_8505);
or U10620 (N_10620,N_7579,N_7827);
or U10621 (N_10621,N_6022,N_6894);
nand U10622 (N_10622,N_8134,N_7158);
or U10623 (N_10623,N_9121,N_6829);
xor U10624 (N_10624,N_5977,N_8110);
nor U10625 (N_10625,N_5404,N_9397);
nand U10626 (N_10626,N_5492,N_5259);
and U10627 (N_10627,N_6980,N_6391);
xor U10628 (N_10628,N_7654,N_7230);
nand U10629 (N_10629,N_8409,N_9848);
xnor U10630 (N_10630,N_9015,N_8051);
nand U10631 (N_10631,N_7612,N_6581);
nor U10632 (N_10632,N_6132,N_7982);
or U10633 (N_10633,N_8670,N_9564);
xor U10634 (N_10634,N_7366,N_7202);
nor U10635 (N_10635,N_8659,N_8715);
and U10636 (N_10636,N_7593,N_8071);
xor U10637 (N_10637,N_7020,N_5660);
nand U10638 (N_10638,N_7577,N_7601);
xor U10639 (N_10639,N_8749,N_5906);
nor U10640 (N_10640,N_5647,N_5869);
or U10641 (N_10641,N_6775,N_7720);
nand U10642 (N_10642,N_9973,N_5097);
xnor U10643 (N_10643,N_8922,N_6532);
and U10644 (N_10644,N_7242,N_7642);
nand U10645 (N_10645,N_5450,N_6494);
nand U10646 (N_10646,N_9840,N_8215);
nor U10647 (N_10647,N_8550,N_6580);
xnor U10648 (N_10648,N_7404,N_7387);
nand U10649 (N_10649,N_5688,N_9472);
or U10650 (N_10650,N_9748,N_6035);
nand U10651 (N_10651,N_6766,N_5819);
or U10652 (N_10652,N_5864,N_9029);
xor U10653 (N_10653,N_7711,N_7990);
or U10654 (N_10654,N_7985,N_6028);
nor U10655 (N_10655,N_5573,N_7303);
xor U10656 (N_10656,N_8668,N_7776);
and U10657 (N_10657,N_8011,N_9402);
nor U10658 (N_10658,N_8604,N_9484);
or U10659 (N_10659,N_8037,N_6013);
nor U10660 (N_10660,N_8776,N_6405);
or U10661 (N_10661,N_9634,N_8097);
and U10662 (N_10662,N_6718,N_6502);
nor U10663 (N_10663,N_7040,N_7005);
or U10664 (N_10664,N_7707,N_6136);
xor U10665 (N_10665,N_7252,N_6684);
nand U10666 (N_10666,N_7274,N_6648);
nor U10667 (N_10667,N_9653,N_7704);
xor U10668 (N_10668,N_8260,N_6957);
nand U10669 (N_10669,N_5386,N_9255);
nand U10670 (N_10670,N_8927,N_8421);
xnor U10671 (N_10671,N_9207,N_5027);
nor U10672 (N_10672,N_5623,N_5249);
or U10673 (N_10673,N_8942,N_7396);
nor U10674 (N_10674,N_9626,N_9130);
or U10675 (N_10675,N_6311,N_9837);
xnor U10676 (N_10676,N_7860,N_6162);
nand U10677 (N_10677,N_7539,N_5122);
xnor U10678 (N_10678,N_9314,N_5105);
nand U10679 (N_10679,N_8474,N_8054);
and U10680 (N_10680,N_5137,N_5535);
and U10681 (N_10681,N_8937,N_9813);
xor U10682 (N_10682,N_7843,N_5485);
xnor U10683 (N_10683,N_7790,N_6071);
or U10684 (N_10684,N_7470,N_7581);
xor U10685 (N_10685,N_8119,N_9013);
and U10686 (N_10686,N_8355,N_5921);
xor U10687 (N_10687,N_7683,N_9482);
nor U10688 (N_10688,N_7615,N_7355);
and U10689 (N_10689,N_6759,N_9202);
xnor U10690 (N_10690,N_5718,N_6787);
and U10691 (N_10691,N_6890,N_5480);
nor U10692 (N_10692,N_9447,N_5384);
nand U10693 (N_10693,N_9076,N_6260);
and U10694 (N_10694,N_7801,N_6296);
or U10695 (N_10695,N_5483,N_5854);
nand U10696 (N_10696,N_8249,N_5071);
nand U10697 (N_10697,N_9023,N_8452);
nand U10698 (N_10698,N_9928,N_7537);
or U10699 (N_10699,N_6041,N_9772);
xor U10700 (N_10700,N_9968,N_8376);
xor U10701 (N_10701,N_5251,N_6297);
and U10702 (N_10702,N_7523,N_7281);
or U10703 (N_10703,N_6270,N_6994);
nor U10704 (N_10704,N_7548,N_5433);
nor U10705 (N_10705,N_8433,N_7785);
or U10706 (N_10706,N_7482,N_6636);
and U10707 (N_10707,N_7151,N_6789);
nor U10708 (N_10708,N_9050,N_8487);
and U10709 (N_10709,N_6306,N_9432);
and U10710 (N_10710,N_8490,N_9544);
or U10711 (N_10711,N_8693,N_7658);
nand U10712 (N_10712,N_5516,N_6323);
or U10713 (N_10713,N_6528,N_9644);
and U10714 (N_10714,N_5653,N_9263);
xnor U10715 (N_10715,N_6239,N_6724);
nand U10716 (N_10716,N_8728,N_5228);
nand U10717 (N_10717,N_9195,N_6017);
xor U10718 (N_10718,N_5733,N_6948);
and U10719 (N_10719,N_9878,N_7594);
nor U10720 (N_10720,N_5737,N_5552);
nand U10721 (N_10721,N_7184,N_7119);
and U10722 (N_10722,N_9682,N_8799);
xnor U10723 (N_10723,N_9017,N_5032);
or U10724 (N_10724,N_6651,N_7900);
xor U10725 (N_10725,N_5172,N_7948);
nand U10726 (N_10726,N_9630,N_6015);
xor U10727 (N_10727,N_7197,N_7923);
nor U10728 (N_10728,N_8384,N_6128);
nor U10729 (N_10729,N_5613,N_6204);
and U10730 (N_10730,N_9745,N_9554);
and U10731 (N_10731,N_9690,N_5729);
xor U10732 (N_10732,N_6744,N_7199);
nand U10733 (N_10733,N_9933,N_8366);
and U10734 (N_10734,N_8457,N_8382);
and U10735 (N_10735,N_5751,N_6983);
and U10736 (N_10736,N_8591,N_9965);
nand U10737 (N_10737,N_9947,N_6594);
xnor U10738 (N_10738,N_7963,N_9435);
and U10739 (N_10739,N_8905,N_7367);
or U10740 (N_10740,N_8347,N_7447);
nor U10741 (N_10741,N_5565,N_5707);
xnor U10742 (N_10742,N_8199,N_5590);
nand U10743 (N_10743,N_8640,N_9710);
nand U10744 (N_10744,N_9449,N_9274);
xor U10745 (N_10745,N_8687,N_5180);
and U10746 (N_10746,N_5389,N_6705);
nor U10747 (N_10747,N_5312,N_5540);
or U10748 (N_10748,N_8796,N_8139);
xor U10749 (N_10749,N_7449,N_8602);
xnor U10750 (N_10750,N_6673,N_8507);
nand U10751 (N_10751,N_6662,N_6224);
nand U10752 (N_10752,N_7462,N_8731);
or U10753 (N_10753,N_8262,N_5392);
xor U10754 (N_10754,N_5536,N_6067);
or U10755 (N_10755,N_9197,N_6091);
nand U10756 (N_10756,N_8929,N_6697);
nor U10757 (N_10757,N_7329,N_5374);
nor U10758 (N_10758,N_9063,N_6540);
xnor U10759 (N_10759,N_7938,N_9018);
xor U10760 (N_10760,N_7361,N_9503);
xor U10761 (N_10761,N_5654,N_6085);
and U10762 (N_10762,N_5935,N_6981);
nand U10763 (N_10763,N_6150,N_9687);
nor U10764 (N_10764,N_9725,N_6531);
or U10765 (N_10765,N_5791,N_5094);
xor U10766 (N_10766,N_5053,N_7236);
nor U10767 (N_10767,N_9720,N_7461);
xor U10768 (N_10768,N_9110,N_8864);
or U10769 (N_10769,N_5563,N_9786);
nand U10770 (N_10770,N_7188,N_7015);
nor U10771 (N_10771,N_7606,N_5336);
nand U10772 (N_10772,N_9719,N_9595);
or U10773 (N_10773,N_5808,N_6396);
xor U10774 (N_10774,N_8065,N_6315);
or U10775 (N_10775,N_7434,N_9043);
nor U10776 (N_10776,N_6993,N_5630);
and U10777 (N_10777,N_7547,N_8669);
nand U10778 (N_10778,N_7718,N_9948);
xor U10779 (N_10779,N_5693,N_9094);
xnor U10780 (N_10780,N_8039,N_6507);
or U10781 (N_10781,N_5123,N_8501);
or U10782 (N_10782,N_7970,N_8820);
nor U10783 (N_10783,N_6418,N_8521);
nor U10784 (N_10784,N_7944,N_6909);
and U10785 (N_10785,N_7770,N_8798);
nor U10786 (N_10786,N_9145,N_6519);
nor U10787 (N_10787,N_8663,N_8572);
xnor U10788 (N_10788,N_7148,N_6801);
xnor U10789 (N_10789,N_6206,N_8954);
nand U10790 (N_10790,N_7108,N_8073);
xnor U10791 (N_10791,N_5350,N_9187);
nor U10792 (N_10792,N_9090,N_7940);
nor U10793 (N_10793,N_7864,N_5157);
nor U10794 (N_10794,N_7004,N_7936);
and U10795 (N_10795,N_6676,N_6087);
nand U10796 (N_10796,N_8159,N_7797);
or U10797 (N_10797,N_6003,N_6797);
nand U10798 (N_10798,N_7068,N_7740);
nand U10799 (N_10799,N_7332,N_7996);
and U10800 (N_10800,N_8440,N_6431);
and U10801 (N_10801,N_9031,N_5271);
nand U10802 (N_10802,N_6133,N_9898);
and U10803 (N_10803,N_7320,N_5835);
and U10804 (N_10804,N_9457,N_7065);
or U10805 (N_10805,N_6783,N_6370);
nor U10806 (N_10806,N_5135,N_8089);
and U10807 (N_10807,N_5128,N_6809);
or U10808 (N_10808,N_6301,N_6717);
nand U10809 (N_10809,N_8697,N_8496);
or U10810 (N_10810,N_5475,N_6924);
and U10811 (N_10811,N_6897,N_7110);
or U10812 (N_10812,N_9210,N_6855);
xor U10813 (N_10813,N_6304,N_5175);
nor U10814 (N_10814,N_7235,N_6982);
nand U10815 (N_10815,N_5677,N_7870);
and U10816 (N_10816,N_7109,N_7600);
nor U10817 (N_10817,N_7267,N_6956);
and U10818 (N_10818,N_9120,N_9688);
nand U10819 (N_10819,N_5283,N_6101);
and U10820 (N_10820,N_8125,N_5984);
nand U10821 (N_10821,N_8308,N_6509);
nand U10822 (N_10822,N_6062,N_5193);
or U10823 (N_10823,N_7777,N_7407);
or U10824 (N_10824,N_9829,N_5504);
nor U10825 (N_10825,N_7412,N_7056);
xor U10826 (N_10826,N_7623,N_8155);
nand U10827 (N_10827,N_7209,N_6820);
xor U10828 (N_10828,N_9072,N_8479);
or U10829 (N_10829,N_6286,N_9466);
and U10830 (N_10830,N_7551,N_9036);
xor U10831 (N_10831,N_9937,N_5749);
or U10832 (N_10832,N_8045,N_7496);
or U10833 (N_10833,N_7403,N_7515);
nor U10834 (N_10834,N_5712,N_9873);
or U10835 (N_10835,N_9375,N_8024);
xor U10836 (N_10836,N_6973,N_9701);
nand U10837 (N_10837,N_8369,N_9643);
nor U10838 (N_10838,N_8455,N_6792);
and U10839 (N_10839,N_8739,N_7957);
xnor U10840 (N_10840,N_8405,N_5937);
nor U10841 (N_10841,N_8015,N_8792);
nor U10842 (N_10842,N_8719,N_9087);
nand U10843 (N_10843,N_6093,N_7009);
and U10844 (N_10844,N_6382,N_6867);
and U10845 (N_10845,N_9333,N_6731);
xnor U10846 (N_10846,N_8438,N_5224);
nand U10847 (N_10847,N_8223,N_7529);
xnor U10848 (N_10848,N_8492,N_7115);
nand U10849 (N_10849,N_9984,N_5676);
xnor U10850 (N_10850,N_5555,N_5752);
nand U10851 (N_10851,N_9052,N_8908);
nand U10852 (N_10852,N_7816,N_9738);
nor U10853 (N_10853,N_5855,N_8885);
nand U10854 (N_10854,N_6882,N_8599);
and U10855 (N_10855,N_5133,N_8248);
and U10856 (N_10856,N_9647,N_6501);
nand U10857 (N_10857,N_8701,N_8581);
nand U10858 (N_10858,N_9146,N_7111);
xor U10859 (N_10859,N_5829,N_6438);
nand U10860 (N_10860,N_8252,N_9659);
and U10861 (N_10861,N_8635,N_5511);
xor U10862 (N_10862,N_7278,N_6055);
or U10863 (N_10863,N_6356,N_6533);
or U10864 (N_10864,N_5393,N_6081);
or U10865 (N_10865,N_6988,N_7443);
or U10866 (N_10866,N_7584,N_8321);
or U10867 (N_10867,N_9797,N_8060);
nand U10868 (N_10868,N_5945,N_6553);
and U10869 (N_10869,N_7300,N_5370);
nand U10870 (N_10870,N_9155,N_5628);
nor U10871 (N_10871,N_5940,N_5892);
or U10872 (N_10872,N_7296,N_5631);
or U10873 (N_10873,N_9832,N_9147);
nor U10874 (N_10874,N_5473,N_9194);
or U10875 (N_10875,N_8370,N_9893);
xnor U10876 (N_10876,N_6720,N_8323);
or U10877 (N_10877,N_7530,N_8028);
nor U10878 (N_10878,N_5147,N_5482);
xnor U10879 (N_10879,N_9814,N_5745);
and U10880 (N_10880,N_9985,N_9824);
nor U10881 (N_10881,N_5442,N_5760);
and U10882 (N_10882,N_6111,N_5512);
xnor U10883 (N_10883,N_7761,N_8760);
and U10884 (N_10884,N_8959,N_6077);
or U10885 (N_10885,N_6979,N_9666);
xnor U10886 (N_10886,N_5394,N_9759);
and U10887 (N_10887,N_7077,N_6896);
or U10888 (N_10888,N_7569,N_5476);
or U10889 (N_10889,N_7154,N_9258);
xnor U10890 (N_10890,N_6886,N_8241);
nor U10891 (N_10891,N_8994,N_6902);
nand U10892 (N_10892,N_9971,N_7181);
xor U10893 (N_10893,N_6265,N_9581);
nand U10894 (N_10894,N_9374,N_5486);
nor U10895 (N_10895,N_7906,N_6021);
and U10896 (N_10896,N_6218,N_9491);
and U10897 (N_10897,N_5687,N_6272);
xor U10898 (N_10898,N_9297,N_5978);
xnor U10899 (N_10899,N_9209,N_9779);
and U10900 (N_10900,N_7578,N_7371);
xnor U10901 (N_10901,N_7534,N_8514);
xor U10902 (N_10902,N_6690,N_5509);
nor U10903 (N_10903,N_8990,N_5489);
or U10904 (N_10904,N_7605,N_6878);
or U10905 (N_10905,N_7047,N_7834);
xor U10906 (N_10906,N_7826,N_8672);
and U10907 (N_10907,N_6641,N_6806);
nor U10908 (N_10908,N_6108,N_8768);
or U10909 (N_10909,N_6620,N_5904);
or U10910 (N_10910,N_6287,N_6070);
xnor U10911 (N_10911,N_6461,N_5671);
xor U10912 (N_10912,N_9733,N_6558);
xnor U10913 (N_10913,N_9876,N_8754);
xor U10914 (N_10914,N_8725,N_5478);
xnor U10915 (N_10915,N_6278,N_7568);
nor U10916 (N_10916,N_7053,N_9465);
nand U10917 (N_10917,N_7892,N_5125);
and U10918 (N_10918,N_5431,N_9262);
and U10919 (N_10919,N_6152,N_9205);
or U10920 (N_10920,N_5261,N_5988);
and U10921 (N_10921,N_8350,N_9753);
nor U10922 (N_10922,N_6455,N_8006);
nor U10923 (N_10923,N_9359,N_5328);
or U10924 (N_10924,N_7682,N_7139);
and U10925 (N_10925,N_9562,N_7800);
and U10926 (N_10926,N_9191,N_8290);
xnor U10927 (N_10927,N_7226,N_6240);
or U10928 (N_10928,N_7478,N_8932);
nand U10929 (N_10929,N_9388,N_8649);
nor U10930 (N_10930,N_7964,N_6049);
nand U10931 (N_10931,N_7114,N_6654);
nand U10932 (N_10932,N_7195,N_6938);
xor U10933 (N_10933,N_8306,N_8272);
nor U10934 (N_10934,N_6790,N_9942);
xnor U10935 (N_10935,N_8892,N_9773);
or U10936 (N_10936,N_9438,N_6653);
or U10937 (N_10937,N_7792,N_6360);
and U10938 (N_10938,N_5170,N_6203);
or U10939 (N_10939,N_8753,N_7048);
and U10940 (N_10940,N_5001,N_9042);
or U10941 (N_10941,N_9785,N_6042);
xor U10942 (N_10942,N_7335,N_7318);
and U10943 (N_10943,N_9487,N_6279);
and U10944 (N_10944,N_5742,N_7730);
or U10945 (N_10945,N_6413,N_6060);
nand U10946 (N_10946,N_7025,N_6685);
or U10947 (N_10947,N_8352,N_6804);
or U10948 (N_10948,N_8101,N_8377);
and U10949 (N_10949,N_8906,N_6453);
xor U10950 (N_10950,N_6606,N_9489);
or U10951 (N_10951,N_8251,N_8983);
nand U10952 (N_10952,N_9641,N_9558);
or U10953 (N_10953,N_5739,N_8503);
xnor U10954 (N_10954,N_5724,N_7133);
nor U10955 (N_10955,N_6749,N_8960);
and U10956 (N_10956,N_5777,N_6961);
nor U10957 (N_10957,N_6310,N_6214);
nand U10958 (N_10958,N_5139,N_9953);
or U10959 (N_10959,N_8644,N_7428);
or U10960 (N_10960,N_7472,N_6244);
nand U10961 (N_10961,N_5422,N_8064);
xnor U10962 (N_10962,N_6795,N_9776);
and U10963 (N_10963,N_7409,N_6039);
nor U10964 (N_10964,N_9272,N_7613);
nand U10965 (N_10965,N_6868,N_6303);
nor U10966 (N_10966,N_7198,N_6618);
or U10967 (N_10967,N_9116,N_5430);
nand U10968 (N_10968,N_9033,N_5887);
xnor U10969 (N_10969,N_9010,N_9593);
and U10970 (N_10970,N_6106,N_8189);
nor U10971 (N_10971,N_9815,N_9660);
xnor U10972 (N_10972,N_9875,N_7631);
nor U10973 (N_10973,N_5314,N_6569);
xnor U10974 (N_10974,N_5886,N_5447);
and U10975 (N_10975,N_8847,N_9450);
nor U10976 (N_10976,N_7737,N_5807);
nand U10977 (N_10977,N_7360,N_8210);
and U10978 (N_10978,N_8558,N_9956);
and U10979 (N_10979,N_6780,N_6406);
nand U10980 (N_10980,N_5091,N_7965);
nand U10981 (N_10981,N_8483,N_9890);
nor U10982 (N_10982,N_8454,N_5365);
and U10983 (N_10983,N_8411,N_5994);
nor U10984 (N_10984,N_8400,N_5824);
and U10985 (N_10985,N_5227,N_6812);
nand U10986 (N_10986,N_5440,N_9068);
xnor U10987 (N_10987,N_8044,N_5810);
xnor U10988 (N_10988,N_6351,N_7120);
nand U10989 (N_10989,N_7430,N_8962);
nand U10990 (N_10990,N_6094,N_7894);
xnor U10991 (N_10991,N_8839,N_5307);
or U10992 (N_10992,N_8146,N_6332);
or U10993 (N_10993,N_5943,N_9729);
or U10994 (N_10994,N_7945,N_7421);
nor U10995 (N_10995,N_7564,N_7991);
nand U10996 (N_10996,N_7405,N_9141);
nor U10997 (N_10997,N_8538,N_7806);
nand U10998 (N_10998,N_8722,N_9541);
nand U10999 (N_10999,N_7506,N_5597);
and U11000 (N_11000,N_9954,N_8589);
or U11001 (N_11001,N_9744,N_5926);
nor U11002 (N_11002,N_9340,N_8208);
xnor U11003 (N_11003,N_5025,N_7460);
nor U11004 (N_11004,N_9613,N_8005);
or U11005 (N_11005,N_7839,N_7876);
nor U11006 (N_11006,N_8232,N_8723);
xnor U11007 (N_11007,N_9332,N_5830);
or U11008 (N_11008,N_8726,N_7835);
nor U11009 (N_11009,N_8416,N_9925);
nor U11010 (N_11010,N_8475,N_5987);
and U11011 (N_11011,N_7595,N_9067);
nor U11012 (N_11012,N_5789,N_6796);
and U11013 (N_11013,N_5758,N_9418);
xnor U11014 (N_11014,N_5612,N_8516);
and U11015 (N_11015,N_9097,N_7441);
and U11016 (N_11016,N_5167,N_8522);
xor U11017 (N_11017,N_7735,N_8921);
nor U11018 (N_11018,N_8325,N_7424);
or U11019 (N_11019,N_6688,N_7960);
xor U11020 (N_11020,N_7193,N_7836);
and U11021 (N_11021,N_5562,N_6230);
and U11022 (N_11022,N_8164,N_8476);
and U11023 (N_11023,N_9412,N_5119);
nand U11024 (N_11024,N_9499,N_6949);
and U11025 (N_11025,N_8020,N_5454);
or U11026 (N_11026,N_5530,N_7164);
and U11027 (N_11027,N_9253,N_8019);
xnor U11028 (N_11028,N_6877,N_8244);
and U11029 (N_11029,N_7819,N_6220);
or U11030 (N_11030,N_9809,N_5549);
xor U11031 (N_11031,N_6754,N_7846);
nor U11032 (N_11032,N_9821,N_8949);
nand U11033 (N_11033,N_6004,N_9328);
and U11034 (N_11034,N_7100,N_7050);
nand U11035 (N_11035,N_7039,N_5576);
and U11036 (N_11036,N_5773,N_8958);
nor U11037 (N_11037,N_8336,N_5406);
xnor U11038 (N_11038,N_9810,N_7106);
xor U11039 (N_11039,N_6416,N_5235);
nand U11040 (N_11040,N_7381,N_8082);
or U11041 (N_11041,N_8364,N_5106);
and U11042 (N_11042,N_7967,N_9721);
and U11043 (N_11043,N_6928,N_7531);
nor U11044 (N_11044,N_8481,N_6851);
and U11045 (N_11045,N_8972,N_6079);
or U11046 (N_11046,N_7553,N_9513);
and U11047 (N_11047,N_7351,N_7622);
or U11048 (N_11048,N_5991,N_9727);
xnor U11049 (N_11049,N_8563,N_8292);
or U11050 (N_11050,N_7160,N_9180);
and U11051 (N_11051,N_9442,N_7171);
nand U11052 (N_11052,N_6762,N_9069);
nor U11053 (N_11053,N_8417,N_7261);
nor U11054 (N_11054,N_9697,N_9452);
or U11055 (N_11055,N_7203,N_9575);
or U11056 (N_11056,N_8775,N_8360);
and U11057 (N_11057,N_8555,N_6889);
or U11058 (N_11058,N_7343,N_5464);
nor U11059 (N_11059,N_9213,N_6842);
nor U11060 (N_11060,N_9680,N_9468);
nand U11061 (N_11061,N_9625,N_6379);
nand U11062 (N_11062,N_5882,N_5308);
and U11063 (N_11063,N_9863,N_8530);
nand U11064 (N_11064,N_8995,N_7562);
xor U11065 (N_11065,N_9250,N_7081);
nand U11066 (N_11066,N_8036,N_9711);
and U11067 (N_11067,N_9238,N_7962);
xnor U11068 (N_11068,N_6630,N_8822);
nand U11069 (N_11069,N_5215,N_9805);
and U11070 (N_11070,N_9441,N_6076);
xor U11071 (N_11071,N_7314,N_7984);
or U11072 (N_11072,N_6115,N_9533);
nor U11073 (N_11073,N_7545,N_9842);
xor U11074 (N_11074,N_7752,N_6184);
or U11075 (N_11075,N_6856,N_6645);
or U11076 (N_11076,N_7766,N_6476);
and U11077 (N_11077,N_5528,N_8040);
xnor U11078 (N_11078,N_8485,N_8743);
nand U11079 (N_11079,N_8806,N_5371);
nand U11080 (N_11080,N_7112,N_8430);
nand U11081 (N_11081,N_7304,N_5355);
and U11082 (N_11082,N_8396,N_8614);
xor U11083 (N_11083,N_8460,N_9223);
xor U11084 (N_11084,N_7821,N_8043);
xor U11085 (N_11085,N_9594,N_9676);
and U11086 (N_11086,N_6824,N_7297);
xnor U11087 (N_11087,N_7143,N_5099);
nand U11088 (N_11088,N_9443,N_9967);
nor U11089 (N_11089,N_5665,N_8228);
xor U11090 (N_11090,N_6590,N_5495);
xnor U11091 (N_11091,N_9046,N_6358);
or U11092 (N_11092,N_8613,N_5250);
or U11093 (N_11093,N_6646,N_8301);
xnor U11094 (N_11094,N_5177,N_8917);
and U11095 (N_11095,N_8893,N_5583);
or U11096 (N_11096,N_9601,N_5488);
nand U11097 (N_11097,N_5900,N_7365);
nor U11098 (N_11098,N_7765,N_9804);
nor U11099 (N_11099,N_6127,N_9819);
xnor U11100 (N_11100,N_9070,N_8095);
and U11101 (N_11101,N_7976,N_5037);
and U11102 (N_11102,N_8880,N_9901);
nor U11103 (N_11103,N_6170,N_6871);
or U11104 (N_11104,N_9222,N_7913);
or U11105 (N_11105,N_7525,N_9632);
nor U11106 (N_11106,N_5989,N_7713);
and U11107 (N_11107,N_7429,N_5684);
nor U11108 (N_11108,N_7211,N_6318);
or U11109 (N_11109,N_6793,N_5253);
xor U11110 (N_11110,N_5713,N_8042);
nor U11111 (N_11111,N_9568,N_8935);
xnor U11112 (N_11112,N_6593,N_5052);
and U11113 (N_11113,N_8554,N_8128);
nor U11114 (N_11114,N_9543,N_5732);
or U11115 (N_11115,N_9523,N_9448);
nor U11116 (N_11116,N_5643,N_7795);
or U11117 (N_11117,N_9661,N_6770);
nor U11118 (N_11118,N_8643,N_7867);
nand U11119 (N_11119,N_9823,N_7284);
nor U11120 (N_11120,N_6320,N_5056);
xor U11121 (N_11121,N_8213,N_5443);
nor U11122 (N_11122,N_6512,N_5714);
xor U11123 (N_11123,N_9714,N_8132);
nand U11124 (N_11124,N_5303,N_6929);
nand U11125 (N_11125,N_6112,N_9456);
nor U11126 (N_11126,N_7519,N_5165);
and U11127 (N_11127,N_6425,N_9151);
or U11128 (N_11128,N_6337,N_9244);
nand U11129 (N_11129,N_6216,N_6639);
xor U11130 (N_11130,N_5413,N_6375);
nand U11131 (N_11131,N_6727,N_8059);
or U11132 (N_11132,N_8075,N_9309);
nor U11133 (N_11133,N_7285,N_6420);
nand U11134 (N_11134,N_8689,N_6609);
or U11135 (N_11135,N_6904,N_9427);
and U11136 (N_11136,N_7308,N_7754);
nor U11137 (N_11137,N_6281,N_7927);
or U11138 (N_11138,N_9454,N_9387);
or U11139 (N_11139,N_7510,N_5260);
and U11140 (N_11140,N_6513,N_7516);
or U11141 (N_11141,N_9611,N_8666);
nand U11142 (N_11142,N_8150,N_5474);
xnor U11143 (N_11143,N_5717,N_7125);
xor U11144 (N_11144,N_8463,N_8078);
nand U11145 (N_11145,N_8354,N_5589);
nor U11146 (N_11146,N_5063,N_6183);
nor U11147 (N_11147,N_7357,N_6799);
and U11148 (N_11148,N_8265,N_7486);
xnor U11149 (N_11149,N_6833,N_9060);
xnor U11150 (N_11150,N_5514,N_6069);
nand U11151 (N_11151,N_6564,N_7993);
nor U11152 (N_11152,N_6322,N_6181);
nand U11153 (N_11153,N_8610,N_5722);
or U11154 (N_11154,N_8540,N_7950);
nand U11155 (N_11155,N_6078,N_5767);
and U11156 (N_11156,N_9362,N_6621);
or U11157 (N_11157,N_7911,N_6499);
and U11158 (N_11158,N_6289,N_6536);
or U11159 (N_11159,N_9536,N_7337);
nor U11160 (N_11160,N_9004,N_7645);
and U11161 (N_11161,N_9527,N_5899);
nor U11162 (N_11162,N_7353,N_7789);
xor U11163 (N_11163,N_7392,N_9913);
nor U11164 (N_11164,N_6864,N_7473);
and U11165 (N_11165,N_9437,N_6044);
nor U11166 (N_11166,N_9577,N_7781);
nor U11167 (N_11167,N_8218,N_8074);
nor U11168 (N_11168,N_9945,N_8948);
and U11169 (N_11169,N_8813,N_6368);
nand U11170 (N_11170,N_9529,N_5679);
or U11171 (N_11171,N_8304,N_9578);
and U11172 (N_11172,N_9066,N_6365);
xnor U11173 (N_11173,N_6029,N_6551);
nand U11174 (N_11174,N_5054,N_5046);
and U11175 (N_11175,N_6192,N_5109);
nand U11176 (N_11176,N_7088,N_7567);
or U11177 (N_11177,N_6090,N_8066);
xnor U11178 (N_11178,N_7260,N_6422);
nand U11179 (N_11179,N_6616,N_6176);
nand U11180 (N_11180,N_8933,N_7893);
and U11181 (N_11181,N_7722,N_5985);
or U11182 (N_11182,N_6123,N_8853);
nand U11183 (N_11183,N_6207,N_8662);
or U11184 (N_11184,N_7397,N_8004);
nand U11185 (N_11185,N_8978,N_7708);
nor U11186 (N_11186,N_8708,N_6421);
nand U11187 (N_11187,N_7794,N_5031);
nand U11188 (N_11188,N_6312,N_5659);
or U11189 (N_11189,N_9605,N_7697);
xor U11190 (N_11190,N_9907,N_8227);
nand U11191 (N_11191,N_9275,N_7206);
nor U11192 (N_11192,N_8096,N_5527);
and U11193 (N_11193,N_8779,N_9859);
or U11194 (N_11194,N_6134,N_8404);
nand U11195 (N_11195,N_6426,N_8401);
nand U11196 (N_11196,N_9622,N_5064);
nand U11197 (N_11197,N_7187,N_7196);
and U11198 (N_11198,N_6247,N_7784);
or U11199 (N_11199,N_7117,N_5289);
and U11200 (N_11200,N_8963,N_6038);
or U11201 (N_11201,N_7302,N_7087);
nand U11202 (N_11202,N_8577,N_7728);
nand U11203 (N_11203,N_7833,N_7748);
and U11204 (N_11204,N_7021,N_5821);
or U11205 (N_11205,N_7830,N_7248);
nand U11206 (N_11206,N_7259,N_5962);
nor U11207 (N_11207,N_6159,N_8425);
nand U11208 (N_11208,N_9126,N_7691);
xnor U11209 (N_11209,N_5333,N_6704);
nor U11210 (N_11210,N_8209,N_9138);
xor U11211 (N_11211,N_7454,N_9857);
nor U11212 (N_11212,N_6515,N_7352);
nor U11213 (N_11213,N_8348,N_9566);
nor U11214 (N_11214,N_5151,N_8797);
xor U11215 (N_11215,N_6437,N_8219);
or U11216 (N_11216,N_6677,N_8499);
nand U11217 (N_11217,N_7330,N_8378);
nor U11218 (N_11218,N_6602,N_7636);
nor U11219 (N_11219,N_8258,N_5917);
or U11220 (N_11220,N_5407,N_7137);
xnor U11221 (N_11221,N_8090,N_5553);
xnor U11222 (N_11222,N_6319,N_8500);
xnor U11223 (N_11223,N_9166,N_5418);
xor U11224 (N_11224,N_9548,N_7895);
nor U11225 (N_11225,N_8627,N_7775);
and U11226 (N_11226,N_5138,N_6237);
nand U11227 (N_11227,N_8777,N_8965);
xnor U11228 (N_11228,N_6354,N_9930);
nand U11229 (N_11229,N_9656,N_9831);
or U11230 (N_11230,N_5743,N_5068);
and U11231 (N_11231,N_8804,N_6803);
and U11232 (N_11232,N_8309,N_9830);
xnor U11233 (N_11233,N_8870,N_7495);
and U11234 (N_11234,N_8351,N_6600);
nand U11235 (N_11235,N_9794,N_7878);
nand U11236 (N_11236,N_6940,N_6410);
nor U11237 (N_11237,N_5214,N_9234);
and U11238 (N_11238,N_9988,N_8912);
xnor U11239 (N_11239,N_7095,N_7439);
or U11240 (N_11240,N_8419,N_8470);
or U11241 (N_11241,N_5827,N_9203);
and U11242 (N_11242,N_9694,N_9256);
nor U11243 (N_11243,N_9266,N_9346);
xor U11244 (N_11244,N_9352,N_5231);
nand U11245 (N_11245,N_7256,N_6895);
xnor U11246 (N_11246,N_5976,N_7406);
and U11247 (N_11247,N_8233,N_5658);
or U11248 (N_11248,N_6862,N_7881);
nand U11249 (N_11249,N_9532,N_6975);
xor U11250 (N_11250,N_6852,N_8175);
nor U11251 (N_11251,N_7512,N_6603);
nand U11252 (N_11252,N_9406,N_8283);
nand U11253 (N_11253,N_6950,N_8524);
xor U11254 (N_11254,N_7354,N_7868);
or U11255 (N_11255,N_5934,N_8867);
xnor U11256 (N_11256,N_8632,N_8729);
nor U11257 (N_11257,N_8116,N_6188);
nor U11258 (N_11258,N_9758,N_7866);
nand U11259 (N_11259,N_6485,N_5757);
and U11260 (N_11260,N_5341,N_5544);
nor U11261 (N_11261,N_7063,N_5896);
and U11262 (N_11262,N_8795,N_9799);
xor U11263 (N_11263,N_9806,N_9106);
xnor U11264 (N_11264,N_8578,N_5736);
nand U11265 (N_11265,N_5682,N_5615);
xor U11266 (N_11266,N_9735,N_5858);
xor U11267 (N_11267,N_6559,N_5672);
or U11268 (N_11268,N_6342,N_5038);
xnor U11269 (N_11269,N_9061,N_6552);
and U11270 (N_11270,N_6215,N_5792);
xor U11271 (N_11271,N_6943,N_8426);
xor U11272 (N_11272,N_7698,N_5022);
and U11273 (N_11273,N_9044,N_7453);
xor U11274 (N_11274,N_8886,N_9444);
xor U11275 (N_11275,N_9716,N_8609);
and U11276 (N_11276,N_8875,N_8941);
xnor U11277 (N_11277,N_6632,N_8319);
and U11278 (N_11278,N_7885,N_9767);
and U11279 (N_11279,N_5219,N_5938);
or U11280 (N_11280,N_8767,N_7307);
nand U11281 (N_11281,N_6923,N_5237);
xnor U11282 (N_11282,N_8345,N_8413);
nand U11283 (N_11283,N_9344,N_6355);
xnor U11284 (N_11284,N_9852,N_8810);
and U11285 (N_11285,N_5444,N_6876);
nor U11286 (N_11286,N_8264,N_9552);
and U11287 (N_11287,N_9737,N_7550);
and U11288 (N_11288,N_6427,N_9278);
and U11289 (N_11289,N_7469,N_9198);
xor U11290 (N_11290,N_5644,N_5338);
xor U11291 (N_11291,N_8170,N_8472);
xor U11292 (N_11292,N_7287,N_5344);
and U11293 (N_11293,N_6872,N_9386);
nor U11294 (N_11294,N_6284,N_7904);
and U11295 (N_11295,N_6622,N_8141);
or U11296 (N_11296,N_6687,N_5098);
or U11297 (N_11297,N_7146,N_7756);
nand U11298 (N_11298,N_9981,N_5661);
or U11299 (N_11299,N_8242,N_8821);
xnor U11300 (N_11300,N_9751,N_6748);
nor U11301 (N_11301,N_7739,N_8910);
xnor U11302 (N_11302,N_7734,N_7426);
xor U11303 (N_11303,N_7994,N_5694);
xor U11304 (N_11304,N_7847,N_6412);
or U11305 (N_11305,N_7974,N_7660);
and U11306 (N_11306,N_9793,N_6441);
nand U11307 (N_11307,N_8204,N_6072);
and U11308 (N_11308,N_8680,N_6841);
xnor U11309 (N_11309,N_6407,N_9327);
and U11310 (N_11310,N_6672,N_6543);
or U11311 (N_11311,N_7554,N_5868);
nor U11312 (N_11312,N_5706,N_8118);
xnor U11313 (N_11313,N_5292,N_8786);
xnor U11314 (N_11314,N_7054,N_8593);
or U11315 (N_11315,N_9420,N_5893);
or U11316 (N_11316,N_9424,N_9251);
or U11317 (N_11317,N_5621,N_6554);
and U11318 (N_11318,N_9508,N_8394);
nor U11319 (N_11319,N_8616,N_6348);
nand U11320 (N_11320,N_7517,N_6147);
and U11321 (N_11321,N_8067,N_5129);
xnor U11322 (N_11322,N_5663,N_8235);
nand U11323 (N_11323,N_7166,N_6043);
nor U11324 (N_11324,N_5727,N_7481);
nand U11325 (N_11325,N_7182,N_8641);
nand U11326 (N_11326,N_5569,N_7665);
nor U11327 (N_11327,N_6596,N_7549);
and U11328 (N_11328,N_5880,N_6965);
and U11329 (N_11329,N_8432,N_8133);
and U11330 (N_11330,N_7977,N_9870);
nor U11331 (N_11331,N_9781,N_6936);
and U11332 (N_11332,N_5501,N_5853);
nor U11333 (N_11333,N_5302,N_9675);
or U11334 (N_11334,N_8676,N_9670);
nor U11335 (N_11335,N_5453,N_9579);
xnor U11336 (N_11336,N_5319,N_6848);
xor U11337 (N_11337,N_9269,N_5116);
xnor U11338 (N_11338,N_8163,N_5471);
nand U11339 (N_11339,N_5217,N_7772);
nand U11340 (N_11340,N_8970,N_6189);
and U11341 (N_11341,N_9098,N_5635);
nor U11342 (N_11342,N_8545,N_9963);
or U11343 (N_11343,N_6741,N_5587);
xor U11344 (N_11344,N_5487,N_8944);
nor U11345 (N_11345,N_5929,N_6178);
and U11346 (N_11346,N_9525,N_8812);
xnor U11347 (N_11347,N_5812,N_5967);
nand U11348 (N_11348,N_9312,N_5045);
nand U11349 (N_11349,N_9349,N_8771);
nor U11350 (N_11350,N_9321,N_8811);
xnor U11351 (N_11351,N_8447,N_8137);
nand U11352 (N_11352,N_6526,N_8829);
xnor U11353 (N_11353,N_8212,N_8539);
nand U11354 (N_11354,N_5774,N_7620);
and U11355 (N_11355,N_6729,N_5357);
nand U11356 (N_11356,N_9705,N_9987);
nand U11357 (N_11357,N_6057,N_8099);
nor U11358 (N_11358,N_5225,N_7749);
nand U11359 (N_11359,N_7755,N_6267);
nor U11360 (N_11360,N_8898,N_8575);
nand U11361 (N_11361,N_9940,N_5616);
nand U11362 (N_11362,N_8547,N_8618);
or U11363 (N_11363,N_5278,N_5849);
xnor U11364 (N_11364,N_5970,N_7592);
nor U11365 (N_11365,N_5069,N_6958);
xor U11366 (N_11366,N_7052,N_9381);
nor U11367 (N_11367,N_6668,N_8053);
xor U11368 (N_11368,N_9284,N_9228);
or U11369 (N_11369,N_7333,N_5150);
nor U11370 (N_11370,N_6031,N_7786);
and U11371 (N_11371,N_9109,N_5076);
and U11372 (N_11372,N_5335,N_8996);
xor U11373 (N_11373,N_5008,N_5915);
or U11374 (N_11374,N_5470,N_7128);
or U11375 (N_11375,N_5229,N_9348);
xor U11376 (N_11376,N_6444,N_8480);
xor U11377 (N_11377,N_7035,N_8337);
nand U11378 (N_11378,N_8190,N_7241);
nand U11379 (N_11379,N_5903,N_8205);
nor U11380 (N_11380,N_7463,N_5267);
nand U11381 (N_11381,N_8685,N_5149);
xor U11382 (N_11382,N_7703,N_5691);
xor U11383 (N_11383,N_8845,N_7168);
nand U11384 (N_11384,N_8302,N_7057);
xor U11385 (N_11385,N_5783,N_8774);
and U11386 (N_11386,N_5205,N_8682);
and U11387 (N_11387,N_5208,N_5818);
and U11388 (N_11388,N_8631,N_5681);
or U11389 (N_11389,N_8625,N_9966);
xor U11390 (N_11390,N_8863,N_8720);
xor U11391 (N_11391,N_6487,N_7007);
nor U11392 (N_11392,N_8865,N_5841);
and U11393 (N_11393,N_6520,N_5506);
xnor U11394 (N_11394,N_7062,N_5387);
and U11395 (N_11395,N_5995,N_6324);
or U11396 (N_11396,N_5972,N_6210);
and U11397 (N_11397,N_7069,N_9939);
nand U11398 (N_11398,N_6953,N_7299);
or U11399 (N_11399,N_6208,N_6492);
nand U11400 (N_11400,N_7738,N_5957);
nand U11401 (N_11401,N_6142,N_5186);
or U11402 (N_11402,N_7436,N_5315);
and U11403 (N_11403,N_8628,N_6693);
nand U11404 (N_11404,N_9627,N_5154);
nor U11405 (N_11405,N_8427,N_7079);
nand U11406 (N_11406,N_5153,N_8177);
xor U11407 (N_11407,N_9260,N_7768);
nor U11408 (N_11408,N_6541,N_7505);
or U11409 (N_11409,N_8160,N_7045);
and U11410 (N_11410,N_5513,N_6213);
or U11411 (N_11411,N_8192,N_7317);
nor U11412 (N_11412,N_9866,N_9674);
xnor U11413 (N_11413,N_8456,N_5196);
xnor U11414 (N_11414,N_7859,N_7282);
or U11415 (N_11415,N_5421,N_9467);
and U11416 (N_11416,N_9990,N_7275);
xor U11417 (N_11417,N_9555,N_8226);
xnor U11418 (N_11418,N_7212,N_7070);
xnor U11419 (N_11419,N_7619,N_8343);
and U11420 (N_11420,N_7702,N_5564);
xnor U11421 (N_11421,N_5925,N_8891);
or U11422 (N_11422,N_9176,N_9219);
nand U11423 (N_11423,N_6408,N_8086);
xor U11424 (N_11424,N_8909,N_5185);
xor U11425 (N_11425,N_5065,N_6874);
xnor U11426 (N_11426,N_9698,N_8817);
nor U11427 (N_11427,N_8498,N_6921);
or U11428 (N_11428,N_8667,N_8494);
or U11429 (N_11429,N_6737,N_9331);
or U11430 (N_11430,N_9782,N_6960);
or U11431 (N_11431,N_5372,N_8769);
xnor U11432 (N_11432,N_9247,N_9858);
nor U11433 (N_11433,N_7729,N_5507);
nand U11434 (N_11434,N_8651,N_7107);
or U11435 (N_11435,N_6140,N_7144);
and U11436 (N_11436,N_6156,N_9896);
or U11437 (N_11437,N_7150,N_7916);
nand U11438 (N_11438,N_6084,N_7032);
and U11439 (N_11439,N_9281,N_7163);
or U11440 (N_11440,N_9908,N_7672);
and U11441 (N_11441,N_8211,N_7200);
or U11442 (N_11442,N_6338,N_5041);
nor U11443 (N_11443,N_7090,N_8434);
xnor U11444 (N_11444,N_9073,N_6388);
nor U11445 (N_11445,N_6317,N_7321);
nor U11446 (N_11446,N_9777,N_5863);
or U11447 (N_11447,N_7014,N_7509);
nor U11448 (N_11448,N_6735,N_6158);
xnor U11449 (N_11449,N_6756,N_9257);
xor U11450 (N_11450,N_7074,N_5358);
and U11451 (N_11451,N_9934,N_6164);
and U11452 (N_11452,N_5121,N_9330);
xnor U11453 (N_11453,N_6881,N_5043);
nor U11454 (N_11454,N_9240,N_6666);
nor U11455 (N_11455,N_9277,N_8458);
and U11456 (N_11456,N_9924,N_5881);
xnor U11457 (N_11457,N_9071,N_5873);
xnor U11458 (N_11458,N_9563,N_6883);
xnor U11459 (N_11459,N_9335,N_5313);
nor U11460 (N_11460,N_7745,N_6986);
nand U11461 (N_11461,N_6832,N_8293);
nand U11462 (N_11462,N_8243,N_5624);
nor U11463 (N_11463,N_6879,N_8270);
or U11464 (N_11464,N_8881,N_9872);
nor U11465 (N_11465,N_5521,N_8619);
nand U11466 (N_11466,N_8121,N_9016);
and U11467 (N_11467,N_7129,N_7935);
or U11468 (N_11468,N_7399,N_7479);
nor U11469 (N_11469,N_9868,N_7323);
nor U11470 (N_11470,N_6460,N_5238);
and U11471 (N_11471,N_8989,N_6275);
nor U11472 (N_11472,N_9483,N_9648);
and U11473 (N_11473,N_6667,N_6931);
xor U11474 (N_11474,N_5294,N_8069);
or U11475 (N_11475,N_5828,N_7747);
or U11476 (N_11476,N_9123,N_8488);
nand U11477 (N_11477,N_7131,N_8314);
nor U11478 (N_11478,N_8733,N_8879);
and U11479 (N_11479,N_8010,N_7043);
xnor U11480 (N_11480,N_9567,N_9783);
xor U11481 (N_11481,N_7452,N_9339);
nor U11482 (N_11482,N_5455,N_8752);
or U11483 (N_11483,N_7073,N_9342);
or U11484 (N_11484,N_8757,N_6892);
xnor U11485 (N_11485,N_7369,N_8114);
and U11486 (N_11486,N_6000,N_8816);
nand U11487 (N_11487,N_7101,N_5786);
or U11488 (N_11488,N_5246,N_8462);
or U11489 (N_11489,N_5911,N_9633);
or U11490 (N_11490,N_9134,N_7071);
nor U11491 (N_11491,N_6572,N_7344);
nor U11492 (N_11492,N_6805,N_5850);
nor U11493 (N_11493,N_6774,N_8273);
and U11494 (N_11494,N_9618,N_8149);
xnor U11495 (N_11495,N_7813,N_7648);
or U11496 (N_11496,N_8638,N_7147);
xnor U11497 (N_11497,N_8398,N_6714);
or U11498 (N_11498,N_9818,N_6398);
and U11499 (N_11499,N_9542,N_9530);
nand U11500 (N_11500,N_8049,N_7223);
xor U11501 (N_11501,N_9834,N_6821);
nor U11502 (N_11502,N_8136,N_9642);
xor U11503 (N_11503,N_8654,N_9756);
nand U11504 (N_11504,N_5463,N_8088);
xor U11505 (N_11505,N_8181,N_7229);
or U11506 (N_11506,N_5575,N_7566);
nand U11507 (N_11507,N_5034,N_7102);
nor U11508 (N_11508,N_8854,N_9986);
and U11509 (N_11509,N_8171,N_8320);
nor U11510 (N_11510,N_8955,N_7845);
xnor U11511 (N_11511,N_9936,N_5039);
and U11512 (N_11512,N_5859,N_7882);
nor U11513 (N_11513,N_6836,N_5322);
nand U11514 (N_11514,N_7723,N_7917);
xnor U11515 (N_11515,N_9080,N_8647);
nand U11516 (N_11516,N_7558,N_7552);
or U11517 (N_11517,N_5708,N_5885);
nand U11518 (N_11518,N_9728,N_5840);
nor U11519 (N_11519,N_8977,N_9706);
nor U11520 (N_11520,N_5345,N_7383);
nor U11521 (N_11521,N_5689,N_5160);
and U11522 (N_11522,N_6045,N_8590);
and U11523 (N_11523,N_8951,N_8869);
nor U11524 (N_11524,N_7721,N_6393);
xnor U11525 (N_11525,N_6066,N_9519);
or U11526 (N_11526,N_9867,N_5762);
nor U11527 (N_11527,N_9405,N_9931);
nand U11528 (N_11528,N_8025,N_9142);
and U11529 (N_11529,N_9391,N_6734);
nand U11530 (N_11530,N_5537,N_5969);
or U11531 (N_11531,N_6905,N_8842);
nor U11532 (N_11532,N_6249,N_9617);
nand U11533 (N_11533,N_5916,N_9909);
xor U11534 (N_11534,N_8185,N_6703);
xnor U11535 (N_11535,N_6990,N_7488);
xor U11536 (N_11536,N_9534,N_8278);
or U11537 (N_11537,N_9672,N_7695);
nor U11538 (N_11538,N_6363,N_7310);
or U11539 (N_11539,N_9361,N_7798);
nor U11540 (N_11540,N_6490,N_5176);
nand U11541 (N_11541,N_9604,N_7774);
nand U11542 (N_11542,N_6366,N_8694);
nand U11543 (N_11543,N_6135,N_7640);
and U11544 (N_11544,N_9214,N_6915);
or U11545 (N_11545,N_9199,N_9667);
xor U11546 (N_11546,N_9905,N_9232);
nor U11547 (N_11547,N_9475,N_7008);
and U11548 (N_11548,N_5522,N_8596);
and U11549 (N_11549,N_5941,N_6331);
and U11550 (N_11550,N_8982,N_5162);
and U11551 (N_11551,N_5702,N_9075);
xnor U11552 (N_11552,N_6901,N_7912);
nor U11553 (N_11553,N_8130,N_9229);
nand U11554 (N_11554,N_8191,N_9958);
nand U11555 (N_11555,N_9811,N_6430);
nor U11556 (N_11556,N_8580,N_5199);
or U11557 (N_11557,N_8645,N_8195);
or U11558 (N_11558,N_5966,N_8250);
xnor U11559 (N_11559,N_5202,N_5140);
xor U11560 (N_11560,N_9526,N_9730);
nand U11561 (N_11561,N_7013,N_8918);
nand U11562 (N_11562,N_8634,N_7218);
nor U11563 (N_11563,N_8158,N_5223);
nand U11564 (N_11564,N_9723,N_5080);
or U11565 (N_11565,N_8736,N_7716);
xnor U11566 (N_11566,N_9383,N_8688);
or U11567 (N_11567,N_5951,N_8142);
nor U11568 (N_11568,N_9171,N_6185);
nand U11569 (N_11569,N_9559,N_5730);
nor U11570 (N_11570,N_9576,N_9610);
and U11571 (N_11571,N_7788,N_7855);
xnor U11572 (N_11572,N_5936,N_8284);
or U11573 (N_11573,N_9311,N_5062);
or U11574 (N_11574,N_9488,N_6634);
nand U11575 (N_11575,N_8327,N_7759);
nand U11576 (N_11576,N_9101,N_8569);
nor U11577 (N_11577,N_9040,N_6568);
or U11578 (N_11578,N_5255,N_5321);
nor U11579 (N_11579,N_5875,N_6586);
and U11580 (N_11580,N_7863,N_7706);
nand U11581 (N_11581,N_8229,N_7565);
or U11582 (N_11582,N_9307,N_9860);
xor U11583 (N_11583,N_7127,N_6180);
or U11584 (N_11584,N_6574,N_6030);
xnor U11585 (N_11585,N_5997,N_9874);
nand U11586 (N_11586,N_8407,N_5342);
xor U11587 (N_11587,N_9572,N_8268);
nand U11588 (N_11588,N_6006,N_9645);
nor U11589 (N_11589,N_9996,N_5953);
and U11590 (N_11590,N_6415,N_7066);
nand U11591 (N_11591,N_5368,N_9108);
and U11592 (N_11592,N_8115,N_7162);
or U11593 (N_11593,N_7105,N_8874);
nor U11594 (N_11594,N_6061,N_5092);
and U11595 (N_11595,N_5340,N_5272);
xor U11596 (N_11596,N_5585,N_5204);
and U11597 (N_11597,N_7817,N_7956);
xor U11598 (N_11598,N_8424,N_6295);
nand U11599 (N_11599,N_6089,N_7328);
nand U11600 (N_11600,N_8586,N_9012);
nand U11601 (N_11601,N_5716,N_8373);
nand U11602 (N_11602,N_7910,N_5144);
nor U11603 (N_11603,N_8684,N_8732);
xor U11604 (N_11604,N_9384,N_9609);
nand U11605 (N_11605,N_6007,N_5856);
nand U11606 (N_11606,N_8104,N_8387);
xor U11607 (N_11607,N_5426,N_9798);
xor U11608 (N_11608,N_5768,N_9902);
nor U11609 (N_11609,N_7466,N_7179);
nand U11610 (N_11610,N_9371,N_6068);
and U11611 (N_11611,N_8562,N_7586);
and U11612 (N_11612,N_5343,N_6472);
and U11613 (N_11613,N_5588,N_9739);
xnor U11614 (N_11614,N_7603,N_9517);
and U11615 (N_11615,N_7217,N_7629);
nor U11616 (N_11616,N_8890,N_8671);
xor U11617 (N_11617,N_5163,N_9396);
xnor U11618 (N_11618,N_6865,N_9174);
or U11619 (N_11619,N_9619,N_7896);
or U11620 (N_11620,N_9591,N_6193);
xnor U11621 (N_11621,N_9212,N_8844);
nand U11622 (N_11622,N_6449,N_8259);
or U11623 (N_11623,N_5673,N_8145);
xor U11624 (N_11624,N_9157,N_5220);
or U11625 (N_11625,N_7520,N_9919);
nor U11626 (N_11626,N_8513,N_8092);
xnor U11627 (N_11627,N_6811,N_6925);
nand U11628 (N_11628,N_6837,N_7402);
nor U11629 (N_11629,N_7560,N_5166);
and U11630 (N_11630,N_7262,N_6432);
nor U11631 (N_11631,N_5493,N_6280);
or U11632 (N_11632,N_7664,N_7555);
nor U11633 (N_11633,N_8916,N_5814);
nor U11634 (N_11634,N_6987,N_5330);
xnor U11635 (N_11635,N_6105,N_8261);
nor U11636 (N_11636,N_9390,N_9888);
or U11637 (N_11637,N_5686,N_9178);
nand U11638 (N_11638,N_6849,N_5083);
xnor U11639 (N_11639,N_9304,N_9960);
nor U11640 (N_11640,N_7340,N_6664);
or U11641 (N_11641,N_7474,N_9479);
nor U11642 (N_11642,N_6933,N_6888);
or U11643 (N_11643,N_5913,N_9382);
nor U11644 (N_11644,N_8592,N_8123);
nor U11645 (N_11645,N_6629,N_6439);
nand U11646 (N_11646,N_9301,N_6334);
xor U11647 (N_11647,N_5964,N_6951);
and U11648 (N_11648,N_6175,N_5058);
nor U11649 (N_11649,N_5113,N_9426);
xnor U11650 (N_11650,N_9784,N_8712);
or U11651 (N_11651,N_6414,N_8675);
or U11652 (N_11652,N_8946,N_7998);
nor U11653 (N_11653,N_9894,N_8529);
nor U11654 (N_11654,N_9816,N_7029);
nand U11655 (N_11655,N_9170,N_5209);
nand U11656 (N_11656,N_6255,N_6475);
xor U11657 (N_11657,N_9434,N_8557);
or U11658 (N_11658,N_9393,N_8832);
nand U11659 (N_11659,N_5026,N_8217);
and U11660 (N_11660,N_9296,N_8056);
nand U11661 (N_11661,N_9431,N_6828);
and U11662 (N_11662,N_6802,N_9341);
or U11663 (N_11663,N_9149,N_5266);
xnor U11664 (N_11664,N_6012,N_8017);
and U11665 (N_11665,N_6386,N_6922);
or U11666 (N_11666,N_7583,N_6571);
or U11667 (N_11667,N_6578,N_6765);
nor U11668 (N_11668,N_5766,N_6104);
nand U11669 (N_11669,N_7093,N_7591);
nor U11670 (N_11670,N_8976,N_9158);
and U11671 (N_11671,N_6716,N_5412);
nand U11672 (N_11672,N_9788,N_6374);
or U11673 (N_11673,N_5481,N_7391);
or U11674 (N_11674,N_6493,N_6462);
and U11675 (N_11675,N_5741,N_8707);
xnor U11676 (N_11676,N_5603,N_9167);
or U11677 (N_11677,N_6345,N_7425);
nand U11678 (N_11678,N_6544,N_6486);
or U11679 (N_11679,N_9334,N_9159);
and U11680 (N_11680,N_8615,N_9855);
xor U11681 (N_11681,N_9746,N_8956);
and U11682 (N_11682,N_5390,N_7644);
xnor U11683 (N_11683,N_8704,N_9227);
xnor U11684 (N_11684,N_8334,N_7767);
and U11685 (N_11685,N_6985,N_6604);
and U11686 (N_11686,N_8477,N_9133);
or U11687 (N_11687,N_6767,N_9132);
xor U11688 (N_11688,N_7671,N_8127);
nand U11689 (N_11689,N_8860,N_6095);
nand U11690 (N_11690,N_9620,N_7975);
nor U11691 (N_11691,N_8974,N_9150);
and U11692 (N_11692,N_9055,N_8442);
nand U11693 (N_11693,N_5602,N_7067);
and U11694 (N_11694,N_9731,N_9962);
and U11695 (N_11695,N_7590,N_6728);
nor U11696 (N_11696,N_5198,N_8168);
nor U11697 (N_11697,N_9224,N_8789);
and U11698 (N_11698,N_9689,N_6173);
nor U11699 (N_11699,N_6340,N_8877);
and U11700 (N_11700,N_7245,N_8431);
nor U11701 (N_11701,N_9474,N_5801);
nand U11702 (N_11702,N_7104,N_8784);
nor U11703 (N_11703,N_6643,N_8998);
and U11704 (N_11704,N_7588,N_6330);
nor U11705 (N_11705,N_6605,N_5216);
and U11706 (N_11706,N_6436,N_5960);
xor U11707 (N_11707,N_5872,N_8077);
nor U11708 (N_11708,N_9498,N_6946);
nor U11709 (N_11709,N_6350,N_7688);
nor U11710 (N_11710,N_7475,N_8718);
or U11711 (N_11711,N_6816,N_7919);
xor U11712 (N_11712,N_8021,N_9131);
and U11713 (N_11713,N_5700,N_8225);
xnor U11714 (N_11714,N_6466,N_7822);
and U11715 (N_11715,N_7389,N_8815);
and U11716 (N_11716,N_9654,N_8984);
or U11717 (N_11717,N_6656,N_5115);
nand U11718 (N_11718,N_7423,N_6471);
xor U11719 (N_11719,N_7394,N_8661);
nand U11720 (N_11720,N_6329,N_8543);
or U11721 (N_11721,N_9512,N_9750);
xnor U11722 (N_11722,N_8371,N_9520);
or U11723 (N_11723,N_9215,N_5383);
or U11724 (N_11724,N_5538,N_6970);
or U11725 (N_11725,N_7156,N_5401);
xnor U11726 (N_11726,N_5417,N_6614);
nand U11727 (N_11727,N_7459,N_7961);
xor U11728 (N_11728,N_5279,N_8340);
nand U11729 (N_11729,N_9316,N_9879);
xnor U11730 (N_11730,N_5388,N_8286);
xor U11731 (N_11731,N_5169,N_7170);
or U11732 (N_11732,N_8124,N_8518);
or U11733 (N_11733,N_6686,N_6129);
and U11734 (N_11734,N_6561,N_5543);
or U11735 (N_11735,N_6034,N_9317);
xnor U11736 (N_11736,N_8294,N_6505);
nand U11737 (N_11737,N_6290,N_9125);
or U11738 (N_11738,N_7573,N_5181);
and U11739 (N_11739,N_8202,N_7780);
nand U11740 (N_11740,N_5574,N_7437);
nand U11741 (N_11741,N_9775,N_8913);
and U11742 (N_11742,N_9254,N_8247);
nand U11743 (N_11743,N_5318,N_5804);
and U11744 (N_11744,N_9325,N_7677);
nor U11745 (N_11745,N_9970,N_8584);
xor U11746 (N_11746,N_9650,N_5622);
nor U11747 (N_11747,N_6171,N_8103);
xor U11748 (N_11748,N_7239,N_8266);
nand U11749 (N_11749,N_6341,N_8714);
and U11750 (N_11750,N_8231,N_6292);
nand U11751 (N_11751,N_5754,N_8144);
xor U11752 (N_11752,N_5845,N_7322);
or U11753 (N_11753,N_9607,N_9045);
nand U11754 (N_11754,N_9403,N_5211);
xor U11755 (N_11755,N_8836,N_9394);
and U11756 (N_11756,N_5028,N_7083);
xor U11757 (N_11757,N_8117,N_7382);
and U11758 (N_11758,N_8342,N_8594);
xor U11759 (N_11759,N_7898,N_7610);
xnor U11760 (N_11760,N_7901,N_7851);
nand U11761 (N_11761,N_5136,N_6972);
nand U11762 (N_11762,N_8084,N_9220);
nand U11763 (N_11763,N_7924,N_6746);
or U11764 (N_11764,N_9769,N_9796);
nand U11765 (N_11765,N_6245,N_7724);
nor U11766 (N_11766,N_9514,N_5143);
xnor U11767 (N_11767,N_5402,N_5605);
nand U11768 (N_11768,N_6491,N_5782);
xnor U11769 (N_11769,N_6903,N_8818);
xor U11770 (N_11770,N_6268,N_9573);
and U11771 (N_11771,N_7585,N_5971);
xor U11772 (N_11772,N_8410,N_9471);
nor U11773 (N_11773,N_7484,N_5499);
or U11774 (N_11774,N_6149,N_7225);
xor U11775 (N_11775,N_8642,N_7969);
nand U11776 (N_11776,N_7840,N_8234);
or U11777 (N_11777,N_8988,N_8239);
xnor U11778 (N_11778,N_7673,N_7811);
xnor U11779 (N_11779,N_5195,N_8617);
nor U11780 (N_11780,N_5769,N_6758);
or U11781 (N_11781,N_8335,N_6109);
nor U11782 (N_11782,N_5287,N_7175);
nand U11783 (N_11783,N_5182,N_5823);
and U11784 (N_11784,N_9640,N_9006);
and U11785 (N_11785,N_7884,N_6764);
nor U11786 (N_11786,N_5332,N_5638);
xor U11787 (N_11787,N_8841,N_5838);
xor U11788 (N_11788,N_8657,N_6992);
nor U11789 (N_11789,N_7779,N_8236);
or U11790 (N_11790,N_6096,N_6719);
and U11791 (N_11791,N_5963,N_8807);
xnor U11792 (N_11792,N_9477,N_9580);
xnor U11793 (N_11793,N_7871,N_7999);
xor U11794 (N_11794,N_6463,N_6964);
xnor U11795 (N_11795,N_7224,N_9980);
nand U11796 (N_11796,N_5770,N_6397);
xnor U11797 (N_11797,N_7377,N_5579);
or U11798 (N_11798,N_6730,N_5363);
xor U11799 (N_11799,N_9473,N_6826);
or U11800 (N_11800,N_6782,N_5409);
or U11801 (N_11801,N_8764,N_5103);
nor U11802 (N_11802,N_9032,N_7832);
or U11803 (N_11803,N_7971,N_7818);
nor U11804 (N_11804,N_5029,N_5297);
or U11805 (N_11805,N_8740,N_6619);
nor U11806 (N_11806,N_5351,N_9820);
nor U11807 (N_11807,N_6945,N_9143);
and U11808 (N_11808,N_6110,N_9982);
xnor U11809 (N_11809,N_6102,N_5005);
xor U11810 (N_11810,N_5639,N_8003);
or U11811 (N_11811,N_8437,N_7676);
nor U11812 (N_11812,N_9763,N_5391);
xnor U11813 (N_11813,N_9049,N_9124);
xnor U11814 (N_11814,N_9378,N_5061);
xnor U11815 (N_11815,N_5558,N_7204);
nand U11816 (N_11816,N_9478,N_6875);
or U11817 (N_11817,N_6635,N_5825);
or U11818 (N_11818,N_6232,N_7006);
nand U11819 (N_11819,N_5520,N_5146);
nand U11820 (N_11820,N_6591,N_8423);
xor U11821 (N_11821,N_9118,N_5364);
or U11822 (N_11822,N_7309,N_9078);
and U11823 (N_11823,N_8947,N_6745);
nor U11824 (N_11824,N_7502,N_8193);
nand U11825 (N_11825,N_7632,N_9590);
nand U11826 (N_11826,N_6773,N_5755);
xnor U11827 (N_11827,N_8683,N_6768);
or U11828 (N_11828,N_6146,N_9074);
nor U11829 (N_11829,N_8093,N_5093);
nand U11830 (N_11830,N_8300,N_6555);
nor U11831 (N_11831,N_9569,N_8605);
nand U11832 (N_11832,N_9459,N_5897);
nand U11833 (N_11833,N_9062,N_7400);
and U11834 (N_11834,N_7134,N_5458);
nand U11835 (N_11835,N_8316,N_9165);
xor U11836 (N_11836,N_7393,N_7621);
nand U11837 (N_11837,N_9395,N_6399);
or U11838 (N_11838,N_6019,N_9795);
or U11839 (N_11839,N_7220,N_8154);
nand U11840 (N_11840,N_6145,N_8203);
or U11841 (N_11841,N_5410,N_7778);
nor U11842 (N_11842,N_5016,N_5194);
xor U11843 (N_11843,N_9445,N_6454);
nand U11844 (N_11844,N_6258,N_5126);
or U11845 (N_11845,N_5735,N_8928);
nand U11846 (N_11846,N_8379,N_5375);
nor U11847 (N_11847,N_6954,N_6857);
nor U11848 (N_11848,N_7269,N_9692);
or U11849 (N_11849,N_8276,N_7498);
xnor U11850 (N_11850,N_8000,N_9978);
nor U11851 (N_11851,N_7637,N_8987);
nor U11852 (N_11852,N_5437,N_9323);
or U11853 (N_11853,N_9365,N_8484);
nor U11854 (N_11854,N_5190,N_7918);
or U11855 (N_11855,N_6538,N_5518);
xnor U11856 (N_11856,N_9587,N_9655);
xnor U11857 (N_11857,N_8368,N_9218);
or U11858 (N_11858,N_7458,N_8940);
or U11859 (N_11859,N_9236,N_6191);
xor U11860 (N_11860,N_9367,N_9268);
or U11861 (N_11861,N_5870,N_8568);
and U11862 (N_11862,N_7643,N_7420);
and U11863 (N_11863,N_9762,N_8856);
and U11864 (N_11864,N_6390,N_9713);
nor U11865 (N_11865,N_9369,N_6937);
nor U11866 (N_11866,N_9364,N_5568);
nor U11867 (N_11867,N_5503,N_9678);
nand U11868 (N_11868,N_6898,N_7455);
nor U11869 (N_11869,N_9686,N_6166);
nand U11870 (N_11870,N_9741,N_5168);
xor U11871 (N_11871,N_9299,N_5188);
and U11872 (N_11872,N_6131,N_7356);
xor U11873 (N_11873,N_8072,N_8883);
xnor U11874 (N_11874,N_9248,N_6866);
nand U11875 (N_11875,N_5632,N_9295);
and U11876 (N_11876,N_9521,N_6167);
nor U11877 (N_11877,N_8681,N_7543);
xnor U11878 (N_11878,N_7678,N_8275);
and U11879 (N_11879,N_6827,N_5523);
nor U11880 (N_11880,N_5414,N_9539);
or U11881 (N_11881,N_6750,N_5703);
xnor U11882 (N_11882,N_8257,N_7995);
nor U11883 (N_11883,N_9481,N_8761);
nand U11884 (N_11884,N_6073,N_7757);
or U11885 (N_11885,N_9511,N_6367);
and U11886 (N_11886,N_6989,N_7312);
and U11887 (N_11887,N_7897,N_7169);
xor U11888 (N_11888,N_9051,N_9366);
nand U11889 (N_11889,N_5704,N_6839);
nor U11890 (N_11890,N_5557,N_7135);
nor U11891 (N_11891,N_5248,N_6114);
and U11892 (N_11892,N_8925,N_8408);
xor U11893 (N_11893,N_6906,N_6316);
or U11894 (N_11894,N_9338,N_6075);
and U11895 (N_11895,N_7027,N_7313);
nor U11896 (N_11896,N_5577,N_7268);
and U11897 (N_11897,N_8085,N_9160);
nand U11898 (N_11898,N_7227,N_7521);
or U11899 (N_11899,N_5491,N_9356);
or U11900 (N_11900,N_5992,N_7416);
or U11901 (N_11901,N_6327,N_5500);
or U11902 (N_11902,N_9100,N_6254);
xor U11903 (N_11903,N_7879,N_8823);
nor U11904 (N_11904,N_9206,N_6182);
or U11905 (N_11905,N_6860,N_8915);
xor U11906 (N_11906,N_8222,N_6253);
nor U11907 (N_11907,N_5400,N_8512);
and U11908 (N_11908,N_9528,N_9764);
nand U11909 (N_11909,N_6234,N_8802);
nand U11910 (N_11910,N_7141,N_5674);
and U11911 (N_11911,N_6529,N_9380);
or U11912 (N_11912,N_9093,N_9430);
or U11913 (N_11913,N_5781,N_5753);
nor U11914 (N_11914,N_5243,N_7626);
or U11915 (N_11915,N_8016,N_8772);
and U11916 (N_11916,N_9886,N_6459);
nand U11917 (N_11917,N_6037,N_5675);
and U11918 (N_11918,N_5710,N_6092);
nor U11919 (N_11919,N_7189,N_7607);
nand U11920 (N_11920,N_5857,N_6235);
nand U11921 (N_11921,N_7877,N_6701);
xor U11922 (N_11922,N_6542,N_6757);
nor U11923 (N_11923,N_5070,N_6723);
and U11924 (N_11924,N_7662,N_7435);
nor U11925 (N_11925,N_6511,N_7570);
or U11926 (N_11926,N_9154,N_7346);
nand U11927 (N_11927,N_5633,N_8678);
nor U11928 (N_11928,N_8091,N_5747);
nand U11929 (N_11929,N_6781,N_6753);
nand U11930 (N_11930,N_9724,N_6419);
nor U11931 (N_11931,N_7824,N_5582);
xor U11932 (N_11932,N_8553,N_5634);
or U11933 (N_11933,N_6201,N_5664);
xor U11934 (N_11934,N_6395,N_8985);
or U11935 (N_11935,N_9373,N_6694);
or U11936 (N_11936,N_8363,N_7675);
nand U11937 (N_11937,N_7290,N_7378);
xnor U11938 (N_11938,N_7257,N_9574);
nor U11939 (N_11939,N_5961,N_9914);
nor U11940 (N_11940,N_8493,N_7011);
or U11941 (N_11941,N_5428,N_5785);
nor U11942 (N_11942,N_6611,N_9531);
and U11943 (N_11943,N_5230,N_9944);
and U11944 (N_11944,N_8297,N_5379);
and U11945 (N_11945,N_7580,N_6481);
and U11946 (N_11946,N_7051,N_6409);
and U11947 (N_11947,N_9950,N_5748);
or U11948 (N_11948,N_9376,N_7253);
nand U11949 (N_11949,N_7793,N_8254);
nand U11950 (N_11950,N_7177,N_7295);
nor U11951 (N_11951,N_7411,N_9768);
xnor U11952 (N_11952,N_8109,N_5081);
nor U11953 (N_11953,N_7410,N_5451);
nor U11954 (N_11954,N_8033,N_8344);
nand U11955 (N_11955,N_9300,N_8783);
nand U11956 (N_11956,N_6083,N_5438);
xnor U11957 (N_11957,N_6482,N_6099);
xnor U11958 (N_11958,N_5498,N_7638);
and U11959 (N_11959,N_7888,N_5356);
nand U11960 (N_11960,N_6577,N_6098);
nor U11961 (N_11961,N_9326,N_5651);
nand U11962 (N_11962,N_8571,N_9470);
nor U11963 (N_11963,N_9551,N_8353);
xnor U11964 (N_11964,N_6383,N_6863);
nor U11965 (N_11965,N_5221,N_5179);
xnor U11966 (N_11966,N_5876,N_9800);
xor U11967 (N_11967,N_5118,N_5164);
nand U11968 (N_11968,N_5325,N_6478);
nand U11969 (N_11969,N_7719,N_8080);
nand U11970 (N_11970,N_9501,N_5948);
xor U11971 (N_11971,N_5360,N_6086);
and U11972 (N_11972,N_5050,N_6930);
nor U11973 (N_11973,N_7385,N_8826);
xor U11974 (N_11974,N_5636,N_6194);
and U11975 (N_11975,N_7294,N_9657);
nand U11976 (N_11976,N_6815,N_8583);
nand U11977 (N_11977,N_8851,N_7072);
and U11978 (N_11978,N_6916,N_5738);
or U11979 (N_11979,N_6584,N_5996);
xnor U11980 (N_11980,N_5329,N_6302);
nand U11981 (N_11981,N_5309,N_5397);
nand U11982 (N_11982,N_6282,N_9900);
or U11983 (N_11983,N_9221,N_9190);
xnor U11984 (N_11984,N_6566,N_9057);
or U11985 (N_11985,N_6263,N_9028);
and U11986 (N_11986,N_6205,N_6050);
and U11987 (N_11987,N_7326,N_9421);
and U11988 (N_11988,N_8548,N_6187);
or U11989 (N_11989,N_6506,N_8113);
nand U11990 (N_11990,N_7172,N_7933);
and U11991 (N_11991,N_8696,N_9712);
nand U11992 (N_11992,N_7712,N_9496);
or U11993 (N_11993,N_7680,N_5003);
nor U11994 (N_11994,N_7207,N_7608);
and U11995 (N_11995,N_7350,N_8001);
nor U11996 (N_11996,N_7769,N_9606);
and U11997 (N_11997,N_8741,N_8332);
or U11998 (N_11998,N_5598,N_7231);
xor U11999 (N_11999,N_8052,N_6798);
nand U12000 (N_12000,N_6307,N_6222);
or U12001 (N_12001,N_6565,N_7852);
or U12002 (N_12002,N_6198,N_6944);
and U12003 (N_12003,N_6844,N_9856);
xor U12004 (N_12004,N_8365,N_6575);
or U12005 (N_12005,N_6381,N_7480);
and U12006 (N_12006,N_9095,N_7844);
xor U12007 (N_12007,N_9704,N_7928);
nand U12008 (N_12008,N_5290,N_5990);
and U12009 (N_12009,N_5066,N_6784);
and U12010 (N_12010,N_9961,N_8793);
xnor U12011 (N_12011,N_8791,N_5142);
nor U12012 (N_12012,N_5416,N_9964);
or U12013 (N_12013,N_7535,N_8648);
or U12014 (N_12014,N_7444,N_6451);
nand U12015 (N_12015,N_8157,N_5117);
and U12016 (N_12016,N_7264,N_7571);
or U12017 (N_12017,N_8748,N_6500);
nor U12018 (N_12018,N_5222,N_9877);
and U12019 (N_12019,N_6680,N_6679);
or U12020 (N_12020,N_9083,N_8271);
and U12021 (N_12021,N_5826,N_9490);
nor U12022 (N_12022,N_5457,N_9408);
or U12023 (N_12023,N_9993,N_9399);
and U12024 (N_12024,N_5901,N_6036);
and U12025 (N_12025,N_5852,N_8002);
nand U12026 (N_12026,N_7513,N_7136);
nor U12027 (N_12027,N_8871,N_7727);
and U12028 (N_12028,N_6548,N_7641);
and U12029 (N_12029,N_8986,N_6259);
nor U12030 (N_12030,N_7451,N_5912);
nand U12031 (N_12031,N_5550,N_6861);
or U12032 (N_12032,N_9817,N_8710);
nand U12033 (N_12033,N_6747,N_9949);
and U12034 (N_12034,N_5517,N_7988);
xor U12035 (N_12035,N_7503,N_5698);
or U12036 (N_12036,N_9658,N_8449);
or U12037 (N_12037,N_5709,N_5715);
nor U12038 (N_12038,N_7118,N_8766);
nand U12039 (N_12039,N_7471,N_8014);
nor U12040 (N_12040,N_7934,N_6660);
or U12041 (N_12041,N_6243,N_5192);
or U12042 (N_12042,N_7733,N_9553);
and U12043 (N_12043,N_5212,N_5396);
xor U12044 (N_12044,N_6699,N_5646);
and U12045 (N_12045,N_9849,N_7753);
and U12046 (N_12046,N_7799,N_6671);
xnor U12047 (N_12047,N_8653,N_9952);
xor U12048 (N_12048,N_7635,N_9500);
xnor U12049 (N_12049,N_7841,N_9177);
and U12050 (N_12050,N_5524,N_8312);
and U12051 (N_12051,N_9828,N_7873);
and U12052 (N_12052,N_7222,N_9599);
nor U12053 (N_12053,N_7627,N_9419);
nor U12054 (N_12054,N_9770,N_6695);
xor U12055 (N_12055,N_8305,N_8511);
or U12056 (N_12056,N_6601,N_5955);
and U12057 (N_12057,N_6484,N_6371);
and U12058 (N_12058,N_6567,N_6959);
xnor U12059 (N_12059,N_7098,N_7255);
and U12060 (N_12060,N_8650,N_7926);
xor U12061 (N_12061,N_5865,N_6202);
nor U12062 (N_12062,N_5171,N_9935);
nand U12063 (N_12063,N_6583,N_9246);
or U12064 (N_12064,N_7883,N_8041);
or U12065 (N_12065,N_8238,N_5744);
nand U12066 (N_12066,N_9320,N_9231);
and U12067 (N_12067,N_5423,N_8600);
xor U12068 (N_12068,N_5082,N_9695);
or U12069 (N_12069,N_6377,N_5019);
nand U12070 (N_12070,N_6196,N_8464);
nand U12071 (N_12071,N_8359,N_8838);
or U12072 (N_12072,N_7082,N_8727);
xnor U12073 (N_12073,N_6384,N_7889);
or U12074 (N_12074,N_8887,N_7715);
nor U12075 (N_12075,N_5779,N_8824);
or U12076 (N_12076,N_8298,N_6681);
nand U12077 (N_12077,N_8009,N_7710);
and U12078 (N_12078,N_7771,N_8435);
xnor U12079 (N_12079,N_7997,N_9596);
or U12080 (N_12080,N_9079,N_9148);
nand U12081 (N_12081,N_9677,N_5108);
nand U12082 (N_12082,N_5241,N_6498);
nand U12083 (N_12083,N_7589,N_5531);
xnor U12084 (N_12084,N_8151,N_7611);
or U12085 (N_12085,N_8465,N_5089);
nand U12086 (N_12086,N_6740,N_8108);
xor U12087 (N_12087,N_5800,N_9460);
or U12088 (N_12088,N_8030,N_5806);
nor U12089 (N_12089,N_5765,N_7324);
nor U12090 (N_12090,N_5974,N_8422);
nor U12091 (N_12091,N_6225,N_8525);
and U12092 (N_12092,N_5477,N_6402);
nor U12093 (N_12093,N_6976,N_5581);
nand U12094 (N_12094,N_5018,N_9699);
nand U12095 (N_12095,N_7849,N_7415);
nand U12096 (N_12096,N_5610,N_8852);
or U12097 (N_12097,N_9583,N_6434);
and U12098 (N_12098,N_8945,N_9014);
nand U12099 (N_12099,N_5337,N_7650);
or U12100 (N_12100,N_6624,N_5515);
nand U12101 (N_12101,N_8143,N_6009);
xnor U12102 (N_12102,N_7247,N_5648);
or U12103 (N_12103,N_5087,N_6563);
xor U12104 (N_12104,N_8535,N_8156);
nand U12105 (N_12105,N_6056,N_8221);
nor U12106 (N_12106,N_7494,N_7699);
nor U12107 (N_12107,N_6835,N_6674);
and U12108 (N_12108,N_7732,N_8747);
or U12109 (N_12109,N_8311,N_6615);
xnor U12110 (N_12110,N_8237,N_7692);
or U12111 (N_12111,N_7701,N_6228);
or U12112 (N_12112,N_9835,N_8705);
or U12113 (N_12113,N_8081,N_9407);
nor U12114 (N_12114,N_7651,N_8083);
or U12115 (N_12115,N_9747,N_9038);
nor U12116 (N_12116,N_8981,N_5306);
nor U12117 (N_12117,N_8055,N_6233);
or U12118 (N_12118,N_5073,N_6113);
xnor U12119 (N_12119,N_9895,N_5460);
xor U12120 (N_12120,N_9059,N_7705);
or U12121 (N_12121,N_5268,N_6908);
or U12122 (N_12122,N_5441,N_6313);
or U12123 (N_12123,N_9916,N_7828);
nand U12124 (N_12124,N_7861,N_5618);
xnor U12125 (N_12125,N_7121,N_5156);
nor U12126 (N_12126,N_5270,N_7375);
and U12127 (N_12127,N_6817,N_8717);
xnor U12128 (N_12128,N_8035,N_9385);
xor U12129 (N_12129,N_5469,N_8828);
or U12130 (N_12130,N_8533,N_7653);
nand U12131 (N_12131,N_8428,N_8061);
and U12132 (N_12132,N_9778,N_5534);
or U12133 (N_12133,N_8588,N_7276);
or U12134 (N_12134,N_6626,N_7234);
or U12135 (N_12135,N_6715,N_6291);
nor U12136 (N_12136,N_7782,N_5609);
and U12137 (N_12137,N_6435,N_7807);
nand U12138 (N_12138,N_8200,N_7628);
and U12139 (N_12139,N_6241,N_5650);
and U12140 (N_12140,N_5656,N_7763);
nand U12141 (N_12141,N_8900,N_6174);
and U12142 (N_12142,N_6456,N_9495);
nor U12143 (N_12143,N_9267,N_6819);
nor U12144 (N_12144,N_7440,N_8902);
nor U12145 (N_12145,N_8835,N_9464);
and U12146 (N_12146,N_6650,N_7805);
nor U12147 (N_12147,N_9825,N_8691);
or U12148 (N_12148,N_9927,N_9977);
or U12149 (N_12149,N_8787,N_8699);
nand U12150 (N_12150,N_9322,N_6652);
nand U12151 (N_12151,N_7003,N_8418);
nand U12152 (N_12152,N_9736,N_9476);
and U12153 (N_12153,N_6539,N_8573);
and U12154 (N_12154,N_6919,N_6266);
and U12155 (N_12155,N_9237,N_6428);
xnor U12156 (N_12156,N_5317,N_9843);
nor U12157 (N_12157,N_7725,N_7646);
and U12158 (N_12158,N_7633,N_8800);
and U12159 (N_12159,N_9844,N_8652);
nand U12160 (N_12160,N_5526,N_8034);
nand U12161 (N_12161,N_7190,N_7363);
nand U12162 (N_12162,N_6195,N_7142);
xor U12163 (N_12163,N_6595,N_6378);
or U12164 (N_12164,N_9401,N_5572);
nand U12165 (N_12165,N_8361,N_8058);
and U12166 (N_12166,N_9054,N_6293);
or U12167 (N_12167,N_6221,N_8780);
xor U12168 (N_12168,N_7258,N_6598);
or U12169 (N_12169,N_7598,N_7336);
nor U12170 (N_12170,N_8391,N_8068);
nand U12171 (N_12171,N_8606,N_6658);
or U12172 (N_12172,N_6534,N_8322);
xnor U12173 (N_12173,N_6231,N_9516);
or U12174 (N_12174,N_6587,N_5844);
nand U12175 (N_12175,N_7031,N_8709);
or U12176 (N_12176,N_7292,N_9929);
or U12177 (N_12177,N_7280,N_5021);
xnor U12178 (N_12178,N_7559,N_8997);
xor U12179 (N_12179,N_6698,N_6997);
and U12180 (N_12180,N_8526,N_8664);
nor U12181 (N_12181,N_7331,N_7853);
nor U12182 (N_12182,N_6999,N_6364);
nor U12183 (N_12183,N_7647,N_9826);
nor U12184 (N_12184,N_9041,N_5419);
nand U12185 (N_12185,N_9034,N_6623);
nor U12186 (N_12186,N_5311,N_8357);
and U12187 (N_12187,N_7709,N_6711);
nor U12188 (N_12188,N_6547,N_6579);
nor U12189 (N_12189,N_9112,N_7038);
xnor U12190 (N_12190,N_9355,N_7909);
and U12191 (N_12191,N_5011,N_9906);
nand U12192 (N_12192,N_7700,N_7837);
xor U12193 (N_12193,N_6517,N_9615);
nor U12194 (N_12194,N_7173,N_5600);
or U12195 (N_12195,N_9510,N_9904);
xor U12196 (N_12196,N_9099,N_6880);
nand U12197 (N_12197,N_5939,N_8636);
nor U12198 (N_12198,N_6772,N_6357);
or U12199 (N_12199,N_7001,N_5304);
and U12200 (N_12200,N_9975,N_9291);
xor U12201 (N_12201,N_5787,N_9310);
xor U12202 (N_12202,N_8022,N_7398);
nor U12203 (N_12203,N_7946,N_9603);
nand U12204 (N_12204,N_7094,N_9722);
nand U12205 (N_12205,N_7359,N_8735);
xor U12206 (N_12206,N_9685,N_9943);
xnor U12207 (N_12207,N_7887,N_9011);
xnor U12208 (N_12208,N_5291,N_7542);
and U12209 (N_12209,N_5276,N_9998);
xor U12210 (N_12210,N_8899,N_8381);
and U12211 (N_12211,N_9889,N_9313);
or U12212 (N_12212,N_7931,N_9077);
nor U12213 (N_12213,N_5662,N_6722);
xnor U12214 (N_12214,N_9853,N_6910);
nor U12215 (N_12215,N_5446,N_5014);
xnor U12216 (N_12216,N_9377,N_5809);
or U12217 (N_12217,N_6126,N_6800);
xnor U12218 (N_12218,N_5642,N_5822);
nor U12219 (N_12219,N_7113,N_8502);
nand U12220 (N_12220,N_7250,N_7485);
and U12221 (N_12221,N_8843,N_9957);
or U12222 (N_12222,N_6470,N_7092);
or U12223 (N_12223,N_5159,N_7630);
and U12224 (N_12224,N_7270,N_7060);
xnor U12225 (N_12225,N_7376,N_9976);
nand U12226 (N_12226,N_5788,N_8528);
nor U12227 (N_12227,N_8803,N_8519);
and U12228 (N_12228,N_7587,N_8390);
or U12229 (N_12229,N_5434,N_9193);
nor U12230 (N_12230,N_7417,N_7514);
and U12231 (N_12231,N_8630,N_9480);
or U12232 (N_12232,N_9053,N_7905);
and U12233 (N_12233,N_5655,N_5275);
or U12234 (N_12234,N_9308,N_9127);
nor U12235 (N_12235,N_5832,N_6403);
xor U12236 (N_12236,N_6389,N_8878);
or U12237 (N_12237,N_6352,N_8560);
nand U12238 (N_12238,N_8167,N_5979);
nand U12239 (N_12239,N_8759,N_6169);
nand U12240 (N_12240,N_5382,N_8048);
or U12241 (N_12241,N_5436,N_5131);
nand U12242 (N_12242,N_5778,N_6637);
and U12243 (N_12243,N_8473,N_9433);
or U12244 (N_12244,N_7815,N_6424);
and U12245 (N_12245,N_5931,N_9992);
nand U12246 (N_12246,N_7064,N_6065);
nand U12247 (N_12247,N_7657,N_6570);
and U12248 (N_12248,N_8950,N_7319);
and U12249 (N_12249,N_8861,N_8310);
nor U12250 (N_12250,N_6387,N_6692);
xor U12251 (N_12251,N_6064,N_7228);
nand U12252 (N_12252,N_6810,N_8105);
nand U12253 (N_12253,N_8999,N_8607);
nor U12254 (N_12254,N_9932,N_9709);
and U12255 (N_12255,N_5130,N_7493);
and U12256 (N_12256,N_7808,N_5924);
and U12257 (N_12257,N_6336,N_8857);
nand U12258 (N_12258,N_9273,N_7533);
nor U12259 (N_12259,N_8660,N_9140);
xor U12260 (N_12260,N_9024,N_9812);
nand U12261 (N_12261,N_9105,N_9351);
or U12262 (N_12262,N_5746,N_5468);
nand U12263 (N_12263,N_5701,N_6161);
and U12264 (N_12264,N_9693,N_8188);
nand U12265 (N_12265,N_5667,N_5889);
and U12266 (N_12266,N_9742,N_8827);
or U12267 (N_12267,N_9602,N_8046);
xor U12268 (N_12268,N_5914,N_9184);
nor U12269 (N_12269,N_9862,N_8330);
and U12270 (N_12270,N_7639,N_9208);
xnor U12271 (N_12271,N_6670,N_7010);
nor U12272 (N_12272,N_6262,N_6589);
and U12273 (N_12273,N_8126,N_7186);
or U12274 (N_12274,N_5668,N_9217);
or U12275 (N_12275,N_6597,N_5930);
and U12276 (N_12276,N_5756,N_5466);
nand U12277 (N_12277,N_7370,N_8443);
nand U12278 (N_12278,N_8094,N_8148);
nand U12279 (N_12279,N_8106,N_5611);
and U12280 (N_12280,N_6429,N_6628);
nor U12281 (N_12281,N_8724,N_7527);
xnor U12282 (N_12282,N_8392,N_7492);
or U12283 (N_12283,N_8279,N_7617);
xor U12284 (N_12284,N_5218,N_7408);
and U12285 (N_12285,N_7751,N_7908);
nor U12286 (N_12286,N_5055,N_7973);
nor U12287 (N_12287,N_6530,N_6024);
or U12288 (N_12288,N_9665,N_6226);
or U12289 (N_12289,N_5348,N_7954);
nor U12290 (N_12290,N_7205,N_5049);
nor U12291 (N_12291,N_7457,N_9598);
nand U12292 (N_12292,N_7338,N_9560);
nand U12293 (N_12293,N_7341,N_9181);
nand U12294 (N_12294,N_9509,N_9614);
and U12295 (N_12295,N_9343,N_5982);
nand U12296 (N_12296,N_6423,N_7490);
xor U12297 (N_12297,N_8858,N_6477);
and U12298 (N_12298,N_5252,N_9494);
or U12299 (N_12299,N_7652,N_6963);
or U12300 (N_12300,N_8884,N_8317);
nand U12301 (N_12301,N_7238,N_7036);
or U12302 (N_12302,N_5652,N_9265);
or U12303 (N_12303,N_7384,N_9808);
nand U12304 (N_12304,N_7561,N_9915);
nor U12305 (N_12305,N_7130,N_7544);
nand U12306 (N_12306,N_5846,N_8711);
nor U12307 (N_12307,N_5100,N_6223);
nor U12308 (N_12308,N_6458,N_7670);
or U12309 (N_12309,N_9497,N_5380);
or U12310 (N_12310,N_6947,N_6046);
nor U12311 (N_12311,N_9882,N_5907);
xor U12312 (N_12312,N_8186,N_8882);
and U12313 (N_12313,N_9279,N_6546);
nand U12314 (N_12314,N_8966,N_5533);
or U12315 (N_12315,N_7325,N_7215);
nor U12316 (N_12316,N_5432,N_9293);
or U12317 (N_12317,N_6047,N_5657);
and U12318 (N_12318,N_7655,N_9910);
xnor U12319 (N_12319,N_7448,N_6373);
nor U12320 (N_12320,N_9423,N_5956);
nor U12321 (N_12321,N_5983,N_7022);
or U12322 (N_12322,N_8903,N_7266);
nand U12323 (N_12323,N_9585,N_7002);
or U12324 (N_12324,N_6807,N_6627);
nand U12325 (N_12325,N_9881,N_5265);
nor U12326 (N_12326,N_7000,N_7499);
nor U12327 (N_12327,N_5998,N_6518);
nor U12328 (N_12328,N_5346,N_9005);
nand U12329 (N_12329,N_9280,N_9179);
xor U12330 (N_12330,N_6321,N_6640);
nand U12331 (N_12331,N_9379,N_9865);
nand U12332 (N_12332,N_7214,N_7825);
or U12333 (N_12333,N_5775,N_8129);
xnor U12334 (N_12334,N_5608,N_9854);
nand U12335 (N_12335,N_5696,N_7301);
or U12336 (N_12336,N_9951,N_5942);
xor U12337 (N_12337,N_5299,N_9921);
nor U12338 (N_12338,N_9787,N_5986);
xnor U12339 (N_12339,N_6713,N_5057);
nand U12340 (N_12340,N_7501,N_6610);
or U12341 (N_12341,N_7930,N_8174);
nand U12342 (N_12342,N_5051,N_5566);
and U12343 (N_12343,N_6665,N_8333);
and U12344 (N_12344,N_8758,N_9185);
nand U12345 (N_12345,N_5720,N_7373);
xnor U12346 (N_12346,N_7465,N_5124);
or U12347 (N_12347,N_5909,N_6887);
xor U12348 (N_12348,N_6504,N_8329);
nor U12349 (N_12349,N_8968,N_8734);
and U12350 (N_12350,N_5626,N_6496);
or U12351 (N_12351,N_5206,N_6706);
xor U12352 (N_12352,N_7854,N_7055);
nor U12353 (N_12353,N_5867,N_8441);
xor U12354 (N_12354,N_5213,N_6347);
nand U12355 (N_12355,N_6400,N_6853);
and U12356 (N_12356,N_8403,N_9037);
xor U12357 (N_12357,N_7511,N_8220);
nand U12358 (N_12358,N_7576,N_6468);
nor U12359 (N_12359,N_7080,N_9506);
nand U12360 (N_12360,N_6978,N_8703);
nor U12361 (N_12361,N_7422,N_9168);
nor U12362 (N_12362,N_9743,N_5820);
or U12363 (N_12363,N_8608,N_8814);
nor U12364 (N_12364,N_6521,N_9637);
nand U12365 (N_12365,N_5980,N_5601);
xnor U12366 (N_12366,N_9535,N_8834);
xor U12367 (N_12367,N_7477,N_8888);
xor U12368 (N_12368,N_8808,N_8561);
xor U12369 (N_12369,N_5114,N_6550);
xnor U12370 (N_12370,N_8566,N_9766);
nand U12371 (N_12371,N_8267,N_6700);
nor U12372 (N_12372,N_8744,N_7272);
nor U12373 (N_12373,N_6328,N_6830);
nor U12374 (N_12374,N_5173,N_5385);
or U12375 (N_12375,N_7497,N_8536);
nand U12376 (N_12376,N_6447,N_5561);
nor U12377 (N_12377,N_6858,N_6172);
nor U12378 (N_12378,N_7661,N_5843);
and U12379 (N_12379,N_5075,N_7856);
and U12380 (N_12380,N_9392,N_8556);
and U12381 (N_12381,N_6661,N_9570);
and U12382 (N_12382,N_5429,N_9991);
nand U12383 (N_12383,N_5044,N_6252);
or U12384 (N_12384,N_9586,N_8904);
xor U12385 (N_12385,N_5927,N_7433);
nor U12386 (N_12386,N_9492,N_5815);
nor U12387 (N_12387,N_8459,N_7306);
or U12388 (N_12388,N_9649,N_6480);
nand U12389 (N_12389,N_5541,N_5293);
and U12390 (N_12390,N_8782,N_6846);
xnor U12391 (N_12391,N_8819,N_8621);
xnor U12392 (N_12392,N_6333,N_8038);
or U12393 (N_12393,N_8506,N_5952);
and U12394 (N_12394,N_9357,N_9003);
nor U12395 (N_12395,N_8062,N_6573);
or U12396 (N_12396,N_5790,N_5420);
nand U12397 (N_12397,N_5240,N_8050);
or U12398 (N_12398,N_5895,N_8746);
and U12399 (N_12399,N_7983,N_8751);
xor U12400 (N_12400,N_9283,N_7233);
or U12401 (N_12401,N_9995,N_5085);
nor U12402 (N_12402,N_8326,N_5281);
nor U12403 (N_12403,N_6659,N_5959);
or U12404 (N_12404,N_8070,N_6117);
nor U12405 (N_12405,N_7240,N_7116);
nand U12406 (N_12406,N_9801,N_7814);
nand U12407 (N_12407,N_7858,N_8162);
and U12408 (N_12408,N_7966,N_7528);
xor U12409 (N_12409,N_9792,N_7764);
xnor U12410 (N_12410,N_5200,N_8023);
xor U12411 (N_12411,N_6966,N_7419);
and U12412 (N_12412,N_7649,N_9752);
nor U12413 (N_12413,N_5269,N_9156);
and U12414 (N_12414,N_9972,N_9115);
xor U12415 (N_12415,N_7124,N_5725);
or U12416 (N_12416,N_9085,N_7717);
and U12417 (N_12417,N_8637,N_5197);
nor U12418 (N_12418,N_6465,N_6063);
nor U12419 (N_12419,N_9515,N_8277);
xnor U12420 (N_12420,N_5670,N_8112);
nor U12421 (N_12421,N_9651,N_5592);
xnor U12422 (N_12422,N_8491,N_9001);
nor U12423 (N_12423,N_8582,N_9671);
and U12424 (N_12424,N_6103,N_7251);
nand U12425 (N_12425,N_9439,N_8920);
nand U12426 (N_12426,N_8467,N_9225);
nor U12427 (N_12427,N_5805,N_8153);
or U12428 (N_12428,N_6027,N_6033);
and U12429 (N_12429,N_5560,N_8399);
and U12430 (N_12430,N_8029,N_5461);
xnor U12431 (N_12431,N_5102,N_8207);
xor U12432 (N_12432,N_5866,N_7541);
nor U12433 (N_12433,N_7857,N_5617);
or U12434 (N_12434,N_8943,N_5040);
xor U12435 (N_12435,N_5112,N_6148);
or U12436 (N_12436,N_9922,N_9416);
or U12437 (N_12437,N_5334,N_8931);
or U12438 (N_12438,N_9662,N_8895);
nor U12439 (N_12439,N_6696,N_7669);
and U12440 (N_12440,N_8570,N_9425);
or U12441 (N_12441,N_6163,N_8730);
nand U12442 (N_12442,N_6385,N_9549);
nand U12443 (N_12443,N_9137,N_7311);
nand U12444 (N_12444,N_7024,N_5796);
xnor U12445 (N_12445,N_6791,N_8914);
nor U12446 (N_12446,N_5048,N_9584);
xor U12447 (N_12447,N_6585,N_9201);
and U12448 (N_12448,N_7046,N_9241);
and U12449 (N_12449,N_8388,N_9708);
and U12450 (N_12450,N_9463,N_6144);
nand U12451 (N_12451,N_5158,N_7802);
xnor U12452 (N_12452,N_8969,N_5519);
nand U12453 (N_12453,N_5189,N_5695);
nand U12454 (N_12454,N_6755,N_9912);
nor U12455 (N_12455,N_6691,N_6655);
nor U12456 (N_12456,N_6669,N_5373);
nand U12457 (N_12457,N_7327,N_6361);
nand U12458 (N_12458,N_5923,N_8395);
and U12459 (N_12459,N_8517,N_5408);
nor U12460 (N_12460,N_7616,N_7980);
nand U12461 (N_12461,N_5067,N_7947);
nand U12462 (N_12462,N_6120,N_6657);
nand U12463 (N_12463,N_9136,N_5101);
xnor U12464 (N_12464,N_9315,N_9774);
xor U12465 (N_12465,N_5851,N_8926);
nand U12466 (N_12466,N_7277,N_6576);
or U12467 (N_12467,N_9186,N_8291);
nor U12468 (N_12468,N_5362,N_7379);
or U12469 (N_12469,N_5232,N_6822);
nand U12470 (N_12470,N_6299,N_5894);
xnor U12471 (N_12471,N_8026,N_5006);
nand U12472 (N_12472,N_5813,N_8967);
and U12473 (N_12473,N_9027,N_8018);
nor U12474 (N_12474,N_6404,N_9833);
nor U12475 (N_12475,N_9969,N_9026);
and U12476 (N_12476,N_9292,N_8849);
nor U12477 (N_12477,N_9760,N_8100);
nand U12478 (N_12478,N_6786,N_7291);
and U12479 (N_12479,N_5888,N_7981);
nor U12480 (N_12480,N_6139,N_7689);
nand U12481 (N_12481,N_7208,N_8178);
and U12482 (N_12482,N_7823,N_8280);
nand U12483 (N_12483,N_9771,N_8537);
nor U12484 (N_12484,N_5567,N_7237);
and U12485 (N_12485,N_5649,N_9092);
nor U12486 (N_12486,N_7084,N_5326);
nand U12487 (N_12487,N_6190,N_9233);
or U12488 (N_12488,N_8971,N_5879);
nor U12489 (N_12489,N_8173,N_9469);
nand U12490 (N_12490,N_9162,N_8794);
xor U12491 (N_12491,N_5532,N_8992);
nand U12492 (N_12492,N_7582,N_5459);
and U12493 (N_12493,N_6831,N_8331);
or U12494 (N_12494,N_6326,N_7602);
or U12495 (N_12495,N_5310,N_8850);
xnor U12496 (N_12496,N_5002,N_7216);
nor U12497 (N_12497,N_7279,N_8397);
and U12498 (N_12498,N_7978,N_8201);
nand U12499 (N_12499,N_6211,N_9887);
xnor U12500 (N_12500,N_8784,N_9182);
nor U12501 (N_12501,N_7054,N_6907);
and U12502 (N_12502,N_7700,N_9243);
nand U12503 (N_12503,N_5222,N_7087);
nand U12504 (N_12504,N_9053,N_9496);
and U12505 (N_12505,N_5304,N_8037);
nand U12506 (N_12506,N_7172,N_9054);
nand U12507 (N_12507,N_7287,N_9889);
nor U12508 (N_12508,N_6257,N_6884);
and U12509 (N_12509,N_7572,N_6106);
and U12510 (N_12510,N_9986,N_6994);
and U12511 (N_12511,N_7749,N_8479);
nor U12512 (N_12512,N_7211,N_6946);
or U12513 (N_12513,N_7784,N_8151);
nor U12514 (N_12514,N_7073,N_6336);
xor U12515 (N_12515,N_7313,N_6890);
nand U12516 (N_12516,N_5226,N_5630);
or U12517 (N_12517,N_8588,N_9642);
xor U12518 (N_12518,N_8652,N_6380);
and U12519 (N_12519,N_8604,N_8984);
and U12520 (N_12520,N_9150,N_6280);
xnor U12521 (N_12521,N_8529,N_7955);
nor U12522 (N_12522,N_6138,N_9693);
nand U12523 (N_12523,N_8630,N_8288);
and U12524 (N_12524,N_9563,N_7449);
nand U12525 (N_12525,N_9281,N_7314);
nand U12526 (N_12526,N_9634,N_7753);
and U12527 (N_12527,N_6526,N_5574);
nand U12528 (N_12528,N_9574,N_6255);
nor U12529 (N_12529,N_6282,N_7654);
xnor U12530 (N_12530,N_7804,N_7938);
nor U12531 (N_12531,N_5943,N_6901);
nor U12532 (N_12532,N_7944,N_8735);
xnor U12533 (N_12533,N_5650,N_5335);
and U12534 (N_12534,N_6544,N_6482);
and U12535 (N_12535,N_7009,N_7126);
nor U12536 (N_12536,N_8037,N_7617);
xor U12537 (N_12537,N_9085,N_5781);
or U12538 (N_12538,N_6610,N_5488);
xor U12539 (N_12539,N_8039,N_8498);
xor U12540 (N_12540,N_9140,N_8791);
and U12541 (N_12541,N_5293,N_6210);
or U12542 (N_12542,N_8094,N_6225);
or U12543 (N_12543,N_9592,N_6278);
and U12544 (N_12544,N_5258,N_8439);
and U12545 (N_12545,N_9391,N_9421);
and U12546 (N_12546,N_6948,N_6310);
nand U12547 (N_12547,N_7719,N_6968);
nor U12548 (N_12548,N_8139,N_6862);
nor U12549 (N_12549,N_9789,N_8657);
and U12550 (N_12550,N_7347,N_5132);
nor U12551 (N_12551,N_9075,N_9146);
xnor U12552 (N_12552,N_9787,N_7122);
nor U12553 (N_12553,N_9955,N_7281);
xor U12554 (N_12554,N_5200,N_6339);
and U12555 (N_12555,N_9967,N_8508);
or U12556 (N_12556,N_5131,N_6540);
nand U12557 (N_12557,N_9696,N_5534);
nor U12558 (N_12558,N_9891,N_9616);
nor U12559 (N_12559,N_5921,N_8171);
nor U12560 (N_12560,N_6649,N_5396);
or U12561 (N_12561,N_9767,N_6016);
nor U12562 (N_12562,N_9473,N_7291);
nand U12563 (N_12563,N_7279,N_5281);
or U12564 (N_12564,N_6983,N_7389);
and U12565 (N_12565,N_9506,N_6838);
nor U12566 (N_12566,N_9034,N_5304);
nand U12567 (N_12567,N_5348,N_7475);
nor U12568 (N_12568,N_9694,N_9897);
xnor U12569 (N_12569,N_8974,N_7387);
nand U12570 (N_12570,N_6827,N_9687);
nand U12571 (N_12571,N_6653,N_5407);
nor U12572 (N_12572,N_6108,N_9222);
nand U12573 (N_12573,N_8993,N_6653);
xor U12574 (N_12574,N_8917,N_7801);
or U12575 (N_12575,N_6822,N_9726);
xor U12576 (N_12576,N_7591,N_6353);
xor U12577 (N_12577,N_6745,N_8883);
nor U12578 (N_12578,N_8284,N_5368);
or U12579 (N_12579,N_7614,N_9836);
nor U12580 (N_12580,N_8533,N_6131);
xor U12581 (N_12581,N_8369,N_5635);
or U12582 (N_12582,N_8765,N_5145);
or U12583 (N_12583,N_8349,N_5201);
nand U12584 (N_12584,N_7145,N_7546);
nand U12585 (N_12585,N_7059,N_7822);
nor U12586 (N_12586,N_7090,N_8966);
nor U12587 (N_12587,N_7453,N_8229);
xnor U12588 (N_12588,N_8003,N_9923);
xor U12589 (N_12589,N_8940,N_9512);
and U12590 (N_12590,N_6591,N_9472);
or U12591 (N_12591,N_5828,N_9317);
or U12592 (N_12592,N_5098,N_7113);
xor U12593 (N_12593,N_8111,N_5137);
xor U12594 (N_12594,N_8250,N_8889);
or U12595 (N_12595,N_8521,N_5438);
or U12596 (N_12596,N_7506,N_6729);
xor U12597 (N_12597,N_8619,N_5369);
and U12598 (N_12598,N_6172,N_6595);
nor U12599 (N_12599,N_5258,N_6995);
nand U12600 (N_12600,N_9648,N_7866);
xnor U12601 (N_12601,N_7528,N_8813);
nor U12602 (N_12602,N_8114,N_9118);
xnor U12603 (N_12603,N_6415,N_6340);
and U12604 (N_12604,N_7646,N_6539);
nor U12605 (N_12605,N_7955,N_7969);
or U12606 (N_12606,N_7765,N_5567);
or U12607 (N_12607,N_5264,N_9946);
nand U12608 (N_12608,N_9011,N_5564);
or U12609 (N_12609,N_7611,N_6475);
xnor U12610 (N_12610,N_9884,N_6103);
nor U12611 (N_12611,N_5997,N_9010);
xor U12612 (N_12612,N_8756,N_6041);
xor U12613 (N_12613,N_7678,N_9053);
and U12614 (N_12614,N_6061,N_6483);
and U12615 (N_12615,N_5951,N_8916);
xnor U12616 (N_12616,N_5669,N_9440);
nor U12617 (N_12617,N_8262,N_8423);
nand U12618 (N_12618,N_9813,N_6111);
nor U12619 (N_12619,N_9230,N_8129);
nand U12620 (N_12620,N_6687,N_9103);
nand U12621 (N_12621,N_9067,N_7341);
nand U12622 (N_12622,N_8014,N_8432);
xnor U12623 (N_12623,N_6565,N_5290);
xnor U12624 (N_12624,N_5239,N_5744);
or U12625 (N_12625,N_5595,N_5421);
nor U12626 (N_12626,N_9591,N_8383);
or U12627 (N_12627,N_6188,N_8219);
xnor U12628 (N_12628,N_8598,N_9017);
nand U12629 (N_12629,N_7869,N_5422);
xor U12630 (N_12630,N_5552,N_9256);
xnor U12631 (N_12631,N_5272,N_7913);
nor U12632 (N_12632,N_7012,N_7088);
nand U12633 (N_12633,N_9600,N_5146);
or U12634 (N_12634,N_9949,N_5382);
nand U12635 (N_12635,N_6594,N_5362);
nand U12636 (N_12636,N_7248,N_6767);
and U12637 (N_12637,N_7010,N_8077);
or U12638 (N_12638,N_7825,N_8114);
and U12639 (N_12639,N_8586,N_5706);
nand U12640 (N_12640,N_9972,N_7515);
and U12641 (N_12641,N_5053,N_7195);
xor U12642 (N_12642,N_8683,N_7752);
nand U12643 (N_12643,N_9652,N_6178);
nor U12644 (N_12644,N_8034,N_7030);
or U12645 (N_12645,N_7600,N_9649);
nand U12646 (N_12646,N_7943,N_7812);
nor U12647 (N_12647,N_5805,N_6779);
nor U12648 (N_12648,N_7564,N_6900);
or U12649 (N_12649,N_9498,N_5904);
or U12650 (N_12650,N_9794,N_5292);
xnor U12651 (N_12651,N_8164,N_6120);
nor U12652 (N_12652,N_5250,N_6665);
xnor U12653 (N_12653,N_7636,N_6452);
xor U12654 (N_12654,N_5864,N_6408);
xnor U12655 (N_12655,N_7660,N_7520);
or U12656 (N_12656,N_7955,N_8731);
nor U12657 (N_12657,N_8362,N_8272);
and U12658 (N_12658,N_9744,N_9189);
nor U12659 (N_12659,N_7328,N_6780);
nor U12660 (N_12660,N_5652,N_5168);
nand U12661 (N_12661,N_9006,N_6579);
nor U12662 (N_12662,N_9571,N_5077);
nand U12663 (N_12663,N_5602,N_5312);
and U12664 (N_12664,N_8976,N_9817);
nor U12665 (N_12665,N_8438,N_6699);
xnor U12666 (N_12666,N_5434,N_7442);
and U12667 (N_12667,N_6685,N_6621);
and U12668 (N_12668,N_7902,N_8519);
nor U12669 (N_12669,N_5070,N_6613);
nand U12670 (N_12670,N_8850,N_8180);
or U12671 (N_12671,N_8473,N_8864);
xor U12672 (N_12672,N_6078,N_5164);
nor U12673 (N_12673,N_5401,N_9499);
nand U12674 (N_12674,N_7167,N_8462);
xor U12675 (N_12675,N_9363,N_5074);
xor U12676 (N_12676,N_8382,N_6018);
xnor U12677 (N_12677,N_8205,N_8804);
and U12678 (N_12678,N_5687,N_9397);
nand U12679 (N_12679,N_9835,N_5898);
nor U12680 (N_12680,N_9168,N_8702);
and U12681 (N_12681,N_9311,N_8740);
xnor U12682 (N_12682,N_7133,N_5546);
nand U12683 (N_12683,N_6318,N_7638);
nor U12684 (N_12684,N_9385,N_9442);
nand U12685 (N_12685,N_7599,N_7492);
nand U12686 (N_12686,N_8180,N_6823);
nand U12687 (N_12687,N_6993,N_9519);
or U12688 (N_12688,N_8220,N_9224);
nand U12689 (N_12689,N_9750,N_7977);
or U12690 (N_12690,N_5587,N_7640);
nand U12691 (N_12691,N_7536,N_9982);
xnor U12692 (N_12692,N_5426,N_9675);
xor U12693 (N_12693,N_7038,N_6696);
or U12694 (N_12694,N_9679,N_9639);
nand U12695 (N_12695,N_5560,N_7028);
nand U12696 (N_12696,N_7404,N_5297);
nor U12697 (N_12697,N_7790,N_5878);
nor U12698 (N_12698,N_7943,N_5442);
xor U12699 (N_12699,N_7367,N_8968);
nand U12700 (N_12700,N_8233,N_6659);
xor U12701 (N_12701,N_9843,N_8033);
or U12702 (N_12702,N_5065,N_8305);
and U12703 (N_12703,N_8642,N_8761);
nand U12704 (N_12704,N_9575,N_6445);
nor U12705 (N_12705,N_8898,N_9696);
xor U12706 (N_12706,N_8858,N_7741);
nor U12707 (N_12707,N_9083,N_8083);
nand U12708 (N_12708,N_5188,N_5518);
and U12709 (N_12709,N_6864,N_5666);
nand U12710 (N_12710,N_8772,N_7999);
nor U12711 (N_12711,N_6240,N_6122);
nor U12712 (N_12712,N_9983,N_9516);
xor U12713 (N_12713,N_9715,N_7153);
and U12714 (N_12714,N_7103,N_9721);
or U12715 (N_12715,N_9256,N_6216);
or U12716 (N_12716,N_8794,N_6292);
xnor U12717 (N_12717,N_5505,N_6731);
nor U12718 (N_12718,N_5830,N_5263);
xor U12719 (N_12719,N_6245,N_5156);
nand U12720 (N_12720,N_7692,N_9471);
xnor U12721 (N_12721,N_7632,N_9727);
xnor U12722 (N_12722,N_5270,N_5898);
and U12723 (N_12723,N_7314,N_6845);
nor U12724 (N_12724,N_9014,N_9389);
or U12725 (N_12725,N_9049,N_8081);
nor U12726 (N_12726,N_8058,N_5873);
or U12727 (N_12727,N_6359,N_6218);
and U12728 (N_12728,N_7093,N_7070);
nand U12729 (N_12729,N_9542,N_7114);
xor U12730 (N_12730,N_7641,N_8692);
nand U12731 (N_12731,N_8228,N_6700);
xnor U12732 (N_12732,N_8387,N_7684);
nand U12733 (N_12733,N_5188,N_9488);
xnor U12734 (N_12734,N_9207,N_5012);
or U12735 (N_12735,N_6582,N_8999);
or U12736 (N_12736,N_7324,N_5497);
nor U12737 (N_12737,N_9537,N_7819);
or U12738 (N_12738,N_6608,N_9645);
xor U12739 (N_12739,N_8268,N_6076);
xor U12740 (N_12740,N_6074,N_8911);
nor U12741 (N_12741,N_5655,N_7802);
or U12742 (N_12742,N_5917,N_8397);
xor U12743 (N_12743,N_8026,N_7722);
nand U12744 (N_12744,N_6681,N_5727);
or U12745 (N_12745,N_7670,N_6828);
nand U12746 (N_12746,N_7042,N_7282);
nor U12747 (N_12747,N_6656,N_6267);
and U12748 (N_12748,N_7895,N_6638);
nor U12749 (N_12749,N_7069,N_7775);
xnor U12750 (N_12750,N_5436,N_5646);
xor U12751 (N_12751,N_8542,N_7199);
and U12752 (N_12752,N_9652,N_6141);
and U12753 (N_12753,N_7237,N_9464);
and U12754 (N_12754,N_6051,N_6581);
nand U12755 (N_12755,N_6696,N_6272);
xor U12756 (N_12756,N_9415,N_8514);
nor U12757 (N_12757,N_9266,N_7699);
and U12758 (N_12758,N_7028,N_8620);
or U12759 (N_12759,N_8157,N_9061);
or U12760 (N_12760,N_7269,N_6980);
nand U12761 (N_12761,N_6469,N_7195);
xnor U12762 (N_12762,N_5920,N_7080);
and U12763 (N_12763,N_7263,N_7278);
nand U12764 (N_12764,N_5809,N_7324);
nand U12765 (N_12765,N_7201,N_7168);
or U12766 (N_12766,N_7127,N_6905);
xnor U12767 (N_12767,N_6591,N_9535);
nor U12768 (N_12768,N_6526,N_9963);
nand U12769 (N_12769,N_5396,N_6561);
and U12770 (N_12770,N_6496,N_5202);
xnor U12771 (N_12771,N_9842,N_7935);
and U12772 (N_12772,N_8825,N_5115);
nor U12773 (N_12773,N_6680,N_6006);
nor U12774 (N_12774,N_5600,N_8003);
nand U12775 (N_12775,N_7811,N_5748);
and U12776 (N_12776,N_9604,N_9581);
nand U12777 (N_12777,N_7883,N_5800);
or U12778 (N_12778,N_5218,N_8494);
and U12779 (N_12779,N_9581,N_8015);
nor U12780 (N_12780,N_7261,N_5119);
xor U12781 (N_12781,N_6839,N_9098);
nand U12782 (N_12782,N_9958,N_8778);
nor U12783 (N_12783,N_6352,N_8326);
nand U12784 (N_12784,N_7816,N_5978);
nand U12785 (N_12785,N_5602,N_7977);
nand U12786 (N_12786,N_5476,N_5158);
xnor U12787 (N_12787,N_9886,N_8433);
nor U12788 (N_12788,N_5151,N_5504);
or U12789 (N_12789,N_5008,N_9876);
nand U12790 (N_12790,N_8290,N_6855);
xor U12791 (N_12791,N_9578,N_9518);
xor U12792 (N_12792,N_9260,N_9263);
nand U12793 (N_12793,N_7473,N_9980);
or U12794 (N_12794,N_9662,N_5533);
and U12795 (N_12795,N_7219,N_5267);
or U12796 (N_12796,N_8551,N_5553);
xnor U12797 (N_12797,N_6580,N_8178);
and U12798 (N_12798,N_5097,N_6247);
and U12799 (N_12799,N_7375,N_8029);
nor U12800 (N_12800,N_5357,N_5423);
xor U12801 (N_12801,N_6895,N_7510);
or U12802 (N_12802,N_8481,N_8330);
or U12803 (N_12803,N_7565,N_7384);
nor U12804 (N_12804,N_9809,N_8220);
nand U12805 (N_12805,N_6857,N_9225);
and U12806 (N_12806,N_7536,N_8412);
and U12807 (N_12807,N_6387,N_6373);
or U12808 (N_12808,N_7080,N_9846);
xor U12809 (N_12809,N_6640,N_8512);
nand U12810 (N_12810,N_7711,N_6243);
xor U12811 (N_12811,N_7603,N_9946);
xnor U12812 (N_12812,N_6801,N_6538);
xnor U12813 (N_12813,N_6287,N_6984);
and U12814 (N_12814,N_9515,N_9083);
and U12815 (N_12815,N_6347,N_7274);
or U12816 (N_12816,N_7703,N_8818);
and U12817 (N_12817,N_7757,N_9083);
nand U12818 (N_12818,N_5183,N_7997);
or U12819 (N_12819,N_5344,N_8357);
and U12820 (N_12820,N_5463,N_5831);
nor U12821 (N_12821,N_7694,N_8548);
xnor U12822 (N_12822,N_9015,N_7809);
nor U12823 (N_12823,N_5590,N_9668);
nor U12824 (N_12824,N_9572,N_7127);
nand U12825 (N_12825,N_9639,N_8833);
or U12826 (N_12826,N_5811,N_8769);
or U12827 (N_12827,N_5902,N_5129);
or U12828 (N_12828,N_7012,N_8594);
nor U12829 (N_12829,N_6432,N_5159);
xnor U12830 (N_12830,N_6897,N_6080);
and U12831 (N_12831,N_5144,N_9132);
xnor U12832 (N_12832,N_5371,N_7675);
nor U12833 (N_12833,N_6591,N_9292);
or U12834 (N_12834,N_7929,N_5933);
nand U12835 (N_12835,N_6642,N_9016);
and U12836 (N_12836,N_5054,N_6962);
xnor U12837 (N_12837,N_9328,N_8347);
and U12838 (N_12838,N_6571,N_9591);
xnor U12839 (N_12839,N_9536,N_6836);
nand U12840 (N_12840,N_6250,N_7635);
nand U12841 (N_12841,N_5823,N_9676);
and U12842 (N_12842,N_9251,N_6713);
or U12843 (N_12843,N_9392,N_8211);
nand U12844 (N_12844,N_8421,N_5391);
nand U12845 (N_12845,N_8439,N_5680);
xor U12846 (N_12846,N_8906,N_8316);
nand U12847 (N_12847,N_6506,N_5161);
or U12848 (N_12848,N_5931,N_6480);
nor U12849 (N_12849,N_7514,N_9765);
and U12850 (N_12850,N_5628,N_8969);
xor U12851 (N_12851,N_5352,N_9844);
nand U12852 (N_12852,N_9334,N_5628);
xnor U12853 (N_12853,N_6949,N_5797);
nand U12854 (N_12854,N_7110,N_9049);
and U12855 (N_12855,N_7293,N_6942);
xnor U12856 (N_12856,N_6135,N_8293);
or U12857 (N_12857,N_5932,N_9793);
nor U12858 (N_12858,N_5571,N_6079);
nand U12859 (N_12859,N_9490,N_9401);
and U12860 (N_12860,N_7328,N_5707);
nand U12861 (N_12861,N_5804,N_6981);
or U12862 (N_12862,N_6886,N_5353);
xor U12863 (N_12863,N_7634,N_9027);
and U12864 (N_12864,N_5093,N_5514);
or U12865 (N_12865,N_5341,N_9829);
nand U12866 (N_12866,N_8834,N_8965);
nor U12867 (N_12867,N_7730,N_7907);
xor U12868 (N_12868,N_6967,N_5293);
nand U12869 (N_12869,N_6476,N_5240);
and U12870 (N_12870,N_6179,N_9740);
nand U12871 (N_12871,N_7051,N_8630);
or U12872 (N_12872,N_5970,N_5033);
xor U12873 (N_12873,N_6571,N_8915);
and U12874 (N_12874,N_5033,N_9129);
xnor U12875 (N_12875,N_6314,N_9404);
or U12876 (N_12876,N_9773,N_9389);
and U12877 (N_12877,N_7024,N_8924);
xnor U12878 (N_12878,N_8036,N_8980);
nand U12879 (N_12879,N_7150,N_9720);
nand U12880 (N_12880,N_6681,N_5071);
nor U12881 (N_12881,N_9939,N_9028);
xnor U12882 (N_12882,N_6859,N_8659);
or U12883 (N_12883,N_9892,N_9583);
nand U12884 (N_12884,N_7480,N_8529);
nor U12885 (N_12885,N_8041,N_9029);
nor U12886 (N_12886,N_8607,N_5529);
and U12887 (N_12887,N_6357,N_8208);
and U12888 (N_12888,N_7159,N_7427);
and U12889 (N_12889,N_7989,N_5728);
nand U12890 (N_12890,N_6600,N_8823);
nor U12891 (N_12891,N_8606,N_7927);
xnor U12892 (N_12892,N_9643,N_5267);
nor U12893 (N_12893,N_7665,N_6461);
nand U12894 (N_12894,N_8191,N_8021);
or U12895 (N_12895,N_8574,N_5366);
or U12896 (N_12896,N_7620,N_9204);
and U12897 (N_12897,N_9776,N_8844);
or U12898 (N_12898,N_5622,N_6469);
xnor U12899 (N_12899,N_7040,N_5050);
nand U12900 (N_12900,N_7778,N_7457);
nor U12901 (N_12901,N_9676,N_9803);
or U12902 (N_12902,N_8225,N_9762);
or U12903 (N_12903,N_9875,N_5440);
nand U12904 (N_12904,N_8362,N_7427);
or U12905 (N_12905,N_6345,N_5037);
nor U12906 (N_12906,N_7144,N_7804);
xor U12907 (N_12907,N_8195,N_8368);
xor U12908 (N_12908,N_7631,N_8698);
xor U12909 (N_12909,N_6082,N_7922);
nor U12910 (N_12910,N_5452,N_7514);
xnor U12911 (N_12911,N_8958,N_9808);
xor U12912 (N_12912,N_7461,N_9316);
nor U12913 (N_12913,N_9707,N_6388);
or U12914 (N_12914,N_5930,N_5024);
nor U12915 (N_12915,N_9817,N_9519);
and U12916 (N_12916,N_9378,N_6366);
and U12917 (N_12917,N_5268,N_7954);
nand U12918 (N_12918,N_8043,N_9412);
or U12919 (N_12919,N_6126,N_6740);
or U12920 (N_12920,N_9881,N_5797);
or U12921 (N_12921,N_8322,N_9808);
and U12922 (N_12922,N_8886,N_9481);
xnor U12923 (N_12923,N_7349,N_5255);
and U12924 (N_12924,N_5000,N_8737);
or U12925 (N_12925,N_7203,N_6078);
xnor U12926 (N_12926,N_9553,N_5529);
or U12927 (N_12927,N_8739,N_7844);
and U12928 (N_12928,N_7396,N_7740);
nor U12929 (N_12929,N_7217,N_7388);
or U12930 (N_12930,N_6135,N_9940);
nor U12931 (N_12931,N_8822,N_7458);
or U12932 (N_12932,N_6864,N_9788);
or U12933 (N_12933,N_6862,N_7199);
nor U12934 (N_12934,N_5175,N_6087);
xnor U12935 (N_12935,N_6985,N_9273);
and U12936 (N_12936,N_6971,N_7472);
nand U12937 (N_12937,N_6717,N_9815);
xor U12938 (N_12938,N_8262,N_5607);
xor U12939 (N_12939,N_5469,N_7418);
nand U12940 (N_12940,N_7779,N_5600);
nand U12941 (N_12941,N_5137,N_9273);
xnor U12942 (N_12942,N_6865,N_8445);
and U12943 (N_12943,N_9368,N_9868);
or U12944 (N_12944,N_5767,N_6517);
and U12945 (N_12945,N_5982,N_9064);
and U12946 (N_12946,N_7512,N_7772);
nand U12947 (N_12947,N_7655,N_6331);
nand U12948 (N_12948,N_6853,N_7104);
nor U12949 (N_12949,N_6760,N_7971);
and U12950 (N_12950,N_5968,N_9878);
nand U12951 (N_12951,N_8457,N_9974);
nor U12952 (N_12952,N_5181,N_6716);
nand U12953 (N_12953,N_9913,N_5697);
and U12954 (N_12954,N_5783,N_7327);
nor U12955 (N_12955,N_8073,N_9851);
xor U12956 (N_12956,N_9080,N_6280);
nor U12957 (N_12957,N_6297,N_6532);
or U12958 (N_12958,N_6171,N_5391);
nand U12959 (N_12959,N_6634,N_8281);
and U12960 (N_12960,N_8136,N_8483);
xor U12961 (N_12961,N_5105,N_9715);
xnor U12962 (N_12962,N_8876,N_9494);
nand U12963 (N_12963,N_8787,N_9003);
or U12964 (N_12964,N_9056,N_8505);
and U12965 (N_12965,N_7923,N_9163);
nor U12966 (N_12966,N_9692,N_5221);
nand U12967 (N_12967,N_6338,N_8073);
or U12968 (N_12968,N_7621,N_7729);
xnor U12969 (N_12969,N_5879,N_9005);
or U12970 (N_12970,N_9654,N_8067);
or U12971 (N_12971,N_6324,N_7911);
nor U12972 (N_12972,N_8101,N_5492);
xor U12973 (N_12973,N_8718,N_8599);
or U12974 (N_12974,N_7137,N_8733);
xor U12975 (N_12975,N_9703,N_7117);
nor U12976 (N_12976,N_7672,N_7353);
and U12977 (N_12977,N_5651,N_8993);
nand U12978 (N_12978,N_6858,N_7503);
xnor U12979 (N_12979,N_8882,N_6761);
and U12980 (N_12980,N_8142,N_8150);
xnor U12981 (N_12981,N_5961,N_5935);
nor U12982 (N_12982,N_8622,N_7090);
nor U12983 (N_12983,N_6394,N_7630);
xor U12984 (N_12984,N_9893,N_7705);
nor U12985 (N_12985,N_7600,N_8440);
and U12986 (N_12986,N_8782,N_5963);
or U12987 (N_12987,N_5417,N_9526);
xnor U12988 (N_12988,N_8150,N_8983);
and U12989 (N_12989,N_6029,N_5567);
or U12990 (N_12990,N_5007,N_9396);
nor U12991 (N_12991,N_5241,N_7542);
nand U12992 (N_12992,N_8369,N_9764);
nand U12993 (N_12993,N_7076,N_9283);
nor U12994 (N_12994,N_5534,N_7091);
and U12995 (N_12995,N_6788,N_9074);
and U12996 (N_12996,N_9505,N_8388);
nand U12997 (N_12997,N_8751,N_7210);
nor U12998 (N_12998,N_6724,N_7277);
nand U12999 (N_12999,N_5249,N_5581);
or U13000 (N_13000,N_7927,N_7546);
nor U13001 (N_13001,N_6739,N_6451);
nor U13002 (N_13002,N_8566,N_5161);
nor U13003 (N_13003,N_7025,N_8309);
xor U13004 (N_13004,N_6760,N_5002);
nor U13005 (N_13005,N_7899,N_7070);
nor U13006 (N_13006,N_5713,N_5640);
or U13007 (N_13007,N_7720,N_6948);
nand U13008 (N_13008,N_6628,N_6411);
nor U13009 (N_13009,N_9462,N_5736);
xnor U13010 (N_13010,N_6439,N_6299);
nor U13011 (N_13011,N_5661,N_9979);
or U13012 (N_13012,N_9036,N_8916);
nand U13013 (N_13013,N_5198,N_7018);
or U13014 (N_13014,N_6403,N_6765);
and U13015 (N_13015,N_5175,N_5872);
and U13016 (N_13016,N_5291,N_5427);
xnor U13017 (N_13017,N_5104,N_9452);
nor U13018 (N_13018,N_8807,N_9627);
nor U13019 (N_13019,N_8346,N_9723);
and U13020 (N_13020,N_8974,N_6611);
nor U13021 (N_13021,N_9986,N_7209);
nand U13022 (N_13022,N_8285,N_7075);
or U13023 (N_13023,N_6516,N_7272);
nor U13024 (N_13024,N_6266,N_9812);
xor U13025 (N_13025,N_7376,N_6459);
and U13026 (N_13026,N_8570,N_8277);
xnor U13027 (N_13027,N_9415,N_8477);
or U13028 (N_13028,N_7855,N_7949);
nand U13029 (N_13029,N_9979,N_9795);
xor U13030 (N_13030,N_7375,N_8740);
nor U13031 (N_13031,N_8145,N_7549);
and U13032 (N_13032,N_5346,N_6819);
or U13033 (N_13033,N_9444,N_9249);
nor U13034 (N_13034,N_9639,N_6378);
nand U13035 (N_13035,N_9303,N_9952);
nor U13036 (N_13036,N_8036,N_6291);
nand U13037 (N_13037,N_8925,N_9431);
and U13038 (N_13038,N_5324,N_5308);
nor U13039 (N_13039,N_5477,N_7213);
nand U13040 (N_13040,N_6202,N_7771);
or U13041 (N_13041,N_9228,N_6459);
and U13042 (N_13042,N_9195,N_9506);
nand U13043 (N_13043,N_6262,N_6800);
nand U13044 (N_13044,N_9683,N_7695);
nor U13045 (N_13045,N_6931,N_6109);
or U13046 (N_13046,N_5565,N_7642);
and U13047 (N_13047,N_9566,N_5894);
nand U13048 (N_13048,N_7251,N_5433);
xnor U13049 (N_13049,N_9842,N_5171);
and U13050 (N_13050,N_9376,N_6782);
xor U13051 (N_13051,N_5782,N_9142);
nor U13052 (N_13052,N_9018,N_6666);
or U13053 (N_13053,N_8922,N_6522);
nand U13054 (N_13054,N_9821,N_8212);
nor U13055 (N_13055,N_7949,N_6123);
and U13056 (N_13056,N_6531,N_9011);
or U13057 (N_13057,N_6927,N_7298);
or U13058 (N_13058,N_7986,N_6814);
nor U13059 (N_13059,N_8471,N_5415);
nand U13060 (N_13060,N_8276,N_8986);
xor U13061 (N_13061,N_7689,N_9108);
and U13062 (N_13062,N_5192,N_9189);
nand U13063 (N_13063,N_6863,N_7251);
or U13064 (N_13064,N_5006,N_7095);
and U13065 (N_13065,N_8177,N_5680);
nand U13066 (N_13066,N_8671,N_6826);
and U13067 (N_13067,N_5096,N_8526);
nand U13068 (N_13068,N_5436,N_6927);
or U13069 (N_13069,N_6165,N_8113);
and U13070 (N_13070,N_6982,N_7911);
and U13071 (N_13071,N_6589,N_7111);
xnor U13072 (N_13072,N_5406,N_9026);
nor U13073 (N_13073,N_8690,N_6722);
xor U13074 (N_13074,N_9907,N_6526);
and U13075 (N_13075,N_8058,N_7160);
nand U13076 (N_13076,N_9141,N_7560);
or U13077 (N_13077,N_8219,N_5266);
nand U13078 (N_13078,N_9203,N_9675);
nand U13079 (N_13079,N_9480,N_8657);
xor U13080 (N_13080,N_8805,N_7352);
or U13081 (N_13081,N_6075,N_7698);
and U13082 (N_13082,N_9263,N_8627);
or U13083 (N_13083,N_7017,N_9134);
or U13084 (N_13084,N_9995,N_7158);
nor U13085 (N_13085,N_6499,N_8442);
xor U13086 (N_13086,N_9362,N_8234);
and U13087 (N_13087,N_8741,N_5325);
or U13088 (N_13088,N_6084,N_5367);
or U13089 (N_13089,N_9850,N_5715);
or U13090 (N_13090,N_7445,N_8561);
and U13091 (N_13091,N_7066,N_7224);
or U13092 (N_13092,N_6360,N_6732);
or U13093 (N_13093,N_6005,N_9528);
nor U13094 (N_13094,N_9462,N_8690);
nand U13095 (N_13095,N_7796,N_8109);
nor U13096 (N_13096,N_9383,N_5809);
nand U13097 (N_13097,N_7814,N_6334);
nand U13098 (N_13098,N_7617,N_5671);
nor U13099 (N_13099,N_5879,N_5154);
nand U13100 (N_13100,N_6738,N_9209);
and U13101 (N_13101,N_7546,N_6332);
nand U13102 (N_13102,N_9236,N_6978);
or U13103 (N_13103,N_5674,N_5857);
nor U13104 (N_13104,N_6408,N_6503);
nor U13105 (N_13105,N_6352,N_9169);
xnor U13106 (N_13106,N_8784,N_9397);
and U13107 (N_13107,N_8467,N_9681);
nand U13108 (N_13108,N_7805,N_6552);
xnor U13109 (N_13109,N_6276,N_5879);
xor U13110 (N_13110,N_6317,N_7138);
xor U13111 (N_13111,N_9733,N_9363);
nand U13112 (N_13112,N_7503,N_9000);
nand U13113 (N_13113,N_5915,N_5923);
or U13114 (N_13114,N_5481,N_6436);
nor U13115 (N_13115,N_7605,N_5630);
and U13116 (N_13116,N_5447,N_5431);
xor U13117 (N_13117,N_7334,N_7685);
nand U13118 (N_13118,N_5050,N_7777);
xnor U13119 (N_13119,N_8695,N_5780);
or U13120 (N_13120,N_6162,N_7941);
and U13121 (N_13121,N_6513,N_8790);
xnor U13122 (N_13122,N_7978,N_8875);
or U13123 (N_13123,N_6990,N_9402);
or U13124 (N_13124,N_8403,N_5343);
and U13125 (N_13125,N_6772,N_5151);
nand U13126 (N_13126,N_6259,N_5433);
and U13127 (N_13127,N_8117,N_6070);
or U13128 (N_13128,N_9571,N_8609);
xnor U13129 (N_13129,N_5269,N_8980);
nor U13130 (N_13130,N_9354,N_5091);
or U13131 (N_13131,N_8194,N_6069);
and U13132 (N_13132,N_8378,N_6830);
and U13133 (N_13133,N_8043,N_9254);
xor U13134 (N_13134,N_7462,N_8270);
and U13135 (N_13135,N_7692,N_8263);
or U13136 (N_13136,N_8646,N_6217);
xnor U13137 (N_13137,N_5224,N_7210);
nand U13138 (N_13138,N_8305,N_8550);
nor U13139 (N_13139,N_9894,N_6919);
xnor U13140 (N_13140,N_6768,N_6338);
or U13141 (N_13141,N_9416,N_9253);
or U13142 (N_13142,N_6972,N_6997);
and U13143 (N_13143,N_8388,N_8878);
nor U13144 (N_13144,N_9055,N_6636);
or U13145 (N_13145,N_8525,N_7410);
nand U13146 (N_13146,N_9106,N_9042);
or U13147 (N_13147,N_7697,N_9224);
and U13148 (N_13148,N_5749,N_8208);
nor U13149 (N_13149,N_7547,N_6730);
and U13150 (N_13150,N_9175,N_9169);
or U13151 (N_13151,N_9845,N_9477);
or U13152 (N_13152,N_5702,N_8713);
nor U13153 (N_13153,N_6826,N_8584);
or U13154 (N_13154,N_5328,N_7443);
xnor U13155 (N_13155,N_6021,N_7130);
and U13156 (N_13156,N_9777,N_5077);
and U13157 (N_13157,N_9415,N_9058);
nor U13158 (N_13158,N_7386,N_8581);
nor U13159 (N_13159,N_8605,N_6492);
nor U13160 (N_13160,N_8525,N_7451);
and U13161 (N_13161,N_9364,N_5690);
nor U13162 (N_13162,N_6240,N_9092);
nand U13163 (N_13163,N_6333,N_8067);
nor U13164 (N_13164,N_9123,N_5189);
xnor U13165 (N_13165,N_9217,N_9423);
nand U13166 (N_13166,N_9569,N_8115);
and U13167 (N_13167,N_5777,N_7336);
nand U13168 (N_13168,N_6061,N_9630);
xnor U13169 (N_13169,N_5256,N_5626);
and U13170 (N_13170,N_8652,N_5340);
xor U13171 (N_13171,N_6004,N_8152);
and U13172 (N_13172,N_7202,N_6707);
and U13173 (N_13173,N_5373,N_5771);
or U13174 (N_13174,N_8959,N_7244);
xor U13175 (N_13175,N_5673,N_6982);
xnor U13176 (N_13176,N_5779,N_8061);
and U13177 (N_13177,N_5171,N_8973);
xor U13178 (N_13178,N_5564,N_8844);
nor U13179 (N_13179,N_5766,N_5602);
and U13180 (N_13180,N_7927,N_8504);
xnor U13181 (N_13181,N_7224,N_8302);
and U13182 (N_13182,N_5880,N_6680);
and U13183 (N_13183,N_9807,N_8657);
nand U13184 (N_13184,N_6454,N_6100);
nand U13185 (N_13185,N_8850,N_9749);
nand U13186 (N_13186,N_5161,N_7992);
xor U13187 (N_13187,N_7316,N_5945);
or U13188 (N_13188,N_7510,N_9173);
nor U13189 (N_13189,N_7462,N_7125);
and U13190 (N_13190,N_5348,N_8210);
nand U13191 (N_13191,N_6589,N_7848);
nor U13192 (N_13192,N_8045,N_6038);
or U13193 (N_13193,N_5963,N_5595);
nand U13194 (N_13194,N_7798,N_9560);
nor U13195 (N_13195,N_5853,N_9507);
nor U13196 (N_13196,N_9835,N_8295);
nand U13197 (N_13197,N_8681,N_6379);
xor U13198 (N_13198,N_7460,N_9107);
or U13199 (N_13199,N_6778,N_7793);
nor U13200 (N_13200,N_7241,N_7048);
nor U13201 (N_13201,N_5780,N_9303);
or U13202 (N_13202,N_5690,N_6927);
nand U13203 (N_13203,N_5505,N_9149);
or U13204 (N_13204,N_8945,N_9882);
xnor U13205 (N_13205,N_7849,N_9747);
or U13206 (N_13206,N_8795,N_5413);
xor U13207 (N_13207,N_8745,N_9749);
nand U13208 (N_13208,N_9511,N_8049);
nor U13209 (N_13209,N_9724,N_9024);
and U13210 (N_13210,N_9654,N_8499);
nand U13211 (N_13211,N_8458,N_7104);
xnor U13212 (N_13212,N_6892,N_7012);
and U13213 (N_13213,N_5082,N_7389);
nor U13214 (N_13214,N_6785,N_5450);
and U13215 (N_13215,N_5526,N_5302);
nor U13216 (N_13216,N_7196,N_7208);
nor U13217 (N_13217,N_8406,N_7970);
and U13218 (N_13218,N_8700,N_5393);
nand U13219 (N_13219,N_9290,N_7956);
and U13220 (N_13220,N_6478,N_9673);
nor U13221 (N_13221,N_7817,N_7044);
xor U13222 (N_13222,N_9381,N_9458);
nor U13223 (N_13223,N_6230,N_8879);
nand U13224 (N_13224,N_7364,N_9499);
and U13225 (N_13225,N_6308,N_8400);
or U13226 (N_13226,N_6186,N_8040);
or U13227 (N_13227,N_8274,N_7534);
and U13228 (N_13228,N_6876,N_8974);
nand U13229 (N_13229,N_7588,N_6670);
or U13230 (N_13230,N_8966,N_6526);
nand U13231 (N_13231,N_5124,N_7591);
and U13232 (N_13232,N_6366,N_9846);
nor U13233 (N_13233,N_8995,N_6918);
xor U13234 (N_13234,N_8114,N_7442);
xor U13235 (N_13235,N_9395,N_5696);
or U13236 (N_13236,N_7859,N_6541);
xor U13237 (N_13237,N_7690,N_8934);
nand U13238 (N_13238,N_5539,N_5827);
xor U13239 (N_13239,N_6890,N_6097);
nand U13240 (N_13240,N_9317,N_6826);
nand U13241 (N_13241,N_8658,N_7469);
or U13242 (N_13242,N_9219,N_8094);
and U13243 (N_13243,N_7367,N_6742);
and U13244 (N_13244,N_7954,N_9337);
or U13245 (N_13245,N_6735,N_5937);
nand U13246 (N_13246,N_7616,N_5076);
or U13247 (N_13247,N_9760,N_6370);
nand U13248 (N_13248,N_7074,N_6006);
xor U13249 (N_13249,N_6193,N_9307);
or U13250 (N_13250,N_9087,N_9806);
and U13251 (N_13251,N_7117,N_9869);
and U13252 (N_13252,N_6717,N_9955);
nor U13253 (N_13253,N_5158,N_6681);
nor U13254 (N_13254,N_9949,N_5974);
nand U13255 (N_13255,N_8279,N_6181);
or U13256 (N_13256,N_7367,N_9442);
and U13257 (N_13257,N_6406,N_8073);
nand U13258 (N_13258,N_6958,N_8634);
nand U13259 (N_13259,N_5450,N_9097);
nor U13260 (N_13260,N_9567,N_9994);
and U13261 (N_13261,N_9026,N_9961);
nand U13262 (N_13262,N_5412,N_6060);
and U13263 (N_13263,N_9462,N_7410);
or U13264 (N_13264,N_8108,N_7368);
nand U13265 (N_13265,N_8944,N_8550);
nand U13266 (N_13266,N_6262,N_5616);
and U13267 (N_13267,N_8184,N_9068);
and U13268 (N_13268,N_9800,N_5629);
xnor U13269 (N_13269,N_8969,N_5927);
and U13270 (N_13270,N_6753,N_9776);
and U13271 (N_13271,N_7437,N_5658);
nand U13272 (N_13272,N_5914,N_7317);
xor U13273 (N_13273,N_8826,N_9512);
xor U13274 (N_13274,N_6127,N_8277);
or U13275 (N_13275,N_9035,N_5681);
or U13276 (N_13276,N_5898,N_6064);
xnor U13277 (N_13277,N_8280,N_9552);
or U13278 (N_13278,N_7608,N_7726);
nor U13279 (N_13279,N_5980,N_7780);
or U13280 (N_13280,N_6724,N_5236);
or U13281 (N_13281,N_7406,N_8297);
nor U13282 (N_13282,N_6199,N_5888);
xor U13283 (N_13283,N_9652,N_7829);
nand U13284 (N_13284,N_5656,N_8433);
nand U13285 (N_13285,N_8057,N_8495);
xor U13286 (N_13286,N_6433,N_5379);
or U13287 (N_13287,N_5077,N_6501);
or U13288 (N_13288,N_5278,N_9904);
xor U13289 (N_13289,N_7454,N_6950);
nand U13290 (N_13290,N_7054,N_7806);
and U13291 (N_13291,N_8272,N_9853);
and U13292 (N_13292,N_5315,N_6222);
and U13293 (N_13293,N_7240,N_9550);
and U13294 (N_13294,N_7937,N_7164);
xnor U13295 (N_13295,N_8298,N_6152);
xnor U13296 (N_13296,N_5347,N_5504);
and U13297 (N_13297,N_6676,N_7280);
and U13298 (N_13298,N_8109,N_8782);
and U13299 (N_13299,N_7869,N_6594);
and U13300 (N_13300,N_8904,N_7713);
or U13301 (N_13301,N_9119,N_6709);
nor U13302 (N_13302,N_5129,N_9309);
nor U13303 (N_13303,N_6121,N_7586);
xor U13304 (N_13304,N_8439,N_6884);
nor U13305 (N_13305,N_5648,N_7774);
and U13306 (N_13306,N_6995,N_6388);
nor U13307 (N_13307,N_7688,N_6963);
and U13308 (N_13308,N_7923,N_5034);
xnor U13309 (N_13309,N_9039,N_7598);
nor U13310 (N_13310,N_7526,N_6812);
nand U13311 (N_13311,N_5265,N_5093);
nand U13312 (N_13312,N_7887,N_6590);
or U13313 (N_13313,N_9351,N_6405);
nor U13314 (N_13314,N_6506,N_6697);
nand U13315 (N_13315,N_9464,N_5862);
and U13316 (N_13316,N_9784,N_9057);
nand U13317 (N_13317,N_9926,N_7667);
nor U13318 (N_13318,N_5554,N_6036);
nor U13319 (N_13319,N_9138,N_7755);
and U13320 (N_13320,N_7093,N_9643);
or U13321 (N_13321,N_6388,N_5452);
xnor U13322 (N_13322,N_9112,N_5642);
nor U13323 (N_13323,N_6682,N_5030);
nor U13324 (N_13324,N_8624,N_6219);
and U13325 (N_13325,N_8671,N_8968);
xnor U13326 (N_13326,N_6050,N_6258);
or U13327 (N_13327,N_5788,N_6477);
or U13328 (N_13328,N_9065,N_7589);
nand U13329 (N_13329,N_8527,N_8611);
nand U13330 (N_13330,N_6042,N_8004);
xor U13331 (N_13331,N_9688,N_5342);
and U13332 (N_13332,N_6456,N_7638);
xnor U13333 (N_13333,N_6231,N_8269);
nor U13334 (N_13334,N_5617,N_9198);
and U13335 (N_13335,N_5756,N_5113);
nor U13336 (N_13336,N_5817,N_6820);
nor U13337 (N_13337,N_9287,N_7900);
xor U13338 (N_13338,N_5460,N_8198);
nor U13339 (N_13339,N_5235,N_5731);
nor U13340 (N_13340,N_8411,N_6682);
nor U13341 (N_13341,N_9213,N_8451);
and U13342 (N_13342,N_9008,N_9972);
xnor U13343 (N_13343,N_8249,N_6727);
nand U13344 (N_13344,N_5841,N_5595);
nand U13345 (N_13345,N_7708,N_5589);
and U13346 (N_13346,N_9935,N_9783);
nand U13347 (N_13347,N_5751,N_9286);
nand U13348 (N_13348,N_9046,N_6098);
nand U13349 (N_13349,N_6686,N_6325);
nor U13350 (N_13350,N_6232,N_5888);
xnor U13351 (N_13351,N_7424,N_5483);
nor U13352 (N_13352,N_6109,N_9292);
xor U13353 (N_13353,N_7408,N_5208);
or U13354 (N_13354,N_8036,N_5405);
nand U13355 (N_13355,N_6429,N_9851);
xnor U13356 (N_13356,N_5114,N_6205);
xor U13357 (N_13357,N_5194,N_7210);
xnor U13358 (N_13358,N_9411,N_7512);
xor U13359 (N_13359,N_6184,N_6305);
or U13360 (N_13360,N_8624,N_7958);
and U13361 (N_13361,N_7309,N_9932);
xor U13362 (N_13362,N_6639,N_9601);
and U13363 (N_13363,N_5946,N_8670);
nand U13364 (N_13364,N_6682,N_7673);
and U13365 (N_13365,N_8890,N_9102);
nor U13366 (N_13366,N_9202,N_8249);
nor U13367 (N_13367,N_9884,N_8280);
xor U13368 (N_13368,N_5456,N_9690);
and U13369 (N_13369,N_7634,N_9422);
and U13370 (N_13370,N_5515,N_9501);
and U13371 (N_13371,N_8169,N_8628);
nor U13372 (N_13372,N_8695,N_6216);
and U13373 (N_13373,N_7667,N_6114);
or U13374 (N_13374,N_5960,N_9577);
xor U13375 (N_13375,N_7862,N_8427);
xor U13376 (N_13376,N_6698,N_8702);
nand U13377 (N_13377,N_8286,N_5391);
nor U13378 (N_13378,N_7120,N_9185);
and U13379 (N_13379,N_5297,N_7307);
and U13380 (N_13380,N_8748,N_8999);
xnor U13381 (N_13381,N_5264,N_6603);
nor U13382 (N_13382,N_9810,N_7679);
nand U13383 (N_13383,N_9083,N_8495);
or U13384 (N_13384,N_6851,N_9150);
or U13385 (N_13385,N_6922,N_9443);
nand U13386 (N_13386,N_9361,N_5955);
nor U13387 (N_13387,N_7475,N_8415);
nor U13388 (N_13388,N_8303,N_5935);
xor U13389 (N_13389,N_7519,N_7371);
nor U13390 (N_13390,N_5850,N_6452);
xor U13391 (N_13391,N_6003,N_8043);
nor U13392 (N_13392,N_7542,N_9861);
or U13393 (N_13393,N_5181,N_9870);
and U13394 (N_13394,N_6655,N_6631);
or U13395 (N_13395,N_6435,N_6330);
or U13396 (N_13396,N_9823,N_8959);
and U13397 (N_13397,N_5092,N_9749);
xnor U13398 (N_13398,N_7538,N_6989);
nand U13399 (N_13399,N_7024,N_5802);
or U13400 (N_13400,N_7235,N_5539);
nor U13401 (N_13401,N_7247,N_7086);
nor U13402 (N_13402,N_8143,N_6523);
or U13403 (N_13403,N_8756,N_6984);
nor U13404 (N_13404,N_6814,N_5446);
xnor U13405 (N_13405,N_7896,N_8238);
nand U13406 (N_13406,N_9981,N_6344);
xnor U13407 (N_13407,N_7311,N_9795);
and U13408 (N_13408,N_6209,N_5749);
or U13409 (N_13409,N_7640,N_5911);
nand U13410 (N_13410,N_7878,N_7998);
or U13411 (N_13411,N_9881,N_7402);
nor U13412 (N_13412,N_5607,N_6958);
nand U13413 (N_13413,N_7936,N_8532);
xnor U13414 (N_13414,N_8449,N_8375);
nand U13415 (N_13415,N_9914,N_9349);
nor U13416 (N_13416,N_5174,N_9222);
xnor U13417 (N_13417,N_5315,N_7635);
xor U13418 (N_13418,N_6757,N_9100);
xor U13419 (N_13419,N_9302,N_5707);
and U13420 (N_13420,N_7272,N_7609);
or U13421 (N_13421,N_5684,N_7544);
nor U13422 (N_13422,N_7087,N_5655);
xor U13423 (N_13423,N_7895,N_6700);
nand U13424 (N_13424,N_7575,N_8836);
nand U13425 (N_13425,N_6782,N_7048);
or U13426 (N_13426,N_6146,N_8202);
nand U13427 (N_13427,N_6567,N_7299);
nor U13428 (N_13428,N_6331,N_6710);
xor U13429 (N_13429,N_8767,N_7211);
nand U13430 (N_13430,N_7371,N_7293);
xnor U13431 (N_13431,N_6540,N_7544);
nor U13432 (N_13432,N_8314,N_8271);
or U13433 (N_13433,N_9764,N_5442);
or U13434 (N_13434,N_6072,N_7806);
and U13435 (N_13435,N_9156,N_9496);
and U13436 (N_13436,N_5888,N_9557);
and U13437 (N_13437,N_7400,N_8039);
nor U13438 (N_13438,N_7697,N_5471);
or U13439 (N_13439,N_8424,N_6925);
and U13440 (N_13440,N_7892,N_9264);
and U13441 (N_13441,N_9422,N_7625);
or U13442 (N_13442,N_7083,N_7809);
xor U13443 (N_13443,N_7253,N_8415);
nor U13444 (N_13444,N_5327,N_7117);
and U13445 (N_13445,N_5023,N_7599);
nor U13446 (N_13446,N_9186,N_5673);
xor U13447 (N_13447,N_7529,N_8710);
and U13448 (N_13448,N_7042,N_6776);
xnor U13449 (N_13449,N_6542,N_6494);
nand U13450 (N_13450,N_9905,N_5355);
xor U13451 (N_13451,N_6067,N_9313);
or U13452 (N_13452,N_5671,N_6981);
and U13453 (N_13453,N_5230,N_6365);
and U13454 (N_13454,N_7553,N_9944);
or U13455 (N_13455,N_8936,N_5358);
xnor U13456 (N_13456,N_7380,N_9701);
xor U13457 (N_13457,N_6348,N_8757);
nand U13458 (N_13458,N_7603,N_8257);
xor U13459 (N_13459,N_6395,N_6769);
and U13460 (N_13460,N_6084,N_6681);
or U13461 (N_13461,N_5452,N_5703);
xor U13462 (N_13462,N_6254,N_6577);
nor U13463 (N_13463,N_7934,N_7695);
xnor U13464 (N_13464,N_8848,N_8394);
or U13465 (N_13465,N_6672,N_9026);
xnor U13466 (N_13466,N_9601,N_7978);
or U13467 (N_13467,N_6328,N_9826);
and U13468 (N_13468,N_8712,N_5259);
nor U13469 (N_13469,N_9476,N_6617);
nor U13470 (N_13470,N_6649,N_5421);
xor U13471 (N_13471,N_8961,N_8810);
xor U13472 (N_13472,N_6317,N_9906);
nor U13473 (N_13473,N_8926,N_6144);
xnor U13474 (N_13474,N_8893,N_6328);
nand U13475 (N_13475,N_9706,N_6893);
nor U13476 (N_13476,N_6908,N_9829);
xor U13477 (N_13477,N_8564,N_6048);
and U13478 (N_13478,N_9465,N_8707);
and U13479 (N_13479,N_5854,N_9232);
nor U13480 (N_13480,N_9148,N_6872);
nand U13481 (N_13481,N_5377,N_6987);
xnor U13482 (N_13482,N_8249,N_7044);
nand U13483 (N_13483,N_6822,N_8059);
and U13484 (N_13484,N_6557,N_8668);
and U13485 (N_13485,N_8302,N_6436);
xnor U13486 (N_13486,N_6195,N_6044);
or U13487 (N_13487,N_9639,N_8838);
nand U13488 (N_13488,N_8914,N_8858);
or U13489 (N_13489,N_6389,N_7556);
nand U13490 (N_13490,N_5775,N_8413);
or U13491 (N_13491,N_8985,N_9957);
or U13492 (N_13492,N_7087,N_9411);
and U13493 (N_13493,N_8501,N_5454);
nand U13494 (N_13494,N_9158,N_6463);
nor U13495 (N_13495,N_8872,N_9772);
and U13496 (N_13496,N_5621,N_5821);
and U13497 (N_13497,N_5613,N_6124);
and U13498 (N_13498,N_9595,N_7584);
xnor U13499 (N_13499,N_7691,N_8183);
or U13500 (N_13500,N_8846,N_5648);
nor U13501 (N_13501,N_8325,N_9208);
xnor U13502 (N_13502,N_9888,N_5662);
nand U13503 (N_13503,N_6664,N_6380);
nand U13504 (N_13504,N_5562,N_6891);
xor U13505 (N_13505,N_6978,N_9508);
nor U13506 (N_13506,N_8944,N_9997);
or U13507 (N_13507,N_7118,N_7034);
nand U13508 (N_13508,N_8021,N_5908);
or U13509 (N_13509,N_5462,N_8635);
xor U13510 (N_13510,N_6515,N_6099);
nor U13511 (N_13511,N_7850,N_5934);
nand U13512 (N_13512,N_6408,N_9770);
xor U13513 (N_13513,N_5281,N_9449);
and U13514 (N_13514,N_8952,N_7976);
and U13515 (N_13515,N_8396,N_7995);
nor U13516 (N_13516,N_8426,N_8827);
or U13517 (N_13517,N_8354,N_9384);
xnor U13518 (N_13518,N_9051,N_7496);
xor U13519 (N_13519,N_6862,N_8988);
or U13520 (N_13520,N_5443,N_5802);
xnor U13521 (N_13521,N_6017,N_7024);
nand U13522 (N_13522,N_5651,N_5433);
or U13523 (N_13523,N_5504,N_8595);
or U13524 (N_13524,N_6045,N_7694);
and U13525 (N_13525,N_9834,N_7482);
or U13526 (N_13526,N_5885,N_7642);
nor U13527 (N_13527,N_7702,N_7802);
nand U13528 (N_13528,N_8993,N_6168);
nor U13529 (N_13529,N_7753,N_8961);
xor U13530 (N_13530,N_8049,N_6311);
nand U13531 (N_13531,N_9890,N_8049);
nand U13532 (N_13532,N_5804,N_9067);
nor U13533 (N_13533,N_7465,N_7985);
and U13534 (N_13534,N_8617,N_6837);
or U13535 (N_13535,N_8106,N_7834);
or U13536 (N_13536,N_9392,N_7207);
or U13537 (N_13537,N_9868,N_8307);
and U13538 (N_13538,N_5244,N_9512);
xnor U13539 (N_13539,N_8997,N_5517);
and U13540 (N_13540,N_7730,N_9260);
xor U13541 (N_13541,N_7457,N_8394);
nor U13542 (N_13542,N_6130,N_7923);
and U13543 (N_13543,N_5349,N_7582);
nand U13544 (N_13544,N_9775,N_6314);
nor U13545 (N_13545,N_9462,N_9886);
xnor U13546 (N_13546,N_5438,N_9759);
and U13547 (N_13547,N_5745,N_5351);
and U13548 (N_13548,N_9085,N_8497);
xnor U13549 (N_13549,N_8984,N_6672);
and U13550 (N_13550,N_6555,N_6920);
xor U13551 (N_13551,N_6001,N_8649);
xnor U13552 (N_13552,N_6214,N_7329);
and U13553 (N_13553,N_5137,N_5282);
nor U13554 (N_13554,N_5051,N_9973);
or U13555 (N_13555,N_8768,N_6579);
nand U13556 (N_13556,N_7569,N_7745);
nand U13557 (N_13557,N_8101,N_8369);
and U13558 (N_13558,N_8113,N_5608);
or U13559 (N_13559,N_5621,N_8602);
or U13560 (N_13560,N_8756,N_5507);
and U13561 (N_13561,N_9673,N_6085);
xnor U13562 (N_13562,N_5319,N_7448);
and U13563 (N_13563,N_6999,N_5737);
xnor U13564 (N_13564,N_5946,N_6916);
nand U13565 (N_13565,N_8785,N_7841);
nand U13566 (N_13566,N_6077,N_5632);
xor U13567 (N_13567,N_5291,N_7254);
xnor U13568 (N_13568,N_6086,N_6006);
nor U13569 (N_13569,N_6105,N_9769);
or U13570 (N_13570,N_9356,N_6586);
and U13571 (N_13571,N_7117,N_6727);
xnor U13572 (N_13572,N_8583,N_5818);
xnor U13573 (N_13573,N_6550,N_9348);
and U13574 (N_13574,N_5464,N_6948);
nand U13575 (N_13575,N_7518,N_7822);
nand U13576 (N_13576,N_9703,N_9484);
and U13577 (N_13577,N_6273,N_5344);
nand U13578 (N_13578,N_8203,N_7184);
nor U13579 (N_13579,N_5890,N_8562);
and U13580 (N_13580,N_5022,N_9101);
nand U13581 (N_13581,N_8722,N_6916);
and U13582 (N_13582,N_6747,N_8052);
or U13583 (N_13583,N_6068,N_9935);
nand U13584 (N_13584,N_9354,N_8406);
xor U13585 (N_13585,N_7575,N_9113);
nor U13586 (N_13586,N_5615,N_6220);
and U13587 (N_13587,N_7078,N_5919);
and U13588 (N_13588,N_7203,N_7442);
nand U13589 (N_13589,N_9789,N_6399);
or U13590 (N_13590,N_6139,N_6729);
or U13591 (N_13591,N_7823,N_7858);
xnor U13592 (N_13592,N_7175,N_6769);
nand U13593 (N_13593,N_7210,N_6010);
xor U13594 (N_13594,N_7449,N_9514);
and U13595 (N_13595,N_6703,N_5360);
xnor U13596 (N_13596,N_9826,N_6972);
nand U13597 (N_13597,N_9029,N_5868);
nand U13598 (N_13598,N_6756,N_5940);
or U13599 (N_13599,N_8542,N_5102);
nor U13600 (N_13600,N_5400,N_8496);
and U13601 (N_13601,N_6445,N_9168);
or U13602 (N_13602,N_9047,N_6401);
or U13603 (N_13603,N_8095,N_6533);
or U13604 (N_13604,N_5390,N_6693);
xor U13605 (N_13605,N_8028,N_9526);
nor U13606 (N_13606,N_8536,N_5180);
xor U13607 (N_13607,N_6035,N_8797);
xor U13608 (N_13608,N_5265,N_9933);
or U13609 (N_13609,N_8118,N_5238);
xor U13610 (N_13610,N_7816,N_7269);
or U13611 (N_13611,N_5846,N_9924);
nand U13612 (N_13612,N_5630,N_6486);
or U13613 (N_13613,N_5234,N_5362);
nor U13614 (N_13614,N_9368,N_5652);
and U13615 (N_13615,N_7177,N_5777);
nand U13616 (N_13616,N_8270,N_5010);
and U13617 (N_13617,N_6355,N_6740);
nand U13618 (N_13618,N_6457,N_8069);
nor U13619 (N_13619,N_8832,N_7411);
nor U13620 (N_13620,N_6496,N_9630);
xor U13621 (N_13621,N_5455,N_5669);
nand U13622 (N_13622,N_6268,N_7483);
or U13623 (N_13623,N_7545,N_8717);
nor U13624 (N_13624,N_5404,N_7324);
xor U13625 (N_13625,N_9529,N_5603);
nor U13626 (N_13626,N_7004,N_5377);
or U13627 (N_13627,N_7754,N_8209);
nor U13628 (N_13628,N_5782,N_5668);
nand U13629 (N_13629,N_7930,N_5132);
or U13630 (N_13630,N_7314,N_9052);
or U13631 (N_13631,N_9976,N_6461);
or U13632 (N_13632,N_6510,N_9660);
and U13633 (N_13633,N_7021,N_6349);
nor U13634 (N_13634,N_7232,N_9139);
xor U13635 (N_13635,N_5736,N_8872);
xnor U13636 (N_13636,N_9301,N_5885);
and U13637 (N_13637,N_7472,N_8977);
nor U13638 (N_13638,N_7379,N_8060);
nand U13639 (N_13639,N_6365,N_5198);
nand U13640 (N_13640,N_9173,N_9093);
nor U13641 (N_13641,N_8562,N_9379);
nor U13642 (N_13642,N_8838,N_6451);
and U13643 (N_13643,N_8321,N_9507);
and U13644 (N_13644,N_7102,N_5041);
nor U13645 (N_13645,N_6510,N_6825);
xnor U13646 (N_13646,N_8297,N_9082);
or U13647 (N_13647,N_5568,N_9927);
and U13648 (N_13648,N_6875,N_6649);
xnor U13649 (N_13649,N_8873,N_8547);
nor U13650 (N_13650,N_9786,N_6620);
and U13651 (N_13651,N_9998,N_9158);
or U13652 (N_13652,N_5792,N_9966);
xor U13653 (N_13653,N_6126,N_7801);
nor U13654 (N_13654,N_7485,N_8212);
nand U13655 (N_13655,N_5864,N_5368);
or U13656 (N_13656,N_5115,N_5220);
nor U13657 (N_13657,N_5801,N_6097);
nor U13658 (N_13658,N_9513,N_7660);
nand U13659 (N_13659,N_5806,N_6555);
nor U13660 (N_13660,N_9400,N_7209);
xnor U13661 (N_13661,N_6588,N_7332);
nor U13662 (N_13662,N_7154,N_9083);
or U13663 (N_13663,N_5058,N_9422);
nor U13664 (N_13664,N_9173,N_5153);
nand U13665 (N_13665,N_5873,N_6699);
xnor U13666 (N_13666,N_6618,N_5387);
or U13667 (N_13667,N_8785,N_9611);
nand U13668 (N_13668,N_7334,N_5299);
nand U13669 (N_13669,N_8803,N_5435);
or U13670 (N_13670,N_7268,N_8884);
or U13671 (N_13671,N_8328,N_6096);
and U13672 (N_13672,N_9840,N_9563);
and U13673 (N_13673,N_7376,N_9388);
nor U13674 (N_13674,N_9993,N_5333);
nand U13675 (N_13675,N_9633,N_9095);
nor U13676 (N_13676,N_7917,N_6604);
and U13677 (N_13677,N_6073,N_6419);
and U13678 (N_13678,N_5209,N_6025);
nor U13679 (N_13679,N_9744,N_5129);
nor U13680 (N_13680,N_9884,N_6070);
nand U13681 (N_13681,N_8523,N_7075);
nand U13682 (N_13682,N_6841,N_6116);
and U13683 (N_13683,N_9296,N_7765);
or U13684 (N_13684,N_5086,N_5889);
nand U13685 (N_13685,N_7845,N_8322);
and U13686 (N_13686,N_7212,N_6935);
and U13687 (N_13687,N_5088,N_7314);
nor U13688 (N_13688,N_6305,N_7517);
nor U13689 (N_13689,N_9902,N_5922);
nor U13690 (N_13690,N_7135,N_8279);
nor U13691 (N_13691,N_9051,N_8873);
nor U13692 (N_13692,N_8523,N_9594);
and U13693 (N_13693,N_5056,N_9428);
nor U13694 (N_13694,N_7154,N_9022);
and U13695 (N_13695,N_8947,N_5529);
and U13696 (N_13696,N_5751,N_6317);
or U13697 (N_13697,N_5208,N_9146);
nand U13698 (N_13698,N_5684,N_5626);
or U13699 (N_13699,N_6948,N_8764);
or U13700 (N_13700,N_6918,N_8226);
nand U13701 (N_13701,N_9019,N_8429);
nand U13702 (N_13702,N_6054,N_8622);
or U13703 (N_13703,N_6404,N_8589);
or U13704 (N_13704,N_9792,N_6844);
nor U13705 (N_13705,N_7276,N_9571);
and U13706 (N_13706,N_7673,N_9767);
or U13707 (N_13707,N_9784,N_5937);
xor U13708 (N_13708,N_9262,N_5493);
nor U13709 (N_13709,N_9662,N_7170);
or U13710 (N_13710,N_7026,N_9521);
and U13711 (N_13711,N_6438,N_5013);
or U13712 (N_13712,N_5086,N_5598);
or U13713 (N_13713,N_8932,N_9892);
xor U13714 (N_13714,N_9987,N_5255);
nor U13715 (N_13715,N_6180,N_5040);
nor U13716 (N_13716,N_8043,N_6933);
nor U13717 (N_13717,N_7334,N_8396);
or U13718 (N_13718,N_8195,N_8874);
nand U13719 (N_13719,N_6732,N_5097);
nand U13720 (N_13720,N_6226,N_6035);
nor U13721 (N_13721,N_5014,N_7525);
xnor U13722 (N_13722,N_5535,N_8840);
nand U13723 (N_13723,N_8202,N_7761);
or U13724 (N_13724,N_8755,N_8260);
xnor U13725 (N_13725,N_5972,N_9390);
xnor U13726 (N_13726,N_9469,N_6450);
nor U13727 (N_13727,N_9455,N_7308);
or U13728 (N_13728,N_5180,N_7186);
nand U13729 (N_13729,N_7368,N_6851);
xnor U13730 (N_13730,N_9483,N_9349);
nand U13731 (N_13731,N_7944,N_6487);
or U13732 (N_13732,N_6533,N_9492);
nor U13733 (N_13733,N_9216,N_7338);
and U13734 (N_13734,N_5462,N_9532);
or U13735 (N_13735,N_7578,N_9940);
nand U13736 (N_13736,N_8742,N_5778);
xor U13737 (N_13737,N_9481,N_9650);
xor U13738 (N_13738,N_8819,N_8940);
or U13739 (N_13739,N_9364,N_6505);
nor U13740 (N_13740,N_9027,N_9880);
nand U13741 (N_13741,N_9399,N_9571);
xor U13742 (N_13742,N_5270,N_6909);
nand U13743 (N_13743,N_8426,N_8993);
or U13744 (N_13744,N_6192,N_7184);
or U13745 (N_13745,N_7805,N_8931);
nand U13746 (N_13746,N_7203,N_7572);
nand U13747 (N_13747,N_8799,N_9873);
or U13748 (N_13748,N_5193,N_9562);
nor U13749 (N_13749,N_9459,N_6721);
and U13750 (N_13750,N_7398,N_6799);
nand U13751 (N_13751,N_9686,N_5777);
and U13752 (N_13752,N_8031,N_5089);
or U13753 (N_13753,N_5340,N_7242);
nand U13754 (N_13754,N_9430,N_5702);
xnor U13755 (N_13755,N_7630,N_6970);
and U13756 (N_13756,N_8844,N_8707);
or U13757 (N_13757,N_7920,N_7562);
nand U13758 (N_13758,N_7479,N_5708);
xnor U13759 (N_13759,N_9205,N_6715);
and U13760 (N_13760,N_8934,N_9894);
xor U13761 (N_13761,N_6691,N_8040);
and U13762 (N_13762,N_6315,N_9795);
and U13763 (N_13763,N_6714,N_7484);
nand U13764 (N_13764,N_6770,N_5171);
nor U13765 (N_13765,N_6580,N_6041);
and U13766 (N_13766,N_8614,N_5792);
or U13767 (N_13767,N_8158,N_7406);
nor U13768 (N_13768,N_9839,N_6521);
nor U13769 (N_13769,N_6760,N_8368);
or U13770 (N_13770,N_9393,N_7282);
nor U13771 (N_13771,N_8355,N_9741);
xnor U13772 (N_13772,N_9631,N_5310);
nor U13773 (N_13773,N_8307,N_7781);
or U13774 (N_13774,N_9335,N_9222);
or U13775 (N_13775,N_5725,N_8986);
and U13776 (N_13776,N_9579,N_8810);
or U13777 (N_13777,N_5846,N_8626);
or U13778 (N_13778,N_6950,N_8834);
xnor U13779 (N_13779,N_6000,N_7214);
nor U13780 (N_13780,N_9888,N_5969);
nor U13781 (N_13781,N_5829,N_9611);
and U13782 (N_13782,N_8560,N_5540);
nor U13783 (N_13783,N_6542,N_7035);
nor U13784 (N_13784,N_9624,N_8091);
nor U13785 (N_13785,N_8033,N_5801);
nor U13786 (N_13786,N_7271,N_5826);
nand U13787 (N_13787,N_6730,N_8542);
xor U13788 (N_13788,N_9361,N_6090);
nor U13789 (N_13789,N_7644,N_6485);
and U13790 (N_13790,N_9573,N_9564);
nor U13791 (N_13791,N_5872,N_6260);
nor U13792 (N_13792,N_6798,N_8228);
xor U13793 (N_13793,N_6292,N_8059);
and U13794 (N_13794,N_8760,N_9099);
or U13795 (N_13795,N_8040,N_6266);
and U13796 (N_13796,N_9136,N_8234);
or U13797 (N_13797,N_5403,N_6259);
xor U13798 (N_13798,N_9471,N_8558);
and U13799 (N_13799,N_5350,N_8440);
or U13800 (N_13800,N_8291,N_7211);
nand U13801 (N_13801,N_8848,N_7508);
nor U13802 (N_13802,N_7592,N_6133);
or U13803 (N_13803,N_7919,N_7703);
or U13804 (N_13804,N_5921,N_8678);
or U13805 (N_13805,N_8277,N_5605);
xor U13806 (N_13806,N_5654,N_6294);
nand U13807 (N_13807,N_9288,N_8560);
and U13808 (N_13808,N_8200,N_7571);
or U13809 (N_13809,N_9306,N_6265);
or U13810 (N_13810,N_8668,N_6327);
or U13811 (N_13811,N_8296,N_5219);
xor U13812 (N_13812,N_8450,N_7671);
or U13813 (N_13813,N_6783,N_6163);
nor U13814 (N_13814,N_8690,N_8219);
or U13815 (N_13815,N_7160,N_5375);
or U13816 (N_13816,N_6135,N_9666);
xnor U13817 (N_13817,N_8529,N_8407);
nand U13818 (N_13818,N_6451,N_7269);
or U13819 (N_13819,N_9800,N_8979);
nand U13820 (N_13820,N_8670,N_8180);
nand U13821 (N_13821,N_5781,N_5444);
and U13822 (N_13822,N_8641,N_6786);
and U13823 (N_13823,N_5917,N_9048);
xor U13824 (N_13824,N_7845,N_9593);
or U13825 (N_13825,N_7970,N_8171);
nor U13826 (N_13826,N_9597,N_6499);
nand U13827 (N_13827,N_7723,N_7619);
nor U13828 (N_13828,N_8865,N_7232);
xnor U13829 (N_13829,N_7593,N_6414);
nand U13830 (N_13830,N_6447,N_5435);
xnor U13831 (N_13831,N_8740,N_9140);
and U13832 (N_13832,N_5084,N_7076);
xor U13833 (N_13833,N_9328,N_9182);
nand U13834 (N_13834,N_6944,N_7010);
or U13835 (N_13835,N_9205,N_7400);
xor U13836 (N_13836,N_6937,N_5931);
xnor U13837 (N_13837,N_6089,N_9309);
and U13838 (N_13838,N_6924,N_7474);
or U13839 (N_13839,N_6320,N_7968);
and U13840 (N_13840,N_6427,N_7731);
nor U13841 (N_13841,N_7433,N_9410);
nor U13842 (N_13842,N_5354,N_9733);
nand U13843 (N_13843,N_5341,N_6204);
nand U13844 (N_13844,N_7248,N_5394);
or U13845 (N_13845,N_8425,N_5241);
nand U13846 (N_13846,N_5858,N_9190);
or U13847 (N_13847,N_8229,N_8339);
xnor U13848 (N_13848,N_9831,N_6555);
nand U13849 (N_13849,N_7120,N_9154);
and U13850 (N_13850,N_5250,N_8785);
xor U13851 (N_13851,N_5134,N_5380);
nand U13852 (N_13852,N_7377,N_5646);
nor U13853 (N_13853,N_6657,N_7635);
nor U13854 (N_13854,N_7141,N_5440);
nand U13855 (N_13855,N_6255,N_9853);
xor U13856 (N_13856,N_9017,N_9733);
xor U13857 (N_13857,N_9680,N_7650);
or U13858 (N_13858,N_9073,N_7671);
xnor U13859 (N_13859,N_9147,N_9825);
xnor U13860 (N_13860,N_8523,N_5285);
or U13861 (N_13861,N_8303,N_8197);
nand U13862 (N_13862,N_5995,N_9885);
xnor U13863 (N_13863,N_6952,N_6494);
nand U13864 (N_13864,N_7087,N_8811);
and U13865 (N_13865,N_9778,N_6381);
nor U13866 (N_13866,N_6517,N_9499);
xnor U13867 (N_13867,N_7505,N_7056);
nand U13868 (N_13868,N_7867,N_6197);
and U13869 (N_13869,N_7860,N_7422);
nor U13870 (N_13870,N_6338,N_7975);
or U13871 (N_13871,N_9717,N_9914);
nand U13872 (N_13872,N_6077,N_9955);
nor U13873 (N_13873,N_5221,N_9574);
or U13874 (N_13874,N_7171,N_9211);
xnor U13875 (N_13875,N_9008,N_5078);
or U13876 (N_13876,N_5763,N_7620);
nand U13877 (N_13877,N_5202,N_5198);
xor U13878 (N_13878,N_6385,N_8847);
xor U13879 (N_13879,N_5046,N_5522);
and U13880 (N_13880,N_5288,N_8922);
xnor U13881 (N_13881,N_5097,N_8208);
nor U13882 (N_13882,N_7705,N_6118);
nor U13883 (N_13883,N_7665,N_9072);
nor U13884 (N_13884,N_5175,N_8474);
and U13885 (N_13885,N_7620,N_7256);
and U13886 (N_13886,N_8120,N_6786);
and U13887 (N_13887,N_6640,N_6312);
and U13888 (N_13888,N_8296,N_9160);
nor U13889 (N_13889,N_5346,N_7645);
nor U13890 (N_13890,N_8887,N_9047);
nor U13891 (N_13891,N_7250,N_9883);
nand U13892 (N_13892,N_8109,N_7637);
and U13893 (N_13893,N_8156,N_9528);
and U13894 (N_13894,N_8542,N_8866);
or U13895 (N_13895,N_8718,N_9820);
nor U13896 (N_13896,N_9295,N_8932);
xor U13897 (N_13897,N_7317,N_7628);
nand U13898 (N_13898,N_9913,N_5682);
nand U13899 (N_13899,N_6001,N_8002);
or U13900 (N_13900,N_6605,N_9986);
nand U13901 (N_13901,N_9509,N_7699);
and U13902 (N_13902,N_9006,N_7696);
nor U13903 (N_13903,N_8472,N_8791);
xor U13904 (N_13904,N_8347,N_5543);
nor U13905 (N_13905,N_6516,N_8207);
xnor U13906 (N_13906,N_8682,N_6189);
and U13907 (N_13907,N_6487,N_8969);
or U13908 (N_13908,N_7098,N_8123);
nand U13909 (N_13909,N_5339,N_7502);
or U13910 (N_13910,N_8264,N_6070);
or U13911 (N_13911,N_6106,N_7482);
nand U13912 (N_13912,N_6639,N_5470);
xor U13913 (N_13913,N_7450,N_5636);
nand U13914 (N_13914,N_5391,N_6154);
and U13915 (N_13915,N_8961,N_9016);
and U13916 (N_13916,N_5551,N_6300);
xnor U13917 (N_13917,N_5876,N_8087);
xnor U13918 (N_13918,N_5447,N_8182);
nor U13919 (N_13919,N_9697,N_8295);
nand U13920 (N_13920,N_7637,N_8285);
nand U13921 (N_13921,N_9700,N_6826);
nor U13922 (N_13922,N_6362,N_8666);
or U13923 (N_13923,N_5220,N_7112);
or U13924 (N_13924,N_7779,N_5323);
and U13925 (N_13925,N_5312,N_5363);
nor U13926 (N_13926,N_7177,N_7077);
or U13927 (N_13927,N_9902,N_8951);
nand U13928 (N_13928,N_8566,N_6854);
and U13929 (N_13929,N_6964,N_5205);
nor U13930 (N_13930,N_7373,N_9056);
nor U13931 (N_13931,N_7189,N_8174);
nor U13932 (N_13932,N_9046,N_6338);
xor U13933 (N_13933,N_8461,N_7881);
and U13934 (N_13934,N_8385,N_5523);
or U13935 (N_13935,N_6370,N_7204);
xnor U13936 (N_13936,N_6431,N_8039);
or U13937 (N_13937,N_7030,N_7674);
xor U13938 (N_13938,N_7914,N_5637);
or U13939 (N_13939,N_7902,N_5999);
xor U13940 (N_13940,N_6983,N_7582);
nand U13941 (N_13941,N_7001,N_5021);
or U13942 (N_13942,N_8160,N_6413);
nand U13943 (N_13943,N_8725,N_5299);
nor U13944 (N_13944,N_9108,N_8722);
or U13945 (N_13945,N_5835,N_5012);
nor U13946 (N_13946,N_6258,N_6075);
nor U13947 (N_13947,N_6434,N_9830);
or U13948 (N_13948,N_9414,N_6574);
or U13949 (N_13949,N_9050,N_9973);
xor U13950 (N_13950,N_8641,N_6318);
xnor U13951 (N_13951,N_6044,N_6230);
nor U13952 (N_13952,N_7519,N_5013);
xor U13953 (N_13953,N_5404,N_8925);
xnor U13954 (N_13954,N_9027,N_9909);
and U13955 (N_13955,N_5100,N_6109);
xnor U13956 (N_13956,N_8791,N_6223);
or U13957 (N_13957,N_8449,N_8197);
nor U13958 (N_13958,N_8547,N_5338);
nor U13959 (N_13959,N_9205,N_5826);
and U13960 (N_13960,N_9472,N_7779);
nand U13961 (N_13961,N_5524,N_8013);
and U13962 (N_13962,N_6101,N_5783);
nand U13963 (N_13963,N_6898,N_5520);
nand U13964 (N_13964,N_8262,N_9416);
nand U13965 (N_13965,N_8877,N_5564);
and U13966 (N_13966,N_7067,N_5672);
xnor U13967 (N_13967,N_8352,N_5321);
xor U13968 (N_13968,N_8334,N_8182);
and U13969 (N_13969,N_7995,N_6041);
xnor U13970 (N_13970,N_7230,N_5957);
and U13971 (N_13971,N_6303,N_8662);
nor U13972 (N_13972,N_8492,N_9762);
xnor U13973 (N_13973,N_7005,N_5443);
nand U13974 (N_13974,N_9539,N_8126);
nand U13975 (N_13975,N_5992,N_9777);
or U13976 (N_13976,N_6789,N_5190);
or U13977 (N_13977,N_8465,N_6656);
nor U13978 (N_13978,N_8828,N_5994);
and U13979 (N_13979,N_8829,N_9837);
and U13980 (N_13980,N_7226,N_8697);
nor U13981 (N_13981,N_8281,N_9075);
nor U13982 (N_13982,N_5320,N_8211);
and U13983 (N_13983,N_8681,N_6988);
or U13984 (N_13984,N_7961,N_5840);
nand U13985 (N_13985,N_6718,N_7194);
and U13986 (N_13986,N_5722,N_5995);
nand U13987 (N_13987,N_9264,N_7659);
xor U13988 (N_13988,N_8071,N_5040);
nand U13989 (N_13989,N_7430,N_9021);
nand U13990 (N_13990,N_6937,N_6059);
nand U13991 (N_13991,N_7984,N_7520);
and U13992 (N_13992,N_8995,N_9077);
nand U13993 (N_13993,N_5092,N_7706);
nor U13994 (N_13994,N_9577,N_8846);
nand U13995 (N_13995,N_7320,N_8657);
xnor U13996 (N_13996,N_6479,N_7867);
nand U13997 (N_13997,N_8879,N_7412);
or U13998 (N_13998,N_6003,N_7578);
nor U13999 (N_13999,N_8241,N_7222);
nor U14000 (N_14000,N_8479,N_9892);
or U14001 (N_14001,N_9862,N_8159);
nand U14002 (N_14002,N_5012,N_8496);
xor U14003 (N_14003,N_5816,N_8143);
nor U14004 (N_14004,N_9715,N_8787);
or U14005 (N_14005,N_6033,N_5201);
or U14006 (N_14006,N_6877,N_8440);
or U14007 (N_14007,N_9528,N_9205);
or U14008 (N_14008,N_5636,N_6103);
xnor U14009 (N_14009,N_5635,N_5234);
and U14010 (N_14010,N_9048,N_9399);
xnor U14011 (N_14011,N_8475,N_9536);
and U14012 (N_14012,N_9345,N_7549);
and U14013 (N_14013,N_5722,N_6214);
nand U14014 (N_14014,N_9308,N_9931);
xnor U14015 (N_14015,N_5092,N_9505);
nor U14016 (N_14016,N_6880,N_7498);
or U14017 (N_14017,N_6354,N_6503);
or U14018 (N_14018,N_7908,N_5932);
or U14019 (N_14019,N_5914,N_9493);
nand U14020 (N_14020,N_9246,N_6309);
nor U14021 (N_14021,N_5762,N_9370);
xor U14022 (N_14022,N_7660,N_9785);
or U14023 (N_14023,N_6446,N_7470);
or U14024 (N_14024,N_7191,N_9382);
or U14025 (N_14025,N_7323,N_8533);
nor U14026 (N_14026,N_5332,N_7001);
xor U14027 (N_14027,N_9055,N_7775);
and U14028 (N_14028,N_5931,N_9076);
nor U14029 (N_14029,N_7920,N_7721);
or U14030 (N_14030,N_6020,N_9487);
and U14031 (N_14031,N_5905,N_7712);
and U14032 (N_14032,N_7599,N_5987);
or U14033 (N_14033,N_8434,N_9615);
nor U14034 (N_14034,N_7320,N_9226);
and U14035 (N_14035,N_7961,N_9115);
or U14036 (N_14036,N_7475,N_7576);
and U14037 (N_14037,N_9400,N_9294);
nor U14038 (N_14038,N_5959,N_8912);
or U14039 (N_14039,N_7068,N_6597);
nand U14040 (N_14040,N_8504,N_9511);
and U14041 (N_14041,N_8035,N_6501);
xor U14042 (N_14042,N_7416,N_5018);
nor U14043 (N_14043,N_8797,N_6308);
xnor U14044 (N_14044,N_9771,N_5935);
or U14045 (N_14045,N_8559,N_7076);
xnor U14046 (N_14046,N_8049,N_7071);
or U14047 (N_14047,N_8049,N_7277);
or U14048 (N_14048,N_7216,N_8891);
and U14049 (N_14049,N_8406,N_9958);
nor U14050 (N_14050,N_6162,N_7714);
or U14051 (N_14051,N_8629,N_5749);
and U14052 (N_14052,N_9531,N_8487);
or U14053 (N_14053,N_8444,N_8024);
and U14054 (N_14054,N_9937,N_6569);
or U14055 (N_14055,N_5544,N_7907);
and U14056 (N_14056,N_5240,N_5079);
or U14057 (N_14057,N_7224,N_5619);
nand U14058 (N_14058,N_6875,N_9626);
or U14059 (N_14059,N_5373,N_6532);
or U14060 (N_14060,N_5217,N_8206);
xnor U14061 (N_14061,N_6868,N_6541);
or U14062 (N_14062,N_9642,N_5824);
nand U14063 (N_14063,N_8377,N_6803);
xor U14064 (N_14064,N_5407,N_7836);
and U14065 (N_14065,N_6031,N_5719);
and U14066 (N_14066,N_7819,N_9738);
xor U14067 (N_14067,N_8781,N_7076);
and U14068 (N_14068,N_9832,N_5932);
and U14069 (N_14069,N_5729,N_6225);
xor U14070 (N_14070,N_6527,N_6383);
or U14071 (N_14071,N_7013,N_6573);
xor U14072 (N_14072,N_5164,N_5569);
nand U14073 (N_14073,N_8198,N_5330);
and U14074 (N_14074,N_9271,N_8370);
nor U14075 (N_14075,N_9011,N_9058);
nand U14076 (N_14076,N_6272,N_8960);
nor U14077 (N_14077,N_9037,N_8783);
and U14078 (N_14078,N_5422,N_5171);
nor U14079 (N_14079,N_6213,N_9803);
nor U14080 (N_14080,N_6427,N_8793);
nor U14081 (N_14081,N_8169,N_5188);
or U14082 (N_14082,N_8314,N_7043);
nand U14083 (N_14083,N_7435,N_6481);
nand U14084 (N_14084,N_5795,N_5490);
xor U14085 (N_14085,N_8464,N_7602);
and U14086 (N_14086,N_5554,N_8493);
xnor U14087 (N_14087,N_5164,N_6888);
or U14088 (N_14088,N_5773,N_6167);
or U14089 (N_14089,N_7886,N_6123);
nor U14090 (N_14090,N_9437,N_6154);
and U14091 (N_14091,N_8793,N_5296);
xnor U14092 (N_14092,N_6584,N_9577);
xnor U14093 (N_14093,N_6198,N_9451);
nand U14094 (N_14094,N_7254,N_9120);
xnor U14095 (N_14095,N_6346,N_8426);
or U14096 (N_14096,N_7350,N_5851);
xor U14097 (N_14097,N_6249,N_9753);
xnor U14098 (N_14098,N_5398,N_5933);
nor U14099 (N_14099,N_8329,N_6855);
and U14100 (N_14100,N_5390,N_5594);
nand U14101 (N_14101,N_8803,N_8960);
or U14102 (N_14102,N_8462,N_7776);
nand U14103 (N_14103,N_7659,N_7708);
and U14104 (N_14104,N_6837,N_6052);
and U14105 (N_14105,N_7490,N_8871);
nand U14106 (N_14106,N_9748,N_8117);
nor U14107 (N_14107,N_6003,N_8611);
xnor U14108 (N_14108,N_5147,N_6471);
nand U14109 (N_14109,N_8911,N_6346);
and U14110 (N_14110,N_9675,N_7502);
or U14111 (N_14111,N_6225,N_5002);
or U14112 (N_14112,N_7311,N_6846);
nand U14113 (N_14113,N_6705,N_8696);
and U14114 (N_14114,N_5611,N_7959);
nand U14115 (N_14115,N_8845,N_7347);
nor U14116 (N_14116,N_7343,N_8860);
or U14117 (N_14117,N_9125,N_8994);
nand U14118 (N_14118,N_5191,N_8747);
xnor U14119 (N_14119,N_6054,N_5685);
nand U14120 (N_14120,N_7972,N_9696);
or U14121 (N_14121,N_7523,N_7484);
or U14122 (N_14122,N_6083,N_9981);
xnor U14123 (N_14123,N_5314,N_8262);
nor U14124 (N_14124,N_5018,N_9910);
and U14125 (N_14125,N_5300,N_5117);
nor U14126 (N_14126,N_5693,N_7689);
or U14127 (N_14127,N_7797,N_8468);
xor U14128 (N_14128,N_6817,N_8021);
xor U14129 (N_14129,N_8421,N_9431);
xnor U14130 (N_14130,N_6661,N_9267);
xor U14131 (N_14131,N_8309,N_9812);
and U14132 (N_14132,N_8406,N_7178);
nand U14133 (N_14133,N_8350,N_9439);
xnor U14134 (N_14134,N_9751,N_8754);
or U14135 (N_14135,N_6193,N_9397);
and U14136 (N_14136,N_6356,N_8265);
xor U14137 (N_14137,N_5594,N_7915);
nor U14138 (N_14138,N_9711,N_9351);
and U14139 (N_14139,N_8973,N_8758);
nor U14140 (N_14140,N_6125,N_9253);
nand U14141 (N_14141,N_9028,N_7110);
nor U14142 (N_14142,N_5806,N_5566);
and U14143 (N_14143,N_7372,N_6940);
nor U14144 (N_14144,N_9307,N_9882);
and U14145 (N_14145,N_8426,N_5024);
nor U14146 (N_14146,N_8448,N_6902);
or U14147 (N_14147,N_9228,N_6393);
or U14148 (N_14148,N_7657,N_8157);
or U14149 (N_14149,N_9465,N_9384);
nor U14150 (N_14150,N_7206,N_7820);
and U14151 (N_14151,N_6869,N_7090);
or U14152 (N_14152,N_5884,N_9414);
and U14153 (N_14153,N_8875,N_7542);
xor U14154 (N_14154,N_5433,N_7727);
and U14155 (N_14155,N_6913,N_8689);
and U14156 (N_14156,N_5641,N_8493);
nand U14157 (N_14157,N_7236,N_7437);
or U14158 (N_14158,N_8874,N_8558);
xnor U14159 (N_14159,N_8413,N_7455);
and U14160 (N_14160,N_8413,N_8279);
nor U14161 (N_14161,N_7170,N_8014);
or U14162 (N_14162,N_6864,N_9073);
or U14163 (N_14163,N_7924,N_5553);
nand U14164 (N_14164,N_9894,N_5294);
or U14165 (N_14165,N_7884,N_5093);
or U14166 (N_14166,N_7578,N_7425);
or U14167 (N_14167,N_8788,N_8912);
nor U14168 (N_14168,N_9098,N_9623);
xor U14169 (N_14169,N_7061,N_8410);
or U14170 (N_14170,N_5277,N_9129);
xor U14171 (N_14171,N_9295,N_5773);
or U14172 (N_14172,N_5988,N_8058);
or U14173 (N_14173,N_7676,N_8514);
and U14174 (N_14174,N_7282,N_5104);
xor U14175 (N_14175,N_6405,N_5372);
nor U14176 (N_14176,N_5107,N_8909);
and U14177 (N_14177,N_9943,N_5689);
nor U14178 (N_14178,N_5117,N_7393);
nor U14179 (N_14179,N_6407,N_5241);
xor U14180 (N_14180,N_5070,N_8514);
xor U14181 (N_14181,N_5557,N_5738);
nand U14182 (N_14182,N_8345,N_8124);
and U14183 (N_14183,N_9473,N_7720);
nand U14184 (N_14184,N_9734,N_7338);
nor U14185 (N_14185,N_7943,N_7904);
or U14186 (N_14186,N_5978,N_5063);
nand U14187 (N_14187,N_6997,N_7398);
nor U14188 (N_14188,N_7390,N_7457);
nor U14189 (N_14189,N_6138,N_7674);
xnor U14190 (N_14190,N_7540,N_9548);
or U14191 (N_14191,N_6870,N_8421);
nand U14192 (N_14192,N_6443,N_5723);
nor U14193 (N_14193,N_7384,N_9478);
xnor U14194 (N_14194,N_8712,N_9984);
or U14195 (N_14195,N_9081,N_5929);
nand U14196 (N_14196,N_8312,N_8644);
xor U14197 (N_14197,N_5387,N_6829);
xor U14198 (N_14198,N_8579,N_6367);
nor U14199 (N_14199,N_5362,N_8584);
nor U14200 (N_14200,N_8537,N_8488);
nor U14201 (N_14201,N_9511,N_8298);
xor U14202 (N_14202,N_7230,N_9448);
and U14203 (N_14203,N_8642,N_5457);
xnor U14204 (N_14204,N_9146,N_7088);
nor U14205 (N_14205,N_5278,N_6001);
and U14206 (N_14206,N_8959,N_5286);
or U14207 (N_14207,N_6504,N_9163);
nor U14208 (N_14208,N_9767,N_7849);
xnor U14209 (N_14209,N_6482,N_5355);
nor U14210 (N_14210,N_5050,N_8127);
or U14211 (N_14211,N_5149,N_9245);
nand U14212 (N_14212,N_7334,N_7778);
or U14213 (N_14213,N_9118,N_6892);
nand U14214 (N_14214,N_9564,N_5834);
and U14215 (N_14215,N_5994,N_8508);
and U14216 (N_14216,N_8507,N_9130);
or U14217 (N_14217,N_5364,N_5555);
nand U14218 (N_14218,N_8559,N_7730);
and U14219 (N_14219,N_9465,N_7828);
xor U14220 (N_14220,N_5672,N_5609);
nor U14221 (N_14221,N_9391,N_7541);
nor U14222 (N_14222,N_7185,N_5206);
nand U14223 (N_14223,N_9899,N_7862);
or U14224 (N_14224,N_6623,N_5521);
nand U14225 (N_14225,N_8575,N_8926);
or U14226 (N_14226,N_8431,N_8600);
and U14227 (N_14227,N_5624,N_5584);
nor U14228 (N_14228,N_7663,N_8832);
and U14229 (N_14229,N_8161,N_5727);
or U14230 (N_14230,N_8403,N_6205);
and U14231 (N_14231,N_9274,N_9616);
and U14232 (N_14232,N_6116,N_9770);
nor U14233 (N_14233,N_9975,N_5519);
or U14234 (N_14234,N_6973,N_7926);
nand U14235 (N_14235,N_9377,N_6182);
nand U14236 (N_14236,N_9904,N_6630);
or U14237 (N_14237,N_8388,N_9965);
or U14238 (N_14238,N_6430,N_7950);
xnor U14239 (N_14239,N_9220,N_7192);
xor U14240 (N_14240,N_7014,N_8561);
or U14241 (N_14241,N_9653,N_8518);
nor U14242 (N_14242,N_5713,N_6080);
nor U14243 (N_14243,N_8463,N_5128);
nand U14244 (N_14244,N_8772,N_9351);
nor U14245 (N_14245,N_9492,N_5764);
nand U14246 (N_14246,N_7348,N_8161);
or U14247 (N_14247,N_9706,N_5861);
or U14248 (N_14248,N_6574,N_6226);
nor U14249 (N_14249,N_5000,N_9442);
nand U14250 (N_14250,N_8918,N_6693);
nor U14251 (N_14251,N_7304,N_6712);
xnor U14252 (N_14252,N_6996,N_9656);
nor U14253 (N_14253,N_9759,N_7009);
or U14254 (N_14254,N_6521,N_6403);
or U14255 (N_14255,N_8475,N_9258);
and U14256 (N_14256,N_7738,N_7235);
or U14257 (N_14257,N_9169,N_9280);
nor U14258 (N_14258,N_7932,N_9125);
nand U14259 (N_14259,N_6102,N_8238);
or U14260 (N_14260,N_7512,N_7026);
xor U14261 (N_14261,N_6559,N_9026);
or U14262 (N_14262,N_8562,N_5934);
xor U14263 (N_14263,N_5166,N_8783);
nor U14264 (N_14264,N_6837,N_6987);
nand U14265 (N_14265,N_7657,N_8682);
or U14266 (N_14266,N_7730,N_5156);
nor U14267 (N_14267,N_5469,N_8898);
or U14268 (N_14268,N_7995,N_5175);
or U14269 (N_14269,N_6972,N_5243);
and U14270 (N_14270,N_6442,N_8566);
and U14271 (N_14271,N_7295,N_8419);
and U14272 (N_14272,N_6857,N_5823);
or U14273 (N_14273,N_9628,N_6875);
nand U14274 (N_14274,N_6615,N_8494);
or U14275 (N_14275,N_7167,N_5409);
or U14276 (N_14276,N_9852,N_7926);
nor U14277 (N_14277,N_7662,N_6618);
nand U14278 (N_14278,N_6041,N_7956);
nand U14279 (N_14279,N_9207,N_6408);
and U14280 (N_14280,N_6874,N_8763);
nand U14281 (N_14281,N_8342,N_9819);
nand U14282 (N_14282,N_6724,N_8926);
nor U14283 (N_14283,N_5373,N_6419);
nor U14284 (N_14284,N_6512,N_5076);
or U14285 (N_14285,N_9115,N_7716);
and U14286 (N_14286,N_8223,N_5407);
xnor U14287 (N_14287,N_7014,N_5214);
xor U14288 (N_14288,N_8730,N_8587);
or U14289 (N_14289,N_6490,N_6759);
and U14290 (N_14290,N_6614,N_8855);
nor U14291 (N_14291,N_7564,N_5058);
and U14292 (N_14292,N_9392,N_8880);
xor U14293 (N_14293,N_5294,N_6180);
or U14294 (N_14294,N_5287,N_6871);
nor U14295 (N_14295,N_7993,N_9423);
and U14296 (N_14296,N_5164,N_9564);
nand U14297 (N_14297,N_9597,N_5663);
xor U14298 (N_14298,N_6672,N_6591);
nor U14299 (N_14299,N_9518,N_7213);
xor U14300 (N_14300,N_6947,N_8825);
nor U14301 (N_14301,N_7439,N_7195);
xnor U14302 (N_14302,N_8430,N_5068);
and U14303 (N_14303,N_8206,N_8316);
or U14304 (N_14304,N_5500,N_6925);
nand U14305 (N_14305,N_8548,N_5867);
nor U14306 (N_14306,N_6527,N_6147);
nand U14307 (N_14307,N_6911,N_7355);
and U14308 (N_14308,N_8579,N_7348);
nor U14309 (N_14309,N_8168,N_8008);
xnor U14310 (N_14310,N_8097,N_5747);
or U14311 (N_14311,N_9128,N_6423);
or U14312 (N_14312,N_7525,N_9873);
nor U14313 (N_14313,N_7397,N_9658);
xor U14314 (N_14314,N_8757,N_5762);
or U14315 (N_14315,N_8901,N_6675);
nand U14316 (N_14316,N_8805,N_5243);
xor U14317 (N_14317,N_9119,N_9917);
or U14318 (N_14318,N_8222,N_8907);
nor U14319 (N_14319,N_7426,N_7196);
nor U14320 (N_14320,N_6143,N_9143);
nor U14321 (N_14321,N_5762,N_8743);
xor U14322 (N_14322,N_9988,N_9574);
and U14323 (N_14323,N_8174,N_5958);
or U14324 (N_14324,N_7683,N_8517);
nor U14325 (N_14325,N_9648,N_8193);
nor U14326 (N_14326,N_5708,N_8220);
nor U14327 (N_14327,N_8313,N_7480);
nor U14328 (N_14328,N_7986,N_9767);
nand U14329 (N_14329,N_7983,N_6020);
nand U14330 (N_14330,N_5164,N_5810);
nor U14331 (N_14331,N_6738,N_5452);
nand U14332 (N_14332,N_6886,N_7082);
nor U14333 (N_14333,N_6462,N_7512);
nand U14334 (N_14334,N_8271,N_6928);
xor U14335 (N_14335,N_6227,N_8688);
nand U14336 (N_14336,N_8261,N_8670);
nand U14337 (N_14337,N_9902,N_6455);
or U14338 (N_14338,N_7045,N_8548);
and U14339 (N_14339,N_8824,N_7478);
nand U14340 (N_14340,N_6885,N_9143);
nor U14341 (N_14341,N_5035,N_7341);
xnor U14342 (N_14342,N_5710,N_8962);
and U14343 (N_14343,N_8143,N_5440);
xor U14344 (N_14344,N_6770,N_5712);
xnor U14345 (N_14345,N_6820,N_5017);
or U14346 (N_14346,N_6868,N_6715);
xor U14347 (N_14347,N_6476,N_9336);
nand U14348 (N_14348,N_7814,N_8514);
and U14349 (N_14349,N_9408,N_5076);
and U14350 (N_14350,N_5869,N_9006);
or U14351 (N_14351,N_8931,N_9980);
or U14352 (N_14352,N_5000,N_7851);
nand U14353 (N_14353,N_9170,N_8160);
nand U14354 (N_14354,N_9859,N_5999);
or U14355 (N_14355,N_5039,N_6567);
xnor U14356 (N_14356,N_6505,N_9298);
and U14357 (N_14357,N_8775,N_6367);
nor U14358 (N_14358,N_8279,N_5229);
xor U14359 (N_14359,N_9457,N_8749);
or U14360 (N_14360,N_8255,N_8653);
nand U14361 (N_14361,N_6099,N_5245);
nand U14362 (N_14362,N_8963,N_9685);
xnor U14363 (N_14363,N_8790,N_5275);
nor U14364 (N_14364,N_9669,N_5703);
xnor U14365 (N_14365,N_8051,N_5518);
or U14366 (N_14366,N_8313,N_6626);
xor U14367 (N_14367,N_8035,N_6607);
and U14368 (N_14368,N_9856,N_8971);
or U14369 (N_14369,N_9853,N_8151);
and U14370 (N_14370,N_6057,N_8088);
and U14371 (N_14371,N_7971,N_8193);
nor U14372 (N_14372,N_8087,N_6656);
xnor U14373 (N_14373,N_6902,N_7260);
or U14374 (N_14374,N_9041,N_7481);
and U14375 (N_14375,N_6465,N_9044);
or U14376 (N_14376,N_9834,N_8732);
and U14377 (N_14377,N_5398,N_9451);
or U14378 (N_14378,N_8766,N_9263);
and U14379 (N_14379,N_6210,N_7770);
nor U14380 (N_14380,N_9737,N_5940);
or U14381 (N_14381,N_9020,N_5078);
or U14382 (N_14382,N_7571,N_8077);
and U14383 (N_14383,N_7101,N_6057);
nand U14384 (N_14384,N_7502,N_9186);
xor U14385 (N_14385,N_6454,N_8688);
and U14386 (N_14386,N_8387,N_7401);
nor U14387 (N_14387,N_7757,N_7437);
or U14388 (N_14388,N_8160,N_9324);
or U14389 (N_14389,N_8259,N_9049);
or U14390 (N_14390,N_7011,N_5598);
and U14391 (N_14391,N_5502,N_6760);
and U14392 (N_14392,N_9489,N_9658);
nand U14393 (N_14393,N_5486,N_7882);
xor U14394 (N_14394,N_6457,N_8769);
nor U14395 (N_14395,N_5144,N_6808);
nand U14396 (N_14396,N_9074,N_8302);
and U14397 (N_14397,N_7535,N_7689);
xor U14398 (N_14398,N_8593,N_8758);
xor U14399 (N_14399,N_8471,N_9262);
nand U14400 (N_14400,N_7020,N_5294);
xor U14401 (N_14401,N_5756,N_6557);
and U14402 (N_14402,N_6240,N_8051);
xor U14403 (N_14403,N_6488,N_7397);
or U14404 (N_14404,N_5830,N_5351);
nor U14405 (N_14405,N_9938,N_8163);
and U14406 (N_14406,N_8764,N_7240);
and U14407 (N_14407,N_8437,N_8546);
nor U14408 (N_14408,N_6984,N_5802);
xnor U14409 (N_14409,N_7630,N_7773);
nand U14410 (N_14410,N_6021,N_6788);
xnor U14411 (N_14411,N_5179,N_5319);
or U14412 (N_14412,N_7529,N_6214);
nor U14413 (N_14413,N_7824,N_9817);
xor U14414 (N_14414,N_6930,N_6482);
and U14415 (N_14415,N_6990,N_9302);
or U14416 (N_14416,N_5769,N_7043);
and U14417 (N_14417,N_5269,N_5615);
xor U14418 (N_14418,N_8155,N_9105);
or U14419 (N_14419,N_5247,N_8095);
nor U14420 (N_14420,N_8797,N_9021);
and U14421 (N_14421,N_7980,N_6015);
and U14422 (N_14422,N_9064,N_6323);
nand U14423 (N_14423,N_5651,N_6513);
or U14424 (N_14424,N_9458,N_9139);
or U14425 (N_14425,N_8678,N_7395);
or U14426 (N_14426,N_6354,N_5404);
xor U14427 (N_14427,N_8958,N_8143);
nand U14428 (N_14428,N_9547,N_5305);
nor U14429 (N_14429,N_8260,N_6137);
and U14430 (N_14430,N_5545,N_8428);
xnor U14431 (N_14431,N_7302,N_9379);
and U14432 (N_14432,N_5826,N_5777);
and U14433 (N_14433,N_5499,N_6380);
nor U14434 (N_14434,N_6401,N_6542);
and U14435 (N_14435,N_9768,N_9493);
nor U14436 (N_14436,N_8561,N_7832);
or U14437 (N_14437,N_8444,N_6097);
nor U14438 (N_14438,N_6979,N_5584);
xor U14439 (N_14439,N_5378,N_7684);
xor U14440 (N_14440,N_5560,N_9387);
and U14441 (N_14441,N_8899,N_5469);
xor U14442 (N_14442,N_7412,N_9731);
xor U14443 (N_14443,N_5015,N_5835);
nand U14444 (N_14444,N_5396,N_6957);
xor U14445 (N_14445,N_6751,N_9049);
xnor U14446 (N_14446,N_6859,N_9456);
and U14447 (N_14447,N_5089,N_7156);
nor U14448 (N_14448,N_8622,N_9015);
nand U14449 (N_14449,N_9547,N_6730);
nor U14450 (N_14450,N_5043,N_7482);
and U14451 (N_14451,N_7646,N_7733);
xnor U14452 (N_14452,N_8470,N_5682);
xnor U14453 (N_14453,N_5793,N_8999);
nand U14454 (N_14454,N_7241,N_8787);
or U14455 (N_14455,N_5866,N_8070);
xor U14456 (N_14456,N_8588,N_9724);
nand U14457 (N_14457,N_7341,N_6749);
and U14458 (N_14458,N_6737,N_8432);
and U14459 (N_14459,N_5428,N_9993);
xnor U14460 (N_14460,N_5268,N_6308);
nor U14461 (N_14461,N_9294,N_6735);
or U14462 (N_14462,N_7729,N_8773);
nand U14463 (N_14463,N_9061,N_5698);
xnor U14464 (N_14464,N_5015,N_7642);
xnor U14465 (N_14465,N_9353,N_9894);
nor U14466 (N_14466,N_6089,N_6356);
nand U14467 (N_14467,N_6014,N_8708);
and U14468 (N_14468,N_9662,N_8753);
nor U14469 (N_14469,N_7692,N_8847);
nand U14470 (N_14470,N_9140,N_8086);
nor U14471 (N_14471,N_5572,N_5995);
xnor U14472 (N_14472,N_9548,N_9376);
or U14473 (N_14473,N_5152,N_5598);
nor U14474 (N_14474,N_9094,N_5433);
nor U14475 (N_14475,N_5179,N_9559);
xor U14476 (N_14476,N_8451,N_5203);
xor U14477 (N_14477,N_9957,N_5573);
nor U14478 (N_14478,N_5923,N_9933);
nand U14479 (N_14479,N_6131,N_8697);
xor U14480 (N_14480,N_7793,N_8286);
nand U14481 (N_14481,N_7098,N_8701);
or U14482 (N_14482,N_6098,N_9873);
xor U14483 (N_14483,N_5221,N_8485);
xnor U14484 (N_14484,N_9132,N_5400);
or U14485 (N_14485,N_9157,N_5338);
nand U14486 (N_14486,N_5739,N_5873);
nor U14487 (N_14487,N_8382,N_7466);
nor U14488 (N_14488,N_6575,N_8940);
xor U14489 (N_14489,N_7436,N_5478);
nand U14490 (N_14490,N_5074,N_6479);
or U14491 (N_14491,N_7042,N_9869);
or U14492 (N_14492,N_8513,N_5610);
nor U14493 (N_14493,N_8350,N_6598);
or U14494 (N_14494,N_6008,N_6068);
or U14495 (N_14495,N_8099,N_5102);
nor U14496 (N_14496,N_7453,N_5721);
xnor U14497 (N_14497,N_5313,N_5113);
and U14498 (N_14498,N_9226,N_5313);
nand U14499 (N_14499,N_6487,N_9653);
xor U14500 (N_14500,N_8193,N_6475);
nor U14501 (N_14501,N_8573,N_6833);
and U14502 (N_14502,N_9229,N_7361);
nor U14503 (N_14503,N_6748,N_6797);
xnor U14504 (N_14504,N_9230,N_6145);
xnor U14505 (N_14505,N_9223,N_8825);
or U14506 (N_14506,N_9080,N_5391);
xnor U14507 (N_14507,N_5490,N_6010);
nor U14508 (N_14508,N_8294,N_9024);
nor U14509 (N_14509,N_5917,N_9885);
or U14510 (N_14510,N_7317,N_9859);
or U14511 (N_14511,N_9507,N_5846);
nand U14512 (N_14512,N_6919,N_5833);
or U14513 (N_14513,N_8634,N_5206);
nor U14514 (N_14514,N_7310,N_6229);
and U14515 (N_14515,N_7076,N_8330);
or U14516 (N_14516,N_9476,N_6394);
nand U14517 (N_14517,N_9780,N_5837);
and U14518 (N_14518,N_8065,N_8915);
and U14519 (N_14519,N_6460,N_8781);
or U14520 (N_14520,N_5918,N_5635);
nand U14521 (N_14521,N_8905,N_7197);
xnor U14522 (N_14522,N_9757,N_7357);
xor U14523 (N_14523,N_6993,N_8623);
and U14524 (N_14524,N_7591,N_8103);
or U14525 (N_14525,N_9488,N_5226);
nand U14526 (N_14526,N_9059,N_7187);
nor U14527 (N_14527,N_6111,N_8294);
nand U14528 (N_14528,N_6258,N_6321);
nand U14529 (N_14529,N_6790,N_7872);
nand U14530 (N_14530,N_7875,N_7894);
xor U14531 (N_14531,N_6861,N_6042);
nand U14532 (N_14532,N_5870,N_7634);
xnor U14533 (N_14533,N_6294,N_7365);
nor U14534 (N_14534,N_6066,N_7511);
xor U14535 (N_14535,N_9614,N_5860);
xor U14536 (N_14536,N_8828,N_9378);
nor U14537 (N_14537,N_6644,N_6954);
and U14538 (N_14538,N_5919,N_7190);
nand U14539 (N_14539,N_8798,N_7099);
and U14540 (N_14540,N_6201,N_9620);
and U14541 (N_14541,N_5000,N_5656);
nand U14542 (N_14542,N_6194,N_5834);
xor U14543 (N_14543,N_5344,N_8153);
xnor U14544 (N_14544,N_7494,N_7326);
or U14545 (N_14545,N_5148,N_5183);
or U14546 (N_14546,N_9220,N_8389);
nor U14547 (N_14547,N_9444,N_7222);
nand U14548 (N_14548,N_6195,N_6446);
nor U14549 (N_14549,N_9525,N_8790);
nor U14550 (N_14550,N_5920,N_5409);
and U14551 (N_14551,N_9236,N_9824);
nand U14552 (N_14552,N_8718,N_7881);
and U14553 (N_14553,N_5148,N_7354);
or U14554 (N_14554,N_7112,N_6504);
xnor U14555 (N_14555,N_8938,N_7060);
xor U14556 (N_14556,N_8855,N_8000);
and U14557 (N_14557,N_6565,N_8869);
nand U14558 (N_14558,N_8700,N_5640);
xor U14559 (N_14559,N_7203,N_6057);
and U14560 (N_14560,N_8854,N_7700);
or U14561 (N_14561,N_6382,N_9613);
nor U14562 (N_14562,N_5329,N_6645);
nor U14563 (N_14563,N_5920,N_5289);
and U14564 (N_14564,N_7463,N_7800);
xnor U14565 (N_14565,N_8591,N_6158);
xnor U14566 (N_14566,N_6407,N_7746);
nor U14567 (N_14567,N_5748,N_8506);
nand U14568 (N_14568,N_9047,N_8105);
nand U14569 (N_14569,N_6747,N_5072);
nor U14570 (N_14570,N_8880,N_7847);
nor U14571 (N_14571,N_5091,N_7256);
and U14572 (N_14572,N_9580,N_9392);
nand U14573 (N_14573,N_8350,N_7112);
xor U14574 (N_14574,N_6404,N_8085);
nor U14575 (N_14575,N_9700,N_8753);
xnor U14576 (N_14576,N_6655,N_9604);
nand U14577 (N_14577,N_7351,N_5526);
or U14578 (N_14578,N_8740,N_7851);
xor U14579 (N_14579,N_5654,N_9889);
and U14580 (N_14580,N_7716,N_9794);
xor U14581 (N_14581,N_8800,N_6859);
xnor U14582 (N_14582,N_6788,N_9410);
xnor U14583 (N_14583,N_6270,N_6644);
and U14584 (N_14584,N_7207,N_7352);
nor U14585 (N_14585,N_8326,N_8878);
nand U14586 (N_14586,N_9716,N_5666);
xnor U14587 (N_14587,N_7511,N_9418);
or U14588 (N_14588,N_6364,N_8070);
and U14589 (N_14589,N_9788,N_9647);
or U14590 (N_14590,N_5991,N_5485);
nand U14591 (N_14591,N_6821,N_6431);
nor U14592 (N_14592,N_9968,N_9980);
nor U14593 (N_14593,N_6461,N_9558);
or U14594 (N_14594,N_8102,N_8412);
and U14595 (N_14595,N_5102,N_5131);
nand U14596 (N_14596,N_5810,N_9034);
and U14597 (N_14597,N_8965,N_8939);
and U14598 (N_14598,N_5789,N_5828);
and U14599 (N_14599,N_7776,N_6331);
nor U14600 (N_14600,N_5392,N_5518);
and U14601 (N_14601,N_8495,N_9444);
xnor U14602 (N_14602,N_6515,N_6157);
nand U14603 (N_14603,N_8993,N_8002);
nand U14604 (N_14604,N_9989,N_6510);
and U14605 (N_14605,N_5393,N_5457);
or U14606 (N_14606,N_5079,N_5793);
and U14607 (N_14607,N_9663,N_9070);
xnor U14608 (N_14608,N_7261,N_7490);
nand U14609 (N_14609,N_6680,N_5073);
nor U14610 (N_14610,N_6552,N_8490);
nand U14611 (N_14611,N_8084,N_9564);
xnor U14612 (N_14612,N_8989,N_9310);
and U14613 (N_14613,N_9943,N_5044);
xnor U14614 (N_14614,N_6201,N_8068);
xnor U14615 (N_14615,N_5008,N_6952);
xnor U14616 (N_14616,N_6205,N_9545);
and U14617 (N_14617,N_7123,N_8894);
nand U14618 (N_14618,N_9960,N_9936);
nor U14619 (N_14619,N_6909,N_7088);
xor U14620 (N_14620,N_8796,N_7773);
nand U14621 (N_14621,N_9411,N_7742);
or U14622 (N_14622,N_7432,N_9124);
and U14623 (N_14623,N_8041,N_6232);
nand U14624 (N_14624,N_6197,N_8227);
nor U14625 (N_14625,N_7041,N_7995);
xor U14626 (N_14626,N_6751,N_8349);
xnor U14627 (N_14627,N_6752,N_8859);
nor U14628 (N_14628,N_6343,N_7979);
nor U14629 (N_14629,N_6328,N_5045);
nand U14630 (N_14630,N_8707,N_7891);
nand U14631 (N_14631,N_7477,N_6213);
or U14632 (N_14632,N_5010,N_7102);
xnor U14633 (N_14633,N_5599,N_6064);
or U14634 (N_14634,N_5016,N_5088);
and U14635 (N_14635,N_9394,N_7178);
and U14636 (N_14636,N_7475,N_7598);
nor U14637 (N_14637,N_8591,N_6200);
and U14638 (N_14638,N_5885,N_5803);
or U14639 (N_14639,N_7331,N_6562);
xor U14640 (N_14640,N_7911,N_5314);
and U14641 (N_14641,N_9386,N_5608);
or U14642 (N_14642,N_9864,N_8551);
nand U14643 (N_14643,N_5350,N_8760);
or U14644 (N_14644,N_6787,N_9683);
nor U14645 (N_14645,N_9284,N_7721);
and U14646 (N_14646,N_8940,N_5441);
nand U14647 (N_14647,N_7186,N_7641);
xor U14648 (N_14648,N_9627,N_7842);
and U14649 (N_14649,N_5763,N_6059);
nand U14650 (N_14650,N_8593,N_5006);
or U14651 (N_14651,N_6517,N_7226);
or U14652 (N_14652,N_8434,N_8535);
xor U14653 (N_14653,N_8954,N_8671);
xnor U14654 (N_14654,N_7614,N_8676);
xnor U14655 (N_14655,N_8425,N_9555);
nand U14656 (N_14656,N_9006,N_6420);
and U14657 (N_14657,N_6495,N_7536);
and U14658 (N_14658,N_8505,N_7498);
or U14659 (N_14659,N_9755,N_9256);
and U14660 (N_14660,N_6823,N_6718);
nand U14661 (N_14661,N_8334,N_5736);
and U14662 (N_14662,N_6712,N_7980);
or U14663 (N_14663,N_9780,N_5600);
or U14664 (N_14664,N_7934,N_6220);
and U14665 (N_14665,N_9571,N_5813);
nand U14666 (N_14666,N_6337,N_9551);
xnor U14667 (N_14667,N_5262,N_7511);
nand U14668 (N_14668,N_9083,N_6984);
nor U14669 (N_14669,N_7936,N_6801);
and U14670 (N_14670,N_7448,N_9696);
xnor U14671 (N_14671,N_5233,N_9454);
and U14672 (N_14672,N_8190,N_9650);
nand U14673 (N_14673,N_9938,N_8143);
or U14674 (N_14674,N_8462,N_6604);
and U14675 (N_14675,N_8759,N_5296);
nor U14676 (N_14676,N_6808,N_9300);
nor U14677 (N_14677,N_9395,N_5300);
xnor U14678 (N_14678,N_8472,N_6454);
and U14679 (N_14679,N_9723,N_5163);
nand U14680 (N_14680,N_9752,N_9679);
nor U14681 (N_14681,N_6225,N_7369);
or U14682 (N_14682,N_6042,N_8093);
and U14683 (N_14683,N_5991,N_5325);
xnor U14684 (N_14684,N_5364,N_7123);
or U14685 (N_14685,N_6999,N_9959);
nor U14686 (N_14686,N_5973,N_9435);
or U14687 (N_14687,N_5946,N_5200);
nor U14688 (N_14688,N_7343,N_9404);
nand U14689 (N_14689,N_7598,N_7532);
nand U14690 (N_14690,N_7710,N_7457);
xnor U14691 (N_14691,N_5950,N_7972);
and U14692 (N_14692,N_5561,N_9146);
nand U14693 (N_14693,N_6309,N_7674);
nand U14694 (N_14694,N_7289,N_9676);
nor U14695 (N_14695,N_9413,N_9639);
and U14696 (N_14696,N_8675,N_8834);
nor U14697 (N_14697,N_6400,N_5458);
nor U14698 (N_14698,N_9643,N_6105);
nand U14699 (N_14699,N_5027,N_8288);
nor U14700 (N_14700,N_9319,N_8450);
or U14701 (N_14701,N_6775,N_6121);
xnor U14702 (N_14702,N_7745,N_6118);
nand U14703 (N_14703,N_9202,N_9393);
xor U14704 (N_14704,N_8364,N_5671);
nor U14705 (N_14705,N_7631,N_7043);
nor U14706 (N_14706,N_9978,N_7249);
or U14707 (N_14707,N_7325,N_6720);
nor U14708 (N_14708,N_8940,N_8209);
xor U14709 (N_14709,N_8031,N_7009);
or U14710 (N_14710,N_9545,N_8169);
xnor U14711 (N_14711,N_6481,N_8031);
nor U14712 (N_14712,N_7732,N_6249);
nand U14713 (N_14713,N_6415,N_6224);
xnor U14714 (N_14714,N_8803,N_8676);
nor U14715 (N_14715,N_6995,N_8541);
xor U14716 (N_14716,N_9233,N_8367);
nand U14717 (N_14717,N_5857,N_6072);
nand U14718 (N_14718,N_6422,N_5650);
and U14719 (N_14719,N_5574,N_7862);
and U14720 (N_14720,N_8097,N_8276);
nor U14721 (N_14721,N_5263,N_8241);
and U14722 (N_14722,N_6363,N_8399);
xnor U14723 (N_14723,N_5194,N_9334);
or U14724 (N_14724,N_7428,N_9832);
xnor U14725 (N_14725,N_9803,N_7113);
and U14726 (N_14726,N_6916,N_5193);
and U14727 (N_14727,N_5361,N_5627);
and U14728 (N_14728,N_7059,N_8408);
and U14729 (N_14729,N_7548,N_8690);
xnor U14730 (N_14730,N_7537,N_8786);
xnor U14731 (N_14731,N_9792,N_6629);
nand U14732 (N_14732,N_5392,N_8993);
nor U14733 (N_14733,N_8777,N_8972);
nand U14734 (N_14734,N_5463,N_8415);
or U14735 (N_14735,N_9513,N_6519);
or U14736 (N_14736,N_7179,N_8306);
nand U14737 (N_14737,N_6322,N_7009);
xnor U14738 (N_14738,N_7151,N_5658);
nand U14739 (N_14739,N_8399,N_7569);
nand U14740 (N_14740,N_8020,N_6416);
or U14741 (N_14741,N_6387,N_6085);
nor U14742 (N_14742,N_6209,N_9915);
xor U14743 (N_14743,N_8860,N_7127);
nand U14744 (N_14744,N_7476,N_6912);
xnor U14745 (N_14745,N_9447,N_8853);
xor U14746 (N_14746,N_8545,N_5841);
nor U14747 (N_14747,N_6261,N_7933);
or U14748 (N_14748,N_9422,N_8832);
xnor U14749 (N_14749,N_5142,N_9640);
xnor U14750 (N_14750,N_8154,N_7406);
nand U14751 (N_14751,N_9839,N_8964);
nor U14752 (N_14752,N_7594,N_7555);
and U14753 (N_14753,N_9647,N_8110);
and U14754 (N_14754,N_9375,N_6999);
and U14755 (N_14755,N_5617,N_7183);
nand U14756 (N_14756,N_5388,N_9701);
nand U14757 (N_14757,N_9190,N_8628);
nor U14758 (N_14758,N_8526,N_9367);
or U14759 (N_14759,N_7471,N_8732);
xnor U14760 (N_14760,N_6836,N_6415);
nand U14761 (N_14761,N_7155,N_6097);
or U14762 (N_14762,N_8669,N_8898);
nor U14763 (N_14763,N_6650,N_5573);
or U14764 (N_14764,N_8850,N_5130);
or U14765 (N_14765,N_9666,N_6642);
nor U14766 (N_14766,N_5171,N_7547);
xor U14767 (N_14767,N_6683,N_5473);
nor U14768 (N_14768,N_7854,N_7369);
nand U14769 (N_14769,N_7875,N_7889);
or U14770 (N_14770,N_5938,N_5091);
and U14771 (N_14771,N_5871,N_9055);
nor U14772 (N_14772,N_6986,N_7153);
and U14773 (N_14773,N_6695,N_7748);
nor U14774 (N_14774,N_7933,N_9262);
and U14775 (N_14775,N_6449,N_6187);
or U14776 (N_14776,N_8508,N_9325);
nor U14777 (N_14777,N_9467,N_5371);
nand U14778 (N_14778,N_7183,N_7718);
nand U14779 (N_14779,N_5733,N_8597);
or U14780 (N_14780,N_5722,N_7570);
nor U14781 (N_14781,N_6896,N_9747);
or U14782 (N_14782,N_8786,N_5792);
and U14783 (N_14783,N_9019,N_6213);
nand U14784 (N_14784,N_8947,N_5247);
or U14785 (N_14785,N_7336,N_6162);
xor U14786 (N_14786,N_9493,N_6320);
xnor U14787 (N_14787,N_7465,N_9405);
xor U14788 (N_14788,N_5199,N_7902);
and U14789 (N_14789,N_9807,N_8706);
xnor U14790 (N_14790,N_6158,N_5003);
or U14791 (N_14791,N_5276,N_6114);
nor U14792 (N_14792,N_6995,N_9744);
xor U14793 (N_14793,N_9878,N_9389);
nand U14794 (N_14794,N_7201,N_7056);
or U14795 (N_14795,N_8492,N_8762);
nand U14796 (N_14796,N_6993,N_9577);
nor U14797 (N_14797,N_5563,N_7335);
nor U14798 (N_14798,N_6401,N_6931);
xnor U14799 (N_14799,N_7155,N_8416);
nand U14800 (N_14800,N_9821,N_8436);
xnor U14801 (N_14801,N_6571,N_8481);
or U14802 (N_14802,N_5912,N_5160);
xor U14803 (N_14803,N_6000,N_7497);
nor U14804 (N_14804,N_8617,N_8866);
and U14805 (N_14805,N_5340,N_6187);
and U14806 (N_14806,N_7761,N_8237);
xor U14807 (N_14807,N_9329,N_6230);
or U14808 (N_14808,N_8201,N_6879);
xor U14809 (N_14809,N_6275,N_9919);
or U14810 (N_14810,N_5795,N_9222);
xnor U14811 (N_14811,N_8448,N_6783);
xnor U14812 (N_14812,N_8806,N_8531);
nand U14813 (N_14813,N_7329,N_6238);
and U14814 (N_14814,N_7813,N_7919);
xor U14815 (N_14815,N_9492,N_5580);
nor U14816 (N_14816,N_5166,N_5417);
nor U14817 (N_14817,N_8764,N_8064);
nand U14818 (N_14818,N_5507,N_8342);
nor U14819 (N_14819,N_7125,N_7391);
xor U14820 (N_14820,N_9773,N_6384);
xor U14821 (N_14821,N_7845,N_9505);
nor U14822 (N_14822,N_6291,N_5406);
xnor U14823 (N_14823,N_8670,N_9172);
nor U14824 (N_14824,N_7899,N_6698);
nor U14825 (N_14825,N_9746,N_5332);
nor U14826 (N_14826,N_8953,N_9827);
nand U14827 (N_14827,N_8522,N_9674);
or U14828 (N_14828,N_9348,N_6194);
and U14829 (N_14829,N_8317,N_5533);
or U14830 (N_14830,N_9922,N_5028);
or U14831 (N_14831,N_7938,N_9975);
nand U14832 (N_14832,N_5934,N_8874);
and U14833 (N_14833,N_6084,N_6073);
and U14834 (N_14834,N_7363,N_7600);
xnor U14835 (N_14835,N_8462,N_8671);
or U14836 (N_14836,N_5332,N_8851);
nand U14837 (N_14837,N_9977,N_7190);
xnor U14838 (N_14838,N_7925,N_6263);
or U14839 (N_14839,N_8886,N_7593);
and U14840 (N_14840,N_5392,N_5674);
xor U14841 (N_14841,N_7125,N_5544);
and U14842 (N_14842,N_7550,N_9272);
xor U14843 (N_14843,N_5105,N_5293);
xor U14844 (N_14844,N_8935,N_8509);
and U14845 (N_14845,N_9241,N_5492);
and U14846 (N_14846,N_8985,N_5331);
xnor U14847 (N_14847,N_7757,N_5181);
and U14848 (N_14848,N_9132,N_5639);
xor U14849 (N_14849,N_5832,N_7735);
xnor U14850 (N_14850,N_7960,N_8853);
xnor U14851 (N_14851,N_7890,N_8220);
nor U14852 (N_14852,N_9242,N_7769);
xnor U14853 (N_14853,N_5634,N_6331);
or U14854 (N_14854,N_7214,N_5330);
xor U14855 (N_14855,N_9009,N_8776);
nand U14856 (N_14856,N_6495,N_8262);
xor U14857 (N_14857,N_8621,N_8667);
xor U14858 (N_14858,N_8184,N_6750);
nor U14859 (N_14859,N_9196,N_8399);
or U14860 (N_14860,N_6164,N_9832);
xor U14861 (N_14861,N_6946,N_7349);
and U14862 (N_14862,N_9642,N_8821);
nor U14863 (N_14863,N_5087,N_5261);
xnor U14864 (N_14864,N_9214,N_9145);
and U14865 (N_14865,N_6797,N_8032);
and U14866 (N_14866,N_5645,N_5597);
nand U14867 (N_14867,N_9998,N_7032);
and U14868 (N_14868,N_7093,N_5076);
nand U14869 (N_14869,N_9195,N_7981);
and U14870 (N_14870,N_6978,N_8788);
nor U14871 (N_14871,N_7004,N_8617);
nand U14872 (N_14872,N_6370,N_9381);
and U14873 (N_14873,N_6327,N_8182);
xor U14874 (N_14874,N_5945,N_5918);
and U14875 (N_14875,N_8875,N_6158);
nor U14876 (N_14876,N_9425,N_8501);
xor U14877 (N_14877,N_7604,N_5807);
and U14878 (N_14878,N_5365,N_9032);
and U14879 (N_14879,N_6699,N_6821);
nand U14880 (N_14880,N_9668,N_9526);
nor U14881 (N_14881,N_7827,N_5997);
or U14882 (N_14882,N_5228,N_7260);
or U14883 (N_14883,N_7873,N_9613);
and U14884 (N_14884,N_9590,N_9441);
and U14885 (N_14885,N_5325,N_5887);
nor U14886 (N_14886,N_7890,N_9516);
and U14887 (N_14887,N_7499,N_7475);
nor U14888 (N_14888,N_7087,N_8565);
xnor U14889 (N_14889,N_5849,N_5405);
nand U14890 (N_14890,N_5955,N_5940);
or U14891 (N_14891,N_7936,N_9090);
nand U14892 (N_14892,N_8896,N_9906);
nand U14893 (N_14893,N_8208,N_6465);
nor U14894 (N_14894,N_9810,N_6560);
and U14895 (N_14895,N_7977,N_9349);
nor U14896 (N_14896,N_5989,N_8874);
nor U14897 (N_14897,N_8954,N_7366);
and U14898 (N_14898,N_5734,N_6893);
nor U14899 (N_14899,N_9005,N_8969);
xnor U14900 (N_14900,N_8934,N_6711);
nor U14901 (N_14901,N_9771,N_6268);
nor U14902 (N_14902,N_5747,N_8183);
nand U14903 (N_14903,N_9128,N_5473);
nand U14904 (N_14904,N_5512,N_9961);
or U14905 (N_14905,N_5040,N_6225);
nor U14906 (N_14906,N_6540,N_6322);
nor U14907 (N_14907,N_9877,N_9220);
nor U14908 (N_14908,N_7678,N_6940);
nand U14909 (N_14909,N_6580,N_7378);
nand U14910 (N_14910,N_5781,N_9588);
and U14911 (N_14911,N_9701,N_7078);
or U14912 (N_14912,N_9434,N_7274);
nor U14913 (N_14913,N_8526,N_8768);
nor U14914 (N_14914,N_8090,N_8863);
and U14915 (N_14915,N_7110,N_6041);
xnor U14916 (N_14916,N_9150,N_6034);
or U14917 (N_14917,N_8729,N_9746);
xor U14918 (N_14918,N_8930,N_7221);
nor U14919 (N_14919,N_8047,N_6280);
xor U14920 (N_14920,N_7325,N_5798);
xor U14921 (N_14921,N_9054,N_7239);
and U14922 (N_14922,N_8597,N_5187);
nor U14923 (N_14923,N_6481,N_7160);
and U14924 (N_14924,N_8388,N_8781);
xor U14925 (N_14925,N_5942,N_8989);
and U14926 (N_14926,N_7092,N_8135);
and U14927 (N_14927,N_8457,N_9407);
or U14928 (N_14928,N_5146,N_5702);
or U14929 (N_14929,N_9552,N_9979);
and U14930 (N_14930,N_7934,N_7120);
or U14931 (N_14931,N_6415,N_6079);
nor U14932 (N_14932,N_9188,N_7733);
or U14933 (N_14933,N_6919,N_6132);
or U14934 (N_14934,N_7891,N_8066);
xor U14935 (N_14935,N_7623,N_5949);
and U14936 (N_14936,N_5170,N_5024);
nand U14937 (N_14937,N_6829,N_7857);
and U14938 (N_14938,N_7642,N_5980);
nor U14939 (N_14939,N_7818,N_8483);
and U14940 (N_14940,N_5702,N_6632);
nand U14941 (N_14941,N_7251,N_5160);
or U14942 (N_14942,N_6398,N_6635);
nor U14943 (N_14943,N_7029,N_7197);
and U14944 (N_14944,N_8184,N_5504);
and U14945 (N_14945,N_6226,N_9237);
nand U14946 (N_14946,N_8030,N_5468);
nor U14947 (N_14947,N_7792,N_7481);
nand U14948 (N_14948,N_7570,N_5041);
or U14949 (N_14949,N_7167,N_5244);
nor U14950 (N_14950,N_5305,N_8844);
and U14951 (N_14951,N_7210,N_6265);
nor U14952 (N_14952,N_9251,N_8654);
nor U14953 (N_14953,N_9047,N_7106);
nor U14954 (N_14954,N_5283,N_6766);
xor U14955 (N_14955,N_6016,N_8347);
or U14956 (N_14956,N_9935,N_6995);
xnor U14957 (N_14957,N_9528,N_8431);
nand U14958 (N_14958,N_9866,N_9207);
or U14959 (N_14959,N_5664,N_8659);
or U14960 (N_14960,N_9121,N_8636);
xnor U14961 (N_14961,N_6270,N_5587);
nand U14962 (N_14962,N_5009,N_5615);
and U14963 (N_14963,N_5144,N_9947);
nand U14964 (N_14964,N_6973,N_5266);
nor U14965 (N_14965,N_7636,N_6230);
xnor U14966 (N_14966,N_8639,N_7571);
nor U14967 (N_14967,N_8575,N_6532);
xor U14968 (N_14968,N_8114,N_5333);
nand U14969 (N_14969,N_6314,N_9995);
nand U14970 (N_14970,N_5264,N_6764);
or U14971 (N_14971,N_9357,N_9329);
nor U14972 (N_14972,N_7169,N_6296);
xor U14973 (N_14973,N_5787,N_8380);
and U14974 (N_14974,N_8188,N_5377);
or U14975 (N_14975,N_7213,N_8435);
xor U14976 (N_14976,N_9033,N_6309);
nor U14977 (N_14977,N_8765,N_9465);
xor U14978 (N_14978,N_8985,N_7955);
nand U14979 (N_14979,N_9942,N_5141);
or U14980 (N_14980,N_8475,N_7968);
nand U14981 (N_14981,N_9313,N_9827);
or U14982 (N_14982,N_8509,N_8298);
or U14983 (N_14983,N_6801,N_5341);
nand U14984 (N_14984,N_7525,N_9501);
and U14985 (N_14985,N_9328,N_9479);
or U14986 (N_14986,N_7926,N_5986);
nand U14987 (N_14987,N_5601,N_9446);
xnor U14988 (N_14988,N_7993,N_6435);
xor U14989 (N_14989,N_9156,N_6702);
or U14990 (N_14990,N_8400,N_6320);
or U14991 (N_14991,N_7918,N_9351);
or U14992 (N_14992,N_6384,N_8791);
xnor U14993 (N_14993,N_9262,N_5632);
nand U14994 (N_14994,N_9276,N_8365);
or U14995 (N_14995,N_5917,N_9786);
nor U14996 (N_14996,N_6284,N_7678);
nor U14997 (N_14997,N_6441,N_9342);
xor U14998 (N_14998,N_5908,N_7378);
nand U14999 (N_14999,N_8241,N_7047);
nand U15000 (N_15000,N_12481,N_11169);
or U15001 (N_15001,N_13145,N_14747);
or U15002 (N_15002,N_10886,N_12131);
and U15003 (N_15003,N_11872,N_10059);
xor U15004 (N_15004,N_13686,N_12896);
or U15005 (N_15005,N_13631,N_14623);
nor U15006 (N_15006,N_11348,N_11894);
nand U15007 (N_15007,N_12462,N_11868);
nor U15008 (N_15008,N_10170,N_12151);
nor U15009 (N_15009,N_12730,N_10576);
nor U15010 (N_15010,N_11573,N_14480);
or U15011 (N_15011,N_12004,N_11426);
nor U15012 (N_15012,N_14404,N_14618);
xnor U15013 (N_15013,N_13041,N_12356);
or U15014 (N_15014,N_10063,N_12621);
nor U15015 (N_15015,N_11567,N_10261);
and U15016 (N_15016,N_12519,N_13839);
or U15017 (N_15017,N_12709,N_12225);
and U15018 (N_15018,N_13914,N_11931);
nand U15019 (N_15019,N_11732,N_13454);
nor U15020 (N_15020,N_11743,N_12988);
nor U15021 (N_15021,N_12699,N_10189);
xor U15022 (N_15022,N_12304,N_14109);
or U15023 (N_15023,N_12647,N_13475);
or U15024 (N_15024,N_13922,N_13432);
or U15025 (N_15025,N_12203,N_13322);
nor U15026 (N_15026,N_12696,N_14691);
nand U15027 (N_15027,N_10270,N_14894);
nand U15028 (N_15028,N_11336,N_14484);
xnor U15029 (N_15029,N_12340,N_10856);
or U15030 (N_15030,N_14372,N_10550);
or U15031 (N_15031,N_13455,N_10068);
or U15032 (N_15032,N_12635,N_14227);
or U15033 (N_15033,N_14123,N_14275);
or U15034 (N_15034,N_10748,N_12438);
nand U15035 (N_15035,N_14394,N_14864);
or U15036 (N_15036,N_14931,N_12666);
and U15037 (N_15037,N_12260,N_13078);
xor U15038 (N_15038,N_13327,N_11941);
nor U15039 (N_15039,N_14065,N_11121);
xnor U15040 (N_15040,N_12570,N_13512);
and U15041 (N_15041,N_13062,N_11350);
nor U15042 (N_15042,N_13148,N_11686);
nand U15043 (N_15043,N_10188,N_12817);
and U15044 (N_15044,N_10530,N_13030);
xor U15045 (N_15045,N_14823,N_13532);
xor U15046 (N_15046,N_11819,N_14285);
xor U15047 (N_15047,N_14925,N_12440);
or U15048 (N_15048,N_10971,N_13996);
xor U15049 (N_15049,N_13192,N_10936);
nor U15050 (N_15050,N_10112,N_13840);
and U15051 (N_15051,N_11440,N_13910);
and U15052 (N_15052,N_10796,N_12807);
xnor U15053 (N_15053,N_13693,N_13184);
nand U15054 (N_15054,N_13518,N_13209);
xnor U15055 (N_15055,N_13575,N_11746);
xnor U15056 (N_15056,N_12913,N_10536);
or U15057 (N_15057,N_11463,N_14100);
or U15058 (N_15058,N_13586,N_10148);
and U15059 (N_15059,N_14322,N_10926);
nand U15060 (N_15060,N_12749,N_12590);
xnor U15061 (N_15061,N_13002,N_13894);
nand U15062 (N_15062,N_12275,N_10488);
nor U15063 (N_15063,N_13499,N_14125);
and U15064 (N_15064,N_12932,N_12092);
xor U15065 (N_15065,N_10772,N_14760);
nand U15066 (N_15066,N_13049,N_11824);
xnor U15067 (N_15067,N_11618,N_10101);
xnor U15068 (N_15068,N_10217,N_10386);
nor U15069 (N_15069,N_14153,N_11934);
nor U15070 (N_15070,N_14082,N_11141);
and U15071 (N_15071,N_12412,N_13177);
or U15072 (N_15072,N_12587,N_10093);
nand U15073 (N_15073,N_12136,N_11881);
and U15074 (N_15074,N_14564,N_11901);
xnor U15075 (N_15075,N_12675,N_12154);
nand U15076 (N_15076,N_12318,N_14406);
and U15077 (N_15077,N_11401,N_12194);
or U15078 (N_15078,N_11837,N_13251);
nand U15079 (N_15079,N_12068,N_12366);
or U15080 (N_15080,N_12762,N_14563);
or U15081 (N_15081,N_10017,N_13605);
nor U15082 (N_15082,N_11533,N_10319);
nor U15083 (N_15083,N_12836,N_11299);
nand U15084 (N_15084,N_11635,N_11237);
nand U15085 (N_15085,N_10794,N_10954);
nand U15086 (N_15086,N_14197,N_10046);
and U15087 (N_15087,N_11825,N_11607);
or U15088 (N_15088,N_14403,N_12985);
nand U15089 (N_15089,N_10763,N_14765);
or U15090 (N_15090,N_10080,N_12704);
nor U15091 (N_15091,N_14458,N_11985);
nand U15092 (N_15092,N_11273,N_12120);
nor U15093 (N_15093,N_14391,N_11430);
xor U15094 (N_15094,N_14980,N_14437);
nand U15095 (N_15095,N_10600,N_13590);
nor U15096 (N_15096,N_12155,N_12622);
nor U15097 (N_15097,N_10825,N_12224);
and U15098 (N_15098,N_13502,N_12303);
nand U15099 (N_15099,N_10991,N_12043);
xnor U15100 (N_15100,N_13055,N_10558);
or U15101 (N_15101,N_14344,N_10943);
nand U15102 (N_15102,N_10168,N_10585);
xnor U15103 (N_15103,N_10218,N_14439);
xor U15104 (N_15104,N_13801,N_10555);
or U15105 (N_15105,N_13008,N_11194);
and U15106 (N_15106,N_10262,N_13153);
and U15107 (N_15107,N_14256,N_12718);
xor U15108 (N_15108,N_13827,N_10908);
nand U15109 (N_15109,N_11779,N_10947);
or U15110 (N_15110,N_14470,N_12143);
or U15111 (N_15111,N_10304,N_11096);
and U15112 (N_15112,N_10404,N_13366);
or U15113 (N_15113,N_11524,N_11285);
xnor U15114 (N_15114,N_10892,N_13608);
nand U15115 (N_15115,N_14853,N_13205);
nor U15116 (N_15116,N_11030,N_14221);
nor U15117 (N_15117,N_12823,N_12517);
nor U15118 (N_15118,N_13888,N_14028);
and U15119 (N_15119,N_10638,N_13353);
and U15120 (N_15120,N_11856,N_12008);
or U15121 (N_15121,N_10653,N_11443);
nor U15122 (N_15122,N_11483,N_12424);
nand U15123 (N_15123,N_14543,N_13882);
and U15124 (N_15124,N_11117,N_14089);
xnor U15125 (N_15125,N_13537,N_11980);
or U15126 (N_15126,N_10269,N_14602);
xnor U15127 (N_15127,N_11723,N_11193);
nor U15128 (N_15128,N_10251,N_13622);
nand U15129 (N_15129,N_13162,N_13529);
nand U15130 (N_15130,N_13956,N_10382);
or U15131 (N_15131,N_12905,N_14388);
nand U15132 (N_15132,N_13032,N_11382);
nor U15133 (N_15133,N_10927,N_13426);
and U15134 (N_15134,N_13955,N_11949);
and U15135 (N_15135,N_14421,N_10734);
nand U15136 (N_15136,N_10108,N_11124);
or U15137 (N_15137,N_13929,N_13083);
and U15138 (N_15138,N_10429,N_10138);
and U15139 (N_15139,N_10456,N_10939);
nor U15140 (N_15140,N_11233,N_10816);
xor U15141 (N_15141,N_10077,N_11606);
and U15142 (N_15142,N_11405,N_14369);
xnor U15143 (N_15143,N_14264,N_10853);
nand U15144 (N_15144,N_12518,N_10460);
nor U15145 (N_15145,N_12236,N_11840);
nand U15146 (N_15146,N_11268,N_14802);
xor U15147 (N_15147,N_14238,N_13399);
xor U15148 (N_15148,N_14375,N_14818);
or U15149 (N_15149,N_13878,N_11017);
xnor U15150 (N_15150,N_11238,N_14808);
and U15151 (N_15151,N_13259,N_11183);
xor U15152 (N_15152,N_13460,N_11329);
or U15153 (N_15153,N_11377,N_12885);
nor U15154 (N_15154,N_13923,N_11530);
or U15155 (N_15155,N_11764,N_14918);
and U15156 (N_15156,N_12186,N_10430);
or U15157 (N_15157,N_12018,N_11178);
and U15158 (N_15158,N_10511,N_11695);
xnor U15159 (N_15159,N_14743,N_14057);
nand U15160 (N_15160,N_13732,N_14333);
nand U15161 (N_15161,N_12610,N_11228);
and U15162 (N_15162,N_13893,N_10512);
nor U15163 (N_15163,N_12710,N_11315);
or U15164 (N_15164,N_13129,N_13506);
nand U15165 (N_15165,N_13900,N_11015);
or U15166 (N_15166,N_11650,N_14142);
nor U15167 (N_15167,N_11526,N_10258);
nor U15168 (N_15168,N_13515,N_13510);
nand U15169 (N_15169,N_12083,N_14888);
nand U15170 (N_15170,N_13376,N_12539);
and U15171 (N_15171,N_11522,N_14967);
or U15172 (N_15172,N_13836,N_13051);
nand U15173 (N_15173,N_14280,N_13727);
xor U15174 (N_15174,N_10125,N_13236);
xnor U15175 (N_15175,N_14638,N_11652);
or U15176 (N_15176,N_13067,N_10703);
and U15177 (N_15177,N_11119,N_13403);
and U15178 (N_15178,N_11133,N_10757);
and U15179 (N_15179,N_10373,N_13271);
xnor U15180 (N_15180,N_13130,N_12331);
or U15181 (N_15181,N_12552,N_11602);
nand U15182 (N_15182,N_11062,N_12797);
nor U15183 (N_15183,N_11927,N_10779);
or U15184 (N_15184,N_13748,N_10995);
and U15185 (N_15185,N_10974,N_13109);
nor U15186 (N_15186,N_11967,N_12222);
xor U15187 (N_15187,N_10279,N_11097);
or U15188 (N_15188,N_14577,N_10829);
or U15189 (N_15189,N_13611,N_12554);
and U15190 (N_15190,N_11977,N_12643);
nand U15191 (N_15191,N_14156,N_10697);
nand U15192 (N_15192,N_11333,N_13398);
and U15193 (N_15193,N_14666,N_12367);
nand U15194 (N_15194,N_10551,N_13930);
and U15195 (N_15195,N_12968,N_12943);
nand U15196 (N_15196,N_11751,N_11323);
nor U15197 (N_15197,N_10399,N_14649);
nor U15198 (N_15198,N_14834,N_14660);
and U15199 (N_15199,N_14007,N_13980);
or U15200 (N_15200,N_14521,N_11231);
nand U15201 (N_15201,N_11266,N_10975);
or U15202 (N_15202,N_13991,N_10053);
nand U15203 (N_15203,N_13451,N_13494);
nor U15204 (N_15204,N_13609,N_11472);
xnor U15205 (N_15205,N_11919,N_12159);
nand U15206 (N_15206,N_12256,N_14667);
or U15207 (N_15207,N_12583,N_14207);
and U15208 (N_15208,N_12626,N_12065);
nand U15209 (N_15209,N_11920,N_13793);
nor U15210 (N_15210,N_10377,N_10543);
nand U15211 (N_15211,N_13504,N_11603);
xor U15212 (N_15212,N_10427,N_12689);
and U15213 (N_15213,N_11074,N_13050);
nor U15214 (N_15214,N_13652,N_10675);
nor U15215 (N_15215,N_13382,N_11519);
and U15216 (N_15216,N_14718,N_10154);
or U15217 (N_15217,N_10143,N_13323);
nand U15218 (N_15218,N_13986,N_14682);
xnor U15219 (N_15219,N_12555,N_13188);
or U15220 (N_15220,N_12110,N_14445);
xor U15221 (N_15221,N_14130,N_13260);
nand U15222 (N_15222,N_10976,N_13722);
xnor U15223 (N_15223,N_10281,N_12197);
xnor U15224 (N_15224,N_12939,N_13054);
nand U15225 (N_15225,N_11031,N_13858);
nor U15226 (N_15226,N_11215,N_11554);
or U15227 (N_15227,N_13121,N_14976);
nor U15228 (N_15228,N_10644,N_10855);
nor U15229 (N_15229,N_13562,N_14038);
and U15230 (N_15230,N_11490,N_10238);
or U15231 (N_15231,N_14454,N_12900);
or U15232 (N_15232,N_13577,N_12594);
or U15233 (N_15233,N_11808,N_11277);
and U15234 (N_15234,N_12764,N_10918);
or U15235 (N_15235,N_10626,N_14008);
nand U15236 (N_15236,N_14027,N_14144);
and U15237 (N_15237,N_11768,N_12287);
xor U15238 (N_15238,N_13289,N_13430);
xor U15239 (N_15239,N_13962,N_14632);
nand U15240 (N_15240,N_14268,N_13337);
nand U15241 (N_15241,N_14979,N_14022);
nand U15242 (N_15242,N_13816,N_11820);
nand U15243 (N_15243,N_11135,N_14756);
nand U15244 (N_15244,N_10335,N_14961);
nand U15245 (N_15245,N_12317,N_14392);
xor U15246 (N_15246,N_11675,N_12319);
and U15247 (N_15247,N_12961,N_10972);
nand U15248 (N_15248,N_13081,N_10219);
or U15249 (N_15249,N_13675,N_10841);
nor U15250 (N_15250,N_14946,N_12867);
and U15251 (N_15251,N_13147,N_12179);
or U15252 (N_15252,N_12919,N_12598);
nand U15253 (N_15253,N_14548,N_10647);
and U15254 (N_15254,N_10612,N_13942);
or U15255 (N_15255,N_11341,N_12861);
and U15256 (N_15256,N_10481,N_14077);
nor U15257 (N_15257,N_10556,N_13901);
nand U15258 (N_15258,N_11905,N_12439);
or U15259 (N_15259,N_10860,N_11950);
xor U15260 (N_15260,N_11151,N_13101);
and U15261 (N_15261,N_10061,N_14825);
and U15262 (N_15262,N_10385,N_11833);
xnor U15263 (N_15263,N_11539,N_10273);
or U15264 (N_15264,N_11057,N_12850);
or U15265 (N_15265,N_13719,N_12830);
nand U15266 (N_15266,N_14235,N_12071);
nand U15267 (N_15267,N_13472,N_14408);
nor U15268 (N_15268,N_11548,N_12551);
nand U15269 (N_15269,N_12390,N_11947);
xnor U15270 (N_15270,N_13250,N_13553);
xor U15271 (N_15271,N_13102,N_14801);
nand U15272 (N_15272,N_14746,N_10826);
and U15273 (N_15273,N_14017,N_14821);
xor U15274 (N_15274,N_13733,N_12278);
or U15275 (N_15275,N_11374,N_11309);
nand U15276 (N_15276,N_10824,N_10256);
and U15277 (N_15277,N_11339,N_14095);
xor U15278 (N_15278,N_13479,N_11297);
and U15279 (N_15279,N_12447,N_14185);
and U15280 (N_15280,N_14795,N_10162);
xnor U15281 (N_15281,N_11729,N_12650);
nand U15282 (N_15282,N_13088,N_13099);
xor U15283 (N_15283,N_12529,N_12640);
nand U15284 (N_15284,N_12577,N_13463);
nor U15285 (N_15285,N_14615,N_10076);
nor U15286 (N_15286,N_10328,N_12756);
and U15287 (N_15287,N_13253,N_14570);
xnor U15288 (N_15288,N_11278,N_11796);
nand U15289 (N_15289,N_14219,N_10532);
xnor U15290 (N_15290,N_13673,N_13073);
or U15291 (N_15291,N_11995,N_11452);
xnor U15292 (N_15292,N_11446,N_10761);
or U15293 (N_15293,N_13482,N_11221);
nor U15294 (N_15294,N_13691,N_14674);
and U15295 (N_15295,N_14798,N_14405);
nor U15296 (N_15296,N_11761,N_10894);
nand U15297 (N_15297,N_14587,N_14449);
xor U15298 (N_15298,N_12538,N_14872);
nor U15299 (N_15299,N_10361,N_12210);
nand U15300 (N_15300,N_10419,N_11496);
or U15301 (N_15301,N_11535,N_11457);
or U15302 (N_15302,N_12283,N_10065);
nor U15303 (N_15303,N_11416,N_11044);
nand U15304 (N_15304,N_13191,N_14242);
xnor U15305 (N_15305,N_12674,N_14401);
and U15306 (N_15306,N_12377,N_14266);
and U15307 (N_15307,N_12133,N_11380);
or U15308 (N_15308,N_11632,N_10352);
or U15309 (N_15309,N_13600,N_13343);
and U15310 (N_15310,N_12661,N_12338);
nor U15311 (N_15311,N_13766,N_11190);
nor U15312 (N_15312,N_14133,N_12314);
nand U15313 (N_15313,N_10833,N_12825);
nand U15314 (N_15314,N_12668,N_12171);
and U15315 (N_15315,N_13898,N_14919);
nor U15316 (N_15316,N_12500,N_12550);
nand U15317 (N_15317,N_14316,N_11906);
or U15318 (N_15318,N_14447,N_11818);
nand U15319 (N_15319,N_10791,N_14892);
nor U15320 (N_15320,N_13347,N_13689);
nand U15321 (N_15321,N_11848,N_13118);
nor U15322 (N_15322,N_13334,N_14049);
nand U15323 (N_15323,N_12032,N_12732);
nor U15324 (N_15324,N_13108,N_10048);
xor U15325 (N_15325,N_12717,N_11714);
or U15326 (N_15326,N_12715,N_13265);
and U15327 (N_15327,N_10648,N_13294);
or U15328 (N_15328,N_14576,N_14610);
or U15329 (N_15329,N_11256,N_13017);
xnor U15330 (N_15330,N_12064,N_11997);
xor U15331 (N_15331,N_10531,N_10760);
and U15332 (N_15332,N_11294,N_10846);
nand U15333 (N_15333,N_13074,N_10229);
or U15334 (N_15334,N_12097,N_12014);
xor U15335 (N_15335,N_14415,N_14260);
or U15336 (N_15336,N_13400,N_14522);
nand U15337 (N_15337,N_11023,N_11574);
or U15338 (N_15338,N_13198,N_10934);
or U15339 (N_15339,N_11930,N_14091);
xor U15340 (N_15340,N_12801,N_10810);
and U15341 (N_15341,N_14354,N_11454);
nor U15342 (N_15342,N_13203,N_14476);
xnor U15343 (N_15343,N_12468,N_13902);
nor U15344 (N_15344,N_10347,N_14005);
or U15345 (N_15345,N_13838,N_12486);
nor U15346 (N_15346,N_13539,N_10009);
xor U15347 (N_15347,N_10838,N_14159);
nor U15348 (N_15348,N_11722,N_10898);
xnor U15349 (N_15349,N_12739,N_13522);
nor U15350 (N_15350,N_10233,N_13240);
and U15351 (N_15351,N_12475,N_12084);
nor U15352 (N_15352,N_11338,N_10446);
xor U15353 (N_15353,N_10114,N_13422);
nand U15354 (N_15354,N_13871,N_13579);
and U15355 (N_15355,N_14757,N_11741);
nor U15356 (N_15356,N_10015,N_10467);
xnor U15357 (N_15357,N_14485,N_13033);
nand U15358 (N_15358,N_14414,N_12307);
or U15359 (N_15359,N_10008,N_13607);
or U15360 (N_15360,N_12364,N_13659);
or U15361 (N_15361,N_14448,N_10274);
and U15362 (N_15362,N_14606,N_13200);
and U15363 (N_15363,N_10663,N_10198);
nand U15364 (N_15364,N_14594,N_10267);
and U15365 (N_15365,N_12003,N_12467);
and U15366 (N_15366,N_11161,N_10331);
nand U15367 (N_15367,N_14353,N_11726);
nor U15368 (N_15368,N_13210,N_10739);
or U15369 (N_15369,N_13790,N_12474);
and U15370 (N_15370,N_14317,N_11489);
nor U15371 (N_15371,N_14318,N_11758);
and U15372 (N_15372,N_11798,N_11710);
xnor U15373 (N_15373,N_14766,N_14814);
nor U15374 (N_15374,N_10503,N_13020);
or U15375 (N_15375,N_12156,N_14964);
xor U15376 (N_15376,N_12332,N_11653);
and U15377 (N_15377,N_14870,N_14172);
xnor U15378 (N_15378,N_12604,N_12129);
or U15379 (N_15379,N_14581,N_11287);
xor U15380 (N_15380,N_14993,N_13096);
xnor U15381 (N_15381,N_10524,N_14323);
or U15382 (N_15382,N_14274,N_10620);
xnor U15383 (N_15383,N_14179,N_12477);
nand U15384 (N_15384,N_12524,N_10097);
nand U15385 (N_15385,N_12031,N_11411);
and U15386 (N_15386,N_14584,N_10078);
nor U15387 (N_15387,N_14407,N_14579);
and U15388 (N_15388,N_11793,N_11054);
nor U15389 (N_15389,N_12306,N_11642);
and U15390 (N_15390,N_12062,N_13320);
and U15391 (N_15391,N_10137,N_14004);
or U15392 (N_15392,N_10422,N_14370);
and U15393 (N_15393,N_13638,N_13392);
nor U15394 (N_15394,N_11663,N_10158);
xor U15395 (N_15395,N_10628,N_14416);
nor U15396 (N_15396,N_11407,N_10574);
and U15397 (N_15397,N_13513,N_10606);
nand U15398 (N_15398,N_10177,N_11082);
xor U15399 (N_15399,N_10397,N_13538);
nand U15400 (N_15400,N_14985,N_13027);
and U15401 (N_15401,N_13796,N_11735);
nor U15402 (N_15402,N_14163,N_13138);
and U15403 (N_15403,N_13446,N_14755);
xor U15404 (N_15404,N_12286,N_11232);
and U15405 (N_15405,N_10131,N_12326);
and U15406 (N_15406,N_13080,N_13468);
or U15407 (N_15407,N_13536,N_10002);
nand U15408 (N_15408,N_12342,N_10603);
or U15409 (N_15409,N_10598,N_11485);
nor U15410 (N_15410,N_11175,N_10725);
nand U15411 (N_15411,N_11511,N_14390);
and U15412 (N_15412,N_11687,N_12104);
or U15413 (N_15413,N_11314,N_10693);
or U15414 (N_15414,N_13977,N_11864);
or U15415 (N_15415,N_10755,N_11900);
xor U15416 (N_15416,N_11406,N_10808);
nand U15417 (N_15417,N_11867,N_11831);
or U15418 (N_15418,N_14510,N_13179);
nor U15419 (N_15419,N_14512,N_10340);
and U15420 (N_15420,N_13808,N_13469);
xnor U15421 (N_15421,N_10042,N_13065);
or U15422 (N_15422,N_11955,N_11842);
nand U15423 (N_15423,N_11200,N_11569);
nor U15424 (N_15424,N_14628,N_14356);
nor U15425 (N_15425,N_14547,N_11581);
nor U15426 (N_15426,N_10907,N_12727);
and U15427 (N_15427,N_12309,N_13321);
xor U15428 (N_15428,N_13842,N_12115);
or U15429 (N_15429,N_12346,N_13953);
and U15430 (N_15430,N_12033,N_14002);
xnor U15431 (N_15431,N_13150,N_13618);
nand U15432 (N_15432,N_10767,N_11384);
or U15433 (N_15433,N_14488,N_13954);
and U15434 (N_15434,N_13069,N_14015);
and U15435 (N_15435,N_10250,N_10707);
xor U15436 (N_15436,N_11925,N_11038);
nor U15437 (N_15437,N_11780,N_14456);
xnor U15438 (N_15438,N_12135,N_13272);
and U15439 (N_15439,N_14284,N_12262);
or U15440 (N_15440,N_12733,N_12231);
or U15441 (N_15441,N_11125,N_13262);
and U15442 (N_15442,N_14203,N_14029);
xnor U15443 (N_15443,N_14758,N_14018);
and U15444 (N_15444,N_11849,N_14882);
nand U15445 (N_15445,N_11694,N_13571);
nand U15446 (N_15446,N_12066,N_12549);
nor U15447 (N_15447,N_13592,N_13225);
xnor U15448 (N_15448,N_11594,N_12230);
or U15449 (N_15449,N_14900,N_11671);
and U15450 (N_15450,N_14889,N_13267);
and U15451 (N_15451,N_13375,N_14878);
and U15452 (N_15452,N_10955,N_11372);
xnor U15453 (N_15453,N_10041,N_11830);
and U15454 (N_15454,N_11560,N_10462);
or U15455 (N_15455,N_13349,N_10669);
and U15456 (N_15456,N_11417,N_11468);
nor U15457 (N_15457,N_10582,N_14187);
and U15458 (N_15458,N_14300,N_13443);
nand U15459 (N_15459,N_14010,N_10196);
xnor U15460 (N_15460,N_10876,N_12653);
xnor U15461 (N_15461,N_14949,N_14271);
nor U15462 (N_15462,N_10726,N_14595);
nand U15463 (N_15463,N_11766,N_10450);
xnor U15464 (N_15464,N_13870,N_14565);
xnor U15465 (N_15465,N_12520,N_12929);
or U15466 (N_15466,N_12617,N_12742);
nor U15467 (N_15467,N_11557,N_12272);
nor U15468 (N_15468,N_11381,N_12748);
xnor U15469 (N_15469,N_10227,N_11212);
nand U15470 (N_15470,N_14434,N_11167);
xnor U15471 (N_15471,N_14116,N_12034);
nand U15472 (N_15472,N_11756,N_12002);
or U15473 (N_15473,N_12016,N_11043);
nand U15474 (N_15474,N_14122,N_12284);
or U15475 (N_15475,N_11879,N_10000);
or U15476 (N_15476,N_10812,N_14191);
xor U15477 (N_15477,N_13306,N_11247);
xnor U15478 (N_15478,N_14475,N_10521);
xnor U15479 (N_15479,N_13133,N_14514);
nor U15480 (N_15480,N_14474,N_11750);
or U15481 (N_15481,N_12242,N_12045);
xor U15482 (N_15482,N_11537,N_12313);
xnor U15483 (N_15483,N_11585,N_14640);
nor U15484 (N_15484,N_10743,N_14947);
nor U15485 (N_15485,N_12976,N_10110);
and U15486 (N_15486,N_14903,N_11841);
or U15487 (N_15487,N_12738,N_14984);
nor U15488 (N_15488,N_10470,N_14815);
xnor U15489 (N_15489,N_11397,N_12023);
nand U15490 (N_15490,N_11656,N_11700);
xor U15491 (N_15491,N_14950,N_14062);
nor U15492 (N_15492,N_11303,N_14128);
and U15493 (N_15493,N_14088,N_11752);
nor U15494 (N_15494,N_11922,N_14960);
nand U15495 (N_15495,N_12781,N_11531);
nor U15496 (N_15496,N_12204,N_11226);
nor U15497 (N_15497,N_11220,N_13667);
and U15498 (N_15498,N_11562,N_11435);
or U15499 (N_15499,N_11680,N_10649);
xor U15500 (N_15500,N_10489,N_11568);
or U15501 (N_15501,N_14217,N_14079);
nand U15502 (N_15502,N_11325,N_12582);
and U15503 (N_15503,N_14811,N_14020);
nand U15504 (N_15504,N_11363,N_10771);
or U15505 (N_15505,N_14986,N_12452);
xor U15506 (N_15506,N_12012,N_12089);
or U15507 (N_15507,N_11769,N_10994);
nand U15508 (N_15508,N_10169,N_14591);
or U15509 (N_15509,N_14701,N_14314);
xnor U15510 (N_15510,N_12389,N_12285);
nor U15511 (N_15511,N_12564,N_13190);
nor U15512 (N_15512,N_13572,N_13224);
or U15513 (N_15513,N_12281,N_10847);
and U15514 (N_15514,N_10494,N_14061);
and U15515 (N_15515,N_14246,N_14675);
nor U15516 (N_15516,N_13478,N_11375);
or U15517 (N_15517,N_11629,N_10339);
nand U15518 (N_15518,N_13325,N_12087);
or U15519 (N_15519,N_11102,N_11252);
xnor U15520 (N_15520,N_14923,N_13874);
xnor U15521 (N_15521,N_14930,N_13486);
nor U15522 (N_15522,N_13489,N_13333);
or U15523 (N_15523,N_11727,N_10026);
and U15524 (N_15524,N_12920,N_14835);
nand U15525 (N_15525,N_13247,N_12579);
xor U15526 (N_15526,N_12890,N_11267);
or U15527 (N_15527,N_12942,N_11893);
and U15528 (N_15528,N_12418,N_13844);
nor U15529 (N_15529,N_12614,N_14865);
and U15530 (N_15530,N_11669,N_14759);
xnor U15531 (N_15531,N_10330,N_10627);
xnor U15532 (N_15532,N_10575,N_11302);
or U15533 (N_15533,N_14282,N_13741);
and U15534 (N_15534,N_14359,N_11870);
or U15535 (N_15535,N_13470,N_14231);
xnor U15536 (N_15536,N_10243,N_10664);
xor U15537 (N_15537,N_10679,N_14549);
nor U15538 (N_15538,N_11450,N_12184);
nand U15539 (N_15539,N_13444,N_10129);
and U15540 (N_15540,N_13829,N_14536);
nor U15541 (N_15541,N_10246,N_11862);
or U15542 (N_15542,N_11116,N_10614);
and U15543 (N_15543,N_10091,N_14803);
xor U15544 (N_15544,N_12734,N_10435);
nor U15545 (N_15545,N_14225,N_10730);
nand U15546 (N_15546,N_12435,N_14902);
or U15547 (N_15547,N_10085,N_11551);
nand U15548 (N_15548,N_10837,N_10220);
or U15549 (N_15549,N_10368,N_12324);
or U15550 (N_15550,N_14212,N_10912);
nand U15551 (N_15551,N_13124,N_11274);
or U15552 (N_15552,N_12523,N_10200);
xor U15553 (N_15553,N_12993,N_10356);
and U15554 (N_15554,N_13125,N_11105);
nor U15555 (N_15555,N_12216,N_10875);
nor U15556 (N_15556,N_12954,N_13402);
and U15557 (N_15557,N_10900,N_12721);
or U15558 (N_15558,N_10075,N_11142);
or U15559 (N_15559,N_14196,N_12865);
nand U15560 (N_15560,N_14827,N_10727);
and U15561 (N_15561,N_11861,N_10504);
nand U15562 (N_15562,N_11822,N_13685);
nor U15563 (N_15563,N_11486,N_10226);
and U15564 (N_15564,N_14035,N_14527);
or U15565 (N_15565,N_13654,N_13594);
and U15566 (N_15566,N_12049,N_12443);
xnor U15567 (N_15567,N_12701,N_12472);
or U15568 (N_15568,N_11419,N_14775);
or U15569 (N_15569,N_13794,N_13799);
nor U15570 (N_15570,N_11932,N_12240);
nand U15571 (N_15571,N_14074,N_12684);
nand U15572 (N_15572,N_13943,N_11179);
nand U15573 (N_15573,N_10484,N_12958);
and U15574 (N_15574,N_13798,N_11286);
and U15575 (N_15575,N_12894,N_10514);
xnor U15576 (N_15576,N_10623,N_13531);
or U15577 (N_15577,N_10146,N_12964);
nand U15578 (N_15578,N_11404,N_12678);
or U15579 (N_15579,N_10706,N_14542);
nand U15580 (N_15580,N_10986,N_11001);
nor U15581 (N_15581,N_14349,N_14328);
nand U15582 (N_15582,N_10139,N_14630);
xor U15583 (N_15583,N_13853,N_13617);
nor U15584 (N_15584,N_12703,N_14267);
nand U15585 (N_15585,N_10223,N_11717);
nand U15586 (N_15586,N_12044,N_13624);
nand U15587 (N_15587,N_10264,N_13231);
xor U15588 (N_15588,N_10333,N_14310);
nor U15589 (N_15589,N_14098,N_12347);
nor U15590 (N_15590,N_13413,N_10120);
nor U15591 (N_15591,N_14753,N_12970);
and U15592 (N_15592,N_12456,N_14511);
or U15593 (N_15593,N_14634,N_14646);
nor U15594 (N_15594,N_10283,N_13155);
nand U15595 (N_15595,N_12515,N_12592);
nor U15596 (N_15596,N_13161,N_10405);
and U15597 (N_15597,N_10951,N_14073);
and U15598 (N_15598,N_12843,N_12426);
and U15599 (N_15599,N_14481,N_10498);
and U15600 (N_15600,N_13007,N_10537);
nand U15601 (N_15601,N_14343,N_12530);
or U15602 (N_15602,N_10228,N_11767);
xor U15603 (N_15603,N_14482,N_13960);
and U15604 (N_15604,N_11201,N_13814);
and U15605 (N_15605,N_10332,N_10864);
xor U15606 (N_15606,N_13180,N_14174);
nand U15607 (N_15607,N_12249,N_12127);
nand U15608 (N_15608,N_11492,N_11366);
nor U15609 (N_15609,N_12241,N_11270);
or U15610 (N_15610,N_10028,N_11982);
xor U15611 (N_15611,N_13809,N_10657);
or U15612 (N_15612,N_12196,N_10859);
and U15613 (N_15613,N_12427,N_11155);
and U15614 (N_15614,N_13567,N_13373);
or U15615 (N_15615,N_11612,N_12209);
nor U15616 (N_15616,N_14789,N_11021);
nand U15617 (N_15617,N_14636,N_13079);
or U15618 (N_15618,N_13487,N_14688);
nor U15619 (N_15619,N_11207,N_10630);
xnor U15620 (N_15620,N_12047,N_12464);
nor U15621 (N_15621,N_11140,N_10966);
xnor U15622 (N_15622,N_13290,N_12048);
and U15623 (N_15623,N_10105,N_13812);
and U15624 (N_15624,N_10501,N_12422);
or U15625 (N_15625,N_12864,N_12292);
nor U15626 (N_15626,N_12527,N_11832);
nor U15627 (N_15627,N_10952,N_12258);
and U15628 (N_15628,N_14042,N_13024);
nand U15629 (N_15629,N_12945,N_11209);
nand U15630 (N_15630,N_14357,N_11217);
xnor U15631 (N_15631,N_12026,N_10353);
or U15632 (N_15632,N_14773,N_12971);
xnor U15633 (N_15633,N_10619,N_12987);
and U15634 (N_15634,N_11093,N_10809);
or U15635 (N_15635,N_11022,N_11655);
and U15636 (N_15636,N_13152,N_13746);
and U15637 (N_15637,N_13726,N_12405);
xor U15638 (N_15638,N_14590,N_13134);
or U15639 (N_15639,N_13710,N_10192);
nand U15640 (N_15640,N_10981,N_13551);
or U15641 (N_15641,N_14337,N_14329);
nor U15642 (N_15642,N_11353,N_12305);
xnor U15643 (N_15643,N_13852,N_13019);
and U15644 (N_15644,N_10642,N_12280);
and U15645 (N_15645,N_13744,N_11622);
nand U15646 (N_15646,N_13661,N_10252);
nor U15647 (N_15647,N_12180,N_14164);
and U15648 (N_15648,N_10118,N_11385);
nand U15649 (N_15649,N_14997,N_10054);
nand U15650 (N_15650,N_14693,N_13009);
xnor U15651 (N_15651,N_11123,N_14836);
nor U15652 (N_15652,N_10712,N_14592);
and U15653 (N_15653,N_12728,N_13031);
nor U15654 (N_15654,N_11176,N_11343);
nand U15655 (N_15655,N_13112,N_11515);
xor U15656 (N_15656,N_14657,N_10622);
nor U15657 (N_15657,N_12176,N_11451);
xor U15658 (N_15658,N_12777,N_14578);
xor U15659 (N_15659,N_11578,N_13706);
and U15660 (N_15660,N_12613,N_12561);
and U15661 (N_15661,N_11418,N_10932);
nor U15662 (N_15662,N_11946,N_12608);
and U15663 (N_15663,N_12161,N_11657);
nor U15664 (N_15664,N_13174,N_12323);
and U15665 (N_15665,N_14555,N_10432);
nor U15666 (N_15666,N_13660,N_11698);
xnor U15667 (N_15667,N_11184,N_11254);
or U15668 (N_15668,N_14609,N_13467);
nor U15669 (N_15669,N_11892,N_12198);
and U15670 (N_15670,N_12392,N_11570);
nor U15671 (N_15671,N_12056,N_14146);
or U15672 (N_15672,N_13248,N_14862);
and U15673 (N_15673,N_11591,N_10580);
nor U15674 (N_15674,N_10421,N_14909);
or U15675 (N_15675,N_10617,N_11067);
and U15676 (N_15676,N_10374,N_10586);
nor U15677 (N_15677,N_11944,N_12189);
xnor U15678 (N_15678,N_12015,N_14053);
and U15679 (N_15679,N_13682,N_13119);
nor U15680 (N_15680,N_12455,N_12784);
and U15681 (N_15681,N_10581,N_10821);
or U15682 (N_15682,N_10024,N_12190);
nor U15683 (N_15683,N_11915,N_10445);
xor U15684 (N_15684,N_11845,N_13704);
and U15685 (N_15685,N_11760,N_10144);
xor U15686 (N_15686,N_10535,N_11805);
and U15687 (N_15687,N_13418,N_13298);
xnor U15688 (N_15688,N_12423,N_11505);
xor U15689 (N_15689,N_12290,N_10423);
nand U15690 (N_15690,N_11494,N_14705);
or U15691 (N_15691,N_13815,N_13543);
nand U15692 (N_15692,N_11371,N_11327);
nor U15693 (N_15693,N_10775,N_12891);
nor U15694 (N_15694,N_12459,N_14011);
nor U15695 (N_15695,N_10050,N_14987);
and U15696 (N_15696,N_10245,N_12802);
nor U15697 (N_15697,N_12251,N_14777);
nor U15698 (N_15698,N_14920,N_13784);
and U15699 (N_15699,N_14771,N_11469);
nand U15700 (N_15700,N_12670,N_14438);
nand U15701 (N_15701,N_14901,N_14237);
or U15702 (N_15702,N_14792,N_13018);
xnor U15703 (N_15703,N_11351,N_14026);
nand U15704 (N_15704,N_10996,N_11170);
xnor U15705 (N_15705,N_14715,N_10458);
or U15706 (N_15706,N_11939,N_13662);
and U15707 (N_15707,N_12813,N_13958);
nand U15708 (N_15708,N_11061,N_14184);
nand U15709 (N_15709,N_12719,N_14240);
nand U15710 (N_15710,N_11628,N_13303);
xnor U15711 (N_15711,N_11400,N_10721);
xor U15712 (N_15712,N_10553,N_13056);
and U15713 (N_15713,N_13246,N_12926);
or U15714 (N_15714,N_13959,N_10548);
or U15715 (N_15715,N_13116,N_10471);
nand U15716 (N_15716,N_10074,N_14540);
xor U15717 (N_15717,N_10795,N_14966);
and U15718 (N_15718,N_10662,N_13982);
nand U15719 (N_15719,N_10398,N_12729);
nand U15720 (N_15720,N_10698,N_11050);
and U15721 (N_15721,N_14031,N_14873);
or U15722 (N_15722,N_13383,N_11601);
xor U15723 (N_15723,N_14139,N_12812);
xor U15724 (N_15724,N_11014,N_10444);
nand U15725 (N_15725,N_10079,N_12562);
or U15726 (N_15726,N_10515,N_12687);
xnor U15727 (N_15727,N_12493,N_14379);
nor U15728 (N_15728,N_13318,N_12754);
or U15729 (N_15729,N_14165,N_11085);
and U15730 (N_15730,N_10916,N_11225);
nand U15731 (N_15731,N_11929,N_10187);
or U15732 (N_15732,N_13003,N_11070);
xor U15733 (N_15733,N_13650,N_10538);
nor U15734 (N_15734,N_14269,N_10241);
nand U15735 (N_15735,N_13692,N_13599);
xor U15736 (N_15736,N_11563,N_13779);
xor U15737 (N_15737,N_13672,N_12498);
nand U15738 (N_15738,N_10082,N_10815);
or U15739 (N_15739,N_12753,N_10213);
or U15740 (N_15740,N_10313,N_11589);
nand U15741 (N_15741,N_10830,N_10272);
or U15742 (N_15742,N_11064,N_11245);
or U15743 (N_15743,N_11185,N_14972);
nand U15744 (N_15744,N_11158,N_11797);
nor U15745 (N_15745,N_10762,N_10799);
and U15746 (N_15746,N_13891,N_12148);
nor U15747 (N_15747,N_10865,N_11361);
and U15748 (N_15748,N_14003,N_14664);
xnor U15749 (N_15749,N_10917,N_14096);
nor U15750 (N_15750,N_14374,N_14286);
xnor U15751 (N_15751,N_14999,N_13381);
nor U15752 (N_15752,N_12007,N_11040);
xor U15753 (N_15753,N_13864,N_10284);
nand U15754 (N_15754,N_14620,N_12348);
xnor U15755 (N_15755,N_14876,N_14831);
nand U15756 (N_15756,N_12743,N_14339);
nand U15757 (N_15757,N_10668,N_14559);
nor U15758 (N_15758,N_10206,N_12150);
and U15759 (N_15759,N_10334,N_13021);
xor U15760 (N_15760,N_14898,N_11637);
and U15761 (N_15761,N_14940,N_12766);
or U15762 (N_15762,N_10615,N_10525);
nand U15763 (N_15763,N_13146,N_14796);
or U15764 (N_15764,N_14585,N_10595);
xor U15765 (N_15765,N_13648,N_12106);
xnor U15766 (N_15766,N_13907,N_13819);
nand U15767 (N_15767,N_10426,N_10699);
nand U15768 (N_15768,N_12878,N_13046);
xor U15769 (N_15769,N_14071,N_10004);
xor U15770 (N_15770,N_13544,N_10178);
nand U15771 (N_15771,N_13831,N_14365);
xnor U15772 (N_15772,N_13584,N_11392);
or U15773 (N_15773,N_13677,N_14430);
nor U15774 (N_15774,N_12659,N_12744);
nand U15775 (N_15775,N_11999,N_13534);
nand U15776 (N_15776,N_12255,N_10171);
nor U15777 (N_15777,N_10889,N_11661);
or U15778 (N_15778,N_12433,N_12826);
nor U15779 (N_15779,N_11005,N_10210);
xnor U15780 (N_15780,N_14000,N_13103);
or U15781 (N_15781,N_11084,N_12384);
nand U15782 (N_15782,N_13904,N_10944);
nor U15783 (N_15783,N_13300,N_12265);
or U15784 (N_15784,N_13496,N_12525);
or U15785 (N_15785,N_11659,N_14912);
xnor U15786 (N_15786,N_13068,N_10977);
nor U15787 (N_15787,N_11358,N_13876);
and U15788 (N_15788,N_11282,N_14847);
or U15789 (N_15789,N_14571,N_12824);
or U15790 (N_15790,N_14102,N_10720);
or U15791 (N_15791,N_13761,N_11550);
and U15792 (N_15792,N_10247,N_11623);
and U15793 (N_15793,N_13564,N_12027);
xnor U15794 (N_15794,N_10802,N_14926);
nor U15795 (N_15795,N_11971,N_14953);
nand U15796 (N_15796,N_10298,N_12660);
nor U15797 (N_15797,N_13787,N_11280);
or U15798 (N_15798,N_13243,N_10651);
nand U15799 (N_15799,N_12722,N_14820);
or U15800 (N_15800,N_14725,N_10672);
xnor U15801 (N_15801,N_14917,N_10940);
nand U15802 (N_15802,N_13754,N_11143);
and U15803 (N_15803,N_12591,N_14099);
or U15804 (N_15804,N_12328,N_12979);
or U15805 (N_15805,N_10811,N_14210);
nor U15806 (N_15806,N_11923,N_12202);
and U15807 (N_15807,N_12485,N_10978);
xor U15808 (N_15808,N_12805,N_14023);
nand U15809 (N_15809,N_11039,N_11099);
nor U15810 (N_15810,N_12693,N_13285);
xor U15811 (N_15811,N_10866,N_12706);
xnor U15812 (N_15812,N_11855,N_11790);
xnor U15813 (N_15813,N_11283,N_12499);
or U15814 (N_15814,N_13040,N_10364);
xnor U15815 (N_15815,N_12030,N_11298);
nor U15816 (N_15816,N_12680,N_12682);
or U15817 (N_15817,N_12917,N_13311);
nand U15818 (N_15818,N_14243,N_10392);
or U15819 (N_15819,N_14507,N_14719);
or U15820 (N_15820,N_13237,N_13409);
or U15821 (N_15821,N_13932,N_14340);
nand U15822 (N_15822,N_12211,N_13437);
or U15823 (N_15823,N_11360,N_13593);
xor U15824 (N_15824,N_11234,N_11787);
nand U15825 (N_15825,N_11275,N_12775);
xnor U15826 (N_15826,N_11402,N_13233);
xnor U15827 (N_15827,N_12245,N_13684);
or U15828 (N_15828,N_12615,N_11834);
or U15829 (N_15829,N_11250,N_12657);
and U15830 (N_15830,N_12076,N_11035);
and U15831 (N_15831,N_13666,N_10505);
nand U15832 (N_15832,N_13731,N_14687);
and U15833 (N_15833,N_11307,N_14346);
nor U15834 (N_15834,N_14707,N_13547);
or U15835 (N_15835,N_13332,N_14752);
xnor U15836 (N_15836,N_13734,N_12491);
nand U15837 (N_15837,N_11978,N_13695);
nor U15838 (N_15838,N_12247,N_13764);
nand U15839 (N_15839,N_10151,N_12227);
or U15840 (N_15840,N_12024,N_12851);
or U15841 (N_15841,N_12293,N_10349);
nand U15842 (N_15842,N_13107,N_12747);
nand U15843 (N_15843,N_11313,N_12910);
nor U15844 (N_15844,N_12182,N_11609);
xor U15845 (N_15845,N_14689,N_14436);
and U15846 (N_15846,N_11777,N_10142);
xor U15847 (N_15847,N_10756,N_10872);
or U15848 (N_15848,N_10321,N_10384);
nand U15849 (N_15849,N_11149,N_13221);
nand U15850 (N_15850,N_10278,N_13011);
nand U15851 (N_15851,N_12847,N_12337);
nor U15852 (N_15852,N_13196,N_10345);
xnor U15853 (N_15853,N_13714,N_10714);
and U15854 (N_15854,N_14068,N_10018);
nor U15855 (N_15855,N_13811,N_11658);
xnor U15856 (N_15856,N_10596,N_13576);
nand U15857 (N_15857,N_10854,N_12859);
nor U15858 (N_15858,N_13063,N_10140);
nor U15859 (N_15859,N_11685,N_13760);
nor U15860 (N_15860,N_13058,N_13277);
nand U15861 (N_15861,N_12877,N_12778);
nor U15862 (N_15862,N_14016,N_11134);
and U15863 (N_15863,N_10359,N_11664);
or U15864 (N_15864,N_14697,N_12420);
nand U15865 (N_15865,N_10546,N_14528);
xor U15866 (N_15866,N_11651,N_11261);
and U15867 (N_15867,N_10350,N_12941);
or U15868 (N_15868,N_11989,N_11028);
or U15869 (N_15869,N_11156,N_10088);
and U15870 (N_15870,N_13554,N_11078);
or U15871 (N_15871,N_11188,N_12982);
or U15872 (N_15872,N_12897,N_13223);
and U15873 (N_15873,N_14951,N_12178);
xnor U15874 (N_15874,N_12821,N_12114);
or U15875 (N_15875,N_12698,N_12157);
and U15876 (N_15876,N_10235,N_13360);
or U15877 (N_15877,N_10563,N_11478);
nor U15878 (N_15878,N_12214,N_10509);
nor U15879 (N_15879,N_13075,N_12914);
nand U15880 (N_15880,N_14148,N_11495);
nand U15881 (N_15881,N_11553,N_14325);
nand U15882 (N_15882,N_10051,N_12090);
or U15883 (N_15883,N_12755,N_11080);
and U15884 (N_15884,N_13535,N_13424);
nand U15885 (N_15885,N_14658,N_10415);
and U15886 (N_15886,N_12301,N_13640);
nor U15887 (N_15887,N_10237,N_14819);
and U15888 (N_15888,N_13495,N_13948);
nor U15889 (N_15889,N_10095,N_11319);
or U15890 (N_15890,N_13847,N_11890);
xor U15891 (N_15891,N_13092,N_14289);
and U15892 (N_15892,N_14168,N_14092);
nor U15893 (N_15893,N_14945,N_11996);
nor U15894 (N_15894,N_11445,N_13340);
xnor U15895 (N_15895,N_13728,N_10181);
nor U15896 (N_15896,N_13197,N_13514);
and U15897 (N_15897,N_10276,N_12185);
nor U15898 (N_15898,N_13757,N_12619);
nand U15899 (N_15899,N_14296,N_13806);
nor U15900 (N_15900,N_13701,N_11009);
nor U15901 (N_15901,N_14738,N_13768);
nor U15902 (N_15902,N_12354,N_13189);
nand U15903 (N_15903,N_14469,N_11503);
or U15904 (N_15904,N_11229,N_14684);
and U15905 (N_15905,N_14412,N_13044);
nand U15906 (N_15906,N_14839,N_10719);
xor U15907 (N_15907,N_10858,N_11497);
or U15908 (N_15908,N_10443,N_13885);
and U15909 (N_15909,N_11059,N_13182);
and U15910 (N_15910,N_11875,N_13708);
xor U15911 (N_15911,N_14575,N_12665);
nand U15912 (N_15912,N_13057,N_14132);
and U15913 (N_15913,N_10067,N_10800);
or U15914 (N_15914,N_14711,N_10312);
or U15915 (N_15915,N_12870,N_13476);
nor U15916 (N_15916,N_11424,N_14201);
xnor U15917 (N_15917,N_12261,N_13288);
and U15918 (N_15918,N_13933,N_13345);
xor U15919 (N_15919,N_12339,N_11011);
or U15920 (N_15920,N_13560,N_13877);
xnor U15921 (N_15921,N_11481,N_10774);
nor U15922 (N_15922,N_12974,N_12909);
xnor U15923 (N_15923,N_14147,N_13548);
xor U15924 (N_15924,N_12250,N_11045);
and U15925 (N_15925,N_12899,N_10677);
or U15926 (N_15926,N_11817,N_14036);
nor U15927 (N_15927,N_13085,N_13045);
xnor U15928 (N_15928,N_12404,N_10570);
nand U15929 (N_15929,N_13585,N_11003);
and U15930 (N_15930,N_10487,N_11019);
nor U15931 (N_15931,N_14994,N_12683);
nor U15932 (N_15932,N_11579,N_10790);
or U15933 (N_15933,N_11036,N_10096);
nand U15934 (N_15934,N_14729,N_14973);
xnor U15935 (N_15935,N_12289,N_12081);
and U15936 (N_15936,N_12951,N_10199);
nand U15937 (N_15937,N_13305,N_11561);
nand U15938 (N_15938,N_14714,N_11556);
xnor U15939 (N_15939,N_10099,N_10737);
or U15940 (N_15940,N_11471,N_13707);
or U15941 (N_15941,N_12395,N_13428);
and U15942 (N_15942,N_13774,N_10817);
nor U15943 (N_15943,N_12414,N_13702);
or U15944 (N_15944,N_12029,N_14586);
or U15945 (N_15945,N_10770,N_10897);
nor U15946 (N_15946,N_11182,N_12580);
xnor U15947 (N_15947,N_13445,N_11731);
and U15948 (N_15948,N_14978,N_14492);
nor U15949 (N_15949,N_10654,N_14234);
or U15950 (N_15950,N_13545,N_10604);
nor U15951 (N_15951,N_14690,N_11498);
nor U15952 (N_15952,N_13047,N_14150);
nor U15953 (N_15953,N_14617,N_14041);
xnor U15954 (N_15954,N_10362,N_14182);
nor U15955 (N_15955,N_11118,N_14642);
xor U15956 (N_15956,N_12644,N_10136);
xnor U15957 (N_15957,N_12862,N_10751);
or U15958 (N_15958,N_11024,N_13082);
nand U15959 (N_15959,N_12898,N_11342);
nor U15960 (N_15960,N_12565,N_10960);
nor U15961 (N_15961,N_10113,N_11504);
and U15962 (N_15962,N_13988,N_14992);
nand U15963 (N_15963,N_11770,N_13690);
or U15964 (N_15964,N_12611,N_13416);
and U15965 (N_15965,N_13817,N_10937);
nand U15966 (N_15966,N_14251,N_14744);
xor U15967 (N_15967,N_12124,N_10631);
xnor U15968 (N_15968,N_13143,N_11438);
nor U15969 (N_15969,N_10735,N_13252);
xnor U15970 (N_15970,N_12263,N_11049);
nor U15971 (N_15971,N_12607,N_10881);
or U15972 (N_15972,N_13903,N_10588);
xor U15973 (N_15973,N_11728,N_11244);
xor U15974 (N_15974,N_11747,N_10436);
and U15975 (N_15975,N_12141,N_12257);
nor U15976 (N_15976,N_12999,N_12288);
xnor U15977 (N_15977,N_12073,N_11516);
nor U15978 (N_15978,N_14491,N_10066);
nand U15979 (N_15979,N_10539,N_12799);
xnor U15980 (N_15980,N_12956,N_10840);
xor U15981 (N_15981,N_12244,N_10957);
or U15982 (N_15982,N_11086,N_13384);
xnor U15983 (N_15983,N_12938,N_14970);
xnor U15984 (N_15984,N_12046,N_13015);
nand U15985 (N_15985,N_14216,N_12557);
xnor U15986 (N_15986,N_13014,N_12079);
xor U15987 (N_15987,N_13245,N_14669);
or U15988 (N_15988,N_13879,N_13395);
nand U15989 (N_15989,N_10839,N_10564);
nor U15990 (N_15990,N_14728,N_14508);
nor U15991 (N_15991,N_11850,N_12600);
or U15992 (N_15992,N_10873,N_13404);
and U15993 (N_15993,N_12569,N_14199);
nand U15994 (N_15994,N_11720,N_12145);
nor U15995 (N_15995,N_13169,N_12432);
xor U15996 (N_15996,N_12536,N_12957);
nor U15997 (N_15997,N_13527,N_11224);
or U15998 (N_15998,N_11888,N_11166);
nor U15999 (N_15999,N_13397,N_14250);
nand U16000 (N_16000,N_14934,N_11972);
or U16001 (N_16001,N_10909,N_13971);
nand U16002 (N_16002,N_12568,N_12193);
or U16003 (N_16003,N_11795,N_12429);
xnor U16004 (N_16004,N_12918,N_14726);
and U16005 (N_16005,N_12981,N_10948);
and U16006 (N_16006,N_11399,N_10686);
and U16007 (N_16007,N_13713,N_11781);
nor U16008 (N_16008,N_12845,N_14513);
and U16009 (N_16009,N_13336,N_13581);
nor U16010 (N_16010,N_14420,N_12880);
nand U16011 (N_16011,N_13072,N_14424);
and U16012 (N_16012,N_11555,N_11320);
nand U16013 (N_16013,N_11583,N_10337);
nor U16014 (N_16014,N_13843,N_13884);
nand U16015 (N_16015,N_13461,N_11055);
or U16016 (N_16016,N_11281,N_13620);
xor U16017 (N_16017,N_11668,N_14741);
nand U16018 (N_16018,N_10924,N_14258);
nand U16019 (N_16019,N_13012,N_11487);
or U16020 (N_16020,N_12393,N_10522);
nor U16021 (N_16021,N_11239,N_12535);
and U16022 (N_16022,N_11634,N_14806);
nand U16023 (N_16023,N_14680,N_11911);
nor U16024 (N_16024,N_12378,N_12077);
nand U16025 (N_16025,N_12990,N_14423);
and U16026 (N_16026,N_11346,N_14192);
nor U16027 (N_16027,N_12741,N_11532);
nor U16028 (N_16028,N_12531,N_14770);
and U16029 (N_16029,N_10542,N_14186);
nand U16030 (N_16030,N_12229,N_11165);
or U16031 (N_16031,N_11763,N_10244);
or U16032 (N_16032,N_13039,N_12428);
or U16033 (N_16033,N_10925,N_11258);
or U16034 (N_16034,N_10010,N_12827);
nor U16035 (N_16035,N_10915,N_12248);
nand U16036 (N_16036,N_14358,N_11037);
or U16037 (N_16037,N_12059,N_10807);
or U16038 (N_16038,N_14568,N_10670);
nand U16039 (N_16039,N_11230,N_11521);
xnor U16040 (N_16040,N_10591,N_10014);
nand U16041 (N_16041,N_13115,N_10234);
nand U16042 (N_16042,N_10056,N_12138);
nor U16043 (N_16043,N_13833,N_13845);
nand U16044 (N_16044,N_14928,N_10369);
nor U16045 (N_16045,N_10587,N_10107);
xnor U16046 (N_16046,N_13623,N_11783);
nand U16047 (N_16047,N_11500,N_13453);
nand U16048 (N_16048,N_11676,N_10084);
or U16049 (N_16049,N_13094,N_11640);
or U16050 (N_16050,N_10263,N_14441);
xor U16051 (N_16051,N_12654,N_12372);
xor U16052 (N_16052,N_14538,N_11882);
xor U16053 (N_16053,N_11110,N_10987);
nand U16054 (N_16054,N_13765,N_12630);
nand U16055 (N_16055,N_12983,N_13788);
and U16056 (N_16056,N_10910,N_11580);
xnor U16057 (N_16057,N_10681,N_13837);
or U16058 (N_16058,N_11321,N_13193);
xor U16059 (N_16059,N_13244,N_12835);
or U16060 (N_16060,N_11639,N_14277);
and U16061 (N_16061,N_10888,N_12996);
or U16062 (N_16062,N_14024,N_10589);
nand U16063 (N_16063,N_12977,N_13915);
nor U16064 (N_16064,N_11127,N_11679);
or U16065 (N_16065,N_13328,N_14259);
xnor U16066 (N_16066,N_11682,N_12625);
xor U16067 (N_16067,N_12967,N_12773);
nor U16068 (N_16068,N_11386,N_14708);
nor U16069 (N_16069,N_13556,N_12490);
or U16070 (N_16070,N_12341,N_14954);
nand U16071 (N_16071,N_11466,N_14428);
or U16072 (N_16072,N_11092,N_10973);
and U16073 (N_16073,N_13367,N_10621);
xor U16074 (N_16074,N_10259,N_12219);
nor U16075 (N_16075,N_10451,N_12872);
nand U16076 (N_16076,N_10029,N_13715);
xor U16077 (N_16077,N_14681,N_12816);
nand U16078 (N_16078,N_12998,N_11444);
nor U16079 (N_16079,N_13220,N_12403);
and U16080 (N_16080,N_10249,N_12596);
or U16081 (N_16081,N_13052,N_11810);
nand U16082 (N_16082,N_10528,N_10111);
nor U16083 (N_16083,N_12759,N_12911);
nand U16084 (N_16084,N_12585,N_13818);
nor U16085 (N_16085,N_14856,N_13105);
nand U16086 (N_16086,N_14398,N_12279);
nor U16087 (N_16087,N_13694,N_13232);
or U16088 (N_16088,N_14616,N_12828);
or U16089 (N_16089,N_12380,N_12768);
nor U16090 (N_16090,N_10899,N_14464);
xnor U16091 (N_16091,N_13994,N_12779);
nor U16092 (N_16092,N_13172,N_10424);
nand U16093 (N_16093,N_12669,N_14442);
nand U16094 (N_16094,N_14890,N_14907);
and U16095 (N_16095,N_13606,N_10135);
xnor U16096 (N_16096,N_10773,N_13477);
or U16097 (N_16097,N_11534,N_13979);
nand U16098 (N_16098,N_11060,N_11540);
xnor U16099 (N_16099,N_13128,N_13950);
or U16100 (N_16100,N_12702,N_10485);
nand U16101 (N_16101,N_12163,N_13449);
or U16102 (N_16102,N_13280,N_14332);
and U16103 (N_16103,N_11518,N_10605);
nor U16104 (N_16104,N_10440,N_10317);
nor U16105 (N_16105,N_10723,N_11173);
xor U16106 (N_16106,N_10718,N_13171);
xor U16107 (N_16107,N_11689,N_10741);
nand U16108 (N_16108,N_14593,N_12705);
nand U16109 (N_16109,N_12478,N_11058);
xor U16110 (N_16110,N_13241,N_14063);
and U16111 (N_16111,N_11235,N_11368);
nor U16112 (N_16112,N_13456,N_11271);
nor U16113 (N_16113,N_10045,N_14083);
nand U16114 (N_16114,N_12421,N_14750);
and U16115 (N_16115,N_12200,N_11641);
or U16116 (N_16116,N_10381,N_13655);
nand U16117 (N_16117,N_10395,N_14355);
and U16118 (N_16118,N_10956,N_12629);
and U16119 (N_16119,N_13773,N_13753);
nand U16120 (N_16120,N_10310,N_13723);
nand U16121 (N_16121,N_13683,N_11943);
xnor U16122 (N_16122,N_12752,N_11396);
nand U16123 (N_16123,N_11572,N_13258);
nand U16124 (N_16124,N_13354,N_12441);
nand U16125 (N_16125,N_14506,N_10689);
xnor U16126 (N_16126,N_13286,N_13957);
xnor U16127 (N_16127,N_10982,N_14678);
nand U16128 (N_16128,N_13917,N_12992);
or U16129 (N_16129,N_10877,N_10464);
nor U16130 (N_16130,N_10660,N_14435);
xor U16131 (N_16131,N_12856,N_12672);
xnor U16132 (N_16132,N_11132,N_13362);
nor U16133 (N_16133,N_13926,N_10793);
nand U16134 (N_16134,N_13473,N_11126);
nor U16135 (N_16135,N_12761,N_11662);
and U16136 (N_16136,N_10207,N_14969);
or U16137 (N_16137,N_12501,N_11393);
nor U16138 (N_16138,N_13410,N_14494);
xor U16139 (N_16139,N_12888,N_14965);
and U16140 (N_16140,N_14341,N_14671);
and U16141 (N_16141,N_13846,N_14209);
nor U16142 (N_16142,N_13541,N_12457);
nand U16143 (N_16143,N_12330,N_10593);
nor U16144 (N_16144,N_11887,N_14143);
or U16145 (N_16145,N_10022,N_13279);
and U16146 (N_16146,N_13679,N_12792);
nand U16147 (N_16147,N_11421,N_10758);
xor U16148 (N_16148,N_14526,N_12349);
or U16149 (N_16149,N_14627,N_12360);
nor U16150 (N_16150,N_14922,N_10294);
or U16151 (N_16151,N_10804,N_14605);
or U16152 (N_16152,N_13737,N_13070);
and U16153 (N_16153,N_12351,N_10938);
xnor U16154 (N_16154,N_13832,N_10040);
or U16155 (N_16155,N_12177,N_13010);
and U16156 (N_16156,N_11227,N_12886);
or U16157 (N_16157,N_14272,N_14550);
and U16158 (N_16158,N_11816,N_14232);
and U16159 (N_16159,N_10584,N_11988);
nand U16160 (N_16160,N_10633,N_14600);
nand U16161 (N_16161,N_12848,N_14731);
and U16162 (N_16162,N_12912,N_14175);
and U16163 (N_16163,N_12274,N_14154);
nand U16164 (N_16164,N_10645,N_12463);
and U16165 (N_16165,N_13293,N_10275);
and U16166 (N_16166,N_13697,N_13729);
nor U16167 (N_16167,N_11264,N_14537);
nor U16168 (N_16168,N_10820,N_14763);
nand U16169 (N_16169,N_14304,N_14409);
nand U16170 (N_16170,N_10523,N_13167);
nand U16171 (N_16171,N_14603,N_11046);
nand U16172 (N_16172,N_10357,N_13735);
nor U16173 (N_16173,N_10650,N_12373);
xor U16174 (N_16174,N_14252,N_13316);
nor U16175 (N_16175,N_14293,N_10299);
xnor U16176 (N_16176,N_11168,N_12963);
nand U16177 (N_16177,N_14446,N_11692);
or U16178 (N_16178,N_12875,N_13736);
or U16179 (N_16179,N_14351,N_12218);
nor U16180 (N_16180,N_10629,N_14695);
xnor U16181 (N_16181,N_13598,N_10508);
or U16182 (N_16182,N_12842,N_14377);
nor U16183 (N_16183,N_11617,N_12335);
xnor U16184 (N_16184,N_11428,N_13093);
and U16185 (N_16185,N_11312,N_10145);
nor U16186 (N_16186,N_11737,N_13588);
nor U16187 (N_16187,N_12259,N_10923);
or U16188 (N_16188,N_10150,N_13139);
nor U16189 (N_16189,N_11597,N_11536);
nor U16190 (N_16190,N_12208,N_13570);
and U16191 (N_16191,N_10476,N_14804);
nand U16192 (N_16192,N_11690,N_11715);
or U16193 (N_16193,N_12700,N_12677);
nand U16194 (N_16194,N_13151,N_14495);
or U16195 (N_16195,N_11821,N_14694);
nor U16196 (N_16196,N_14709,N_12400);
or U16197 (N_16197,N_14866,N_14648);
and U16198 (N_16198,N_11335,N_11016);
nor U16199 (N_16199,N_12849,N_12726);
or U16200 (N_16200,N_14281,N_11839);
xnor U16201 (N_16201,N_12628,N_13149);
nor U16202 (N_16202,N_10842,N_14461);
nand U16203 (N_16203,N_14717,N_14855);
xnor U16204 (N_16204,N_13628,N_12160);
nor U16205 (N_16205,N_11605,N_14780);
nor U16206 (N_16206,N_13035,N_14211);
nand U16207 (N_16207,N_11205,N_13195);
nor U16208 (N_16208,N_10277,N_10867);
xnor U16209 (N_16209,N_12040,N_12072);
xor U16210 (N_16210,N_14320,N_12858);
and U16211 (N_16211,N_12375,N_14845);
nand U16212 (N_16212,N_13457,N_10126);
nand U16213 (N_16213,N_13973,N_10341);
and U16214 (N_16214,N_12540,N_12102);
xnor U16215 (N_16215,N_10782,N_11586);
nand U16216 (N_16216,N_11002,N_14330);
nor U16217 (N_16217,N_11528,N_14013);
or U16218 (N_16218,N_11131,N_12889);
nor U16219 (N_16219,N_13270,N_13117);
and U16220 (N_16220,N_12408,N_12296);
nor U16221 (N_16221,N_14032,N_10288);
nor U16222 (N_16222,N_10577,N_11912);
and U16223 (N_16223,N_10323,N_10625);
or U16224 (N_16224,N_14070,N_12973);
nand U16225 (N_16225,N_11677,N_13759);
xnor U16226 (N_16226,N_13869,N_12690);
and U16227 (N_16227,N_14054,N_11362);
nor U16228 (N_16228,N_11742,N_12321);
nand U16229 (N_16229,N_11415,N_12228);
xnor U16230 (N_16230,N_11042,N_11969);
and U16231 (N_16231,N_10968,N_14641);
and U16232 (N_16232,N_13022,N_12419);
and U16233 (N_16233,N_14704,N_11317);
xnor U16234 (N_16234,N_13613,N_10222);
nor U16235 (N_16235,N_13669,N_10529);
and U16236 (N_16236,N_10740,N_12268);
nand U16237 (N_16237,N_11871,N_13781);
or U16238 (N_16238,N_14817,N_11455);
or U16239 (N_16239,N_12140,N_13084);
and U16240 (N_16240,N_11048,N_14121);
xor U16241 (N_16241,N_10032,N_10901);
and U16242 (N_16242,N_12382,N_12355);
nand U16243 (N_16243,N_13299,N_12852);
or U16244 (N_16244,N_12903,N_14220);
nor U16245 (N_16245,N_11300,N_14515);
xnor U16246 (N_16246,N_12532,N_14413);
nand U16247 (N_16247,N_14473,N_11759);
and U16248 (N_16248,N_14262,N_10367);
nor U16249 (N_16249,N_11153,N_11804);
or U16250 (N_16250,N_11541,N_11387);
xnor U16251 (N_16251,N_13274,N_10240);
and U16252 (N_16252,N_12789,N_14769);
nor U16253 (N_16253,N_10702,N_12758);
or U16254 (N_16254,N_12425,N_13627);
nor U16255 (N_16255,N_14683,N_13725);
nor U16256 (N_16256,N_12793,N_14670);
or U16257 (N_16257,N_14534,N_14913);
or U16258 (N_16258,N_13924,N_12469);
nand U16259 (N_16259,N_12774,N_11613);
nand U16260 (N_16260,N_12188,N_10025);
and U16261 (N_16261,N_12483,N_10179);
xnor U16262 (N_16262,N_13578,N_11414);
nand U16263 (N_16263,N_11926,N_13356);
nor U16264 (N_16264,N_13187,N_12740);
xor U16265 (N_16265,N_14263,N_13987);
and U16266 (N_16266,N_10465,N_14935);
xor U16267 (N_16267,N_12572,N_13688);
xor U16268 (N_16268,N_10358,N_13219);
or U16269 (N_16269,N_12969,N_13342);
nor U16270 (N_16270,N_11649,N_14843);
and U16271 (N_16271,N_14223,N_12098);
and U16272 (N_16272,N_10665,N_14740);
nor U16273 (N_16273,N_12095,N_10437);
and U16274 (N_16274,N_14051,N_10742);
or U16275 (N_16275,N_14893,N_11966);
or U16276 (N_16276,N_13176,N_14410);
xnor U16277 (N_16277,N_11025,N_14597);
nor U16278 (N_16278,N_14001,N_13023);
and U16279 (N_16279,N_11704,N_14288);
nand U16280 (N_16280,N_13122,N_14451);
and U16281 (N_16281,N_11958,N_11265);
or U16282 (N_16282,N_13969,N_10666);
xor U16283 (N_16283,N_11473,N_10106);
or U16284 (N_16284,N_12234,N_12074);
nor U16285 (N_16285,N_11508,N_10953);
and U16286 (N_16286,N_11243,N_13281);
or U16287 (N_16287,N_12308,N_10567);
nor U16288 (N_16288,N_13856,N_11587);
nor U16289 (N_16289,N_12713,N_10766);
or U16290 (N_16290,N_12934,N_14787);
and U16291 (N_16291,N_11914,N_14386);
nand U16292 (N_16292,N_12358,N_12962);
xor U16293 (N_16293,N_14696,N_12874);
or U16294 (N_16294,N_11599,N_11098);
and U16295 (N_16295,N_14503,N_14650);
and U16296 (N_16296,N_11079,N_14247);
and U16297 (N_16297,N_11542,N_10478);
xnor U16298 (N_16298,N_10232,N_14535);
or U16299 (N_16299,N_12916,N_11408);
nand U16300 (N_16300,N_14868,N_11094);
and U16301 (N_16301,N_14044,N_10667);
nand U16302 (N_16302,N_13563,N_10455);
nor U16303 (N_16303,N_14270,N_10412);
and U16304 (N_16304,N_14115,N_13126);
xor U16305 (N_16305,N_11379,N_10885);
nand U16306 (N_16306,N_12504,N_10394);
nor U16307 (N_16307,N_11899,N_12819);
and U16308 (N_16308,N_12980,N_13703);
or U16309 (N_16309,N_13315,N_14842);
nand U16310 (N_16310,N_14698,N_14517);
or U16311 (N_16311,N_11786,N_14261);
nor U16312 (N_16312,N_14652,N_11865);
nor U16313 (N_16313,N_13291,N_11081);
nor U16314 (N_16314,N_14952,N_12567);
or U16315 (N_16315,N_14336,N_10202);
or U16316 (N_16316,N_11475,N_10852);
and U16317 (N_16317,N_13423,N_13698);
and U16318 (N_16318,N_13573,N_14465);
and U16319 (N_16319,N_11316,N_10156);
nor U16320 (N_16320,N_12126,N_12986);
nor U16321 (N_16321,N_10834,N_13700);
nand U16322 (N_16322,N_14807,N_10389);
nor U16323 (N_16323,N_14742,N_13159);
nand U16324 (N_16324,N_14858,N_11523);
and U16325 (N_16325,N_11993,N_12270);
or U16326 (N_16326,N_14629,N_10491);
and U16327 (N_16327,N_11101,N_14989);
xnor U16328 (N_16328,N_10208,N_13227);
nand U16329 (N_16329,N_13792,N_10355);
or U16330 (N_16330,N_13194,N_14551);
xor U16331 (N_16331,N_10684,N_12325);
nor U16332 (N_16332,N_13396,N_10039);
or U16333 (N_16333,N_13519,N_11344);
xnor U16334 (N_16334,N_13530,N_14427);
and U16335 (N_16335,N_14486,N_10599);
nor U16336 (N_16336,N_11332,N_13637);
nor U16337 (N_16337,N_11129,N_13491);
nor U16338 (N_16338,N_10871,N_12566);
nor U16339 (N_16339,N_14090,N_14841);
xor U16340 (N_16340,N_12972,N_11461);
or U16341 (N_16341,N_13604,N_14371);
nand U16342 (N_16342,N_13928,N_10776);
nand U16343 (N_16343,N_10094,N_10788);
or U16344 (N_16344,N_10300,N_12107);
nand U16345 (N_16345,N_10634,N_10011);
xnor U16346 (N_16346,N_13338,N_11854);
nor U16347 (N_16347,N_13222,N_13447);
and U16348 (N_16348,N_11506,N_12206);
or U16349 (N_16349,N_12685,N_12302);
nor U16350 (N_16350,N_10163,N_10729);
or U16351 (N_16351,N_14529,N_12409);
nor U16352 (N_16352,N_10069,N_12581);
xor U16353 (N_16353,N_10710,N_10006);
nor U16354 (N_16354,N_12965,N_10678);
xnor U16355 (N_16355,N_12461,N_14321);
and U16356 (N_16356,N_11242,N_14553);
nand U16357 (N_16357,N_10711,N_13803);
or U16358 (N_16358,N_11251,N_11090);
nand U16359 (N_16359,N_11688,N_14140);
or U16360 (N_16360,N_11776,N_10990);
nand U16361 (N_16361,N_13855,N_11425);
xnor U16362 (N_16362,N_11549,N_14307);
and U16363 (N_16363,N_14462,N_13214);
nor U16364 (N_16364,N_12488,N_10104);
nor U16365 (N_16365,N_13984,N_13106);
and U16366 (N_16366,N_11340,N_11829);
and U16367 (N_16367,N_11484,N_12220);
nand U16368 (N_16368,N_10433,N_12069);
xnor U16369 (N_16369,N_14958,N_11148);
nand U16370 (N_16370,N_10366,N_11191);
xor U16371 (N_16371,N_14908,N_11383);
and U16372 (N_16372,N_10239,N_12201);
and U16373 (N_16373,N_11269,N_10020);
or U16374 (N_16374,N_10016,N_13199);
nand U16375 (N_16375,N_12492,N_13730);
nor U16376 (N_16376,N_10655,N_11643);
or U16377 (N_16377,N_12921,N_12652);
xor U16378 (N_16378,N_10610,N_11365);
or U16379 (N_16379,N_13528,N_11869);
or U16380 (N_16380,N_11477,N_14525);
xor U16381 (N_16381,N_12291,N_14152);
nor U16382 (N_16382,N_12834,N_13111);
nand U16383 (N_16383,N_14292,N_12839);
and U16384 (N_16384,N_10057,N_11157);
nor U16385 (N_16385,N_11844,N_14183);
nor U16386 (N_16386,N_12165,N_14093);
and U16387 (N_16387,N_10882,N_10680);
and U16388 (N_16388,N_14499,N_10049);
xor U16389 (N_16389,N_10037,N_14588);
xor U16390 (N_16390,N_13892,N_10964);
xor U16391 (N_16391,N_12511,N_12365);
nand U16392 (N_16392,N_13004,N_12057);
and U16393 (N_16393,N_14545,N_12769);
xnor U16394 (N_16394,N_11464,N_12873);
nand U16395 (N_16395,N_10021,N_12716);
and U16396 (N_16396,N_14833,N_10979);
nand U16397 (N_16397,N_10819,N_13438);
and U16398 (N_16398,N_11873,N_14117);
nand U16399 (N_16399,N_14279,N_12780);
nor U16400 (N_16400,N_12080,N_12387);
xor U16401 (N_16401,N_13319,N_11851);
nand U16402 (N_16402,N_12695,N_13944);
nand U16403 (N_16403,N_14034,N_12831);
xnor U16404 (N_16404,N_12298,N_12513);
xnor U16405 (N_16405,N_12663,N_10027);
nor U16406 (N_16406,N_10100,N_13521);
nand U16407 (N_16407,N_14363,N_14467);
xnor U16408 (N_16408,N_12808,N_14255);
nor U16409 (N_16409,N_12105,N_13368);
nand U16410 (N_16410,N_11645,N_13632);
nor U16411 (N_16411,N_13670,N_14826);
nand U16412 (N_16412,N_12648,N_10172);
xor U16413 (N_16413,N_11253,N_12386);
nor U16414 (N_16414,N_11103,N_13276);
nand U16415 (N_16415,N_10161,N_13076);
xnor U16416 (N_16416,N_12239,N_13651);
or U16417 (N_16417,N_11018,N_14308);
and U16418 (N_16418,N_10611,N_11423);
xnor U16419 (N_16419,N_11543,N_14631);
nor U16420 (N_16420,N_14315,N_14762);
and U16421 (N_16421,N_10473,N_11575);
nor U16422 (N_16422,N_13615,N_11913);
nor U16423 (N_16423,N_12271,N_11697);
nor U16424 (N_16424,N_13976,N_13429);
and U16425 (N_16425,N_14012,N_12907);
xor U16426 (N_16426,N_12586,N_11089);
xor U16427 (N_16427,N_10768,N_14800);
nor U16428 (N_16428,N_12763,N_13745);
or U16429 (N_16429,N_14135,N_14411);
or U16430 (N_16430,N_11347,N_11290);
xnor U16431 (N_16431,N_10930,N_13465);
xnor U16432 (N_16432,N_12947,N_14176);
and U16433 (N_16433,N_12534,N_14786);
nor U16434 (N_16434,N_14021,N_11047);
and U16435 (N_16435,N_14498,N_14214);
nand U16436 (N_16436,N_12574,N_12955);
nand U16437 (N_16437,N_14381,N_12923);
nor U16438 (N_16438,N_10365,N_12445);
nand U16439 (N_16439,N_12312,N_13771);
xnor U16440 (N_16440,N_13804,N_10700);
nor U16441 (N_16441,N_13480,N_11884);
or U16442 (N_16442,N_13975,N_11588);
nand U16443 (N_16443,N_14959,N_10547);
or U16444 (N_16444,N_10157,N_14248);
nand U16445 (N_16445,N_11210,N_10301);
nand U16446 (N_16446,N_10561,N_13612);
and U16447 (N_16447,N_11113,N_12060);
or U16448 (N_16448,N_13113,N_11112);
and U16449 (N_16449,N_11948,N_13718);
nand U16450 (N_16450,N_13964,N_12638);
or U16451 (N_16451,N_10848,N_13680);
or U16452 (N_16452,N_13098,N_11398);
and U16453 (N_16453,N_13503,N_13166);
nor U16454 (N_16454,N_11033,N_13439);
and U16455 (N_16455,N_14107,N_12333);
or U16456 (N_16456,N_13526,N_14426);
and U16457 (N_16457,N_13273,N_14939);
or U16458 (N_16458,N_11109,N_14081);
nor U16459 (N_16459,N_14194,N_12078);
or U16460 (N_16460,N_14785,N_12391);
and U16461 (N_16461,N_11056,N_11584);
and U16462 (N_16462,N_14039,N_11162);
nand U16463 (N_16463,N_12837,N_11456);
or U16464 (N_16464,N_12787,N_10780);
nand U16465 (N_16465,N_14637,N_13820);
xor U16466 (N_16466,N_14400,N_13938);
nand U16467 (N_16467,N_10736,N_12315);
nand U16468 (N_16468,N_13230,N_14364);
nor U16469 (N_16469,N_10428,N_11111);
xor U16470 (N_16470,N_12480,N_10708);
nand U16471 (N_16471,N_10306,N_11476);
xor U16472 (N_16472,N_10869,N_11984);
xor U16473 (N_16473,N_14963,N_11678);
or U16474 (N_16474,N_13997,N_10309);
or U16475 (N_16475,N_14968,N_13302);
or U16476 (N_16476,N_13671,N_13164);
and U16477 (N_16477,N_10449,N_10609);
nand U16478 (N_16478,N_13542,N_12295);
and U16479 (N_16479,N_10786,N_12000);
nor U16480 (N_16480,N_12505,N_13324);
nor U16481 (N_16481,N_11614,N_12001);
nand U16482 (N_16482,N_12369,N_14661);
nand U16483 (N_16483,N_10594,N_11181);
nand U16484 (N_16484,N_12853,N_11806);
xor U16485 (N_16485,N_12125,N_14444);
nand U16486 (N_16486,N_12297,N_12052);
and U16487 (N_16487,N_10747,N_10265);
nand U16488 (N_16488,N_10072,N_11898);
nor U16489 (N_16489,N_11422,N_10087);
xor U16490 (N_16490,N_12922,N_12376);
nand U16491 (N_16491,N_14854,N_11359);
or U16492 (N_16492,N_13674,N_12925);
or U16493 (N_16493,N_12893,N_14560);
nand U16494 (N_16494,N_14712,N_13433);
nand U16495 (N_16495,N_12254,N_14450);
nor U16496 (N_16496,N_14520,N_10122);
xnor U16497 (N_16497,N_14625,N_10205);
and U16498 (N_16498,N_12166,N_12855);
nand U16499 (N_16499,N_13006,N_14532);
or U16500 (N_16500,N_11964,N_12605);
nor U16501 (N_16501,N_11130,N_13278);
or U16502 (N_16502,N_11052,N_12009);
and U16503 (N_16503,N_14990,N_10887);
xnor U16504 (N_16504,N_12482,N_11921);
xnor U16505 (N_16505,N_13228,N_14060);
xor U16506 (N_16506,N_10883,N_14319);
or U16507 (N_16507,N_14347,N_14598);
nand U16508 (N_16508,N_12416,N_14193);
nand U16509 (N_16509,N_13136,N_11683);
nand U16510 (N_16510,N_14167,N_14505);
or U16511 (N_16511,N_13767,N_12882);
nor U16512 (N_16512,N_14198,N_10297);
nor U16513 (N_16513,N_13645,N_12948);
and U16514 (N_16514,N_11434,N_14119);
and U16515 (N_16515,N_12215,N_14501);
and U16516 (N_16516,N_14635,N_11289);
nand U16517 (N_16517,N_12736,N_13064);
or U16518 (N_16518,N_12612,N_10315);
xnor U16519 (N_16519,N_13346,N_12949);
and U16520 (N_16520,N_10764,N_12450);
nor U16521 (N_16521,N_13974,N_14367);
nor U16522 (N_16522,N_11942,N_11437);
and U16523 (N_16523,N_13466,N_13985);
nand U16524 (N_16524,N_10409,N_13037);
nor U16525 (N_16525,N_10013,N_12020);
nand U16526 (N_16526,N_10813,N_10469);
or U16527 (N_16527,N_13301,N_11137);
or U16528 (N_16528,N_13587,N_13493);
and U16529 (N_16529,N_13235,N_10351);
and U16530 (N_16530,N_10195,N_10480);
nand U16531 (N_16531,N_12542,N_11782);
nand U16532 (N_16532,N_12745,N_10590);
xnor U16533 (N_16533,N_12359,N_10661);
nor U16534 (N_16534,N_10197,N_11771);
or U16535 (N_16535,N_13160,N_11886);
nor U16536 (N_16536,N_12506,N_12495);
nand U16537 (N_16537,N_11843,N_11013);
xnor U16538 (N_16538,N_13264,N_12751);
and U16539 (N_16539,N_11453,N_10946);
or U16540 (N_16540,N_12123,N_13100);
xnor U16541 (N_16541,N_11177,N_11981);
or U16542 (N_16542,N_12553,N_13249);
or U16543 (N_16543,N_10878,N_10055);
and U16544 (N_16544,N_10980,N_13658);
and U16545 (N_16545,N_10342,N_13890);
xnor U16546 (N_16546,N_13038,N_12863);
nor U16547 (N_16547,N_12959,N_13998);
or U16548 (N_16548,N_11378,N_12363);
nor U16549 (N_16549,N_13095,N_13580);
and U16550 (N_16550,N_11187,N_12563);
and U16551 (N_16551,N_11106,N_14810);
and U16552 (N_16552,N_14809,N_13387);
and U16553 (N_16553,N_11403,N_12028);
or U16554 (N_16554,N_12712,N_10579);
xor U16555 (N_16555,N_10165,N_13059);
xor U16556 (N_16556,N_13501,N_10801);
nand U16557 (N_16557,N_11740,N_11620);
or U16558 (N_16558,N_10752,N_13552);
nor U16559 (N_16559,N_13887,N_10400);
or U16560 (N_16560,N_11895,N_12294);
nand U16561 (N_16561,N_14647,N_14138);
or U16562 (N_16562,N_10388,N_13895);
nand U16563 (N_16563,N_11410,N_13391);
xnor U16564 (N_16564,N_11334,N_11724);
or U16565 (N_16565,N_14776,N_12205);
xor U16566 (N_16566,N_13268,N_12785);
xnor U16567 (N_16567,N_14112,N_10420);
nor U16568 (N_16568,N_14886,N_13742);
xor U16569 (N_16569,N_13363,N_11794);
or U16570 (N_16570,N_12276,N_14911);
or U16571 (N_16571,N_13601,N_10086);
xnor U16572 (N_16572,N_13436,N_10236);
and U16573 (N_16573,N_13314,N_12997);
xnor U16574 (N_16574,N_14583,N_13386);
or U16575 (N_16575,N_11876,N_14162);
and U16576 (N_16576,N_13440,N_12269);
nor U16577 (N_16577,N_10224,N_11718);
xor U16578 (N_16578,N_11507,N_12760);
or U16579 (N_16579,N_12396,N_12093);
xor U16580 (N_16580,N_11968,N_14897);
xor U16581 (N_16581,N_13657,N_11885);
nand U16582 (N_16582,N_11924,N_11791);
xnor U16583 (N_16583,N_11091,N_11041);
or U16584 (N_16584,N_10411,N_14557);
or U16585 (N_16585,N_13507,N_10516);
xnor U16586 (N_16586,N_13310,N_14941);
xor U16587 (N_16587,N_10513,N_11891);
and U16588 (N_16588,N_10696,N_10640);
nand U16589 (N_16589,N_13137,N_14988);
or U16590 (N_16590,N_11745,N_14639);
nand U16591 (N_16591,N_12994,N_13906);
and U16592 (N_16592,N_13785,N_13626);
or U16593 (N_16593,N_14345,N_12883);
nor U16594 (N_16594,N_10062,N_13896);
xor U16595 (N_16595,N_11691,N_10896);
and U16596 (N_16596,N_13275,N_12869);
nor U16597 (N_16597,N_11636,N_10448);
and U16598 (N_16598,N_14504,N_11800);
xnor U16599 (N_16599,N_14104,N_10468);
nand U16600 (N_16600,N_11160,N_12149);
xnor U16601 (N_16601,N_12334,N_14927);
xor U16602 (N_16602,N_13558,N_10999);
and U16603 (N_16603,N_13813,N_14326);
xnor U16604 (N_16604,N_11813,N_13559);
nor U16605 (N_16605,N_11293,N_12471);
nand U16606 (N_16606,N_14072,N_14417);
nor U16607 (N_16607,N_11590,N_12820);
and U16608 (N_16608,N_14118,N_11493);
nand U16609 (N_16609,N_13341,N_14047);
nand U16610 (N_16610,N_11626,N_14869);
or U16611 (N_16611,N_14710,N_14278);
and U16612 (N_16612,N_12545,N_14453);
xnor U16613 (N_16613,N_14124,N_12343);
or U16614 (N_16614,N_12489,N_12833);
or U16615 (N_16615,N_10906,N_10064);
xor U16616 (N_16616,N_11736,N_14463);
and U16617 (N_16617,N_10777,N_10822);
xnor U16618 (N_16618,N_12593,N_12415);
xor U16619 (N_16619,N_12299,N_13208);
or U16620 (N_16620,N_12507,N_10692);
or U16621 (N_16621,N_13533,N_10185);
nand U16622 (N_16622,N_12879,N_13780);
nor U16623 (N_16623,N_13287,N_11792);
nand U16624 (N_16624,N_12442,N_14867);
and U16625 (N_16625,N_13186,N_11928);
nand U16626 (N_16626,N_12658,N_11482);
xor U16627 (N_16627,N_10314,N_14025);
nand U16628 (N_16628,N_14686,N_14059);
xor U16629 (N_16629,N_13361,N_14685);
nand U16630 (N_16630,N_12841,N_11956);
or U16631 (N_16631,N_14043,N_11219);
or U16632 (N_16632,N_11666,N_10526);
nand U16633 (N_16633,N_10961,N_11431);
and U16634 (N_16634,N_11940,N_14478);
nor U16635 (N_16635,N_12765,N_10119);
nand U16636 (N_16636,N_12639,N_13865);
xnor U16637 (N_16637,N_11604,N_10089);
nor U16638 (N_16638,N_13331,N_12162);
or U16639 (N_16639,N_13699,N_14276);
nand U16640 (N_16640,N_10133,N_12623);
nor U16641 (N_16641,N_10835,N_13485);
nand U16642 (N_16642,N_13610,N_13937);
or U16643 (N_16643,N_12311,N_12496);
nand U16644 (N_16644,N_11284,N_13913);
nand U16645 (N_16645,N_13881,N_10387);
or U16646 (N_16646,N_12735,N_14566);
or U16647 (N_16647,N_13500,N_12243);
xor U16648 (N_16648,N_12904,N_14948);
and U16649 (N_16649,N_13269,N_11774);
nor U16650 (N_16650,N_12673,N_12444);
and U16651 (N_16651,N_13908,N_10383);
nand U16652 (N_16652,N_14141,N_13516);
and U16653 (N_16653,N_10346,N_14938);
nor U16654 (N_16654,N_12832,N_14306);
xnor U16655 (N_16655,N_10043,N_13216);
and U16656 (N_16656,N_10750,N_13206);
xnor U16657 (N_16657,N_10305,N_11202);
and U16658 (N_16658,N_12212,N_12101);
nand U16659 (N_16659,N_11292,N_10683);
or U16660 (N_16660,N_14171,N_11772);
or U16661 (N_16661,N_11621,N_11488);
xor U16662 (N_16662,N_13897,N_10724);
nor U16663 (N_16663,N_13880,N_13417);
and U16664 (N_16664,N_14614,N_10378);
and U16665 (N_16665,N_10271,N_12329);
and U16666 (N_16666,N_13940,N_13042);
or U16667 (N_16667,N_13989,N_13775);
nor U16668 (N_16668,N_10935,N_14624);
xnor U16669 (N_16669,N_12646,N_13574);
xnor U16670 (N_16670,N_10159,N_11196);
xnor U16671 (N_16671,N_10344,N_10914);
xor U16672 (N_16672,N_10701,N_14703);
nand U16673 (N_16673,N_12061,N_10656);
and U16674 (N_16674,N_13854,N_10490);
or U16675 (N_16675,N_11525,N_11773);
and U16676 (N_16676,N_14929,N_14076);
nor U16677 (N_16677,N_11552,N_13005);
or U16678 (N_16678,N_11199,N_10507);
nand U16679 (N_16679,N_11236,N_14048);
nand U16680 (N_16680,N_14662,N_14253);
and U16681 (N_16681,N_14851,N_12543);
nand U16682 (N_16682,N_12800,N_10214);
xor U16683 (N_16683,N_14779,N_10336);
xor U16684 (N_16684,N_11373,N_14828);
or U16685 (N_16685,N_11076,N_10406);
xor U16686 (N_16686,N_14905,N_10783);
nand U16687 (N_16687,N_12694,N_10789);
and U16688 (N_16688,N_13308,N_10327);
nand U16689 (N_16689,N_11577,N_13716);
and U16690 (N_16690,N_10749,N_11716);
xor U16691 (N_16691,N_13566,N_11788);
nand U16692 (N_16692,N_11260,N_13173);
xnor U16693 (N_16693,N_10231,N_13899);
and U16694 (N_16694,N_10676,N_14254);
nor U16695 (N_16695,N_11593,N_13705);
nor U16696 (N_16696,N_12788,N_10709);
nor U16697 (N_16697,N_10438,N_11370);
nor U16698 (N_16698,N_11965,N_13525);
nand U16699 (N_16699,N_14975,N_10733);
nand U16700 (N_16700,N_14302,N_10769);
and U16701 (N_16701,N_13717,N_12776);
nor U16702 (N_16702,N_11730,N_13217);
or U16703 (N_16703,N_14202,N_11288);
nor U16704 (N_16704,N_13786,N_12119);
and U16705 (N_16705,N_13616,N_10044);
nand U16706 (N_16706,N_11857,N_12128);
and U16707 (N_16707,N_10308,N_12041);
or U16708 (N_16708,N_11203,N_13411);
nor U16709 (N_16709,N_12006,N_11811);
xnor U16710 (N_16710,N_14105,N_14129);
and U16711 (N_16711,N_10190,N_11953);
xor U16712 (N_16712,N_13165,N_11935);
xor U16713 (N_16713,N_11513,N_10945);
nand U16714 (N_16714,N_12892,N_14724);
nor U16715 (N_16715,N_12013,N_12021);
nand U16716 (N_16716,N_11328,N_13335);
nor U16717 (N_16717,N_14110,N_12353);
xor U16718 (N_16718,N_13614,N_11863);
or U16719 (N_16719,N_12025,N_11546);
xor U16720 (N_16720,N_10565,N_13204);
nand U16721 (N_16721,N_14348,N_12512);
or U16722 (N_16722,N_13945,N_11828);
nand U16723 (N_16723,N_10997,N_11801);
nor U16724 (N_16724,N_12327,N_13135);
and U16725 (N_16725,N_12430,N_13863);
nor U16726 (N_16726,N_13261,N_14730);
xnor U16727 (N_16727,N_10534,N_12173);
xor U16728 (N_16728,N_13540,N_11933);
or U16729 (N_16729,N_14533,N_12067);
nand U16730 (N_16730,N_12503,N_12575);
xnor U16731 (N_16731,N_11582,N_12578);
and U16732 (N_16732,N_10674,N_10688);
and U16733 (N_16733,N_11128,N_14479);
nand U16734 (N_16734,N_14875,N_13664);
nor U16735 (N_16735,N_12144,N_11413);
and U16736 (N_16736,N_10360,N_14573);
and U16737 (N_16737,N_14679,N_12035);
xor U16738 (N_16738,N_13295,N_13756);
nand U16739 (N_16739,N_10255,N_11192);
xnor U16740 (N_16740,N_11114,N_12937);
and U16741 (N_16741,N_10441,N_12484);
nand U16742 (N_16742,N_11611,N_13995);
xor U16743 (N_16743,N_11352,N_10363);
or U16744 (N_16744,N_12175,N_11544);
nor U16745 (N_16745,N_11272,N_14291);
and U16746 (N_16746,N_11020,N_12984);
xnor U16747 (N_16747,N_11702,N_12576);
xor U16748 (N_16748,N_13296,N_10375);
or U16749 (N_16749,N_14863,N_14830);
nand U16750 (N_16750,N_11520,N_10844);
or U16751 (N_16751,N_14772,N_14397);
nand U16752 (N_16752,N_12142,N_12310);
or U16753 (N_16753,N_12434,N_12146);
and U16754 (N_16754,N_13797,N_13509);
or U16755 (N_16755,N_13830,N_14178);
or U16756 (N_16756,N_14601,N_10691);
and U16757 (N_16757,N_10182,N_14218);
nor U16758 (N_16758,N_12887,N_13025);
nand U16759 (N_16759,N_11246,N_11749);
nand U16760 (N_16760,N_10639,N_13834);
nand U16761 (N_16761,N_11186,N_10286);
nand U16762 (N_16762,N_11838,N_12609);
or U16763 (N_16763,N_12924,N_14829);
xnor U16764 (N_16764,N_14523,N_10658);
nand U16765 (N_16765,N_12791,N_13202);
nor U16766 (N_16766,N_12011,N_10967);
xnor U16767 (N_16767,N_11672,N_14204);
nor U16768 (N_16768,N_14335,N_13523);
nand U16769 (N_16769,N_14531,N_14904);
or U16770 (N_16770,N_11122,N_11208);
or U16771 (N_16771,N_11051,N_11753);
and U16772 (N_16772,N_14956,N_11310);
or U16773 (N_16773,N_10541,N_10569);
nand U16774 (N_16774,N_13990,N_11670);
xor U16775 (N_16775,N_11907,N_13097);
or U16776 (N_16776,N_14396,N_10950);
or U16777 (N_16777,N_11240,N_12345);
nand U16778 (N_16778,N_12796,N_13284);
and U16779 (N_16779,N_12410,N_13569);
nor U16780 (N_16780,N_12686,N_14832);
or U16781 (N_16781,N_12645,N_14387);
and U16782 (N_16782,N_14037,N_10109);
nand U16783 (N_16783,N_11846,N_11835);
nor U16784 (N_16784,N_10324,N_10874);
and U16785 (N_16785,N_14380,N_11802);
and U16786 (N_16786,N_11558,N_10379);
xor U16787 (N_16787,N_14312,N_10608);
nand U16788 (N_16788,N_12978,N_13886);
nor U16789 (N_16789,N_12725,N_12509);
xor U16790 (N_16790,N_13939,N_12397);
nor U16791 (N_16791,N_10920,N_12829);
nor U16792 (N_16792,N_11172,N_10173);
xor U16793 (N_16793,N_10071,N_11600);
and U16794 (N_16794,N_10266,N_13158);
and U16795 (N_16795,N_10152,N_12708);
or U16796 (N_16796,N_12927,N_12803);
or U16797 (N_16797,N_14885,N_12671);
or U16798 (N_16798,N_10805,N_12054);
nand U16799 (N_16799,N_12344,N_13132);
xor U16800 (N_16800,N_13826,N_10155);
nand U16801 (N_16801,N_13421,N_12627);
nor U16802 (N_16802,N_11147,N_13795);
or U16803 (N_16803,N_11983,N_14459);
or U16804 (N_16804,N_11171,N_14895);
nor U16805 (N_16805,N_11908,N_14861);
nor U16806 (N_16806,N_13912,N_12497);
or U16807 (N_16807,N_10268,N_13805);
nand U16808 (N_16808,N_10759,N_12818);
nand U16809 (N_16809,N_10671,N_11592);
and U16810 (N_16810,N_14790,N_13000);
and U16811 (N_16811,N_11896,N_14846);
nor U16812 (N_16812,N_10744,N_10390);
and U16813 (N_16813,N_11708,N_14009);
or U16814 (N_16814,N_10492,N_12199);
nand U16815 (N_16815,N_10785,N_13970);
nor U16816 (N_16816,N_14078,N_13999);
or U16817 (N_16817,N_11739,N_12368);
and U16818 (N_16818,N_13687,N_14303);
nor U16819 (N_16819,N_10452,N_14713);
nor U16820 (N_16820,N_10376,N_13941);
nand U16821 (N_16821,N_14094,N_11638);
and U16822 (N_16822,N_10123,N_13653);
nand U16823 (N_16823,N_13442,N_13358);
nand U16824 (N_16824,N_10931,N_14824);
or U16825 (N_16825,N_12273,N_10891);
nor U16826 (N_16826,N_11705,N_12641);
nor U16827 (N_16827,N_11936,N_13471);
and U16828 (N_16828,N_14177,N_10407);
or U16829 (N_16829,N_14228,N_12584);
nand U16830 (N_16830,N_13860,N_13364);
and U16831 (N_16831,N_12091,N_12446);
nand U16832 (N_16832,N_14654,N_13297);
xnor U16833 (N_16833,N_12139,N_13963);
and U16834 (N_16834,N_11432,N_14519);
nor U16835 (N_16835,N_13053,N_10851);
nand U16836 (N_16836,N_12253,N_12449);
xnor U16837 (N_16837,N_10687,N_13555);
or U16838 (N_16838,N_13755,N_14418);
nor U16839 (N_16839,N_10921,N_11877);
nor U16840 (N_16840,N_13401,N_14567);
nor U16841 (N_16841,N_11765,N_12522);
nand U16842 (N_16842,N_12871,N_10343);
nand U16843 (N_16843,N_12465,N_13001);
xnor U16844 (N_16844,N_12192,N_10083);
or U16845 (N_16845,N_11065,N_14784);
xor U16846 (N_16846,N_12798,N_14493);
and U16847 (N_16847,N_11775,N_10070);
xnor U16848 (N_16848,N_11087,N_14206);
nor U16849 (N_16849,N_14229,N_13825);
nor U16850 (N_16850,N_13508,N_12476);
nand U16851 (N_16851,N_13524,N_10035);
xor U16852 (N_16852,N_14502,N_13743);
xnor U16853 (N_16853,N_14215,N_12854);
xnor U16854 (N_16854,N_14443,N_10003);
and U16855 (N_16855,N_12526,N_10969);
nand U16856 (N_16856,N_14389,N_13978);
xnor U16857 (N_16857,N_14169,N_11389);
or U16858 (N_16858,N_13875,N_10149);
and U16859 (N_16859,N_10836,N_10527);
xor U16860 (N_16860,N_10845,N_11214);
nor U16861 (N_16861,N_12960,N_11754);
and U16862 (N_16862,N_14236,N_10147);
nand U16863 (N_16863,N_13549,N_13520);
and U16864 (N_16864,N_13565,N_11815);
and U16865 (N_16865,N_10963,N_11357);
nand U16866 (N_16866,N_11545,N_11987);
and U16867 (N_16867,N_11598,N_13255);
nor U16868 (N_16868,N_13229,N_11330);
or U16869 (N_16869,N_13355,N_13927);
or U16870 (N_16870,N_12121,N_10592);
xor U16871 (N_16871,N_14991,N_14633);
nand U16872 (N_16872,N_11973,N_12195);
and U16873 (N_16873,N_10453,N_14393);
nand U16874 (N_16874,N_11077,N_11812);
and U16875 (N_16875,N_11100,N_12935);
or U16876 (N_16876,N_14368,N_13369);
or U16877 (N_16877,N_10254,N_11367);
nor U16878 (N_16878,N_10993,N_12320);
and U16879 (N_16879,N_12050,N_10959);
xnor U16880 (N_16880,N_13591,N_13961);
and U16881 (N_16881,N_11063,N_14805);
or U16882 (N_16882,N_12264,N_14158);
or U16883 (N_16883,N_11889,N_14324);
nor U16884 (N_16884,N_11394,N_10868);
xor U16885 (N_16885,N_13459,N_13385);
and U16886 (N_16886,N_10329,N_13721);
nand U16887 (N_16887,N_12277,N_12679);
and U16888 (N_16888,N_10497,N_10566);
or U16889 (N_16889,N_10454,N_11447);
nand U16890 (N_16890,N_11376,N_11860);
nand U16891 (N_16891,N_10862,N_11388);
nor U16892 (N_16892,N_14069,N_13484);
nor U16893 (N_16893,N_13696,N_12411);
nand U16894 (N_16894,N_10038,N_14816);
or U16895 (N_16895,N_10371,N_10134);
or U16896 (N_16896,N_10380,N_14932);
nand U16897 (N_16897,N_13916,N_12113);
and U16898 (N_16898,N_10023,N_14645);
and U16899 (N_16899,N_10831,N_10463);
or U16900 (N_16900,N_10007,N_10402);
nor U16901 (N_16901,N_14350,N_10797);
nor U16902 (N_16902,N_12931,N_10212);
xnor U16903 (N_16903,N_13851,N_13091);
and U16904 (N_16904,N_10983,N_12991);
nand U16905 (N_16905,N_10019,N_10166);
xor U16906 (N_16906,N_14874,N_10554);
or U16907 (N_16907,N_10204,N_10005);
and U16908 (N_16908,N_14019,N_13968);
nor U16909 (N_16909,N_13120,N_13762);
and U16910 (N_16910,N_12692,N_10102);
and U16911 (N_16911,N_10784,N_14287);
nand U16912 (N_16912,N_12226,N_13920);
and U16913 (N_16913,N_14342,N_14723);
nand U16914 (N_16914,N_10201,N_11195);
nor U16915 (N_16915,N_14080,N_14663);
nand U16916 (N_16916,N_10466,N_11725);
xor U16917 (N_16917,N_10602,N_10034);
nor U16918 (N_16918,N_12881,N_13263);
and U16919 (N_16919,N_14665,N_14213);
xor U16920 (N_16920,N_14891,N_12370);
or U16921 (N_16921,N_11571,N_13740);
nor U16922 (N_16922,N_10540,N_13211);
and U16923 (N_16923,N_12589,N_13568);
or U16924 (N_16924,N_11918,N_14619);
nand U16925 (N_16925,N_12085,N_12042);
nor U16926 (N_16926,N_14157,N_10781);
nor U16927 (N_16927,N_14097,N_12437);
xor U16928 (N_16928,N_12667,N_13921);
xor U16929 (N_16929,N_14781,N_10903);
or U16930 (N_16930,N_12750,N_11684);
nand U16931 (N_16931,N_11654,N_14101);
and U16932 (N_16932,N_13077,N_11616);
and U16933 (N_16933,N_10372,N_14338);
or U16934 (N_16934,N_14782,N_12100);
and U16935 (N_16935,N_13778,N_10439);
or U16936 (N_16936,N_11462,N_11827);
or U16937 (N_16937,N_11755,N_11785);
nor U16938 (N_16938,N_11324,N_13016);
xnor U16939 (N_16939,N_13034,N_11667);
or U16940 (N_16940,N_11395,N_14974);
or U16941 (N_16941,N_13857,N_10180);
xor U16942 (N_16942,N_10474,N_11150);
nor U16943 (N_16943,N_14331,N_11075);
nand U16944 (N_16944,N_12866,N_12966);
and U16945 (N_16945,N_12772,N_13344);
and U16946 (N_16946,N_10311,N_13389);
and U16947 (N_16947,N_13724,N_12168);
nand U16948 (N_16948,N_10391,N_11647);
or U16949 (N_16949,N_14075,N_12908);
nand U16950 (N_16950,N_11990,N_10186);
or U16951 (N_16951,N_11733,N_12169);
and U16952 (N_16952,N_13772,N_13090);
nand U16953 (N_16953,N_13557,N_14582);
or U16954 (N_16954,N_13800,N_14844);
and U16955 (N_16955,N_14561,N_10414);
and U16956 (N_16956,N_14727,N_10568);
and U16957 (N_16957,N_13156,N_10704);
or U16958 (N_16958,N_13992,N_12546);
nand U16959 (N_16959,N_10717,N_12860);
and U16960 (N_16960,N_13492,N_14230);
and U16961 (N_16961,N_14541,N_14362);
nand U16962 (N_16962,N_12548,N_13668);
nor U16963 (N_16963,N_10557,N_12238);
or U16964 (N_16964,N_14982,N_13490);
nand U16965 (N_16965,N_14837,N_10732);
or U16966 (N_16966,N_12316,N_10447);
nand U16967 (N_16967,N_11957,N_12466);
or U16968 (N_16968,N_13441,N_13393);
xor U16969 (N_16969,N_10203,N_11499);
xnor U16970 (N_16970,N_10442,N_13738);
or U16971 (N_16971,N_13408,N_10905);
or U16972 (N_16972,N_14906,N_13824);
nor U16973 (N_16973,N_10303,N_14702);
nand U16974 (N_16974,N_14748,N_10879);
xnor U16975 (N_16975,N_10942,N_13720);
nor U16976 (N_16976,N_10753,N_14936);
xnor U16977 (N_16977,N_13427,N_12352);
xnor U16978 (N_16978,N_14086,N_13866);
and U16979 (N_16979,N_14244,N_12170);
or U16980 (N_16980,N_11433,N_10731);
xor U16981 (N_16981,N_12995,N_11701);
nand U16982 (N_16982,N_14848,N_12217);
nor U16983 (N_16983,N_14720,N_14376);
nand U16984 (N_16984,N_10132,N_14433);
or U16985 (N_16985,N_11807,N_13619);
and U16986 (N_16986,N_10601,N_10348);
nand U16987 (N_16987,N_11010,N_11559);
nand U16988 (N_16988,N_11970,N_11565);
nand U16989 (N_16989,N_14500,N_13822);
and U16990 (N_16990,N_14452,N_14677);
xor U16991 (N_16991,N_12470,N_12840);
or U16992 (N_16992,N_13641,N_10295);
or U16993 (N_16993,N_14222,N_12431);
xnor U16994 (N_16994,N_12055,N_10098);
and U16995 (N_16995,N_13183,N_13889);
or U16996 (N_16996,N_12844,N_12036);
and U16997 (N_16997,N_10694,N_13234);
and U16998 (N_16998,N_11107,N_10849);
nand U16999 (N_16999,N_12786,N_11349);
nand U17000 (N_17000,N_13634,N_12187);
nand U17001 (N_17001,N_11163,N_13061);
nor U17002 (N_17002,N_14552,N_10124);
xnor U17003 (N_17003,N_10418,N_14604);
nor U17004 (N_17004,N_13751,N_13326);
or U17005 (N_17005,N_14046,N_11596);
nor U17006 (N_17006,N_11249,N_14840);
xor U17007 (N_17007,N_13905,N_14487);
xnor U17008 (N_17008,N_11699,N_13769);
and U17009 (N_17009,N_11331,N_10030);
nand U17010 (N_17010,N_13828,N_13370);
nand U17011 (N_17011,N_10636,N_10092);
xor U17012 (N_17012,N_11748,N_13918);
xor U17013 (N_17013,N_11066,N_14208);
and U17014 (N_17014,N_13966,N_13621);
and U17015 (N_17015,N_13872,N_12388);
and U17016 (N_17016,N_10922,N_11345);
nor U17017 (N_17017,N_13141,N_14180);
nor U17018 (N_17018,N_10573,N_14468);
and U17019 (N_17019,N_10242,N_12022);
xnor U17020 (N_17020,N_13175,N_11674);
or U17021 (N_17021,N_13431,N_10248);
xor U17022 (N_17022,N_11008,N_14327);
or U17023 (N_17023,N_11673,N_13309);
or U17024 (N_17024,N_14490,N_14849);
and U17025 (N_17025,N_10320,N_14981);
and U17026 (N_17026,N_12588,N_10613);
nor U17027 (N_17027,N_13394,N_14656);
and U17028 (N_17028,N_10001,N_11073);
and U17029 (N_17029,N_10496,N_12406);
and U17030 (N_17030,N_10828,N_10618);
nand U17031 (N_17031,N_13110,N_12794);
xnor U17032 (N_17032,N_10814,N_10738);
or U17033 (N_17033,N_13936,N_12361);
or U17034 (N_17034,N_11409,N_12906);
nor U17035 (N_17035,N_13789,N_14860);
nor U17036 (N_17036,N_10322,N_14653);
xnor U17037 (N_17037,N_11427,N_10052);
and U17038 (N_17038,N_10457,N_10479);
nor U17039 (N_17039,N_11951,N_12134);
and U17040 (N_17040,N_11960,N_11693);
and U17041 (N_17041,N_12122,N_10495);
or U17042 (N_17042,N_13861,N_13420);
xnor U17043 (N_17043,N_14524,N_11897);
xnor U17044 (N_17044,N_12010,N_13635);
nor U17045 (N_17045,N_14497,N_14402);
and U17046 (N_17046,N_13665,N_11991);
nor U17047 (N_17047,N_11391,N_13163);
nand U17048 (N_17048,N_14611,N_14539);
nor U17049 (N_17049,N_12681,N_11441);
and U17050 (N_17050,N_12606,N_13242);
xor U17051 (N_17051,N_14460,N_14915);
and U17052 (N_17052,N_11305,N_10985);
nand U17053 (N_17053,N_14111,N_14884);
or U17054 (N_17054,N_14651,N_10517);
xor U17055 (N_17055,N_11814,N_11104);
xnor U17056 (N_17056,N_14937,N_13390);
and U17057 (N_17057,N_11216,N_14190);
xor U17058 (N_17058,N_12809,N_11304);
xnor U17059 (N_17059,N_14736,N_12094);
nor U17060 (N_17060,N_12637,N_14050);
nor U17061 (N_17061,N_11071,N_12381);
nand U17062 (N_17062,N_12458,N_14151);
and U17063 (N_17063,N_11115,N_13848);
nor U17064 (N_17064,N_14774,N_13807);
nand U17065 (N_17065,N_13841,N_12362);
xor U17066 (N_17066,N_10607,N_13178);
xor U17067 (N_17067,N_13371,N_10798);
or U17068 (N_17068,N_13919,N_14233);
nand U17069 (N_17069,N_13419,N_13212);
xnor U17070 (N_17070,N_10090,N_10338);
or U17071 (N_17071,N_13412,N_14283);
nor U17072 (N_17072,N_10475,N_13312);
nor U17073 (N_17073,N_10510,N_14067);
and U17074 (N_17074,N_12172,N_12571);
nor U17075 (N_17075,N_12082,N_10659);
nand U17076 (N_17076,N_12946,N_13849);
or U17077 (N_17077,N_14516,N_11108);
and U17078 (N_17078,N_13123,N_12537);
nand U17079 (N_17079,N_13625,N_11514);
nand U17080 (N_17080,N_10583,N_12112);
nand U17081 (N_17081,N_14265,N_12398);
nor U17082 (N_17082,N_11517,N_13407);
nor U17083 (N_17083,N_11152,N_14294);
nor U17084 (N_17084,N_10307,N_11027);
nand U17085 (N_17085,N_11034,N_11198);
nand U17086 (N_17086,N_11916,N_13087);
nor U17087 (N_17087,N_13435,N_10929);
xnor U17088 (N_17088,N_13181,N_10302);
or U17089 (N_17089,N_10949,N_13663);
nand U17090 (N_17090,N_12502,N_14596);
xor U17091 (N_17091,N_11954,N_10941);
nor U17092 (N_17092,N_11318,N_14113);
nand U17093 (N_17093,N_14422,N_10652);
xor U17094 (N_17094,N_11909,N_11068);
and U17095 (N_17095,N_12902,N_14998);
or U17096 (N_17096,N_12282,N_14643);
and U17097 (N_17097,N_14066,N_10673);
and U17098 (N_17098,N_10209,N_12558);
and U17099 (N_17099,N_12664,N_12037);
and U17100 (N_17100,N_11276,N_11826);
and U17101 (N_17101,N_11709,N_12933);
xor U17102 (N_17102,N_11337,N_14739);
or U17103 (N_17103,N_10292,N_13282);
or U17104 (N_17104,N_12901,N_11412);
xnor U17105 (N_17105,N_11211,N_14673);
nand U17106 (N_17106,N_12636,N_14226);
or U17107 (N_17107,N_13226,N_14145);
or U17108 (N_17108,N_14205,N_10904);
nand U17109 (N_17109,N_14033,N_14477);
or U17110 (N_17110,N_12757,N_11976);
xor U17111 (N_17111,N_10296,N_12508);
or U17112 (N_17112,N_13711,N_11648);
nor U17113 (N_17113,N_11439,N_13352);
xnor U17114 (N_17114,N_12930,N_14161);
and U17115 (N_17115,N_14298,N_14996);
and U17116 (N_17116,N_10519,N_12814);
and U17117 (N_17117,N_11595,N_13868);
nand U17118 (N_17118,N_11975,N_12117);
nand U17119 (N_17119,N_11174,N_11139);
xor U17120 (N_17120,N_14793,N_13256);
nand U17121 (N_17121,N_14799,N_10713);
nor U17122 (N_17122,N_10559,N_12953);
xnor U17123 (N_17123,N_14385,N_14120);
nor U17124 (N_17124,N_14301,N_12039);
xor U17125 (N_17125,N_12473,N_11356);
or U17126 (N_17126,N_13909,N_11904);
nor U17127 (N_17127,N_14160,N_10408);
nand U17128 (N_17128,N_14788,N_10506);
xnor U17129 (N_17129,N_10486,N_10103);
or U17130 (N_17130,N_12767,N_14108);
and U17131 (N_17131,N_12510,N_14360);
nand U17132 (N_17132,N_12944,N_12624);
nand U17133 (N_17133,N_11083,N_14668);
nor U17134 (N_17134,N_11222,N_11665);
nand U17135 (N_17135,N_13405,N_12385);
and U17136 (N_17136,N_12417,N_14544);
nor U17137 (N_17137,N_12857,N_10193);
nand U17138 (N_17138,N_12514,N_11072);
xor U17139 (N_17139,N_12810,N_14943);
xnor U17140 (N_17140,N_10403,N_10175);
or U17141 (N_17141,N_14944,N_11218);
and U17142 (N_17142,N_11719,N_10073);
or U17143 (N_17143,N_12975,N_13676);
nand U17144 (N_17144,N_12374,N_11301);
and U17145 (N_17145,N_13238,N_14838);
nor U17146 (N_17146,N_10141,N_12846);
nand U17147 (N_17147,N_10425,N_11006);
nor U17148 (N_17148,N_10646,N_13170);
xor U17149 (N_17149,N_12556,N_10870);
nor U17150 (N_17150,N_14556,N_10850);
or U17151 (N_17151,N_14751,N_11937);
xnor U17152 (N_17152,N_10290,N_10167);
or U17153 (N_17153,N_14877,N_12620);
nand U17154 (N_17154,N_11138,N_11706);
nor U17155 (N_17155,N_14224,N_11809);
and U17156 (N_17156,N_14188,N_13517);
xor U17157 (N_17157,N_13925,N_10988);
nor U17158 (N_17158,N_12267,N_11296);
or U17159 (N_17159,N_14313,N_11566);
xor U17160 (N_17160,N_14764,N_13131);
xnor U17161 (N_17161,N_11262,N_11069);
and U17162 (N_17162,N_13630,N_11095);
nand U17163 (N_17163,N_14607,N_10843);
nor U17164 (N_17164,N_13071,N_13758);
xnor U17165 (N_17165,N_12697,N_11610);
xor U17166 (N_17166,N_12649,N_12191);
nor U17167 (N_17167,N_12181,N_12383);
xor U17168 (N_17168,N_10287,N_13681);
or U17169 (N_17169,N_13983,N_11145);
xor U17170 (N_17170,N_13380,N_13911);
and U17171 (N_17171,N_12714,N_11241);
and U17172 (N_17172,N_11164,N_12266);
nor U17173 (N_17173,N_14822,N_12711);
xor U17174 (N_17174,N_11527,N_14859);
and U17175 (N_17175,N_13603,N_10289);
xnor U17176 (N_17176,N_10911,N_11625);
and U17177 (N_17177,N_13330,N_12811);
or U17178 (N_17178,N_11974,N_13378);
and U17179 (N_17179,N_10216,N_12401);
nor U17180 (N_17180,N_11713,N_11448);
xnor U17181 (N_17181,N_14378,N_10401);
and U17182 (N_17182,N_10998,N_12223);
and U17183 (N_17183,N_10544,N_11874);
xnor U17184 (N_17184,N_12547,N_10572);
nand U17185 (N_17185,N_14871,N_10291);
xor U17186 (N_17186,N_12454,N_13931);
xor U17187 (N_17187,N_14644,N_12221);
nor U17188 (N_17188,N_10832,N_14084);
nand U17189 (N_17189,N_10823,N_11986);
or U17190 (N_17190,N_10325,N_14136);
xnor U17191 (N_17191,N_13935,N_12213);
or U17192 (N_17192,N_10326,N_14055);
or U17193 (N_17193,N_12790,N_13835);
nand U17194 (N_17194,N_12516,N_11880);
nor U17195 (N_17195,N_14706,N_14466);
xnor U17196 (N_17196,N_14114,N_11631);
nor U17197 (N_17197,N_14692,N_14432);
and U17198 (N_17198,N_10461,N_12936);
or U17199 (N_17199,N_11479,N_12618);
and U17200 (N_17200,N_10746,N_12088);
nor U17201 (N_17201,N_10533,N_14812);
nand U17202 (N_17202,N_14030,N_11144);
xnor U17203 (N_17203,N_14014,N_12451);
or U17204 (N_17204,N_14309,N_12691);
nor U17205 (N_17205,N_10722,N_10857);
nor U17206 (N_17206,N_13678,N_13365);
nor U17207 (N_17207,N_14791,N_10253);
nand U17208 (N_17208,N_12634,N_12950);
nand U17209 (N_17209,N_13372,N_14933);
nand U17210 (N_17210,N_14734,N_14056);
nor U17211 (N_17211,N_14425,N_13185);
nand U17212 (N_17212,N_13629,N_13357);
nor U17213 (N_17213,N_10695,N_13013);
nor U17214 (N_17214,N_12099,N_14896);
and U17215 (N_17215,N_10962,N_13802);
or U17216 (N_17216,N_14761,N_12782);
nand U17217 (N_17217,N_11644,N_12038);
nand U17218 (N_17218,N_13060,N_12237);
or U17219 (N_17219,N_13951,N_14612);
nand U17220 (N_17220,N_10520,N_13511);
nand U17221 (N_17221,N_13458,N_12235);
or U17222 (N_17222,N_11784,N_10502);
and U17223 (N_17223,N_11707,N_14794);
xor U17224 (N_17224,N_11660,N_13776);
or U17225 (N_17225,N_13450,N_11470);
nand U17226 (N_17226,N_11459,N_12560);
nor U17227 (N_17227,N_13498,N_11502);
xnor U17228 (N_17228,N_12063,N_14257);
nand U17229 (N_17229,N_12533,N_10396);
xnor U17230 (N_17230,N_13647,N_11480);
xor U17231 (N_17231,N_12058,N_10549);
and U17232 (N_17232,N_12232,N_10933);
or U17233 (N_17233,N_14737,N_10499);
or U17234 (N_17234,N_11938,N_11257);
nand U17235 (N_17235,N_12153,N_11961);
nand U17236 (N_17236,N_12111,N_12895);
xor U17237 (N_17237,N_13464,N_10260);
and U17238 (N_17238,N_10410,N_12494);
or U17239 (N_17239,N_14569,N_10280);
and U17240 (N_17240,N_12371,N_11248);
nor U17241 (N_17241,N_11823,N_14957);
and U17242 (N_17242,N_12707,N_14914);
xnor U17243 (N_17243,N_14299,N_13207);
xnor U17244 (N_17244,N_12783,N_11436);
and U17245 (N_17245,N_14052,N_13168);
nand U17246 (N_17246,N_10545,N_13946);
xor U17247 (N_17247,N_11053,N_10880);
nor U17248 (N_17248,N_11711,N_10913);
and U17249 (N_17249,N_13406,N_10184);
nand U17250 (N_17250,N_10803,N_13709);
nor U17251 (N_17251,N_14721,N_11369);
or U17252 (N_17252,N_10483,N_13739);
xnor U17253 (N_17253,N_13777,N_13747);
nand U17254 (N_17254,N_11295,N_13505);
nand U17255 (N_17255,N_14166,N_10211);
or U17256 (N_17256,N_12130,N_14181);
nand U17257 (N_17257,N_14006,N_10293);
and U17258 (N_17258,N_10637,N_14334);
nand U17259 (N_17259,N_13712,N_13374);
nand U17260 (N_17260,N_14881,N_13483);
xor U17261 (N_17261,N_14245,N_13029);
nand U17262 (N_17262,N_10632,N_12940);
or U17263 (N_17263,N_14297,N_13215);
xor U17264 (N_17264,N_12070,N_12651);
or U17265 (N_17265,N_14749,N_13201);
and U17266 (N_17266,N_14471,N_13474);
nor U17267 (N_17267,N_13213,N_12806);
and U17268 (N_17268,N_14085,N_14910);
and U17269 (N_17269,N_10477,N_14880);
and U17270 (N_17270,N_10861,N_13597);
and U17271 (N_17271,N_13752,N_12989);
and U17272 (N_17272,N_10685,N_11279);
or U17273 (N_17273,N_12723,N_14295);
nor U17274 (N_17274,N_10413,N_13497);
or U17275 (N_17275,N_14305,N_12655);
or U17276 (N_17276,N_12868,N_13596);
and U17277 (N_17277,N_10863,N_10127);
or U17278 (N_17278,N_13379,N_11354);
or U17279 (N_17279,N_14700,N_13448);
xnor U17280 (N_17280,N_14131,N_14942);
or U17281 (N_17281,N_13642,N_10431);
xor U17282 (N_17282,N_14384,N_13972);
xnor U17283 (N_17283,N_12688,N_13351);
or U17284 (N_17284,N_14395,N_12118);
or U17285 (N_17285,N_12399,N_12075);
nand U17286 (N_17286,N_10616,N_14429);
nand U17287 (N_17287,N_14440,N_14195);
nor U17288 (N_17288,N_13304,N_11491);
nor U17289 (N_17289,N_12019,N_11959);
and U17290 (N_17290,N_12109,N_11945);
xor U17291 (N_17291,N_13452,N_10183);
nand U17292 (N_17292,N_10434,N_10081);
or U17293 (N_17293,N_12601,N_11615);
nand U17294 (N_17294,N_12479,N_13415);
and U17295 (N_17295,N_11910,N_10215);
and U17296 (N_17296,N_13348,N_10624);
nor U17297 (N_17297,N_11853,N_14924);
xor U17298 (N_17298,N_10153,N_14699);
and U17299 (N_17299,N_10121,N_12051);
or U17300 (N_17300,N_14134,N_13636);
and U17301 (N_17301,N_11004,N_11847);
or U17302 (N_17302,N_10787,N_12116);
xor U17303 (N_17303,N_11998,N_14613);
xnor U17304 (N_17304,N_11721,N_13144);
or U17305 (N_17305,N_14352,N_12876);
and U17306 (N_17306,N_14126,N_11836);
xor U17307 (N_17307,N_14916,N_14716);
xor U17308 (N_17308,N_10641,N_14149);
and U17309 (N_17309,N_14621,N_10033);
or U17310 (N_17310,N_13550,N_14087);
or U17311 (N_17311,N_11646,N_10116);
nand U17312 (N_17312,N_10174,N_13048);
nor U17313 (N_17313,N_13028,N_12599);
and U17314 (N_17314,N_10778,N_13218);
nand U17315 (N_17315,N_14058,N_11308);
nand U17316 (N_17316,N_14155,N_12336);
xor U17317 (N_17317,N_11326,N_12573);
nor U17318 (N_17318,N_10902,N_12771);
nor U17319 (N_17319,N_10230,N_13750);
xnor U17320 (N_17320,N_14879,N_10884);
nand U17321 (N_17321,N_14419,N_12676);
nand U17322 (N_17322,N_11963,N_10928);
nor U17323 (N_17323,N_14977,N_13749);
and U17324 (N_17324,N_11213,N_13043);
or U17325 (N_17325,N_14173,N_11734);
or U17326 (N_17326,N_13157,N_10221);
nand U17327 (N_17327,N_14455,N_12633);
and U17328 (N_17328,N_11390,N_13546);
nor U17329 (N_17329,N_12086,N_10643);
nor U17330 (N_17330,N_14655,N_14574);
nor U17331 (N_17331,N_11962,N_12394);
nand U17332 (N_17332,N_12137,N_10992);
nand U17333 (N_17333,N_14311,N_12597);
xnor U17334 (N_17334,N_14659,N_11510);
nand U17335 (N_17335,N_10117,N_14921);
xnor U17336 (N_17336,N_10058,N_14676);
nand U17337 (N_17337,N_13140,N_10827);
xor U17338 (N_17338,N_10036,N_14732);
xor U17339 (N_17339,N_13595,N_13257);
nor U17340 (N_17340,N_11311,N_13952);
nand U17341 (N_17341,N_13949,N_13850);
or U17342 (N_17342,N_12108,N_12103);
and U17343 (N_17343,N_13821,N_10393);
or U17344 (N_17344,N_12815,N_10257);
or U17345 (N_17345,N_10560,N_13862);
xnor U17346 (N_17346,N_14530,N_12158);
and U17347 (N_17347,N_14589,N_10370);
and U17348 (N_17348,N_11465,N_11429);
nand U17349 (N_17349,N_12017,N_12804);
nand U17350 (N_17350,N_11458,N_13639);
or U17351 (N_17351,N_10164,N_13791);
or U17352 (N_17352,N_12724,N_12357);
or U17353 (N_17353,N_11712,N_13947);
nor U17354 (N_17354,N_14599,N_13602);
nor U17355 (N_17355,N_13254,N_14189);
nand U17356 (N_17356,N_13434,N_11538);
xor U17357 (N_17357,N_14899,N_14170);
nand U17358 (N_17358,N_14103,N_14472);
xnor U17359 (N_17359,N_13154,N_11154);
xnor U17360 (N_17360,N_13317,N_12167);
nor U17361 (N_17361,N_10416,N_12413);
nor U17362 (N_17362,N_11627,N_13783);
nand U17363 (N_17363,N_13488,N_11197);
and U17364 (N_17364,N_13656,N_12207);
or U17365 (N_17365,N_12952,N_13377);
xor U17366 (N_17366,N_13649,N_12407);
nand U17367 (N_17367,N_11442,N_10191);
nor U17368 (N_17368,N_10225,N_13425);
nand U17369 (N_17369,N_14239,N_10635);
xnor U17370 (N_17370,N_14580,N_12053);
or U17371 (N_17371,N_14496,N_11364);
or U17372 (N_17372,N_10060,N_14883);
nor U17373 (N_17373,N_12602,N_14754);
nand U17374 (N_17374,N_11762,N_11029);
xnor U17375 (N_17375,N_14735,N_11449);
nor U17376 (N_17376,N_10354,N_12884);
or U17377 (N_17377,N_10518,N_13086);
or U17378 (N_17378,N_14045,N_12521);
nand U17379 (N_17379,N_11799,N_14745);
and U17380 (N_17380,N_13823,N_11501);
nor U17381 (N_17381,N_14857,N_12436);
nor U17382 (N_17382,N_13782,N_11789);
and U17383 (N_17383,N_11000,N_14366);
nand U17384 (N_17384,N_11322,N_11420);
nand U17385 (N_17385,N_13127,N_11223);
and U17386 (N_17386,N_10893,N_12720);
and U17387 (N_17387,N_12746,N_10597);
xor U17388 (N_17388,N_11564,N_14431);
and U17389 (N_17389,N_10047,N_14983);
or U17390 (N_17390,N_14768,N_13388);
nor U17391 (N_17391,N_10705,N_13114);
xor U17392 (N_17392,N_13643,N_13867);
and U17393 (N_17393,N_14064,N_14626);
xnor U17394 (N_17394,N_11120,N_12838);
xnor U17395 (N_17395,N_10115,N_14382);
xor U17396 (N_17396,N_11509,N_10472);
nor U17397 (N_17397,N_13770,N_10562);
or U17398 (N_17398,N_10128,N_11026);
nand U17399 (N_17399,N_11529,N_14373);
nand U17400 (N_17400,N_14558,N_10031);
and U17401 (N_17401,N_13883,N_11159);
and U17402 (N_17402,N_13481,N_13633);
xor U17403 (N_17403,N_11992,N_11633);
and U17404 (N_17404,N_12559,N_10958);
nor U17405 (N_17405,N_10806,N_12453);
or U17406 (N_17406,N_11355,N_11608);
nor U17407 (N_17407,N_12246,N_10690);
xnor U17408 (N_17408,N_12132,N_11859);
nand U17409 (N_17409,N_12300,N_12544);
nor U17410 (N_17410,N_12656,N_13589);
nand U17411 (N_17411,N_10316,N_14813);
and U17412 (N_17412,N_13066,N_11189);
nor U17413 (N_17413,N_14546,N_12528);
or U17414 (N_17414,N_10012,N_10716);
nand U17415 (N_17415,N_12642,N_12005);
xnor U17416 (N_17416,N_12915,N_11883);
xnor U17417 (N_17417,N_11858,N_14767);
nor U17418 (N_17418,N_10176,N_13561);
nor U17419 (N_17419,N_14483,N_13350);
xnor U17420 (N_17420,N_14361,N_11136);
and U17421 (N_17421,N_14887,N_12322);
or U17422 (N_17422,N_10682,N_12616);
and U17423 (N_17423,N_10970,N_12402);
or U17424 (N_17424,N_12147,N_14399);
nor U17425 (N_17425,N_12164,N_12174);
and U17426 (N_17426,N_14200,N_11474);
or U17427 (N_17427,N_13266,N_10919);
nand U17428 (N_17428,N_11460,N_11291);
and U17429 (N_17429,N_13967,N_12460);
nand U17430 (N_17430,N_13462,N_10160);
xnor U17431 (N_17431,N_14249,N_14733);
xnor U17432 (N_17432,N_12448,N_10792);
nand U17433 (N_17433,N_13339,N_13329);
and U17434 (N_17434,N_14622,N_11630);
and U17435 (N_17435,N_13036,N_13313);
nor U17436 (N_17436,N_14778,N_12632);
nor U17437 (N_17437,N_11255,N_12795);
or U17438 (N_17438,N_13283,N_10282);
nand U17439 (N_17439,N_11994,N_14852);
nand U17440 (N_17440,N_11206,N_14850);
or U17441 (N_17441,N_11180,N_12096);
or U17442 (N_17442,N_12928,N_13583);
or U17443 (N_17443,N_11032,N_10130);
nand U17444 (N_17444,N_13026,N_14562);
or U17445 (N_17445,N_11467,N_11703);
xnor U17446 (N_17446,N_11866,N_10965);
or U17447 (N_17447,N_12770,N_11204);
nor U17448 (N_17448,N_10194,N_12822);
xor U17449 (N_17449,N_11306,N_14971);
xor U17450 (N_17450,N_14518,N_12379);
and U17451 (N_17451,N_10493,N_11259);
or U17452 (N_17452,N_11852,N_14106);
xnor U17453 (N_17453,N_12603,N_10459);
nand U17454 (N_17454,N_11012,N_11917);
nor U17455 (N_17455,N_11088,N_13239);
nor U17456 (N_17456,N_11007,N_12541);
nor U17457 (N_17457,N_10482,N_13582);
or U17458 (N_17458,N_10818,N_14127);
xnor U17459 (N_17459,N_13965,N_10715);
and U17460 (N_17460,N_13934,N_11738);
xor U17461 (N_17461,N_10417,N_13859);
or U17462 (N_17462,N_11744,N_12487);
nor U17463 (N_17463,N_11624,N_14290);
or U17464 (N_17464,N_10571,N_13810);
nor U17465 (N_17465,N_13981,N_11757);
xnor U17466 (N_17466,N_14383,N_12631);
and U17467 (N_17467,N_12350,N_13307);
and U17468 (N_17468,N_13644,N_14137);
nor U17469 (N_17469,N_14273,N_13873);
or U17470 (N_17470,N_13142,N_12595);
xnor U17471 (N_17471,N_11263,N_12731);
nand U17472 (N_17472,N_11979,N_13763);
nor U17473 (N_17473,N_11878,N_11146);
and U17474 (N_17474,N_12233,N_12662);
nor U17475 (N_17475,N_14241,N_11952);
or U17476 (N_17476,N_12152,N_11512);
nand U17477 (N_17477,N_14955,N_12183);
or U17478 (N_17478,N_11902,N_11547);
xnor U17479 (N_17479,N_14457,N_11778);
and U17480 (N_17480,N_10895,N_10318);
or U17481 (N_17481,N_14489,N_14040);
or U17482 (N_17482,N_10754,N_13359);
or U17483 (N_17483,N_11696,N_13292);
or U17484 (N_17484,N_14572,N_14797);
nand U17485 (N_17485,N_14672,N_11803);
nor U17486 (N_17486,N_10285,N_13104);
nand U17487 (N_17487,N_12252,N_10578);
or U17488 (N_17488,N_11903,N_10552);
nand U17489 (N_17489,N_11619,N_14608);
nand U17490 (N_17490,N_13089,N_13414);
and U17491 (N_17491,N_14995,N_14554);
or U17492 (N_17492,N_11576,N_14722);
nand U17493 (N_17493,N_10500,N_13646);
nand U17494 (N_17494,N_10745,N_13993);
or U17495 (N_17495,N_10728,N_14962);
xor U17496 (N_17496,N_10984,N_12737);
and U17497 (N_17497,N_10765,N_14783);
xnor U17498 (N_17498,N_10890,N_14509);
nor U17499 (N_17499,N_11681,N_10989);
xnor U17500 (N_17500,N_12455,N_10426);
xor U17501 (N_17501,N_13437,N_11067);
xnor U17502 (N_17502,N_14885,N_12166);
and U17503 (N_17503,N_10676,N_12687);
xnor U17504 (N_17504,N_14975,N_10860);
nand U17505 (N_17505,N_13434,N_11046);
or U17506 (N_17506,N_10979,N_10429);
and U17507 (N_17507,N_10294,N_10184);
nor U17508 (N_17508,N_11745,N_14236);
xnor U17509 (N_17509,N_11884,N_11148);
or U17510 (N_17510,N_14952,N_14372);
or U17511 (N_17511,N_11162,N_14637);
and U17512 (N_17512,N_12171,N_14642);
nor U17513 (N_17513,N_10895,N_12162);
and U17514 (N_17514,N_11875,N_12060);
nand U17515 (N_17515,N_12651,N_13893);
and U17516 (N_17516,N_14110,N_12827);
or U17517 (N_17517,N_12030,N_10197);
nor U17518 (N_17518,N_13210,N_13401);
xor U17519 (N_17519,N_11420,N_13062);
xor U17520 (N_17520,N_14827,N_13943);
xnor U17521 (N_17521,N_11712,N_11787);
nor U17522 (N_17522,N_11902,N_11323);
or U17523 (N_17523,N_14030,N_10741);
or U17524 (N_17524,N_11012,N_13834);
xor U17525 (N_17525,N_10566,N_12213);
or U17526 (N_17526,N_12602,N_12277);
or U17527 (N_17527,N_14201,N_11300);
xnor U17528 (N_17528,N_12998,N_14543);
or U17529 (N_17529,N_12133,N_12207);
nor U17530 (N_17530,N_13393,N_11414);
and U17531 (N_17531,N_14221,N_12993);
nand U17532 (N_17532,N_12257,N_11852);
and U17533 (N_17533,N_14536,N_12581);
xor U17534 (N_17534,N_13825,N_13813);
xor U17535 (N_17535,N_14881,N_13198);
and U17536 (N_17536,N_13019,N_11575);
xor U17537 (N_17537,N_14178,N_12938);
and U17538 (N_17538,N_10464,N_10799);
and U17539 (N_17539,N_12436,N_12941);
and U17540 (N_17540,N_13039,N_10629);
or U17541 (N_17541,N_12045,N_14436);
nand U17542 (N_17542,N_13529,N_11627);
nor U17543 (N_17543,N_11632,N_11631);
or U17544 (N_17544,N_14379,N_13898);
and U17545 (N_17545,N_11678,N_14124);
or U17546 (N_17546,N_11252,N_10618);
nand U17547 (N_17547,N_12383,N_10024);
and U17548 (N_17548,N_10369,N_12013);
xor U17549 (N_17549,N_14422,N_11660);
nand U17550 (N_17550,N_11065,N_14819);
nor U17551 (N_17551,N_11450,N_14307);
nor U17552 (N_17552,N_11521,N_14527);
nor U17553 (N_17553,N_13803,N_10296);
and U17554 (N_17554,N_12325,N_11270);
and U17555 (N_17555,N_13173,N_12153);
nand U17556 (N_17556,N_14569,N_12333);
or U17557 (N_17557,N_11657,N_10296);
nand U17558 (N_17558,N_12096,N_11355);
xnor U17559 (N_17559,N_14160,N_11281);
nand U17560 (N_17560,N_10019,N_14228);
xor U17561 (N_17561,N_13114,N_14983);
and U17562 (N_17562,N_13589,N_11968);
xor U17563 (N_17563,N_12562,N_14818);
xnor U17564 (N_17564,N_11008,N_10446);
nor U17565 (N_17565,N_13469,N_12758);
xor U17566 (N_17566,N_14317,N_11911);
xor U17567 (N_17567,N_13447,N_11472);
nor U17568 (N_17568,N_12675,N_10939);
or U17569 (N_17569,N_10557,N_10346);
and U17570 (N_17570,N_10839,N_12591);
nand U17571 (N_17571,N_11736,N_13912);
or U17572 (N_17572,N_11821,N_12650);
nor U17573 (N_17573,N_14640,N_11055);
and U17574 (N_17574,N_11131,N_12188);
nor U17575 (N_17575,N_11091,N_11116);
nor U17576 (N_17576,N_11131,N_11033);
and U17577 (N_17577,N_13058,N_11268);
nand U17578 (N_17578,N_12649,N_12245);
nand U17579 (N_17579,N_13572,N_12258);
nand U17580 (N_17580,N_10624,N_14429);
xor U17581 (N_17581,N_12640,N_11249);
nand U17582 (N_17582,N_13052,N_11433);
xor U17583 (N_17583,N_10636,N_10287);
nor U17584 (N_17584,N_13994,N_11337);
nand U17585 (N_17585,N_14105,N_10810);
or U17586 (N_17586,N_13319,N_13454);
xnor U17587 (N_17587,N_12013,N_11994);
and U17588 (N_17588,N_13012,N_11149);
xor U17589 (N_17589,N_12480,N_11778);
nand U17590 (N_17590,N_14571,N_14887);
or U17591 (N_17591,N_11149,N_12117);
and U17592 (N_17592,N_10270,N_10714);
nor U17593 (N_17593,N_13572,N_10518);
xnor U17594 (N_17594,N_12286,N_14621);
xor U17595 (N_17595,N_10773,N_13705);
nor U17596 (N_17596,N_11147,N_11866);
xor U17597 (N_17597,N_14648,N_10511);
nor U17598 (N_17598,N_12683,N_13326);
and U17599 (N_17599,N_14703,N_14148);
nor U17600 (N_17600,N_13146,N_10065);
or U17601 (N_17601,N_14604,N_11051);
xnor U17602 (N_17602,N_10607,N_10312);
nand U17603 (N_17603,N_14929,N_11460);
and U17604 (N_17604,N_12651,N_13277);
nand U17605 (N_17605,N_14130,N_12320);
and U17606 (N_17606,N_12947,N_13875);
xnor U17607 (N_17607,N_14231,N_10387);
or U17608 (N_17608,N_14811,N_12960);
or U17609 (N_17609,N_11486,N_12702);
nor U17610 (N_17610,N_14447,N_12736);
or U17611 (N_17611,N_12557,N_10206);
nand U17612 (N_17612,N_10211,N_13272);
nand U17613 (N_17613,N_13715,N_13315);
or U17614 (N_17614,N_13628,N_14412);
or U17615 (N_17615,N_11076,N_12427);
xnor U17616 (N_17616,N_12416,N_11848);
and U17617 (N_17617,N_10107,N_10841);
xor U17618 (N_17618,N_13754,N_10751);
xor U17619 (N_17619,N_10818,N_13126);
nand U17620 (N_17620,N_13753,N_11089);
nand U17621 (N_17621,N_14178,N_13999);
xor U17622 (N_17622,N_11328,N_10084);
nand U17623 (N_17623,N_11132,N_14376);
and U17624 (N_17624,N_12104,N_11514);
nor U17625 (N_17625,N_14614,N_11149);
nand U17626 (N_17626,N_10395,N_11401);
or U17627 (N_17627,N_14767,N_12478);
xnor U17628 (N_17628,N_10489,N_10337);
xnor U17629 (N_17629,N_10814,N_10290);
nand U17630 (N_17630,N_10350,N_11598);
or U17631 (N_17631,N_11583,N_14862);
nor U17632 (N_17632,N_11906,N_10746);
nand U17633 (N_17633,N_13553,N_13793);
nor U17634 (N_17634,N_10096,N_11524);
and U17635 (N_17635,N_12251,N_12543);
and U17636 (N_17636,N_14358,N_13100);
or U17637 (N_17637,N_13519,N_10205);
nand U17638 (N_17638,N_13582,N_14806);
nor U17639 (N_17639,N_14930,N_13234);
and U17640 (N_17640,N_14287,N_11150);
and U17641 (N_17641,N_12884,N_10828);
and U17642 (N_17642,N_13198,N_13861);
xnor U17643 (N_17643,N_12907,N_10262);
nor U17644 (N_17644,N_14799,N_10285);
nand U17645 (N_17645,N_11229,N_10962);
nor U17646 (N_17646,N_11957,N_12650);
xnor U17647 (N_17647,N_14674,N_12049);
nor U17648 (N_17648,N_13666,N_14768);
nand U17649 (N_17649,N_10042,N_11290);
nor U17650 (N_17650,N_11056,N_12465);
nor U17651 (N_17651,N_11399,N_13398);
nand U17652 (N_17652,N_12377,N_12337);
nand U17653 (N_17653,N_13572,N_13521);
xor U17654 (N_17654,N_14194,N_11641);
and U17655 (N_17655,N_14233,N_13866);
xor U17656 (N_17656,N_11339,N_13468);
nor U17657 (N_17657,N_14828,N_11934);
and U17658 (N_17658,N_14225,N_10919);
nor U17659 (N_17659,N_14823,N_13912);
xor U17660 (N_17660,N_13544,N_14408);
nand U17661 (N_17661,N_12609,N_12620);
nand U17662 (N_17662,N_14021,N_10113);
nand U17663 (N_17663,N_14384,N_14692);
xnor U17664 (N_17664,N_14482,N_14267);
xnor U17665 (N_17665,N_11402,N_12204);
nor U17666 (N_17666,N_14148,N_11683);
and U17667 (N_17667,N_11349,N_10650);
xnor U17668 (N_17668,N_12724,N_10777);
or U17669 (N_17669,N_10636,N_13583);
nand U17670 (N_17670,N_14616,N_14662);
xor U17671 (N_17671,N_14060,N_10413);
xor U17672 (N_17672,N_12631,N_11175);
nand U17673 (N_17673,N_11845,N_14776);
and U17674 (N_17674,N_12512,N_10133);
nor U17675 (N_17675,N_12112,N_13944);
and U17676 (N_17676,N_14994,N_14372);
and U17677 (N_17677,N_10815,N_13619);
or U17678 (N_17678,N_13520,N_11876);
or U17679 (N_17679,N_10295,N_14436);
nor U17680 (N_17680,N_13501,N_12468);
or U17681 (N_17681,N_10952,N_10889);
xor U17682 (N_17682,N_11446,N_10183);
xor U17683 (N_17683,N_13073,N_14840);
nor U17684 (N_17684,N_13348,N_14283);
or U17685 (N_17685,N_13141,N_13171);
and U17686 (N_17686,N_12336,N_11436);
nor U17687 (N_17687,N_14924,N_12512);
or U17688 (N_17688,N_13949,N_11780);
or U17689 (N_17689,N_12205,N_12088);
nor U17690 (N_17690,N_12986,N_12176);
nor U17691 (N_17691,N_14825,N_14606);
and U17692 (N_17692,N_11164,N_10763);
xnor U17693 (N_17693,N_13035,N_10136);
or U17694 (N_17694,N_10287,N_11244);
or U17695 (N_17695,N_13058,N_11535);
nand U17696 (N_17696,N_10746,N_10828);
xnor U17697 (N_17697,N_12530,N_12639);
xor U17698 (N_17698,N_12825,N_13132);
or U17699 (N_17699,N_10067,N_10886);
nor U17700 (N_17700,N_14214,N_11999);
nor U17701 (N_17701,N_14662,N_12651);
or U17702 (N_17702,N_11583,N_11023);
xor U17703 (N_17703,N_14795,N_10488);
and U17704 (N_17704,N_10445,N_13100);
xnor U17705 (N_17705,N_13452,N_13809);
or U17706 (N_17706,N_11054,N_11206);
nand U17707 (N_17707,N_11400,N_10488);
xor U17708 (N_17708,N_11519,N_11786);
or U17709 (N_17709,N_11481,N_11880);
or U17710 (N_17710,N_11366,N_12022);
or U17711 (N_17711,N_12851,N_12266);
xor U17712 (N_17712,N_12717,N_14485);
and U17713 (N_17713,N_11013,N_11832);
and U17714 (N_17714,N_13167,N_14417);
nor U17715 (N_17715,N_11748,N_10806);
and U17716 (N_17716,N_13777,N_10677);
nor U17717 (N_17717,N_12130,N_13503);
and U17718 (N_17718,N_14978,N_10054);
nand U17719 (N_17719,N_12880,N_10640);
nor U17720 (N_17720,N_14830,N_10229);
xnor U17721 (N_17721,N_13531,N_10512);
or U17722 (N_17722,N_11568,N_14773);
nor U17723 (N_17723,N_13396,N_12640);
and U17724 (N_17724,N_11421,N_12940);
or U17725 (N_17725,N_11494,N_11667);
and U17726 (N_17726,N_12562,N_10554);
nand U17727 (N_17727,N_12815,N_13444);
nor U17728 (N_17728,N_12983,N_10161);
and U17729 (N_17729,N_13522,N_13028);
xnor U17730 (N_17730,N_11195,N_12687);
xor U17731 (N_17731,N_11771,N_11823);
xnor U17732 (N_17732,N_14821,N_14160);
nor U17733 (N_17733,N_11404,N_14476);
nand U17734 (N_17734,N_13375,N_12982);
and U17735 (N_17735,N_11374,N_14814);
and U17736 (N_17736,N_14208,N_14004);
and U17737 (N_17737,N_10309,N_12976);
nand U17738 (N_17738,N_14388,N_14296);
and U17739 (N_17739,N_13914,N_11877);
xnor U17740 (N_17740,N_13283,N_14937);
xor U17741 (N_17741,N_12987,N_11229);
nand U17742 (N_17742,N_14088,N_12525);
nor U17743 (N_17743,N_11597,N_10603);
or U17744 (N_17744,N_12409,N_13456);
or U17745 (N_17745,N_12715,N_11448);
xor U17746 (N_17746,N_10711,N_11901);
or U17747 (N_17747,N_14869,N_11827);
nand U17748 (N_17748,N_10309,N_13139);
nor U17749 (N_17749,N_14789,N_10873);
nor U17750 (N_17750,N_14790,N_11387);
nand U17751 (N_17751,N_13331,N_10514);
nand U17752 (N_17752,N_11239,N_11069);
or U17753 (N_17753,N_13683,N_14003);
and U17754 (N_17754,N_11724,N_10080);
xnor U17755 (N_17755,N_13495,N_10202);
nand U17756 (N_17756,N_12479,N_11856);
or U17757 (N_17757,N_14209,N_13946);
and U17758 (N_17758,N_14093,N_10062);
nor U17759 (N_17759,N_13652,N_14668);
nor U17760 (N_17760,N_14756,N_13406);
nor U17761 (N_17761,N_11956,N_13360);
nor U17762 (N_17762,N_10851,N_13247);
nand U17763 (N_17763,N_11460,N_12006);
xor U17764 (N_17764,N_13668,N_14549);
and U17765 (N_17765,N_13746,N_13115);
and U17766 (N_17766,N_12032,N_13570);
xor U17767 (N_17767,N_11834,N_10045);
nor U17768 (N_17768,N_14496,N_13081);
xnor U17769 (N_17769,N_11824,N_14048);
or U17770 (N_17770,N_14161,N_14794);
and U17771 (N_17771,N_11193,N_10458);
nor U17772 (N_17772,N_14332,N_12581);
xor U17773 (N_17773,N_10745,N_12992);
nor U17774 (N_17774,N_13127,N_11389);
and U17775 (N_17775,N_14383,N_13787);
nor U17776 (N_17776,N_10540,N_12036);
and U17777 (N_17777,N_11123,N_13346);
nor U17778 (N_17778,N_13075,N_12466);
and U17779 (N_17779,N_14119,N_10080);
nor U17780 (N_17780,N_13561,N_10685);
nand U17781 (N_17781,N_12076,N_13258);
nor U17782 (N_17782,N_12895,N_13336);
and U17783 (N_17783,N_13677,N_11549);
nand U17784 (N_17784,N_10105,N_14724);
nand U17785 (N_17785,N_11367,N_10642);
and U17786 (N_17786,N_14118,N_11585);
and U17787 (N_17787,N_14684,N_14501);
xnor U17788 (N_17788,N_14537,N_11234);
and U17789 (N_17789,N_13852,N_14345);
and U17790 (N_17790,N_14622,N_14764);
or U17791 (N_17791,N_11371,N_14478);
xor U17792 (N_17792,N_10646,N_14346);
nor U17793 (N_17793,N_13425,N_12717);
and U17794 (N_17794,N_11494,N_14129);
or U17795 (N_17795,N_11186,N_11490);
or U17796 (N_17796,N_10757,N_14029);
or U17797 (N_17797,N_10012,N_11177);
nor U17798 (N_17798,N_13910,N_12086);
and U17799 (N_17799,N_11931,N_12127);
and U17800 (N_17800,N_11128,N_14123);
xnor U17801 (N_17801,N_11751,N_12647);
nand U17802 (N_17802,N_13926,N_14087);
xor U17803 (N_17803,N_13477,N_14508);
and U17804 (N_17804,N_12500,N_11857);
xnor U17805 (N_17805,N_10074,N_11425);
and U17806 (N_17806,N_12549,N_11935);
nand U17807 (N_17807,N_13380,N_13062);
or U17808 (N_17808,N_12665,N_10304);
nor U17809 (N_17809,N_10884,N_10723);
nand U17810 (N_17810,N_11445,N_10648);
and U17811 (N_17811,N_14185,N_10314);
and U17812 (N_17812,N_12446,N_13700);
nand U17813 (N_17813,N_13304,N_12289);
and U17814 (N_17814,N_14320,N_11879);
and U17815 (N_17815,N_12329,N_13198);
or U17816 (N_17816,N_14905,N_13856);
nor U17817 (N_17817,N_12355,N_11578);
nand U17818 (N_17818,N_10770,N_11961);
nor U17819 (N_17819,N_13297,N_14077);
or U17820 (N_17820,N_13970,N_14311);
nand U17821 (N_17821,N_14044,N_13865);
xnor U17822 (N_17822,N_10775,N_11061);
or U17823 (N_17823,N_14568,N_12336);
nand U17824 (N_17824,N_11724,N_12942);
nor U17825 (N_17825,N_14376,N_11196);
xnor U17826 (N_17826,N_10079,N_10819);
and U17827 (N_17827,N_13816,N_11117);
and U17828 (N_17828,N_10161,N_13874);
and U17829 (N_17829,N_10757,N_10787);
xnor U17830 (N_17830,N_14257,N_11546);
and U17831 (N_17831,N_12640,N_14660);
xor U17832 (N_17832,N_11370,N_13301);
nand U17833 (N_17833,N_14987,N_13929);
or U17834 (N_17834,N_11969,N_14076);
and U17835 (N_17835,N_13707,N_12783);
or U17836 (N_17836,N_12423,N_11094);
and U17837 (N_17837,N_12716,N_13146);
xnor U17838 (N_17838,N_13026,N_14055);
or U17839 (N_17839,N_14398,N_14376);
nand U17840 (N_17840,N_11028,N_13441);
xnor U17841 (N_17841,N_12553,N_14527);
or U17842 (N_17842,N_11478,N_12262);
xor U17843 (N_17843,N_14673,N_12464);
nor U17844 (N_17844,N_14371,N_13139);
and U17845 (N_17845,N_12906,N_12784);
nor U17846 (N_17846,N_14255,N_12271);
xor U17847 (N_17847,N_13111,N_13741);
nand U17848 (N_17848,N_10819,N_12735);
and U17849 (N_17849,N_12443,N_14031);
nand U17850 (N_17850,N_12713,N_11363);
nand U17851 (N_17851,N_12535,N_10082);
xor U17852 (N_17852,N_13180,N_12580);
nand U17853 (N_17853,N_11164,N_12188);
nor U17854 (N_17854,N_10805,N_11798);
nor U17855 (N_17855,N_14436,N_12565);
or U17856 (N_17856,N_13786,N_14865);
and U17857 (N_17857,N_10448,N_12287);
nand U17858 (N_17858,N_12575,N_10963);
and U17859 (N_17859,N_14348,N_12519);
nand U17860 (N_17860,N_12244,N_14775);
and U17861 (N_17861,N_13727,N_13001);
nor U17862 (N_17862,N_14820,N_11271);
or U17863 (N_17863,N_14251,N_14545);
xnor U17864 (N_17864,N_10414,N_10551);
or U17865 (N_17865,N_11190,N_14949);
xor U17866 (N_17866,N_13597,N_14706);
nand U17867 (N_17867,N_12348,N_11420);
nand U17868 (N_17868,N_14988,N_14334);
nor U17869 (N_17869,N_11956,N_11886);
and U17870 (N_17870,N_12665,N_13070);
nand U17871 (N_17871,N_10838,N_10848);
nor U17872 (N_17872,N_13693,N_13561);
xnor U17873 (N_17873,N_13620,N_14787);
or U17874 (N_17874,N_14997,N_13390);
nand U17875 (N_17875,N_12218,N_12950);
xnor U17876 (N_17876,N_11061,N_14325);
nor U17877 (N_17877,N_12829,N_11549);
or U17878 (N_17878,N_10423,N_14643);
nand U17879 (N_17879,N_10408,N_10822);
xnor U17880 (N_17880,N_14513,N_11671);
or U17881 (N_17881,N_13390,N_12071);
nand U17882 (N_17882,N_13641,N_12417);
or U17883 (N_17883,N_14292,N_14475);
or U17884 (N_17884,N_11469,N_12716);
xnor U17885 (N_17885,N_10504,N_10422);
nand U17886 (N_17886,N_12368,N_14267);
or U17887 (N_17887,N_11828,N_10464);
or U17888 (N_17888,N_11103,N_11088);
nor U17889 (N_17889,N_10270,N_11276);
nand U17890 (N_17890,N_10057,N_13032);
and U17891 (N_17891,N_14968,N_14748);
xnor U17892 (N_17892,N_10294,N_14307);
or U17893 (N_17893,N_11984,N_14263);
nor U17894 (N_17894,N_12250,N_10849);
nand U17895 (N_17895,N_12761,N_12103);
nor U17896 (N_17896,N_13372,N_11721);
nand U17897 (N_17897,N_14246,N_14784);
nand U17898 (N_17898,N_13163,N_10734);
or U17899 (N_17899,N_11571,N_11490);
or U17900 (N_17900,N_11806,N_12063);
xor U17901 (N_17901,N_12068,N_13001);
or U17902 (N_17902,N_10661,N_14623);
or U17903 (N_17903,N_12270,N_11052);
or U17904 (N_17904,N_11006,N_10808);
xor U17905 (N_17905,N_11867,N_10671);
xor U17906 (N_17906,N_13560,N_14211);
or U17907 (N_17907,N_12564,N_14562);
and U17908 (N_17908,N_10983,N_14088);
nand U17909 (N_17909,N_11493,N_14000);
nor U17910 (N_17910,N_13744,N_12807);
nand U17911 (N_17911,N_14389,N_10239);
xor U17912 (N_17912,N_13806,N_11383);
xnor U17913 (N_17913,N_10592,N_13067);
or U17914 (N_17914,N_13477,N_12369);
nand U17915 (N_17915,N_10543,N_14708);
nand U17916 (N_17916,N_14847,N_12851);
nor U17917 (N_17917,N_10430,N_11255);
and U17918 (N_17918,N_13489,N_12809);
nor U17919 (N_17919,N_13801,N_13669);
and U17920 (N_17920,N_12883,N_13835);
nand U17921 (N_17921,N_11042,N_14093);
or U17922 (N_17922,N_10134,N_12354);
nand U17923 (N_17923,N_10013,N_10223);
or U17924 (N_17924,N_11290,N_11858);
nand U17925 (N_17925,N_14254,N_12611);
nor U17926 (N_17926,N_14794,N_11936);
xor U17927 (N_17927,N_10560,N_11916);
xnor U17928 (N_17928,N_11765,N_14084);
nor U17929 (N_17929,N_13773,N_11005);
or U17930 (N_17930,N_12029,N_12490);
or U17931 (N_17931,N_14622,N_10345);
nor U17932 (N_17932,N_13061,N_13641);
nor U17933 (N_17933,N_10182,N_10269);
or U17934 (N_17934,N_13671,N_13769);
xnor U17935 (N_17935,N_14198,N_12904);
nand U17936 (N_17936,N_12749,N_10098);
nand U17937 (N_17937,N_12555,N_10778);
or U17938 (N_17938,N_10090,N_14233);
nand U17939 (N_17939,N_14746,N_12776);
xnor U17940 (N_17940,N_14569,N_14001);
and U17941 (N_17941,N_11525,N_14271);
and U17942 (N_17942,N_13542,N_10363);
nand U17943 (N_17943,N_14948,N_11717);
nor U17944 (N_17944,N_11309,N_13446);
nand U17945 (N_17945,N_10051,N_14739);
and U17946 (N_17946,N_11286,N_12892);
and U17947 (N_17947,N_12571,N_11308);
xor U17948 (N_17948,N_11903,N_12172);
xor U17949 (N_17949,N_12476,N_12783);
xor U17950 (N_17950,N_13826,N_10559);
nand U17951 (N_17951,N_12911,N_14555);
nand U17952 (N_17952,N_12165,N_10026);
or U17953 (N_17953,N_12629,N_14897);
xor U17954 (N_17954,N_11629,N_10791);
nor U17955 (N_17955,N_10427,N_12741);
nor U17956 (N_17956,N_13521,N_13582);
or U17957 (N_17957,N_11963,N_12653);
and U17958 (N_17958,N_12041,N_14374);
or U17959 (N_17959,N_14268,N_13628);
or U17960 (N_17960,N_10806,N_14265);
nand U17961 (N_17961,N_10506,N_10196);
and U17962 (N_17962,N_13062,N_12283);
xor U17963 (N_17963,N_12038,N_10336);
and U17964 (N_17964,N_10229,N_12402);
nand U17965 (N_17965,N_12106,N_12083);
and U17966 (N_17966,N_11868,N_12130);
nand U17967 (N_17967,N_13703,N_13691);
nor U17968 (N_17968,N_10778,N_10506);
and U17969 (N_17969,N_11687,N_11714);
nand U17970 (N_17970,N_10981,N_11513);
nand U17971 (N_17971,N_11119,N_14308);
nand U17972 (N_17972,N_12043,N_11000);
xor U17973 (N_17973,N_13037,N_11652);
or U17974 (N_17974,N_10277,N_13209);
nand U17975 (N_17975,N_11747,N_11734);
nand U17976 (N_17976,N_13458,N_10998);
nand U17977 (N_17977,N_13868,N_13367);
or U17978 (N_17978,N_10527,N_13503);
nor U17979 (N_17979,N_10610,N_13729);
nand U17980 (N_17980,N_12539,N_11176);
and U17981 (N_17981,N_10695,N_14557);
xnor U17982 (N_17982,N_11097,N_12770);
nor U17983 (N_17983,N_10754,N_11333);
or U17984 (N_17984,N_12537,N_11700);
nand U17985 (N_17985,N_12379,N_13358);
or U17986 (N_17986,N_12327,N_11877);
xnor U17987 (N_17987,N_10894,N_10091);
and U17988 (N_17988,N_13274,N_12195);
nor U17989 (N_17989,N_13895,N_11268);
nand U17990 (N_17990,N_11347,N_11482);
or U17991 (N_17991,N_11275,N_12158);
nor U17992 (N_17992,N_10920,N_12681);
nand U17993 (N_17993,N_14982,N_10828);
and U17994 (N_17994,N_14395,N_11115);
nand U17995 (N_17995,N_14771,N_13677);
xnor U17996 (N_17996,N_10180,N_14558);
and U17997 (N_17997,N_14601,N_11447);
or U17998 (N_17998,N_13175,N_12260);
or U17999 (N_17999,N_10356,N_14203);
nand U18000 (N_18000,N_12526,N_12159);
nand U18001 (N_18001,N_10107,N_14415);
and U18002 (N_18002,N_10679,N_13425);
nand U18003 (N_18003,N_12780,N_13500);
xnor U18004 (N_18004,N_11332,N_12722);
nor U18005 (N_18005,N_12399,N_11971);
nor U18006 (N_18006,N_10299,N_10574);
nor U18007 (N_18007,N_14493,N_14092);
and U18008 (N_18008,N_11472,N_11845);
nand U18009 (N_18009,N_10541,N_12772);
nor U18010 (N_18010,N_11210,N_11070);
nor U18011 (N_18011,N_14650,N_11553);
nor U18012 (N_18012,N_14070,N_12772);
xnor U18013 (N_18013,N_10367,N_13766);
or U18014 (N_18014,N_10337,N_14519);
nand U18015 (N_18015,N_14253,N_12003);
or U18016 (N_18016,N_14817,N_10788);
and U18017 (N_18017,N_10221,N_11715);
and U18018 (N_18018,N_11201,N_14149);
xor U18019 (N_18019,N_11502,N_12554);
nor U18020 (N_18020,N_11412,N_13486);
nor U18021 (N_18021,N_14893,N_14010);
xor U18022 (N_18022,N_14082,N_14153);
xnor U18023 (N_18023,N_10176,N_13088);
nand U18024 (N_18024,N_10557,N_11352);
or U18025 (N_18025,N_12018,N_14644);
nand U18026 (N_18026,N_11241,N_11904);
or U18027 (N_18027,N_11085,N_12527);
or U18028 (N_18028,N_13701,N_10406);
and U18029 (N_18029,N_10868,N_10495);
nand U18030 (N_18030,N_14092,N_13007);
nand U18031 (N_18031,N_10271,N_11271);
and U18032 (N_18032,N_14982,N_10164);
or U18033 (N_18033,N_13997,N_14821);
nor U18034 (N_18034,N_10352,N_10618);
nor U18035 (N_18035,N_13354,N_14267);
or U18036 (N_18036,N_12235,N_10782);
or U18037 (N_18037,N_11713,N_11747);
nor U18038 (N_18038,N_10508,N_10366);
nor U18039 (N_18039,N_12551,N_13482);
and U18040 (N_18040,N_10134,N_11613);
or U18041 (N_18041,N_14604,N_14780);
nand U18042 (N_18042,N_13080,N_13525);
nand U18043 (N_18043,N_13603,N_11698);
nor U18044 (N_18044,N_13874,N_10859);
and U18045 (N_18045,N_12578,N_12420);
or U18046 (N_18046,N_13341,N_13904);
nand U18047 (N_18047,N_13717,N_14923);
and U18048 (N_18048,N_10476,N_12328);
nor U18049 (N_18049,N_12223,N_12315);
and U18050 (N_18050,N_10449,N_12729);
or U18051 (N_18051,N_10595,N_13785);
and U18052 (N_18052,N_10176,N_14923);
xnor U18053 (N_18053,N_11849,N_11562);
xor U18054 (N_18054,N_14584,N_14909);
or U18055 (N_18055,N_10924,N_10427);
nor U18056 (N_18056,N_13328,N_13000);
xnor U18057 (N_18057,N_13435,N_13828);
nand U18058 (N_18058,N_14212,N_14437);
nor U18059 (N_18059,N_14039,N_10283);
nand U18060 (N_18060,N_10720,N_14797);
nor U18061 (N_18061,N_13400,N_13840);
and U18062 (N_18062,N_11187,N_11759);
nand U18063 (N_18063,N_12424,N_12006);
nor U18064 (N_18064,N_12390,N_13999);
nor U18065 (N_18065,N_12482,N_11353);
nand U18066 (N_18066,N_12153,N_10479);
nand U18067 (N_18067,N_14137,N_10905);
and U18068 (N_18068,N_12752,N_10237);
nand U18069 (N_18069,N_14311,N_11499);
or U18070 (N_18070,N_13009,N_14582);
nor U18071 (N_18071,N_10206,N_11660);
nand U18072 (N_18072,N_12511,N_14766);
nand U18073 (N_18073,N_11177,N_14088);
nand U18074 (N_18074,N_14594,N_14690);
nor U18075 (N_18075,N_13501,N_14079);
xor U18076 (N_18076,N_13948,N_10448);
nand U18077 (N_18077,N_14685,N_12697);
nand U18078 (N_18078,N_12971,N_13438);
nand U18079 (N_18079,N_11865,N_14747);
xor U18080 (N_18080,N_11869,N_13311);
xor U18081 (N_18081,N_10891,N_11856);
and U18082 (N_18082,N_11682,N_10424);
or U18083 (N_18083,N_13870,N_10939);
or U18084 (N_18084,N_11309,N_11420);
nor U18085 (N_18085,N_14174,N_12529);
nand U18086 (N_18086,N_11901,N_11895);
and U18087 (N_18087,N_13923,N_14928);
nor U18088 (N_18088,N_12794,N_12006);
xnor U18089 (N_18089,N_10848,N_10877);
nand U18090 (N_18090,N_12086,N_12272);
or U18091 (N_18091,N_10515,N_11115);
and U18092 (N_18092,N_12061,N_14228);
xor U18093 (N_18093,N_10615,N_11857);
and U18094 (N_18094,N_13446,N_12035);
xor U18095 (N_18095,N_12531,N_11868);
or U18096 (N_18096,N_14203,N_12126);
xor U18097 (N_18097,N_14527,N_13633);
or U18098 (N_18098,N_11229,N_12412);
xnor U18099 (N_18099,N_11807,N_11095);
xor U18100 (N_18100,N_10342,N_12963);
and U18101 (N_18101,N_11967,N_10981);
xor U18102 (N_18102,N_13773,N_11909);
nor U18103 (N_18103,N_13923,N_10500);
or U18104 (N_18104,N_11078,N_11763);
and U18105 (N_18105,N_14571,N_13469);
nand U18106 (N_18106,N_10191,N_14233);
or U18107 (N_18107,N_12250,N_10444);
or U18108 (N_18108,N_11767,N_12272);
xnor U18109 (N_18109,N_12512,N_12262);
xnor U18110 (N_18110,N_12814,N_12996);
or U18111 (N_18111,N_13577,N_11649);
nand U18112 (N_18112,N_14859,N_10190);
or U18113 (N_18113,N_10660,N_12680);
or U18114 (N_18114,N_12913,N_11364);
xnor U18115 (N_18115,N_10228,N_10706);
or U18116 (N_18116,N_10591,N_12849);
xor U18117 (N_18117,N_11499,N_12218);
and U18118 (N_18118,N_11333,N_10375);
or U18119 (N_18119,N_13189,N_11745);
nand U18120 (N_18120,N_14280,N_12641);
or U18121 (N_18121,N_14713,N_12978);
nand U18122 (N_18122,N_11714,N_13203);
nand U18123 (N_18123,N_11274,N_11278);
nor U18124 (N_18124,N_10177,N_12342);
xor U18125 (N_18125,N_14695,N_12950);
or U18126 (N_18126,N_13854,N_10148);
and U18127 (N_18127,N_10621,N_13023);
and U18128 (N_18128,N_11912,N_12595);
nor U18129 (N_18129,N_13151,N_12750);
nor U18130 (N_18130,N_13964,N_14932);
nand U18131 (N_18131,N_10461,N_14132);
nor U18132 (N_18132,N_11575,N_12583);
nor U18133 (N_18133,N_12337,N_14771);
nor U18134 (N_18134,N_13503,N_13297);
and U18135 (N_18135,N_12240,N_10819);
nor U18136 (N_18136,N_13135,N_11650);
nand U18137 (N_18137,N_10535,N_14943);
xor U18138 (N_18138,N_13637,N_13416);
or U18139 (N_18139,N_10366,N_12264);
and U18140 (N_18140,N_14677,N_13647);
or U18141 (N_18141,N_13839,N_13570);
nor U18142 (N_18142,N_10113,N_11892);
and U18143 (N_18143,N_12668,N_11321);
nand U18144 (N_18144,N_10128,N_12302);
nand U18145 (N_18145,N_10985,N_12343);
nand U18146 (N_18146,N_11763,N_10776);
and U18147 (N_18147,N_10894,N_13059);
nor U18148 (N_18148,N_10302,N_12653);
xor U18149 (N_18149,N_14639,N_12708);
and U18150 (N_18150,N_13201,N_13764);
or U18151 (N_18151,N_13873,N_12608);
nand U18152 (N_18152,N_14561,N_13959);
or U18153 (N_18153,N_14199,N_10287);
nand U18154 (N_18154,N_10812,N_14994);
xor U18155 (N_18155,N_13987,N_12662);
and U18156 (N_18156,N_10118,N_13652);
xnor U18157 (N_18157,N_11688,N_12403);
nor U18158 (N_18158,N_13856,N_11754);
nor U18159 (N_18159,N_14301,N_13517);
and U18160 (N_18160,N_12317,N_14924);
or U18161 (N_18161,N_12927,N_10414);
and U18162 (N_18162,N_12843,N_13401);
and U18163 (N_18163,N_10661,N_14329);
and U18164 (N_18164,N_14057,N_10946);
nand U18165 (N_18165,N_13290,N_13257);
nor U18166 (N_18166,N_12800,N_12030);
or U18167 (N_18167,N_14282,N_10178);
and U18168 (N_18168,N_14221,N_14470);
nand U18169 (N_18169,N_12328,N_11713);
nor U18170 (N_18170,N_10350,N_14934);
or U18171 (N_18171,N_12270,N_14413);
nor U18172 (N_18172,N_11572,N_11703);
nor U18173 (N_18173,N_12333,N_12545);
or U18174 (N_18174,N_14014,N_12259);
nand U18175 (N_18175,N_12845,N_12786);
nand U18176 (N_18176,N_10659,N_10270);
nand U18177 (N_18177,N_11646,N_11280);
xnor U18178 (N_18178,N_14075,N_14457);
xor U18179 (N_18179,N_12561,N_10165);
and U18180 (N_18180,N_11245,N_12937);
or U18181 (N_18181,N_13601,N_14587);
and U18182 (N_18182,N_10450,N_11886);
and U18183 (N_18183,N_10376,N_11678);
or U18184 (N_18184,N_13936,N_11767);
nand U18185 (N_18185,N_13042,N_11864);
and U18186 (N_18186,N_14217,N_10116);
nor U18187 (N_18187,N_10290,N_10789);
and U18188 (N_18188,N_10189,N_10413);
and U18189 (N_18189,N_12423,N_14828);
xnor U18190 (N_18190,N_14868,N_13320);
or U18191 (N_18191,N_12716,N_10485);
nor U18192 (N_18192,N_11575,N_14197);
nand U18193 (N_18193,N_13177,N_10067);
and U18194 (N_18194,N_13269,N_10369);
or U18195 (N_18195,N_12583,N_11057);
and U18196 (N_18196,N_14986,N_12544);
nor U18197 (N_18197,N_11901,N_10264);
xor U18198 (N_18198,N_10015,N_13649);
or U18199 (N_18199,N_10490,N_13857);
nand U18200 (N_18200,N_12011,N_12937);
nor U18201 (N_18201,N_13152,N_11270);
xor U18202 (N_18202,N_11293,N_14647);
nor U18203 (N_18203,N_11441,N_10850);
nand U18204 (N_18204,N_12781,N_10105);
xor U18205 (N_18205,N_14740,N_12152);
nor U18206 (N_18206,N_14143,N_13166);
or U18207 (N_18207,N_13251,N_10842);
nand U18208 (N_18208,N_13976,N_10657);
or U18209 (N_18209,N_14351,N_12927);
or U18210 (N_18210,N_12980,N_11812);
nand U18211 (N_18211,N_14255,N_12000);
xor U18212 (N_18212,N_14984,N_14480);
or U18213 (N_18213,N_11131,N_12803);
nor U18214 (N_18214,N_14924,N_13518);
or U18215 (N_18215,N_14763,N_14999);
and U18216 (N_18216,N_13793,N_13057);
nor U18217 (N_18217,N_12168,N_13912);
and U18218 (N_18218,N_13589,N_11266);
nor U18219 (N_18219,N_14066,N_12355);
and U18220 (N_18220,N_14586,N_10131);
or U18221 (N_18221,N_14156,N_10663);
nand U18222 (N_18222,N_11870,N_10695);
nor U18223 (N_18223,N_13608,N_10521);
nor U18224 (N_18224,N_12589,N_14066);
nor U18225 (N_18225,N_10028,N_14354);
or U18226 (N_18226,N_12039,N_13306);
or U18227 (N_18227,N_13248,N_14694);
nand U18228 (N_18228,N_12210,N_11997);
nor U18229 (N_18229,N_11036,N_14310);
nor U18230 (N_18230,N_14075,N_11838);
xnor U18231 (N_18231,N_14687,N_11687);
xnor U18232 (N_18232,N_14238,N_13698);
nand U18233 (N_18233,N_10496,N_10468);
and U18234 (N_18234,N_10147,N_13576);
nor U18235 (N_18235,N_14000,N_14134);
or U18236 (N_18236,N_14394,N_13024);
and U18237 (N_18237,N_11761,N_10786);
xnor U18238 (N_18238,N_10437,N_12179);
or U18239 (N_18239,N_10324,N_11524);
xnor U18240 (N_18240,N_14614,N_12317);
nand U18241 (N_18241,N_12556,N_10080);
nor U18242 (N_18242,N_10261,N_12179);
nand U18243 (N_18243,N_12659,N_12449);
nand U18244 (N_18244,N_14173,N_11494);
nand U18245 (N_18245,N_12061,N_14130);
or U18246 (N_18246,N_13891,N_13305);
or U18247 (N_18247,N_11214,N_11494);
and U18248 (N_18248,N_10088,N_11497);
nor U18249 (N_18249,N_14757,N_11040);
nand U18250 (N_18250,N_10980,N_14099);
and U18251 (N_18251,N_14788,N_12989);
and U18252 (N_18252,N_11329,N_10632);
xnor U18253 (N_18253,N_12927,N_13517);
nand U18254 (N_18254,N_13895,N_10677);
and U18255 (N_18255,N_14315,N_14833);
nor U18256 (N_18256,N_13301,N_11894);
xnor U18257 (N_18257,N_11705,N_14275);
or U18258 (N_18258,N_14897,N_14113);
nor U18259 (N_18259,N_11553,N_11607);
nand U18260 (N_18260,N_12291,N_12896);
and U18261 (N_18261,N_12181,N_11397);
xor U18262 (N_18262,N_11528,N_10914);
and U18263 (N_18263,N_10955,N_11187);
nand U18264 (N_18264,N_14392,N_11584);
and U18265 (N_18265,N_12607,N_13668);
or U18266 (N_18266,N_11797,N_11291);
nor U18267 (N_18267,N_14045,N_14988);
and U18268 (N_18268,N_13640,N_13262);
and U18269 (N_18269,N_14239,N_14553);
xor U18270 (N_18270,N_10358,N_14021);
or U18271 (N_18271,N_10142,N_14232);
xnor U18272 (N_18272,N_12663,N_10594);
and U18273 (N_18273,N_13586,N_12680);
xor U18274 (N_18274,N_12723,N_14831);
and U18275 (N_18275,N_14710,N_12909);
xor U18276 (N_18276,N_10304,N_13842);
xnor U18277 (N_18277,N_14850,N_12238);
nand U18278 (N_18278,N_11488,N_14210);
xnor U18279 (N_18279,N_12276,N_12046);
nand U18280 (N_18280,N_12311,N_14736);
nand U18281 (N_18281,N_14980,N_14200);
xor U18282 (N_18282,N_14037,N_13361);
nand U18283 (N_18283,N_11310,N_14869);
nand U18284 (N_18284,N_10836,N_10940);
xor U18285 (N_18285,N_11641,N_12918);
or U18286 (N_18286,N_10268,N_14173);
xnor U18287 (N_18287,N_10837,N_10662);
xnor U18288 (N_18288,N_11650,N_14846);
xor U18289 (N_18289,N_11495,N_12818);
xor U18290 (N_18290,N_11403,N_10327);
nor U18291 (N_18291,N_14926,N_14999);
or U18292 (N_18292,N_11362,N_12318);
nor U18293 (N_18293,N_10738,N_13152);
xor U18294 (N_18294,N_12227,N_10159);
or U18295 (N_18295,N_14728,N_11574);
nor U18296 (N_18296,N_10799,N_11305);
nand U18297 (N_18297,N_11038,N_13244);
nand U18298 (N_18298,N_12774,N_10216);
or U18299 (N_18299,N_13018,N_12554);
nor U18300 (N_18300,N_12252,N_11666);
nor U18301 (N_18301,N_14685,N_13974);
and U18302 (N_18302,N_12807,N_12927);
and U18303 (N_18303,N_12177,N_12400);
nand U18304 (N_18304,N_11556,N_13611);
xor U18305 (N_18305,N_12652,N_11534);
nor U18306 (N_18306,N_10736,N_13628);
and U18307 (N_18307,N_10045,N_10777);
nor U18308 (N_18308,N_12642,N_13955);
nor U18309 (N_18309,N_12297,N_14970);
nand U18310 (N_18310,N_11569,N_13593);
or U18311 (N_18311,N_11667,N_10165);
xnor U18312 (N_18312,N_11952,N_13952);
xnor U18313 (N_18313,N_12655,N_12339);
nor U18314 (N_18314,N_14939,N_12355);
and U18315 (N_18315,N_12892,N_11246);
or U18316 (N_18316,N_12477,N_10579);
xnor U18317 (N_18317,N_11607,N_12194);
nor U18318 (N_18318,N_13642,N_10963);
nor U18319 (N_18319,N_14529,N_14964);
or U18320 (N_18320,N_14147,N_14929);
or U18321 (N_18321,N_13635,N_11726);
or U18322 (N_18322,N_11487,N_12934);
or U18323 (N_18323,N_13840,N_13489);
nor U18324 (N_18324,N_12441,N_12354);
or U18325 (N_18325,N_12939,N_12012);
and U18326 (N_18326,N_11935,N_10948);
and U18327 (N_18327,N_11467,N_10176);
and U18328 (N_18328,N_11695,N_11972);
xor U18329 (N_18329,N_10926,N_10051);
or U18330 (N_18330,N_10465,N_13698);
xor U18331 (N_18331,N_10408,N_14402);
and U18332 (N_18332,N_10600,N_13762);
nand U18333 (N_18333,N_14768,N_13050);
and U18334 (N_18334,N_10944,N_13400);
or U18335 (N_18335,N_11179,N_12943);
or U18336 (N_18336,N_11066,N_14815);
xnor U18337 (N_18337,N_10069,N_11544);
or U18338 (N_18338,N_10802,N_12467);
nand U18339 (N_18339,N_11410,N_13261);
xor U18340 (N_18340,N_13941,N_14096);
xnor U18341 (N_18341,N_12144,N_14049);
nand U18342 (N_18342,N_12871,N_12450);
nand U18343 (N_18343,N_10519,N_11639);
nand U18344 (N_18344,N_10985,N_14684);
and U18345 (N_18345,N_12427,N_13345);
nor U18346 (N_18346,N_12206,N_11601);
or U18347 (N_18347,N_13357,N_11222);
xor U18348 (N_18348,N_12067,N_13022);
xnor U18349 (N_18349,N_11948,N_14180);
and U18350 (N_18350,N_11325,N_14178);
or U18351 (N_18351,N_14434,N_11200);
or U18352 (N_18352,N_10551,N_14768);
nor U18353 (N_18353,N_10313,N_10478);
nand U18354 (N_18354,N_14523,N_10161);
or U18355 (N_18355,N_10988,N_10559);
nand U18356 (N_18356,N_12395,N_13854);
nor U18357 (N_18357,N_11801,N_10317);
or U18358 (N_18358,N_10433,N_12578);
xnor U18359 (N_18359,N_14247,N_13526);
xnor U18360 (N_18360,N_14484,N_11658);
nor U18361 (N_18361,N_13637,N_12054);
and U18362 (N_18362,N_10348,N_10983);
or U18363 (N_18363,N_10190,N_10749);
xnor U18364 (N_18364,N_10069,N_13305);
and U18365 (N_18365,N_14312,N_13641);
or U18366 (N_18366,N_14515,N_12971);
xnor U18367 (N_18367,N_11268,N_10837);
or U18368 (N_18368,N_11338,N_13262);
or U18369 (N_18369,N_13067,N_13326);
nor U18370 (N_18370,N_13774,N_12296);
nand U18371 (N_18371,N_10443,N_10710);
xnor U18372 (N_18372,N_14190,N_10903);
nand U18373 (N_18373,N_11033,N_11626);
or U18374 (N_18374,N_14246,N_14471);
nand U18375 (N_18375,N_11671,N_14987);
xnor U18376 (N_18376,N_12253,N_13200);
nand U18377 (N_18377,N_11131,N_10140);
and U18378 (N_18378,N_13177,N_14837);
nand U18379 (N_18379,N_11808,N_13066);
and U18380 (N_18380,N_11151,N_11679);
xor U18381 (N_18381,N_11541,N_13533);
or U18382 (N_18382,N_14491,N_14354);
or U18383 (N_18383,N_10803,N_10264);
or U18384 (N_18384,N_12419,N_10213);
nand U18385 (N_18385,N_13690,N_10954);
or U18386 (N_18386,N_12914,N_10325);
nor U18387 (N_18387,N_10042,N_10588);
nand U18388 (N_18388,N_11187,N_12149);
nor U18389 (N_18389,N_13432,N_11685);
and U18390 (N_18390,N_14131,N_11471);
xor U18391 (N_18391,N_10952,N_14976);
xnor U18392 (N_18392,N_11215,N_12677);
xor U18393 (N_18393,N_12127,N_13233);
nand U18394 (N_18394,N_11791,N_13869);
nor U18395 (N_18395,N_14670,N_10204);
xor U18396 (N_18396,N_13821,N_14443);
or U18397 (N_18397,N_10088,N_12082);
xor U18398 (N_18398,N_12155,N_14701);
xnor U18399 (N_18399,N_13837,N_13898);
xnor U18400 (N_18400,N_11048,N_11368);
xor U18401 (N_18401,N_12761,N_12748);
and U18402 (N_18402,N_13789,N_14582);
or U18403 (N_18403,N_12328,N_11257);
xor U18404 (N_18404,N_10304,N_12327);
nand U18405 (N_18405,N_11047,N_12972);
xor U18406 (N_18406,N_10582,N_14191);
nor U18407 (N_18407,N_14028,N_11181);
nor U18408 (N_18408,N_10244,N_10790);
or U18409 (N_18409,N_14582,N_13617);
xnor U18410 (N_18410,N_10342,N_10492);
nand U18411 (N_18411,N_12564,N_14637);
xnor U18412 (N_18412,N_14798,N_10673);
nor U18413 (N_18413,N_11768,N_11725);
nor U18414 (N_18414,N_14960,N_12292);
or U18415 (N_18415,N_11486,N_11317);
nand U18416 (N_18416,N_13494,N_10658);
xnor U18417 (N_18417,N_12391,N_11566);
xor U18418 (N_18418,N_10210,N_10177);
and U18419 (N_18419,N_12058,N_11750);
nor U18420 (N_18420,N_11185,N_14034);
or U18421 (N_18421,N_12742,N_11498);
nand U18422 (N_18422,N_12419,N_11999);
xor U18423 (N_18423,N_14158,N_11345);
xor U18424 (N_18424,N_11017,N_13021);
or U18425 (N_18425,N_14884,N_11041);
nor U18426 (N_18426,N_12099,N_14568);
nand U18427 (N_18427,N_13944,N_10631);
xnor U18428 (N_18428,N_11200,N_14600);
or U18429 (N_18429,N_10243,N_13774);
or U18430 (N_18430,N_11637,N_14270);
or U18431 (N_18431,N_13992,N_14938);
and U18432 (N_18432,N_12625,N_14363);
nor U18433 (N_18433,N_12263,N_12253);
or U18434 (N_18434,N_14131,N_12681);
nand U18435 (N_18435,N_13239,N_11541);
nand U18436 (N_18436,N_12323,N_10067);
or U18437 (N_18437,N_12359,N_11090);
nand U18438 (N_18438,N_13783,N_14613);
nor U18439 (N_18439,N_13154,N_13166);
nor U18440 (N_18440,N_11141,N_12941);
nor U18441 (N_18441,N_12221,N_10465);
or U18442 (N_18442,N_11993,N_11193);
or U18443 (N_18443,N_14952,N_12798);
or U18444 (N_18444,N_11822,N_14206);
or U18445 (N_18445,N_14570,N_12674);
nand U18446 (N_18446,N_13111,N_13244);
or U18447 (N_18447,N_13090,N_12122);
or U18448 (N_18448,N_12620,N_12060);
xor U18449 (N_18449,N_10064,N_13179);
and U18450 (N_18450,N_12286,N_12244);
xor U18451 (N_18451,N_11447,N_14096);
xnor U18452 (N_18452,N_13025,N_12123);
nand U18453 (N_18453,N_13661,N_12669);
and U18454 (N_18454,N_12591,N_12439);
or U18455 (N_18455,N_12243,N_13198);
nor U18456 (N_18456,N_14934,N_10825);
nand U18457 (N_18457,N_10567,N_14307);
and U18458 (N_18458,N_10608,N_14825);
nor U18459 (N_18459,N_14708,N_13357);
nand U18460 (N_18460,N_14498,N_13356);
xor U18461 (N_18461,N_11311,N_11959);
xor U18462 (N_18462,N_14692,N_10765);
and U18463 (N_18463,N_11090,N_12850);
xor U18464 (N_18464,N_11524,N_12789);
nand U18465 (N_18465,N_11604,N_11561);
and U18466 (N_18466,N_10574,N_10931);
or U18467 (N_18467,N_11380,N_11566);
and U18468 (N_18468,N_14812,N_10159);
and U18469 (N_18469,N_12396,N_12427);
or U18470 (N_18470,N_13818,N_14450);
and U18471 (N_18471,N_14032,N_12131);
or U18472 (N_18472,N_13099,N_10977);
xnor U18473 (N_18473,N_13904,N_10941);
and U18474 (N_18474,N_13659,N_11204);
nand U18475 (N_18475,N_14221,N_14870);
xnor U18476 (N_18476,N_10442,N_13568);
and U18477 (N_18477,N_11602,N_13723);
nand U18478 (N_18478,N_10276,N_14688);
or U18479 (N_18479,N_11525,N_14874);
nor U18480 (N_18480,N_12233,N_10180);
xor U18481 (N_18481,N_12342,N_10932);
nand U18482 (N_18482,N_13970,N_12915);
and U18483 (N_18483,N_10029,N_13223);
and U18484 (N_18484,N_11838,N_12780);
or U18485 (N_18485,N_13607,N_13038);
nand U18486 (N_18486,N_11463,N_14079);
and U18487 (N_18487,N_14790,N_11710);
or U18488 (N_18488,N_10633,N_11162);
xor U18489 (N_18489,N_10937,N_14624);
nor U18490 (N_18490,N_10219,N_14666);
or U18491 (N_18491,N_13606,N_13051);
xnor U18492 (N_18492,N_10227,N_14696);
nor U18493 (N_18493,N_12537,N_10311);
nor U18494 (N_18494,N_14258,N_13633);
nand U18495 (N_18495,N_10498,N_11446);
and U18496 (N_18496,N_10579,N_11933);
or U18497 (N_18497,N_12816,N_13351);
nand U18498 (N_18498,N_13251,N_10712);
nor U18499 (N_18499,N_13835,N_10143);
and U18500 (N_18500,N_11907,N_14345);
or U18501 (N_18501,N_12983,N_10221);
nand U18502 (N_18502,N_11223,N_11831);
and U18503 (N_18503,N_11174,N_14170);
nand U18504 (N_18504,N_11507,N_11474);
nand U18505 (N_18505,N_10301,N_11088);
and U18506 (N_18506,N_13762,N_11598);
nand U18507 (N_18507,N_11927,N_10372);
and U18508 (N_18508,N_10446,N_12295);
or U18509 (N_18509,N_13252,N_13978);
nor U18510 (N_18510,N_12590,N_13395);
xor U18511 (N_18511,N_10179,N_11921);
and U18512 (N_18512,N_14279,N_10621);
xor U18513 (N_18513,N_10957,N_10284);
and U18514 (N_18514,N_12926,N_14123);
xor U18515 (N_18515,N_13076,N_12753);
nand U18516 (N_18516,N_11377,N_12746);
nand U18517 (N_18517,N_11005,N_12032);
and U18518 (N_18518,N_11140,N_10377);
and U18519 (N_18519,N_10444,N_13540);
xor U18520 (N_18520,N_14929,N_11793);
nor U18521 (N_18521,N_14223,N_13377);
xor U18522 (N_18522,N_13402,N_13751);
and U18523 (N_18523,N_13616,N_13427);
nor U18524 (N_18524,N_13704,N_10402);
or U18525 (N_18525,N_11127,N_12582);
or U18526 (N_18526,N_12918,N_13605);
nand U18527 (N_18527,N_14040,N_13172);
xnor U18528 (N_18528,N_11584,N_12415);
and U18529 (N_18529,N_10217,N_12712);
nand U18530 (N_18530,N_13780,N_14272);
xnor U18531 (N_18531,N_12557,N_14798);
and U18532 (N_18532,N_12915,N_13280);
nor U18533 (N_18533,N_12108,N_11843);
or U18534 (N_18534,N_12712,N_11392);
nor U18535 (N_18535,N_10772,N_11420);
nand U18536 (N_18536,N_12461,N_10299);
and U18537 (N_18537,N_14051,N_12571);
nand U18538 (N_18538,N_11383,N_12551);
or U18539 (N_18539,N_12593,N_10043);
xor U18540 (N_18540,N_14268,N_10772);
and U18541 (N_18541,N_14752,N_11640);
or U18542 (N_18542,N_14825,N_13071);
nor U18543 (N_18543,N_13312,N_14802);
xnor U18544 (N_18544,N_14802,N_10641);
nor U18545 (N_18545,N_13334,N_12384);
and U18546 (N_18546,N_13376,N_14022);
nand U18547 (N_18547,N_14336,N_11482);
xor U18548 (N_18548,N_13542,N_13796);
or U18549 (N_18549,N_10987,N_12209);
or U18550 (N_18550,N_12740,N_13747);
nor U18551 (N_18551,N_13091,N_13407);
nand U18552 (N_18552,N_12811,N_14712);
nor U18553 (N_18553,N_13833,N_12561);
or U18554 (N_18554,N_13324,N_11116);
and U18555 (N_18555,N_13378,N_10156);
or U18556 (N_18556,N_14729,N_12294);
nand U18557 (N_18557,N_12691,N_10064);
nor U18558 (N_18558,N_11341,N_11943);
and U18559 (N_18559,N_12666,N_11349);
and U18560 (N_18560,N_14973,N_11879);
nand U18561 (N_18561,N_13921,N_14273);
nor U18562 (N_18562,N_12490,N_13148);
nor U18563 (N_18563,N_10196,N_10168);
nor U18564 (N_18564,N_12134,N_11194);
and U18565 (N_18565,N_10327,N_11586);
nand U18566 (N_18566,N_11886,N_14394);
xnor U18567 (N_18567,N_13179,N_13465);
xor U18568 (N_18568,N_12717,N_14679);
nor U18569 (N_18569,N_13784,N_13004);
nor U18570 (N_18570,N_12618,N_14138);
nand U18571 (N_18571,N_14350,N_12597);
or U18572 (N_18572,N_11258,N_13363);
nor U18573 (N_18573,N_13401,N_11706);
and U18574 (N_18574,N_14689,N_10392);
xnor U18575 (N_18575,N_12342,N_13274);
nor U18576 (N_18576,N_14732,N_11047);
nand U18577 (N_18577,N_13235,N_13774);
or U18578 (N_18578,N_13634,N_12834);
nand U18579 (N_18579,N_13442,N_12024);
xor U18580 (N_18580,N_13682,N_14120);
or U18581 (N_18581,N_11410,N_14062);
xnor U18582 (N_18582,N_11913,N_11062);
and U18583 (N_18583,N_13721,N_14639);
nand U18584 (N_18584,N_13924,N_14341);
nor U18585 (N_18585,N_13920,N_11281);
xor U18586 (N_18586,N_12293,N_10295);
xor U18587 (N_18587,N_10041,N_11879);
nand U18588 (N_18588,N_11209,N_10366);
nor U18589 (N_18589,N_14653,N_13430);
and U18590 (N_18590,N_12122,N_10231);
and U18591 (N_18591,N_11060,N_14468);
xnor U18592 (N_18592,N_14041,N_14201);
nor U18593 (N_18593,N_13284,N_13904);
nand U18594 (N_18594,N_12352,N_13266);
and U18595 (N_18595,N_12023,N_11697);
nand U18596 (N_18596,N_13056,N_12362);
and U18597 (N_18597,N_10826,N_12065);
and U18598 (N_18598,N_13823,N_10407);
and U18599 (N_18599,N_11301,N_10172);
or U18600 (N_18600,N_14321,N_13438);
xor U18601 (N_18601,N_14116,N_13348);
nor U18602 (N_18602,N_14144,N_13059);
nor U18603 (N_18603,N_14190,N_13791);
or U18604 (N_18604,N_10598,N_10044);
nor U18605 (N_18605,N_11120,N_10437);
and U18606 (N_18606,N_11596,N_12286);
xnor U18607 (N_18607,N_10364,N_14417);
nand U18608 (N_18608,N_13817,N_13806);
or U18609 (N_18609,N_10507,N_10706);
xor U18610 (N_18610,N_10978,N_13880);
and U18611 (N_18611,N_13796,N_11572);
xnor U18612 (N_18612,N_12354,N_10615);
xor U18613 (N_18613,N_12063,N_10998);
and U18614 (N_18614,N_14986,N_10917);
nor U18615 (N_18615,N_10150,N_10468);
nor U18616 (N_18616,N_11287,N_14791);
or U18617 (N_18617,N_10539,N_11988);
nand U18618 (N_18618,N_12702,N_14557);
xor U18619 (N_18619,N_13899,N_12866);
and U18620 (N_18620,N_13478,N_14789);
or U18621 (N_18621,N_10814,N_14128);
and U18622 (N_18622,N_14838,N_11871);
nor U18623 (N_18623,N_14315,N_12119);
and U18624 (N_18624,N_13777,N_12435);
or U18625 (N_18625,N_10515,N_14274);
nand U18626 (N_18626,N_14803,N_13499);
xnor U18627 (N_18627,N_10118,N_13516);
nand U18628 (N_18628,N_13128,N_11397);
nor U18629 (N_18629,N_10662,N_12688);
nor U18630 (N_18630,N_12368,N_10934);
and U18631 (N_18631,N_10638,N_13260);
nand U18632 (N_18632,N_10607,N_14745);
or U18633 (N_18633,N_13334,N_14427);
or U18634 (N_18634,N_13290,N_12052);
nand U18635 (N_18635,N_12642,N_11827);
xor U18636 (N_18636,N_12147,N_14033);
and U18637 (N_18637,N_10120,N_12205);
xnor U18638 (N_18638,N_13134,N_14451);
nor U18639 (N_18639,N_13103,N_12455);
nor U18640 (N_18640,N_10239,N_12644);
xor U18641 (N_18641,N_11335,N_14425);
or U18642 (N_18642,N_12667,N_10073);
nor U18643 (N_18643,N_12220,N_12519);
xnor U18644 (N_18644,N_12927,N_10082);
nand U18645 (N_18645,N_11181,N_13198);
xnor U18646 (N_18646,N_14421,N_14311);
nand U18647 (N_18647,N_14129,N_10025);
nor U18648 (N_18648,N_10142,N_10824);
nand U18649 (N_18649,N_14360,N_14594);
xnor U18650 (N_18650,N_13352,N_10492);
xnor U18651 (N_18651,N_10491,N_14346);
and U18652 (N_18652,N_10018,N_10402);
nor U18653 (N_18653,N_11334,N_10562);
xnor U18654 (N_18654,N_10781,N_11834);
xor U18655 (N_18655,N_14069,N_11544);
or U18656 (N_18656,N_10852,N_12415);
or U18657 (N_18657,N_12581,N_10781);
or U18658 (N_18658,N_11586,N_13788);
or U18659 (N_18659,N_11039,N_13923);
nor U18660 (N_18660,N_14984,N_13002);
nand U18661 (N_18661,N_10804,N_11265);
and U18662 (N_18662,N_13766,N_11472);
nand U18663 (N_18663,N_10415,N_14655);
and U18664 (N_18664,N_13775,N_11349);
nand U18665 (N_18665,N_11110,N_13254);
and U18666 (N_18666,N_14802,N_13573);
and U18667 (N_18667,N_14298,N_11201);
or U18668 (N_18668,N_12344,N_11429);
xnor U18669 (N_18669,N_11214,N_12098);
xor U18670 (N_18670,N_13706,N_13365);
and U18671 (N_18671,N_14950,N_13293);
nor U18672 (N_18672,N_12088,N_13964);
and U18673 (N_18673,N_12980,N_12774);
nor U18674 (N_18674,N_12278,N_10608);
xor U18675 (N_18675,N_13656,N_11056);
xor U18676 (N_18676,N_14033,N_12500);
and U18677 (N_18677,N_13179,N_14637);
and U18678 (N_18678,N_10946,N_11384);
nor U18679 (N_18679,N_10309,N_14472);
nand U18680 (N_18680,N_11748,N_14919);
nor U18681 (N_18681,N_10536,N_12901);
nor U18682 (N_18682,N_11063,N_10836);
xor U18683 (N_18683,N_12034,N_13430);
xor U18684 (N_18684,N_13676,N_13257);
nor U18685 (N_18685,N_13031,N_12451);
nand U18686 (N_18686,N_11707,N_12609);
nor U18687 (N_18687,N_13278,N_10772);
or U18688 (N_18688,N_12406,N_12880);
or U18689 (N_18689,N_12177,N_10862);
or U18690 (N_18690,N_10355,N_14180);
xor U18691 (N_18691,N_11848,N_13352);
nand U18692 (N_18692,N_13865,N_10655);
and U18693 (N_18693,N_10082,N_10821);
nand U18694 (N_18694,N_14486,N_13869);
or U18695 (N_18695,N_11382,N_13135);
or U18696 (N_18696,N_13850,N_12644);
nor U18697 (N_18697,N_11008,N_11988);
xnor U18698 (N_18698,N_12836,N_12360);
nand U18699 (N_18699,N_11228,N_11818);
nand U18700 (N_18700,N_11580,N_14879);
or U18701 (N_18701,N_11034,N_14944);
nor U18702 (N_18702,N_11068,N_13759);
and U18703 (N_18703,N_14379,N_13415);
nor U18704 (N_18704,N_14688,N_10920);
and U18705 (N_18705,N_13413,N_12712);
or U18706 (N_18706,N_11686,N_13232);
nand U18707 (N_18707,N_12600,N_12387);
nor U18708 (N_18708,N_14593,N_13040);
and U18709 (N_18709,N_14799,N_11502);
xnor U18710 (N_18710,N_11204,N_10478);
xor U18711 (N_18711,N_14142,N_11647);
and U18712 (N_18712,N_10833,N_11254);
nor U18713 (N_18713,N_12584,N_13999);
nand U18714 (N_18714,N_14910,N_12525);
xnor U18715 (N_18715,N_13031,N_11993);
or U18716 (N_18716,N_10347,N_14152);
or U18717 (N_18717,N_14671,N_10905);
and U18718 (N_18718,N_12479,N_10155);
nor U18719 (N_18719,N_10651,N_11986);
xor U18720 (N_18720,N_11611,N_11194);
or U18721 (N_18721,N_14506,N_11640);
nor U18722 (N_18722,N_10235,N_10407);
xor U18723 (N_18723,N_13195,N_13825);
xnor U18724 (N_18724,N_14657,N_14305);
nor U18725 (N_18725,N_14584,N_14520);
nand U18726 (N_18726,N_11948,N_13231);
nor U18727 (N_18727,N_10362,N_11796);
or U18728 (N_18728,N_11988,N_12190);
xnor U18729 (N_18729,N_13495,N_11953);
xnor U18730 (N_18730,N_13755,N_12953);
or U18731 (N_18731,N_13032,N_12026);
xor U18732 (N_18732,N_12502,N_13227);
nand U18733 (N_18733,N_11639,N_12547);
and U18734 (N_18734,N_11009,N_10022);
nand U18735 (N_18735,N_14895,N_10757);
nor U18736 (N_18736,N_12954,N_12906);
and U18737 (N_18737,N_14438,N_14212);
or U18738 (N_18738,N_14805,N_14730);
nor U18739 (N_18739,N_13551,N_13558);
nand U18740 (N_18740,N_11710,N_14287);
nor U18741 (N_18741,N_12729,N_11167);
and U18742 (N_18742,N_13006,N_10067);
or U18743 (N_18743,N_10000,N_14956);
or U18744 (N_18744,N_11723,N_12453);
nand U18745 (N_18745,N_14611,N_10967);
and U18746 (N_18746,N_11831,N_12259);
nor U18747 (N_18747,N_12295,N_12434);
nor U18748 (N_18748,N_14230,N_13251);
xnor U18749 (N_18749,N_12707,N_10259);
nand U18750 (N_18750,N_10312,N_13330);
or U18751 (N_18751,N_12237,N_12366);
nor U18752 (N_18752,N_12043,N_10638);
nand U18753 (N_18753,N_10411,N_10461);
nor U18754 (N_18754,N_12287,N_14678);
nand U18755 (N_18755,N_13008,N_11958);
xnor U18756 (N_18756,N_12036,N_14496);
xnor U18757 (N_18757,N_10070,N_13858);
and U18758 (N_18758,N_14998,N_11690);
or U18759 (N_18759,N_12652,N_12278);
nor U18760 (N_18760,N_10972,N_10824);
and U18761 (N_18761,N_14086,N_12713);
nand U18762 (N_18762,N_11787,N_13158);
nor U18763 (N_18763,N_12195,N_12410);
nand U18764 (N_18764,N_14050,N_10472);
xnor U18765 (N_18765,N_14287,N_14188);
nand U18766 (N_18766,N_10665,N_11411);
nor U18767 (N_18767,N_10675,N_10975);
xnor U18768 (N_18768,N_11461,N_11183);
nand U18769 (N_18769,N_11513,N_11330);
nand U18770 (N_18770,N_12140,N_11211);
or U18771 (N_18771,N_11084,N_13164);
nand U18772 (N_18772,N_12116,N_14644);
nand U18773 (N_18773,N_13670,N_10949);
xnor U18774 (N_18774,N_14050,N_14877);
nor U18775 (N_18775,N_10671,N_14140);
and U18776 (N_18776,N_10830,N_13693);
or U18777 (N_18777,N_13412,N_12705);
and U18778 (N_18778,N_14583,N_10426);
nor U18779 (N_18779,N_10209,N_13898);
and U18780 (N_18780,N_13753,N_12693);
and U18781 (N_18781,N_13747,N_14053);
nor U18782 (N_18782,N_13391,N_11068);
nor U18783 (N_18783,N_10145,N_14464);
or U18784 (N_18784,N_13701,N_13952);
or U18785 (N_18785,N_14409,N_10766);
xnor U18786 (N_18786,N_12798,N_13169);
or U18787 (N_18787,N_13971,N_13894);
nor U18788 (N_18788,N_13902,N_13990);
or U18789 (N_18789,N_12397,N_14046);
nor U18790 (N_18790,N_10618,N_13218);
nand U18791 (N_18791,N_12953,N_10332);
nor U18792 (N_18792,N_12448,N_13931);
or U18793 (N_18793,N_11816,N_14457);
or U18794 (N_18794,N_12183,N_10349);
and U18795 (N_18795,N_13197,N_11713);
and U18796 (N_18796,N_14448,N_14537);
nor U18797 (N_18797,N_14755,N_11688);
nand U18798 (N_18798,N_14791,N_12129);
and U18799 (N_18799,N_13777,N_12627);
xnor U18800 (N_18800,N_12854,N_13272);
nand U18801 (N_18801,N_13181,N_13432);
or U18802 (N_18802,N_10058,N_12293);
and U18803 (N_18803,N_12830,N_11467);
xor U18804 (N_18804,N_10963,N_12482);
nor U18805 (N_18805,N_13193,N_10936);
and U18806 (N_18806,N_13198,N_12257);
nand U18807 (N_18807,N_10485,N_10484);
or U18808 (N_18808,N_13151,N_12872);
or U18809 (N_18809,N_14176,N_10336);
or U18810 (N_18810,N_12873,N_12052);
xor U18811 (N_18811,N_12728,N_11680);
nor U18812 (N_18812,N_12093,N_10018);
and U18813 (N_18813,N_11249,N_11891);
or U18814 (N_18814,N_12761,N_10659);
xnor U18815 (N_18815,N_12146,N_14661);
nor U18816 (N_18816,N_10904,N_12754);
or U18817 (N_18817,N_11109,N_11616);
or U18818 (N_18818,N_14474,N_10589);
nor U18819 (N_18819,N_12803,N_11514);
and U18820 (N_18820,N_13328,N_11843);
nor U18821 (N_18821,N_11717,N_13166);
or U18822 (N_18822,N_13855,N_10916);
nand U18823 (N_18823,N_14002,N_13110);
or U18824 (N_18824,N_14361,N_11377);
and U18825 (N_18825,N_10471,N_12667);
nor U18826 (N_18826,N_14696,N_14568);
nand U18827 (N_18827,N_13931,N_12572);
and U18828 (N_18828,N_13403,N_10343);
xnor U18829 (N_18829,N_11105,N_12625);
and U18830 (N_18830,N_13713,N_11595);
xnor U18831 (N_18831,N_11550,N_10326);
nand U18832 (N_18832,N_12165,N_12701);
or U18833 (N_18833,N_10824,N_13005);
or U18834 (N_18834,N_10324,N_13014);
nor U18835 (N_18835,N_11067,N_10094);
or U18836 (N_18836,N_12409,N_10267);
or U18837 (N_18837,N_10924,N_13835);
nor U18838 (N_18838,N_13074,N_10982);
xor U18839 (N_18839,N_14792,N_14986);
xnor U18840 (N_18840,N_12147,N_11658);
xnor U18841 (N_18841,N_12251,N_12598);
or U18842 (N_18842,N_10979,N_12131);
xor U18843 (N_18843,N_12519,N_14677);
xor U18844 (N_18844,N_11168,N_11485);
nand U18845 (N_18845,N_12768,N_11472);
xnor U18846 (N_18846,N_14655,N_10257);
and U18847 (N_18847,N_10642,N_14290);
nor U18848 (N_18848,N_10093,N_12473);
nor U18849 (N_18849,N_11671,N_11212);
nand U18850 (N_18850,N_12072,N_14872);
xor U18851 (N_18851,N_13519,N_13752);
nor U18852 (N_18852,N_11936,N_13368);
xor U18853 (N_18853,N_11237,N_10497);
nand U18854 (N_18854,N_11925,N_10529);
nand U18855 (N_18855,N_10906,N_12167);
nor U18856 (N_18856,N_12340,N_12956);
or U18857 (N_18857,N_13046,N_13476);
xnor U18858 (N_18858,N_14955,N_14761);
or U18859 (N_18859,N_12815,N_12038);
nand U18860 (N_18860,N_13689,N_10685);
xnor U18861 (N_18861,N_11853,N_10165);
xor U18862 (N_18862,N_14591,N_12646);
nand U18863 (N_18863,N_10151,N_13255);
xor U18864 (N_18864,N_10688,N_14781);
and U18865 (N_18865,N_11462,N_14784);
or U18866 (N_18866,N_10111,N_13423);
or U18867 (N_18867,N_14141,N_12293);
nor U18868 (N_18868,N_14562,N_11674);
xor U18869 (N_18869,N_10400,N_11354);
nand U18870 (N_18870,N_11936,N_12023);
nor U18871 (N_18871,N_11570,N_14221);
nand U18872 (N_18872,N_14498,N_14669);
nand U18873 (N_18873,N_12529,N_12819);
nor U18874 (N_18874,N_11543,N_12275);
and U18875 (N_18875,N_12822,N_14707);
and U18876 (N_18876,N_14195,N_11916);
or U18877 (N_18877,N_14314,N_12881);
or U18878 (N_18878,N_14961,N_10020);
xnor U18879 (N_18879,N_10875,N_10059);
nor U18880 (N_18880,N_11270,N_14985);
xor U18881 (N_18881,N_14739,N_13122);
or U18882 (N_18882,N_12910,N_12515);
or U18883 (N_18883,N_10705,N_12043);
xor U18884 (N_18884,N_12908,N_12144);
nand U18885 (N_18885,N_10160,N_14145);
nand U18886 (N_18886,N_13422,N_10869);
nor U18887 (N_18887,N_10007,N_13609);
nand U18888 (N_18888,N_11846,N_10274);
nor U18889 (N_18889,N_11876,N_12750);
xnor U18890 (N_18890,N_11359,N_11490);
and U18891 (N_18891,N_13315,N_13931);
nor U18892 (N_18892,N_14380,N_13121);
or U18893 (N_18893,N_11911,N_10260);
xnor U18894 (N_18894,N_12883,N_13812);
or U18895 (N_18895,N_14330,N_10135);
nand U18896 (N_18896,N_13798,N_13037);
nor U18897 (N_18897,N_14559,N_11479);
nor U18898 (N_18898,N_11397,N_11161);
nand U18899 (N_18899,N_12876,N_10328);
and U18900 (N_18900,N_14239,N_14551);
and U18901 (N_18901,N_12151,N_11602);
nor U18902 (N_18902,N_14578,N_10826);
xnor U18903 (N_18903,N_13222,N_14152);
or U18904 (N_18904,N_14180,N_13998);
and U18905 (N_18905,N_11835,N_13360);
nand U18906 (N_18906,N_12743,N_14520);
or U18907 (N_18907,N_13921,N_13177);
and U18908 (N_18908,N_13401,N_12355);
xor U18909 (N_18909,N_10856,N_10877);
and U18910 (N_18910,N_11045,N_11093);
xnor U18911 (N_18911,N_10011,N_14199);
nand U18912 (N_18912,N_10227,N_11360);
or U18913 (N_18913,N_11700,N_14672);
nor U18914 (N_18914,N_14250,N_14420);
xnor U18915 (N_18915,N_14916,N_10294);
or U18916 (N_18916,N_11366,N_13358);
nor U18917 (N_18917,N_10213,N_12641);
and U18918 (N_18918,N_10289,N_10697);
and U18919 (N_18919,N_10865,N_13372);
nand U18920 (N_18920,N_12860,N_12169);
or U18921 (N_18921,N_13373,N_10055);
and U18922 (N_18922,N_14146,N_14483);
nand U18923 (N_18923,N_11433,N_14674);
and U18924 (N_18924,N_12043,N_13035);
xnor U18925 (N_18925,N_13935,N_12870);
xor U18926 (N_18926,N_12537,N_12762);
nand U18927 (N_18927,N_10300,N_10599);
nor U18928 (N_18928,N_13836,N_11746);
nor U18929 (N_18929,N_12935,N_13258);
and U18930 (N_18930,N_13540,N_12341);
nor U18931 (N_18931,N_13048,N_10829);
or U18932 (N_18932,N_14848,N_11422);
xnor U18933 (N_18933,N_12204,N_11573);
or U18934 (N_18934,N_11903,N_13569);
nor U18935 (N_18935,N_12871,N_11756);
xnor U18936 (N_18936,N_10661,N_11619);
xor U18937 (N_18937,N_12370,N_12778);
nor U18938 (N_18938,N_13783,N_11802);
or U18939 (N_18939,N_12204,N_12012);
and U18940 (N_18940,N_14147,N_11412);
xnor U18941 (N_18941,N_10041,N_10072);
nor U18942 (N_18942,N_13157,N_14033);
nand U18943 (N_18943,N_10478,N_14353);
xor U18944 (N_18944,N_14399,N_14468);
nor U18945 (N_18945,N_11641,N_14328);
or U18946 (N_18946,N_10836,N_10910);
nor U18947 (N_18947,N_14072,N_10858);
and U18948 (N_18948,N_14162,N_14183);
or U18949 (N_18949,N_10610,N_11899);
and U18950 (N_18950,N_14958,N_11621);
nor U18951 (N_18951,N_14607,N_11013);
and U18952 (N_18952,N_13846,N_14683);
or U18953 (N_18953,N_13374,N_11976);
and U18954 (N_18954,N_10560,N_11564);
nand U18955 (N_18955,N_12259,N_10585);
nand U18956 (N_18956,N_14560,N_10858);
and U18957 (N_18957,N_14224,N_13908);
nand U18958 (N_18958,N_14717,N_12888);
nor U18959 (N_18959,N_14891,N_14734);
xnor U18960 (N_18960,N_13304,N_14599);
xor U18961 (N_18961,N_10337,N_13146);
nand U18962 (N_18962,N_10820,N_10674);
nand U18963 (N_18963,N_10459,N_11160);
or U18964 (N_18964,N_12613,N_14823);
and U18965 (N_18965,N_10369,N_10193);
xnor U18966 (N_18966,N_12618,N_13755);
and U18967 (N_18967,N_12338,N_12879);
nor U18968 (N_18968,N_14056,N_11739);
and U18969 (N_18969,N_13694,N_14490);
nand U18970 (N_18970,N_13343,N_10321);
xor U18971 (N_18971,N_13881,N_11184);
nand U18972 (N_18972,N_12452,N_14641);
xor U18973 (N_18973,N_13890,N_11460);
xor U18974 (N_18974,N_11374,N_13365);
and U18975 (N_18975,N_12132,N_13968);
nor U18976 (N_18976,N_10921,N_14893);
or U18977 (N_18977,N_14154,N_13599);
and U18978 (N_18978,N_14792,N_14968);
and U18979 (N_18979,N_13857,N_10561);
and U18980 (N_18980,N_10237,N_10148);
xor U18981 (N_18981,N_10601,N_12015);
xnor U18982 (N_18982,N_13759,N_12977);
and U18983 (N_18983,N_13947,N_14129);
and U18984 (N_18984,N_10925,N_13644);
nand U18985 (N_18985,N_12203,N_10814);
xnor U18986 (N_18986,N_11456,N_10892);
and U18987 (N_18987,N_12961,N_10569);
nor U18988 (N_18988,N_10852,N_13677);
xor U18989 (N_18989,N_12519,N_14425);
nor U18990 (N_18990,N_13718,N_11097);
nand U18991 (N_18991,N_10057,N_10564);
nor U18992 (N_18992,N_10351,N_10807);
and U18993 (N_18993,N_11457,N_11720);
nand U18994 (N_18994,N_11619,N_11898);
nor U18995 (N_18995,N_13352,N_10193);
or U18996 (N_18996,N_13706,N_13317);
nor U18997 (N_18997,N_11010,N_14020);
and U18998 (N_18998,N_13488,N_14838);
and U18999 (N_18999,N_12069,N_10130);
or U19000 (N_19000,N_12773,N_12751);
and U19001 (N_19001,N_14106,N_11054);
xor U19002 (N_19002,N_12376,N_13105);
or U19003 (N_19003,N_10796,N_10713);
nand U19004 (N_19004,N_10624,N_13683);
nor U19005 (N_19005,N_12692,N_14164);
and U19006 (N_19006,N_11086,N_12528);
nor U19007 (N_19007,N_12088,N_14803);
xnor U19008 (N_19008,N_10963,N_12191);
and U19009 (N_19009,N_10988,N_14226);
xor U19010 (N_19010,N_13937,N_14787);
xor U19011 (N_19011,N_13548,N_12334);
nor U19012 (N_19012,N_14980,N_11615);
nor U19013 (N_19013,N_11317,N_10805);
and U19014 (N_19014,N_11092,N_12448);
or U19015 (N_19015,N_11556,N_12294);
or U19016 (N_19016,N_12713,N_14471);
nor U19017 (N_19017,N_12875,N_11699);
nor U19018 (N_19018,N_13664,N_13055);
or U19019 (N_19019,N_12586,N_10092);
or U19020 (N_19020,N_12435,N_14000);
nor U19021 (N_19021,N_13700,N_14815);
or U19022 (N_19022,N_11931,N_12188);
nor U19023 (N_19023,N_13198,N_11710);
nand U19024 (N_19024,N_11236,N_10267);
or U19025 (N_19025,N_10657,N_14182);
xnor U19026 (N_19026,N_10917,N_10707);
and U19027 (N_19027,N_14980,N_10757);
nor U19028 (N_19028,N_10166,N_11771);
nor U19029 (N_19029,N_14585,N_11023);
or U19030 (N_19030,N_14920,N_11783);
or U19031 (N_19031,N_10024,N_14359);
and U19032 (N_19032,N_14475,N_12406);
xor U19033 (N_19033,N_11388,N_11371);
nand U19034 (N_19034,N_10211,N_14127);
xor U19035 (N_19035,N_10658,N_11385);
xnor U19036 (N_19036,N_10973,N_13584);
nand U19037 (N_19037,N_10955,N_12609);
xnor U19038 (N_19038,N_12684,N_13507);
or U19039 (N_19039,N_13726,N_13464);
nor U19040 (N_19040,N_12189,N_11183);
xor U19041 (N_19041,N_10389,N_13955);
or U19042 (N_19042,N_12509,N_12668);
or U19043 (N_19043,N_11201,N_11249);
xor U19044 (N_19044,N_11340,N_14242);
and U19045 (N_19045,N_12507,N_13620);
nor U19046 (N_19046,N_10526,N_10170);
or U19047 (N_19047,N_11231,N_11286);
nor U19048 (N_19048,N_14282,N_14648);
nand U19049 (N_19049,N_11539,N_14219);
and U19050 (N_19050,N_13727,N_10425);
nor U19051 (N_19051,N_11016,N_12321);
nand U19052 (N_19052,N_13033,N_10136);
xor U19053 (N_19053,N_13134,N_11261);
or U19054 (N_19054,N_13193,N_13703);
nor U19055 (N_19055,N_13981,N_12188);
xnor U19056 (N_19056,N_14367,N_14287);
or U19057 (N_19057,N_10875,N_14789);
and U19058 (N_19058,N_14849,N_12468);
xor U19059 (N_19059,N_12798,N_13142);
or U19060 (N_19060,N_13817,N_12936);
or U19061 (N_19061,N_12258,N_12605);
xnor U19062 (N_19062,N_13093,N_13471);
and U19063 (N_19063,N_12907,N_11589);
xnor U19064 (N_19064,N_10988,N_11932);
or U19065 (N_19065,N_13946,N_10703);
and U19066 (N_19066,N_11270,N_13499);
or U19067 (N_19067,N_14051,N_13033);
or U19068 (N_19068,N_14180,N_13874);
and U19069 (N_19069,N_10972,N_14035);
nor U19070 (N_19070,N_14362,N_12921);
nor U19071 (N_19071,N_11478,N_11135);
and U19072 (N_19072,N_10614,N_11069);
or U19073 (N_19073,N_10102,N_14770);
nand U19074 (N_19074,N_13330,N_10921);
and U19075 (N_19075,N_10042,N_11349);
nand U19076 (N_19076,N_12384,N_10952);
and U19077 (N_19077,N_10322,N_14371);
or U19078 (N_19078,N_11624,N_14112);
and U19079 (N_19079,N_10325,N_13326);
xnor U19080 (N_19080,N_12783,N_11471);
xnor U19081 (N_19081,N_11055,N_12779);
xor U19082 (N_19082,N_13900,N_13491);
xor U19083 (N_19083,N_11930,N_11764);
nand U19084 (N_19084,N_13569,N_10275);
nand U19085 (N_19085,N_13969,N_13487);
nand U19086 (N_19086,N_13454,N_14888);
xnor U19087 (N_19087,N_14188,N_10354);
nand U19088 (N_19088,N_12744,N_12448);
nor U19089 (N_19089,N_12973,N_12557);
nand U19090 (N_19090,N_12391,N_14019);
nand U19091 (N_19091,N_12233,N_12620);
nand U19092 (N_19092,N_14813,N_10401);
or U19093 (N_19093,N_11842,N_12664);
xnor U19094 (N_19094,N_11316,N_10062);
nand U19095 (N_19095,N_12017,N_11027);
xnor U19096 (N_19096,N_11032,N_11896);
nand U19097 (N_19097,N_10609,N_12156);
nand U19098 (N_19098,N_12383,N_11556);
and U19099 (N_19099,N_13826,N_13036);
and U19100 (N_19100,N_12838,N_12786);
and U19101 (N_19101,N_14053,N_11044);
xor U19102 (N_19102,N_12002,N_11932);
nand U19103 (N_19103,N_14295,N_12021);
nor U19104 (N_19104,N_14897,N_14483);
nor U19105 (N_19105,N_12662,N_10521);
nor U19106 (N_19106,N_14078,N_10013);
or U19107 (N_19107,N_13290,N_12604);
xnor U19108 (N_19108,N_13993,N_10595);
nor U19109 (N_19109,N_11163,N_13097);
xnor U19110 (N_19110,N_12511,N_10766);
nand U19111 (N_19111,N_12458,N_11773);
xor U19112 (N_19112,N_12933,N_11078);
nor U19113 (N_19113,N_13808,N_13645);
nand U19114 (N_19114,N_12683,N_10157);
and U19115 (N_19115,N_12422,N_11820);
nand U19116 (N_19116,N_14123,N_13391);
and U19117 (N_19117,N_11664,N_14346);
nand U19118 (N_19118,N_11271,N_11789);
xnor U19119 (N_19119,N_10702,N_12646);
nand U19120 (N_19120,N_11254,N_10019);
xnor U19121 (N_19121,N_11404,N_13333);
and U19122 (N_19122,N_13767,N_11100);
nand U19123 (N_19123,N_11949,N_13911);
or U19124 (N_19124,N_14291,N_14195);
or U19125 (N_19125,N_13841,N_14798);
xor U19126 (N_19126,N_12205,N_13430);
or U19127 (N_19127,N_14994,N_13087);
nand U19128 (N_19128,N_11135,N_11106);
nor U19129 (N_19129,N_13990,N_14541);
xnor U19130 (N_19130,N_12807,N_13413);
or U19131 (N_19131,N_11747,N_13944);
xor U19132 (N_19132,N_14662,N_13528);
xor U19133 (N_19133,N_13479,N_11933);
nand U19134 (N_19134,N_12410,N_14759);
nand U19135 (N_19135,N_14135,N_12236);
nor U19136 (N_19136,N_13884,N_10945);
xnor U19137 (N_19137,N_11131,N_13944);
and U19138 (N_19138,N_13225,N_12527);
or U19139 (N_19139,N_13539,N_14602);
nor U19140 (N_19140,N_13766,N_10514);
and U19141 (N_19141,N_13809,N_14669);
and U19142 (N_19142,N_11756,N_14818);
xnor U19143 (N_19143,N_14548,N_10770);
or U19144 (N_19144,N_13661,N_10051);
and U19145 (N_19145,N_11234,N_12192);
nor U19146 (N_19146,N_11922,N_11429);
or U19147 (N_19147,N_11595,N_11971);
or U19148 (N_19148,N_13051,N_10737);
nor U19149 (N_19149,N_11292,N_12216);
or U19150 (N_19150,N_12344,N_10098);
nor U19151 (N_19151,N_14424,N_13892);
nor U19152 (N_19152,N_12257,N_13400);
or U19153 (N_19153,N_14856,N_11634);
or U19154 (N_19154,N_11898,N_10562);
nand U19155 (N_19155,N_10124,N_14352);
nor U19156 (N_19156,N_14717,N_13639);
or U19157 (N_19157,N_11265,N_12914);
nand U19158 (N_19158,N_10940,N_10045);
or U19159 (N_19159,N_13334,N_10512);
nor U19160 (N_19160,N_13776,N_10601);
or U19161 (N_19161,N_11363,N_13381);
nand U19162 (N_19162,N_10165,N_11443);
nand U19163 (N_19163,N_10944,N_12432);
or U19164 (N_19164,N_12309,N_10966);
nor U19165 (N_19165,N_13246,N_10189);
or U19166 (N_19166,N_10698,N_12585);
nand U19167 (N_19167,N_10329,N_14178);
and U19168 (N_19168,N_10690,N_13870);
nor U19169 (N_19169,N_14966,N_12741);
xnor U19170 (N_19170,N_10897,N_10204);
xor U19171 (N_19171,N_12878,N_12713);
or U19172 (N_19172,N_10415,N_12686);
or U19173 (N_19173,N_12261,N_13472);
nand U19174 (N_19174,N_11879,N_13119);
nand U19175 (N_19175,N_10859,N_11906);
or U19176 (N_19176,N_11682,N_14613);
and U19177 (N_19177,N_10394,N_13708);
or U19178 (N_19178,N_13693,N_10120);
xor U19179 (N_19179,N_11578,N_12847);
nor U19180 (N_19180,N_12023,N_14229);
xor U19181 (N_19181,N_11412,N_11740);
xnor U19182 (N_19182,N_11724,N_10676);
and U19183 (N_19183,N_10725,N_12732);
nor U19184 (N_19184,N_13591,N_14124);
and U19185 (N_19185,N_11489,N_14710);
xor U19186 (N_19186,N_11526,N_14183);
xnor U19187 (N_19187,N_12860,N_12422);
and U19188 (N_19188,N_12677,N_14420);
nor U19189 (N_19189,N_10677,N_12609);
and U19190 (N_19190,N_10327,N_10362);
or U19191 (N_19191,N_13718,N_12041);
and U19192 (N_19192,N_14744,N_13478);
xnor U19193 (N_19193,N_10843,N_13293);
or U19194 (N_19194,N_10561,N_13272);
xnor U19195 (N_19195,N_14150,N_10113);
and U19196 (N_19196,N_13941,N_11068);
nor U19197 (N_19197,N_11183,N_11044);
nand U19198 (N_19198,N_13795,N_12563);
or U19199 (N_19199,N_12530,N_10681);
nor U19200 (N_19200,N_10860,N_13090);
nor U19201 (N_19201,N_12557,N_11445);
nor U19202 (N_19202,N_10870,N_11787);
nand U19203 (N_19203,N_13134,N_12484);
nor U19204 (N_19204,N_10498,N_13954);
nand U19205 (N_19205,N_12658,N_13854);
and U19206 (N_19206,N_13121,N_11397);
or U19207 (N_19207,N_11672,N_14225);
nand U19208 (N_19208,N_13538,N_13516);
xor U19209 (N_19209,N_14063,N_10324);
nor U19210 (N_19210,N_11437,N_12116);
or U19211 (N_19211,N_12742,N_14563);
xor U19212 (N_19212,N_11121,N_12215);
and U19213 (N_19213,N_12802,N_11358);
or U19214 (N_19214,N_12743,N_14308);
or U19215 (N_19215,N_10310,N_12856);
and U19216 (N_19216,N_10767,N_13938);
nand U19217 (N_19217,N_12237,N_11893);
nor U19218 (N_19218,N_13235,N_10514);
xnor U19219 (N_19219,N_13606,N_13801);
and U19220 (N_19220,N_13053,N_14224);
xnor U19221 (N_19221,N_14847,N_14447);
and U19222 (N_19222,N_12088,N_12173);
nand U19223 (N_19223,N_10633,N_11359);
or U19224 (N_19224,N_12944,N_14335);
nor U19225 (N_19225,N_11324,N_10010);
nor U19226 (N_19226,N_12064,N_14889);
or U19227 (N_19227,N_10404,N_12069);
or U19228 (N_19228,N_12537,N_13083);
nor U19229 (N_19229,N_10733,N_13063);
xnor U19230 (N_19230,N_10097,N_11100);
and U19231 (N_19231,N_11528,N_11414);
xor U19232 (N_19232,N_13425,N_13755);
nand U19233 (N_19233,N_14270,N_14045);
or U19234 (N_19234,N_13203,N_12920);
nand U19235 (N_19235,N_13361,N_11757);
and U19236 (N_19236,N_13107,N_14939);
and U19237 (N_19237,N_10702,N_11437);
and U19238 (N_19238,N_14657,N_10377);
and U19239 (N_19239,N_14267,N_14257);
and U19240 (N_19240,N_10750,N_12385);
or U19241 (N_19241,N_13588,N_10697);
nand U19242 (N_19242,N_12261,N_11860);
nand U19243 (N_19243,N_10762,N_11030);
nand U19244 (N_19244,N_12220,N_10213);
nor U19245 (N_19245,N_12797,N_14023);
or U19246 (N_19246,N_14924,N_12297);
or U19247 (N_19247,N_13802,N_12067);
nand U19248 (N_19248,N_11439,N_12693);
xor U19249 (N_19249,N_14057,N_14102);
xor U19250 (N_19250,N_14448,N_12327);
and U19251 (N_19251,N_14128,N_12780);
xnor U19252 (N_19252,N_13228,N_14919);
and U19253 (N_19253,N_12321,N_14249);
nor U19254 (N_19254,N_12748,N_10177);
xnor U19255 (N_19255,N_11472,N_12334);
xnor U19256 (N_19256,N_14872,N_14453);
xor U19257 (N_19257,N_11831,N_10082);
xnor U19258 (N_19258,N_13996,N_14228);
and U19259 (N_19259,N_12102,N_11506);
xor U19260 (N_19260,N_14640,N_14312);
nor U19261 (N_19261,N_11483,N_11320);
nand U19262 (N_19262,N_13637,N_13128);
xnor U19263 (N_19263,N_14567,N_12260);
and U19264 (N_19264,N_14546,N_12304);
and U19265 (N_19265,N_13065,N_11276);
xnor U19266 (N_19266,N_11744,N_14104);
xnor U19267 (N_19267,N_14628,N_10553);
nand U19268 (N_19268,N_10035,N_10693);
nor U19269 (N_19269,N_13520,N_13246);
and U19270 (N_19270,N_10080,N_12803);
nand U19271 (N_19271,N_10291,N_14307);
or U19272 (N_19272,N_10501,N_11217);
and U19273 (N_19273,N_13697,N_11101);
or U19274 (N_19274,N_10425,N_10602);
xnor U19275 (N_19275,N_12545,N_11287);
and U19276 (N_19276,N_10982,N_10510);
nand U19277 (N_19277,N_13313,N_11540);
nand U19278 (N_19278,N_10033,N_11544);
and U19279 (N_19279,N_14063,N_11215);
nor U19280 (N_19280,N_13167,N_10859);
nand U19281 (N_19281,N_12982,N_13734);
nor U19282 (N_19282,N_10069,N_12371);
and U19283 (N_19283,N_11692,N_12907);
xnor U19284 (N_19284,N_13057,N_13988);
nand U19285 (N_19285,N_14707,N_11110);
nand U19286 (N_19286,N_10462,N_14814);
xnor U19287 (N_19287,N_12762,N_12586);
or U19288 (N_19288,N_10474,N_10710);
nor U19289 (N_19289,N_10172,N_13343);
or U19290 (N_19290,N_10530,N_11428);
xnor U19291 (N_19291,N_10126,N_12809);
nand U19292 (N_19292,N_11661,N_13252);
nand U19293 (N_19293,N_13140,N_14576);
nor U19294 (N_19294,N_12988,N_10449);
xor U19295 (N_19295,N_14840,N_14144);
or U19296 (N_19296,N_10300,N_10618);
and U19297 (N_19297,N_12491,N_10264);
or U19298 (N_19298,N_11763,N_14253);
and U19299 (N_19299,N_11906,N_11454);
and U19300 (N_19300,N_12805,N_13480);
and U19301 (N_19301,N_10858,N_12194);
nor U19302 (N_19302,N_14600,N_12151);
and U19303 (N_19303,N_12767,N_13904);
or U19304 (N_19304,N_14871,N_14615);
nand U19305 (N_19305,N_12100,N_13216);
and U19306 (N_19306,N_14926,N_14376);
and U19307 (N_19307,N_11460,N_12802);
nand U19308 (N_19308,N_14247,N_12483);
or U19309 (N_19309,N_10954,N_13508);
nand U19310 (N_19310,N_13339,N_13170);
or U19311 (N_19311,N_12247,N_10191);
and U19312 (N_19312,N_11563,N_10566);
nand U19313 (N_19313,N_10321,N_12927);
nor U19314 (N_19314,N_10788,N_14068);
or U19315 (N_19315,N_12703,N_14211);
nand U19316 (N_19316,N_14894,N_12516);
nand U19317 (N_19317,N_14727,N_14715);
or U19318 (N_19318,N_14042,N_10384);
nor U19319 (N_19319,N_13770,N_10367);
nand U19320 (N_19320,N_10179,N_13940);
nand U19321 (N_19321,N_11759,N_10072);
xor U19322 (N_19322,N_10585,N_13978);
and U19323 (N_19323,N_10294,N_14503);
nor U19324 (N_19324,N_11875,N_11039);
and U19325 (N_19325,N_10770,N_13890);
xor U19326 (N_19326,N_13366,N_13572);
nor U19327 (N_19327,N_12640,N_10130);
xor U19328 (N_19328,N_13381,N_12143);
or U19329 (N_19329,N_13225,N_11456);
and U19330 (N_19330,N_11111,N_10352);
or U19331 (N_19331,N_10419,N_11245);
xnor U19332 (N_19332,N_13410,N_13541);
nand U19333 (N_19333,N_12610,N_12359);
xnor U19334 (N_19334,N_11934,N_12281);
or U19335 (N_19335,N_12479,N_14896);
and U19336 (N_19336,N_12262,N_10734);
or U19337 (N_19337,N_14103,N_12893);
and U19338 (N_19338,N_14256,N_14219);
xor U19339 (N_19339,N_13137,N_14504);
or U19340 (N_19340,N_14705,N_14148);
and U19341 (N_19341,N_11004,N_11661);
nand U19342 (N_19342,N_13613,N_14785);
nand U19343 (N_19343,N_10524,N_10462);
nand U19344 (N_19344,N_11526,N_12598);
or U19345 (N_19345,N_12785,N_11627);
xor U19346 (N_19346,N_10693,N_11144);
or U19347 (N_19347,N_13470,N_14275);
xor U19348 (N_19348,N_10429,N_10314);
and U19349 (N_19349,N_14231,N_13272);
or U19350 (N_19350,N_13981,N_10282);
nand U19351 (N_19351,N_13925,N_13086);
nand U19352 (N_19352,N_12358,N_11295);
and U19353 (N_19353,N_12074,N_13582);
or U19354 (N_19354,N_14424,N_13338);
and U19355 (N_19355,N_10861,N_12462);
nand U19356 (N_19356,N_14253,N_12332);
xnor U19357 (N_19357,N_12956,N_10351);
xor U19358 (N_19358,N_13992,N_13640);
xnor U19359 (N_19359,N_13738,N_11557);
nor U19360 (N_19360,N_12314,N_11149);
and U19361 (N_19361,N_12094,N_11629);
xnor U19362 (N_19362,N_11366,N_10860);
xnor U19363 (N_19363,N_14745,N_10304);
or U19364 (N_19364,N_14529,N_12828);
or U19365 (N_19365,N_14264,N_14873);
and U19366 (N_19366,N_10372,N_14157);
and U19367 (N_19367,N_12693,N_13954);
and U19368 (N_19368,N_10774,N_14021);
and U19369 (N_19369,N_14418,N_14464);
and U19370 (N_19370,N_10428,N_11495);
or U19371 (N_19371,N_10877,N_11829);
nand U19372 (N_19372,N_11752,N_14889);
xor U19373 (N_19373,N_10282,N_13477);
nor U19374 (N_19374,N_14711,N_11158);
nand U19375 (N_19375,N_13670,N_12129);
nor U19376 (N_19376,N_12853,N_13324);
or U19377 (N_19377,N_10782,N_11683);
nor U19378 (N_19378,N_10204,N_12355);
or U19379 (N_19379,N_11226,N_11179);
nand U19380 (N_19380,N_13288,N_11086);
and U19381 (N_19381,N_13498,N_10160);
nand U19382 (N_19382,N_14839,N_11791);
nand U19383 (N_19383,N_13203,N_12365);
xor U19384 (N_19384,N_12872,N_14160);
nor U19385 (N_19385,N_10570,N_12386);
xor U19386 (N_19386,N_12206,N_11445);
nand U19387 (N_19387,N_14405,N_12053);
nor U19388 (N_19388,N_10562,N_11080);
or U19389 (N_19389,N_12876,N_12571);
or U19390 (N_19390,N_12206,N_11177);
or U19391 (N_19391,N_11906,N_14117);
or U19392 (N_19392,N_10290,N_12572);
and U19393 (N_19393,N_10501,N_13619);
nand U19394 (N_19394,N_10267,N_13292);
or U19395 (N_19395,N_12035,N_11366);
xnor U19396 (N_19396,N_10439,N_13107);
and U19397 (N_19397,N_10185,N_14185);
nand U19398 (N_19398,N_11583,N_13935);
nand U19399 (N_19399,N_11604,N_12303);
and U19400 (N_19400,N_11704,N_13179);
nand U19401 (N_19401,N_12426,N_12707);
and U19402 (N_19402,N_13476,N_11287);
and U19403 (N_19403,N_13626,N_10013);
nand U19404 (N_19404,N_12911,N_10232);
or U19405 (N_19405,N_11742,N_12540);
and U19406 (N_19406,N_13552,N_14198);
nor U19407 (N_19407,N_10423,N_14695);
or U19408 (N_19408,N_14102,N_10688);
nand U19409 (N_19409,N_11042,N_11140);
and U19410 (N_19410,N_13408,N_12042);
and U19411 (N_19411,N_14002,N_14393);
nor U19412 (N_19412,N_11646,N_12645);
nand U19413 (N_19413,N_10562,N_13133);
xor U19414 (N_19414,N_10593,N_14532);
nand U19415 (N_19415,N_13066,N_12404);
and U19416 (N_19416,N_12335,N_11534);
xor U19417 (N_19417,N_10655,N_13282);
xor U19418 (N_19418,N_14590,N_12871);
or U19419 (N_19419,N_12044,N_11476);
and U19420 (N_19420,N_12071,N_12674);
nor U19421 (N_19421,N_13249,N_14465);
and U19422 (N_19422,N_11381,N_12166);
and U19423 (N_19423,N_10512,N_12515);
xor U19424 (N_19424,N_13189,N_12008);
or U19425 (N_19425,N_12406,N_11830);
xnor U19426 (N_19426,N_14030,N_13181);
xnor U19427 (N_19427,N_11422,N_14247);
nand U19428 (N_19428,N_11568,N_14899);
nand U19429 (N_19429,N_11926,N_10619);
and U19430 (N_19430,N_10881,N_14120);
nor U19431 (N_19431,N_10972,N_14503);
or U19432 (N_19432,N_14890,N_12125);
nand U19433 (N_19433,N_14553,N_11954);
or U19434 (N_19434,N_14537,N_13840);
or U19435 (N_19435,N_10508,N_11087);
nor U19436 (N_19436,N_14926,N_12912);
xor U19437 (N_19437,N_13217,N_14410);
or U19438 (N_19438,N_14614,N_10705);
nor U19439 (N_19439,N_10685,N_10346);
nand U19440 (N_19440,N_13451,N_11153);
or U19441 (N_19441,N_14048,N_11405);
xor U19442 (N_19442,N_10076,N_12212);
nor U19443 (N_19443,N_11362,N_12802);
nand U19444 (N_19444,N_10072,N_14061);
xor U19445 (N_19445,N_14593,N_13857);
nand U19446 (N_19446,N_14808,N_14596);
and U19447 (N_19447,N_10843,N_11430);
or U19448 (N_19448,N_14608,N_13082);
nand U19449 (N_19449,N_14458,N_11304);
nor U19450 (N_19450,N_14762,N_11001);
nand U19451 (N_19451,N_11059,N_14823);
nor U19452 (N_19452,N_10951,N_12233);
and U19453 (N_19453,N_10740,N_13957);
nor U19454 (N_19454,N_13369,N_12610);
or U19455 (N_19455,N_14264,N_12535);
xor U19456 (N_19456,N_14247,N_12873);
and U19457 (N_19457,N_11775,N_11820);
nor U19458 (N_19458,N_12200,N_13830);
or U19459 (N_19459,N_11237,N_10667);
or U19460 (N_19460,N_10303,N_10106);
nor U19461 (N_19461,N_13891,N_10467);
and U19462 (N_19462,N_13461,N_11081);
xor U19463 (N_19463,N_14776,N_11693);
and U19464 (N_19464,N_14039,N_14512);
and U19465 (N_19465,N_11593,N_13970);
and U19466 (N_19466,N_10855,N_11151);
nor U19467 (N_19467,N_10304,N_12139);
xor U19468 (N_19468,N_12885,N_11360);
xor U19469 (N_19469,N_11928,N_14618);
nand U19470 (N_19470,N_12227,N_14484);
nor U19471 (N_19471,N_12841,N_13919);
or U19472 (N_19472,N_12722,N_13020);
xnor U19473 (N_19473,N_10078,N_11951);
nor U19474 (N_19474,N_10963,N_11766);
and U19475 (N_19475,N_11855,N_11363);
or U19476 (N_19476,N_14627,N_10028);
nand U19477 (N_19477,N_11040,N_11448);
nor U19478 (N_19478,N_11006,N_12054);
or U19479 (N_19479,N_11393,N_12065);
nand U19480 (N_19480,N_12806,N_10919);
and U19481 (N_19481,N_13622,N_14011);
xnor U19482 (N_19482,N_10333,N_13288);
nand U19483 (N_19483,N_11538,N_11042);
or U19484 (N_19484,N_14629,N_11886);
xor U19485 (N_19485,N_14346,N_14088);
nand U19486 (N_19486,N_12922,N_12053);
nand U19487 (N_19487,N_11406,N_12026);
nor U19488 (N_19488,N_13901,N_11619);
and U19489 (N_19489,N_11629,N_10160);
and U19490 (N_19490,N_11567,N_10969);
nor U19491 (N_19491,N_14041,N_12509);
nand U19492 (N_19492,N_10578,N_14898);
xor U19493 (N_19493,N_13445,N_10231);
nand U19494 (N_19494,N_11912,N_12979);
nand U19495 (N_19495,N_13622,N_12707);
or U19496 (N_19496,N_10847,N_10401);
and U19497 (N_19497,N_13325,N_10610);
or U19498 (N_19498,N_11508,N_13726);
or U19499 (N_19499,N_10987,N_11561);
xnor U19500 (N_19500,N_10212,N_10622);
nor U19501 (N_19501,N_10959,N_10862);
or U19502 (N_19502,N_12065,N_11685);
and U19503 (N_19503,N_10717,N_11944);
and U19504 (N_19504,N_12174,N_12958);
xor U19505 (N_19505,N_11422,N_12785);
or U19506 (N_19506,N_11885,N_10613);
or U19507 (N_19507,N_14785,N_10848);
or U19508 (N_19508,N_10713,N_10148);
and U19509 (N_19509,N_14492,N_10958);
xor U19510 (N_19510,N_14281,N_14372);
xnor U19511 (N_19511,N_14349,N_14063);
or U19512 (N_19512,N_12723,N_10740);
nor U19513 (N_19513,N_12878,N_11056);
xor U19514 (N_19514,N_13481,N_12211);
or U19515 (N_19515,N_14878,N_10373);
and U19516 (N_19516,N_13342,N_14312);
nand U19517 (N_19517,N_11670,N_14607);
or U19518 (N_19518,N_13869,N_14209);
nand U19519 (N_19519,N_11770,N_12662);
and U19520 (N_19520,N_13654,N_11781);
and U19521 (N_19521,N_13540,N_11922);
nor U19522 (N_19522,N_11050,N_10555);
nand U19523 (N_19523,N_13842,N_10645);
or U19524 (N_19524,N_11405,N_12137);
nor U19525 (N_19525,N_13379,N_11428);
and U19526 (N_19526,N_10057,N_12444);
and U19527 (N_19527,N_10482,N_13534);
or U19528 (N_19528,N_13360,N_12348);
nand U19529 (N_19529,N_12749,N_13679);
nand U19530 (N_19530,N_12713,N_12485);
nor U19531 (N_19531,N_14582,N_11774);
xnor U19532 (N_19532,N_13660,N_11359);
xnor U19533 (N_19533,N_10428,N_10218);
and U19534 (N_19534,N_12956,N_10502);
nor U19535 (N_19535,N_12571,N_12435);
nand U19536 (N_19536,N_13840,N_14604);
and U19537 (N_19537,N_11897,N_12640);
and U19538 (N_19538,N_10027,N_13119);
nor U19539 (N_19539,N_10433,N_11540);
nor U19540 (N_19540,N_11415,N_13197);
xor U19541 (N_19541,N_11754,N_13785);
or U19542 (N_19542,N_13461,N_10600);
or U19543 (N_19543,N_10222,N_14357);
and U19544 (N_19544,N_13953,N_14972);
xnor U19545 (N_19545,N_13841,N_10452);
nor U19546 (N_19546,N_11890,N_12561);
and U19547 (N_19547,N_11929,N_13128);
and U19548 (N_19548,N_11362,N_14891);
nand U19549 (N_19549,N_14584,N_13493);
and U19550 (N_19550,N_11023,N_11298);
xnor U19551 (N_19551,N_11683,N_10392);
nand U19552 (N_19552,N_10275,N_10871);
and U19553 (N_19553,N_12200,N_14288);
nor U19554 (N_19554,N_12564,N_11387);
and U19555 (N_19555,N_13016,N_12392);
xor U19556 (N_19556,N_10088,N_11214);
and U19557 (N_19557,N_12639,N_10816);
and U19558 (N_19558,N_11450,N_12605);
and U19559 (N_19559,N_12542,N_12841);
xor U19560 (N_19560,N_10139,N_14847);
xnor U19561 (N_19561,N_11983,N_13827);
xnor U19562 (N_19562,N_12485,N_13067);
and U19563 (N_19563,N_12928,N_10160);
nand U19564 (N_19564,N_10673,N_11153);
and U19565 (N_19565,N_13791,N_13060);
nand U19566 (N_19566,N_12459,N_13251);
or U19567 (N_19567,N_13202,N_12097);
xnor U19568 (N_19568,N_12498,N_11697);
nand U19569 (N_19569,N_14209,N_11716);
or U19570 (N_19570,N_13738,N_11604);
or U19571 (N_19571,N_12115,N_12473);
and U19572 (N_19572,N_10574,N_12332);
xor U19573 (N_19573,N_12480,N_13285);
nor U19574 (N_19574,N_12251,N_10057);
nand U19575 (N_19575,N_13173,N_11675);
nand U19576 (N_19576,N_10963,N_14470);
nand U19577 (N_19577,N_10608,N_14659);
nor U19578 (N_19578,N_13326,N_12177);
xor U19579 (N_19579,N_10035,N_13241);
or U19580 (N_19580,N_10540,N_11341);
xor U19581 (N_19581,N_13491,N_13071);
xnor U19582 (N_19582,N_12469,N_12802);
and U19583 (N_19583,N_14112,N_13953);
xnor U19584 (N_19584,N_10536,N_10146);
xnor U19585 (N_19585,N_12738,N_12909);
nand U19586 (N_19586,N_14520,N_11380);
nor U19587 (N_19587,N_13224,N_12545);
and U19588 (N_19588,N_14159,N_13243);
nor U19589 (N_19589,N_10672,N_14444);
nor U19590 (N_19590,N_10152,N_12410);
nor U19591 (N_19591,N_13947,N_10632);
xor U19592 (N_19592,N_12058,N_12525);
and U19593 (N_19593,N_13413,N_13817);
or U19594 (N_19594,N_13161,N_13250);
nand U19595 (N_19595,N_11516,N_13166);
xnor U19596 (N_19596,N_11819,N_12370);
nand U19597 (N_19597,N_12566,N_10613);
and U19598 (N_19598,N_14138,N_13551);
nor U19599 (N_19599,N_11266,N_13678);
nor U19600 (N_19600,N_11113,N_11966);
and U19601 (N_19601,N_10225,N_13000);
nor U19602 (N_19602,N_12379,N_10454);
nor U19603 (N_19603,N_13427,N_13386);
nand U19604 (N_19604,N_11285,N_11631);
or U19605 (N_19605,N_11570,N_13812);
nor U19606 (N_19606,N_10988,N_10535);
nor U19607 (N_19607,N_11552,N_11138);
nor U19608 (N_19608,N_12420,N_14694);
nor U19609 (N_19609,N_12863,N_14375);
nor U19610 (N_19610,N_14259,N_13975);
and U19611 (N_19611,N_10339,N_11656);
nor U19612 (N_19612,N_10389,N_11136);
xnor U19613 (N_19613,N_10979,N_13465);
nand U19614 (N_19614,N_13243,N_14471);
nor U19615 (N_19615,N_11221,N_12259);
nor U19616 (N_19616,N_14889,N_11338);
nor U19617 (N_19617,N_10697,N_11148);
xor U19618 (N_19618,N_12393,N_14161);
and U19619 (N_19619,N_13215,N_12438);
xor U19620 (N_19620,N_10947,N_11602);
or U19621 (N_19621,N_12706,N_10935);
nor U19622 (N_19622,N_11699,N_13594);
nor U19623 (N_19623,N_12825,N_11270);
nand U19624 (N_19624,N_10154,N_12786);
and U19625 (N_19625,N_10263,N_11290);
or U19626 (N_19626,N_11096,N_14512);
xor U19627 (N_19627,N_12027,N_14719);
nand U19628 (N_19628,N_12041,N_10885);
nor U19629 (N_19629,N_13848,N_10177);
nand U19630 (N_19630,N_10419,N_10320);
and U19631 (N_19631,N_14077,N_11942);
and U19632 (N_19632,N_12242,N_11637);
and U19633 (N_19633,N_12090,N_13885);
xnor U19634 (N_19634,N_13274,N_14663);
nand U19635 (N_19635,N_10439,N_13731);
and U19636 (N_19636,N_11241,N_10192);
xor U19637 (N_19637,N_11876,N_11092);
nand U19638 (N_19638,N_12264,N_11944);
nand U19639 (N_19639,N_10021,N_10512);
or U19640 (N_19640,N_11835,N_11216);
xnor U19641 (N_19641,N_12025,N_11915);
nor U19642 (N_19642,N_14309,N_14639);
or U19643 (N_19643,N_12985,N_12463);
and U19644 (N_19644,N_10017,N_14258);
xnor U19645 (N_19645,N_13310,N_14432);
xor U19646 (N_19646,N_12503,N_13501);
or U19647 (N_19647,N_12838,N_13496);
nor U19648 (N_19648,N_11274,N_12164);
nand U19649 (N_19649,N_14943,N_12832);
nor U19650 (N_19650,N_10718,N_14959);
or U19651 (N_19651,N_14909,N_14689);
nand U19652 (N_19652,N_13176,N_14407);
nand U19653 (N_19653,N_12950,N_14885);
nor U19654 (N_19654,N_10103,N_12893);
and U19655 (N_19655,N_10332,N_10601);
and U19656 (N_19656,N_13504,N_11183);
and U19657 (N_19657,N_12591,N_13474);
and U19658 (N_19658,N_11578,N_11639);
nor U19659 (N_19659,N_11404,N_12348);
nor U19660 (N_19660,N_13422,N_13094);
xor U19661 (N_19661,N_14784,N_12987);
nand U19662 (N_19662,N_14517,N_12672);
nand U19663 (N_19663,N_13022,N_14696);
and U19664 (N_19664,N_10760,N_13227);
xnor U19665 (N_19665,N_14325,N_10665);
nand U19666 (N_19666,N_14692,N_10305);
nand U19667 (N_19667,N_13616,N_13354);
nand U19668 (N_19668,N_10074,N_11035);
xnor U19669 (N_19669,N_10927,N_11483);
or U19670 (N_19670,N_10300,N_14775);
nand U19671 (N_19671,N_10139,N_11454);
nand U19672 (N_19672,N_13182,N_10867);
nor U19673 (N_19673,N_11143,N_14987);
xor U19674 (N_19674,N_11940,N_13819);
nor U19675 (N_19675,N_14272,N_10849);
and U19676 (N_19676,N_12457,N_10130);
and U19677 (N_19677,N_14513,N_12761);
nor U19678 (N_19678,N_12701,N_10746);
nand U19679 (N_19679,N_12225,N_14601);
nor U19680 (N_19680,N_10014,N_14788);
or U19681 (N_19681,N_13382,N_12276);
or U19682 (N_19682,N_10929,N_13943);
xor U19683 (N_19683,N_11173,N_14394);
nand U19684 (N_19684,N_10567,N_11864);
xor U19685 (N_19685,N_13184,N_12588);
and U19686 (N_19686,N_14173,N_10864);
and U19687 (N_19687,N_12310,N_13824);
and U19688 (N_19688,N_13417,N_13390);
nor U19689 (N_19689,N_12579,N_10089);
or U19690 (N_19690,N_10914,N_12438);
xnor U19691 (N_19691,N_11098,N_14612);
nand U19692 (N_19692,N_11533,N_13957);
nand U19693 (N_19693,N_10842,N_13697);
xnor U19694 (N_19694,N_12840,N_11423);
and U19695 (N_19695,N_12399,N_13589);
and U19696 (N_19696,N_11749,N_14606);
nor U19697 (N_19697,N_10794,N_11024);
xor U19698 (N_19698,N_14230,N_10289);
or U19699 (N_19699,N_13550,N_14624);
nand U19700 (N_19700,N_11962,N_10644);
or U19701 (N_19701,N_11786,N_14679);
nand U19702 (N_19702,N_11481,N_14597);
nand U19703 (N_19703,N_13797,N_14933);
nand U19704 (N_19704,N_14056,N_11570);
and U19705 (N_19705,N_10999,N_11083);
nor U19706 (N_19706,N_12049,N_14215);
or U19707 (N_19707,N_13028,N_11523);
or U19708 (N_19708,N_10753,N_13975);
nand U19709 (N_19709,N_11332,N_12466);
nor U19710 (N_19710,N_13237,N_14608);
nor U19711 (N_19711,N_13004,N_12445);
nor U19712 (N_19712,N_10721,N_12198);
nor U19713 (N_19713,N_14664,N_14520);
nand U19714 (N_19714,N_12502,N_11789);
and U19715 (N_19715,N_10660,N_10861);
nand U19716 (N_19716,N_14864,N_12576);
nand U19717 (N_19717,N_11397,N_12382);
or U19718 (N_19718,N_10235,N_10647);
xnor U19719 (N_19719,N_14158,N_12821);
nand U19720 (N_19720,N_13838,N_12541);
or U19721 (N_19721,N_14277,N_12098);
or U19722 (N_19722,N_13511,N_11886);
nor U19723 (N_19723,N_10897,N_10086);
nor U19724 (N_19724,N_10594,N_12246);
nand U19725 (N_19725,N_13852,N_10726);
nor U19726 (N_19726,N_14067,N_10940);
and U19727 (N_19727,N_12684,N_13736);
or U19728 (N_19728,N_14243,N_13421);
and U19729 (N_19729,N_11777,N_12747);
and U19730 (N_19730,N_12317,N_13533);
and U19731 (N_19731,N_11831,N_12781);
nand U19732 (N_19732,N_14134,N_14859);
and U19733 (N_19733,N_12969,N_11567);
nor U19734 (N_19734,N_11279,N_10173);
or U19735 (N_19735,N_11789,N_12720);
or U19736 (N_19736,N_13587,N_13911);
or U19737 (N_19737,N_13114,N_10350);
or U19738 (N_19738,N_14223,N_14163);
or U19739 (N_19739,N_14406,N_14291);
or U19740 (N_19740,N_13394,N_12350);
nor U19741 (N_19741,N_11917,N_14820);
xor U19742 (N_19742,N_13267,N_14093);
or U19743 (N_19743,N_11179,N_10551);
xor U19744 (N_19744,N_14692,N_13536);
nor U19745 (N_19745,N_11425,N_10903);
and U19746 (N_19746,N_12385,N_10377);
xor U19747 (N_19747,N_11241,N_11381);
xor U19748 (N_19748,N_13762,N_13331);
nand U19749 (N_19749,N_10076,N_13321);
and U19750 (N_19750,N_12759,N_12894);
or U19751 (N_19751,N_11909,N_12382);
xor U19752 (N_19752,N_12208,N_14186);
or U19753 (N_19753,N_11186,N_12654);
nor U19754 (N_19754,N_10865,N_14093);
and U19755 (N_19755,N_11598,N_12051);
nor U19756 (N_19756,N_11497,N_14714);
nor U19757 (N_19757,N_12210,N_11184);
or U19758 (N_19758,N_12809,N_12432);
nand U19759 (N_19759,N_11012,N_11075);
or U19760 (N_19760,N_13131,N_10425);
and U19761 (N_19761,N_13755,N_11799);
nor U19762 (N_19762,N_11273,N_14118);
and U19763 (N_19763,N_10171,N_10053);
and U19764 (N_19764,N_12670,N_12514);
nand U19765 (N_19765,N_11344,N_10166);
or U19766 (N_19766,N_11065,N_12424);
xor U19767 (N_19767,N_12807,N_14822);
xor U19768 (N_19768,N_10895,N_10856);
xnor U19769 (N_19769,N_12666,N_10556);
and U19770 (N_19770,N_11924,N_11944);
or U19771 (N_19771,N_12565,N_13502);
and U19772 (N_19772,N_13042,N_13058);
or U19773 (N_19773,N_14388,N_14571);
and U19774 (N_19774,N_14042,N_14318);
or U19775 (N_19775,N_12251,N_14889);
nand U19776 (N_19776,N_14299,N_14060);
or U19777 (N_19777,N_10971,N_11787);
nor U19778 (N_19778,N_13936,N_10340);
nand U19779 (N_19779,N_14200,N_14701);
nor U19780 (N_19780,N_13604,N_12007);
nor U19781 (N_19781,N_11188,N_13555);
xnor U19782 (N_19782,N_10909,N_12420);
nand U19783 (N_19783,N_12396,N_13643);
nand U19784 (N_19784,N_14066,N_14514);
and U19785 (N_19785,N_11174,N_14945);
xor U19786 (N_19786,N_11608,N_12979);
nor U19787 (N_19787,N_14055,N_12408);
xnor U19788 (N_19788,N_11987,N_12970);
and U19789 (N_19789,N_12429,N_11357);
nand U19790 (N_19790,N_13411,N_10392);
nor U19791 (N_19791,N_13947,N_11485);
nand U19792 (N_19792,N_11554,N_13285);
nor U19793 (N_19793,N_10088,N_12634);
xor U19794 (N_19794,N_10041,N_14355);
xor U19795 (N_19795,N_14417,N_10705);
xor U19796 (N_19796,N_14254,N_11624);
and U19797 (N_19797,N_12299,N_12267);
xor U19798 (N_19798,N_11069,N_14421);
nor U19799 (N_19799,N_13035,N_13936);
nand U19800 (N_19800,N_10328,N_13035);
xnor U19801 (N_19801,N_11072,N_13995);
nor U19802 (N_19802,N_11640,N_10243);
xnor U19803 (N_19803,N_13448,N_10240);
or U19804 (N_19804,N_13360,N_14680);
xor U19805 (N_19805,N_11952,N_12239);
and U19806 (N_19806,N_13322,N_10963);
xnor U19807 (N_19807,N_14499,N_14062);
and U19808 (N_19808,N_13512,N_14282);
or U19809 (N_19809,N_10352,N_11348);
nor U19810 (N_19810,N_14171,N_14354);
xor U19811 (N_19811,N_12810,N_13373);
and U19812 (N_19812,N_11689,N_10901);
xor U19813 (N_19813,N_10132,N_12331);
nand U19814 (N_19814,N_11130,N_11206);
xor U19815 (N_19815,N_12077,N_14028);
nand U19816 (N_19816,N_10623,N_14950);
nor U19817 (N_19817,N_12622,N_13579);
or U19818 (N_19818,N_11112,N_10974);
nor U19819 (N_19819,N_11057,N_12678);
xor U19820 (N_19820,N_11248,N_11476);
nor U19821 (N_19821,N_12729,N_11060);
nand U19822 (N_19822,N_10874,N_14770);
nand U19823 (N_19823,N_14100,N_10683);
nor U19824 (N_19824,N_10709,N_13213);
and U19825 (N_19825,N_10274,N_13321);
or U19826 (N_19826,N_10227,N_11504);
xor U19827 (N_19827,N_12525,N_11839);
xor U19828 (N_19828,N_11117,N_14946);
nand U19829 (N_19829,N_14331,N_11862);
nand U19830 (N_19830,N_10042,N_10202);
nand U19831 (N_19831,N_13894,N_11175);
or U19832 (N_19832,N_13853,N_11520);
and U19833 (N_19833,N_11457,N_14040);
nand U19834 (N_19834,N_13946,N_10504);
or U19835 (N_19835,N_12681,N_14687);
nor U19836 (N_19836,N_12278,N_13763);
nand U19837 (N_19837,N_12275,N_10175);
or U19838 (N_19838,N_13925,N_14951);
xnor U19839 (N_19839,N_14649,N_12068);
nor U19840 (N_19840,N_10193,N_12702);
xor U19841 (N_19841,N_14567,N_14282);
or U19842 (N_19842,N_12555,N_10075);
or U19843 (N_19843,N_12287,N_12803);
and U19844 (N_19844,N_12817,N_10872);
or U19845 (N_19845,N_14546,N_11697);
nand U19846 (N_19846,N_11484,N_12390);
nand U19847 (N_19847,N_12444,N_12920);
xnor U19848 (N_19848,N_14419,N_10056);
xor U19849 (N_19849,N_14936,N_13422);
and U19850 (N_19850,N_14139,N_10217);
xnor U19851 (N_19851,N_10665,N_14371);
nand U19852 (N_19852,N_10709,N_10569);
and U19853 (N_19853,N_10614,N_11362);
or U19854 (N_19854,N_11268,N_14396);
and U19855 (N_19855,N_10101,N_10415);
xor U19856 (N_19856,N_12558,N_10284);
or U19857 (N_19857,N_12043,N_14855);
xnor U19858 (N_19858,N_14613,N_12806);
nand U19859 (N_19859,N_14333,N_10714);
nor U19860 (N_19860,N_13412,N_13148);
nand U19861 (N_19861,N_11707,N_14988);
and U19862 (N_19862,N_11655,N_14024);
nor U19863 (N_19863,N_13034,N_11331);
nand U19864 (N_19864,N_12717,N_11492);
nor U19865 (N_19865,N_10029,N_10499);
xnor U19866 (N_19866,N_14556,N_12882);
or U19867 (N_19867,N_14912,N_14800);
nand U19868 (N_19868,N_12762,N_13963);
and U19869 (N_19869,N_11617,N_13581);
and U19870 (N_19870,N_10259,N_13757);
xor U19871 (N_19871,N_12861,N_10231);
nand U19872 (N_19872,N_12687,N_13272);
xnor U19873 (N_19873,N_14406,N_11755);
and U19874 (N_19874,N_10417,N_12416);
xnor U19875 (N_19875,N_13460,N_14908);
or U19876 (N_19876,N_14202,N_10067);
and U19877 (N_19877,N_11884,N_13108);
and U19878 (N_19878,N_13044,N_14928);
or U19879 (N_19879,N_13349,N_13212);
nand U19880 (N_19880,N_14791,N_12577);
and U19881 (N_19881,N_14514,N_12114);
nor U19882 (N_19882,N_10526,N_10754);
nor U19883 (N_19883,N_12072,N_13882);
nor U19884 (N_19884,N_14574,N_12551);
nor U19885 (N_19885,N_10296,N_13184);
nand U19886 (N_19886,N_13031,N_14447);
nor U19887 (N_19887,N_12085,N_14830);
nor U19888 (N_19888,N_14723,N_12777);
or U19889 (N_19889,N_12669,N_12679);
nor U19890 (N_19890,N_10878,N_10137);
nor U19891 (N_19891,N_14504,N_12580);
or U19892 (N_19892,N_12384,N_10448);
nor U19893 (N_19893,N_12488,N_10214);
or U19894 (N_19894,N_12743,N_12973);
nor U19895 (N_19895,N_13152,N_11634);
or U19896 (N_19896,N_13955,N_11813);
xor U19897 (N_19897,N_12594,N_13829);
or U19898 (N_19898,N_10285,N_10241);
nor U19899 (N_19899,N_12569,N_13542);
xnor U19900 (N_19900,N_10214,N_14200);
and U19901 (N_19901,N_11567,N_12626);
xor U19902 (N_19902,N_12698,N_10635);
and U19903 (N_19903,N_11822,N_10461);
xnor U19904 (N_19904,N_12657,N_11320);
or U19905 (N_19905,N_14991,N_14265);
nand U19906 (N_19906,N_10611,N_14153);
nor U19907 (N_19907,N_13382,N_14706);
or U19908 (N_19908,N_11580,N_13157);
and U19909 (N_19909,N_10648,N_13437);
nor U19910 (N_19910,N_14920,N_13645);
nor U19911 (N_19911,N_14969,N_13164);
nand U19912 (N_19912,N_14218,N_12112);
nor U19913 (N_19913,N_10489,N_12692);
nand U19914 (N_19914,N_14576,N_10683);
nand U19915 (N_19915,N_10263,N_10288);
xor U19916 (N_19916,N_14101,N_11684);
and U19917 (N_19917,N_11276,N_11899);
nand U19918 (N_19918,N_13023,N_12282);
or U19919 (N_19919,N_12897,N_12679);
xnor U19920 (N_19920,N_10876,N_11764);
nor U19921 (N_19921,N_14124,N_12267);
xor U19922 (N_19922,N_13264,N_11767);
or U19923 (N_19923,N_12467,N_10672);
or U19924 (N_19924,N_13271,N_13765);
and U19925 (N_19925,N_10038,N_12615);
xor U19926 (N_19926,N_14562,N_12163);
xnor U19927 (N_19927,N_11804,N_12207);
and U19928 (N_19928,N_10557,N_12910);
or U19929 (N_19929,N_12118,N_10466);
nand U19930 (N_19930,N_14000,N_11012);
nor U19931 (N_19931,N_10396,N_10761);
nor U19932 (N_19932,N_12705,N_12649);
nand U19933 (N_19933,N_11300,N_13206);
and U19934 (N_19934,N_14863,N_13140);
or U19935 (N_19935,N_10992,N_10722);
xor U19936 (N_19936,N_13028,N_13266);
nor U19937 (N_19937,N_13370,N_11887);
nor U19938 (N_19938,N_10886,N_12716);
and U19939 (N_19939,N_12014,N_14470);
and U19940 (N_19940,N_13691,N_11736);
nand U19941 (N_19941,N_13286,N_11334);
or U19942 (N_19942,N_11834,N_14685);
nor U19943 (N_19943,N_14981,N_12574);
xnor U19944 (N_19944,N_11316,N_10136);
nor U19945 (N_19945,N_14629,N_12538);
or U19946 (N_19946,N_10011,N_12629);
and U19947 (N_19947,N_14175,N_14168);
xor U19948 (N_19948,N_11438,N_11750);
or U19949 (N_19949,N_10808,N_12530);
xor U19950 (N_19950,N_12442,N_10642);
nor U19951 (N_19951,N_11031,N_12773);
nor U19952 (N_19952,N_14185,N_10102);
and U19953 (N_19953,N_14938,N_11886);
nand U19954 (N_19954,N_14531,N_10692);
or U19955 (N_19955,N_10871,N_13840);
xnor U19956 (N_19956,N_13287,N_13045);
or U19957 (N_19957,N_14278,N_14700);
xor U19958 (N_19958,N_13346,N_13831);
nand U19959 (N_19959,N_13542,N_13745);
nor U19960 (N_19960,N_13843,N_11282);
xnor U19961 (N_19961,N_13749,N_14144);
nand U19962 (N_19962,N_13699,N_11687);
and U19963 (N_19963,N_14988,N_13946);
or U19964 (N_19964,N_14333,N_12229);
and U19965 (N_19965,N_14983,N_14787);
nand U19966 (N_19966,N_10152,N_14010);
nor U19967 (N_19967,N_14254,N_14391);
nor U19968 (N_19968,N_14591,N_13964);
and U19969 (N_19969,N_10369,N_11929);
nand U19970 (N_19970,N_10727,N_11338);
and U19971 (N_19971,N_14924,N_10138);
nor U19972 (N_19972,N_13207,N_10075);
and U19973 (N_19973,N_13818,N_13136);
nand U19974 (N_19974,N_10189,N_14785);
xor U19975 (N_19975,N_12135,N_13551);
and U19976 (N_19976,N_12795,N_13704);
nor U19977 (N_19977,N_11410,N_11113);
xor U19978 (N_19978,N_10951,N_10814);
nand U19979 (N_19979,N_11211,N_11782);
and U19980 (N_19980,N_10274,N_13274);
nor U19981 (N_19981,N_12829,N_10804);
nor U19982 (N_19982,N_13932,N_14426);
and U19983 (N_19983,N_13065,N_10421);
and U19984 (N_19984,N_13272,N_13235);
nand U19985 (N_19985,N_10925,N_11441);
nor U19986 (N_19986,N_14751,N_13253);
or U19987 (N_19987,N_10600,N_10689);
xnor U19988 (N_19988,N_13698,N_14117);
and U19989 (N_19989,N_10229,N_14686);
xor U19990 (N_19990,N_11432,N_10622);
nand U19991 (N_19991,N_13833,N_11174);
nor U19992 (N_19992,N_12093,N_14567);
nand U19993 (N_19993,N_13698,N_12186);
or U19994 (N_19994,N_12526,N_14848);
nor U19995 (N_19995,N_10948,N_11905);
nor U19996 (N_19996,N_11727,N_10150);
nand U19997 (N_19997,N_11803,N_12746);
or U19998 (N_19998,N_10896,N_11480);
nor U19999 (N_19999,N_13811,N_11462);
and UO_0 (O_0,N_17061,N_16129);
nand UO_1 (O_1,N_15750,N_17871);
or UO_2 (O_2,N_18566,N_18662);
or UO_3 (O_3,N_15509,N_19633);
or UO_4 (O_4,N_18868,N_17227);
and UO_5 (O_5,N_17882,N_17694);
nor UO_6 (O_6,N_18444,N_18796);
nor UO_7 (O_7,N_18733,N_16297);
nand UO_8 (O_8,N_19872,N_18339);
and UO_9 (O_9,N_16888,N_16689);
nor UO_10 (O_10,N_15963,N_15342);
xnor UO_11 (O_11,N_15320,N_16156);
and UO_12 (O_12,N_19319,N_18888);
nand UO_13 (O_13,N_18192,N_18001);
or UO_14 (O_14,N_18772,N_15127);
or UO_15 (O_15,N_15887,N_16456);
nand UO_16 (O_16,N_17373,N_19599);
nor UO_17 (O_17,N_16474,N_19969);
xnor UO_18 (O_18,N_18659,N_19860);
nand UO_19 (O_19,N_19728,N_18619);
xnor UO_20 (O_20,N_15197,N_18926);
xnor UO_21 (O_21,N_16414,N_15852);
and UO_22 (O_22,N_17708,N_15224);
nor UO_23 (O_23,N_17327,N_16558);
nand UO_24 (O_24,N_17656,N_19799);
nor UO_25 (O_25,N_16669,N_16730);
xnor UO_26 (O_26,N_17617,N_16963);
nor UO_27 (O_27,N_17726,N_18626);
nor UO_28 (O_28,N_16366,N_15591);
and UO_29 (O_29,N_15986,N_17429);
or UO_30 (O_30,N_18488,N_19168);
and UO_31 (O_31,N_19592,N_17719);
and UO_32 (O_32,N_16548,N_18138);
nor UO_33 (O_33,N_17401,N_15882);
xor UO_34 (O_34,N_16684,N_18225);
or UO_35 (O_35,N_17380,N_15310);
and UO_36 (O_36,N_17321,N_19097);
xor UO_37 (O_37,N_15816,N_19219);
nor UO_38 (O_38,N_19618,N_16628);
or UO_39 (O_39,N_15713,N_16819);
and UO_40 (O_40,N_19119,N_15794);
and UO_41 (O_41,N_16429,N_18264);
or UO_42 (O_42,N_15215,N_16069);
nand UO_43 (O_43,N_17104,N_16728);
xor UO_44 (O_44,N_15548,N_17734);
nor UO_45 (O_45,N_15235,N_19296);
nor UO_46 (O_46,N_19626,N_15672);
nor UO_47 (O_47,N_18840,N_16394);
xor UO_48 (O_48,N_15427,N_19444);
or UO_49 (O_49,N_17875,N_17998);
nor UO_50 (O_50,N_18473,N_16216);
nor UO_51 (O_51,N_19758,N_15468);
nor UO_52 (O_52,N_19501,N_19896);
and UO_53 (O_53,N_16640,N_17736);
and UO_54 (O_54,N_17986,N_15451);
nand UO_55 (O_55,N_16504,N_16149);
or UO_56 (O_56,N_18308,N_15677);
nor UO_57 (O_57,N_19297,N_16946);
or UO_58 (O_58,N_15329,N_18597);
nor UO_59 (O_59,N_15757,N_18744);
nand UO_60 (O_60,N_19063,N_19265);
xor UO_61 (O_61,N_16421,N_19846);
or UO_62 (O_62,N_15179,N_16067);
nor UO_63 (O_63,N_17535,N_18025);
nand UO_64 (O_64,N_19263,N_17443);
xnor UO_65 (O_65,N_16341,N_16844);
xnor UO_66 (O_66,N_17696,N_16180);
nand UO_67 (O_67,N_19649,N_16228);
nor UO_68 (O_68,N_15169,N_18393);
xnor UO_69 (O_69,N_17755,N_16713);
and UO_70 (O_70,N_15970,N_19900);
nand UO_71 (O_71,N_15174,N_18831);
nand UO_72 (O_72,N_15878,N_18305);
nor UO_73 (O_73,N_18203,N_17873);
nand UO_74 (O_74,N_17156,N_15621);
and UO_75 (O_75,N_16092,N_16993);
xor UO_76 (O_76,N_19556,N_15643);
xnor UO_77 (O_77,N_18380,N_18923);
and UO_78 (O_78,N_15168,N_18751);
or UO_79 (O_79,N_18351,N_18104);
or UO_80 (O_80,N_19164,N_16376);
nand UO_81 (O_81,N_18412,N_15270);
xor UO_82 (O_82,N_19103,N_19762);
nand UO_83 (O_83,N_16039,N_17878);
nor UO_84 (O_84,N_19970,N_16931);
nor UO_85 (O_85,N_15132,N_17364);
or UO_86 (O_86,N_16295,N_18016);
and UO_87 (O_87,N_19137,N_19777);
nor UO_88 (O_88,N_16837,N_17682);
xnor UO_89 (O_89,N_16289,N_16442);
nor UO_90 (O_90,N_15438,N_15292);
nand UO_91 (O_91,N_18310,N_17253);
nor UO_92 (O_92,N_18902,N_16758);
or UO_93 (O_93,N_17490,N_17032);
nor UO_94 (O_94,N_15200,N_15130);
nand UO_95 (O_95,N_16538,N_19014);
or UO_96 (O_96,N_18789,N_17823);
xor UO_97 (O_97,N_15767,N_17125);
nand UO_98 (O_98,N_19174,N_19347);
and UO_99 (O_99,N_15546,N_17495);
nor UO_100 (O_100,N_16094,N_19867);
nand UO_101 (O_101,N_17920,N_15289);
or UO_102 (O_102,N_17711,N_17833);
or UO_103 (O_103,N_17685,N_15908);
nand UO_104 (O_104,N_16311,N_19515);
nor UO_105 (O_105,N_17519,N_17663);
nor UO_106 (O_106,N_19227,N_19722);
or UO_107 (O_107,N_16405,N_18188);
or UO_108 (O_108,N_19432,N_18767);
and UO_109 (O_109,N_18136,N_18642);
nor UO_110 (O_110,N_18986,N_17994);
nand UO_111 (O_111,N_16162,N_16170);
nand UO_112 (O_112,N_17573,N_19800);
xnor UO_113 (O_113,N_15349,N_15964);
xnor UO_114 (O_114,N_18937,N_17971);
or UO_115 (O_115,N_16920,N_15830);
nor UO_116 (O_116,N_16412,N_17187);
or UO_117 (O_117,N_17133,N_16072);
and UO_118 (O_118,N_16594,N_15516);
and UO_119 (O_119,N_16360,N_19476);
xnor UO_120 (O_120,N_16491,N_17805);
nor UO_121 (O_121,N_16921,N_19731);
and UO_122 (O_122,N_15293,N_16877);
nor UO_123 (O_123,N_19978,N_15976);
nand UO_124 (O_124,N_17139,N_16042);
nand UO_125 (O_125,N_16747,N_16817);
nor UO_126 (O_126,N_17594,N_16773);
nand UO_127 (O_127,N_19909,N_17623);
nor UO_128 (O_128,N_18839,N_16232);
nor UO_129 (O_129,N_18852,N_15135);
nand UO_130 (O_130,N_19999,N_15424);
nor UO_131 (O_131,N_16202,N_19849);
xor UO_132 (O_132,N_15573,N_18559);
or UO_133 (O_133,N_17802,N_16799);
and UO_134 (O_134,N_17636,N_17856);
nor UO_135 (O_135,N_15782,N_17138);
nand UO_136 (O_136,N_17453,N_18518);
or UO_137 (O_137,N_19165,N_16936);
nor UO_138 (O_138,N_17190,N_17000);
and UO_139 (O_139,N_18703,N_15785);
nand UO_140 (O_140,N_19315,N_18190);
nand UO_141 (O_141,N_15711,N_19436);
nand UO_142 (O_142,N_18011,N_17079);
nor UO_143 (O_143,N_18830,N_19200);
or UO_144 (O_144,N_16134,N_17911);
nor UO_145 (O_145,N_16871,N_15699);
nand UO_146 (O_146,N_18069,N_17953);
xnor UO_147 (O_147,N_16978,N_15260);
or UO_148 (O_148,N_15212,N_17848);
nand UO_149 (O_149,N_19630,N_16961);
nand UO_150 (O_150,N_16624,N_18030);
and UO_151 (O_151,N_17722,N_17258);
or UO_152 (O_152,N_19552,N_17390);
nand UO_153 (O_153,N_17358,N_19182);
nand UO_154 (O_154,N_17967,N_16862);
and UO_155 (O_155,N_19875,N_17431);
nand UO_156 (O_156,N_16509,N_16501);
nand UO_157 (O_157,N_15993,N_19897);
or UO_158 (O_158,N_19175,N_16288);
and UO_159 (O_159,N_15651,N_17929);
or UO_160 (O_160,N_17626,N_17646);
xor UO_161 (O_161,N_17306,N_16841);
xor UO_162 (O_162,N_16079,N_15796);
and UO_163 (O_163,N_19636,N_16868);
nor UO_164 (O_164,N_19449,N_17416);
or UO_165 (O_165,N_15141,N_17164);
and UO_166 (O_166,N_19146,N_18342);
or UO_167 (O_167,N_18194,N_18664);
and UO_168 (O_168,N_19820,N_17314);
and UO_169 (O_169,N_16448,N_19864);
or UO_170 (O_170,N_16802,N_18955);
nor UO_171 (O_171,N_17154,N_16241);
and UO_172 (O_172,N_18427,N_18898);
nor UO_173 (O_173,N_17531,N_19268);
nor UO_174 (O_174,N_18794,N_17940);
nand UO_175 (O_175,N_18279,N_15601);
xnor UO_176 (O_176,N_15556,N_15091);
nor UO_177 (O_177,N_18777,N_18019);
xor UO_178 (O_178,N_17886,N_19941);
and UO_179 (O_179,N_15491,N_16701);
xor UO_180 (O_180,N_17662,N_18552);
and UO_181 (O_181,N_15754,N_17447);
nand UO_182 (O_182,N_16245,N_16714);
and UO_183 (O_183,N_19631,N_19356);
xor UO_184 (O_184,N_18099,N_19621);
xor UO_185 (O_185,N_17415,N_16830);
nand UO_186 (O_186,N_16183,N_19904);
or UO_187 (O_187,N_18110,N_16056);
nor UO_188 (O_188,N_16043,N_15394);
and UO_189 (O_189,N_19027,N_19131);
or UO_190 (O_190,N_18423,N_17192);
and UO_191 (O_191,N_16858,N_17089);
xor UO_192 (O_192,N_19015,N_16801);
and UO_193 (O_193,N_16275,N_16842);
nor UO_194 (O_194,N_18887,N_15925);
and UO_195 (O_195,N_18845,N_19306);
and UO_196 (O_196,N_17420,N_17843);
or UO_197 (O_197,N_16726,N_16242);
nor UO_198 (O_198,N_17555,N_16780);
nor UO_199 (O_199,N_17015,N_16471);
and UO_200 (O_200,N_16172,N_16519);
and UO_201 (O_201,N_15783,N_15679);
nor UO_202 (O_202,N_16497,N_18798);
and UO_203 (O_203,N_17883,N_16573);
and UO_204 (O_204,N_19398,N_16195);
nor UO_205 (O_205,N_19725,N_16075);
xor UO_206 (O_206,N_18086,N_17821);
nand UO_207 (O_207,N_19123,N_19199);
or UO_208 (O_208,N_17224,N_18547);
and UO_209 (O_209,N_19405,N_18804);
and UO_210 (O_210,N_17509,N_16576);
nand UO_211 (O_211,N_17100,N_17203);
nor UO_212 (O_212,N_17868,N_16850);
xnor UO_213 (O_213,N_15935,N_17537);
or UO_214 (O_214,N_15447,N_18646);
nor UO_215 (O_215,N_19925,N_19384);
nor UO_216 (O_216,N_15612,N_17333);
nor UO_217 (O_217,N_15371,N_18343);
nor UO_218 (O_218,N_18551,N_16586);
or UO_219 (O_219,N_17146,N_17254);
and UO_220 (O_220,N_17432,N_19968);
nand UO_221 (O_221,N_19850,N_16510);
nand UO_222 (O_222,N_17903,N_17572);
and UO_223 (O_223,N_18161,N_19043);
nand UO_224 (O_224,N_15356,N_18519);
xnor UO_225 (O_225,N_15345,N_15561);
and UO_226 (O_226,N_19658,N_19775);
nor UO_227 (O_227,N_18482,N_16419);
or UO_228 (O_228,N_17220,N_18876);
nor UO_229 (O_229,N_16688,N_15518);
nand UO_230 (O_230,N_17579,N_15862);
and UO_231 (O_231,N_18449,N_15937);
or UO_232 (O_232,N_19557,N_18006);
and UO_233 (O_233,N_18152,N_15961);
nor UO_234 (O_234,N_16818,N_16331);
and UO_235 (O_235,N_17480,N_19450);
xnor UO_236 (O_236,N_19637,N_18486);
and UO_237 (O_237,N_15918,N_17941);
or UO_238 (O_238,N_17942,N_18940);
xor UO_239 (O_239,N_18358,N_16828);
and UO_240 (O_240,N_17632,N_15088);
nor UO_241 (O_241,N_16437,N_16080);
nor UO_242 (O_242,N_18394,N_17650);
nand UO_243 (O_243,N_15812,N_19150);
or UO_244 (O_244,N_17024,N_19908);
nor UO_245 (O_245,N_18347,N_19118);
and UO_246 (O_246,N_17408,N_16106);
nand UO_247 (O_247,N_15245,N_17062);
or UO_248 (O_248,N_18023,N_17135);
xor UO_249 (O_249,N_17150,N_18354);
and UO_250 (O_250,N_19838,N_15121);
nand UO_251 (O_251,N_15528,N_17691);
nor UO_252 (O_252,N_17282,N_18718);
or UO_253 (O_253,N_16439,N_18630);
and UO_254 (O_254,N_17445,N_16846);
or UO_255 (O_255,N_17144,N_17811);
and UO_256 (O_256,N_17645,N_18509);
nor UO_257 (O_257,N_16220,N_17859);
nand UO_258 (O_258,N_18866,N_17093);
and UO_259 (O_259,N_17174,N_16483);
or UO_260 (O_260,N_18277,N_19172);
or UO_261 (O_261,N_17864,N_15302);
or UO_262 (O_262,N_19163,N_17238);
nand UO_263 (O_263,N_19509,N_15641);
nor UO_264 (O_264,N_16024,N_17785);
or UO_265 (O_265,N_17905,N_17588);
or UO_266 (O_266,N_19525,N_19357);
or UO_267 (O_267,N_18971,N_15319);
and UO_268 (O_268,N_17344,N_18149);
nor UO_269 (O_269,N_18345,N_17030);
nand UO_270 (O_270,N_17397,N_19977);
or UO_271 (O_271,N_18314,N_15682);
or UO_272 (O_272,N_15664,N_17777);
nand UO_273 (O_273,N_18182,N_16813);
nor UO_274 (O_274,N_18123,N_15746);
xnor UO_275 (O_275,N_16292,N_17749);
and UO_276 (O_276,N_16757,N_17350);
xor UO_277 (O_277,N_15741,N_19489);
nand UO_278 (O_278,N_17807,N_18102);
xor UO_279 (O_279,N_15572,N_18439);
and UO_280 (O_280,N_16947,N_16348);
nand UO_281 (O_281,N_15763,N_18784);
nor UO_282 (O_282,N_18383,N_17155);
xor UO_283 (O_283,N_17710,N_18369);
xor UO_284 (O_284,N_19302,N_17659);
nand UO_285 (O_285,N_19305,N_18927);
and UO_286 (O_286,N_17092,N_18403);
xor UO_287 (O_287,N_15244,N_16998);
nand UO_288 (O_288,N_15483,N_19346);
nand UO_289 (O_289,N_18298,N_16416);
or UO_290 (O_290,N_15275,N_17747);
and UO_291 (O_291,N_18531,N_16005);
nand UO_292 (O_292,N_19821,N_19481);
xnor UO_293 (O_293,N_18679,N_19575);
and UO_294 (O_294,N_17892,N_15416);
and UO_295 (O_295,N_18272,N_19311);
xor UO_296 (O_296,N_16972,N_18827);
and UO_297 (O_297,N_15287,N_17219);
nor UO_298 (O_298,N_18032,N_15103);
nor UO_299 (O_299,N_17493,N_15510);
or UO_300 (O_300,N_18991,N_18478);
nor UO_301 (O_301,N_17614,N_19158);
or UO_302 (O_302,N_18649,N_17007);
or UO_303 (O_303,N_19811,N_15718);
or UO_304 (O_304,N_19454,N_15537);
or UO_305 (O_305,N_19529,N_19778);
nor UO_306 (O_306,N_18811,N_18132);
nand UO_307 (O_307,N_17809,N_18385);
nor UO_308 (O_308,N_19120,N_18931);
nand UO_309 (O_309,N_15737,N_16975);
nand UO_310 (O_310,N_19370,N_19570);
or UO_311 (O_311,N_16002,N_18037);
and UO_312 (O_312,N_16602,N_19526);
nand UO_313 (O_313,N_17775,N_15213);
or UO_314 (O_314,N_18027,N_16309);
xnor UO_315 (O_315,N_17675,N_19524);
xnor UO_316 (O_316,N_18134,N_18217);
nor UO_317 (O_317,N_17247,N_19816);
nand UO_318 (O_318,N_15061,N_19228);
or UO_319 (O_319,N_17198,N_16897);
and UO_320 (O_320,N_17326,N_17608);
nor UO_321 (O_321,N_19870,N_19781);
xor UO_322 (O_322,N_19966,N_15017);
nand UO_323 (O_323,N_19535,N_19886);
xor UO_324 (O_324,N_16776,N_18526);
nand UO_325 (O_325,N_17888,N_19303);
and UO_326 (O_326,N_16387,N_18140);
and UO_327 (O_327,N_16646,N_17370);
or UO_328 (O_328,N_15700,N_19061);
and UO_329 (O_329,N_16909,N_16110);
or UO_330 (O_330,N_19076,N_18606);
nand UO_331 (O_331,N_17251,N_16784);
xnor UO_332 (O_332,N_18489,N_16938);
xnor UO_333 (O_333,N_17399,N_18049);
or UO_334 (O_334,N_19500,N_17467);
xnor UO_335 (O_335,N_19056,N_18881);
xnor UO_336 (O_336,N_18332,N_17474);
or UO_337 (O_337,N_18558,N_18651);
nor UO_338 (O_338,N_17464,N_16383);
nor UO_339 (O_339,N_16770,N_15240);
nor UO_340 (O_340,N_15488,N_17386);
and UO_341 (O_341,N_19282,N_15997);
or UO_342 (O_342,N_16091,N_16582);
nand UO_343 (O_343,N_16789,N_15467);
nand UO_344 (O_344,N_16898,N_19736);
or UO_345 (O_345,N_16599,N_15881);
xnor UO_346 (O_346,N_18833,N_18713);
nand UO_347 (O_347,N_16382,N_19367);
nand UO_348 (O_348,N_16767,N_19766);
or UO_349 (O_349,N_19134,N_17462);
or UO_350 (O_350,N_15237,N_16107);
xor UO_351 (O_351,N_15665,N_17305);
nand UO_352 (O_352,N_15579,N_16652);
nor UO_353 (O_353,N_19609,N_16286);
nor UO_354 (O_354,N_16659,N_15716);
nor UO_355 (O_355,N_15723,N_17378);
nand UO_356 (O_356,N_18079,N_17653);
nand UO_357 (O_357,N_19154,N_15075);
xor UO_358 (O_358,N_16555,N_19666);
or UO_359 (O_359,N_19537,N_15396);
nor UO_360 (O_360,N_19375,N_16973);
or UO_361 (O_361,N_18131,N_16450);
xor UO_362 (O_362,N_16151,N_17217);
and UO_363 (O_363,N_17698,N_15800);
nor UO_364 (O_364,N_19815,N_19075);
or UO_365 (O_365,N_16375,N_16399);
nor UO_366 (O_366,N_16215,N_19596);
xor UO_367 (O_367,N_15032,N_17835);
nor UO_368 (O_368,N_19771,N_15125);
and UO_369 (O_369,N_16211,N_17793);
nand UO_370 (O_370,N_16154,N_17779);
xnor UO_371 (O_371,N_15703,N_19993);
and UO_372 (O_372,N_17229,N_16261);
or UO_373 (O_373,N_17652,N_18253);
xnor UO_374 (O_374,N_18842,N_16160);
nand UO_375 (O_375,N_16675,N_15740);
xor UO_376 (O_376,N_15325,N_16223);
nand UO_377 (O_377,N_18832,N_19624);
and UO_378 (O_378,N_19519,N_17392);
or UO_379 (O_379,N_17893,N_17564);
and UO_380 (O_380,N_18126,N_16690);
and UO_381 (O_381,N_16847,N_15369);
nor UO_382 (O_382,N_19170,N_18075);
nor UO_383 (O_383,N_15652,N_16230);
xor UO_384 (O_384,N_18870,N_18769);
nor UO_385 (O_385,N_15704,N_18850);
nor UO_386 (O_386,N_19536,N_15046);
and UO_387 (O_387,N_18108,N_19066);
xor UO_388 (O_388,N_15454,N_18492);
or UO_389 (O_389,N_17362,N_17409);
or UO_390 (O_390,N_16262,N_19413);
and UO_391 (O_391,N_18648,N_15972);
or UO_392 (O_392,N_19299,N_19916);
or UO_393 (O_393,N_15460,N_16627);
and UO_394 (O_394,N_16709,N_15252);
xnor UO_395 (O_395,N_15093,N_18460);
nand UO_396 (O_396,N_17484,N_18917);
xor UO_397 (O_397,N_18307,N_18490);
xor UO_398 (O_398,N_18618,N_17520);
and UO_399 (O_399,N_18252,N_18976);
and UO_400 (O_400,N_18501,N_19512);
and UO_401 (O_401,N_15522,N_15306);
or UO_402 (O_402,N_17186,N_18184);
or UO_403 (O_403,N_18377,N_15692);
nand UO_404 (O_404,N_15904,N_18637);
or UO_405 (O_405,N_16607,N_19924);
nor UO_406 (O_406,N_19180,N_18595);
xnor UO_407 (O_407,N_18109,N_19833);
or UO_408 (O_408,N_18062,N_18838);
and UO_409 (O_409,N_17438,N_19054);
nor UO_410 (O_410,N_15012,N_16617);
or UO_411 (O_411,N_19612,N_15629);
nor UO_412 (O_412,N_18259,N_16873);
nand UO_413 (O_413,N_18877,N_19579);
and UO_414 (O_414,N_17025,N_15562);
or UO_415 (O_415,N_15199,N_18410);
nand UO_416 (O_416,N_15734,N_19337);
xnor UO_417 (O_417,N_16994,N_15907);
or UO_418 (O_418,N_17348,N_16164);
or UO_419 (O_419,N_16906,N_17945);
nor UO_420 (O_420,N_19452,N_17609);
nand UO_421 (O_421,N_18384,N_17611);
xor UO_422 (O_422,N_15089,N_16953);
and UO_423 (O_423,N_17988,N_18523);
nand UO_424 (O_424,N_16677,N_16400);
nand UO_425 (O_425,N_15957,N_15967);
xor UO_426 (O_426,N_16775,N_16795);
nand UO_427 (O_427,N_15863,N_15571);
and UO_428 (O_428,N_18399,N_17357);
nor UO_429 (O_429,N_17271,N_19179);
or UO_430 (O_430,N_17371,N_16086);
or UO_431 (O_431,N_15831,N_18938);
and UO_432 (O_432,N_19005,N_15321);
and UO_433 (O_433,N_15818,N_16832);
and UO_434 (O_434,N_18116,N_15685);
or UO_435 (O_435,N_15045,N_16966);
or UO_436 (O_436,N_16664,N_17366);
xor UO_437 (O_437,N_15962,N_18414);
nor UO_438 (O_438,N_15638,N_19546);
or UO_439 (O_439,N_15466,N_16014);
and UO_440 (O_440,N_18943,N_18056);
xor UO_441 (O_441,N_15849,N_16809);
and UO_442 (O_442,N_16001,N_17185);
xor UO_443 (O_443,N_15544,N_18568);
or UO_444 (O_444,N_15081,N_15854);
nor UO_445 (O_445,N_17754,N_16074);
nand UO_446 (O_446,N_15706,N_18204);
nand UO_447 (O_447,N_19274,N_17745);
and UO_448 (O_448,N_16219,N_15382);
or UO_449 (O_449,N_16161,N_18306);
or UO_450 (O_450,N_16903,N_15404);
xor UO_451 (O_451,N_16284,N_16374);
xor UO_452 (O_452,N_17634,N_18783);
nand UO_453 (O_453,N_19205,N_19521);
nand UO_454 (O_454,N_15667,N_19402);
and UO_455 (O_455,N_17750,N_18819);
nand UO_456 (O_456,N_15539,N_15196);
nor UO_457 (O_457,N_16886,N_16385);
xor UO_458 (O_458,N_17435,N_19745);
nand UO_459 (O_459,N_18437,N_17442);
and UO_460 (O_460,N_19110,N_17161);
xor UO_461 (O_461,N_15719,N_15910);
and UO_462 (O_462,N_18304,N_17345);
and UO_463 (O_463,N_17310,N_17620);
or UO_464 (O_464,N_19258,N_19819);
nand UO_465 (O_465,N_19757,N_19243);
or UO_466 (O_466,N_18258,N_19892);
nor UO_467 (O_467,N_15549,N_18934);
xnor UO_468 (O_468,N_17506,N_19514);
nand UO_469 (O_469,N_16427,N_18456);
and UO_470 (O_470,N_17616,N_15847);
nor UO_471 (O_471,N_19955,N_18706);
or UO_472 (O_472,N_15949,N_15592);
and UO_473 (O_473,N_17915,N_15362);
xnor UO_474 (O_474,N_17980,N_17771);
xor UO_475 (O_475,N_17746,N_17126);
nor UO_476 (O_476,N_17695,N_15005);
and UO_477 (O_477,N_19871,N_18269);
and UO_478 (O_478,N_18781,N_16189);
and UO_479 (O_479,N_16463,N_18643);
and UO_480 (O_480,N_19349,N_17112);
nand UO_481 (O_481,N_17550,N_18335);
nor UO_482 (O_482,N_19652,N_15469);
nand UO_483 (O_483,N_19338,N_19458);
nor UO_484 (O_484,N_18546,N_16484);
nor UO_485 (O_485,N_18998,N_16955);
nor UO_486 (O_486,N_16453,N_19001);
nand UO_487 (O_487,N_17455,N_17987);
nor UO_488 (O_488,N_19988,N_16535);
nand UO_489 (O_489,N_18033,N_17773);
or UO_490 (O_490,N_17195,N_16143);
and UO_491 (O_491,N_17127,N_17958);
xor UO_492 (O_492,N_15026,N_18333);
nand UO_493 (O_493,N_17323,N_18951);
xor UO_494 (O_494,N_17796,N_16979);
xor UO_495 (O_495,N_19495,N_17393);
and UO_496 (O_496,N_17738,N_15870);
nand UO_497 (O_497,N_17273,N_15600);
and UO_498 (O_498,N_15662,N_16735);
xor UO_499 (O_499,N_19430,N_17813);
or UO_500 (O_500,N_15298,N_15894);
nand UO_501 (O_501,N_17119,N_19604);
or UO_502 (O_502,N_15303,N_16697);
xnor UO_503 (O_503,N_19606,N_19009);
nand UO_504 (O_504,N_15037,N_15411);
xnor UO_505 (O_505,N_18814,N_17851);
nand UO_506 (O_506,N_15414,N_15233);
and UO_507 (O_507,N_16849,N_16715);
xnor UO_508 (O_508,N_16939,N_15911);
or UO_509 (O_509,N_18266,N_19921);
and UO_510 (O_510,N_16486,N_17463);
nor UO_511 (O_511,N_18729,N_19973);
xor UO_512 (O_512,N_18324,N_17130);
nand UO_513 (O_513,N_17351,N_18973);
xor UO_514 (O_514,N_15258,N_18688);
or UO_515 (O_515,N_19396,N_18891);
nor UO_516 (O_516,N_17517,N_18135);
xnor UO_517 (O_517,N_16506,N_15959);
xor UO_518 (O_518,N_15047,N_19162);
nand UO_519 (O_519,N_16796,N_17648);
or UO_520 (O_520,N_16481,N_19159);
nor UO_521 (O_521,N_17256,N_17365);
and UO_522 (O_522,N_15691,N_18766);
and UO_523 (O_523,N_15124,N_15269);
xor UO_524 (O_524,N_19478,N_18848);
and UO_525 (O_525,N_16203,N_17159);
or UO_526 (O_526,N_18367,N_16132);
xnor UO_527 (O_527,N_19749,N_17989);
nand UO_528 (O_528,N_18301,N_17975);
nor UO_529 (O_529,N_16036,N_16199);
nand UO_530 (O_530,N_15550,N_19468);
xor UO_531 (O_531,N_19408,N_17402);
nand UO_532 (O_532,N_19720,N_16622);
nand UO_533 (O_533,N_16226,N_16983);
nor UO_534 (O_534,N_18319,N_18073);
nor UO_535 (O_535,N_19212,N_15128);
nand UO_536 (O_536,N_16155,N_18912);
and UO_537 (O_537,N_18294,N_19576);
nor UO_538 (O_538,N_19036,N_17922);
nand UO_539 (O_539,N_19855,N_15065);
nor UO_540 (O_540,N_18443,N_18496);
xor UO_541 (O_541,N_16520,N_17976);
xor UO_542 (O_542,N_15113,N_19744);
and UO_543 (O_543,N_15268,N_18901);
xor UO_544 (O_544,N_17901,N_19682);
nor UO_545 (O_545,N_19412,N_16698);
and UO_546 (O_546,N_15049,N_17867);
nand UO_547 (O_547,N_16512,N_16120);
nor UO_548 (O_548,N_19353,N_19880);
or UO_549 (O_549,N_15279,N_18953);
nand UO_550 (O_550,N_15238,N_15209);
and UO_551 (O_551,N_15627,N_18323);
and UO_552 (O_552,N_18747,N_19868);
nand UO_553 (O_553,N_15464,N_16674);
or UO_554 (O_554,N_15577,N_15106);
and UO_555 (O_555,N_15575,N_17448);
or UO_556 (O_556,N_16338,N_18010);
and UO_557 (O_557,N_17121,N_19292);
and UO_558 (O_558,N_16181,N_19010);
nor UO_559 (O_559,N_19035,N_17814);
nand UO_560 (O_560,N_16461,N_15825);
nand UO_561 (O_561,N_16639,N_17483);
and UO_562 (O_562,N_18522,N_19256);
or UO_563 (O_563,N_17436,N_18682);
or UO_564 (O_564,N_19835,N_15928);
xnor UO_565 (O_565,N_17346,N_16736);
or UO_566 (O_566,N_15297,N_16071);
nand UO_567 (O_567,N_19992,N_19181);
nor UO_568 (O_568,N_15402,N_17596);
nand UO_569 (O_569,N_19240,N_15946);
or UO_570 (O_570,N_15291,N_18710);
nor UO_571 (O_571,N_18990,N_19091);
or UO_572 (O_572,N_15519,N_16089);
and UO_573 (O_573,N_19153,N_15256);
nand UO_574 (O_574,N_18196,N_15410);
nor UO_575 (O_575,N_19696,N_18156);
nand UO_576 (O_576,N_17619,N_18540);
xor UO_577 (O_577,N_15285,N_16514);
or UO_578 (O_578,N_15377,N_15066);
nor UO_579 (O_579,N_18617,N_17374);
nor UO_580 (O_580,N_17101,N_18871);
nand UO_581 (O_581,N_17668,N_18422);
xnor UO_582 (O_582,N_18514,N_19129);
nor UO_583 (O_583,N_19157,N_16320);
and UO_584 (O_584,N_17456,N_15458);
xor UO_585 (O_585,N_16373,N_19828);
nor UO_586 (O_586,N_15457,N_19374);
or UO_587 (O_587,N_15038,N_17532);
or UO_588 (O_588,N_19271,N_16657);
nor UO_589 (O_589,N_17783,N_17065);
nand UO_590 (O_590,N_18441,N_17129);
xor UO_591 (O_591,N_18186,N_15618);
xnor UO_592 (O_592,N_16136,N_17457);
xnor UO_593 (O_593,N_18353,N_18334);
and UO_594 (O_594,N_15450,N_18061);
xor UO_595 (O_595,N_15606,N_19281);
or UO_596 (O_596,N_15018,N_15347);
nor UO_597 (O_597,N_15554,N_17658);
and UO_598 (O_598,N_18803,N_18031);
nand UO_599 (O_599,N_18318,N_17961);
and UO_600 (O_600,N_18130,N_15253);
xor UO_601 (O_601,N_19020,N_16312);
xnor UO_602 (O_602,N_16719,N_15363);
or UO_603 (O_603,N_19837,N_15950);
nand UO_604 (O_604,N_18229,N_18287);
nand UO_605 (O_605,N_16330,N_17897);
and UO_606 (O_606,N_17004,N_15840);
nor UO_607 (O_607,N_17959,N_17876);
and UO_608 (O_608,N_15117,N_15324);
nor UO_609 (O_609,N_15952,N_17476);
and UO_610 (O_610,N_18448,N_15234);
xnor UO_611 (O_611,N_15202,N_18137);
nor UO_612 (O_612,N_19318,N_19204);
and UO_613 (O_613,N_18281,N_17951);
nor UO_614 (O_614,N_18612,N_17152);
nor UO_615 (O_615,N_18533,N_19090);
or UO_616 (O_616,N_19710,N_17137);
nor UO_617 (O_617,N_16269,N_19543);
and UO_618 (O_618,N_15846,N_15218);
nand UO_619 (O_619,N_18059,N_19462);
nor UO_620 (O_620,N_15728,N_16587);
or UO_621 (O_621,N_18704,N_16815);
or UO_622 (O_622,N_17842,N_19112);
nor UO_623 (O_623,N_18732,N_16691);
xnor UO_624 (O_624,N_18549,N_16264);
or UO_625 (O_625,N_16378,N_18903);
or UO_626 (O_626,N_17799,N_18067);
or UO_627 (O_627,N_17689,N_17720);
xnor UO_628 (O_628,N_17369,N_17797);
xnor UO_629 (O_629,N_17672,N_15039);
nor UO_630 (O_630,N_19039,N_18735);
nor UO_631 (O_631,N_16390,N_16707);
or UO_632 (O_632,N_19278,N_15397);
xor UO_633 (O_633,N_15055,N_17028);
or UO_634 (O_634,N_16742,N_15514);
nand UO_635 (O_635,N_17836,N_16901);
nor UO_636 (O_636,N_15383,N_17712);
nor UO_637 (O_637,N_15936,N_15058);
and UO_638 (O_638,N_16141,N_16294);
nand UO_639 (O_639,N_16859,N_18689);
and UO_640 (O_640,N_19840,N_15193);
nor UO_641 (O_641,N_18942,N_17057);
or UO_642 (O_642,N_16857,N_15105);
nor UO_643 (O_643,N_19931,N_17635);
nor UO_644 (O_644,N_18026,N_16793);
or UO_645 (O_645,N_15008,N_15797);
and UO_646 (O_646,N_18401,N_19747);
or UO_647 (O_647,N_19903,N_17741);
or UO_648 (O_648,N_16984,N_15368);
or UO_649 (O_649,N_18273,N_16413);
and UO_650 (O_650,N_16518,N_16085);
or UO_651 (O_651,N_15336,N_17414);
nand UO_652 (O_652,N_19586,N_16508);
or UO_653 (O_653,N_19601,N_18212);
nor UO_654 (O_654,N_18890,N_15229);
nand UO_655 (O_655,N_15358,N_16642);
nor UO_656 (O_656,N_18530,N_17269);
nand UO_657 (O_657,N_17534,N_19826);
nand UO_658 (O_658,N_19613,N_19049);
and UO_659 (O_659,N_18093,N_18265);
xor UO_660 (O_660,N_15249,N_15418);
xor UO_661 (O_661,N_19189,N_18621);
nor UO_662 (O_662,N_19208,N_15978);
and UO_663 (O_663,N_17486,N_15670);
xnor UO_664 (O_664,N_19812,N_16515);
nand UO_665 (O_665,N_15595,N_16050);
and UO_666 (O_666,N_15987,N_17218);
nand UO_667 (O_667,N_19445,N_18256);
nand UO_668 (O_668,N_17514,N_19383);
nor UO_669 (O_669,N_17914,N_15547);
xnor UO_670 (O_670,N_17487,N_19595);
or UO_671 (O_671,N_16418,N_19520);
and UO_672 (O_672,N_16123,N_17968);
and UO_673 (O_673,N_19480,N_15380);
and UO_674 (O_674,N_16571,N_18763);
or UO_675 (O_675,N_17728,N_19293);
xnor UO_676 (O_676,N_19422,N_15909);
xor UO_677 (O_677,N_17740,N_18650);
and UO_678 (O_678,N_17473,N_16462);
xnor UO_679 (O_679,N_16073,N_17010);
nand UO_680 (O_680,N_15512,N_18981);
and UO_681 (O_681,N_19627,N_15778);
nand UO_682 (O_682,N_18210,N_16502);
or UO_683 (O_683,N_19249,N_18691);
or UO_684 (O_684,N_16748,N_18446);
and UO_685 (O_685,N_15666,N_15674);
and UO_686 (O_686,N_19312,N_15774);
nor UO_687 (O_687,N_15272,N_17047);
and UO_688 (O_688,N_19028,N_16169);
xnor UO_689 (O_689,N_19272,N_15151);
and UO_690 (O_690,N_16325,N_16435);
nor UO_691 (O_691,N_15087,N_16217);
nor UO_692 (O_692,N_18677,N_17600);
or UO_693 (O_693,N_16140,N_15861);
nand UO_694 (O_694,N_15111,N_16152);
nor UO_695 (O_695,N_19729,N_19960);
nand UO_696 (O_696,N_19152,N_17311);
nor UO_697 (O_697,N_18640,N_16574);
or UO_698 (O_698,N_16304,N_15628);
and UO_699 (O_699,N_19106,N_18235);
or UO_700 (O_700,N_16671,N_16750);
or UO_701 (O_701,N_16221,N_16589);
xor UO_702 (O_702,N_15343,N_18487);
nor UO_703 (O_703,N_15932,N_15599);
or UO_704 (O_704,N_15323,N_19395);
xnor UO_705 (O_705,N_16369,N_16824);
xnor UO_706 (O_706,N_19308,N_17589);
nand UO_707 (O_707,N_18320,N_18100);
nand UO_708 (O_708,N_18695,N_18183);
nor UO_709 (O_709,N_19214,N_18722);
and UO_710 (O_710,N_15570,N_16334);
and UO_711 (O_711,N_15955,N_16166);
nand UO_712 (O_712,N_15790,N_19477);
nand UO_713 (O_713,N_17936,N_17250);
and UO_714 (O_714,N_19703,N_16612);
nand UO_715 (O_715,N_16090,N_19264);
nor UO_716 (O_716,N_18736,N_16620);
nand UO_717 (O_717,N_16608,N_16825);
and UO_718 (O_718,N_17513,N_16493);
or UO_719 (O_719,N_19578,N_15431);
xnor UO_720 (O_720,N_19608,N_19964);
nor UO_721 (O_721,N_17325,N_16266);
nand UO_722 (O_722,N_18734,N_19597);
xor UO_723 (O_723,N_18762,N_16762);
and UO_724 (O_724,N_16306,N_15832);
nand UO_725 (O_725,N_16310,N_15221);
xor UO_726 (O_726,N_17628,N_18963);
and UO_727 (O_727,N_18669,N_15143);
or UO_728 (O_728,N_16760,N_19330);
or UO_729 (O_729,N_16206,N_18344);
or UO_730 (O_730,N_16783,N_18476);
xor UO_731 (O_731,N_18378,N_19994);
nand UO_732 (O_732,N_17637,N_15793);
nor UO_733 (O_733,N_19810,N_19280);
and UO_734 (O_734,N_18106,N_16167);
or UO_735 (O_735,N_19972,N_18537);
nor UO_736 (O_736,N_15673,N_18162);
xnor UO_737 (O_737,N_19138,N_18166);
nor UO_738 (O_738,N_16996,N_19976);
nor UO_739 (O_739,N_15697,N_18153);
and UO_740 (O_740,N_18060,N_16367);
nand UO_741 (O_741,N_19332,N_17977);
xor UO_742 (O_742,N_19244,N_18171);
nand UO_743 (O_743,N_17048,N_17204);
nor UO_744 (O_744,N_19327,N_17902);
nor UO_745 (O_745,N_16637,N_17870);
nand UO_746 (O_746,N_17206,N_15413);
nor UO_747 (O_747,N_18907,N_16389);
or UO_748 (O_748,N_15455,N_18816);
or UO_749 (O_749,N_18286,N_17160);
xnor UO_750 (O_750,N_19888,N_17496);
nand UO_751 (O_751,N_19753,N_19410);
and UO_752 (O_752,N_16173,N_15180);
or UO_753 (O_753,N_19217,N_18668);
or UO_754 (O_754,N_17776,N_17770);
nand UO_755 (O_755,N_18363,N_17827);
and UO_756 (O_756,N_15408,N_19155);
nand UO_757 (O_757,N_18261,N_18303);
nor UO_758 (O_758,N_18635,N_17955);
and UO_759 (O_759,N_18242,N_15806);
nor UO_760 (O_760,N_17136,N_18224);
nor UO_761 (O_761,N_19926,N_19692);
nor UO_762 (O_762,N_19373,N_17546);
nand UO_763 (O_763,N_15759,N_15201);
nor UO_764 (O_764,N_16423,N_19233);
xnor UO_765 (O_765,N_18582,N_19130);
nand UO_766 (O_766,N_17979,N_16872);
xnor UO_767 (O_767,N_19752,N_17272);
nor UO_768 (O_768,N_15581,N_19084);
xnor UO_769 (O_769,N_19975,N_16287);
or UO_770 (O_770,N_19492,N_15056);
or UO_771 (O_771,N_15698,N_19640);
or UO_772 (O_772,N_16654,N_16733);
xnor UO_773 (O_773,N_18930,N_17787);
nor UO_774 (O_774,N_18944,N_19059);
nor UO_775 (O_775,N_18536,N_18663);
nand UO_776 (O_776,N_16579,N_17622);
and UO_777 (O_777,N_18278,N_18882);
xnor UO_778 (O_778,N_19246,N_19260);
xnor UO_779 (O_779,N_17477,N_19196);
or UO_780 (O_780,N_19379,N_18292);
xnor UO_781 (O_781,N_19853,N_19143);
and UO_782 (O_782,N_18268,N_17299);
xnor UO_783 (O_783,N_19754,N_19085);
nor UO_784 (O_784,N_19467,N_18090);
or UO_785 (O_785,N_18593,N_18505);
nor UO_786 (O_786,N_18255,N_18563);
nand UO_787 (O_787,N_18864,N_18909);
xor UO_788 (O_788,N_18957,N_16239);
nor UO_789 (O_789,N_15749,N_19502);
nand UO_790 (O_790,N_15789,N_18658);
nor UO_791 (O_791,N_15984,N_19698);
or UO_792 (O_792,N_16663,N_17918);
nand UO_793 (O_793,N_18232,N_16208);
nor UO_794 (O_794,N_19475,N_19709);
nand UO_795 (O_795,N_17303,N_16082);
xor UO_796 (O_796,N_15499,N_19750);
nor UO_797 (O_797,N_19026,N_16951);
nand UO_798 (O_798,N_17525,N_16398);
or UO_799 (O_799,N_17418,N_19171);
nor UO_800 (O_800,N_19530,N_17804);
xnor UO_801 (O_801,N_18216,N_19767);
nor UO_802 (O_802,N_16592,N_15247);
xnor UO_803 (O_803,N_17759,N_19560);
nor UO_804 (O_804,N_16267,N_17717);
xnor UO_805 (O_805,N_16908,N_15420);
and UO_806 (O_806,N_16771,N_18283);
and UO_807 (O_807,N_19922,N_18916);
nor UO_808 (O_808,N_16557,N_17504);
nand UO_809 (O_809,N_19806,N_16563);
xnor UO_810 (O_810,N_18556,N_17845);
and UO_811 (O_811,N_17544,N_16907);
and UO_812 (O_812,N_16614,N_15025);
nor UO_813 (O_813,N_15054,N_19072);
and UO_814 (O_814,N_19646,N_16363);
and UO_815 (O_815,N_17688,N_17577);
and UO_816 (O_816,N_18472,N_16718);
xor UO_817 (O_817,N_16803,N_19080);
nor UO_818 (O_818,N_15552,N_18761);
xor UO_819 (O_819,N_16982,N_15817);
xor UO_820 (O_820,N_15211,N_17937);
and UO_821 (O_821,N_17151,N_17163);
nand UO_822 (O_822,N_17016,N_15788);
and UO_823 (O_823,N_16218,N_15333);
xor UO_824 (O_824,N_16470,N_16712);
and UO_825 (O_825,N_19394,N_15619);
or UO_826 (O_826,N_16345,N_19951);
nand UO_827 (O_827,N_19564,N_18007);
xnor UO_828 (O_828,N_15426,N_17116);
or UO_829 (O_829,N_16534,N_15611);
or UO_830 (O_830,N_19429,N_19469);
nand UO_831 (O_831,N_15650,N_15567);
nor UO_832 (O_832,N_17073,N_19291);
nand UO_833 (O_833,N_19858,N_15316);
nand UO_834 (O_834,N_15184,N_19588);
xnor UO_835 (O_835,N_16516,N_15332);
xnor UO_836 (O_836,N_18584,N_19194);
or UO_837 (O_837,N_15028,N_18918);
xor UO_838 (O_838,N_19759,N_15634);
or UO_839 (O_839,N_16711,N_18778);
xnor UO_840 (O_840,N_17367,N_15934);
and UO_841 (O_841,N_18128,N_17286);
nor UO_842 (O_842,N_17424,N_15640);
nor UO_843 (O_843,N_18873,N_17761);
or UO_844 (O_844,N_15295,N_17231);
nand UO_845 (O_845,N_15485,N_15178);
nand UO_846 (O_846,N_18267,N_19600);
nor UO_847 (O_847,N_19795,N_19987);
xnor UO_848 (O_848,N_15053,N_15086);
nand UO_849 (O_849,N_18238,N_16000);
and UO_850 (O_850,N_19648,N_15744);
nand UO_851 (O_851,N_15079,N_16034);
nor UO_852 (O_852,N_18774,N_15036);
xor UO_853 (O_853,N_15386,N_16756);
or UO_854 (O_854,N_16393,N_19314);
nor UO_855 (O_855,N_19057,N_19653);
nor UO_856 (O_856,N_16561,N_18498);
xor UO_857 (O_857,N_18555,N_19829);
and UO_858 (O_858,N_16618,N_17714);
or UO_859 (O_859,N_16335,N_16028);
nand UO_860 (O_860,N_16554,N_18857);
or UO_861 (O_861,N_18936,N_19300);
or UO_862 (O_862,N_15877,N_17255);
nor UO_863 (O_863,N_17124,N_15009);
xor UO_864 (O_864,N_19527,N_17739);
and UO_865 (O_865,N_15517,N_16710);
and UO_866 (O_866,N_17142,N_19433);
and UO_867 (O_867,N_15622,N_16687);
xnor UO_868 (O_868,N_18039,N_17673);
or UO_869 (O_869,N_19187,N_15644);
or UO_870 (O_870,N_18680,N_18897);
nand UO_871 (O_871,N_17363,N_16603);
nand UO_872 (O_872,N_17221,N_17235);
nor UO_873 (O_873,N_18096,N_18600);
nor UO_874 (O_874,N_16408,N_15299);
or UO_875 (O_875,N_19400,N_15011);
and UO_876 (O_876,N_17789,N_18198);
nand UO_877 (O_877,N_18158,N_18296);
and UO_878 (O_878,N_19611,N_16882);
nand UO_879 (O_879,N_17304,N_17638);
xor UO_880 (O_880,N_17417,N_16210);
nand UO_881 (O_881,N_18425,N_19178);
nor UO_882 (O_882,N_15434,N_19505);
and UO_883 (O_883,N_15929,N_15232);
and UO_884 (O_884,N_15884,N_16455);
xor UO_885 (O_885,N_18101,N_19760);
nand UO_886 (O_886,N_15864,N_18391);
nor UO_887 (O_887,N_18189,N_15078);
xnor UO_888 (O_888,N_17970,N_16163);
xnor UO_889 (O_889,N_16426,N_15352);
xor UO_890 (O_890,N_18755,N_15083);
nand UO_891 (O_891,N_18661,N_15243);
nand UO_892 (O_892,N_15762,N_19679);
xnor UO_893 (O_893,N_17732,N_16362);
nand UO_894 (O_894,N_15945,N_18200);
and UO_895 (O_895,N_15610,N_15158);
nor UO_896 (O_896,N_17296,N_16943);
or UO_897 (O_897,N_18929,N_15912);
or UO_898 (O_898,N_17289,N_16727);
or UO_899 (O_899,N_19683,N_15288);
xor UO_900 (O_900,N_19531,N_17018);
and UO_901 (O_901,N_17894,N_18406);
nor UO_902 (O_902,N_15776,N_19733);
nor UO_903 (O_903,N_16204,N_18020);
xnor UO_904 (O_904,N_15974,N_19632);
xnor UO_905 (O_905,N_16317,N_17294);
xor UO_906 (O_906,N_19004,N_18701);
nor UO_907 (O_907,N_19532,N_19025);
xor UO_908 (O_908,N_19431,N_18660);
and UO_909 (O_909,N_17713,N_19674);
and UO_910 (O_910,N_19340,N_18094);
xor UO_911 (O_911,N_17459,N_19563);
nand UO_912 (O_912,N_18312,N_19414);
nor UO_913 (O_913,N_16323,N_17815);
nand UO_914 (O_914,N_17935,N_18579);
nor UO_915 (O_915,N_18880,N_19738);
nand UO_916 (O_916,N_17995,N_18438);
nor UO_917 (O_917,N_18675,N_15470);
nor UO_918 (O_918,N_16840,N_16649);
and UO_919 (O_919,N_15421,N_17316);
xor UO_920 (O_920,N_19559,N_18702);
nor UO_921 (O_921,N_15980,N_16808);
xnor UO_922 (O_922,N_19466,N_19697);
or UO_923 (O_923,N_18904,N_16918);
or UO_924 (O_924,N_15717,N_16621);
and UO_925 (O_925,N_16804,N_19496);
or UO_926 (O_926,N_15101,N_15236);
and UO_927 (O_927,N_19770,N_19298);
and UO_928 (O_928,N_17082,N_15085);
xor UO_929 (O_929,N_16807,N_16878);
nand UO_930 (O_930,N_18571,N_17500);
nand UO_931 (O_931,N_16593,N_15290);
or UO_932 (O_932,N_15335,N_19539);
xor UO_933 (O_933,N_19856,N_19499);
nand UO_934 (O_934,N_18491,N_17064);
or UO_935 (O_935,N_18357,N_19561);
xor UO_936 (O_936,N_15558,N_19695);
nor UO_937 (O_937,N_15835,N_15656);
or UO_938 (O_938,N_15374,N_16755);
nand UO_939 (O_939,N_15021,N_17189);
and UO_940 (O_940,N_17960,N_15676);
nand UO_941 (O_941,N_17890,N_19136);
xor UO_942 (O_942,N_18066,N_15165);
or UO_943 (O_943,N_15659,N_17242);
nand UO_944 (O_944,N_16032,N_19508);
nor UO_945 (O_945,N_18201,N_19464);
nor UO_946 (O_946,N_15484,N_16359);
xnor UO_947 (O_947,N_15261,N_15696);
and UO_948 (O_948,N_16960,N_16884);
xnor UO_949 (O_949,N_17439,N_15157);
or UO_950 (O_950,N_16848,N_16104);
and UO_951 (O_951,N_18696,N_16128);
and UO_952 (O_952,N_18996,N_19907);
xnor UO_953 (O_953,N_19748,N_16396);
or UO_954 (O_954,N_17022,N_18510);
xor UO_955 (O_955,N_16786,N_16404);
xor UO_956 (O_956,N_19177,N_18036);
nand UO_957 (O_957,N_16403,N_15889);
and UO_958 (O_958,N_19362,N_16891);
or UO_959 (O_959,N_17468,N_15906);
or UO_960 (O_960,N_16948,N_17681);
nor UO_961 (O_961,N_16271,N_17751);
and UO_962 (O_962,N_16498,N_19250);
nand UO_963 (O_963,N_17342,N_19320);
nor UO_964 (O_964,N_15100,N_15219);
nand UO_965 (O_965,N_15775,N_15405);
and UO_966 (O_966,N_19203,N_16022);
nor UO_967 (O_967,N_19190,N_18084);
and UO_968 (O_968,N_18855,N_15505);
and UO_969 (O_969,N_18119,N_15092);
and UO_970 (O_970,N_18115,N_19459);
and UO_971 (O_971,N_15205,N_15489);
nand UO_972 (O_972,N_18822,N_15446);
xnor UO_973 (O_973,N_17180,N_15094);
nor UO_974 (O_974,N_19050,N_15381);
nor UO_975 (O_975,N_17153,N_15551);
nand UO_976 (O_976,N_16670,N_17389);
and UO_977 (O_977,N_15400,N_18768);
xor UO_978 (O_978,N_18222,N_16158);
xnor UO_979 (O_979,N_15015,N_18453);
nand UO_980 (O_980,N_15617,N_17539);
xnor UO_981 (O_981,N_17898,N_18418);
or UO_982 (O_982,N_19407,N_18231);
nand UO_983 (O_983,N_16395,N_17930);
or UO_984 (O_984,N_15883,N_19497);
nand UO_985 (O_985,N_15482,N_19876);
nand UO_986 (O_986,N_16411,N_15895);
nand UO_987 (O_987,N_17706,N_15341);
nor UO_988 (O_988,N_18008,N_17169);
and UO_989 (O_989,N_19844,N_18471);
or UO_990 (O_990,N_16703,N_15071);
nand UO_991 (O_991,N_15543,N_17077);
xor UO_992 (O_992,N_15137,N_15865);
and UO_993 (O_993,N_17838,N_17410);
and UO_994 (O_994,N_16078,N_17215);
and UO_995 (O_995,N_18241,N_19368);
xor UO_996 (O_996,N_18779,N_17071);
nand UO_997 (O_997,N_15441,N_17332);
nor UO_998 (O_998,N_16610,N_15331);
and UO_999 (O_999,N_16702,N_16685);
xor UO_1000 (O_1000,N_17090,N_18539);
nor UO_1001 (O_1001,N_17200,N_19676);
or UO_1002 (O_1002,N_19290,N_16546);
or UO_1003 (O_1003,N_15387,N_19418);
and UO_1004 (O_1004,N_17946,N_19209);
nand UO_1005 (O_1005,N_18234,N_15436);
nor UO_1006 (O_1006,N_16792,N_18208);
xnor UO_1007 (O_1007,N_18731,N_15177);
nor UO_1008 (O_1008,N_18074,N_17384);
nand UO_1009 (O_1009,N_18035,N_15583);
xor UO_1010 (O_1010,N_17226,N_17680);
nand UO_1011 (O_1011,N_18495,N_17005);
nand UO_1012 (O_1012,N_18257,N_16990);
or UO_1013 (O_1013,N_17592,N_19382);
and UO_1014 (O_1014,N_16099,N_18395);
nor UO_1015 (O_1015,N_15442,N_18997);
or UO_1016 (O_1016,N_15393,N_15433);
and UO_1017 (O_1017,N_18608,N_18068);
nand UO_1018 (O_1018,N_17808,N_18170);
nand UO_1019 (O_1019,N_16253,N_17411);
xnor UO_1020 (O_1020,N_19037,N_18178);
xor UO_1021 (O_1021,N_19494,N_18029);
nor UO_1022 (O_1022,N_16914,N_16384);
xnor UO_1023 (O_1023,N_15553,N_17337);
nor UO_1024 (O_1024,N_16785,N_16541);
nor UO_1025 (O_1025,N_18538,N_17099);
nand UO_1026 (O_1026,N_17508,N_19934);
and UO_1027 (O_1027,N_16894,N_15156);
and UO_1028 (O_1028,N_15933,N_17315);
nor UO_1029 (O_1029,N_19236,N_19540);
and UO_1030 (O_1030,N_17629,N_15828);
xnor UO_1031 (O_1031,N_18905,N_15999);
xnor UO_1032 (O_1032,N_19098,N_18674);
nand UO_1033 (O_1033,N_18694,N_19008);
nand UO_1034 (O_1034,N_16259,N_16246);
nor UO_1035 (O_1035,N_17563,N_15034);
and UO_1036 (O_1036,N_18185,N_15977);
xnor UO_1037 (O_1037,N_15948,N_18854);
xnor UO_1038 (O_1038,N_15175,N_15471);
and UO_1039 (O_1039,N_15888,N_19681);
xnor UO_1040 (O_1040,N_17527,N_19465);
or UO_1041 (O_1041,N_16929,N_17441);
xnor UO_1042 (O_1042,N_16811,N_18993);
or UO_1043 (O_1043,N_16102,N_18681);
nor UO_1044 (O_1044,N_19642,N_17049);
or UO_1045 (O_1045,N_17469,N_17828);
xor UO_1046 (O_1046,N_15152,N_19997);
nor UO_1047 (O_1047,N_17216,N_18432);
nand UO_1048 (O_1048,N_17427,N_18451);
nand UO_1049 (O_1049,N_17381,N_18910);
nand UO_1050 (O_1050,N_18226,N_19404);
nand UO_1051 (O_1051,N_18147,N_18177);
nor UO_1052 (O_1052,N_17492,N_17536);
or UO_1053 (O_1053,N_15492,N_15751);
nor UO_1054 (O_1054,N_18773,N_15266);
xor UO_1055 (O_1055,N_19573,N_16349);
or UO_1056 (O_1056,N_15756,N_15116);
xnor UO_1057 (O_1057,N_16744,N_17816);
nor UO_1058 (O_1058,N_15474,N_15104);
and UO_1059 (O_1059,N_19142,N_18052);
and UO_1060 (O_1060,N_15780,N_17853);
and UO_1061 (O_1061,N_15695,N_16477);
nand UO_1062 (O_1062,N_16679,N_16440);
nor UO_1063 (O_1063,N_18125,N_19116);
or UO_1064 (O_1064,N_17063,N_15392);
xor UO_1065 (O_1065,N_15502,N_18911);
nor UO_1066 (O_1066,N_15326,N_15251);
and UO_1067 (O_1067,N_15752,N_15144);
nand UO_1068 (O_1068,N_17565,N_15148);
and UO_1069 (O_1069,N_16580,N_16182);
nand UO_1070 (O_1070,N_16769,N_17162);
or UO_1071 (O_1071,N_19568,N_18844);
nor UO_1072 (O_1072,N_19044,N_19147);
xnor UO_1073 (O_1073,N_18984,N_16797);
nor UO_1074 (O_1074,N_15278,N_19016);
nand UO_1075 (O_1075,N_19485,N_15023);
xnor UO_1076 (O_1076,N_18442,N_16178);
nor UO_1077 (O_1077,N_18639,N_19550);
nand UO_1078 (O_1078,N_19077,N_18337);
nand UO_1079 (O_1079,N_19761,N_19774);
or UO_1080 (O_1080,N_18215,N_16095);
nor UO_1081 (O_1081,N_19776,N_17679);
or UO_1082 (O_1082,N_19797,N_19789);
and UO_1083 (O_1083,N_15203,N_17602);
nand UO_1084 (O_1084,N_19276,N_18575);
nand UO_1085 (O_1085,N_19574,N_17426);
xor UO_1086 (O_1086,N_19912,N_17283);
and UO_1087 (O_1087,N_15048,N_16240);
xor UO_1088 (O_1088,N_17131,N_15810);
or UO_1089 (O_1089,N_17277,N_15379);
xor UO_1090 (O_1090,N_18719,N_17981);
nor UO_1091 (O_1091,N_16256,N_16604);
nand UO_1092 (O_1092,N_15971,N_18028);
nor UO_1093 (O_1093,N_16125,N_17552);
nor UO_1094 (O_1094,N_16542,N_19585);
and UO_1095 (O_1095,N_17655,N_19701);
nor UO_1096 (O_1096,N_15027,N_17599);
or UO_1097 (O_1097,N_17639,N_16749);
nand UO_1098 (O_1098,N_16017,N_19511);
and UO_1099 (O_1099,N_18169,N_19425);
and UO_1100 (O_1100,N_17693,N_18862);
nand UO_1101 (O_1101,N_18018,N_18790);
and UO_1102 (O_1102,N_16944,N_16119);
nor UO_1103 (O_1103,N_17541,N_16305);
nor UO_1104 (O_1104,N_18921,N_19732);
or UO_1105 (O_1105,N_19798,N_18463);
xor UO_1106 (O_1106,N_17511,N_15689);
nand UO_1107 (O_1107,N_18081,N_16725);
nand UO_1108 (O_1108,N_17965,N_15853);
nor UO_1109 (O_1109,N_19714,N_16851);
and UO_1110 (O_1110,N_17281,N_17395);
xnor UO_1111 (O_1111,N_16029,N_19665);
nor UO_1112 (O_1112,N_18133,N_16791);
xor UO_1113 (O_1113,N_18293,N_19948);
xor UO_1114 (O_1114,N_19773,N_17404);
nand UO_1115 (O_1115,N_15969,N_17569);
nor UO_1116 (O_1116,N_16444,N_19023);
or UO_1117 (O_1117,N_18249,N_16458);
and UO_1118 (O_1118,N_16315,N_15159);
xor UO_1119 (O_1119,N_17928,N_16577);
nor UO_1120 (O_1120,N_19723,N_16523);
or UO_1121 (O_1121,N_19804,N_17491);
nor UO_1122 (O_1122,N_16704,N_15766);
nor UO_1123 (O_1123,N_18118,N_16625);
nand UO_1124 (O_1124,N_16431,N_15559);
xor UO_1125 (O_1125,N_18408,N_15850);
xor UO_1126 (O_1126,N_18676,N_17263);
nand UO_1127 (O_1127,N_18624,N_16357);
xor UO_1128 (O_1128,N_15805,N_17298);
nor UO_1129 (O_1129,N_19898,N_19135);
nand UO_1130 (O_1130,N_19266,N_16992);
or UO_1131 (O_1131,N_18987,N_16794);
nand UO_1132 (O_1132,N_18005,N_15898);
or UO_1133 (O_1133,N_18569,N_17505);
nor UO_1134 (O_1134,N_16572,N_16740);
xnor UO_1135 (O_1135,N_17810,N_18826);
xor UO_1136 (O_1136,N_16111,N_16616);
and UO_1137 (O_1137,N_17264,N_17615);
and UO_1138 (O_1138,N_19380,N_16539);
or UO_1139 (O_1139,N_15207,N_18154);
xnor UO_1140 (O_1140,N_17194,N_17102);
and UO_1141 (O_1141,N_19986,N_19620);
nor UO_1142 (O_1142,N_16902,N_19786);
or UO_1143 (O_1143,N_15900,N_16694);
or UO_1144 (O_1144,N_17379,N_16781);
or UO_1145 (O_1145,N_19191,N_17764);
and UO_1146 (O_1146,N_16234,N_17122);
xnor UO_1147 (O_1147,N_18828,N_18014);
or UO_1148 (O_1148,N_15099,N_19783);
or UO_1149 (O_1149,N_15226,N_15425);
xnor UO_1150 (O_1150,N_15892,N_19487);
nor UO_1151 (O_1151,N_17268,N_17078);
xor UO_1152 (O_1152,N_19041,N_15167);
nand UO_1153 (O_1153,N_16115,N_17803);
xnor UO_1154 (O_1154,N_16971,N_15378);
xor UO_1155 (O_1155,N_17507,N_17425);
nand UO_1156 (O_1156,N_17690,N_17145);
nand UO_1157 (O_1157,N_17499,N_16696);
nor UO_1158 (O_1158,N_18348,N_16934);
and UO_1159 (O_1159,N_18992,N_17270);
or UO_1160 (O_1160,N_16301,N_16096);
nor UO_1161 (O_1161,N_18548,N_17974);
nand UO_1162 (O_1162,N_18528,N_16601);
and UO_1163 (O_1163,N_15688,N_15623);
nand UO_1164 (O_1164,N_18206,N_19401);
nor UO_1165 (O_1165,N_18381,N_19655);
and UO_1166 (O_1166,N_19046,N_16145);
and UO_1167 (O_1167,N_19392,N_18878);
nor UO_1168 (O_1168,N_16536,N_16238);
nor UO_1169 (O_1169,N_19887,N_17001);
or UO_1170 (O_1170,N_18129,N_16889);
and UO_1171 (O_1171,N_18802,N_18513);
nand UO_1172 (O_1172,N_19558,N_17701);
nand UO_1173 (O_1173,N_18561,N_17489);
or UO_1174 (O_1174,N_18858,N_18820);
nor UO_1175 (O_1175,N_18570,N_15496);
xor UO_1176 (O_1176,N_17278,N_18683);
or UO_1177 (O_1177,N_18670,N_17860);
nand UO_1178 (O_1178,N_16782,N_17966);
nand UO_1179 (O_1179,N_16475,N_19743);
or UO_1180 (O_1180,N_19148,N_16329);
and UO_1181 (O_1181,N_16131,N_18527);
and UO_1182 (O_1182,N_16489,N_17840);
and UO_1183 (O_1183,N_18288,N_19788);
or UO_1184 (O_1184,N_15930,N_15905);
or UO_1185 (O_1185,N_15160,N_17566);
xor UO_1186 (O_1186,N_18290,N_17885);
xor UO_1187 (O_1187,N_19645,N_17191);
nor UO_1188 (O_1188,N_16452,N_16159);
and UO_1189 (O_1189,N_19184,N_16343);
nand UO_1190 (O_1190,N_18053,N_16070);
nor UO_1191 (O_1191,N_16600,N_17874);
nor UO_1192 (O_1192,N_18968,N_19488);
nand UO_1193 (O_1193,N_17674,N_19906);
and UO_1194 (O_1194,N_17096,N_17085);
nor UO_1195 (O_1195,N_16469,N_15307);
nand UO_1196 (O_1196,N_19359,N_15953);
nand UO_1197 (O_1197,N_15403,N_18500);
nor UO_1198 (O_1198,N_17479,N_18466);
nor UO_1199 (O_1199,N_15584,N_16093);
nor UO_1200 (O_1200,N_18435,N_15114);
nor UO_1201 (O_1201,N_17904,N_17666);
or UO_1202 (O_1202,N_19528,N_19996);
or UO_1203 (O_1203,N_19437,N_18771);
xnor UO_1204 (O_1204,N_16945,N_15527);
xnor UO_1205 (O_1205,N_16428,N_18512);
nor UO_1206 (O_1206,N_18524,N_15003);
or UO_1207 (O_1207,N_19079,N_18516);
nand UO_1208 (O_1208,N_16821,N_18808);
or UO_1209 (O_1209,N_17575,N_16650);
and UO_1210 (O_1210,N_19594,N_17598);
nand UO_1211 (O_1211,N_16282,N_18837);
or UO_1212 (O_1212,N_19686,N_16340);
and UO_1213 (O_1213,N_15589,N_19325);
xnor UO_1214 (O_1214,N_18707,N_15947);
nor UO_1215 (O_1215,N_18698,N_16314);
and UO_1216 (O_1216,N_15609,N_15646);
nor UO_1217 (O_1217,N_15765,N_17471);
xnor UO_1218 (O_1218,N_17538,N_16611);
or UO_1219 (O_1219,N_18725,N_17670);
nand UO_1220 (O_1220,N_15926,N_18338);
nor UO_1221 (O_1221,N_16451,N_19572);
or UO_1222 (O_1222,N_15340,N_15694);
and UO_1223 (O_1223,N_16647,N_18085);
or UO_1224 (O_1224,N_16959,N_18818);
xor UO_1225 (O_1225,N_18187,N_18469);
xor UO_1226 (O_1226,N_15526,N_18003);
and UO_1227 (O_1227,N_16212,N_19424);
nand UO_1228 (O_1228,N_17228,N_17671);
or UO_1229 (O_1229,N_19998,N_18825);
nand UO_1230 (O_1230,N_15110,N_19193);
nor UO_1231 (O_1231,N_15795,N_18360);
nor UO_1232 (O_1232,N_16912,N_15597);
nand UO_1233 (O_1233,N_18985,N_15531);
xnor UO_1234 (O_1234,N_19307,N_17385);
xnor UO_1235 (O_1235,N_18560,N_15678);
nor UO_1236 (O_1236,N_17193,N_16997);
nand UO_1237 (O_1237,N_16503,N_19517);
and UO_1238 (O_1238,N_17225,N_17866);
and UO_1239 (O_1239,N_16525,N_18043);
nand UO_1240 (O_1240,N_15569,N_18390);
nand UO_1241 (O_1241,N_17700,N_16524);
nand UO_1242 (O_1242,N_18091,N_17997);
nand UO_1243 (O_1243,N_19890,N_18233);
and UO_1244 (O_1244,N_18021,N_18142);
nor UO_1245 (O_1245,N_18089,N_16021);
or UO_1246 (O_1246,N_19241,N_19128);
nand UO_1247 (O_1247,N_15041,N_16752);
and UO_1248 (O_1248,N_15311,N_18587);
nand UO_1249 (O_1249,N_19259,N_18077);
or UO_1250 (O_1250,N_15533,N_17451);
nor UO_1251 (O_1251,N_17449,N_19188);
xor UO_1252 (O_1252,N_18738,N_15875);
nand UO_1253 (O_1253,N_18665,N_19003);
xnor UO_1254 (O_1254,N_16105,N_18440);
xnor UO_1255 (O_1255,N_16505,N_15250);
xnor UO_1256 (O_1256,N_16564,N_16097);
and UO_1257 (O_1257,N_17715,N_15385);
and UO_1258 (O_1258,N_17292,N_18585);
xor UO_1259 (O_1259,N_19393,N_15714);
nor UO_1260 (O_1260,N_18572,N_15459);
nor UO_1261 (O_1261,N_16084,N_19238);
xor UO_1262 (O_1262,N_17683,N_16626);
nand UO_1263 (O_1263,N_19739,N_18885);
nor UO_1264 (O_1264,N_17724,N_19088);
and UO_1265 (O_1265,N_17921,N_19122);
nor UO_1266 (O_1266,N_17849,N_19202);
or UO_1267 (O_1267,N_16839,N_19397);
or UO_1268 (O_1268,N_18562,N_18227);
xnor UO_1269 (O_1269,N_17197,N_17240);
nand UO_1270 (O_1270,N_17952,N_16940);
nor UO_1271 (O_1271,N_15494,N_17992);
and UO_1272 (O_1272,N_16526,N_19341);
xnor UO_1273 (O_1273,N_18709,N_19763);
nor UO_1274 (O_1274,N_15560,N_17590);
xor UO_1275 (O_1275,N_18748,N_18329);
nand UO_1276 (O_1276,N_15419,N_16866);
or UO_1277 (O_1277,N_17630,N_17498);
nor UO_1278 (O_1278,N_19693,N_17084);
nor UO_1279 (O_1279,N_15772,N_18686);
nor UO_1280 (O_1280,N_19929,N_16252);
nor UO_1281 (O_1281,N_17210,N_18071);
nand UO_1282 (O_1282,N_19176,N_19685);
nor UO_1283 (O_1283,N_15858,N_16753);
nor UO_1284 (O_1284,N_17110,N_19254);
nor UO_1285 (O_1285,N_15481,N_19689);
xor UO_1286 (O_1286,N_17792,N_18325);
xor UO_1287 (O_1287,N_18787,N_19195);
and UO_1288 (O_1288,N_19484,N_17038);
xor UO_1289 (O_1289,N_19082,N_18209);
and UO_1290 (O_1290,N_15726,N_16560);
xnor UO_1291 (O_1291,N_19827,N_18775);
or UO_1292 (O_1292,N_19032,N_17067);
nand UO_1293 (O_1293,N_15954,N_16302);
nor UO_1294 (O_1294,N_16778,N_19971);
and UO_1295 (O_1295,N_18202,N_16651);
or UO_1296 (O_1296,N_15648,N_19351);
nor UO_1297 (O_1297,N_17884,N_18175);
and UO_1298 (O_1298,N_16655,N_18065);
xnor UO_1299 (O_1299,N_18413,N_15327);
nor UO_1300 (O_1300,N_19756,N_19166);
nor UO_1301 (O_1301,N_17798,N_16806);
nor UO_1302 (O_1302,N_19657,N_16124);
nor UO_1303 (O_1303,N_16004,N_16787);
and UO_1304 (O_1304,N_18541,N_16328);
xor UO_1305 (O_1305,N_18723,N_19950);
nand UO_1306 (O_1306,N_16243,N_19420);
and UO_1307 (O_1307,N_16062,N_19331);
xor UO_1308 (O_1308,N_16300,N_18673);
and UO_1309 (O_1309,N_19854,N_15478);
or UO_1310 (O_1310,N_19051,N_19124);
nor UO_1311 (O_1311,N_16222,N_18554);
or UO_1312 (O_1312,N_16540,N_16492);
xor UO_1313 (O_1313,N_16058,N_18300);
nand UO_1314 (O_1314,N_15098,N_19342);
or UO_1315 (O_1315,N_18464,N_19694);
xor UO_1316 (O_1316,N_16883,N_16135);
or UO_1317 (O_1317,N_16147,N_18113);
nor UO_1318 (O_1318,N_18791,N_15873);
and UO_1319 (O_1319,N_15836,N_17302);
nor UO_1320 (O_1320,N_15568,N_18913);
or UO_1321 (O_1321,N_17756,N_18302);
xnor UO_1322 (O_1322,N_15276,N_16648);
nor UO_1323 (O_1323,N_17699,N_15996);
or UO_1324 (O_1324,N_15661,N_19021);
xor UO_1325 (O_1325,N_17889,N_19095);
and UO_1326 (O_1326,N_16368,N_19913);
nor UO_1327 (O_1327,N_18172,N_18711);
nand UO_1328 (O_1328,N_18022,N_17280);
or UO_1329 (O_1329,N_18237,N_18892);
or UO_1330 (O_1330,N_17612,N_15574);
nor UO_1331 (O_1331,N_18228,N_16969);
xor UO_1332 (O_1332,N_18409,N_19716);
xnor UO_1333 (O_1333,N_15308,N_16336);
or UO_1334 (O_1334,N_19232,N_15708);
or UO_1335 (O_1335,N_15040,N_18730);
nor UO_1336 (O_1336,N_19764,N_15350);
and UO_1337 (O_1337,N_18309,N_19427);
xnor UO_1338 (O_1338,N_15183,N_19719);
nor UO_1339 (O_1339,N_18690,N_16213);
nand UO_1340 (O_1340,N_16875,N_17601);
and UO_1341 (O_1341,N_19717,N_18392);
nor UO_1342 (O_1342,N_16494,N_15344);
or UO_1343 (O_1343,N_17301,N_16507);
nand UO_1344 (O_1344,N_19704,N_17173);
or UO_1345 (O_1345,N_16693,N_15487);
nor UO_1346 (O_1346,N_17091,N_18157);
nor UO_1347 (O_1347,N_15044,N_15824);
or UO_1348 (O_1348,N_18479,N_17458);
or UO_1349 (O_1349,N_17627,N_15603);
xor UO_1350 (O_1350,N_18327,N_17606);
xor UO_1351 (O_1351,N_15684,N_18230);
nor UO_1352 (O_1352,N_17748,N_17669);
xor UO_1353 (O_1353,N_19078,N_17098);
nand UO_1354 (O_1354,N_19213,N_16705);
or UO_1355 (O_1355,N_16040,N_15538);
or UO_1356 (O_1356,N_17704,N_19239);
or UO_1357 (O_1357,N_15598,N_19831);
nor UO_1358 (O_1358,N_15513,N_16865);
nor UO_1359 (O_1359,N_15042,N_16356);
xnor UO_1360 (O_1360,N_16417,N_17105);
or UO_1361 (O_1361,N_17274,N_19647);
xnor UO_1362 (O_1362,N_15283,N_16422);
and UO_1363 (O_1363,N_17260,N_19581);
xnor UO_1364 (O_1364,N_17276,N_18002);
nand UO_1365 (O_1365,N_18364,N_18450);
or UO_1366 (O_1366,N_17338,N_18977);
or UO_1367 (O_1367,N_18379,N_15890);
and UO_1368 (O_1368,N_19151,N_18900);
xor UO_1369 (O_1369,N_15647,N_15136);
nor UO_1370 (O_1370,N_19328,N_18740);
nand UO_1371 (O_1371,N_16037,N_18693);
nand UO_1372 (O_1372,N_17526,N_19946);
or UO_1373 (O_1373,N_18970,N_17752);
xor UO_1374 (O_1374,N_17072,N_18785);
nand UO_1375 (O_1375,N_19956,N_17382);
xnor UO_1376 (O_1376,N_15192,N_18920);
xnor UO_1377 (O_1377,N_19018,N_16441);
nor UO_1378 (O_1378,N_16774,N_18484);
or UO_1379 (O_1379,N_19354,N_16270);
or UO_1380 (O_1380,N_15013,N_15173);
nor UO_1381 (O_1381,N_18497,N_19286);
nor UO_1382 (O_1382,N_15982,N_15095);
nor UO_1383 (O_1383,N_15430,N_15823);
nand UO_1384 (O_1384,N_18397,N_19654);
nor UO_1385 (O_1385,N_16397,N_15096);
xor UO_1386 (O_1386,N_15080,N_18431);
xor UO_1387 (O_1387,N_19030,N_19471);
or UO_1388 (O_1388,N_15265,N_17753);
or UO_1389 (O_1389,N_17597,N_15274);
xor UO_1390 (O_1390,N_16754,N_16313);
or UO_1391 (O_1391,N_15820,N_19038);
nor UO_1392 (O_1392,N_19641,N_16198);
xor UO_1393 (O_1393,N_17113,N_18447);
nor UO_1394 (O_1394,N_18382,N_17181);
xnor UO_1395 (O_1395,N_18801,N_17472);
and UO_1396 (O_1396,N_16499,N_18494);
and UO_1397 (O_1397,N_16468,N_15145);
nand UO_1398 (O_1398,N_18313,N_15490);
nor UO_1399 (O_1399,N_16459,N_19895);
nand UO_1400 (O_1400,N_16559,N_18797);
xnor UO_1401 (O_1401,N_16823,N_17021);
nand UO_1402 (O_1402,N_17230,N_15006);
nor UO_1403 (O_1403,N_19183,N_18687);
nor UO_1404 (O_1404,N_17019,N_17081);
xnor UO_1405 (O_1405,N_18529,N_18812);
or UO_1406 (O_1406,N_16402,N_15375);
nand UO_1407 (O_1407,N_17654,N_16544);
and UO_1408 (O_1408,N_19253,N_16635);
or UO_1409 (O_1409,N_15062,N_16904);
nand UO_1410 (O_1410,N_15366,N_17069);
nand UO_1411 (O_1411,N_15605,N_18070);
and UO_1412 (O_1412,N_16087,N_18720);
nor UO_1413 (O_1413,N_16168,N_18080);
and UO_1414 (O_1414,N_16308,N_16584);
and UO_1415 (O_1415,N_17757,N_17703);
and UO_1416 (O_1416,N_16739,N_16517);
nand UO_1417 (O_1417,N_16829,N_18054);
nor UO_1418 (O_1418,N_17881,N_15108);
or UO_1419 (O_1419,N_15613,N_15555);
xor UO_1420 (O_1420,N_19226,N_18274);
nor UO_1421 (O_1421,N_19441,N_18370);
and UO_1422 (O_1422,N_19567,N_18805);
and UO_1423 (O_1423,N_15851,N_18631);
xor UO_1424 (O_1424,N_18786,N_19885);
and UO_1425 (O_1425,N_18328,N_18753);
nand UO_1426 (O_1426,N_18127,N_17847);
or UO_1427 (O_1427,N_15614,N_19058);
or UO_1428 (O_1428,N_16545,N_18105);
and UO_1429 (O_1429,N_18326,N_18972);
xor UO_1430 (O_1430,N_16763,N_18557);
or UO_1431 (O_1431,N_19447,N_19735);
nor UO_1432 (O_1432,N_18362,N_18009);
nand UO_1433 (O_1433,N_19294,N_15876);
and UO_1434 (O_1434,N_16466,N_19882);
nand UO_1435 (O_1435,N_17578,N_15070);
or UO_1436 (O_1436,N_16409,N_19185);
and UO_1437 (O_1437,N_16729,N_19099);
nand UO_1438 (O_1438,N_19952,N_19457);
nor UO_1439 (O_1439,N_17865,N_18613);
xor UO_1440 (O_1440,N_18411,N_18821);
and UO_1441 (O_1441,N_15162,N_16327);
or UO_1442 (O_1442,N_18477,N_18965);
nand UO_1443 (O_1443,N_17233,N_17182);
or UO_1444 (O_1444,N_17241,N_18428);
and UO_1445 (O_1445,N_16148,N_19917);
nor UO_1446 (O_1446,N_16528,N_15057);
and UO_1447 (O_1447,N_16935,N_19211);
xor UO_1448 (O_1448,N_15444,N_17428);
xnor UO_1449 (O_1449,N_16432,N_19474);
or UO_1450 (O_1450,N_17963,N_15859);
nand UO_1451 (O_1451,N_18507,N_15339);
or UO_1452 (O_1452,N_19740,N_16950);
xor UO_1453 (O_1453,N_19390,N_17591);
nand UO_1454 (O_1454,N_19335,N_15724);
nor UO_1455 (O_1455,N_16977,N_18960);
or UO_1456 (O_1456,N_18220,N_17621);
or UO_1457 (O_1457,N_17721,N_17956);
or UO_1458 (O_1458,N_16922,N_17087);
and UO_1459 (O_1459,N_18263,N_17910);
nand UO_1460 (O_1460,N_18426,N_17039);
or UO_1461 (O_1461,N_17300,N_16244);
and UO_1462 (O_1462,N_19461,N_15693);
and UO_1463 (O_1463,N_15401,N_16500);
xnor UO_1464 (O_1464,N_15133,N_18420);
nand UO_1465 (O_1465,N_16011,N_19503);
or UO_1466 (O_1466,N_17324,N_15428);
nor UO_1467 (O_1467,N_15074,N_18863);
and UO_1468 (O_1468,N_19965,N_16798);
xnor UO_1469 (O_1469,N_19958,N_17031);
nand UO_1470 (O_1470,N_15960,N_18322);
nand UO_1471 (O_1471,N_19007,N_15154);
nor UO_1472 (O_1472,N_17312,N_16322);
xor UO_1473 (O_1473,N_15389,N_17340);
nor UO_1474 (O_1474,N_15161,N_16547);
and UO_1475 (O_1475,N_18445,N_17343);
nand UO_1476 (O_1476,N_17737,N_19107);
and UO_1477 (O_1477,N_19635,N_16678);
or UO_1478 (O_1478,N_16430,N_15871);
or UO_1479 (O_1479,N_15437,N_19809);
and UO_1480 (O_1480,N_18853,N_17396);
and UO_1481 (O_1481,N_16673,N_18721);
or UO_1482 (O_1482,N_15658,N_16388);
xor UO_1483 (O_1483,N_15545,N_18508);
and UO_1484 (O_1484,N_16048,N_19782);
nor UO_1485 (O_1485,N_17909,N_15262);
and UO_1486 (O_1486,N_19724,N_17059);
nand UO_1487 (O_1487,N_18218,N_15463);
and UO_1488 (O_1488,N_19006,N_19944);
or UO_1489 (O_1489,N_18485,N_15257);
and UO_1490 (O_1490,N_18656,N_17051);
or UO_1491 (O_1491,N_15827,N_19069);
or UO_1492 (O_1492,N_19989,N_19842);
and UO_1493 (O_1493,N_15588,N_17108);
and UO_1494 (O_1494,N_18847,N_15188);
or UO_1495 (O_1495,N_16578,N_18849);
xor UO_1496 (O_1496,N_15364,N_15566);
nand UO_1497 (O_1497,N_16911,N_15166);
nor UO_1498 (O_1498,N_16531,N_15732);
and UO_1499 (O_1499,N_17931,N_16065);
nor UO_1500 (O_1500,N_18214,N_17009);
or UO_1501 (O_1501,N_17727,N_18051);
nand UO_1502 (O_1502,N_18727,N_17388);
nand UO_1503 (O_1503,N_17148,N_19959);
and UO_1504 (O_1504,N_15222,N_19832);
xor UO_1505 (O_1505,N_18894,N_18739);
nand UO_1506 (O_1506,N_18666,N_15317);
nor UO_1507 (O_1507,N_19160,N_18758);
nand UO_1508 (O_1508,N_18180,N_15227);
xor UO_1509 (O_1509,N_15296,N_17559);
xor UO_1510 (O_1510,N_18017,N_17927);
nor UO_1511 (O_1511,N_19438,N_18594);
nor UO_1512 (O_1512,N_15523,N_15150);
xnor UO_1513 (O_1513,N_15155,N_16165);
xor UO_1514 (O_1514,N_16122,N_19000);
and UO_1515 (O_1515,N_19507,N_17172);
xnor UO_1516 (O_1516,N_18050,N_19261);
or UO_1517 (O_1517,N_15022,N_16855);
xnor UO_1518 (O_1518,N_19583,N_18764);
and UO_1519 (O_1519,N_15839,N_17686);
nand UO_1520 (O_1520,N_17076,N_15314);
nor UO_1521 (O_1521,N_19780,N_19316);
nand UO_1522 (O_1522,N_17433,N_16676);
xnor UO_1523 (O_1523,N_15220,N_15353);
nor UO_1524 (O_1524,N_19242,N_15979);
and UO_1525 (O_1525,N_17938,N_15636);
or UO_1526 (O_1526,N_18083,N_16970);
nand UO_1527 (O_1527,N_16566,N_19216);
nand UO_1528 (O_1528,N_18928,N_19186);
nand UO_1529 (O_1529,N_19834,N_18879);
nor UO_1530 (O_1530,N_16598,N_18436);
nor UO_1531 (O_1531,N_19343,N_15943);
xnor UO_1532 (O_1532,N_17510,N_17097);
or UO_1533 (O_1533,N_16361,N_19247);
xnor UO_1534 (O_1534,N_19045,N_17781);
or UO_1535 (O_1535,N_15920,N_16919);
xnor UO_1536 (O_1536,N_15367,N_18906);
or UO_1537 (O_1537,N_17561,N_17854);
xnor UO_1538 (O_1538,N_19869,N_19741);
or UO_1539 (O_1539,N_16465,N_15370);
xor UO_1540 (O_1540,N_19399,N_18603);
nand UO_1541 (O_1541,N_19668,N_18590);
nor UO_1542 (O_1542,N_17406,N_18553);
xor UO_1543 (O_1543,N_18728,N_19878);
or UO_1544 (O_1544,N_18817,N_19453);
nor UO_1545 (O_1545,N_16027,N_19223);
or UO_1546 (O_1546,N_17716,N_19680);
nor UO_1547 (O_1547,N_15281,N_17387);
and UO_1548 (O_1548,N_18645,N_17485);
nand UO_1549 (O_1549,N_15163,N_16605);
and UO_1550 (O_1550,N_17978,N_16567);
nand UO_1551 (O_1551,N_18638,N_16629);
or UO_1552 (O_1552,N_15190,N_18652);
nand UO_1553 (O_1553,N_16721,N_19149);
nor UO_1554 (O_1554,N_18657,N_15388);
nand UO_1555 (O_1555,N_17766,N_16991);
or UO_1556 (O_1556,N_18024,N_15576);
nand UO_1557 (O_1557,N_18946,N_16734);
and UO_1558 (O_1558,N_16680,N_15917);
or UO_1559 (O_1559,N_17196,N_17820);
xor UO_1560 (O_1560,N_19705,N_15035);
xnor UO_1561 (O_1561,N_16874,N_16179);
nor UO_1562 (O_1562,N_16142,N_16144);
nand UO_1563 (O_1563,N_17050,N_19042);
nor UO_1564 (O_1564,N_17586,N_19545);
nand UO_1565 (O_1565,N_18632,N_19930);
or UO_1566 (O_1566,N_16038,N_17114);
nor UO_1567 (O_1567,N_18352,N_17567);
and UO_1568 (O_1568,N_17819,N_15722);
and UO_1569 (O_1569,N_16303,N_17991);
nor UO_1570 (O_1570,N_18165,N_15995);
and UO_1571 (O_1571,N_16224,N_19891);
xor UO_1572 (O_1572,N_19851,N_19548);
or UO_1573 (O_1573,N_17275,N_19101);
nor UO_1574 (O_1574,N_15769,N_18517);
nand UO_1575 (O_1575,N_19634,N_16941);
or UO_1576 (O_1576,N_16171,N_15231);
xor UO_1577 (O_1577,N_15761,N_15758);
or UO_1578 (O_1578,N_19918,N_16879);
nor UO_1579 (O_1579,N_19490,N_15312);
nor UO_1580 (O_1580,N_17234,N_19662);
and UO_1581 (O_1581,N_18373,N_19207);
xor UO_1582 (O_1582,N_19411,N_19460);
nand UO_1583 (O_1583,N_16350,N_18470);
or UO_1584 (O_1584,N_15443,N_15686);
and UO_1585 (O_1585,N_19945,N_15084);
xnor UO_1586 (O_1586,N_16553,N_16177);
nor UO_1587 (O_1587,N_19117,N_17368);
and UO_1588 (O_1588,N_18251,N_19866);
or UO_1589 (O_1589,N_17318,N_19598);
xnor UO_1590 (O_1590,N_19818,N_15204);
nor UO_1591 (O_1591,N_16746,N_19660);
or UO_1592 (O_1592,N_19889,N_19310);
nor UO_1593 (O_1593,N_16041,N_19108);
xor UO_1594 (O_1594,N_19210,N_19498);
or UO_1595 (O_1595,N_19638,N_17570);
nand UO_1596 (O_1596,N_15791,N_15477);
or UO_1597 (O_1597,N_17557,N_16826);
nor UO_1598 (O_1598,N_17603,N_19691);
nand UO_1599 (O_1599,N_19385,N_19639);
nand UO_1600 (O_1600,N_15131,N_17763);
nor UO_1601 (O_1601,N_16585,N_15615);
or UO_1602 (O_1602,N_17943,N_19360);
or UO_1603 (O_1603,N_19672,N_19792);
nand UO_1604 (O_1604,N_19671,N_16910);
and UO_1605 (O_1605,N_16401,N_16044);
nand UO_1606 (O_1606,N_18483,N_17066);
nand UO_1607 (O_1607,N_18502,N_17285);
nand UO_1608 (O_1608,N_15313,N_19565);
and UO_1609 (O_1609,N_19173,N_15813);
xor UO_1610 (O_1610,N_17891,N_18417);
and UO_1611 (O_1611,N_16954,N_17265);
nand UO_1612 (O_1612,N_16812,N_16917);
or UO_1613 (O_1613,N_15412,N_17248);
nand UO_1614 (O_1614,N_19442,N_19161);
nor UO_1615 (O_1615,N_15267,N_17624);
or UO_1616 (O_1616,N_16899,N_15515);
nand UO_1617 (O_1617,N_17587,N_17767);
xor UO_1618 (O_1618,N_17574,N_17466);
nor UO_1619 (O_1619,N_15897,N_19435);
and UO_1620 (O_1620,N_17768,N_17657);
or UO_1621 (O_1621,N_15924,N_18776);
or UO_1622 (O_1622,N_17697,N_17329);
nor UO_1623 (O_1623,N_18330,N_18792);
nor UO_1624 (O_1624,N_19861,N_16054);
nor UO_1625 (O_1625,N_16583,N_17134);
or UO_1626 (O_1626,N_19628,N_16827);
nand UO_1627 (O_1627,N_18745,N_16716);
nand UO_1628 (O_1628,N_15097,N_19947);
or UO_1629 (O_1629,N_16641,N_18465);
or UO_1630 (O_1630,N_18015,N_16989);
nor UO_1631 (O_1631,N_15811,N_18407);
xnor UO_1632 (O_1632,N_18978,N_15815);
nor UO_1633 (O_1633,N_18949,N_18883);
nor UO_1634 (O_1634,N_17899,N_17252);
and UO_1635 (O_1635,N_18179,N_17361);
xnor UO_1636 (O_1636,N_18633,N_16009);
or UO_1637 (O_1637,N_16699,N_15452);
nand UO_1638 (O_1638,N_15781,N_17045);
xnor UO_1639 (O_1639,N_19603,N_15195);
or UO_1640 (O_1640,N_15773,N_17518);
xor UO_1641 (O_1641,N_16708,N_19541);
and UO_1642 (O_1642,N_17171,N_15771);
or UO_1643 (O_1643,N_15337,N_19287);
xor UO_1644 (O_1644,N_16116,N_15742);
and UO_1645 (O_1645,N_17585,N_17284);
and UO_1646 (O_1646,N_18592,N_18372);
nand UO_1647 (O_1647,N_17625,N_16026);
or UO_1648 (O_1648,N_16653,N_15346);
nor UO_1649 (O_1649,N_19406,N_16995);
and UO_1650 (O_1650,N_17786,N_18163);
xor UO_1651 (O_1651,N_19388,N_17718);
nand UO_1652 (O_1652,N_17095,N_15082);
nand UO_1653 (O_1653,N_15076,N_19623);
and UO_1654 (O_1654,N_19730,N_18047);
or UO_1655 (O_1655,N_17925,N_15886);
nand UO_1656 (O_1656,N_15721,N_19156);
nor UO_1657 (O_1657,N_16965,N_18705);
nand UO_1658 (O_1658,N_16205,N_17023);
and UO_1659 (O_1659,N_17837,N_17070);
and UO_1660 (O_1660,N_19852,N_15031);
xor UO_1661 (O_1661,N_16636,N_17482);
xnor UO_1662 (O_1662,N_19220,N_19104);
and UO_1663 (O_1663,N_15225,N_15189);
nor UO_1664 (O_1664,N_15747,N_17437);
and UO_1665 (O_1665,N_15284,N_16339);
nand UO_1666 (O_1666,N_17582,N_17812);
and UO_1667 (O_1667,N_16391,N_16496);
or UO_1668 (O_1668,N_18462,N_16052);
nor UO_1669 (O_1669,N_19448,N_19070);
nand UO_1670 (O_1670,N_19713,N_15857);
nor UO_1671 (O_1671,N_18048,N_15064);
nand UO_1672 (O_1672,N_16207,N_15899);
or UO_1673 (O_1673,N_15981,N_18896);
or UO_1674 (O_1674,N_17863,N_18647);
and UO_1675 (O_1675,N_15194,N_15186);
xor UO_1676 (O_1676,N_19389,N_15951);
nor UO_1677 (O_1677,N_16860,N_19555);
xnor UO_1678 (O_1678,N_17839,N_16088);
nor UO_1679 (O_1679,N_17107,N_17454);
and UO_1680 (O_1680,N_15051,N_18285);
xor UO_1681 (O_1681,N_15435,N_15010);
xnor UO_1682 (O_1682,N_16332,N_15921);
nor UO_1683 (O_1683,N_15809,N_17287);
nor UO_1684 (O_1684,N_18168,N_17651);
nor UO_1685 (O_1685,N_16630,N_17497);
and UO_1686 (O_1686,N_19419,N_19012);
nand UO_1687 (O_1687,N_18289,N_15351);
or UO_1688 (O_1688,N_18356,N_16645);
or UO_1689 (O_1689,N_18389,N_19772);
nand UO_1690 (O_1690,N_17013,N_17103);
and UO_1691 (O_1691,N_15361,N_15530);
and UO_1692 (O_1692,N_19391,N_18155);
or UO_1693 (O_1693,N_16672,N_19491);
or UO_1694 (O_1694,N_15594,N_15230);
xor UO_1695 (O_1695,N_17576,N_18493);
and UO_1696 (O_1696,N_16644,N_16682);
xnor UO_1697 (O_1697,N_18899,N_15273);
nand UO_1698 (O_1698,N_16109,N_19052);
nor UO_1699 (O_1699,N_19081,N_15030);
nor UO_1700 (O_1700,N_19825,N_18924);
and UO_1701 (O_1701,N_19440,N_18419);
nand UO_1702 (O_1702,N_19663,N_19381);
nor UO_1703 (O_1703,N_17080,N_15590);
and UO_1704 (O_1704,N_18933,N_15263);
and UO_1705 (O_1705,N_18583,N_15939);
and UO_1706 (O_1706,N_19807,N_16666);
xor UO_1707 (O_1707,N_16833,N_17778);
nand UO_1708 (O_1708,N_19102,N_16958);
and UO_1709 (O_1709,N_15498,N_17267);
nor UO_1710 (O_1710,N_17516,N_17877);
nor UO_1711 (O_1711,N_15246,N_18939);
and UO_1712 (O_1712,N_15060,N_15497);
nor UO_1713 (O_1713,N_15360,N_15879);
xnor UO_1714 (O_1714,N_19862,N_19074);
xor UO_1715 (O_1715,N_17709,N_16013);
xnor UO_1716 (O_1716,N_17376,N_15315);
xor UO_1717 (O_1717,N_16596,N_18359);
or UO_1718 (O_1718,N_17434,N_17641);
and UO_1719 (O_1719,N_18692,N_16025);
and UO_1720 (O_1720,N_17237,N_19277);
nor UO_1721 (O_1721,N_17355,N_16478);
xor UO_1722 (O_1722,N_17916,N_16415);
nand UO_1723 (O_1723,N_16764,N_15223);
or UO_1724 (O_1724,N_18746,N_15983);
and UO_1725 (O_1725,N_19823,N_16723);
or UO_1726 (O_1726,N_18622,N_16420);
and UO_1727 (O_1727,N_16260,N_15998);
or UO_1728 (O_1728,N_19708,N_15938);
xor UO_1729 (O_1729,N_18387,N_19218);
and UO_1730 (O_1730,N_19125,N_17832);
and UO_1731 (O_1731,N_16342,N_16225);
and UO_1732 (O_1732,N_18103,N_15635);
and UO_1733 (O_1733,N_18402,N_15248);
xnor UO_1734 (O_1734,N_18474,N_19669);
xnor UO_1735 (O_1735,N_19841,N_19304);
nor UO_1736 (O_1736,N_15479,N_18544);
nor UO_1737 (O_1737,N_16745,N_17400);
xor UO_1738 (O_1738,N_17954,N_18336);
nand UO_1739 (O_1739,N_15931,N_18752);
nor UO_1740 (O_1740,N_15301,N_19019);
nand UO_1741 (O_1741,N_17037,N_19472);
nand UO_1742 (O_1742,N_17128,N_17083);
or UO_1743 (O_1743,N_15407,N_16933);
nor UO_1744 (O_1744,N_19991,N_18284);
nor UO_1745 (O_1745,N_18700,N_16298);
nor UO_1746 (O_1746,N_19064,N_17692);
and UO_1747 (O_1747,N_15727,N_18851);
xor UO_1748 (O_1748,N_17908,N_19230);
and UO_1749 (O_1749,N_19938,N_18580);
nor UO_1750 (O_1750,N_15653,N_18213);
xnor UO_1751 (O_1751,N_15792,N_18236);
xor UO_1752 (O_1752,N_15563,N_17394);
and UO_1753 (O_1753,N_16845,N_18644);
nor UO_1754 (O_1754,N_16588,N_19350);
nand UO_1755 (O_1755,N_17618,N_18480);
and UO_1756 (O_1756,N_19141,N_17855);
nor UO_1757 (O_1757,N_16299,N_18159);
or UO_1758 (O_1758,N_19071,N_19252);
xnor UO_1759 (O_1759,N_18499,N_19127);
xor UO_1760 (O_1760,N_18122,N_16473);
or UO_1761 (O_1761,N_19667,N_18609);
or UO_1762 (O_1762,N_15000,N_16916);
or UO_1763 (O_1763,N_18299,N_16008);
xnor UO_1764 (O_1764,N_18297,N_16575);
xor UO_1765 (O_1765,N_17742,N_16146);
nand UO_1766 (O_1766,N_19801,N_19863);
nor UO_1767 (O_1767,N_17560,N_17677);
nand UO_1768 (O_1768,N_18967,N_15787);
nand UO_1769 (O_1769,N_15768,N_17923);
or UO_1770 (O_1770,N_19547,N_19324);
nor UO_1771 (O_1771,N_16913,N_15390);
nand UO_1772 (O_1772,N_18672,N_16737);
and UO_1773 (O_1773,N_15868,N_16354);
xor UO_1774 (O_1774,N_15019,N_17403);
and UO_1775 (O_1775,N_16864,N_16634);
xor UO_1776 (O_1776,N_19295,N_18521);
or UO_1777 (O_1777,N_15149,N_19473);
or UO_1778 (O_1778,N_17056,N_19995);
nor UO_1779 (O_1779,N_15501,N_16835);
nand UO_1780 (O_1780,N_17758,N_19289);
nand UO_1781 (O_1781,N_19229,N_18627);
nand UO_1782 (O_1782,N_17957,N_17232);
and UO_1783 (O_1783,N_17887,N_17730);
nand UO_1784 (O_1784,N_19339,N_19463);
nor UO_1785 (O_1785,N_16661,N_18174);
and UO_1786 (O_1786,N_19911,N_19910);
and UO_1787 (O_1787,N_15690,N_15808);
and UO_1788 (O_1788,N_19198,N_16273);
nand UO_1789 (O_1789,N_17794,N_18239);
and UO_1790 (O_1790,N_16915,N_15657);
and UO_1791 (O_1791,N_19313,N_18371);
or UO_1792 (O_1792,N_16595,N_18211);
xor UO_1793 (O_1793,N_18737,N_15902);
nand UO_1794 (O_1794,N_16838,N_19915);
and UO_1795 (O_1795,N_17239,N_19656);
nand UO_1796 (O_1796,N_18717,N_17143);
nand UO_1797 (O_1797,N_16522,N_16012);
nand UO_1798 (O_1798,N_16352,N_17006);
nand UO_1799 (O_1799,N_17202,N_18271);
nor UO_1800 (O_1800,N_15541,N_16126);
or UO_1801 (O_1801,N_18421,N_17488);
nor UO_1802 (O_1802,N_17858,N_15738);
nand UO_1803 (O_1803,N_15994,N_15739);
xor UO_1804 (O_1804,N_18386,N_15506);
or UO_1805 (O_1805,N_18511,N_18975);
and UO_1806 (O_1806,N_16822,N_19967);
nor UO_1807 (O_1807,N_16380,N_18461);
or UO_1808 (O_1808,N_16521,N_18434);
and UO_1809 (O_1809,N_18823,N_18321);
xnor UO_1810 (O_1810,N_19584,N_19751);
nand UO_1811 (O_1811,N_18111,N_15626);
xnor UO_1812 (O_1812,N_16285,N_15844);
or UO_1813 (O_1813,N_17335,N_16974);
nor UO_1814 (O_1814,N_16192,N_19060);
xnor UO_1815 (O_1815,N_18962,N_15429);
nor UO_1816 (O_1816,N_17356,N_17907);
nand UO_1817 (O_1817,N_18577,N_17313);
nor UO_1818 (O_1818,N_16527,N_19712);
and UO_1819 (O_1819,N_19482,N_16472);
xnor UO_1820 (O_1820,N_15259,N_17644);
or UO_1821 (O_1821,N_18205,N_17262);
and UO_1822 (O_1822,N_17279,N_19619);
or UO_1823 (O_1823,N_19839,N_19980);
nor UO_1824 (O_1824,N_17529,N_16197);
and UO_1825 (O_1825,N_18243,N_19673);
nor UO_1826 (O_1826,N_16856,N_19847);
and UO_1827 (O_1827,N_19092,N_16407);
and UO_1828 (O_1828,N_18961,N_15472);
xor UO_1829 (O_1829,N_17440,N_17184);
and UO_1830 (O_1830,N_17729,N_18191);
nand UO_1831 (O_1831,N_19065,N_17607);
and UO_1832 (O_1832,N_17841,N_17246);
xor UO_1833 (O_1833,N_17643,N_18124);
and UO_1834 (O_1834,N_19848,N_19087);
and UO_1835 (O_1835,N_17475,N_18346);
xor UO_1836 (O_1836,N_15903,N_19784);
nor UO_1837 (O_1837,N_16035,N_19372);
and UO_1838 (O_1838,N_15423,N_15476);
nand UO_1839 (O_1839,N_17012,N_15777);
xor UO_1840 (O_1840,N_17984,N_17733);
and UO_1841 (O_1841,N_16957,N_16255);
xor UO_1842 (O_1842,N_16543,N_17017);
or UO_1843 (O_1843,N_19048,N_16987);
xor UO_1844 (O_1844,N_17568,N_18861);
nor UO_1845 (O_1845,N_18806,N_16923);
xor UO_1846 (O_1846,N_19813,N_17571);
nor UO_1847 (O_1847,N_16967,N_19990);
nor UO_1848 (O_1848,N_19167,N_15798);
nand UO_1849 (O_1849,N_17177,N_17109);
or UO_1850 (O_1850,N_15359,N_19348);
xor UO_1851 (O_1851,N_17055,N_19364);
and UO_1852 (O_1852,N_17244,N_15338);
nor UO_1853 (O_1853,N_15334,N_17830);
nand UO_1854 (O_1854,N_15944,N_17354);
or UO_1855 (O_1855,N_18567,N_16570);
or UO_1856 (O_1856,N_17661,N_17033);
and UO_1857 (O_1857,N_17132,N_17178);
nand UO_1858 (O_1858,N_16805,N_16658);
or UO_1859 (O_1859,N_16937,N_16250);
xor UO_1860 (O_1860,N_18629,N_16190);
nor UO_1861 (O_1861,N_17545,N_17774);
nand UO_1862 (O_1862,N_17201,N_15422);
or UO_1863 (O_1863,N_18034,N_19421);
nand UO_1864 (O_1864,N_17157,N_19571);
nand UO_1865 (O_1865,N_17259,N_16656);
or UO_1866 (O_1866,N_16511,N_16139);
nor UO_1867 (O_1867,N_15409,N_19787);
xor UO_1868 (O_1868,N_17896,N_19371);
nand UO_1869 (O_1869,N_19309,N_16932);
xnor UO_1870 (O_1870,N_16117,N_19726);
xnor UO_1871 (O_1871,N_18246,N_18716);
nand UO_1872 (O_1872,N_17542,N_17199);
xnor UO_1873 (O_1873,N_19549,N_17784);
nor UO_1874 (O_1874,N_18800,N_15755);
and UO_1875 (O_1875,N_18219,N_17188);
and UO_1876 (O_1876,N_18616,N_16777);
nor UO_1877 (O_1877,N_19245,N_17223);
and UO_1878 (O_1878,N_16861,N_17919);
and UO_1879 (O_1879,N_17556,N_17769);
and UO_1880 (O_1880,N_19479,N_16263);
xor UO_1881 (O_1881,N_17002,N_17633);
nor UO_1882 (O_1882,N_19982,N_19062);
or UO_1883 (O_1883,N_16057,N_17665);
xor UO_1884 (O_1884,N_15654,N_17450);
nand UO_1885 (O_1885,N_15720,N_19139);
and UO_1886 (O_1886,N_18799,N_16768);
xor UO_1887 (O_1887,N_18542,N_19943);
xor UO_1888 (O_1888,N_16344,N_18416);
or UO_1889 (O_1889,N_16485,N_15585);
nand UO_1890 (O_1890,N_15891,N_19983);
nor UO_1891 (O_1891,N_16893,N_15208);
nand UO_1892 (O_1892,N_16438,N_15596);
xnor UO_1893 (O_1893,N_17212,N_19115);
nor UO_1894 (O_1894,N_15625,N_18807);
nor UO_1895 (O_1895,N_15893,N_15593);
nor UO_1896 (O_1896,N_15300,N_19483);
or UO_1897 (O_1897,N_17353,N_18475);
and UO_1898 (O_1898,N_18715,N_16247);
nand UO_1899 (O_1899,N_15869,N_15834);
and UO_1900 (O_1900,N_15254,N_18331);
nor UO_1901 (O_1901,N_19428,N_19939);
nand UO_1902 (O_1902,N_16077,N_15841);
xor UO_1903 (O_1903,N_15185,N_15357);
nor UO_1904 (O_1904,N_16476,N_17339);
nand UO_1905 (O_1905,N_16949,N_15007);
or UO_1906 (O_1906,N_15988,N_18455);
nor UO_1907 (O_1907,N_16188,N_17317);
and UO_1908 (O_1908,N_19516,N_19363);
and UO_1909 (O_1909,N_16063,N_18809);
nor UO_1910 (O_1910,N_16843,N_17540);
nor UO_1911 (O_1911,N_16549,N_17879);
nand UO_1912 (O_1912,N_19845,N_15985);
and UO_1913 (O_1913,N_19086,N_17664);
and UO_1914 (O_1914,N_16810,N_18935);
nand UO_1915 (O_1915,N_19659,N_18671);
xnor UO_1916 (O_1916,N_17850,N_17834);
or UO_1917 (O_1917,N_16371,N_19269);
xnor UO_1918 (O_1918,N_17906,N_16532);
or UO_1919 (O_1919,N_17917,N_18604);
xor UO_1920 (O_1920,N_15914,N_19790);
and UO_1921 (O_1921,N_16291,N_19553);
nand UO_1922 (O_1922,N_15786,N_16019);
xnor UO_1923 (O_1923,N_19905,N_17421);
nand UO_1924 (O_1924,N_17900,N_16467);
xnor UO_1925 (O_1925,N_18415,N_16434);
and UO_1926 (O_1926,N_18097,N_18248);
or UO_1927 (O_1927,N_16999,N_19661);
and UO_1928 (O_1928,N_15760,N_18349);
and UO_1929 (O_1929,N_17707,N_16101);
nor UO_1930 (O_1930,N_17762,N_16321);
or UO_1931 (O_1931,N_18925,N_18589);
nand UO_1932 (O_1932,N_16942,N_15540);
xnor UO_1933 (O_1933,N_15176,N_16081);
nand UO_1934 (O_1934,N_17236,N_17580);
xor UO_1935 (O_1935,N_17605,N_16045);
and UO_1936 (O_1936,N_19984,N_15837);
xor UO_1937 (O_1937,N_17423,N_18270);
nand UO_1938 (O_1938,N_17554,N_19962);
or UO_1939 (O_1939,N_18076,N_18146);
or UO_1940 (O_1940,N_17502,N_15181);
nor UO_1941 (O_1941,N_17523,N_19352);
nor UO_1942 (O_1942,N_15565,N_17214);
nand UO_1943 (O_1943,N_15129,N_16706);
xnor UO_1944 (O_1944,N_16358,N_16643);
nor UO_1945 (O_1945,N_17029,N_17932);
xor UO_1946 (O_1946,N_19644,N_16076);
and UO_1947 (O_1947,N_18607,N_15582);
xor UO_1948 (O_1948,N_19329,N_17543);
and UO_1949 (O_1949,N_18262,N_17291);
or UO_1950 (O_1950,N_15146,N_19957);
nor UO_1951 (O_1951,N_16061,N_16895);
and UO_1952 (O_1952,N_18950,N_15271);
or UO_1953 (O_1953,N_18193,N_16720);
xnor UO_1954 (O_1954,N_15286,N_18757);
or UO_1955 (O_1955,N_16447,N_19690);
xor UO_1956 (O_1956,N_19443,N_16010);
xor UO_1957 (O_1957,N_17950,N_15187);
nor UO_1958 (O_1958,N_17205,N_19928);
xor UO_1959 (O_1959,N_16381,N_18598);
xnor UO_1960 (O_1960,N_15294,N_16049);
and UO_1961 (O_1961,N_16731,N_15354);
nand UO_1962 (O_1962,N_15171,N_17948);
or UO_1963 (O_1963,N_18989,N_19093);
nor UO_1964 (O_1964,N_18742,N_18042);
nand UO_1965 (O_1965,N_18223,N_17391);
or UO_1966 (O_1966,N_18834,N_16174);
xnor UO_1967 (O_1967,N_19979,N_19355);
nand UO_1968 (O_1968,N_17293,N_15799);
xnor UO_1969 (O_1969,N_17869,N_18782);
and UO_1970 (O_1970,N_17822,N_17249);
nor UO_1971 (O_1971,N_15753,N_18150);
and UO_1972 (O_1972,N_18240,N_16337);
or UO_1973 (O_1973,N_15504,N_18197);
nor UO_1974 (O_1974,N_15586,N_16552);
and UO_1975 (O_1975,N_19055,N_17933);
xor UO_1976 (O_1976,N_18121,N_16137);
xnor UO_1977 (O_1977,N_17166,N_16138);
xor UO_1978 (O_1978,N_19522,N_17014);
xor UO_1979 (O_1979,N_15164,N_15731);
nor UO_1980 (O_1980,N_17731,N_19940);
xor UO_1981 (O_1981,N_19377,N_15669);
or UO_1982 (O_1982,N_18889,N_18573);
nand UO_1983 (O_1983,N_19779,N_19416);
or UO_1984 (O_1984,N_18614,N_18481);
xnor UO_1985 (O_1985,N_15829,N_17844);
nand UO_1986 (O_1986,N_19376,N_16443);
or UO_1987 (O_1987,N_16108,N_19715);
nor UO_1988 (O_1988,N_16766,N_15645);
nor UO_1989 (O_1989,N_15001,N_15448);
nor UO_1990 (O_1990,N_18164,N_19518);
and UO_1991 (O_1991,N_19024,N_17075);
nand UO_1992 (O_1992,N_15867,N_15916);
nor UO_1993 (O_1993,N_15923,N_18254);
nand UO_1994 (O_1994,N_16490,N_16283);
xor UO_1995 (O_1995,N_15123,N_15940);
or UO_1996 (O_1996,N_16018,N_19927);
and UO_1997 (O_1997,N_17604,N_18078);
and UO_1998 (O_1998,N_15529,N_16926);
and UO_1999 (O_1999,N_17852,N_15842);
nand UO_2000 (O_2000,N_16016,N_18063);
and UO_2001 (O_2001,N_15822,N_15304);
and UO_2002 (O_2002,N_19857,N_17829);
or UO_2003 (O_2003,N_19255,N_16280);
nand UO_2004 (O_2004,N_17743,N_16185);
xnor UO_2005 (O_2005,N_16194,N_17880);
nand UO_2006 (O_2006,N_19361,N_18829);
or UO_2007 (O_2007,N_19022,N_18250);
nand UO_2008 (O_2008,N_15134,N_15607);
or UO_2009 (O_2009,N_19201,N_19105);
xnor UO_2010 (O_2010,N_18534,N_16623);
nand UO_2011 (O_2011,N_19769,N_17307);
xnor UO_2012 (O_2012,N_16692,N_17801);
xnor UO_2013 (O_2013,N_16098,N_18221);
xnor UO_2014 (O_2014,N_15745,N_15821);
nand UO_2015 (O_2015,N_18365,N_17944);
or UO_2016 (O_2016,N_17444,N_19711);
nor UO_2017 (O_2017,N_19109,N_16820);
xor UO_2018 (O_2018,N_18699,N_17678);
or UO_2019 (O_2019,N_19029,N_15002);
and UO_2020 (O_2020,N_16433,N_17947);
or UO_2021 (O_2021,N_16852,N_16293);
nand UO_2022 (O_2022,N_19651,N_17772);
nor UO_2023 (O_2023,N_18836,N_18922);
or UO_2024 (O_2024,N_18954,N_18181);
xnor UO_2025 (O_2025,N_19802,N_19935);
or UO_2026 (O_2026,N_16296,N_15503);
nor UO_2027 (O_2027,N_16157,N_19675);
nor UO_2028 (O_2028,N_17631,N_17913);
and UO_2029 (O_2029,N_15063,N_19894);
or UO_2030 (O_2030,N_17817,N_16237);
or UO_2031 (O_2031,N_17398,N_18653);
xor UO_2032 (O_2032,N_16186,N_18915);
xnor UO_2033 (O_2033,N_17993,N_15826);
xor UO_2034 (O_2034,N_16324,N_16006);
nor UO_2035 (O_2035,N_19899,N_18045);
nor UO_2036 (O_2036,N_16930,N_18749);
nor UO_2037 (O_2037,N_15508,N_18282);
xor UO_2038 (O_2038,N_15580,N_17147);
and UO_2039 (O_2039,N_16457,N_16015);
nand UO_2040 (O_2040,N_18057,N_15029);
or UO_2041 (O_2041,N_15730,N_18741);
nor UO_2042 (O_2042,N_15465,N_16281);
nand UO_2043 (O_2043,N_18964,N_19901);
nor UO_2044 (O_2044,N_19805,N_18139);
xnor UO_2045 (O_2045,N_18098,N_16274);
xnor UO_2046 (O_2046,N_16537,N_15417);
nor UO_2047 (O_2047,N_15965,N_19132);
nand UO_2048 (O_2048,N_16355,N_17478);
or UO_2049 (O_2049,N_18948,N_18980);
nand UO_2050 (O_2050,N_19727,N_19589);
nand UO_2051 (O_2051,N_16277,N_18865);
nand UO_2052 (O_2052,N_16724,N_19446);
or UO_2053 (O_2053,N_15668,N_18167);
and UO_2054 (O_2054,N_16033,N_18173);
or UO_2055 (O_2055,N_18400,N_17412);
nor UO_2056 (O_2056,N_15440,N_18361);
nand UO_2057 (O_2057,N_17725,N_19423);
nor UO_2058 (O_2058,N_17551,N_15630);
or UO_2059 (O_2059,N_15073,N_19067);
nor UO_2060 (O_2060,N_17320,N_16976);
nor UO_2061 (O_2061,N_16887,N_17165);
nand UO_2062 (O_2062,N_19251,N_15521);
nor UO_2063 (O_2063,N_16257,N_18655);
nor UO_2064 (O_2064,N_17949,N_19791);
or UO_2065 (O_2065,N_15122,N_15118);
nand UO_2066 (O_2066,N_18999,N_15915);
nand UO_2067 (O_2067,N_17117,N_15807);
xnor UO_2068 (O_2068,N_17939,N_19936);
or UO_2069 (O_2069,N_17562,N_16885);
nor UO_2070 (O_2070,N_15557,N_19879);
xor UO_2071 (O_2071,N_19920,N_16613);
and UO_2072 (O_2072,N_16031,N_18145);
or UO_2073 (O_2073,N_15784,N_19225);
and UO_2074 (O_2074,N_18040,N_17548);
nor UO_2075 (O_2075,N_15004,N_18872);
or UO_2076 (O_2076,N_17011,N_18875);
and UO_2077 (O_2077,N_16379,N_18144);
nand UO_2078 (O_2078,N_17826,N_18952);
or UO_2079 (O_2079,N_16047,N_15043);
nand UO_2080 (O_2080,N_17857,N_16279);
or UO_2081 (O_2081,N_19625,N_19285);
or UO_2082 (O_2082,N_16928,N_15277);
xor UO_2083 (O_2083,N_18317,N_18982);
and UO_2084 (O_2084,N_15399,N_18586);
nor UO_2085 (O_2085,N_15680,N_15475);
nor UO_2086 (O_2086,N_15802,N_16986);
and UO_2087 (O_2087,N_19326,N_15748);
or UO_2088 (O_2088,N_19615,N_19688);
and UO_2089 (O_2089,N_18429,N_17512);
nand UO_2090 (O_2090,N_16229,N_15507);
nand UO_2091 (O_2091,N_15495,N_15520);
or UO_2092 (O_2092,N_18867,N_19013);
xnor UO_2093 (O_2093,N_16184,N_15956);
nor UO_2094 (O_2094,N_16265,N_16236);
nand UO_2095 (O_2095,N_19843,N_16683);
nor UO_2096 (O_2096,N_19954,N_18148);
xor UO_2097 (O_2097,N_18247,N_16007);
nor UO_2098 (O_2098,N_16896,N_19830);
or UO_2099 (O_2099,N_15216,N_15642);
or UO_2100 (O_2100,N_16214,N_19808);
nor UO_2101 (O_2101,N_19591,N_19768);
and UO_2102 (O_2102,N_15398,N_19197);
and UO_2103 (O_2103,N_17094,N_18295);
or UO_2104 (O_2104,N_19985,N_17026);
xor UO_2105 (O_2105,N_19096,N_15725);
nand UO_2106 (O_2106,N_15330,N_19836);
nand UO_2107 (O_2107,N_18454,N_16551);
and UO_2108 (O_2108,N_18708,N_17422);
xnor UO_2109 (O_2109,N_17647,N_18467);
nor UO_2110 (O_2110,N_17336,N_18199);
nand UO_2111 (O_2111,N_16562,N_17141);
and UO_2112 (O_2112,N_18064,N_18207);
nand UO_2113 (O_2113,N_16258,N_16853);
xor UO_2114 (O_2114,N_18276,N_17593);
xnor UO_2115 (O_2115,N_18055,N_16254);
or UO_2116 (O_2116,N_19334,N_16790);
xor UO_2117 (O_2117,N_16751,N_17595);
xnor UO_2118 (O_2118,N_19336,N_17243);
or UO_2119 (O_2119,N_16881,N_19169);
xor UO_2120 (O_2120,N_18724,N_17460);
or UO_2121 (O_2121,N_16068,N_19262);
nor UO_2122 (O_2122,N_17183,N_18770);
nor UO_2123 (O_2123,N_16530,N_19073);
or UO_2124 (O_2124,N_15453,N_18795);
and UO_2125 (O_2125,N_16436,N_18038);
xnor UO_2126 (O_2126,N_19551,N_16480);
nor UO_2127 (O_2127,N_17824,N_15913);
xnor UO_2128 (O_2128,N_15395,N_16854);
or UO_2129 (O_2129,N_16235,N_19942);
xnor UO_2130 (O_2130,N_16083,N_15804);
and UO_2131 (O_2131,N_16176,N_17969);
and UO_2132 (O_2132,N_15305,N_18350);
nand UO_2133 (O_2133,N_19902,N_19643);
or UO_2134 (O_2134,N_18058,N_17581);
and UO_2135 (O_2135,N_18576,N_19893);
or UO_2136 (O_2136,N_18605,N_15109);
nor UO_2137 (O_2137,N_17788,N_18565);
or UO_2138 (O_2138,N_18974,N_18151);
and UO_2139 (O_2139,N_15770,N_16968);
nor UO_2140 (O_2140,N_18087,N_16425);
or UO_2141 (O_2141,N_16153,N_19607);
nand UO_2142 (O_2142,N_15182,N_19224);
and UO_2143 (O_2143,N_19650,N_18092);
or UO_2144 (O_2144,N_19587,N_16487);
and UO_2145 (O_2145,N_17168,N_18520);
xor UO_2146 (O_2146,N_18856,N_15919);
or UO_2147 (O_2147,N_17118,N_15348);
or UO_2148 (O_2148,N_15391,N_15866);
and UO_2149 (O_2149,N_15922,N_18983);
and UO_2150 (O_2150,N_18636,N_18966);
nor UO_2151 (O_2151,N_19874,N_15604);
nand UO_2152 (O_2152,N_15439,N_15120);
nor UO_2153 (O_2153,N_19317,N_19451);
nor UO_2154 (O_2154,N_16892,N_18793);
and UO_2155 (O_2155,N_19914,N_15242);
and UO_2156 (O_2156,N_15848,N_19822);
nor UO_2157 (O_2157,N_15632,N_17027);
and UO_2158 (O_2158,N_16590,N_17446);
nor UO_2159 (O_2159,N_16631,N_17790);
nor UO_2160 (O_2160,N_17359,N_17179);
xnor UO_2161 (O_2161,N_15874,N_19215);
nand UO_2162 (O_2162,N_16632,N_15210);
and UO_2163 (O_2163,N_15282,N_19493);
and UO_2164 (O_2164,N_15534,N_16717);
or UO_2165 (O_2165,N_18628,N_18013);
nand UO_2166 (O_2166,N_19409,N_19542);
or UO_2167 (O_2167,N_16175,N_15255);
or UO_2168 (O_2168,N_16981,N_18601);
xnor UO_2169 (O_2169,N_16668,N_15710);
xor UO_2170 (O_2170,N_18141,N_18678);
and UO_2171 (O_2171,N_18697,N_17501);
xor UO_2172 (O_2172,N_19011,N_18503);
or UO_2173 (O_2173,N_18143,N_15142);
nor UO_2174 (O_2174,N_16765,N_16606);
nand UO_2175 (O_2175,N_19417,N_16985);
nand UO_2176 (O_2176,N_17158,N_18012);
nor UO_2177 (O_2177,N_19670,N_17818);
nand UO_2178 (O_2178,N_18979,N_16732);
xnor UO_2179 (O_2179,N_19706,N_17723);
nor UO_2180 (O_2180,N_17347,N_19378);
nor UO_2181 (O_2181,N_16326,N_19881);
nand UO_2182 (O_2182,N_17167,N_17452);
nand UO_2183 (O_2183,N_19034,N_16964);
or UO_2184 (O_2184,N_17465,N_17999);
nor UO_2185 (O_2185,N_15445,N_16834);
nand UO_2186 (O_2186,N_16209,N_15172);
or UO_2187 (O_2187,N_16319,N_19222);
nand UO_2188 (O_2188,N_17533,N_17985);
xnor UO_2189 (O_2189,N_15050,N_15843);
and UO_2190 (O_2190,N_18914,N_18341);
nor UO_2191 (O_2191,N_19144,N_19231);
or UO_2192 (O_2192,N_16365,N_19718);
xor UO_2193 (O_2193,N_18072,N_16660);
nand UO_2194 (O_2194,N_19617,N_19235);
nor UO_2195 (O_2195,N_19333,N_15801);
or UO_2196 (O_2196,N_15372,N_19533);
nand UO_2197 (O_2197,N_17470,N_18874);
or UO_2198 (O_2198,N_17040,N_18884);
and UO_2199 (O_2199,N_18959,N_17405);
nor UO_2200 (O_2200,N_16386,N_19884);
and UO_2201 (O_2201,N_18841,N_19664);
or UO_2202 (O_2202,N_16290,N_16406);
nand UO_2203 (O_2203,N_18311,N_17996);
xnor UO_2204 (O_2204,N_16638,N_17046);
nor UO_2205 (O_2205,N_15631,N_16772);
nor UO_2206 (O_2206,N_16249,N_19083);
and UO_2207 (O_2207,N_18095,N_16268);
and UO_2208 (O_2208,N_16619,N_15973);
xor UO_2209 (O_2209,N_19486,N_19742);
and UO_2210 (O_2210,N_15624,N_17042);
and UO_2211 (O_2211,N_15328,N_16364);
or UO_2212 (O_2212,N_17494,N_15702);
xnor UO_2213 (O_2213,N_15701,N_18543);
or UO_2214 (O_2214,N_18743,N_16233);
and UO_2215 (O_2215,N_16201,N_16681);
nor UO_2216 (O_2216,N_19114,N_19981);
nand UO_2217 (O_2217,N_17524,N_18176);
and UO_2218 (O_2218,N_18615,N_16318);
nand UO_2219 (O_2219,N_16925,N_17261);
xor UO_2220 (O_2220,N_19699,N_18726);
xnor UO_2221 (O_2221,N_17211,N_18919);
nand UO_2222 (O_2222,N_19883,N_19605);
and UO_2223 (O_2223,N_16529,N_19582);
nand UO_2224 (O_2224,N_18120,N_15663);
nand UO_2225 (O_2225,N_19322,N_19919);
xnor UO_2226 (O_2226,N_15968,N_19426);
nor UO_2227 (O_2227,N_15814,N_16609);
or UO_2228 (O_2228,N_16114,N_16495);
nand UO_2229 (O_2229,N_18988,N_17780);
and UO_2230 (O_2230,N_19094,N_19345);
and UO_2231 (O_2231,N_15587,N_16870);
and UO_2232 (O_2232,N_15147,N_15992);
nor UO_2233 (O_2233,N_16191,N_17558);
and UO_2234 (O_2234,N_18846,N_18860);
nand UO_2235 (O_2235,N_15927,N_18958);
and UO_2236 (O_2236,N_16927,N_16127);
or UO_2237 (O_2237,N_18545,N_16187);
nand UO_2238 (O_2238,N_15990,N_17640);
and UO_2239 (O_2239,N_19687,N_15415);
nand UO_2240 (O_2240,N_15633,N_16353);
nor UO_2241 (O_2241,N_19033,N_17872);
or UO_2242 (O_2242,N_15845,N_18760);
nand UO_2243 (O_2243,N_17702,N_19814);
nand UO_2244 (O_2244,N_16351,N_16112);
xor UO_2245 (O_2245,N_18759,N_15989);
and UO_2246 (O_2246,N_17924,N_18260);
nor UO_2247 (O_2247,N_18813,N_19275);
or UO_2248 (O_2248,N_15901,N_17245);
or UO_2249 (O_2249,N_18433,N_15068);
nor UO_2250 (O_2250,N_17744,N_16900);
and UO_2251 (O_2251,N_15264,N_15112);
nand UO_2252 (O_2252,N_19323,N_18835);
xor UO_2253 (O_2253,N_18815,N_19279);
or UO_2254 (O_2254,N_16410,N_18452);
xnor UO_2255 (O_2255,N_18574,N_18275);
xor UO_2256 (O_2256,N_16836,N_18969);
or UO_2257 (O_2257,N_15855,N_17111);
xnor UO_2258 (O_2258,N_16193,N_15024);
xnor UO_2259 (O_2259,N_18366,N_15712);
or UO_2260 (O_2260,N_17341,N_18588);
xnor UO_2261 (O_2261,N_17895,N_18714);
nor UO_2262 (O_2262,N_16051,N_17068);
nand UO_2263 (O_2263,N_18810,N_15681);
nand UO_2264 (O_2264,N_18602,N_19544);
nor UO_2265 (O_2265,N_16556,N_17120);
and UO_2266 (O_2266,N_18780,N_16003);
and UO_2267 (O_2267,N_18430,N_19386);
nor UO_2268 (O_2268,N_17003,N_16200);
nor UO_2269 (O_2269,N_18404,N_19937);
xnor UO_2270 (O_2270,N_19785,N_15687);
and UO_2271 (O_2271,N_19358,N_15660);
and UO_2272 (O_2272,N_17140,N_18824);
nand UO_2273 (O_2273,N_15880,N_15153);
and UO_2274 (O_2274,N_19534,N_15461);
and UO_2275 (O_2275,N_19923,N_18107);
xor UO_2276 (O_2276,N_16479,N_17308);
nand UO_2277 (O_2277,N_17522,N_19932);
nor UO_2278 (O_2278,N_17610,N_18945);
or UO_2279 (O_2279,N_17020,N_18046);
xnor UO_2280 (O_2280,N_17295,N_17667);
nand UO_2281 (O_2281,N_15542,N_18641);
and UO_2282 (O_2282,N_19089,N_17058);
nor UO_2283 (O_2283,N_16055,N_18044);
or UO_2284 (O_2284,N_17086,N_18535);
nand UO_2285 (O_2285,N_17515,N_18947);
and UO_2286 (O_2286,N_16424,N_15511);
xor UO_2287 (O_2287,N_18625,N_19234);
or UO_2288 (O_2288,N_19755,N_19873);
nand UO_2289 (O_2289,N_18599,N_16831);
nor UO_2290 (O_2290,N_15280,N_19403);
xnor UO_2291 (O_2291,N_17334,N_16347);
or UO_2292 (O_2292,N_19273,N_19523);
xnor UO_2293 (O_2293,N_18376,N_17735);
xor UO_2294 (O_2294,N_17054,N_16392);
xor UO_2295 (O_2295,N_15365,N_19387);
nand UO_2296 (O_2296,N_15067,N_16150);
nand UO_2297 (O_2297,N_16231,N_15966);
xor UO_2298 (O_2298,N_15119,N_16800);
nand UO_2299 (O_2299,N_15069,N_19629);
and UO_2300 (O_2300,N_16059,N_18041);
and UO_2301 (O_2301,N_17962,N_17549);
nor UO_2302 (O_2302,N_19053,N_15059);
nand UO_2303 (O_2303,N_17035,N_15683);
nand UO_2304 (O_2304,N_17149,N_15524);
or UO_2305 (O_2305,N_16880,N_18506);
xnor UO_2306 (O_2306,N_15107,N_17584);
or UO_2307 (O_2307,N_17791,N_19301);
nand UO_2308 (O_2308,N_19746,N_16759);
nor UO_2309 (O_2309,N_18112,N_15376);
or UO_2310 (O_2310,N_16370,N_16615);
or UO_2311 (O_2311,N_17044,N_17207);
nand UO_2312 (O_2312,N_17964,N_16743);
and UO_2313 (O_2313,N_18195,N_15655);
nand UO_2314 (O_2314,N_19859,N_17765);
nand UO_2315 (O_2315,N_16890,N_19040);
nand UO_2316 (O_2316,N_15052,N_18525);
and UO_2317 (O_2317,N_17349,N_19140);
nand UO_2318 (O_2318,N_19538,N_17208);
nor UO_2319 (O_2319,N_15072,N_17209);
xor UO_2320 (O_2320,N_16667,N_19974);
nand UO_2321 (O_2321,N_18458,N_17503);
nand UO_2322 (O_2322,N_16333,N_19113);
nor UO_2323 (O_2323,N_17806,N_19126);
or UO_2324 (O_2324,N_19793,N_18712);
nand UO_2325 (O_2325,N_18941,N_16272);
or UO_2326 (O_2326,N_18368,N_15838);
nand UO_2327 (O_2327,N_18895,N_15140);
xor UO_2328 (O_2328,N_19610,N_16307);
and UO_2329 (O_2329,N_16482,N_19145);
xor UO_2330 (O_2330,N_16565,N_19248);
nor UO_2331 (O_2331,N_16788,N_19721);
nor UO_2332 (O_2332,N_17106,N_19877);
xor UO_2333 (O_2333,N_18611,N_15241);
nand UO_2334 (O_2334,N_18956,N_17036);
nand UO_2335 (O_2335,N_19803,N_16533);
and UO_2336 (O_2336,N_16372,N_17377);
or UO_2337 (O_2337,N_19700,N_17309);
nand UO_2338 (O_2338,N_16133,N_15214);
and UO_2339 (O_2339,N_18374,N_17319);
nor UO_2340 (O_2340,N_15637,N_18532);
nand UO_2341 (O_2341,N_18591,N_15764);
or UO_2342 (O_2342,N_15536,N_16030);
nor UO_2343 (O_2343,N_15991,N_16278);
nand UO_2344 (O_2344,N_18788,N_19237);
and UO_2345 (O_2345,N_18610,N_18765);
and UO_2346 (O_2346,N_15016,N_17973);
or UO_2347 (O_2347,N_15532,N_19707);
nand UO_2348 (O_2348,N_15608,N_16446);
or UO_2349 (O_2349,N_15384,N_16488);
nor UO_2350 (O_2350,N_17288,N_19366);
nand UO_2351 (O_2351,N_19949,N_17407);
nor UO_2352 (O_2352,N_16863,N_15856);
nor UO_2353 (O_2353,N_17170,N_16460);
or UO_2354 (O_2354,N_19470,N_16227);
or UO_2355 (O_2355,N_19824,N_15020);
and UO_2356 (O_2356,N_15456,N_15355);
and UO_2357 (O_2357,N_16662,N_19737);
xor UO_2358 (O_2358,N_15462,N_19288);
nand UO_2359 (O_2359,N_17060,N_19121);
nor UO_2360 (O_2360,N_16591,N_17266);
nor UO_2361 (O_2361,N_18843,N_18578);
and UO_2362 (O_2362,N_19506,N_16464);
nor UO_2363 (O_2363,N_15090,N_15449);
or UO_2364 (O_2364,N_17800,N_19321);
and UO_2365 (O_2365,N_16597,N_18750);
nand UO_2366 (O_2366,N_15958,N_15743);
or UO_2367 (O_2367,N_15707,N_17034);
xnor UO_2368 (O_2368,N_18654,N_15715);
xor UO_2369 (O_2369,N_15102,N_18316);
and UO_2370 (O_2370,N_19702,N_18667);
or UO_2371 (O_2371,N_19283,N_18596);
xnor UO_2372 (O_2372,N_18623,N_19133);
or UO_2373 (O_2373,N_17008,N_16346);
nand UO_2374 (O_2374,N_17676,N_19017);
nor UO_2375 (O_2375,N_18082,N_17330);
and UO_2376 (O_2376,N_15941,N_16513);
nor UO_2377 (O_2377,N_18004,N_15975);
or UO_2378 (O_2378,N_18088,N_19047);
nand UO_2379 (O_2379,N_18859,N_17825);
nor UO_2380 (O_2380,N_16952,N_15500);
and UO_2381 (O_2381,N_19602,N_16980);
or UO_2382 (O_2382,N_15525,N_17088);
nor UO_2383 (O_2383,N_16060,N_18375);
xor UO_2384 (O_2384,N_15819,N_19865);
and UO_2385 (O_2385,N_17613,N_17642);
or UO_2386 (O_2386,N_18620,N_19267);
nand UO_2387 (O_2387,N_18160,N_18886);
nor UO_2388 (O_2388,N_16121,N_16377);
nor UO_2389 (O_2389,N_15860,N_17972);
and UO_2390 (O_2390,N_16761,N_16276);
nand UO_2391 (O_2391,N_15639,N_19817);
xnor UO_2392 (O_2392,N_15942,N_18396);
and UO_2393 (O_2393,N_17430,N_16665);
xor UO_2394 (O_2394,N_16064,N_15191);
xnor UO_2395 (O_2395,N_17074,N_17521);
or UO_2396 (O_2396,N_15872,N_16445);
nor UO_2397 (O_2397,N_18244,N_15170);
xnor UO_2398 (O_2398,N_18995,N_15649);
xnor UO_2399 (O_2399,N_17934,N_15705);
xnor UO_2400 (O_2400,N_15675,N_19002);
nand UO_2401 (O_2401,N_16816,N_19031);
nor UO_2402 (O_2402,N_19221,N_16316);
nor UO_2403 (O_2403,N_18117,N_17705);
nand UO_2404 (O_2404,N_19953,N_17041);
or UO_2405 (O_2405,N_19562,N_16568);
nand UO_2406 (O_2406,N_17257,N_17290);
or UO_2407 (O_2407,N_17795,N_15473);
nand UO_2408 (O_2408,N_17687,N_15318);
or UO_2409 (O_2409,N_16103,N_18581);
xnor UO_2410 (O_2410,N_18245,N_18315);
or UO_2411 (O_2411,N_15033,N_19344);
or UO_2412 (O_2412,N_19100,N_15115);
or UO_2413 (O_2413,N_18994,N_15616);
xnor UO_2414 (O_2414,N_16988,N_17175);
nor UO_2415 (O_2415,N_19622,N_16118);
nand UO_2416 (O_2416,N_15602,N_18564);
or UO_2417 (O_2417,N_15014,N_18405);
or UO_2418 (O_2418,N_16130,N_18355);
or UO_2419 (O_2419,N_16738,N_18634);
or UO_2420 (O_2420,N_15139,N_17760);
nand UO_2421 (O_2421,N_18468,N_17413);
xnor UO_2422 (O_2422,N_15729,N_19580);
or UO_2423 (O_2423,N_19933,N_19554);
or UO_2424 (O_2424,N_15885,N_17547);
and UO_2425 (O_2425,N_17861,N_17222);
nand UO_2426 (O_2426,N_16100,N_19796);
or UO_2427 (O_2427,N_17990,N_17053);
nor UO_2428 (O_2428,N_19257,N_15198);
and UO_2429 (O_2429,N_18457,N_17115);
or UO_2430 (O_2430,N_16066,N_17352);
and UO_2431 (O_2431,N_15896,N_18908);
nor UO_2432 (O_2432,N_17982,N_19684);
nor UO_2433 (O_2433,N_19569,N_15735);
or UO_2434 (O_2434,N_19765,N_17530);
nand UO_2435 (O_2435,N_15564,N_18280);
xor UO_2436 (O_2436,N_19616,N_15432);
or UO_2437 (O_2437,N_17331,N_15578);
and UO_2438 (O_2438,N_16869,N_17831);
nand UO_2439 (O_2439,N_17213,N_17684);
nand UO_2440 (O_2440,N_18398,N_19590);
xor UO_2441 (O_2441,N_16046,N_17926);
or UO_2442 (O_2442,N_19192,N_16876);
and UO_2443 (O_2443,N_19963,N_19369);
and UO_2444 (O_2444,N_17782,N_17528);
or UO_2445 (O_2445,N_17123,N_18684);
xnor UO_2446 (O_2446,N_15803,N_19455);
and UO_2447 (O_2447,N_18550,N_17052);
xor UO_2448 (O_2448,N_18459,N_15620);
or UO_2449 (O_2449,N_16722,N_19593);
and UO_2450 (O_2450,N_18388,N_18504);
nand UO_2451 (O_2451,N_19439,N_18754);
nor UO_2452 (O_2452,N_19677,N_15733);
nand UO_2453 (O_2453,N_17660,N_19068);
or UO_2454 (O_2454,N_15228,N_15486);
and UO_2455 (O_2455,N_17583,N_16251);
xor UO_2456 (O_2456,N_19614,N_15206);
or UO_2457 (O_2457,N_19734,N_16053);
xor UO_2458 (O_2458,N_18932,N_19434);
nor UO_2459 (O_2459,N_18756,N_17983);
nor UO_2460 (O_2460,N_16956,N_17912);
xor UO_2461 (O_2461,N_17481,N_16700);
nor UO_2462 (O_2462,N_18000,N_17328);
nor UO_2463 (O_2463,N_17322,N_18685);
and UO_2464 (O_2464,N_17383,N_19504);
xor UO_2465 (O_2465,N_15779,N_16020);
nand UO_2466 (O_2466,N_16924,N_18340);
xor UO_2467 (O_2467,N_17419,N_17043);
xor UO_2468 (O_2468,N_16550,N_17176);
or UO_2469 (O_2469,N_16248,N_16023);
nor UO_2470 (O_2470,N_18114,N_15322);
and UO_2471 (O_2471,N_15736,N_15373);
or UO_2472 (O_2472,N_16779,N_15493);
nand UO_2473 (O_2473,N_16449,N_17375);
xor UO_2474 (O_2474,N_19510,N_16686);
nand UO_2475 (O_2475,N_17372,N_17297);
and UO_2476 (O_2476,N_18424,N_15239);
xor UO_2477 (O_2477,N_17553,N_15709);
nor UO_2478 (O_2478,N_16113,N_19111);
and UO_2479 (O_2479,N_16741,N_19415);
and UO_2480 (O_2480,N_16569,N_16454);
xor UO_2481 (O_2481,N_16633,N_15077);
nand UO_2482 (O_2482,N_15309,N_19206);
or UO_2483 (O_2483,N_19270,N_15406);
and UO_2484 (O_2484,N_15138,N_19365);
and UO_2485 (O_2485,N_17461,N_16196);
or UO_2486 (O_2486,N_16867,N_17649);
or UO_2487 (O_2487,N_19456,N_17360);
xor UO_2488 (O_2488,N_19678,N_16695);
or UO_2489 (O_2489,N_19513,N_15217);
nand UO_2490 (O_2490,N_15671,N_15480);
xnor UO_2491 (O_2491,N_19566,N_15833);
or UO_2492 (O_2492,N_19961,N_18291);
nand UO_2493 (O_2493,N_15535,N_18869);
xor UO_2494 (O_2494,N_15126,N_18515);
and UO_2495 (O_2495,N_16814,N_19577);
and UO_2496 (O_2496,N_19284,N_16905);
nor UO_2497 (O_2497,N_19794,N_18893);
xor UO_2498 (O_2498,N_16581,N_17846);
and UO_2499 (O_2499,N_16962,N_17862);
endmodule