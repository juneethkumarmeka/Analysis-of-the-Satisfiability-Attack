module basic_1500_15000_2000_10_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_863,In_1116);
and U1 (N_1,In_1248,In_1444);
and U2 (N_2,In_208,In_521);
and U3 (N_3,In_1351,In_670);
and U4 (N_4,In_390,In_1000);
or U5 (N_5,In_1473,In_482);
or U6 (N_6,In_150,In_1382);
and U7 (N_7,In_745,In_725);
nand U8 (N_8,In_317,In_1172);
xnor U9 (N_9,In_665,In_251);
xnor U10 (N_10,In_597,In_420);
and U11 (N_11,In_851,In_905);
and U12 (N_12,In_447,In_1145);
or U13 (N_13,In_1421,In_331);
and U14 (N_14,In_523,In_51);
nor U15 (N_15,In_1061,In_12);
nor U16 (N_16,In_1214,In_245);
and U17 (N_17,In_387,In_1235);
nand U18 (N_18,In_1087,In_256);
nor U19 (N_19,In_1494,In_835);
or U20 (N_20,In_1230,In_1260);
or U21 (N_21,In_781,In_288);
nor U22 (N_22,In_1150,In_870);
nand U23 (N_23,In_549,In_1224);
or U24 (N_24,In_620,In_684);
nor U25 (N_25,In_797,In_363);
and U26 (N_26,In_398,In_951);
nor U27 (N_27,In_747,In_201);
or U28 (N_28,In_1204,In_1162);
and U29 (N_29,In_602,In_623);
xor U30 (N_30,In_581,In_31);
nor U31 (N_31,In_27,In_1328);
xnor U32 (N_32,In_802,In_667);
or U33 (N_33,In_631,In_1412);
xor U34 (N_34,In_71,In_485);
and U35 (N_35,In_1231,In_1472);
or U36 (N_36,In_715,In_593);
or U37 (N_37,In_840,In_646);
nor U38 (N_38,In_1269,In_791);
xor U39 (N_39,In_176,In_1228);
and U40 (N_40,In_663,In_1447);
xnor U41 (N_41,In_780,In_926);
or U42 (N_42,In_1071,In_1176);
nor U43 (N_43,In_1363,In_291);
nand U44 (N_44,In_1155,In_768);
or U45 (N_45,In_461,In_930);
nand U46 (N_46,In_968,In_472);
nand U47 (N_47,In_20,In_462);
nand U48 (N_48,In_592,In_219);
nand U49 (N_49,In_458,In_1372);
and U50 (N_50,In_1487,In_757);
and U51 (N_51,In_992,In_850);
and U52 (N_52,In_1140,In_721);
nand U53 (N_53,In_1385,In_1236);
nand U54 (N_54,In_87,In_24);
and U55 (N_55,In_407,In_409);
nor U56 (N_56,In_1278,In_22);
or U57 (N_57,In_1316,In_531);
nor U58 (N_58,In_1416,In_886);
nand U59 (N_59,In_321,In_1027);
nand U60 (N_60,In_855,In_1126);
or U61 (N_61,In_963,In_869);
nand U62 (N_62,In_465,In_1080);
and U63 (N_63,In_532,In_46);
nor U64 (N_64,In_1139,In_805);
nand U65 (N_65,In_812,In_308);
nand U66 (N_66,In_625,In_591);
nand U67 (N_67,In_217,In_1264);
and U68 (N_68,In_1420,In_1350);
or U69 (N_69,In_686,In_235);
nand U70 (N_70,In_243,In_421);
nand U71 (N_71,In_312,In_1059);
or U72 (N_72,In_494,In_873);
nand U73 (N_73,In_1365,In_867);
and U74 (N_74,In_1037,In_1057);
or U75 (N_75,In_1445,In_691);
nand U76 (N_76,In_965,In_538);
xnor U77 (N_77,In_1356,In_760);
xor U78 (N_78,In_698,In_818);
or U79 (N_79,In_400,In_1299);
nand U80 (N_80,In_1418,In_18);
nand U81 (N_81,In_191,In_1040);
and U82 (N_82,In_1178,In_672);
or U83 (N_83,In_52,In_103);
and U84 (N_84,In_1437,In_1068);
and U85 (N_85,In_1076,In_1318);
nor U86 (N_86,In_634,In_1022);
and U87 (N_87,In_222,In_1098);
or U88 (N_88,In_875,In_542);
nor U89 (N_89,In_1013,In_811);
or U90 (N_90,In_594,In_403);
and U91 (N_91,In_975,In_1435);
nand U92 (N_92,In_1451,In_799);
or U93 (N_93,In_834,In_1307);
or U94 (N_94,In_789,In_1294);
and U95 (N_95,In_1141,In_1067);
or U96 (N_96,In_709,In_260);
and U97 (N_97,In_493,In_34);
nor U98 (N_98,In_211,In_419);
or U99 (N_99,In_615,In_1189);
nand U100 (N_100,In_1404,In_837);
xor U101 (N_101,In_1481,In_983);
nor U102 (N_102,In_771,In_174);
xor U103 (N_103,In_1195,In_434);
and U104 (N_104,In_268,In_856);
xor U105 (N_105,In_242,In_406);
and U106 (N_106,In_184,In_891);
and U107 (N_107,In_569,In_1092);
nor U108 (N_108,In_1193,In_1387);
xnor U109 (N_109,In_329,In_806);
and U110 (N_110,In_72,In_1099);
or U111 (N_111,In_498,In_512);
or U112 (N_112,In_756,In_673);
nand U113 (N_113,In_880,In_861);
or U114 (N_114,In_391,In_820);
and U115 (N_115,In_383,In_127);
xor U116 (N_116,In_415,In_1005);
and U117 (N_117,In_207,In_53);
xnor U118 (N_118,In_294,In_567);
nand U119 (N_119,In_919,In_755);
and U120 (N_120,In_682,In_727);
nand U121 (N_121,In_169,In_636);
and U122 (N_122,In_69,In_733);
and U123 (N_123,In_1077,In_1241);
and U124 (N_124,In_1011,In_19);
or U125 (N_125,In_424,In_871);
nand U126 (N_126,In_293,In_442);
nor U127 (N_127,In_492,In_1492);
and U128 (N_128,In_681,In_1237);
and U129 (N_129,In_1456,In_1053);
nor U130 (N_130,In_888,In_689);
and U131 (N_131,In_878,In_642);
or U132 (N_132,In_601,In_111);
xor U133 (N_133,In_254,In_647);
nor U134 (N_134,In_119,In_428);
or U135 (N_135,In_333,In_860);
nand U136 (N_136,In_1166,In_833);
xnor U137 (N_137,In_612,In_423);
and U138 (N_138,In_702,In_964);
and U139 (N_139,In_595,In_1215);
nor U140 (N_140,In_884,In_1045);
or U141 (N_141,In_785,In_379);
xnor U142 (N_142,In_1253,In_801);
and U143 (N_143,In_1428,In_1336);
nor U144 (N_144,In_1280,In_1194);
or U145 (N_145,In_788,In_611);
and U146 (N_146,In_1100,In_556);
nor U147 (N_147,In_352,In_987);
or U148 (N_148,In_345,In_528);
nor U149 (N_149,In_619,In_438);
nor U150 (N_150,In_326,In_373);
or U151 (N_151,In_814,In_659);
and U152 (N_152,In_603,In_927);
and U153 (N_153,In_1314,In_393);
or U154 (N_154,In_1374,In_1199);
nand U155 (N_155,In_454,In_325);
nor U156 (N_156,In_165,In_1364);
nor U157 (N_157,In_969,In_1273);
nor U158 (N_158,In_418,In_1020);
nor U159 (N_159,In_874,In_94);
and U160 (N_160,In_1168,In_1149);
nand U161 (N_161,In_262,In_209);
and U162 (N_162,In_147,In_649);
or U163 (N_163,In_1466,In_144);
nand U164 (N_164,In_680,In_723);
nor U165 (N_165,In_82,In_705);
xnor U166 (N_166,In_1187,In_309);
xor U167 (N_167,In_269,In_481);
or U168 (N_168,In_365,In_893);
or U169 (N_169,In_1008,In_513);
and U170 (N_170,In_526,In_118);
nand U171 (N_171,In_1030,In_998);
nor U172 (N_172,In_414,In_822);
nand U173 (N_173,In_1287,In_1300);
and U174 (N_174,In_1461,In_131);
or U175 (N_175,In_1165,In_44);
nand U176 (N_176,In_1433,In_920);
nand U177 (N_177,In_1422,In_786);
and U178 (N_178,In_714,In_979);
nor U179 (N_179,In_938,In_1380);
or U180 (N_180,In_4,In_973);
or U181 (N_181,In_707,In_123);
or U182 (N_182,In_1198,In_562);
nor U183 (N_183,In_218,In_941);
and U184 (N_184,In_370,In_300);
xor U185 (N_185,In_784,In_782);
and U186 (N_186,In_807,In_947);
and U187 (N_187,In_110,In_502);
and U188 (N_188,In_1448,In_519);
or U189 (N_189,In_988,In_399);
or U190 (N_190,In_486,In_233);
xnor U191 (N_191,In_922,In_130);
or U192 (N_192,In_1467,In_1396);
nor U193 (N_193,In_183,In_1244);
xnor U194 (N_194,In_1001,In_1170);
and U195 (N_195,In_923,In_463);
and U196 (N_196,In_1026,In_1161);
nor U197 (N_197,In_221,In_1460);
nor U198 (N_198,In_479,In_473);
xor U199 (N_199,In_607,In_742);
and U200 (N_200,In_1086,In_1229);
nor U201 (N_201,In_292,In_999);
nand U202 (N_202,In_152,In_314);
xnor U203 (N_203,In_720,In_831);
nand U204 (N_204,In_410,In_982);
and U205 (N_205,In_662,In_441);
nand U206 (N_206,In_739,In_1185);
xor U207 (N_207,In_496,In_357);
nand U208 (N_208,In_948,In_204);
or U209 (N_209,In_1180,In_1296);
and U210 (N_210,In_605,In_1457);
nand U211 (N_211,In_1,In_1257);
xor U212 (N_212,In_263,In_1075);
nor U213 (N_213,In_1325,In_358);
or U214 (N_214,In_859,In_692);
nor U215 (N_215,In_1388,In_303);
or U216 (N_216,In_589,In_676);
and U217 (N_217,In_772,In_5);
nand U218 (N_218,In_192,In_289);
nor U219 (N_219,In_576,In_232);
or U220 (N_220,In_1003,In_145);
nand U221 (N_221,In_1341,In_1312);
and U222 (N_222,In_841,In_1393);
nor U223 (N_223,In_36,In_70);
nand U224 (N_224,In_42,In_285);
nand U225 (N_225,In_1154,In_981);
or U226 (N_226,In_1277,In_344);
nand U227 (N_227,In_1190,In_558);
nor U228 (N_228,In_181,In_536);
or U229 (N_229,In_537,In_1137);
nand U230 (N_230,In_1389,In_504);
and U231 (N_231,In_474,In_560);
or U232 (N_232,In_1063,In_223);
nand U233 (N_233,In_1018,In_25);
xor U234 (N_234,In_741,In_779);
or U235 (N_235,In_1395,In_1345);
nor U236 (N_236,In_1271,In_89);
nor U237 (N_237,In_656,In_417);
nor U238 (N_238,In_777,In_1335);
nand U239 (N_239,In_350,In_330);
nand U240 (N_240,In_1223,In_641);
or U241 (N_241,In_41,In_1413);
and U242 (N_242,In_1147,In_316);
nor U243 (N_243,In_224,In_477);
nand U244 (N_244,In_578,In_516);
nor U245 (N_245,In_252,In_1376);
or U246 (N_246,In_1475,In_92);
or U247 (N_247,In_543,In_896);
or U248 (N_248,In_1232,In_1004);
and U249 (N_249,In_1101,In_135);
nor U250 (N_250,In_586,In_246);
nand U251 (N_251,In_228,In_1169);
and U252 (N_252,In_501,In_206);
nor U253 (N_253,In_313,In_753);
xnor U254 (N_254,In_1471,In_1245);
nor U255 (N_255,In_187,In_138);
nand U256 (N_256,In_1156,In_1306);
xor U257 (N_257,In_237,In_1219);
and U258 (N_258,In_264,In_270);
nor U259 (N_259,In_770,In_311);
nor U260 (N_260,In_155,In_540);
or U261 (N_261,In_448,In_1405);
and U262 (N_262,In_962,In_1483);
nor U263 (N_263,In_1449,In_1305);
and U264 (N_264,In_186,In_397);
nand U265 (N_265,In_276,In_813);
nand U266 (N_266,In_1209,In_1477);
nand U267 (N_267,In_160,In_126);
or U268 (N_268,In_342,In_510);
and U269 (N_269,In_1375,In_136);
or U270 (N_270,In_487,In_584);
and U271 (N_271,In_825,In_112);
xnor U272 (N_272,In_1031,In_28);
nor U273 (N_273,In_335,In_710);
nand U274 (N_274,In_552,In_57);
nand U275 (N_275,In_1122,In_956);
and U276 (N_276,In_1208,In_445);
nand U277 (N_277,In_240,In_1286);
nor U278 (N_278,In_958,In_76);
xor U279 (N_279,In_1485,In_944);
nand U280 (N_280,In_748,In_1390);
or U281 (N_281,In_1465,In_1233);
or U282 (N_282,In_1346,In_328);
nor U283 (N_283,In_1499,In_713);
xor U284 (N_284,In_1359,In_161);
nor U285 (N_285,In_1173,In_1213);
or U286 (N_286,In_1496,In_1119);
or U287 (N_287,In_1308,In_568);
nand U288 (N_288,In_514,In_283);
or U289 (N_289,In_253,In_480);
and U290 (N_290,In_933,In_1491);
or U291 (N_291,In_509,In_347);
nand U292 (N_292,In_1054,In_1403);
and U293 (N_293,In_384,In_341);
nand U294 (N_294,In_942,In_970);
nand U295 (N_295,In_386,In_1065);
nand U296 (N_296,In_1398,In_1157);
nand U297 (N_297,In_1073,In_443);
nor U298 (N_298,In_1493,In_173);
nor U299 (N_299,In_1047,In_376);
nor U300 (N_300,In_96,In_1041);
and U301 (N_301,In_1486,In_868);
nand U302 (N_302,In_1497,In_431);
and U303 (N_303,In_736,In_1419);
or U304 (N_304,In_348,In_669);
nor U305 (N_305,In_250,In_892);
or U306 (N_306,In_915,In_395);
nor U307 (N_307,In_225,In_1247);
nor U308 (N_308,In_1109,In_364);
nor U309 (N_309,In_2,In_282);
nand U310 (N_310,In_1105,In_1112);
or U311 (N_311,In_449,In_547);
xor U312 (N_312,In_166,In_1361);
xor U313 (N_313,In_703,In_924);
nand U314 (N_314,In_1323,In_1039);
nand U315 (N_315,In_769,In_446);
or U316 (N_316,In_1117,In_643);
nand U317 (N_317,In_404,In_1329);
or U318 (N_318,In_320,In_887);
nor U319 (N_319,In_453,In_78);
nand U320 (N_320,In_864,In_83);
nand U321 (N_321,In_1060,In_815);
nor U322 (N_322,In_1453,In_142);
nor U323 (N_323,In_56,In_1250);
nor U324 (N_324,In_29,In_62);
or U325 (N_325,In_66,In_14);
or U326 (N_326,In_792,In_503);
xnor U327 (N_327,In_137,In_995);
or U328 (N_328,In_1094,In_1479);
nand U329 (N_329,In_978,In_1123);
or U330 (N_330,In_129,In_158);
nor U331 (N_331,In_939,In_1354);
or U332 (N_332,In_737,In_1035);
nand U333 (N_333,In_534,In_13);
nand U334 (N_334,In_630,In_912);
or U335 (N_335,In_889,In_832);
and U336 (N_336,In_554,In_1164);
nand U337 (N_337,In_381,In_1009);
nor U338 (N_338,In_683,In_382);
nand U339 (N_339,In_359,In_84);
nand U340 (N_340,In_934,In_1295);
nor U341 (N_341,In_1051,In_296);
nor U342 (N_342,In_993,In_1095);
xor U343 (N_343,In_258,In_249);
nand U344 (N_344,In_93,In_1128);
and U345 (N_345,In_708,In_1344);
nor U346 (N_346,In_1282,In_179);
or U347 (N_347,In_315,In_203);
xor U348 (N_348,In_172,In_1196);
nor U349 (N_349,In_1072,In_125);
or U350 (N_350,In_1489,In_1043);
or U351 (N_351,In_946,In_336);
nor U352 (N_352,In_377,In_1333);
and U353 (N_353,In_214,In_356);
xor U354 (N_354,In_1238,In_729);
and U355 (N_355,In_844,In_1070);
or U356 (N_356,In_566,In_764);
nand U357 (N_357,In_724,In_1243);
nor U358 (N_358,In_338,In_695);
nor U359 (N_359,In_1339,In_1242);
nand U360 (N_360,In_1066,In_101);
nor U361 (N_361,In_1177,In_728);
and U362 (N_362,In_437,In_985);
and U363 (N_363,In_193,In_925);
or U364 (N_364,In_162,In_1482);
xnor U365 (N_365,In_425,In_1021);
nor U366 (N_366,In_932,In_3);
nand U367 (N_367,In_1462,In_1332);
nand U368 (N_368,In_456,In_396);
and U369 (N_369,In_1082,In_64);
nand U370 (N_370,In_1484,In_865);
and U371 (N_371,In_694,In_73);
nand U372 (N_372,In_1124,In_272);
xnor U373 (N_373,In_1091,In_750);
or U374 (N_374,In_106,In_937);
nand U375 (N_375,In_1221,In_1337);
and U376 (N_376,In_1069,In_1401);
nand U377 (N_377,In_986,In_1006);
nand U378 (N_378,In_1443,In_685);
nand U379 (N_379,In_522,In_353);
nor U380 (N_380,In_967,In_133);
or U381 (N_381,In_128,In_1476);
and U382 (N_382,In_796,In_427);
or U383 (N_383,In_327,In_115);
or U384 (N_384,In_32,In_862);
xnor U385 (N_385,In_824,In_239);
nor U386 (N_386,In_1304,In_744);
nand U387 (N_387,In_1158,In_234);
xnor U388 (N_388,In_1352,In_95);
or U389 (N_389,In_433,In_1136);
or U390 (N_390,In_557,In_402);
xnor U391 (N_391,In_148,In_977);
xor U392 (N_392,In_687,In_1255);
nand U393 (N_393,In_11,In_1015);
and U394 (N_394,In_238,In_900);
and U395 (N_395,In_306,In_241);
or U396 (N_396,In_38,In_972);
and U397 (N_397,In_26,In_104);
and U398 (N_398,In_277,In_1159);
nor U399 (N_399,In_196,In_337);
or U400 (N_400,In_650,In_185);
nand U401 (N_401,In_787,In_700);
or U402 (N_402,In_199,In_518);
nor U403 (N_403,In_717,In_608);
and U404 (N_404,In_99,In_153);
or U405 (N_405,In_284,In_483);
or U406 (N_406,In_897,In_1267);
nor U407 (N_407,In_100,In_1417);
nor U408 (N_408,In_960,In_1407);
nand U409 (N_409,In_75,In_1016);
nor U410 (N_410,In_244,In_940);
nor U411 (N_411,In_1202,In_163);
xnor U412 (N_412,In_1118,In_1406);
and U413 (N_413,In_819,In_1355);
nand U414 (N_414,In_170,In_140);
nand U415 (N_415,In_0,In_810);
or U416 (N_416,In_935,In_30);
or U417 (N_417,In_1254,In_866);
or U418 (N_418,In_902,In_1302);
nor U419 (N_419,In_91,In_735);
and U420 (N_420,In_911,In_1490);
nor U421 (N_421,In_74,In_846);
nand U422 (N_422,In_1024,In_936);
and U423 (N_423,In_658,In_1369);
xnor U424 (N_424,In_1120,In_1285);
or U425 (N_425,In_712,In_490);
nor U426 (N_426,In_279,In_690);
or U427 (N_427,In_1210,In_1038);
xor U428 (N_428,In_1436,In_460);
nor U429 (N_429,In_633,In_696);
and U430 (N_430,In_1130,In_33);
or U431 (N_431,In_1362,In_8);
xor U432 (N_432,In_1450,In_1033);
xor U433 (N_433,In_849,In_943);
nor U434 (N_434,In_180,In_899);
nor U435 (N_435,In_457,In_495);
xnor U436 (N_436,In_90,In_614);
or U437 (N_437,In_339,In_994);
nand U438 (N_438,In_167,In_561);
nand U439 (N_439,In_903,In_175);
and U440 (N_440,In_61,In_1029);
or U441 (N_441,In_108,In_1348);
nor U442 (N_442,In_440,In_565);
nor U443 (N_443,In_1430,In_226);
xor U444 (N_444,In_551,In_21);
or U445 (N_445,In_68,In_898);
and U446 (N_446,In_535,In_1415);
nand U447 (N_447,In_39,In_957);
nand U448 (N_448,In_1034,In_1452);
nor U449 (N_449,In_1058,In_699);
xnor U450 (N_450,In_231,In_579);
or U451 (N_451,In_908,In_1266);
nor U452 (N_452,In_388,In_1427);
and U453 (N_453,In_913,In_349);
nand U454 (N_454,In_1259,In_385);
and U455 (N_455,In_555,In_334);
and U456 (N_456,In_1439,In_966);
nand U457 (N_457,In_79,In_1272);
nor U458 (N_458,In_1290,In_1347);
or U459 (N_459,In_1197,In_918);
or U460 (N_460,In_1133,In_953);
and U461 (N_461,In_1478,In_754);
nor U462 (N_462,In_392,In_508);
and U463 (N_463,In_287,In_929);
nor U464 (N_464,In_1377,In_1032);
or U465 (N_465,In_550,In_732);
nand U466 (N_466,In_389,In_580);
and U467 (N_467,In_40,In_1373);
nor U468 (N_468,In_1056,In_794);
nor U469 (N_469,In_134,In_1459);
and U470 (N_470,In_247,In_1078);
or U471 (N_471,In_734,In_854);
or U472 (N_472,In_677,In_716);
or U473 (N_473,In_1276,In_997);
or U474 (N_474,In_1309,In_1438);
nand U475 (N_475,In_657,In_259);
or U476 (N_476,In_117,In_674);
nand U477 (N_477,In_573,In_1146);
and U478 (N_478,In_1227,In_1426);
or U479 (N_479,In_302,In_470);
nor U480 (N_480,In_1463,In_1144);
nand U481 (N_481,In_1188,In_1283);
nor U482 (N_482,In_577,In_1275);
nor U483 (N_483,In_1182,In_845);
nand U484 (N_484,In_1392,In_63);
or U485 (N_485,In_146,In_1132);
nand U486 (N_486,In_858,In_1424);
xnor U487 (N_487,In_1081,In_622);
nor U488 (N_488,In_1249,In_178);
or U489 (N_489,In_80,In_1370);
or U490 (N_490,In_1181,In_996);
xnor U491 (N_491,In_1050,In_954);
nor U492 (N_492,In_752,In_114);
nor U493 (N_493,In_297,In_761);
or U494 (N_494,In_711,In_749);
and U495 (N_495,In_821,In_1343);
and U496 (N_496,In_299,In_58);
or U497 (N_497,In_1135,In_151);
nand U498 (N_498,In_1320,In_1175);
nor U499 (N_499,In_1488,In_471);
and U500 (N_500,In_107,In_582);
xor U501 (N_501,In_416,In_1474);
nand U502 (N_502,In_1322,In_1310);
or U503 (N_503,In_767,In_515);
nor U504 (N_504,In_1358,In_1319);
nor U505 (N_505,In_413,In_1455);
xnor U506 (N_506,In_606,In_624);
xor U507 (N_507,In_1432,In_1074);
nand U508 (N_508,In_539,In_1252);
nand U509 (N_509,In_766,In_961);
nor U510 (N_510,In_200,In_1206);
nand U511 (N_511,In_343,In_368);
or U512 (N_512,In_394,In_452);
and U513 (N_513,In_189,In_1104);
nand U514 (N_514,In_322,In_808);
and U515 (N_515,In_1256,In_301);
nand U516 (N_516,In_763,In_1148);
and U517 (N_517,In_1293,In_290);
xor U518 (N_518,In_1317,In_916);
or U519 (N_519,In_1184,In_1469);
nor U520 (N_520,In_652,In_1324);
and U521 (N_521,In_765,In_197);
xnor U522 (N_522,In_1263,In_444);
and U523 (N_523,In_1225,In_617);
nor U524 (N_524,In_590,In_618);
or U525 (N_525,In_1429,In_469);
or U526 (N_526,In_35,In_429);
nand U527 (N_527,In_1131,In_116);
or U528 (N_528,In_668,In_16);
or U529 (N_529,In_1089,In_54);
nand U530 (N_530,In_1106,In_817);
or U531 (N_531,In_455,In_1349);
nand U532 (N_532,In_271,In_459);
xor U533 (N_533,In_827,In_989);
nand U534 (N_534,In_596,In_212);
and U535 (N_535,In_583,In_697);
nand U536 (N_536,In_848,In_157);
xor U537 (N_537,In_909,In_693);
and U538 (N_538,In_828,In_273);
nand U539 (N_539,In_882,In_974);
nand U540 (N_540,In_182,In_660);
and U541 (N_541,In_77,In_1454);
or U542 (N_542,In_451,In_1366);
and U543 (N_543,In_1313,In_613);
nor U544 (N_544,In_793,In_1281);
nand U545 (N_545,In_88,In_910);
or U546 (N_546,In_361,In_265);
or U547 (N_547,In_1153,In_637);
nor U548 (N_548,In_1291,In_210);
nand U549 (N_549,In_491,In_450);
or U550 (N_550,In_798,In_23);
nand U551 (N_551,In_230,In_639);
xor U552 (N_552,In_267,In_190);
and U553 (N_553,In_1397,In_1191);
or U554 (N_554,In_411,In_654);
and U555 (N_555,In_430,In_432);
nand U556 (N_556,In_1226,In_778);
nor U557 (N_557,In_1240,In_215);
nor U558 (N_558,In_876,In_375);
nand U559 (N_559,In_758,In_628);
nor U560 (N_560,In_775,In_307);
xnor U561 (N_561,In_48,In_81);
and U562 (N_562,In_906,In_529);
nor U563 (N_563,In_853,In_1234);
or U564 (N_564,In_1391,In_1064);
nor U565 (N_565,In_371,In_610);
nor U566 (N_566,In_1179,In_227);
nand U567 (N_567,In_236,In_527);
or U568 (N_568,In_530,In_484);
xnor U569 (N_569,In_1402,In_804);
or U570 (N_570,In_1384,In_1470);
nand U571 (N_571,In_648,In_826);
or U572 (N_572,In_1042,In_546);
nor U573 (N_573,In_664,In_97);
or U574 (N_574,In_274,In_1127);
and U575 (N_575,In_1251,In_1381);
and U576 (N_576,In_1371,In_372);
and U577 (N_577,In_790,In_517);
or U578 (N_578,In_816,In_857);
and U579 (N_579,In_360,In_45);
nand U580 (N_580,In_1399,In_621);
nand U581 (N_581,In_759,In_901);
nand U582 (N_582,In_9,In_1134);
and U583 (N_583,In_1110,In_1331);
nor U584 (N_584,In_1083,In_1174);
xor U585 (N_585,In_800,In_945);
or U586 (N_586,In_914,In_852);
nand U587 (N_587,In_783,In_159);
nor U588 (N_588,In_378,In_638);
or U589 (N_589,In_1113,In_1186);
nor U590 (N_590,In_563,In_229);
nand U591 (N_591,In_587,In_1268);
nand U592 (N_592,In_1115,In_559);
nor U593 (N_593,In_164,In_533);
nand U594 (N_594,In_49,In_1468);
or U595 (N_595,In_1284,In_1311);
nand U596 (N_596,In_497,In_1216);
nor U597 (N_597,In_1353,In_980);
xnor U598 (N_598,In_885,In_1097);
nor U599 (N_599,In_1142,In_195);
or U600 (N_600,In_139,In_1017);
nand U601 (N_601,In_553,In_1357);
nand U602 (N_602,In_511,In_401);
or U603 (N_603,In_1152,In_609);
or U604 (N_604,In_1103,In_1379);
and U605 (N_605,In_102,In_564);
and U606 (N_606,In_1192,In_931);
and U607 (N_607,In_1207,In_1222);
or U608 (N_608,In_883,In_1446);
and U609 (N_609,In_507,In_362);
nand U610 (N_610,In_585,In_43);
and U611 (N_611,In_1368,In_1414);
xnor U612 (N_612,In_220,In_1036);
nor U613 (N_613,In_950,In_1002);
and U614 (N_614,In_332,In_679);
nor U615 (N_615,In_1431,In_1315);
nor U616 (N_616,In_59,In_1423);
or U617 (N_617,In_1084,In_213);
nand U618 (N_618,In_1400,In_575);
xor U619 (N_619,In_478,In_120);
nor U620 (N_620,In_124,In_952);
nand U621 (N_621,In_629,In_666);
xor U622 (N_622,In_1211,In_109);
or U623 (N_623,In_836,In_1171);
or U624 (N_624,In_105,In_1297);
nand U625 (N_625,In_1088,In_1340);
nor U626 (N_626,In_475,In_55);
xor U627 (N_627,In_1326,In_890);
or U628 (N_628,In_304,In_85);
nand U629 (N_629,In_917,In_499);
nor U630 (N_630,In_1023,In_1338);
or U631 (N_631,In_1048,In_50);
or U632 (N_632,In_743,In_1408);
nand U633 (N_633,In_644,In_426);
nor U634 (N_634,In_143,In_839);
nand U635 (N_635,In_1025,In_15);
nand U636 (N_636,In_86,In_310);
xor U637 (N_637,In_412,In_541);
xnor U638 (N_638,In_1010,In_635);
or U639 (N_639,In_202,In_188);
or U640 (N_640,In_1062,In_1129);
nand U641 (N_641,In_65,In_795);
or U642 (N_642,In_1205,In_1378);
nor U643 (N_643,In_113,In_1246);
and U644 (N_644,In_1409,In_520);
and U645 (N_645,In_380,In_1383);
xor U646 (N_646,In_645,In_1049);
nand U647 (N_647,In_632,In_1434);
nor U648 (N_648,In_829,In_1218);
and U649 (N_649,In_1270,In_678);
and U650 (N_650,In_1200,In_548);
nor U651 (N_651,In_627,In_1108);
nand U652 (N_652,In_604,In_1410);
xnor U653 (N_653,In_60,In_340);
and U654 (N_654,In_281,In_991);
nand U655 (N_655,In_984,In_959);
and U656 (N_656,In_803,In_701);
nand U657 (N_657,In_671,In_651);
xnor U658 (N_658,In_843,In_1125);
or U659 (N_659,In_67,In_205);
and U660 (N_660,In_928,In_842);
nand U661 (N_661,In_661,In_1342);
or U662 (N_662,In_408,In_907);
nand U663 (N_663,In_319,In_435);
nand U664 (N_664,In_1096,In_1292);
and U665 (N_665,In_286,In_570);
or U666 (N_666,In_809,In_730);
xnor U667 (N_667,In_525,In_6);
nand U668 (N_668,In_1012,In_655);
nand U669 (N_669,In_488,In_1386);
or U670 (N_670,In_298,In_1262);
xor U671 (N_671,In_616,In_838);
or U672 (N_672,In_588,In_1289);
nor U673 (N_673,In_132,In_894);
nor U674 (N_674,In_718,In_1138);
xor U675 (N_675,In_726,In_168);
nor U676 (N_676,In_1046,In_1163);
or U677 (N_677,In_467,In_198);
and U678 (N_678,In_572,In_1288);
nor U679 (N_679,In_154,In_872);
nor U680 (N_680,In_7,In_369);
or U681 (N_681,In_505,In_1258);
nor U682 (N_682,In_156,In_405);
nor U683 (N_683,In_1044,In_1330);
and U684 (N_684,In_1114,In_1143);
nand U685 (N_685,In_1334,In_774);
nor U686 (N_686,In_1327,In_706);
and U687 (N_687,In_466,In_1220);
and U688 (N_688,In_1212,In_598);
nand U689 (N_689,In_422,In_468);
nand U690 (N_690,In_1093,In_1239);
nand U691 (N_691,In_1102,In_1367);
nand U692 (N_692,In_1090,In_830);
nor U693 (N_693,In_675,In_847);
nor U694 (N_694,In_1301,In_921);
xnor U695 (N_695,In_881,In_275);
and U696 (N_696,In_1303,In_1203);
nand U697 (N_697,In_374,In_476);
and U698 (N_698,In_1360,In_740);
nor U699 (N_699,In_10,In_305);
nor U700 (N_700,In_904,In_599);
or U701 (N_701,In_324,In_626);
nor U702 (N_702,In_1183,In_1498);
or U703 (N_703,In_261,In_1464);
or U704 (N_704,In_949,In_1121);
or U705 (N_705,In_1014,In_877);
nand U706 (N_706,In_1217,In_1298);
or U707 (N_707,In_489,In_171);
xnor U708 (N_708,In_1458,In_823);
nor U709 (N_709,In_1052,In_255);
or U710 (N_710,In_1411,In_318);
nand U711 (N_711,In_47,In_1440);
nand U712 (N_712,In_141,In_248);
xor U713 (N_713,In_506,In_354);
and U714 (N_714,In_971,In_955);
nand U715 (N_715,In_545,In_1394);
and U716 (N_716,In_1265,In_976);
or U717 (N_717,In_688,In_1321);
nor U718 (N_718,In_879,In_776);
or U719 (N_719,In_544,In_37);
or U720 (N_720,In_346,In_500);
or U721 (N_721,In_746,In_355);
nor U722 (N_722,In_1055,In_574);
nand U723 (N_723,In_1279,In_1201);
nand U724 (N_724,In_351,In_366);
and U725 (N_725,In_1085,In_266);
or U726 (N_726,In_1019,In_524);
or U727 (N_727,In_1079,In_722);
or U728 (N_728,In_194,In_323);
nor U729 (N_729,In_895,In_719);
nor U730 (N_730,In_1274,In_738);
and U731 (N_731,In_177,In_1160);
xnor U732 (N_732,In_600,In_257);
nor U733 (N_733,In_149,In_1425);
nor U734 (N_734,In_751,In_773);
nor U735 (N_735,In_1480,In_439);
nor U736 (N_736,In_1028,In_98);
nor U737 (N_737,In_278,In_1107);
nor U738 (N_738,In_1167,In_731);
xnor U739 (N_739,In_1441,In_436);
nand U740 (N_740,In_640,In_1151);
and U741 (N_741,In_216,In_295);
nor U742 (N_742,In_1442,In_762);
xor U743 (N_743,In_704,In_280);
or U744 (N_744,In_1495,In_1007);
nor U745 (N_745,In_653,In_121);
nand U746 (N_746,In_1261,In_367);
nor U747 (N_747,In_571,In_17);
or U748 (N_748,In_990,In_1111);
and U749 (N_749,In_122,In_464);
or U750 (N_750,In_1369,In_1170);
nand U751 (N_751,In_811,In_566);
nor U752 (N_752,In_291,In_1006);
nor U753 (N_753,In_312,In_165);
and U754 (N_754,In_679,In_506);
xor U755 (N_755,In_411,In_243);
nor U756 (N_756,In_318,In_563);
and U757 (N_757,In_395,In_107);
xnor U758 (N_758,In_1192,In_668);
nand U759 (N_759,In_1293,In_529);
xor U760 (N_760,In_1410,In_1470);
and U761 (N_761,In_1130,In_1270);
xor U762 (N_762,In_817,In_276);
nand U763 (N_763,In_1028,In_239);
nand U764 (N_764,In_1284,In_234);
or U765 (N_765,In_1190,In_964);
nor U766 (N_766,In_117,In_1224);
and U767 (N_767,In_1309,In_449);
or U768 (N_768,In_960,In_903);
or U769 (N_769,In_195,In_470);
nand U770 (N_770,In_17,In_128);
nor U771 (N_771,In_346,In_1275);
or U772 (N_772,In_747,In_46);
nand U773 (N_773,In_1009,In_805);
nor U774 (N_774,In_157,In_533);
and U775 (N_775,In_1408,In_541);
nand U776 (N_776,In_74,In_1024);
xor U777 (N_777,In_758,In_1047);
and U778 (N_778,In_1288,In_1290);
nand U779 (N_779,In_473,In_1249);
and U780 (N_780,In_416,In_1157);
and U781 (N_781,In_57,In_1411);
nand U782 (N_782,In_1,In_985);
and U783 (N_783,In_231,In_597);
and U784 (N_784,In_1110,In_1140);
xor U785 (N_785,In_785,In_1174);
or U786 (N_786,In_1435,In_1446);
or U787 (N_787,In_1229,In_221);
nand U788 (N_788,In_1093,In_893);
nand U789 (N_789,In_279,In_541);
or U790 (N_790,In_723,In_150);
nor U791 (N_791,In_491,In_1353);
and U792 (N_792,In_153,In_668);
and U793 (N_793,In_486,In_920);
xnor U794 (N_794,In_1341,In_259);
or U795 (N_795,In_286,In_467);
nor U796 (N_796,In_207,In_886);
or U797 (N_797,In_1478,In_1472);
nand U798 (N_798,In_750,In_414);
or U799 (N_799,In_448,In_1303);
nand U800 (N_800,In_732,In_1053);
nor U801 (N_801,In_1056,In_1349);
or U802 (N_802,In_720,In_1289);
nand U803 (N_803,In_1298,In_1211);
nor U804 (N_804,In_589,In_985);
and U805 (N_805,In_214,In_366);
xor U806 (N_806,In_216,In_474);
nand U807 (N_807,In_595,In_1308);
nand U808 (N_808,In_1095,In_547);
nor U809 (N_809,In_163,In_101);
nand U810 (N_810,In_1362,In_1364);
or U811 (N_811,In_653,In_779);
and U812 (N_812,In_109,In_846);
or U813 (N_813,In_716,In_1255);
nor U814 (N_814,In_543,In_273);
or U815 (N_815,In_781,In_542);
nand U816 (N_816,In_2,In_479);
or U817 (N_817,In_308,In_167);
nor U818 (N_818,In_613,In_679);
nor U819 (N_819,In_1366,In_352);
and U820 (N_820,In_1346,In_318);
nand U821 (N_821,In_401,In_944);
xnor U822 (N_822,In_1105,In_1162);
or U823 (N_823,In_596,In_1245);
and U824 (N_824,In_549,In_595);
nor U825 (N_825,In_910,In_613);
nor U826 (N_826,In_258,In_1032);
nand U827 (N_827,In_742,In_1351);
nand U828 (N_828,In_304,In_1371);
and U829 (N_829,In_164,In_238);
nand U830 (N_830,In_852,In_1310);
nand U831 (N_831,In_1217,In_1337);
or U832 (N_832,In_1312,In_972);
nor U833 (N_833,In_488,In_1302);
nand U834 (N_834,In_47,In_1253);
nor U835 (N_835,In_1145,In_1304);
nand U836 (N_836,In_345,In_772);
nand U837 (N_837,In_878,In_1206);
nand U838 (N_838,In_112,In_1493);
or U839 (N_839,In_1355,In_950);
xor U840 (N_840,In_1039,In_1220);
and U841 (N_841,In_229,In_848);
or U842 (N_842,In_639,In_1315);
nor U843 (N_843,In_546,In_1145);
and U844 (N_844,In_700,In_371);
nand U845 (N_845,In_1499,In_1157);
and U846 (N_846,In_887,In_403);
or U847 (N_847,In_1181,In_549);
nor U848 (N_848,In_1254,In_1466);
or U849 (N_849,In_735,In_684);
xnor U850 (N_850,In_1041,In_454);
nor U851 (N_851,In_215,In_467);
or U852 (N_852,In_417,In_1236);
and U853 (N_853,In_562,In_743);
and U854 (N_854,In_1465,In_1294);
and U855 (N_855,In_412,In_31);
nor U856 (N_856,In_630,In_742);
and U857 (N_857,In_265,In_1096);
nor U858 (N_858,In_1140,In_344);
and U859 (N_859,In_799,In_465);
and U860 (N_860,In_308,In_1275);
nand U861 (N_861,In_739,In_6);
and U862 (N_862,In_1107,In_62);
or U863 (N_863,In_220,In_939);
xnor U864 (N_864,In_368,In_170);
nand U865 (N_865,In_866,In_1111);
xnor U866 (N_866,In_74,In_272);
or U867 (N_867,In_424,In_978);
or U868 (N_868,In_90,In_191);
nand U869 (N_869,In_508,In_714);
nand U870 (N_870,In_811,In_224);
or U871 (N_871,In_1093,In_673);
nor U872 (N_872,In_715,In_997);
and U873 (N_873,In_1058,In_875);
nand U874 (N_874,In_684,In_781);
nand U875 (N_875,In_859,In_328);
nand U876 (N_876,In_823,In_593);
nand U877 (N_877,In_678,In_1050);
and U878 (N_878,In_1213,In_629);
or U879 (N_879,In_866,In_503);
xor U880 (N_880,In_1126,In_588);
nor U881 (N_881,In_1294,In_904);
or U882 (N_882,In_743,In_246);
or U883 (N_883,In_568,In_156);
and U884 (N_884,In_741,In_45);
nand U885 (N_885,In_360,In_822);
or U886 (N_886,In_553,In_193);
and U887 (N_887,In_588,In_1495);
or U888 (N_888,In_299,In_439);
or U889 (N_889,In_787,In_499);
nand U890 (N_890,In_522,In_1422);
or U891 (N_891,In_527,In_1008);
nor U892 (N_892,In_23,In_369);
and U893 (N_893,In_739,In_764);
or U894 (N_894,In_824,In_1322);
nor U895 (N_895,In_1178,In_1248);
and U896 (N_896,In_153,In_714);
nand U897 (N_897,In_656,In_428);
or U898 (N_898,In_532,In_563);
nand U899 (N_899,In_1480,In_526);
xnor U900 (N_900,In_1117,In_613);
nor U901 (N_901,In_289,In_1492);
and U902 (N_902,In_326,In_1398);
xnor U903 (N_903,In_1033,In_320);
or U904 (N_904,In_99,In_456);
or U905 (N_905,In_518,In_957);
and U906 (N_906,In_261,In_1108);
and U907 (N_907,In_421,In_582);
or U908 (N_908,In_1209,In_73);
nand U909 (N_909,In_961,In_1292);
nand U910 (N_910,In_464,In_1478);
or U911 (N_911,In_61,In_525);
or U912 (N_912,In_1310,In_587);
nor U913 (N_913,In_459,In_1344);
nor U914 (N_914,In_1055,In_153);
nor U915 (N_915,In_151,In_353);
or U916 (N_916,In_731,In_1277);
nand U917 (N_917,In_1423,In_1230);
and U918 (N_918,In_21,In_412);
nand U919 (N_919,In_1082,In_1270);
nand U920 (N_920,In_1054,In_360);
nand U921 (N_921,In_1360,In_370);
or U922 (N_922,In_1331,In_435);
or U923 (N_923,In_1038,In_1129);
nor U924 (N_924,In_297,In_727);
and U925 (N_925,In_1479,In_1170);
nand U926 (N_926,In_856,In_1209);
nand U927 (N_927,In_1438,In_1077);
nor U928 (N_928,In_553,In_1232);
or U929 (N_929,In_352,In_1307);
xor U930 (N_930,In_683,In_728);
nor U931 (N_931,In_558,In_727);
or U932 (N_932,In_514,In_474);
or U933 (N_933,In_545,In_1328);
or U934 (N_934,In_1448,In_1368);
and U935 (N_935,In_156,In_1392);
or U936 (N_936,In_658,In_42);
or U937 (N_937,In_1030,In_1069);
nand U938 (N_938,In_576,In_115);
nand U939 (N_939,In_636,In_560);
nor U940 (N_940,In_200,In_299);
nand U941 (N_941,In_1492,In_1440);
xor U942 (N_942,In_1088,In_874);
nand U943 (N_943,In_1388,In_103);
or U944 (N_944,In_898,In_361);
nor U945 (N_945,In_673,In_1171);
nor U946 (N_946,In_817,In_629);
and U947 (N_947,In_102,In_1329);
nand U948 (N_948,In_1178,In_90);
and U949 (N_949,In_1362,In_350);
and U950 (N_950,In_1383,In_659);
nand U951 (N_951,In_127,In_466);
nand U952 (N_952,In_495,In_534);
nand U953 (N_953,In_45,In_818);
or U954 (N_954,In_1290,In_747);
nand U955 (N_955,In_964,In_915);
nand U956 (N_956,In_273,In_780);
nand U957 (N_957,In_1053,In_1274);
or U958 (N_958,In_1013,In_136);
or U959 (N_959,In_525,In_1010);
or U960 (N_960,In_1099,In_1189);
and U961 (N_961,In_1123,In_159);
or U962 (N_962,In_432,In_100);
or U963 (N_963,In_1497,In_757);
nor U964 (N_964,In_1118,In_606);
nor U965 (N_965,In_896,In_957);
or U966 (N_966,In_556,In_500);
nor U967 (N_967,In_835,In_704);
xor U968 (N_968,In_482,In_1108);
and U969 (N_969,In_919,In_1126);
or U970 (N_970,In_661,In_1121);
nor U971 (N_971,In_1224,In_1338);
nor U972 (N_972,In_1041,In_395);
and U973 (N_973,In_1476,In_786);
or U974 (N_974,In_525,In_1091);
or U975 (N_975,In_1407,In_844);
or U976 (N_976,In_1414,In_792);
nand U977 (N_977,In_571,In_1280);
nor U978 (N_978,In_1342,In_657);
nand U979 (N_979,In_1120,In_467);
nor U980 (N_980,In_1445,In_314);
or U981 (N_981,In_494,In_715);
nand U982 (N_982,In_852,In_451);
or U983 (N_983,In_1087,In_802);
nor U984 (N_984,In_940,In_668);
xor U985 (N_985,In_1037,In_1440);
and U986 (N_986,In_1118,In_796);
nand U987 (N_987,In_73,In_1497);
or U988 (N_988,In_1411,In_758);
or U989 (N_989,In_696,In_62);
nor U990 (N_990,In_246,In_713);
nor U991 (N_991,In_417,In_387);
and U992 (N_992,In_1490,In_76);
nand U993 (N_993,In_884,In_699);
nor U994 (N_994,In_476,In_35);
and U995 (N_995,In_842,In_542);
nand U996 (N_996,In_770,In_327);
nor U997 (N_997,In_13,In_1112);
and U998 (N_998,In_966,In_771);
or U999 (N_999,In_840,In_1347);
nor U1000 (N_1000,In_450,In_966);
and U1001 (N_1001,In_598,In_673);
and U1002 (N_1002,In_1048,In_408);
xnor U1003 (N_1003,In_675,In_55);
nor U1004 (N_1004,In_357,In_335);
or U1005 (N_1005,In_931,In_440);
xor U1006 (N_1006,In_309,In_506);
nor U1007 (N_1007,In_357,In_1139);
and U1008 (N_1008,In_128,In_1054);
or U1009 (N_1009,In_253,In_1473);
nand U1010 (N_1010,In_794,In_876);
nor U1011 (N_1011,In_590,In_1273);
nand U1012 (N_1012,In_869,In_565);
xor U1013 (N_1013,In_1113,In_178);
nand U1014 (N_1014,In_709,In_1438);
nor U1015 (N_1015,In_1489,In_99);
or U1016 (N_1016,In_1411,In_252);
nand U1017 (N_1017,In_504,In_1409);
nand U1018 (N_1018,In_1122,In_1019);
or U1019 (N_1019,In_1103,In_15);
nand U1020 (N_1020,In_431,In_1391);
and U1021 (N_1021,In_356,In_862);
or U1022 (N_1022,In_135,In_528);
and U1023 (N_1023,In_500,In_83);
and U1024 (N_1024,In_697,In_490);
nor U1025 (N_1025,In_1415,In_663);
and U1026 (N_1026,In_1049,In_1469);
nor U1027 (N_1027,In_1427,In_1086);
and U1028 (N_1028,In_1412,In_1079);
nand U1029 (N_1029,In_331,In_670);
and U1030 (N_1030,In_716,In_633);
nor U1031 (N_1031,In_1226,In_1411);
or U1032 (N_1032,In_1446,In_471);
and U1033 (N_1033,In_1079,In_696);
nor U1034 (N_1034,In_156,In_940);
nor U1035 (N_1035,In_824,In_569);
nand U1036 (N_1036,In_701,In_41);
nor U1037 (N_1037,In_1325,In_1330);
nand U1038 (N_1038,In_577,In_1179);
xor U1039 (N_1039,In_660,In_96);
or U1040 (N_1040,In_1281,In_929);
or U1041 (N_1041,In_588,In_254);
and U1042 (N_1042,In_1455,In_861);
nand U1043 (N_1043,In_365,In_1194);
and U1044 (N_1044,In_529,In_1348);
or U1045 (N_1045,In_1282,In_1164);
nand U1046 (N_1046,In_266,In_1077);
nand U1047 (N_1047,In_982,In_15);
or U1048 (N_1048,In_460,In_32);
nor U1049 (N_1049,In_473,In_591);
nand U1050 (N_1050,In_389,In_221);
or U1051 (N_1051,In_9,In_1332);
nand U1052 (N_1052,In_1169,In_918);
nand U1053 (N_1053,In_338,In_766);
and U1054 (N_1054,In_525,In_499);
nand U1055 (N_1055,In_386,In_892);
and U1056 (N_1056,In_680,In_1310);
nand U1057 (N_1057,In_793,In_88);
nand U1058 (N_1058,In_270,In_1283);
and U1059 (N_1059,In_271,In_580);
nand U1060 (N_1060,In_406,In_86);
and U1061 (N_1061,In_777,In_461);
nand U1062 (N_1062,In_1222,In_1271);
nor U1063 (N_1063,In_398,In_1228);
nand U1064 (N_1064,In_735,In_1298);
nor U1065 (N_1065,In_594,In_259);
nand U1066 (N_1066,In_120,In_1299);
nor U1067 (N_1067,In_1134,In_339);
and U1068 (N_1068,In_1103,In_941);
xor U1069 (N_1069,In_282,In_199);
xnor U1070 (N_1070,In_927,In_171);
nand U1071 (N_1071,In_1025,In_689);
xor U1072 (N_1072,In_331,In_1178);
nand U1073 (N_1073,In_223,In_3);
nor U1074 (N_1074,In_719,In_633);
or U1075 (N_1075,In_624,In_1229);
and U1076 (N_1076,In_38,In_265);
and U1077 (N_1077,In_958,In_755);
or U1078 (N_1078,In_979,In_1390);
nor U1079 (N_1079,In_259,In_488);
and U1080 (N_1080,In_1170,In_1097);
and U1081 (N_1081,In_284,In_1326);
or U1082 (N_1082,In_41,In_1067);
and U1083 (N_1083,In_376,In_209);
or U1084 (N_1084,In_615,In_858);
and U1085 (N_1085,In_4,In_990);
nand U1086 (N_1086,In_1141,In_384);
or U1087 (N_1087,In_687,In_578);
or U1088 (N_1088,In_1384,In_480);
nand U1089 (N_1089,In_620,In_467);
or U1090 (N_1090,In_1441,In_938);
nor U1091 (N_1091,In_1487,In_859);
xor U1092 (N_1092,In_570,In_113);
nor U1093 (N_1093,In_574,In_1371);
and U1094 (N_1094,In_1289,In_793);
or U1095 (N_1095,In_1237,In_1498);
and U1096 (N_1096,In_692,In_742);
or U1097 (N_1097,In_394,In_1261);
nand U1098 (N_1098,In_32,In_774);
nor U1099 (N_1099,In_997,In_862);
or U1100 (N_1100,In_346,In_778);
and U1101 (N_1101,In_1368,In_883);
nor U1102 (N_1102,In_756,In_261);
and U1103 (N_1103,In_640,In_1287);
and U1104 (N_1104,In_980,In_15);
or U1105 (N_1105,In_674,In_1112);
or U1106 (N_1106,In_37,In_1130);
or U1107 (N_1107,In_1095,In_49);
and U1108 (N_1108,In_731,In_168);
and U1109 (N_1109,In_337,In_1076);
nand U1110 (N_1110,In_1197,In_187);
xnor U1111 (N_1111,In_281,In_1498);
xor U1112 (N_1112,In_416,In_1461);
nor U1113 (N_1113,In_1042,In_1013);
and U1114 (N_1114,In_716,In_1137);
nand U1115 (N_1115,In_1496,In_813);
or U1116 (N_1116,In_904,In_862);
nor U1117 (N_1117,In_593,In_306);
nand U1118 (N_1118,In_819,In_98);
nand U1119 (N_1119,In_1356,In_865);
nand U1120 (N_1120,In_1199,In_323);
nor U1121 (N_1121,In_1105,In_1341);
nand U1122 (N_1122,In_1314,In_44);
and U1123 (N_1123,In_403,In_448);
and U1124 (N_1124,In_599,In_381);
or U1125 (N_1125,In_1471,In_239);
nor U1126 (N_1126,In_1475,In_594);
xnor U1127 (N_1127,In_1486,In_111);
or U1128 (N_1128,In_1370,In_182);
or U1129 (N_1129,In_37,In_1469);
and U1130 (N_1130,In_462,In_705);
nor U1131 (N_1131,In_956,In_1460);
nand U1132 (N_1132,In_597,In_1427);
nor U1133 (N_1133,In_1409,In_1201);
and U1134 (N_1134,In_1378,In_255);
or U1135 (N_1135,In_853,In_1115);
nor U1136 (N_1136,In_857,In_1312);
nand U1137 (N_1137,In_410,In_1437);
nor U1138 (N_1138,In_508,In_1444);
or U1139 (N_1139,In_544,In_911);
and U1140 (N_1140,In_778,In_967);
and U1141 (N_1141,In_219,In_711);
and U1142 (N_1142,In_350,In_1119);
nor U1143 (N_1143,In_285,In_1398);
nand U1144 (N_1144,In_459,In_1439);
and U1145 (N_1145,In_372,In_1097);
or U1146 (N_1146,In_461,In_1343);
nand U1147 (N_1147,In_1116,In_494);
nand U1148 (N_1148,In_478,In_90);
nand U1149 (N_1149,In_466,In_1355);
and U1150 (N_1150,In_45,In_428);
or U1151 (N_1151,In_1034,In_562);
nor U1152 (N_1152,In_221,In_394);
and U1153 (N_1153,In_476,In_993);
and U1154 (N_1154,In_1265,In_402);
nor U1155 (N_1155,In_313,In_594);
xor U1156 (N_1156,In_475,In_19);
nand U1157 (N_1157,In_348,In_1270);
and U1158 (N_1158,In_997,In_310);
and U1159 (N_1159,In_362,In_1204);
or U1160 (N_1160,In_525,In_1221);
xor U1161 (N_1161,In_1076,In_1048);
or U1162 (N_1162,In_938,In_574);
or U1163 (N_1163,In_756,In_383);
and U1164 (N_1164,In_1453,In_1045);
and U1165 (N_1165,In_1473,In_883);
or U1166 (N_1166,In_1104,In_137);
and U1167 (N_1167,In_944,In_365);
nand U1168 (N_1168,In_454,In_1061);
or U1169 (N_1169,In_975,In_1207);
xor U1170 (N_1170,In_1261,In_1099);
or U1171 (N_1171,In_951,In_891);
and U1172 (N_1172,In_1127,In_619);
or U1173 (N_1173,In_633,In_91);
xnor U1174 (N_1174,In_143,In_419);
nand U1175 (N_1175,In_734,In_1221);
nor U1176 (N_1176,In_1200,In_998);
or U1177 (N_1177,In_58,In_1220);
or U1178 (N_1178,In_1346,In_1350);
or U1179 (N_1179,In_1193,In_631);
or U1180 (N_1180,In_363,In_247);
nand U1181 (N_1181,In_324,In_1346);
nand U1182 (N_1182,In_482,In_500);
and U1183 (N_1183,In_301,In_374);
nand U1184 (N_1184,In_510,In_950);
xnor U1185 (N_1185,In_576,In_715);
or U1186 (N_1186,In_1386,In_922);
or U1187 (N_1187,In_291,In_1087);
nand U1188 (N_1188,In_1310,In_443);
and U1189 (N_1189,In_1414,In_1381);
nand U1190 (N_1190,In_67,In_105);
or U1191 (N_1191,In_930,In_1050);
nor U1192 (N_1192,In_979,In_346);
or U1193 (N_1193,In_109,In_204);
xnor U1194 (N_1194,In_1338,In_697);
and U1195 (N_1195,In_554,In_1137);
nor U1196 (N_1196,In_1138,In_139);
nor U1197 (N_1197,In_997,In_1437);
or U1198 (N_1198,In_549,In_905);
xnor U1199 (N_1199,In_1044,In_552);
or U1200 (N_1200,In_122,In_1359);
or U1201 (N_1201,In_1133,In_687);
and U1202 (N_1202,In_1046,In_1274);
nand U1203 (N_1203,In_149,In_557);
nand U1204 (N_1204,In_944,In_632);
or U1205 (N_1205,In_362,In_503);
nand U1206 (N_1206,In_489,In_1369);
nor U1207 (N_1207,In_1365,In_986);
or U1208 (N_1208,In_857,In_1408);
nor U1209 (N_1209,In_573,In_1472);
nand U1210 (N_1210,In_933,In_1065);
nand U1211 (N_1211,In_286,In_823);
or U1212 (N_1212,In_160,In_129);
nor U1213 (N_1213,In_1459,In_1372);
and U1214 (N_1214,In_1277,In_909);
nand U1215 (N_1215,In_406,In_541);
and U1216 (N_1216,In_688,In_1458);
nor U1217 (N_1217,In_677,In_506);
xor U1218 (N_1218,In_65,In_1405);
nand U1219 (N_1219,In_777,In_1284);
nand U1220 (N_1220,In_14,In_1394);
and U1221 (N_1221,In_1309,In_1258);
and U1222 (N_1222,In_1334,In_374);
nor U1223 (N_1223,In_635,In_853);
nor U1224 (N_1224,In_53,In_1278);
nor U1225 (N_1225,In_1183,In_679);
xnor U1226 (N_1226,In_845,In_722);
nand U1227 (N_1227,In_934,In_65);
xor U1228 (N_1228,In_76,In_603);
and U1229 (N_1229,In_774,In_148);
or U1230 (N_1230,In_265,In_927);
nor U1231 (N_1231,In_139,In_697);
and U1232 (N_1232,In_256,In_889);
nor U1233 (N_1233,In_603,In_554);
nor U1234 (N_1234,In_1150,In_1425);
nand U1235 (N_1235,In_1081,In_111);
and U1236 (N_1236,In_467,In_1032);
and U1237 (N_1237,In_1449,In_385);
nor U1238 (N_1238,In_766,In_1156);
or U1239 (N_1239,In_982,In_480);
nand U1240 (N_1240,In_128,In_1305);
nand U1241 (N_1241,In_663,In_1116);
nand U1242 (N_1242,In_1089,In_1440);
nand U1243 (N_1243,In_1497,In_1205);
and U1244 (N_1244,In_1451,In_103);
nor U1245 (N_1245,In_837,In_1174);
nor U1246 (N_1246,In_117,In_350);
and U1247 (N_1247,In_1209,In_1396);
or U1248 (N_1248,In_1251,In_539);
and U1249 (N_1249,In_1459,In_192);
or U1250 (N_1250,In_206,In_617);
nor U1251 (N_1251,In_992,In_1088);
nand U1252 (N_1252,In_902,In_665);
or U1253 (N_1253,In_152,In_826);
or U1254 (N_1254,In_490,In_654);
nand U1255 (N_1255,In_499,In_163);
nor U1256 (N_1256,In_587,In_735);
nand U1257 (N_1257,In_1166,In_596);
nand U1258 (N_1258,In_719,In_19);
nor U1259 (N_1259,In_1153,In_462);
or U1260 (N_1260,In_993,In_594);
nand U1261 (N_1261,In_420,In_1161);
nand U1262 (N_1262,In_1488,In_81);
or U1263 (N_1263,In_671,In_1332);
nand U1264 (N_1264,In_374,In_358);
nand U1265 (N_1265,In_389,In_428);
nor U1266 (N_1266,In_1168,In_599);
and U1267 (N_1267,In_187,In_1328);
and U1268 (N_1268,In_1495,In_446);
and U1269 (N_1269,In_690,In_165);
xor U1270 (N_1270,In_480,In_977);
and U1271 (N_1271,In_1420,In_1425);
nand U1272 (N_1272,In_1489,In_562);
or U1273 (N_1273,In_194,In_247);
nand U1274 (N_1274,In_312,In_1107);
or U1275 (N_1275,In_627,In_157);
and U1276 (N_1276,In_1227,In_139);
nor U1277 (N_1277,In_302,In_136);
nor U1278 (N_1278,In_116,In_252);
xnor U1279 (N_1279,In_961,In_839);
and U1280 (N_1280,In_1237,In_37);
and U1281 (N_1281,In_425,In_1093);
and U1282 (N_1282,In_1338,In_1034);
nand U1283 (N_1283,In_1186,In_1020);
nand U1284 (N_1284,In_1349,In_765);
or U1285 (N_1285,In_1190,In_1391);
and U1286 (N_1286,In_344,In_106);
or U1287 (N_1287,In_334,In_789);
and U1288 (N_1288,In_592,In_850);
and U1289 (N_1289,In_1373,In_419);
xnor U1290 (N_1290,In_740,In_12);
nor U1291 (N_1291,In_762,In_177);
or U1292 (N_1292,In_223,In_535);
nand U1293 (N_1293,In_808,In_661);
nand U1294 (N_1294,In_1276,In_1282);
and U1295 (N_1295,In_824,In_1341);
nand U1296 (N_1296,In_882,In_1128);
and U1297 (N_1297,In_1076,In_737);
or U1298 (N_1298,In_533,In_713);
or U1299 (N_1299,In_258,In_503);
nor U1300 (N_1300,In_1255,In_1364);
and U1301 (N_1301,In_1481,In_1178);
xnor U1302 (N_1302,In_825,In_74);
nor U1303 (N_1303,In_1073,In_1403);
or U1304 (N_1304,In_929,In_1456);
nand U1305 (N_1305,In_64,In_663);
or U1306 (N_1306,In_197,In_1437);
nand U1307 (N_1307,In_568,In_1017);
nand U1308 (N_1308,In_1274,In_0);
or U1309 (N_1309,In_462,In_1430);
and U1310 (N_1310,In_1055,In_888);
and U1311 (N_1311,In_258,In_31);
nor U1312 (N_1312,In_102,In_559);
nand U1313 (N_1313,In_324,In_364);
nor U1314 (N_1314,In_935,In_878);
and U1315 (N_1315,In_1457,In_1018);
nor U1316 (N_1316,In_1243,In_1146);
nand U1317 (N_1317,In_1081,In_219);
nand U1318 (N_1318,In_1127,In_889);
nand U1319 (N_1319,In_1422,In_1472);
and U1320 (N_1320,In_725,In_290);
or U1321 (N_1321,In_351,In_1109);
nor U1322 (N_1322,In_908,In_572);
or U1323 (N_1323,In_1143,In_1352);
xnor U1324 (N_1324,In_711,In_163);
nor U1325 (N_1325,In_959,In_14);
nor U1326 (N_1326,In_777,In_586);
nand U1327 (N_1327,In_676,In_1264);
or U1328 (N_1328,In_483,In_1174);
and U1329 (N_1329,In_901,In_771);
nand U1330 (N_1330,In_952,In_1446);
nor U1331 (N_1331,In_929,In_523);
and U1332 (N_1332,In_987,In_815);
and U1333 (N_1333,In_996,In_865);
nor U1334 (N_1334,In_1219,In_1304);
nor U1335 (N_1335,In_936,In_64);
or U1336 (N_1336,In_1305,In_1387);
or U1337 (N_1337,In_93,In_391);
nand U1338 (N_1338,In_166,In_1175);
nand U1339 (N_1339,In_1225,In_1110);
nor U1340 (N_1340,In_1266,In_1126);
nand U1341 (N_1341,In_1131,In_142);
xnor U1342 (N_1342,In_1000,In_148);
nor U1343 (N_1343,In_930,In_1022);
nor U1344 (N_1344,In_995,In_1051);
and U1345 (N_1345,In_1360,In_718);
nand U1346 (N_1346,In_1242,In_467);
nand U1347 (N_1347,In_1074,In_158);
and U1348 (N_1348,In_110,In_684);
or U1349 (N_1349,In_264,In_900);
and U1350 (N_1350,In_1161,In_9);
or U1351 (N_1351,In_668,In_319);
and U1352 (N_1352,In_442,In_599);
xnor U1353 (N_1353,In_1319,In_651);
nand U1354 (N_1354,In_530,In_437);
or U1355 (N_1355,In_1290,In_1469);
nor U1356 (N_1356,In_508,In_898);
xnor U1357 (N_1357,In_827,In_115);
nand U1358 (N_1358,In_397,In_146);
or U1359 (N_1359,In_78,In_689);
nor U1360 (N_1360,In_388,In_1467);
xnor U1361 (N_1361,In_1337,In_1046);
nand U1362 (N_1362,In_844,In_537);
and U1363 (N_1363,In_815,In_416);
or U1364 (N_1364,In_798,In_35);
xnor U1365 (N_1365,In_491,In_323);
nor U1366 (N_1366,In_1429,In_258);
nor U1367 (N_1367,In_242,In_1364);
and U1368 (N_1368,In_659,In_1345);
or U1369 (N_1369,In_258,In_254);
or U1370 (N_1370,In_1403,In_274);
and U1371 (N_1371,In_252,In_1312);
nand U1372 (N_1372,In_1066,In_228);
nor U1373 (N_1373,In_1362,In_1045);
and U1374 (N_1374,In_482,In_1464);
nor U1375 (N_1375,In_256,In_164);
nor U1376 (N_1376,In_498,In_588);
nand U1377 (N_1377,In_541,In_1222);
nand U1378 (N_1378,In_861,In_442);
or U1379 (N_1379,In_311,In_710);
nor U1380 (N_1380,In_957,In_1318);
or U1381 (N_1381,In_136,In_489);
nor U1382 (N_1382,In_722,In_680);
or U1383 (N_1383,In_433,In_1184);
and U1384 (N_1384,In_653,In_31);
nand U1385 (N_1385,In_510,In_1165);
nor U1386 (N_1386,In_1136,In_307);
nor U1387 (N_1387,In_705,In_963);
or U1388 (N_1388,In_378,In_1410);
and U1389 (N_1389,In_1439,In_1191);
xnor U1390 (N_1390,In_1416,In_1390);
nand U1391 (N_1391,In_1319,In_988);
nor U1392 (N_1392,In_1338,In_667);
and U1393 (N_1393,In_946,In_1251);
nand U1394 (N_1394,In_728,In_1296);
or U1395 (N_1395,In_168,In_1140);
nor U1396 (N_1396,In_661,In_618);
xor U1397 (N_1397,In_463,In_1476);
nand U1398 (N_1398,In_158,In_483);
and U1399 (N_1399,In_495,In_378);
nor U1400 (N_1400,In_70,In_960);
or U1401 (N_1401,In_983,In_159);
nor U1402 (N_1402,In_703,In_646);
and U1403 (N_1403,In_1324,In_558);
and U1404 (N_1404,In_284,In_1377);
and U1405 (N_1405,In_759,In_1002);
or U1406 (N_1406,In_591,In_21);
or U1407 (N_1407,In_626,In_636);
and U1408 (N_1408,In_210,In_1343);
or U1409 (N_1409,In_972,In_437);
xor U1410 (N_1410,In_931,In_589);
nor U1411 (N_1411,In_1398,In_150);
and U1412 (N_1412,In_1285,In_630);
nand U1413 (N_1413,In_1039,In_729);
nor U1414 (N_1414,In_1452,In_823);
nand U1415 (N_1415,In_145,In_377);
nor U1416 (N_1416,In_1323,In_1069);
and U1417 (N_1417,In_1100,In_1157);
nand U1418 (N_1418,In_1366,In_1096);
nand U1419 (N_1419,In_737,In_1203);
nor U1420 (N_1420,In_537,In_1330);
nor U1421 (N_1421,In_1453,In_1468);
nor U1422 (N_1422,In_488,In_1229);
or U1423 (N_1423,In_998,In_158);
and U1424 (N_1424,In_1330,In_1299);
nor U1425 (N_1425,In_719,In_243);
nor U1426 (N_1426,In_924,In_1272);
and U1427 (N_1427,In_31,In_1493);
nand U1428 (N_1428,In_739,In_650);
nor U1429 (N_1429,In_1032,In_398);
and U1430 (N_1430,In_643,In_234);
nor U1431 (N_1431,In_1481,In_933);
and U1432 (N_1432,In_200,In_84);
and U1433 (N_1433,In_262,In_1266);
nand U1434 (N_1434,In_434,In_1283);
or U1435 (N_1435,In_1414,In_796);
nand U1436 (N_1436,In_589,In_338);
nand U1437 (N_1437,In_934,In_254);
nor U1438 (N_1438,In_1258,In_19);
nand U1439 (N_1439,In_958,In_657);
nor U1440 (N_1440,In_968,In_513);
and U1441 (N_1441,In_740,In_1036);
or U1442 (N_1442,In_235,In_1475);
nand U1443 (N_1443,In_1482,In_213);
or U1444 (N_1444,In_601,In_890);
xnor U1445 (N_1445,In_1394,In_768);
or U1446 (N_1446,In_871,In_527);
nor U1447 (N_1447,In_1336,In_1072);
and U1448 (N_1448,In_1237,In_34);
nand U1449 (N_1449,In_303,In_152);
xor U1450 (N_1450,In_439,In_1101);
nor U1451 (N_1451,In_1499,In_1084);
nand U1452 (N_1452,In_1333,In_1063);
nor U1453 (N_1453,In_497,In_1151);
nand U1454 (N_1454,In_963,In_1010);
nand U1455 (N_1455,In_1073,In_890);
or U1456 (N_1456,In_778,In_1166);
or U1457 (N_1457,In_829,In_933);
and U1458 (N_1458,In_1146,In_184);
nor U1459 (N_1459,In_149,In_515);
and U1460 (N_1460,In_1284,In_887);
nor U1461 (N_1461,In_1321,In_727);
or U1462 (N_1462,In_150,In_1134);
and U1463 (N_1463,In_63,In_461);
and U1464 (N_1464,In_683,In_1435);
nor U1465 (N_1465,In_1248,In_1227);
and U1466 (N_1466,In_948,In_1022);
xor U1467 (N_1467,In_910,In_473);
nand U1468 (N_1468,In_766,In_41);
or U1469 (N_1469,In_1277,In_958);
nand U1470 (N_1470,In_1461,In_1206);
nor U1471 (N_1471,In_922,In_743);
nor U1472 (N_1472,In_264,In_488);
and U1473 (N_1473,In_199,In_768);
nor U1474 (N_1474,In_998,In_1417);
nor U1475 (N_1475,In_969,In_39);
xnor U1476 (N_1476,In_865,In_767);
and U1477 (N_1477,In_149,In_353);
and U1478 (N_1478,In_102,In_1362);
or U1479 (N_1479,In_82,In_561);
nor U1480 (N_1480,In_648,In_1185);
nor U1481 (N_1481,In_619,In_507);
nand U1482 (N_1482,In_290,In_582);
xnor U1483 (N_1483,In_447,In_1314);
or U1484 (N_1484,In_962,In_938);
and U1485 (N_1485,In_524,In_632);
nor U1486 (N_1486,In_1024,In_1009);
nor U1487 (N_1487,In_862,In_89);
and U1488 (N_1488,In_429,In_22);
nand U1489 (N_1489,In_977,In_1211);
nor U1490 (N_1490,In_285,In_1460);
nor U1491 (N_1491,In_827,In_721);
nand U1492 (N_1492,In_513,In_1195);
xor U1493 (N_1493,In_616,In_1408);
nand U1494 (N_1494,In_725,In_497);
and U1495 (N_1495,In_569,In_37);
nor U1496 (N_1496,In_1089,In_1106);
xor U1497 (N_1497,In_281,In_1213);
xnor U1498 (N_1498,In_620,In_243);
and U1499 (N_1499,In_310,In_1209);
and U1500 (N_1500,N_207,N_412);
nor U1501 (N_1501,N_1182,N_711);
or U1502 (N_1502,N_437,N_347);
nand U1503 (N_1503,N_384,N_730);
nor U1504 (N_1504,N_1415,N_953);
nor U1505 (N_1505,N_909,N_866);
nand U1506 (N_1506,N_910,N_714);
and U1507 (N_1507,N_978,N_1356);
nor U1508 (N_1508,N_1303,N_475);
nand U1509 (N_1509,N_980,N_1154);
nor U1510 (N_1510,N_115,N_441);
nor U1511 (N_1511,N_511,N_98);
nand U1512 (N_1512,N_774,N_1073);
nand U1513 (N_1513,N_884,N_18);
xnor U1514 (N_1514,N_1011,N_416);
and U1515 (N_1515,N_863,N_941);
and U1516 (N_1516,N_244,N_1165);
nor U1517 (N_1517,N_868,N_1321);
or U1518 (N_1518,N_531,N_1202);
nand U1519 (N_1519,N_930,N_1206);
xor U1520 (N_1520,N_638,N_1169);
and U1521 (N_1521,N_1163,N_718);
or U1522 (N_1522,N_522,N_1148);
and U1523 (N_1523,N_908,N_630);
and U1524 (N_1524,N_423,N_251);
and U1525 (N_1525,N_390,N_462);
or U1526 (N_1526,N_1194,N_794);
or U1527 (N_1527,N_1125,N_1292);
xnor U1528 (N_1528,N_440,N_450);
or U1529 (N_1529,N_698,N_839);
xnor U1530 (N_1530,N_518,N_681);
or U1531 (N_1531,N_742,N_969);
nand U1532 (N_1532,N_713,N_229);
xor U1533 (N_1533,N_1328,N_999);
or U1534 (N_1534,N_444,N_199);
nor U1535 (N_1535,N_596,N_302);
and U1536 (N_1536,N_1105,N_1254);
nor U1537 (N_1537,N_250,N_1121);
or U1538 (N_1538,N_466,N_300);
and U1539 (N_1539,N_110,N_1484);
and U1540 (N_1540,N_248,N_1079);
nor U1541 (N_1541,N_791,N_926);
and U1542 (N_1542,N_650,N_121);
nor U1543 (N_1543,N_1382,N_493);
or U1544 (N_1544,N_525,N_385);
xnor U1545 (N_1545,N_396,N_337);
and U1546 (N_1546,N_11,N_1210);
nor U1547 (N_1547,N_1358,N_407);
nor U1548 (N_1548,N_82,N_778);
nor U1549 (N_1549,N_776,N_338);
nand U1550 (N_1550,N_558,N_585);
nor U1551 (N_1551,N_619,N_867);
or U1552 (N_1552,N_798,N_1039);
xnor U1553 (N_1553,N_325,N_451);
nor U1554 (N_1554,N_777,N_335);
and U1555 (N_1555,N_286,N_1315);
xor U1556 (N_1556,N_67,N_34);
or U1557 (N_1557,N_436,N_590);
nor U1558 (N_1558,N_743,N_478);
and U1559 (N_1559,N_758,N_1471);
nor U1560 (N_1560,N_214,N_497);
nand U1561 (N_1561,N_262,N_1000);
or U1562 (N_1562,N_1343,N_963);
nor U1563 (N_1563,N_1304,N_329);
nand U1564 (N_1564,N_973,N_61);
or U1565 (N_1565,N_1115,N_123);
nand U1566 (N_1566,N_1008,N_636);
and U1567 (N_1567,N_1024,N_1272);
and U1568 (N_1568,N_130,N_405);
nor U1569 (N_1569,N_529,N_484);
nor U1570 (N_1570,N_1139,N_156);
nor U1571 (N_1571,N_660,N_1312);
nand U1572 (N_1572,N_879,N_945);
and U1573 (N_1573,N_306,N_534);
nor U1574 (N_1574,N_445,N_516);
nor U1575 (N_1575,N_775,N_595);
nand U1576 (N_1576,N_65,N_1371);
nand U1577 (N_1577,N_1112,N_1232);
or U1578 (N_1578,N_551,N_751);
nand U1579 (N_1579,N_747,N_369);
nand U1580 (N_1580,N_266,N_1166);
nand U1581 (N_1581,N_885,N_108);
or U1582 (N_1582,N_618,N_1111);
xnor U1583 (N_1583,N_716,N_1342);
and U1584 (N_1584,N_284,N_376);
xor U1585 (N_1585,N_557,N_899);
xnor U1586 (N_1586,N_1069,N_208);
nor U1587 (N_1587,N_1249,N_1239);
xnor U1588 (N_1588,N_318,N_1241);
or U1589 (N_1589,N_152,N_195);
and U1590 (N_1590,N_189,N_1458);
nand U1591 (N_1591,N_297,N_165);
nor U1592 (N_1592,N_95,N_797);
or U1593 (N_1593,N_750,N_196);
nand U1594 (N_1594,N_1215,N_962);
nor U1595 (N_1595,N_280,N_901);
and U1596 (N_1596,N_1089,N_1047);
nor U1597 (N_1597,N_952,N_1393);
nand U1598 (N_1598,N_896,N_243);
or U1599 (N_1599,N_1357,N_786);
and U1600 (N_1600,N_1481,N_245);
nand U1601 (N_1601,N_161,N_363);
nand U1602 (N_1602,N_1493,N_721);
nor U1603 (N_1603,N_129,N_366);
nor U1604 (N_1604,N_174,N_1301);
and U1605 (N_1605,N_1435,N_348);
xnor U1606 (N_1606,N_1270,N_771);
or U1607 (N_1607,N_27,N_998);
nor U1608 (N_1608,N_223,N_52);
xnor U1609 (N_1609,N_762,N_1346);
nor U1610 (N_1610,N_173,N_640);
xor U1611 (N_1611,N_455,N_308);
nand U1612 (N_1612,N_674,N_1457);
nor U1613 (N_1613,N_1242,N_904);
nand U1614 (N_1614,N_676,N_1437);
and U1615 (N_1615,N_468,N_625);
xnor U1616 (N_1616,N_274,N_1098);
nand U1617 (N_1617,N_712,N_1055);
or U1618 (N_1618,N_1281,N_1205);
or U1619 (N_1619,N_517,N_809);
and U1620 (N_1620,N_1175,N_486);
nand U1621 (N_1621,N_611,N_184);
nor U1622 (N_1622,N_1302,N_148);
nor U1623 (N_1623,N_1289,N_1368);
or U1624 (N_1624,N_1428,N_133);
and U1625 (N_1625,N_545,N_843);
nor U1626 (N_1626,N_1220,N_496);
nor U1627 (N_1627,N_205,N_501);
xnor U1628 (N_1628,N_175,N_279);
nand U1629 (N_1629,N_1200,N_1018);
nand U1630 (N_1630,N_819,N_857);
xnor U1631 (N_1631,N_773,N_1153);
nand U1632 (N_1632,N_305,N_1385);
nand U1633 (N_1633,N_1106,N_659);
or U1634 (N_1634,N_996,N_513);
and U1635 (N_1635,N_967,N_188);
nor U1636 (N_1636,N_1225,N_204);
and U1637 (N_1637,N_219,N_116);
xnor U1638 (N_1638,N_1258,N_1355);
nor U1639 (N_1639,N_1235,N_1454);
nor U1640 (N_1640,N_19,N_137);
nor U1641 (N_1641,N_586,N_893);
nor U1642 (N_1642,N_1447,N_955);
nand U1643 (N_1643,N_781,N_1275);
xor U1644 (N_1644,N_1196,N_275);
and U1645 (N_1645,N_1353,N_71);
or U1646 (N_1646,N_1077,N_120);
or U1647 (N_1647,N_1429,N_1188);
xnor U1648 (N_1648,N_21,N_160);
or U1649 (N_1649,N_815,N_0);
and U1650 (N_1650,N_111,N_601);
or U1651 (N_1651,N_1142,N_499);
or U1652 (N_1652,N_1341,N_26);
nand U1653 (N_1653,N_1020,N_291);
and U1654 (N_1654,N_1218,N_770);
and U1655 (N_1655,N_271,N_520);
nand U1656 (N_1656,N_902,N_1465);
nor U1657 (N_1657,N_1143,N_1134);
xor U1658 (N_1658,N_1237,N_991);
and U1659 (N_1659,N_324,N_974);
or U1660 (N_1660,N_944,N_479);
nand U1661 (N_1661,N_727,N_1063);
xnor U1662 (N_1662,N_483,N_1229);
or U1663 (N_1663,N_1045,N_487);
nand U1664 (N_1664,N_965,N_326);
nor U1665 (N_1665,N_512,N_372);
nor U1666 (N_1666,N_1460,N_629);
or U1667 (N_1667,N_594,N_14);
or U1668 (N_1668,N_992,N_850);
xor U1669 (N_1669,N_1442,N_72);
and U1670 (N_1670,N_510,N_1414);
xor U1671 (N_1671,N_805,N_634);
nand U1672 (N_1672,N_702,N_1226);
and U1673 (N_1673,N_1347,N_1168);
and U1674 (N_1674,N_959,N_972);
nor U1675 (N_1675,N_1036,N_270);
nand U1676 (N_1676,N_1244,N_624);
nand U1677 (N_1677,N_888,N_1431);
nand U1678 (N_1678,N_39,N_1262);
nor U1679 (N_1679,N_246,N_310);
xor U1680 (N_1680,N_443,N_10);
nor U1681 (N_1681,N_1388,N_894);
xnor U1682 (N_1682,N_535,N_51);
nor U1683 (N_1683,N_321,N_1391);
or U1684 (N_1684,N_332,N_482);
nand U1685 (N_1685,N_737,N_380);
and U1686 (N_1686,N_540,N_767);
or U1687 (N_1687,N_656,N_1082);
nand U1688 (N_1688,N_494,N_1441);
xnor U1689 (N_1689,N_89,N_821);
nand U1690 (N_1690,N_1472,N_150);
nor U1691 (N_1691,N_1479,N_1161);
nand U1692 (N_1692,N_217,N_807);
or U1693 (N_1693,N_544,N_315);
nor U1694 (N_1694,N_690,N_1495);
nand U1695 (N_1695,N_1470,N_485);
nor U1696 (N_1696,N_799,N_203);
nor U1697 (N_1697,N_1023,N_1030);
or U1698 (N_1698,N_1297,N_426);
nand U1699 (N_1699,N_1221,N_180);
nand U1700 (N_1700,N_1392,N_1141);
nand U1701 (N_1701,N_1359,N_1029);
and U1702 (N_1702,N_1213,N_1497);
nand U1703 (N_1703,N_938,N_228);
and U1704 (N_1704,N_951,N_446);
xor U1705 (N_1705,N_345,N_740);
or U1706 (N_1706,N_126,N_1027);
or U1707 (N_1707,N_114,N_745);
or U1708 (N_1708,N_355,N_361);
nand U1709 (N_1709,N_400,N_587);
and U1710 (N_1710,N_1394,N_1070);
nor U1711 (N_1711,N_556,N_1267);
and U1712 (N_1712,N_401,N_1138);
nand U1713 (N_1713,N_1440,N_593);
and U1714 (N_1714,N_685,N_564);
and U1715 (N_1715,N_382,N_1041);
or U1716 (N_1716,N_1491,N_1124);
nor U1717 (N_1717,N_1410,N_1318);
or U1718 (N_1718,N_1376,N_1260);
nand U1719 (N_1719,N_686,N_294);
or U1720 (N_1720,N_1240,N_688);
or U1721 (N_1721,N_46,N_500);
or U1722 (N_1722,N_1379,N_76);
or U1723 (N_1723,N_411,N_1311);
nand U1724 (N_1724,N_782,N_830);
nand U1725 (N_1725,N_198,N_81);
nor U1726 (N_1726,N_859,N_167);
or U1727 (N_1727,N_177,N_1155);
xor U1728 (N_1728,N_66,N_929);
and U1729 (N_1729,N_1286,N_779);
xor U1730 (N_1730,N_151,N_232);
nor U1731 (N_1731,N_1212,N_981);
and U1732 (N_1732,N_652,N_386);
nand U1733 (N_1733,N_925,N_362);
nor U1734 (N_1734,N_261,N_1372);
xnor U1735 (N_1735,N_74,N_1425);
nand U1736 (N_1736,N_808,N_371);
nand U1737 (N_1737,N_268,N_1436);
xnor U1738 (N_1738,N_273,N_873);
or U1739 (N_1739,N_1060,N_1120);
nor U1740 (N_1740,N_124,N_1373);
nand U1741 (N_1741,N_299,N_615);
nand U1742 (N_1742,N_768,N_1322);
or U1743 (N_1743,N_1421,N_1462);
nand U1744 (N_1744,N_60,N_643);
nor U1745 (N_1745,N_84,N_1145);
nand U1746 (N_1746,N_733,N_260);
nand U1747 (N_1747,N_637,N_1181);
nor U1748 (N_1748,N_1207,N_1477);
nand U1749 (N_1749,N_480,N_827);
and U1750 (N_1750,N_1264,N_1012);
nor U1751 (N_1751,N_367,N_724);
xnor U1752 (N_1752,N_706,N_1107);
nor U1753 (N_1753,N_612,N_1445);
or U1754 (N_1754,N_55,N_506);
or U1755 (N_1755,N_134,N_1004);
nor U1756 (N_1756,N_142,N_420);
nor U1757 (N_1757,N_920,N_934);
and U1758 (N_1758,N_766,N_1052);
or U1759 (N_1759,N_30,N_990);
or U1760 (N_1760,N_106,N_1149);
nor U1761 (N_1761,N_796,N_828);
nand U1762 (N_1762,N_616,N_536);
and U1763 (N_1763,N_703,N_1014);
xnor U1764 (N_1764,N_387,N_741);
nor U1765 (N_1765,N_464,N_806);
or U1766 (N_1766,N_1019,N_240);
nor U1767 (N_1767,N_633,N_1050);
or U1768 (N_1768,N_651,N_69);
or U1769 (N_1769,N_90,N_603);
nor U1770 (N_1770,N_679,N_1320);
nor U1771 (N_1771,N_1305,N_561);
or U1772 (N_1772,N_1405,N_892);
or U1773 (N_1773,N_1480,N_614);
xnor U1774 (N_1774,N_85,N_1354);
xor U1775 (N_1775,N_495,N_1430);
xor U1776 (N_1776,N_3,N_298);
nand U1777 (N_1777,N_453,N_789);
nand U1778 (N_1778,N_935,N_7);
and U1779 (N_1779,N_1310,N_1246);
nand U1780 (N_1780,N_97,N_1093);
nor U1781 (N_1781,N_169,N_811);
and U1782 (N_1782,N_1257,N_565);
nand U1783 (N_1783,N_54,N_833);
and U1784 (N_1784,N_442,N_1494);
xnor U1785 (N_1785,N_414,N_190);
or U1786 (N_1786,N_307,N_622);
or U1787 (N_1787,N_961,N_1193);
nand U1788 (N_1788,N_257,N_1174);
or U1789 (N_1789,N_1432,N_1411);
nor U1790 (N_1790,N_627,N_960);
and U1791 (N_1791,N_939,N_872);
nor U1792 (N_1792,N_572,N_870);
nand U1793 (N_1793,N_79,N_1015);
and U1794 (N_1794,N_209,N_547);
nand U1795 (N_1795,N_1486,N_289);
nor U1796 (N_1796,N_1033,N_176);
or U1797 (N_1797,N_258,N_818);
and U1798 (N_1798,N_1406,N_1048);
and U1799 (N_1799,N_1236,N_431);
nand U1800 (N_1800,N_105,N_122);
or U1801 (N_1801,N_657,N_1279);
or U1802 (N_1802,N_249,N_1488);
xor U1803 (N_1803,N_201,N_56);
nand U1804 (N_1804,N_182,N_140);
nor U1805 (N_1805,N_1467,N_340);
nand U1806 (N_1806,N_906,N_296);
or U1807 (N_1807,N_17,N_1103);
and U1808 (N_1808,N_507,N_937);
nand U1809 (N_1809,N_1101,N_1043);
nand U1810 (N_1810,N_1327,N_38);
or U1811 (N_1811,N_845,N_555);
nand U1812 (N_1812,N_1072,N_319);
or U1813 (N_1813,N_581,N_1475);
nand U1814 (N_1814,N_829,N_234);
or U1815 (N_1815,N_322,N_438);
nand U1816 (N_1816,N_989,N_1046);
nor U1817 (N_1817,N_823,N_589);
nor U1818 (N_1818,N_1243,N_871);
and U1819 (N_1819,N_1197,N_765);
and U1820 (N_1820,N_1485,N_1351);
xnor U1821 (N_1821,N_1126,N_567);
nor U1822 (N_1822,N_1028,N_1438);
and U1823 (N_1823,N_64,N_552);
or U1824 (N_1824,N_1150,N_311);
and U1825 (N_1825,N_1177,N_966);
and U1826 (N_1826,N_623,N_881);
nand U1827 (N_1827,N_1058,N_725);
xor U1828 (N_1828,N_736,N_433);
xor U1829 (N_1829,N_639,N_695);
nand U1830 (N_1830,N_1031,N_342);
or U1831 (N_1831,N_127,N_530);
and U1832 (N_1832,N_793,N_617);
xor U1833 (N_1833,N_1295,N_1152);
or U1834 (N_1834,N_215,N_1147);
and U1835 (N_1835,N_986,N_157);
and U1836 (N_1836,N_379,N_672);
and U1837 (N_1837,N_202,N_705);
or U1838 (N_1838,N_943,N_192);
or U1839 (N_1839,N_269,N_699);
nor U1840 (N_1840,N_864,N_381);
nor U1841 (N_1841,N_119,N_1131);
and U1842 (N_1842,N_502,N_47);
and U1843 (N_1843,N_971,N_521);
and U1844 (N_1844,N_312,N_350);
nor U1845 (N_1845,N_149,N_1066);
and U1846 (N_1846,N_566,N_1451);
xor U1847 (N_1847,N_1104,N_48);
xnor U1848 (N_1848,N_792,N_1132);
or U1849 (N_1849,N_508,N_194);
xnor U1850 (N_1850,N_31,N_1336);
nor U1851 (N_1851,N_1418,N_252);
nand U1852 (N_1852,N_764,N_210);
nor U1853 (N_1853,N_950,N_738);
nor U1854 (N_1854,N_370,N_1309);
and U1855 (N_1855,N_824,N_1287);
and U1856 (N_1856,N_383,N_206);
nand U1857 (N_1857,N_1350,N_23);
or U1858 (N_1858,N_936,N_1146);
and U1859 (N_1859,N_877,N_1276);
nand U1860 (N_1860,N_1171,N_976);
xor U1861 (N_1861,N_1054,N_1209);
or U1862 (N_1862,N_1071,N_1159);
or U1863 (N_1863,N_422,N_20);
xnor U1864 (N_1864,N_221,N_1378);
and U1865 (N_1865,N_1059,N_461);
nand U1866 (N_1866,N_358,N_1192);
nor U1867 (N_1867,N_1364,N_836);
nor U1868 (N_1868,N_492,N_1455);
nand U1869 (N_1869,N_1091,N_145);
nand U1870 (N_1870,N_1416,N_220);
nor U1871 (N_1871,N_1306,N_1375);
nand U1872 (N_1872,N_1195,N_942);
and U1873 (N_1873,N_720,N_1231);
xnor U1874 (N_1874,N_351,N_349);
nor U1875 (N_1875,N_15,N_752);
or U1876 (N_1876,N_317,N_354);
nor U1877 (N_1877,N_285,N_1384);
or U1878 (N_1878,N_1298,N_1299);
nor U1879 (N_1879,N_1399,N_684);
nor U1880 (N_1880,N_1238,N_855);
or U1881 (N_1881,N_331,N_117);
nand U1882 (N_1882,N_1398,N_421);
and U1883 (N_1883,N_1496,N_1330);
and U1884 (N_1884,N_86,N_333);
nand U1885 (N_1885,N_406,N_1157);
and U1886 (N_1886,N_1293,N_101);
and U1887 (N_1887,N_598,N_846);
nand U1888 (N_1888,N_236,N_553);
nor U1889 (N_1889,N_293,N_309);
nand U1890 (N_1890,N_680,N_1332);
nor U1891 (N_1891,N_527,N_729);
nand U1892 (N_1892,N_186,N_419);
nand U1893 (N_1893,N_1214,N_940);
and U1894 (N_1894,N_670,N_391);
nand U1895 (N_1895,N_532,N_844);
nor U1896 (N_1896,N_1317,N_1329);
xnor U1897 (N_1897,N_467,N_1268);
xnor U1898 (N_1898,N_822,N_498);
xnor U1899 (N_1899,N_1427,N_895);
nand U1900 (N_1900,N_912,N_922);
and U1901 (N_1901,N_979,N_931);
nor U1902 (N_1902,N_170,N_24);
nor U1903 (N_1903,N_1017,N_399);
nor U1904 (N_1904,N_728,N_1248);
nand U1905 (N_1905,N_689,N_179);
and U1906 (N_1906,N_1040,N_330);
nand U1907 (N_1907,N_99,N_924);
nor U1908 (N_1908,N_216,N_1374);
or U1909 (N_1909,N_550,N_631);
and U1910 (N_1910,N_984,N_983);
nor U1911 (N_1911,N_282,N_1136);
xnor U1912 (N_1912,N_832,N_577);
or U1913 (N_1913,N_837,N_1278);
nor U1914 (N_1914,N_1233,N_424);
and U1915 (N_1915,N_230,N_323);
nor U1916 (N_1916,N_1412,N_118);
or U1917 (N_1917,N_856,N_227);
and U1918 (N_1918,N_238,N_584);
or U1919 (N_1919,N_37,N_138);
nand U1920 (N_1920,N_1360,N_1334);
nor U1921 (N_1921,N_891,N_648);
or U1922 (N_1922,N_543,N_1062);
and U1923 (N_1923,N_887,N_375);
and U1924 (N_1924,N_320,N_897);
nand U1925 (N_1925,N_476,N_1408);
and U1926 (N_1926,N_907,N_1400);
or U1927 (N_1927,N_1010,N_237);
and U1928 (N_1928,N_958,N_814);
and U1929 (N_1929,N_1227,N_570);
nor U1930 (N_1930,N_1397,N_504);
and U1931 (N_1931,N_388,N_430);
and U1932 (N_1932,N_49,N_1273);
nor U1933 (N_1933,N_605,N_574);
nor U1934 (N_1934,N_212,N_353);
nor U1935 (N_1935,N_398,N_235);
nand U1936 (N_1936,N_903,N_505);
or U1937 (N_1937,N_1263,N_715);
nand U1938 (N_1938,N_641,N_490);
nand U1939 (N_1939,N_826,N_700);
or U1940 (N_1940,N_181,N_1296);
nand U1941 (N_1941,N_1032,N_287);
nand U1942 (N_1942,N_928,N_1130);
or U1943 (N_1943,N_772,N_1016);
and U1944 (N_1944,N_1198,N_604);
or U1945 (N_1945,N_346,N_1002);
nand U1946 (N_1946,N_91,N_465);
xor U1947 (N_1947,N_1316,N_57);
nor U1948 (N_1948,N_1224,N_1389);
and U1949 (N_1949,N_327,N_6);
nor U1950 (N_1950,N_187,N_1108);
nor U1951 (N_1951,N_92,N_70);
or U1952 (N_1952,N_459,N_193);
xor U1953 (N_1953,N_880,N_932);
or U1954 (N_1954,N_816,N_946);
nor U1955 (N_1955,N_1127,N_343);
nor U1956 (N_1956,N_1109,N_259);
or U1957 (N_1957,N_949,N_842);
or U1958 (N_1958,N_28,N_1068);
nor U1959 (N_1959,N_143,N_1122);
and U1960 (N_1960,N_447,N_1387);
or U1961 (N_1961,N_1114,N_1478);
xnor U1962 (N_1962,N_434,N_852);
nor U1963 (N_1963,N_1271,N_862);
or U1964 (N_1964,N_1319,N_1366);
or U1965 (N_1965,N_726,N_449);
nor U1966 (N_1966,N_982,N_1449);
and U1967 (N_1967,N_8,N_392);
or U1968 (N_1968,N_1487,N_834);
or U1969 (N_1969,N_609,N_83);
nor U1970 (N_1970,N_1291,N_748);
nor U1971 (N_1971,N_523,N_1474);
nor U1972 (N_1972,N_109,N_890);
nand U1973 (N_1973,N_32,N_673);
or U1974 (N_1974,N_1003,N_933);
or U1975 (N_1975,N_569,N_1075);
or U1976 (N_1976,N_29,N_1219);
or U1977 (N_1977,N_1261,N_1369);
and U1978 (N_1978,N_1468,N_882);
or U1979 (N_1979,N_666,N_146);
or U1980 (N_1980,N_73,N_608);
nor U1981 (N_1981,N_154,N_1088);
nor U1982 (N_1982,N_415,N_103);
nor U1983 (N_1983,N_1083,N_264);
nand U1984 (N_1984,N_1282,N_1026);
nor U1985 (N_1985,N_1056,N_410);
nand U1986 (N_1986,N_77,N_841);
or U1987 (N_1987,N_1118,N_677);
and U1988 (N_1988,N_503,N_239);
and U1989 (N_1989,N_977,N_548);
and U1990 (N_1990,N_1423,N_1404);
or U1991 (N_1991,N_178,N_1084);
nand U1992 (N_1992,N_997,N_755);
or U1993 (N_1993,N_1135,N_1160);
and U1994 (N_1994,N_1483,N_803);
nand U1995 (N_1995,N_1170,N_88);
nor U1996 (N_1996,N_970,N_265);
or U1997 (N_1997,N_78,N_948);
and U1998 (N_1998,N_225,N_344);
nor U1999 (N_1999,N_136,N_377);
and U2000 (N_2000,N_607,N_701);
nor U2001 (N_2001,N_25,N_654);
xnor U2002 (N_2002,N_1167,N_96);
nor U2003 (N_2003,N_1259,N_1476);
and U2004 (N_2004,N_1189,N_1381);
xnor U2005 (N_2005,N_374,N_1380);
nand U2006 (N_2006,N_917,N_472);
or U2007 (N_2007,N_1092,N_1349);
and U2008 (N_2008,N_35,N_112);
nor U2009 (N_2009,N_1172,N_665);
nor U2010 (N_2010,N_644,N_1223);
and U2011 (N_2011,N_272,N_810);
or U2012 (N_2012,N_1461,N_709);
and U2013 (N_2013,N_840,N_364);
or U2014 (N_2014,N_357,N_671);
nor U2015 (N_2015,N_1489,N_290);
and U2016 (N_2016,N_1140,N_255);
nor U2017 (N_2017,N_22,N_93);
nand U2018 (N_2018,N_439,N_213);
or U2019 (N_2019,N_102,N_597);
nor U2020 (N_2020,N_1333,N_785);
or U2021 (N_2021,N_515,N_1419);
nand U2022 (N_2022,N_919,N_172);
nor U2023 (N_2023,N_563,N_964);
and U2024 (N_2024,N_113,N_40);
or U2025 (N_2025,N_800,N_1217);
or U2026 (N_2026,N_1025,N_168);
nor U2027 (N_2027,N_458,N_707);
nor U2028 (N_2028,N_226,N_1323);
nand U2029 (N_2029,N_254,N_403);
nor U2030 (N_2030,N_708,N_1129);
nand U2031 (N_2031,N_549,N_1076);
or U2032 (N_2032,N_1482,N_1211);
xor U2033 (N_2033,N_132,N_838);
and U2034 (N_2034,N_1080,N_1203);
nand U2035 (N_2035,N_848,N_1187);
and U2036 (N_2036,N_861,N_1294);
nand U2037 (N_2037,N_546,N_573);
nor U2038 (N_2038,N_682,N_1022);
nand U2039 (N_2039,N_1424,N_1277);
and U2040 (N_2040,N_1288,N_1390);
and U2041 (N_2041,N_128,N_1123);
nand U2042 (N_2042,N_578,N_1173);
nand U2043 (N_2043,N_393,N_509);
and U2044 (N_2044,N_1178,N_1256);
nor U2045 (N_2045,N_1184,N_62);
or U2046 (N_2046,N_418,N_1191);
or U2047 (N_2047,N_491,N_1090);
and U2048 (N_2048,N_658,N_211);
xor U2049 (N_2049,N_1067,N_739);
nand U2050 (N_2050,N_1097,N_968);
and U2051 (N_2051,N_1006,N_722);
or U2052 (N_2052,N_12,N_267);
nor U2053 (N_2053,N_528,N_1250);
or U2054 (N_2054,N_1164,N_1344);
nor U2055 (N_2055,N_80,N_1377);
xnor U2056 (N_2056,N_191,N_303);
or U2057 (N_2057,N_328,N_1180);
nor U2058 (N_2058,N_394,N_1452);
or U2059 (N_2059,N_147,N_378);
nand U2060 (N_2060,N_1446,N_1201);
and U2061 (N_2061,N_360,N_1456);
nor U2062 (N_2062,N_313,N_519);
nor U2063 (N_2063,N_1339,N_1469);
and U2064 (N_2064,N_921,N_1049);
and U2065 (N_2065,N_975,N_987);
or U2066 (N_2066,N_1252,N_1179);
and U2067 (N_2067,N_1099,N_760);
or U2068 (N_2068,N_473,N_417);
nor U2069 (N_2069,N_457,N_1499);
or U2070 (N_2070,N_645,N_1208);
or U2071 (N_2071,N_668,N_356);
nand U2072 (N_2072,N_474,N_352);
and U2073 (N_2073,N_1086,N_456);
nand U2074 (N_2074,N_813,N_1065);
or U2075 (N_2075,N_704,N_683);
or U2076 (N_2076,N_1396,N_1313);
nand U2077 (N_2077,N_295,N_1269);
and U2078 (N_2078,N_1137,N_1051);
nand U2079 (N_2079,N_1,N_185);
and U2080 (N_2080,N_144,N_1308);
nand U2081 (N_2081,N_1362,N_1128);
or U2082 (N_2082,N_43,N_131);
or U2083 (N_2083,N_1034,N_1087);
and U2084 (N_2084,N_831,N_542);
nand U2085 (N_2085,N_1300,N_642);
or U2086 (N_2086,N_583,N_647);
nor U2087 (N_2087,N_409,N_1352);
and U2088 (N_2088,N_277,N_397);
and U2089 (N_2089,N_1324,N_664);
nand U2090 (N_2090,N_620,N_1367);
nor U2091 (N_2091,N_107,N_783);
and U2092 (N_2092,N_1005,N_59);
nand U2093 (N_2093,N_402,N_1222);
and U2094 (N_2094,N_592,N_1403);
nand U2095 (N_2095,N_749,N_825);
nor U2096 (N_2096,N_693,N_1162);
nand U2097 (N_2097,N_448,N_1439);
nor U2098 (N_2098,N_802,N_1265);
nor U2099 (N_2099,N_359,N_1464);
nor U2100 (N_2100,N_104,N_42);
xnor U2101 (N_2101,N_1348,N_166);
nand U2102 (N_2102,N_278,N_1365);
nand U2103 (N_2103,N_281,N_1245);
xor U2104 (N_2104,N_675,N_579);
or U2105 (N_2105,N_878,N_985);
or U2106 (N_2106,N_197,N_1144);
nand U2107 (N_2107,N_1021,N_1314);
and U2108 (N_2108,N_854,N_541);
xor U2109 (N_2109,N_1156,N_719);
nor U2110 (N_2110,N_757,N_1402);
and U2111 (N_2111,N_1085,N_1094);
nor U2112 (N_2112,N_1283,N_562);
nor U2113 (N_2113,N_1158,N_898);
or U2114 (N_2114,N_1183,N_600);
nand U2115 (N_2115,N_1044,N_1228);
xor U2116 (N_2116,N_50,N_694);
nand U2117 (N_2117,N_538,N_163);
and U2118 (N_2118,N_956,N_316);
nand U2119 (N_2119,N_1417,N_817);
or U2120 (N_2120,N_869,N_162);
nor U2121 (N_2121,N_341,N_591);
nor U2122 (N_2122,N_911,N_1492);
or U2123 (N_2123,N_626,N_847);
xnor U2124 (N_2124,N_865,N_68);
xnor U2125 (N_2125,N_288,N_1064);
nand U2126 (N_2126,N_753,N_224);
and U2127 (N_2127,N_649,N_1466);
or U2128 (N_2128,N_632,N_253);
nand U2129 (N_2129,N_915,N_914);
or U2130 (N_2130,N_432,N_33);
and U2131 (N_2131,N_1117,N_851);
and U2132 (N_2132,N_1042,N_905);
and U2133 (N_2133,N_1363,N_45);
and U2134 (N_2134,N_1426,N_995);
or U2135 (N_2135,N_795,N_155);
xor U2136 (N_2136,N_1420,N_404);
nor U2137 (N_2137,N_53,N_678);
nor U2138 (N_2138,N_628,N_1204);
nor U2139 (N_2139,N_787,N_784);
and U2140 (N_2140,N_1116,N_613);
or U2141 (N_2141,N_655,N_1266);
nor U2142 (N_2142,N_481,N_723);
and U2143 (N_2143,N_1444,N_158);
nand U2144 (N_2144,N_283,N_1401);
nand U2145 (N_2145,N_588,N_1078);
nand U2146 (N_2146,N_4,N_233);
nand U2147 (N_2147,N_804,N_2);
and U2148 (N_2148,N_1013,N_875);
or U2149 (N_2149,N_1234,N_554);
nor U2150 (N_2150,N_769,N_662);
xor U2151 (N_2151,N_756,N_744);
or U2152 (N_2152,N_1386,N_1274);
and U2153 (N_2153,N_1450,N_923);
or U2154 (N_2154,N_1335,N_860);
nand U2155 (N_2155,N_1151,N_1199);
or U2156 (N_2156,N_171,N_276);
nand U2157 (N_2157,N_883,N_1434);
and U2158 (N_2158,N_100,N_454);
nor U2159 (N_2159,N_1253,N_746);
or U2160 (N_2160,N_988,N_947);
or U2161 (N_2161,N_599,N_1413);
and U2162 (N_2162,N_610,N_1009);
nor U2163 (N_2163,N_489,N_470);
or U2164 (N_2164,N_1284,N_1459);
nand U2165 (N_2165,N_304,N_858);
nor U2166 (N_2166,N_425,N_314);
xor U2167 (N_2167,N_141,N_1255);
xor U2168 (N_2168,N_5,N_1053);
nand U2169 (N_2169,N_580,N_560);
and U2170 (N_2170,N_1361,N_87);
or U2171 (N_2171,N_646,N_13);
xor U2172 (N_2172,N_761,N_993);
xor U2173 (N_2173,N_1338,N_1035);
or U2174 (N_2174,N_1230,N_927);
and U2175 (N_2175,N_1433,N_1490);
nor U2176 (N_2176,N_1325,N_717);
nand U2177 (N_2177,N_900,N_477);
nand U2178 (N_2178,N_606,N_732);
and U2179 (N_2179,N_452,N_692);
or U2180 (N_2180,N_153,N_292);
nand U2181 (N_2181,N_218,N_691);
and U2182 (N_2182,N_334,N_1473);
or U2183 (N_2183,N_687,N_395);
nand U2184 (N_2184,N_1453,N_231);
nor U2185 (N_2185,N_801,N_874);
nor U2186 (N_2186,N_222,N_94);
xor U2187 (N_2187,N_731,N_1186);
nor U2188 (N_2188,N_63,N_1037);
or U2189 (N_2189,N_1285,N_621);
and U2190 (N_2190,N_735,N_954);
xnor U2191 (N_2191,N_9,N_435);
nor U2192 (N_2192,N_58,N_1290);
or U2193 (N_2193,N_582,N_514);
or U2194 (N_2194,N_812,N_1443);
xor U2195 (N_2195,N_853,N_1463);
and U2196 (N_2196,N_200,N_571);
and U2197 (N_2197,N_164,N_916);
xor U2198 (N_2198,N_1007,N_533);
nor U2199 (N_2199,N_820,N_526);
nand U2200 (N_2200,N_918,N_663);
nand U2201 (N_2201,N_559,N_602);
and U2202 (N_2202,N_1133,N_1326);
and U2203 (N_2203,N_1422,N_763);
nor U2204 (N_2204,N_16,N_339);
and U2205 (N_2205,N_524,N_1001);
xor U2206 (N_2206,N_242,N_788);
nor U2207 (N_2207,N_1395,N_336);
or U2208 (N_2208,N_1190,N_575);
nand U2209 (N_2209,N_1307,N_365);
or U2210 (N_2210,N_1110,N_913);
nand U2211 (N_2211,N_653,N_957);
nor U2212 (N_2212,N_1407,N_75);
nor U2213 (N_2213,N_790,N_1119);
nand U2214 (N_2214,N_1345,N_754);
nor U2215 (N_2215,N_1095,N_1102);
or U2216 (N_2216,N_710,N_389);
and U2217 (N_2217,N_1383,N_576);
nor U2218 (N_2218,N_635,N_469);
nor U2219 (N_2219,N_368,N_256);
nor U2220 (N_2220,N_1057,N_889);
or U2221 (N_2221,N_1370,N_1081);
xnor U2222 (N_2222,N_1409,N_44);
or U2223 (N_2223,N_696,N_1074);
nand U2224 (N_2224,N_667,N_1331);
and U2225 (N_2225,N_427,N_780);
or U2226 (N_2226,N_1216,N_1038);
and U2227 (N_2227,N_408,N_669);
and U2228 (N_2228,N_1448,N_697);
nand U2229 (N_2229,N_428,N_661);
and U2230 (N_2230,N_886,N_994);
nand U2231 (N_2231,N_1247,N_759);
nand U2232 (N_2232,N_1337,N_373);
nor U2233 (N_2233,N_460,N_247);
and U2234 (N_2234,N_568,N_125);
nor U2235 (N_2235,N_1251,N_849);
nor U2236 (N_2236,N_539,N_429);
nor U2237 (N_2237,N_1113,N_1061);
nand U2238 (N_2238,N_139,N_1340);
nor U2239 (N_2239,N_135,N_1176);
nor U2240 (N_2240,N_471,N_183);
nor U2241 (N_2241,N_734,N_1280);
nor U2242 (N_2242,N_241,N_835);
or U2243 (N_2243,N_36,N_876);
nand U2244 (N_2244,N_488,N_41);
nand U2245 (N_2245,N_159,N_263);
nand U2246 (N_2246,N_1100,N_463);
and U2247 (N_2247,N_1096,N_537);
nand U2248 (N_2248,N_1185,N_301);
nand U2249 (N_2249,N_1498,N_413);
nor U2250 (N_2250,N_769,N_135);
xnor U2251 (N_2251,N_569,N_1133);
or U2252 (N_2252,N_544,N_698);
nand U2253 (N_2253,N_1428,N_1103);
nor U2254 (N_2254,N_250,N_1150);
xor U2255 (N_2255,N_519,N_553);
or U2256 (N_2256,N_1080,N_906);
and U2257 (N_2257,N_747,N_1073);
and U2258 (N_2258,N_1444,N_130);
nor U2259 (N_2259,N_1462,N_555);
or U2260 (N_2260,N_1014,N_799);
xor U2261 (N_2261,N_431,N_1184);
nor U2262 (N_2262,N_946,N_209);
and U2263 (N_2263,N_268,N_340);
xnor U2264 (N_2264,N_3,N_380);
nand U2265 (N_2265,N_1293,N_520);
nand U2266 (N_2266,N_270,N_1303);
nor U2267 (N_2267,N_1121,N_162);
and U2268 (N_2268,N_1061,N_1415);
or U2269 (N_2269,N_588,N_204);
nor U2270 (N_2270,N_1245,N_1057);
nand U2271 (N_2271,N_1272,N_242);
nand U2272 (N_2272,N_1251,N_380);
and U2273 (N_2273,N_779,N_639);
nor U2274 (N_2274,N_67,N_1040);
xor U2275 (N_2275,N_1037,N_1163);
and U2276 (N_2276,N_107,N_669);
and U2277 (N_2277,N_1358,N_196);
or U2278 (N_2278,N_1453,N_245);
or U2279 (N_2279,N_1009,N_258);
and U2280 (N_2280,N_630,N_449);
nand U2281 (N_2281,N_119,N_877);
and U2282 (N_2282,N_1277,N_1048);
nor U2283 (N_2283,N_4,N_978);
or U2284 (N_2284,N_365,N_246);
and U2285 (N_2285,N_99,N_1315);
nand U2286 (N_2286,N_874,N_1045);
nand U2287 (N_2287,N_854,N_774);
nand U2288 (N_2288,N_345,N_1046);
nand U2289 (N_2289,N_840,N_44);
or U2290 (N_2290,N_781,N_1217);
xnor U2291 (N_2291,N_782,N_750);
xor U2292 (N_2292,N_1418,N_1044);
nor U2293 (N_2293,N_1379,N_54);
nand U2294 (N_2294,N_1460,N_1224);
nand U2295 (N_2295,N_666,N_928);
nor U2296 (N_2296,N_1031,N_171);
and U2297 (N_2297,N_1136,N_1328);
nand U2298 (N_2298,N_917,N_693);
nand U2299 (N_2299,N_103,N_1405);
or U2300 (N_2300,N_1034,N_709);
and U2301 (N_2301,N_949,N_504);
and U2302 (N_2302,N_962,N_1244);
nor U2303 (N_2303,N_29,N_1030);
nor U2304 (N_2304,N_230,N_1357);
or U2305 (N_2305,N_1285,N_1104);
nand U2306 (N_2306,N_192,N_1291);
nor U2307 (N_2307,N_869,N_695);
nor U2308 (N_2308,N_555,N_59);
or U2309 (N_2309,N_753,N_826);
nand U2310 (N_2310,N_284,N_175);
nor U2311 (N_2311,N_597,N_169);
xnor U2312 (N_2312,N_1352,N_517);
nor U2313 (N_2313,N_271,N_1307);
and U2314 (N_2314,N_276,N_932);
nor U2315 (N_2315,N_307,N_666);
nor U2316 (N_2316,N_1354,N_519);
and U2317 (N_2317,N_518,N_667);
nand U2318 (N_2318,N_636,N_95);
nand U2319 (N_2319,N_1372,N_1344);
nand U2320 (N_2320,N_284,N_1211);
nand U2321 (N_2321,N_829,N_781);
or U2322 (N_2322,N_783,N_711);
nand U2323 (N_2323,N_771,N_1081);
and U2324 (N_2324,N_882,N_1482);
or U2325 (N_2325,N_1130,N_1318);
or U2326 (N_2326,N_1267,N_787);
nor U2327 (N_2327,N_1073,N_971);
nor U2328 (N_2328,N_613,N_456);
and U2329 (N_2329,N_381,N_1302);
nor U2330 (N_2330,N_48,N_800);
xnor U2331 (N_2331,N_1176,N_102);
and U2332 (N_2332,N_469,N_1099);
or U2333 (N_2333,N_1414,N_32);
nor U2334 (N_2334,N_1262,N_942);
nor U2335 (N_2335,N_915,N_304);
xnor U2336 (N_2336,N_1245,N_1087);
nor U2337 (N_2337,N_635,N_314);
or U2338 (N_2338,N_402,N_665);
xor U2339 (N_2339,N_892,N_1184);
nor U2340 (N_2340,N_66,N_941);
xnor U2341 (N_2341,N_713,N_400);
nor U2342 (N_2342,N_1158,N_864);
nand U2343 (N_2343,N_325,N_1159);
and U2344 (N_2344,N_1208,N_541);
or U2345 (N_2345,N_202,N_1018);
xnor U2346 (N_2346,N_93,N_72);
or U2347 (N_2347,N_666,N_710);
and U2348 (N_2348,N_1279,N_820);
xor U2349 (N_2349,N_455,N_972);
nand U2350 (N_2350,N_392,N_1328);
nor U2351 (N_2351,N_1016,N_1445);
or U2352 (N_2352,N_227,N_896);
and U2353 (N_2353,N_187,N_1035);
xnor U2354 (N_2354,N_1003,N_420);
nor U2355 (N_2355,N_669,N_7);
nor U2356 (N_2356,N_1050,N_149);
or U2357 (N_2357,N_1091,N_473);
xnor U2358 (N_2358,N_1093,N_1243);
and U2359 (N_2359,N_178,N_906);
xor U2360 (N_2360,N_421,N_200);
xnor U2361 (N_2361,N_393,N_222);
or U2362 (N_2362,N_338,N_226);
or U2363 (N_2363,N_1046,N_633);
or U2364 (N_2364,N_55,N_61);
or U2365 (N_2365,N_1152,N_1116);
nand U2366 (N_2366,N_281,N_491);
and U2367 (N_2367,N_1473,N_908);
and U2368 (N_2368,N_542,N_858);
or U2369 (N_2369,N_1059,N_309);
and U2370 (N_2370,N_423,N_628);
xor U2371 (N_2371,N_1245,N_1099);
and U2372 (N_2372,N_790,N_157);
nor U2373 (N_2373,N_899,N_884);
nor U2374 (N_2374,N_1497,N_266);
nand U2375 (N_2375,N_706,N_692);
and U2376 (N_2376,N_538,N_434);
or U2377 (N_2377,N_329,N_635);
or U2378 (N_2378,N_1238,N_1130);
xor U2379 (N_2379,N_1127,N_1085);
nand U2380 (N_2380,N_535,N_516);
nor U2381 (N_2381,N_985,N_210);
nand U2382 (N_2382,N_810,N_370);
or U2383 (N_2383,N_239,N_1390);
and U2384 (N_2384,N_933,N_1410);
nor U2385 (N_2385,N_711,N_57);
nor U2386 (N_2386,N_55,N_1174);
or U2387 (N_2387,N_1118,N_1257);
nand U2388 (N_2388,N_780,N_1291);
and U2389 (N_2389,N_898,N_109);
nor U2390 (N_2390,N_1385,N_678);
nor U2391 (N_2391,N_1060,N_144);
or U2392 (N_2392,N_1068,N_86);
and U2393 (N_2393,N_1293,N_720);
and U2394 (N_2394,N_1488,N_968);
nand U2395 (N_2395,N_1164,N_1461);
nand U2396 (N_2396,N_52,N_311);
and U2397 (N_2397,N_1087,N_1475);
or U2398 (N_2398,N_1259,N_697);
and U2399 (N_2399,N_967,N_1012);
or U2400 (N_2400,N_407,N_518);
and U2401 (N_2401,N_62,N_377);
or U2402 (N_2402,N_1234,N_791);
xor U2403 (N_2403,N_1376,N_1236);
xnor U2404 (N_2404,N_652,N_1476);
nand U2405 (N_2405,N_761,N_622);
nand U2406 (N_2406,N_983,N_1183);
or U2407 (N_2407,N_1004,N_1215);
nor U2408 (N_2408,N_309,N_453);
or U2409 (N_2409,N_1184,N_151);
nand U2410 (N_2410,N_193,N_836);
xor U2411 (N_2411,N_716,N_543);
xnor U2412 (N_2412,N_262,N_990);
nor U2413 (N_2413,N_457,N_19);
xor U2414 (N_2414,N_1264,N_312);
nand U2415 (N_2415,N_1223,N_1104);
or U2416 (N_2416,N_1217,N_714);
or U2417 (N_2417,N_673,N_1451);
and U2418 (N_2418,N_854,N_1020);
and U2419 (N_2419,N_1151,N_1230);
or U2420 (N_2420,N_1384,N_246);
and U2421 (N_2421,N_240,N_1322);
and U2422 (N_2422,N_1133,N_40);
or U2423 (N_2423,N_907,N_453);
nor U2424 (N_2424,N_347,N_1270);
nor U2425 (N_2425,N_626,N_267);
or U2426 (N_2426,N_1046,N_1430);
xor U2427 (N_2427,N_1089,N_420);
nand U2428 (N_2428,N_793,N_905);
and U2429 (N_2429,N_480,N_165);
nand U2430 (N_2430,N_1239,N_150);
nor U2431 (N_2431,N_313,N_111);
nor U2432 (N_2432,N_382,N_989);
nor U2433 (N_2433,N_1103,N_1435);
nand U2434 (N_2434,N_1438,N_936);
or U2435 (N_2435,N_520,N_179);
and U2436 (N_2436,N_1214,N_532);
nor U2437 (N_2437,N_355,N_551);
nand U2438 (N_2438,N_1306,N_220);
xor U2439 (N_2439,N_354,N_16);
or U2440 (N_2440,N_1114,N_567);
nor U2441 (N_2441,N_44,N_358);
nand U2442 (N_2442,N_1331,N_928);
and U2443 (N_2443,N_46,N_185);
or U2444 (N_2444,N_621,N_656);
and U2445 (N_2445,N_410,N_685);
and U2446 (N_2446,N_128,N_888);
xor U2447 (N_2447,N_62,N_267);
or U2448 (N_2448,N_591,N_63);
nand U2449 (N_2449,N_1125,N_354);
nor U2450 (N_2450,N_1231,N_512);
nor U2451 (N_2451,N_634,N_1380);
nand U2452 (N_2452,N_995,N_951);
nand U2453 (N_2453,N_1385,N_1082);
nor U2454 (N_2454,N_252,N_386);
nor U2455 (N_2455,N_356,N_486);
nand U2456 (N_2456,N_1243,N_756);
and U2457 (N_2457,N_1199,N_1402);
or U2458 (N_2458,N_1316,N_612);
and U2459 (N_2459,N_37,N_35);
nand U2460 (N_2460,N_508,N_642);
or U2461 (N_2461,N_92,N_116);
nand U2462 (N_2462,N_429,N_940);
or U2463 (N_2463,N_816,N_1126);
nand U2464 (N_2464,N_1423,N_1228);
nand U2465 (N_2465,N_1251,N_195);
nand U2466 (N_2466,N_909,N_973);
nor U2467 (N_2467,N_1239,N_285);
or U2468 (N_2468,N_47,N_981);
nor U2469 (N_2469,N_264,N_897);
or U2470 (N_2470,N_582,N_271);
or U2471 (N_2471,N_785,N_618);
or U2472 (N_2472,N_1023,N_420);
nand U2473 (N_2473,N_280,N_22);
nand U2474 (N_2474,N_594,N_1285);
nand U2475 (N_2475,N_778,N_307);
nand U2476 (N_2476,N_47,N_1062);
nor U2477 (N_2477,N_60,N_1190);
xor U2478 (N_2478,N_1267,N_46);
nand U2479 (N_2479,N_790,N_663);
and U2480 (N_2480,N_202,N_500);
nor U2481 (N_2481,N_150,N_747);
and U2482 (N_2482,N_1418,N_1427);
nand U2483 (N_2483,N_445,N_910);
nand U2484 (N_2484,N_1414,N_378);
or U2485 (N_2485,N_922,N_699);
and U2486 (N_2486,N_1224,N_523);
and U2487 (N_2487,N_41,N_174);
or U2488 (N_2488,N_1486,N_840);
nand U2489 (N_2489,N_940,N_1205);
nor U2490 (N_2490,N_965,N_837);
nand U2491 (N_2491,N_1478,N_292);
or U2492 (N_2492,N_804,N_1141);
or U2493 (N_2493,N_1057,N_838);
and U2494 (N_2494,N_95,N_67);
or U2495 (N_2495,N_1391,N_862);
or U2496 (N_2496,N_3,N_1133);
nand U2497 (N_2497,N_282,N_1016);
nand U2498 (N_2498,N_1418,N_1269);
and U2499 (N_2499,N_1196,N_523);
xnor U2500 (N_2500,N_1364,N_963);
and U2501 (N_2501,N_1427,N_1159);
nor U2502 (N_2502,N_328,N_132);
nor U2503 (N_2503,N_261,N_1335);
nand U2504 (N_2504,N_349,N_589);
nand U2505 (N_2505,N_152,N_1124);
or U2506 (N_2506,N_520,N_347);
or U2507 (N_2507,N_695,N_1141);
xnor U2508 (N_2508,N_1447,N_1468);
and U2509 (N_2509,N_986,N_745);
or U2510 (N_2510,N_889,N_544);
nand U2511 (N_2511,N_120,N_1340);
nor U2512 (N_2512,N_651,N_647);
and U2513 (N_2513,N_810,N_930);
nor U2514 (N_2514,N_574,N_457);
or U2515 (N_2515,N_1018,N_1375);
nor U2516 (N_2516,N_1161,N_139);
or U2517 (N_2517,N_923,N_963);
nand U2518 (N_2518,N_317,N_906);
nor U2519 (N_2519,N_205,N_415);
xnor U2520 (N_2520,N_1455,N_601);
nand U2521 (N_2521,N_745,N_29);
or U2522 (N_2522,N_1386,N_730);
and U2523 (N_2523,N_1137,N_29);
nand U2524 (N_2524,N_1449,N_61);
nand U2525 (N_2525,N_592,N_322);
nand U2526 (N_2526,N_1025,N_169);
xnor U2527 (N_2527,N_1459,N_530);
or U2528 (N_2528,N_319,N_1404);
or U2529 (N_2529,N_130,N_205);
nand U2530 (N_2530,N_335,N_1344);
nor U2531 (N_2531,N_1378,N_1415);
or U2532 (N_2532,N_1261,N_1252);
or U2533 (N_2533,N_302,N_240);
nor U2534 (N_2534,N_1114,N_1298);
or U2535 (N_2535,N_608,N_541);
nand U2536 (N_2536,N_600,N_335);
nand U2537 (N_2537,N_531,N_1028);
nor U2538 (N_2538,N_1337,N_213);
and U2539 (N_2539,N_518,N_1258);
and U2540 (N_2540,N_482,N_159);
nor U2541 (N_2541,N_847,N_730);
nor U2542 (N_2542,N_997,N_1055);
nor U2543 (N_2543,N_1051,N_1463);
nand U2544 (N_2544,N_1133,N_72);
or U2545 (N_2545,N_1228,N_130);
nand U2546 (N_2546,N_255,N_1417);
nor U2547 (N_2547,N_793,N_1291);
and U2548 (N_2548,N_784,N_536);
nor U2549 (N_2549,N_1164,N_951);
nand U2550 (N_2550,N_1235,N_1241);
and U2551 (N_2551,N_371,N_1091);
and U2552 (N_2552,N_1092,N_1482);
xnor U2553 (N_2553,N_1370,N_208);
nand U2554 (N_2554,N_537,N_284);
nand U2555 (N_2555,N_251,N_326);
and U2556 (N_2556,N_1432,N_890);
nor U2557 (N_2557,N_612,N_301);
nand U2558 (N_2558,N_683,N_226);
or U2559 (N_2559,N_162,N_928);
nand U2560 (N_2560,N_1367,N_139);
xnor U2561 (N_2561,N_538,N_83);
or U2562 (N_2562,N_1148,N_656);
or U2563 (N_2563,N_993,N_1010);
or U2564 (N_2564,N_1185,N_1458);
and U2565 (N_2565,N_512,N_490);
nand U2566 (N_2566,N_637,N_354);
and U2567 (N_2567,N_649,N_832);
and U2568 (N_2568,N_1248,N_1009);
nand U2569 (N_2569,N_897,N_1143);
and U2570 (N_2570,N_478,N_207);
nor U2571 (N_2571,N_37,N_756);
nor U2572 (N_2572,N_983,N_1280);
nor U2573 (N_2573,N_933,N_1164);
or U2574 (N_2574,N_701,N_1108);
and U2575 (N_2575,N_1426,N_503);
or U2576 (N_2576,N_810,N_1034);
nor U2577 (N_2577,N_235,N_633);
and U2578 (N_2578,N_148,N_1198);
nor U2579 (N_2579,N_377,N_626);
xnor U2580 (N_2580,N_1218,N_402);
xnor U2581 (N_2581,N_254,N_949);
and U2582 (N_2582,N_117,N_990);
nor U2583 (N_2583,N_180,N_1416);
nor U2584 (N_2584,N_422,N_171);
nor U2585 (N_2585,N_1158,N_1371);
nand U2586 (N_2586,N_83,N_229);
or U2587 (N_2587,N_661,N_913);
nand U2588 (N_2588,N_278,N_1081);
or U2589 (N_2589,N_687,N_1473);
and U2590 (N_2590,N_115,N_1393);
and U2591 (N_2591,N_1291,N_1380);
and U2592 (N_2592,N_326,N_473);
and U2593 (N_2593,N_1400,N_1493);
nand U2594 (N_2594,N_1003,N_676);
or U2595 (N_2595,N_627,N_540);
and U2596 (N_2596,N_1259,N_180);
nand U2597 (N_2597,N_994,N_1009);
or U2598 (N_2598,N_121,N_1166);
nor U2599 (N_2599,N_179,N_813);
nor U2600 (N_2600,N_400,N_1331);
nand U2601 (N_2601,N_990,N_1400);
nor U2602 (N_2602,N_37,N_1358);
nor U2603 (N_2603,N_1422,N_423);
nand U2604 (N_2604,N_1363,N_1160);
and U2605 (N_2605,N_685,N_289);
and U2606 (N_2606,N_1471,N_675);
nor U2607 (N_2607,N_899,N_138);
nand U2608 (N_2608,N_1462,N_21);
nand U2609 (N_2609,N_270,N_1234);
nor U2610 (N_2610,N_915,N_1229);
nor U2611 (N_2611,N_1411,N_414);
nand U2612 (N_2612,N_1246,N_897);
nor U2613 (N_2613,N_957,N_663);
nor U2614 (N_2614,N_86,N_1391);
and U2615 (N_2615,N_474,N_1148);
nand U2616 (N_2616,N_40,N_720);
or U2617 (N_2617,N_377,N_991);
nor U2618 (N_2618,N_161,N_1154);
or U2619 (N_2619,N_1140,N_805);
nor U2620 (N_2620,N_1138,N_28);
nor U2621 (N_2621,N_23,N_397);
or U2622 (N_2622,N_809,N_617);
nor U2623 (N_2623,N_1117,N_405);
and U2624 (N_2624,N_600,N_1188);
or U2625 (N_2625,N_683,N_1340);
or U2626 (N_2626,N_64,N_454);
and U2627 (N_2627,N_1380,N_1219);
and U2628 (N_2628,N_962,N_1491);
and U2629 (N_2629,N_119,N_84);
nor U2630 (N_2630,N_1005,N_190);
nor U2631 (N_2631,N_483,N_943);
and U2632 (N_2632,N_963,N_344);
or U2633 (N_2633,N_1135,N_747);
nor U2634 (N_2634,N_804,N_1044);
nor U2635 (N_2635,N_1131,N_171);
or U2636 (N_2636,N_980,N_927);
nand U2637 (N_2637,N_1040,N_505);
nor U2638 (N_2638,N_697,N_1188);
xnor U2639 (N_2639,N_182,N_1120);
or U2640 (N_2640,N_469,N_129);
or U2641 (N_2641,N_1480,N_1285);
or U2642 (N_2642,N_970,N_445);
or U2643 (N_2643,N_288,N_829);
nand U2644 (N_2644,N_947,N_831);
xnor U2645 (N_2645,N_1447,N_1240);
and U2646 (N_2646,N_1299,N_1455);
or U2647 (N_2647,N_1241,N_1335);
or U2648 (N_2648,N_460,N_1397);
nor U2649 (N_2649,N_155,N_52);
nand U2650 (N_2650,N_283,N_1369);
or U2651 (N_2651,N_698,N_1079);
xnor U2652 (N_2652,N_1369,N_826);
or U2653 (N_2653,N_1224,N_664);
nand U2654 (N_2654,N_70,N_176);
nor U2655 (N_2655,N_568,N_28);
xor U2656 (N_2656,N_675,N_1474);
nand U2657 (N_2657,N_1287,N_986);
nor U2658 (N_2658,N_459,N_677);
and U2659 (N_2659,N_1346,N_451);
and U2660 (N_2660,N_761,N_179);
and U2661 (N_2661,N_3,N_1006);
and U2662 (N_2662,N_1373,N_921);
nand U2663 (N_2663,N_56,N_835);
nor U2664 (N_2664,N_278,N_239);
xnor U2665 (N_2665,N_993,N_333);
nor U2666 (N_2666,N_714,N_1074);
and U2667 (N_2667,N_367,N_978);
or U2668 (N_2668,N_199,N_335);
and U2669 (N_2669,N_430,N_675);
or U2670 (N_2670,N_594,N_1398);
nand U2671 (N_2671,N_45,N_831);
nor U2672 (N_2672,N_43,N_370);
or U2673 (N_2673,N_964,N_798);
nor U2674 (N_2674,N_644,N_608);
or U2675 (N_2675,N_1046,N_45);
nand U2676 (N_2676,N_1495,N_630);
nand U2677 (N_2677,N_186,N_1313);
or U2678 (N_2678,N_13,N_1055);
and U2679 (N_2679,N_474,N_121);
nor U2680 (N_2680,N_1110,N_696);
and U2681 (N_2681,N_188,N_311);
or U2682 (N_2682,N_1286,N_658);
xnor U2683 (N_2683,N_483,N_1499);
nor U2684 (N_2684,N_1057,N_862);
or U2685 (N_2685,N_1294,N_1108);
nand U2686 (N_2686,N_1350,N_282);
nor U2687 (N_2687,N_742,N_1415);
and U2688 (N_2688,N_1158,N_340);
nand U2689 (N_2689,N_1075,N_88);
or U2690 (N_2690,N_271,N_1477);
nand U2691 (N_2691,N_427,N_1371);
or U2692 (N_2692,N_1189,N_377);
xor U2693 (N_2693,N_541,N_1160);
and U2694 (N_2694,N_114,N_382);
nand U2695 (N_2695,N_964,N_747);
nand U2696 (N_2696,N_591,N_785);
nand U2697 (N_2697,N_486,N_1199);
nand U2698 (N_2698,N_344,N_1192);
nor U2699 (N_2699,N_646,N_253);
and U2700 (N_2700,N_516,N_1001);
nor U2701 (N_2701,N_588,N_84);
or U2702 (N_2702,N_794,N_1395);
and U2703 (N_2703,N_864,N_505);
or U2704 (N_2704,N_267,N_1270);
and U2705 (N_2705,N_1403,N_430);
and U2706 (N_2706,N_1234,N_55);
nand U2707 (N_2707,N_1450,N_1241);
or U2708 (N_2708,N_1481,N_1009);
nand U2709 (N_2709,N_1001,N_1372);
xor U2710 (N_2710,N_1186,N_423);
nand U2711 (N_2711,N_1360,N_1405);
nand U2712 (N_2712,N_54,N_888);
or U2713 (N_2713,N_46,N_262);
nor U2714 (N_2714,N_637,N_215);
xnor U2715 (N_2715,N_488,N_1448);
nand U2716 (N_2716,N_1396,N_1268);
nor U2717 (N_2717,N_282,N_0);
and U2718 (N_2718,N_1359,N_739);
nand U2719 (N_2719,N_1169,N_1498);
nor U2720 (N_2720,N_600,N_475);
nand U2721 (N_2721,N_118,N_285);
nor U2722 (N_2722,N_1100,N_1264);
or U2723 (N_2723,N_135,N_269);
or U2724 (N_2724,N_679,N_1339);
xor U2725 (N_2725,N_246,N_881);
and U2726 (N_2726,N_1443,N_203);
nor U2727 (N_2727,N_565,N_28);
nor U2728 (N_2728,N_1258,N_1064);
xnor U2729 (N_2729,N_1309,N_279);
or U2730 (N_2730,N_445,N_945);
or U2731 (N_2731,N_917,N_1106);
nor U2732 (N_2732,N_476,N_1496);
or U2733 (N_2733,N_1374,N_1387);
nand U2734 (N_2734,N_609,N_1124);
and U2735 (N_2735,N_481,N_330);
or U2736 (N_2736,N_88,N_1062);
nor U2737 (N_2737,N_199,N_385);
nand U2738 (N_2738,N_731,N_739);
or U2739 (N_2739,N_1174,N_699);
and U2740 (N_2740,N_758,N_1251);
nand U2741 (N_2741,N_1156,N_616);
or U2742 (N_2742,N_650,N_1228);
or U2743 (N_2743,N_928,N_908);
and U2744 (N_2744,N_55,N_307);
or U2745 (N_2745,N_1469,N_869);
nand U2746 (N_2746,N_437,N_1391);
and U2747 (N_2747,N_970,N_25);
nand U2748 (N_2748,N_193,N_928);
or U2749 (N_2749,N_1185,N_1157);
nand U2750 (N_2750,N_551,N_77);
nor U2751 (N_2751,N_418,N_1377);
nor U2752 (N_2752,N_1084,N_1386);
nor U2753 (N_2753,N_1440,N_1328);
nand U2754 (N_2754,N_120,N_770);
xnor U2755 (N_2755,N_339,N_546);
nand U2756 (N_2756,N_531,N_1499);
or U2757 (N_2757,N_1031,N_1129);
or U2758 (N_2758,N_289,N_1162);
and U2759 (N_2759,N_1449,N_809);
and U2760 (N_2760,N_517,N_155);
xnor U2761 (N_2761,N_1283,N_1111);
or U2762 (N_2762,N_503,N_189);
and U2763 (N_2763,N_1389,N_788);
nand U2764 (N_2764,N_546,N_813);
xnor U2765 (N_2765,N_723,N_511);
or U2766 (N_2766,N_1115,N_289);
nand U2767 (N_2767,N_770,N_148);
nor U2768 (N_2768,N_122,N_571);
nand U2769 (N_2769,N_482,N_1213);
or U2770 (N_2770,N_176,N_26);
nand U2771 (N_2771,N_217,N_948);
xnor U2772 (N_2772,N_31,N_1012);
xor U2773 (N_2773,N_1401,N_1220);
or U2774 (N_2774,N_891,N_186);
nor U2775 (N_2775,N_1160,N_1155);
nor U2776 (N_2776,N_387,N_124);
and U2777 (N_2777,N_430,N_1235);
and U2778 (N_2778,N_960,N_660);
xor U2779 (N_2779,N_652,N_658);
nand U2780 (N_2780,N_952,N_136);
and U2781 (N_2781,N_1453,N_856);
and U2782 (N_2782,N_905,N_998);
xnor U2783 (N_2783,N_1032,N_100);
and U2784 (N_2784,N_402,N_719);
nor U2785 (N_2785,N_586,N_670);
xor U2786 (N_2786,N_491,N_1343);
nor U2787 (N_2787,N_1132,N_1078);
nor U2788 (N_2788,N_808,N_492);
and U2789 (N_2789,N_1377,N_958);
nand U2790 (N_2790,N_1393,N_412);
and U2791 (N_2791,N_102,N_1481);
nand U2792 (N_2792,N_652,N_1119);
nand U2793 (N_2793,N_635,N_786);
or U2794 (N_2794,N_757,N_1433);
nand U2795 (N_2795,N_622,N_1279);
or U2796 (N_2796,N_877,N_1278);
nor U2797 (N_2797,N_288,N_1276);
nor U2798 (N_2798,N_1271,N_57);
nand U2799 (N_2799,N_399,N_1359);
or U2800 (N_2800,N_1476,N_537);
and U2801 (N_2801,N_1162,N_1025);
and U2802 (N_2802,N_629,N_1322);
or U2803 (N_2803,N_337,N_420);
and U2804 (N_2804,N_835,N_544);
and U2805 (N_2805,N_279,N_754);
or U2806 (N_2806,N_391,N_1094);
nor U2807 (N_2807,N_1137,N_769);
nor U2808 (N_2808,N_278,N_291);
or U2809 (N_2809,N_399,N_1107);
nor U2810 (N_2810,N_1059,N_1484);
nor U2811 (N_2811,N_153,N_1209);
xor U2812 (N_2812,N_1090,N_1201);
xor U2813 (N_2813,N_447,N_20);
xor U2814 (N_2814,N_991,N_138);
and U2815 (N_2815,N_1432,N_824);
nor U2816 (N_2816,N_869,N_693);
or U2817 (N_2817,N_1281,N_975);
nor U2818 (N_2818,N_1022,N_247);
or U2819 (N_2819,N_444,N_1251);
xnor U2820 (N_2820,N_744,N_1023);
and U2821 (N_2821,N_903,N_883);
nor U2822 (N_2822,N_806,N_982);
nand U2823 (N_2823,N_1105,N_1169);
or U2824 (N_2824,N_290,N_1254);
and U2825 (N_2825,N_466,N_562);
or U2826 (N_2826,N_288,N_96);
nor U2827 (N_2827,N_673,N_441);
or U2828 (N_2828,N_750,N_1364);
or U2829 (N_2829,N_111,N_691);
nor U2830 (N_2830,N_817,N_662);
nand U2831 (N_2831,N_1494,N_1313);
nor U2832 (N_2832,N_1355,N_54);
or U2833 (N_2833,N_1422,N_208);
or U2834 (N_2834,N_1489,N_893);
nand U2835 (N_2835,N_820,N_1043);
or U2836 (N_2836,N_681,N_945);
and U2837 (N_2837,N_1161,N_1269);
nand U2838 (N_2838,N_387,N_441);
or U2839 (N_2839,N_1318,N_168);
or U2840 (N_2840,N_41,N_1140);
or U2841 (N_2841,N_1404,N_560);
nor U2842 (N_2842,N_1069,N_919);
or U2843 (N_2843,N_406,N_1202);
xor U2844 (N_2844,N_1465,N_895);
or U2845 (N_2845,N_1454,N_651);
xnor U2846 (N_2846,N_1166,N_157);
and U2847 (N_2847,N_406,N_122);
nor U2848 (N_2848,N_427,N_1043);
or U2849 (N_2849,N_1047,N_1351);
xnor U2850 (N_2850,N_249,N_1184);
nor U2851 (N_2851,N_439,N_1082);
or U2852 (N_2852,N_162,N_487);
xor U2853 (N_2853,N_1300,N_506);
or U2854 (N_2854,N_1137,N_358);
or U2855 (N_2855,N_826,N_554);
xnor U2856 (N_2856,N_940,N_1013);
nand U2857 (N_2857,N_555,N_521);
nor U2858 (N_2858,N_161,N_735);
and U2859 (N_2859,N_557,N_5);
nand U2860 (N_2860,N_855,N_1041);
xor U2861 (N_2861,N_1099,N_763);
nor U2862 (N_2862,N_125,N_919);
nand U2863 (N_2863,N_747,N_251);
or U2864 (N_2864,N_1224,N_1216);
nand U2865 (N_2865,N_126,N_947);
or U2866 (N_2866,N_1394,N_1113);
nor U2867 (N_2867,N_1050,N_340);
nand U2868 (N_2868,N_214,N_896);
or U2869 (N_2869,N_419,N_1052);
nor U2870 (N_2870,N_539,N_966);
xor U2871 (N_2871,N_444,N_70);
nand U2872 (N_2872,N_179,N_668);
nor U2873 (N_2873,N_83,N_1007);
nand U2874 (N_2874,N_953,N_58);
or U2875 (N_2875,N_127,N_334);
or U2876 (N_2876,N_893,N_1207);
and U2877 (N_2877,N_1085,N_146);
nor U2878 (N_2878,N_242,N_884);
xor U2879 (N_2879,N_1420,N_426);
nor U2880 (N_2880,N_555,N_1456);
nand U2881 (N_2881,N_579,N_1200);
and U2882 (N_2882,N_734,N_1387);
and U2883 (N_2883,N_928,N_774);
or U2884 (N_2884,N_998,N_43);
or U2885 (N_2885,N_1459,N_637);
nand U2886 (N_2886,N_518,N_301);
nor U2887 (N_2887,N_552,N_1085);
nor U2888 (N_2888,N_975,N_783);
and U2889 (N_2889,N_1494,N_255);
and U2890 (N_2890,N_539,N_1324);
or U2891 (N_2891,N_1231,N_1217);
nor U2892 (N_2892,N_207,N_1293);
and U2893 (N_2893,N_521,N_1311);
or U2894 (N_2894,N_1338,N_411);
and U2895 (N_2895,N_594,N_1348);
nand U2896 (N_2896,N_1222,N_267);
and U2897 (N_2897,N_104,N_1358);
or U2898 (N_2898,N_330,N_1313);
nor U2899 (N_2899,N_164,N_1463);
xnor U2900 (N_2900,N_1090,N_894);
nor U2901 (N_2901,N_892,N_1108);
nor U2902 (N_2902,N_132,N_179);
nand U2903 (N_2903,N_1040,N_1118);
nand U2904 (N_2904,N_1401,N_1290);
xor U2905 (N_2905,N_455,N_600);
or U2906 (N_2906,N_861,N_1236);
nand U2907 (N_2907,N_563,N_336);
nand U2908 (N_2908,N_1291,N_1372);
xor U2909 (N_2909,N_281,N_777);
and U2910 (N_2910,N_1425,N_37);
nor U2911 (N_2911,N_765,N_1203);
nand U2912 (N_2912,N_269,N_1068);
or U2913 (N_2913,N_1461,N_1029);
and U2914 (N_2914,N_566,N_488);
nand U2915 (N_2915,N_684,N_378);
nor U2916 (N_2916,N_792,N_1248);
nand U2917 (N_2917,N_110,N_150);
or U2918 (N_2918,N_933,N_309);
and U2919 (N_2919,N_1347,N_955);
and U2920 (N_2920,N_458,N_606);
or U2921 (N_2921,N_352,N_680);
or U2922 (N_2922,N_328,N_15);
and U2923 (N_2923,N_75,N_1387);
nor U2924 (N_2924,N_604,N_944);
nor U2925 (N_2925,N_1313,N_1092);
nor U2926 (N_2926,N_525,N_1304);
or U2927 (N_2927,N_1242,N_1440);
or U2928 (N_2928,N_980,N_425);
xnor U2929 (N_2929,N_324,N_1138);
nand U2930 (N_2930,N_115,N_1389);
nand U2931 (N_2931,N_1260,N_256);
or U2932 (N_2932,N_697,N_1064);
and U2933 (N_2933,N_324,N_720);
nor U2934 (N_2934,N_293,N_386);
nand U2935 (N_2935,N_833,N_672);
and U2936 (N_2936,N_619,N_1378);
or U2937 (N_2937,N_367,N_147);
nor U2938 (N_2938,N_1052,N_739);
or U2939 (N_2939,N_708,N_519);
or U2940 (N_2940,N_1452,N_314);
and U2941 (N_2941,N_989,N_939);
nor U2942 (N_2942,N_457,N_993);
or U2943 (N_2943,N_65,N_40);
or U2944 (N_2944,N_1326,N_1355);
nand U2945 (N_2945,N_659,N_411);
or U2946 (N_2946,N_333,N_1124);
or U2947 (N_2947,N_225,N_925);
or U2948 (N_2948,N_47,N_537);
and U2949 (N_2949,N_119,N_1080);
nor U2950 (N_2950,N_1159,N_602);
xor U2951 (N_2951,N_1068,N_903);
nand U2952 (N_2952,N_650,N_1317);
or U2953 (N_2953,N_297,N_282);
xnor U2954 (N_2954,N_849,N_901);
nor U2955 (N_2955,N_1061,N_874);
or U2956 (N_2956,N_1311,N_377);
nand U2957 (N_2957,N_991,N_89);
nand U2958 (N_2958,N_1417,N_1374);
or U2959 (N_2959,N_1369,N_204);
or U2960 (N_2960,N_867,N_96);
or U2961 (N_2961,N_366,N_395);
nor U2962 (N_2962,N_1251,N_1283);
and U2963 (N_2963,N_139,N_537);
nor U2964 (N_2964,N_747,N_1092);
nand U2965 (N_2965,N_92,N_594);
xor U2966 (N_2966,N_699,N_483);
or U2967 (N_2967,N_89,N_1464);
xnor U2968 (N_2968,N_699,N_1176);
xnor U2969 (N_2969,N_231,N_1196);
nand U2970 (N_2970,N_972,N_1217);
nand U2971 (N_2971,N_1195,N_295);
nand U2972 (N_2972,N_948,N_681);
nor U2973 (N_2973,N_1335,N_1404);
or U2974 (N_2974,N_625,N_988);
or U2975 (N_2975,N_1472,N_1128);
nand U2976 (N_2976,N_316,N_225);
or U2977 (N_2977,N_335,N_153);
and U2978 (N_2978,N_1256,N_107);
nand U2979 (N_2979,N_290,N_1344);
and U2980 (N_2980,N_161,N_938);
nor U2981 (N_2981,N_1116,N_1207);
nor U2982 (N_2982,N_701,N_959);
and U2983 (N_2983,N_252,N_965);
nor U2984 (N_2984,N_953,N_794);
xnor U2985 (N_2985,N_1170,N_8);
nand U2986 (N_2986,N_537,N_857);
nor U2987 (N_2987,N_205,N_1137);
nor U2988 (N_2988,N_248,N_1172);
or U2989 (N_2989,N_558,N_1115);
xnor U2990 (N_2990,N_170,N_892);
or U2991 (N_2991,N_1487,N_693);
or U2992 (N_2992,N_350,N_1401);
nor U2993 (N_2993,N_619,N_195);
nand U2994 (N_2994,N_837,N_1399);
and U2995 (N_2995,N_224,N_263);
nor U2996 (N_2996,N_1451,N_1218);
nand U2997 (N_2997,N_899,N_288);
and U2998 (N_2998,N_360,N_828);
or U2999 (N_2999,N_322,N_173);
nor U3000 (N_3000,N_1847,N_1522);
and U3001 (N_3001,N_2532,N_1788);
and U3002 (N_3002,N_2941,N_1911);
nand U3003 (N_3003,N_2015,N_2714);
nand U3004 (N_3004,N_2043,N_1602);
and U3005 (N_3005,N_1883,N_2291);
nand U3006 (N_3006,N_2343,N_2956);
nand U3007 (N_3007,N_1698,N_2873);
nand U3008 (N_3008,N_1694,N_1999);
xnor U3009 (N_3009,N_2233,N_1562);
nand U3010 (N_3010,N_2886,N_1637);
or U3011 (N_3011,N_1786,N_1611);
nand U3012 (N_3012,N_2289,N_2143);
and U3013 (N_3013,N_2960,N_2439);
nand U3014 (N_3014,N_2634,N_2609);
or U3015 (N_3015,N_2925,N_2686);
and U3016 (N_3016,N_2154,N_2536);
and U3017 (N_3017,N_2160,N_1666);
and U3018 (N_3018,N_2818,N_1679);
nand U3019 (N_3019,N_2494,N_2318);
and U3020 (N_3020,N_2017,N_1897);
nand U3021 (N_3021,N_2903,N_2278);
or U3022 (N_3022,N_2817,N_2202);
nand U3023 (N_3023,N_2052,N_2682);
and U3024 (N_3024,N_2210,N_1887);
nand U3025 (N_3025,N_2119,N_1735);
or U3026 (N_3026,N_2431,N_1646);
or U3027 (N_3027,N_2179,N_2685);
and U3028 (N_3028,N_1641,N_2276);
or U3029 (N_3029,N_2997,N_2116);
nor U3030 (N_3030,N_1592,N_2475);
xor U3031 (N_3031,N_2074,N_2470);
nor U3032 (N_3032,N_2772,N_2471);
or U3033 (N_3033,N_1850,N_1524);
xnor U3034 (N_3034,N_2309,N_2665);
or U3035 (N_3035,N_2277,N_1546);
or U3036 (N_3036,N_2527,N_1856);
and U3037 (N_3037,N_1745,N_2888);
xor U3038 (N_3038,N_2385,N_2987);
and U3039 (N_3039,N_2497,N_2166);
and U3040 (N_3040,N_2780,N_2207);
nor U3041 (N_3041,N_1980,N_1722);
or U3042 (N_3042,N_1992,N_2940);
nand U3043 (N_3043,N_1851,N_2484);
nand U3044 (N_3044,N_1998,N_2461);
and U3045 (N_3045,N_2300,N_1908);
nand U3046 (N_3046,N_1560,N_1907);
and U3047 (N_3047,N_1711,N_1793);
or U3048 (N_3048,N_2259,N_2587);
nor U3049 (N_3049,N_2547,N_1703);
nor U3050 (N_3050,N_1542,N_2186);
xor U3051 (N_3051,N_2046,N_2787);
or U3052 (N_3052,N_1586,N_2598);
nand U3053 (N_3053,N_1949,N_2190);
xnor U3054 (N_3054,N_1924,N_2379);
nor U3055 (N_3055,N_2738,N_2007);
nor U3056 (N_3056,N_2813,N_2709);
xnor U3057 (N_3057,N_2773,N_2408);
nand U3058 (N_3058,N_1530,N_1531);
nand U3059 (N_3059,N_1800,N_1579);
nor U3060 (N_3060,N_2150,N_2324);
nand U3061 (N_3061,N_1664,N_1521);
or U3062 (N_3062,N_1649,N_2097);
nor U3063 (N_3063,N_2393,N_2212);
nand U3064 (N_3064,N_1700,N_2244);
or U3065 (N_3065,N_2827,N_2713);
nand U3066 (N_3066,N_2171,N_2495);
nor U3067 (N_3067,N_2287,N_2693);
xnor U3068 (N_3068,N_2863,N_2355);
nand U3069 (N_3069,N_2263,N_1770);
or U3070 (N_3070,N_2703,N_1625);
and U3071 (N_3071,N_1889,N_2783);
nand U3072 (N_3072,N_1619,N_2825);
nor U3073 (N_3073,N_2938,N_2853);
xnor U3074 (N_3074,N_2563,N_2224);
nor U3075 (N_3075,N_2763,N_1598);
or U3076 (N_3076,N_2778,N_2336);
or U3077 (N_3077,N_2782,N_2988);
and U3078 (N_3078,N_2025,N_2103);
and U3079 (N_3079,N_2552,N_2591);
xor U3080 (N_3080,N_2402,N_2188);
nand U3081 (N_3081,N_1667,N_1507);
nand U3082 (N_3082,N_2835,N_2423);
and U3083 (N_3083,N_2846,N_1724);
nand U3084 (N_3084,N_2877,N_2032);
nor U3085 (N_3085,N_2513,N_2478);
or U3086 (N_3086,N_2984,N_2267);
nor U3087 (N_3087,N_2255,N_2468);
nor U3088 (N_3088,N_2584,N_2930);
and U3089 (N_3089,N_2248,N_2361);
nand U3090 (N_3090,N_1600,N_2070);
nor U3091 (N_3091,N_2640,N_2285);
xnor U3092 (N_3092,N_1970,N_2317);
or U3093 (N_3093,N_1606,N_2882);
and U3094 (N_3094,N_1725,N_2392);
and U3095 (N_3095,N_2936,N_2983);
xor U3096 (N_3096,N_2681,N_2365);
or U3097 (N_3097,N_2127,N_2362);
nor U3098 (N_3098,N_2549,N_2384);
and U3099 (N_3099,N_1639,N_2574);
and U3100 (N_3100,N_1953,N_1769);
nor U3101 (N_3101,N_2095,N_2595);
and U3102 (N_3102,N_2252,N_1795);
nand U3103 (N_3103,N_1842,N_2546);
or U3104 (N_3104,N_2991,N_2679);
nor U3105 (N_3105,N_1987,N_2348);
or U3106 (N_3106,N_2486,N_1849);
nor U3107 (N_3107,N_2535,N_1766);
or U3108 (N_3108,N_2001,N_2861);
nand U3109 (N_3109,N_1994,N_2102);
or U3110 (N_3110,N_2680,N_1683);
and U3111 (N_3111,N_2978,N_1653);
nand U3112 (N_3112,N_1807,N_2718);
nand U3113 (N_3113,N_2064,N_1816);
nor U3114 (N_3114,N_1628,N_2373);
nand U3115 (N_3115,N_2342,N_2487);
and U3116 (N_3116,N_1506,N_2316);
nor U3117 (N_3117,N_2899,N_2406);
nor U3118 (N_3118,N_2322,N_1523);
and U3119 (N_3119,N_2488,N_2559);
and U3120 (N_3120,N_2919,N_1848);
or U3121 (N_3121,N_2613,N_1758);
nand U3122 (N_3122,N_1525,N_1968);
nor U3123 (N_3123,N_1729,N_1867);
nand U3124 (N_3124,N_2623,N_2208);
and U3125 (N_3125,N_2751,N_1601);
nand U3126 (N_3126,N_2451,N_1737);
nor U3127 (N_3127,N_1741,N_1659);
or U3128 (N_3128,N_1642,N_1633);
and U3129 (N_3129,N_1686,N_2989);
or U3130 (N_3130,N_2672,N_2193);
and U3131 (N_3131,N_2400,N_1608);
and U3132 (N_3132,N_1803,N_1544);
xor U3133 (N_3133,N_2908,N_1811);
or U3134 (N_3134,N_1916,N_2108);
nor U3135 (N_3135,N_2800,N_2805);
and U3136 (N_3136,N_2555,N_2125);
and U3137 (N_3137,N_2000,N_1858);
nand U3138 (N_3138,N_2652,N_2645);
and U3139 (N_3139,N_2183,N_2567);
and U3140 (N_3140,N_2199,N_2878);
and U3141 (N_3141,N_1767,N_1690);
xor U3142 (N_3142,N_2363,N_1976);
and U3143 (N_3143,N_2616,N_2689);
nor U3144 (N_3144,N_2876,N_1750);
nor U3145 (N_3145,N_2617,N_1549);
nand U3146 (N_3146,N_1901,N_2034);
xnor U3147 (N_3147,N_1699,N_2670);
or U3148 (N_3148,N_1707,N_1840);
and U3149 (N_3149,N_1860,N_2701);
or U3150 (N_3150,N_2858,N_2949);
nand U3151 (N_3151,N_2957,N_1734);
or U3152 (N_3152,N_1588,N_2909);
nor U3153 (N_3153,N_2889,N_2515);
nor U3154 (N_3154,N_2238,N_1863);
xor U3155 (N_3155,N_1581,N_2796);
nor U3156 (N_3156,N_2972,N_2469);
nor U3157 (N_3157,N_2509,N_2086);
nor U3158 (N_3158,N_2091,N_1555);
nand U3159 (N_3159,N_1961,N_1710);
and U3160 (N_3160,N_2364,N_2082);
and U3161 (N_3161,N_2297,N_2409);
and U3162 (N_3162,N_2051,N_1558);
nor U3163 (N_3163,N_1797,N_2624);
or U3164 (N_3164,N_1557,N_1760);
and U3165 (N_3165,N_1564,N_2668);
and U3166 (N_3166,N_2758,N_2955);
nand U3167 (N_3167,N_2979,N_2743);
nor U3168 (N_3168,N_2204,N_2347);
and U3169 (N_3169,N_2662,N_1792);
or U3170 (N_3170,N_1640,N_2162);
nand U3171 (N_3171,N_2820,N_2896);
nor U3172 (N_3172,N_2885,N_2288);
nand U3173 (N_3173,N_1938,N_2739);
nor U3174 (N_3174,N_2059,N_2504);
nor U3175 (N_3175,N_1539,N_2586);
or U3176 (N_3176,N_2554,N_2917);
nand U3177 (N_3177,N_1898,N_1772);
nor U3178 (N_3178,N_2697,N_2657);
nand U3179 (N_3179,N_1744,N_2503);
or U3180 (N_3180,N_1708,N_2575);
nor U3181 (N_3181,N_2664,N_2764);
nand U3182 (N_3182,N_2446,N_2031);
or U3183 (N_3183,N_2087,N_2635);
nor U3184 (N_3184,N_2435,N_2325);
and U3185 (N_3185,N_1752,N_2447);
or U3186 (N_3186,N_1516,N_1895);
or U3187 (N_3187,N_2410,N_2880);
nor U3188 (N_3188,N_2083,N_1775);
and U3189 (N_3189,N_2173,N_2118);
nand U3190 (N_3190,N_2893,N_2557);
and U3191 (N_3191,N_1958,N_2864);
nand U3192 (N_3192,N_2418,N_1782);
or U3193 (N_3193,N_2496,N_1829);
and U3194 (N_3194,N_1723,N_1885);
and U3195 (N_3195,N_2137,N_2067);
xnor U3196 (N_3196,N_1721,N_2310);
nand U3197 (N_3197,N_1991,N_2705);
nor U3198 (N_3198,N_1955,N_2808);
nand U3199 (N_3199,N_2875,N_2594);
nand U3200 (N_3200,N_2601,N_2819);
or U3201 (N_3201,N_1975,N_2089);
nand U3202 (N_3202,N_1764,N_2840);
nand U3203 (N_3203,N_1905,N_2742);
or U3204 (N_3204,N_2740,N_1651);
nor U3205 (N_3205,N_2790,N_2420);
nor U3206 (N_3206,N_2073,N_2553);
and U3207 (N_3207,N_2455,N_2982);
nand U3208 (N_3208,N_2793,N_1878);
or U3209 (N_3209,N_1691,N_1809);
or U3210 (N_3210,N_2352,N_2019);
and U3211 (N_3211,N_2890,N_1616);
xnor U3212 (N_3212,N_2228,N_1550);
or U3213 (N_3213,N_2803,N_2340);
xor U3214 (N_3214,N_2200,N_2101);
nand U3215 (N_3215,N_2229,N_1603);
or U3216 (N_3216,N_2237,N_2608);
nor U3217 (N_3217,N_2964,N_2430);
or U3218 (N_3218,N_1817,N_1892);
and U3219 (N_3219,N_1977,N_2182);
or U3220 (N_3220,N_2528,N_2523);
xor U3221 (N_3221,N_2467,N_1922);
nand U3222 (N_3222,N_2247,N_2192);
or U3223 (N_3223,N_2156,N_2050);
nor U3224 (N_3224,N_2512,N_2194);
or U3225 (N_3225,N_2320,N_2198);
nor U3226 (N_3226,N_2394,N_1584);
and U3227 (N_3227,N_2265,N_2090);
or U3228 (N_3228,N_2438,N_2401);
nand U3229 (N_3229,N_1678,N_1747);
nand U3230 (N_3230,N_2622,N_1835);
nand U3231 (N_3231,N_1548,N_2966);
and U3232 (N_3232,N_1939,N_2568);
nand U3233 (N_3233,N_2845,N_2592);
and U3234 (N_3234,N_2066,N_1573);
and U3235 (N_3235,N_1661,N_2053);
xnor U3236 (N_3236,N_1915,N_1877);
or U3237 (N_3237,N_1853,N_2939);
and U3238 (N_3238,N_2958,N_1732);
nand U3239 (N_3239,N_2830,N_2454);
nand U3240 (N_3240,N_1773,N_2049);
nor U3241 (N_3241,N_1778,N_1652);
and U3242 (N_3242,N_2619,N_2234);
or U3243 (N_3243,N_1636,N_2892);
and U3244 (N_3244,N_2826,N_2728);
and U3245 (N_3245,N_1746,N_2257);
xor U3246 (N_3246,N_2434,N_2735);
nor U3247 (N_3247,N_2950,N_1866);
or U3248 (N_3248,N_2163,N_2596);
nand U3249 (N_3249,N_2719,N_2881);
nor U3250 (N_3250,N_1909,N_1692);
nor U3251 (N_3251,N_1810,N_1605);
nor U3252 (N_3252,N_2387,N_2344);
and U3253 (N_3253,N_2629,N_2147);
nor U3254 (N_3254,N_1820,N_2136);
and U3255 (N_3255,N_1796,N_2823);
or U3256 (N_3256,N_1621,N_1875);
nor U3257 (N_3257,N_1526,N_1701);
or U3258 (N_3258,N_2437,N_2674);
nor U3259 (N_3259,N_1529,N_2804);
xor U3260 (N_3260,N_2610,N_2115);
and U3261 (N_3261,N_1940,N_1804);
or U3262 (N_3262,N_2832,N_1505);
nor U3263 (N_3263,N_1805,N_2911);
nand U3264 (N_3264,N_1501,N_2303);
or U3265 (N_3265,N_2834,N_2542);
and U3266 (N_3266,N_2605,N_2766);
and U3267 (N_3267,N_2928,N_2712);
nor U3268 (N_3268,N_2904,N_2537);
nand U3269 (N_3269,N_1936,N_2124);
and U3270 (N_3270,N_2253,N_2789);
nand U3271 (N_3271,N_2531,N_2391);
and U3272 (N_3272,N_2060,N_2745);
nand U3273 (N_3273,N_2589,N_2040);
xor U3274 (N_3274,N_2453,N_2543);
and U3275 (N_3275,N_2684,N_2837);
nand U3276 (N_3276,N_2581,N_2213);
nor U3277 (N_3277,N_2692,N_2628);
nand U3278 (N_3278,N_2583,N_2510);
nand U3279 (N_3279,N_1715,N_1645);
xor U3280 (N_3280,N_2599,N_1944);
and U3281 (N_3281,N_2891,N_2521);
nor U3282 (N_3282,N_2359,N_2929);
nor U3283 (N_3283,N_2395,N_2544);
nor U3284 (N_3284,N_2273,N_2883);
or U3285 (N_3285,N_2472,N_1827);
nand U3286 (N_3286,N_2900,N_1914);
or U3287 (N_3287,N_2759,N_2731);
nand U3288 (N_3288,N_1671,N_1534);
and U3289 (N_3289,N_1631,N_2164);
and U3290 (N_3290,N_1943,N_2653);
nor U3291 (N_3291,N_2870,N_1731);
xor U3292 (N_3292,N_1563,N_1527);
and U3293 (N_3293,N_1569,N_1865);
or U3294 (N_3294,N_2525,N_1771);
or U3295 (N_3295,N_1882,N_1966);
or U3296 (N_3296,N_1837,N_2573);
nor U3297 (N_3297,N_2305,N_1906);
nand U3298 (N_3298,N_1668,N_1973);
nand U3299 (N_3299,N_2346,N_2639);
nor U3300 (N_3300,N_1647,N_2506);
or U3301 (N_3301,N_1728,N_2068);
or U3302 (N_3302,N_2872,N_2088);
or U3303 (N_3303,N_2129,N_2396);
xor U3304 (N_3304,N_2480,N_2403);
and U3305 (N_3305,N_1540,N_2534);
nor U3306 (N_3306,N_2270,N_2345);
nand U3307 (N_3307,N_2448,N_1547);
and U3308 (N_3308,N_2571,N_2242);
nor U3309 (N_3309,N_1845,N_2153);
nor U3310 (N_3310,N_2860,N_1517);
nor U3311 (N_3311,N_2360,N_2254);
or U3312 (N_3312,N_2945,N_1684);
nand U3313 (N_3313,N_2986,N_2155);
nand U3314 (N_3314,N_2113,N_2367);
xnor U3315 (N_3315,N_1623,N_1918);
nor U3316 (N_3316,N_2181,N_1585);
nand U3317 (N_3317,N_1541,N_2579);
and U3318 (N_3318,N_1514,N_1969);
nand U3319 (N_3319,N_2168,N_2727);
or U3320 (N_3320,N_2501,N_2459);
nand U3321 (N_3321,N_2195,N_1819);
nor U3322 (N_3322,N_1808,N_2120);
xnor U3323 (N_3323,N_2849,N_1537);
nand U3324 (N_3324,N_2282,N_2219);
nand U3325 (N_3325,N_2831,N_2848);
nor U3326 (N_3326,N_2934,N_2868);
nor U3327 (N_3327,N_1655,N_1886);
nor U3328 (N_3328,N_2283,N_2098);
nand U3329 (N_3329,N_2874,N_1689);
and U3330 (N_3330,N_2056,N_1676);
nand U3331 (N_3331,N_2752,N_2272);
xnor U3332 (N_3332,N_2216,N_2676);
nor U3333 (N_3333,N_1902,N_2126);
or U3334 (N_3334,N_2489,N_1654);
nor U3335 (N_3335,N_2922,N_2829);
or U3336 (N_3336,N_1660,N_2667);
or U3337 (N_3337,N_1791,N_1595);
nor U3338 (N_3338,N_2785,N_2262);
nor U3339 (N_3339,N_2951,N_2611);
xnor U3340 (N_3340,N_1995,N_2654);
nand U3341 (N_3341,N_2123,N_2167);
xor U3342 (N_3342,N_2836,N_2398);
xnor U3343 (N_3343,N_2243,N_2669);
nand U3344 (N_3344,N_2944,N_2474);
nor U3345 (N_3345,N_2433,N_2184);
nand U3346 (N_3346,N_2057,N_1846);
or U3347 (N_3347,N_2797,N_1594);
or U3348 (N_3348,N_2811,N_2351);
nor U3349 (N_3349,N_2963,N_2937);
xor U3350 (N_3350,N_2152,N_2197);
and U3351 (N_3351,N_2588,N_2769);
and U3352 (N_3352,N_1511,N_2750);
and U3353 (N_3353,N_2071,N_1823);
nor U3354 (N_3354,N_2240,N_2079);
and U3355 (N_3355,N_2741,N_2476);
nor U3356 (N_3356,N_2295,N_2096);
nor U3357 (N_3357,N_2491,N_1757);
nor U3358 (N_3358,N_1777,N_1774);
nand U3359 (N_3359,N_2341,N_2948);
or U3360 (N_3360,N_2913,N_2801);
and U3361 (N_3361,N_2795,N_1518);
nand U3362 (N_3362,N_2970,N_2161);
and U3363 (N_3363,N_2286,N_2816);
nor U3364 (N_3364,N_2992,N_1825);
nand U3365 (N_3365,N_2648,N_1861);
or U3366 (N_3366,N_2756,N_2481);
nor U3367 (N_3367,N_2696,N_2560);
or U3368 (N_3368,N_2323,N_2335);
nor U3369 (N_3369,N_1612,N_2132);
nand U3370 (N_3370,N_2421,N_2388);
or U3371 (N_3371,N_2349,N_1702);
and U3372 (N_3372,N_2220,N_2405);
nor U3373 (N_3373,N_2256,N_1515);
nand U3374 (N_3374,N_2176,N_2814);
nand U3375 (N_3375,N_2416,N_1552);
nand U3376 (N_3376,N_2702,N_1519);
nor U3377 (N_3377,N_2517,N_1959);
nand U3378 (N_3378,N_2290,N_2027);
nand U3379 (N_3379,N_2570,N_2426);
and U3380 (N_3380,N_2029,N_1838);
nand U3381 (N_3381,N_1751,N_1967);
nand U3382 (N_3382,N_1704,N_1535);
and U3383 (N_3383,N_1556,N_1567);
xnor U3384 (N_3384,N_1665,N_2376);
or U3385 (N_3385,N_2687,N_2671);
and U3386 (N_3386,N_2326,N_2673);
and U3387 (N_3387,N_2650,N_1787);
nor U3388 (N_3388,N_2140,N_2897);
or U3389 (N_3389,N_2799,N_2169);
and U3390 (N_3390,N_2085,N_2768);
nand U3391 (N_3391,N_2294,N_2920);
xnor U3392 (N_3392,N_1806,N_2022);
and U3393 (N_3393,N_1719,N_1925);
and U3394 (N_3394,N_1626,N_2636);
nor U3395 (N_3395,N_2463,N_1785);
or U3396 (N_3396,N_2980,N_2754);
and U3397 (N_3397,N_2660,N_1587);
nand U3398 (N_3398,N_2422,N_2319);
or U3399 (N_3399,N_1833,N_2815);
xnor U3400 (N_3400,N_1609,N_2500);
nor U3401 (N_3401,N_2170,N_2946);
and U3402 (N_3402,N_2397,N_1945);
nand U3403 (N_3403,N_1952,N_2646);
and U3404 (N_3404,N_2602,N_2806);
or U3405 (N_3405,N_1801,N_1635);
and U3406 (N_3406,N_2037,N_2618);
or U3407 (N_3407,N_2969,N_1972);
nand U3408 (N_3408,N_2901,N_1927);
and U3409 (N_3409,N_2869,N_1716);
nor U3410 (N_3410,N_2716,N_2914);
or U3411 (N_3411,N_2466,N_2918);
or U3412 (N_3412,N_2038,N_1739);
and U3413 (N_3413,N_1599,N_1630);
xor U3414 (N_3414,N_1510,N_2732);
nor U3415 (N_3415,N_2514,N_2462);
nand U3416 (N_3416,N_2600,N_2802);
nand U3417 (N_3417,N_2479,N_2271);
and U3418 (N_3418,N_2729,N_2710);
nand U3419 (N_3419,N_2569,N_2722);
or U3420 (N_3420,N_2378,N_2281);
nor U3421 (N_3421,N_1934,N_2312);
and U3422 (N_3422,N_2268,N_2299);
or U3423 (N_3423,N_2093,N_1921);
nor U3424 (N_3424,N_2753,N_2786);
xor U3425 (N_3425,N_2998,N_2308);
and U3426 (N_3426,N_2538,N_2798);
and U3427 (N_3427,N_2971,N_1784);
nand U3428 (N_3428,N_2075,N_1578);
nor U3429 (N_3429,N_1618,N_1673);
nor U3430 (N_3430,N_2044,N_2809);
and U3431 (N_3431,N_2580,N_2065);
or U3432 (N_3432,N_2407,N_2104);
or U3433 (N_3433,N_1828,N_2028);
or U3434 (N_3434,N_1964,N_2725);
nor U3435 (N_3435,N_2339,N_2655);
xor U3436 (N_3436,N_2505,N_2061);
xor U3437 (N_3437,N_2747,N_2372);
xor U3438 (N_3438,N_2307,N_2298);
or U3439 (N_3439,N_2961,N_1545);
nor U3440 (N_3440,N_1755,N_2932);
nand U3441 (N_3441,N_2593,N_1869);
and U3442 (N_3442,N_2690,N_2457);
and U3443 (N_3443,N_2366,N_2562);
nand U3444 (N_3444,N_1963,N_2353);
nand U3445 (N_3445,N_2717,N_1753);
and U3446 (N_3446,N_2099,N_1859);
and U3447 (N_3447,N_2760,N_2857);
nand U3448 (N_3448,N_2943,N_2954);
nand U3449 (N_3449,N_1538,N_1870);
nor U3450 (N_3450,N_2990,N_1662);
xnor U3451 (N_3451,N_2205,N_2187);
nor U3452 (N_3452,N_1593,N_1565);
nor U3453 (N_3453,N_2572,N_2250);
or U3454 (N_3454,N_1960,N_2643);
nand U3455 (N_3455,N_1821,N_2981);
nand U3456 (N_3456,N_2585,N_1738);
nand U3457 (N_3457,N_1988,N_2215);
nor U3458 (N_3458,N_2002,N_2315);
or U3459 (N_3459,N_2625,N_2464);
and U3460 (N_3460,N_1553,N_2959);
xor U3461 (N_3461,N_2952,N_2483);
or U3462 (N_3462,N_2678,N_2301);
nor U3463 (N_3463,N_1956,N_2833);
nand U3464 (N_3464,N_1743,N_2130);
xnor U3465 (N_3465,N_1754,N_2651);
nand U3466 (N_3466,N_2973,N_1622);
or U3467 (N_3467,N_1669,N_1696);
and U3468 (N_3468,N_1843,N_1813);
nor U3469 (N_3469,N_2058,N_1814);
and U3470 (N_3470,N_2511,N_2746);
nor U3471 (N_3471,N_1894,N_2522);
or U3472 (N_3472,N_2558,N_1536);
xnor U3473 (N_3473,N_2445,N_2822);
or U3474 (N_3474,N_2450,N_2924);
or U3475 (N_3475,N_2606,N_2131);
nor U3476 (N_3476,N_2368,N_2906);
nor U3477 (N_3477,N_1985,N_2258);
nand U3478 (N_3478,N_2498,N_1533);
nor U3479 (N_3479,N_1841,N_1607);
nand U3480 (N_3480,N_1768,N_2221);
or U3481 (N_3481,N_2530,N_2011);
nor U3482 (N_3482,N_2627,N_1614);
or U3483 (N_3483,N_2419,N_1670);
or U3484 (N_3484,N_1674,N_2561);
xnor U3485 (N_3485,N_2016,N_1520);
nand U3486 (N_3486,N_2921,N_1857);
nand U3487 (N_3487,N_1954,N_2111);
and U3488 (N_3488,N_2077,N_2477);
nand U3489 (N_3489,N_2045,N_1874);
nand U3490 (N_3490,N_2432,N_2023);
and U3491 (N_3491,N_2761,N_1693);
and U3492 (N_3492,N_1990,N_1798);
nor U3493 (N_3493,N_1629,N_1978);
nor U3494 (N_3494,N_1559,N_1822);
nand U3495 (N_3495,N_1913,N_1643);
nand U3496 (N_3496,N_2374,N_1929);
nand U3497 (N_3497,N_1890,N_2688);
xor U3498 (N_3498,N_2264,N_2916);
nand U3499 (N_3499,N_2533,N_1638);
nand U3500 (N_3500,N_2942,N_1879);
nand U3501 (N_3501,N_1962,N_2867);
or U3502 (N_3502,N_2577,N_2427);
or U3503 (N_3503,N_2706,N_1826);
or U3504 (N_3504,N_2995,N_1617);
nand U3505 (N_3505,N_2371,N_1996);
xor U3506 (N_3506,N_2251,N_2871);
nand U3507 (N_3507,N_1688,N_2284);
or U3508 (N_3508,N_2935,N_1862);
or U3509 (N_3509,N_2781,N_1742);
and U3510 (N_3510,N_1500,N_1718);
nand U3511 (N_3511,N_2603,N_2807);
or U3512 (N_3512,N_2014,N_1910);
or U3513 (N_3513,N_2607,N_1891);
nor U3514 (N_3514,N_1765,N_2413);
and U3515 (N_3515,N_2974,N_2482);
and U3516 (N_3516,N_2621,N_2850);
nand U3517 (N_3517,N_2765,N_2328);
nand U3518 (N_3518,N_2699,N_1965);
and U3519 (N_3519,N_1709,N_2638);
xnor U3520 (N_3520,N_1930,N_2838);
nor U3521 (N_3521,N_1951,N_2821);
nor U3522 (N_3522,N_1852,N_2784);
nor U3523 (N_3523,N_1597,N_2927);
or U3524 (N_3524,N_2810,N_1830);
nand U3525 (N_3525,N_1502,N_2854);
nor U3526 (N_3526,N_2358,N_2683);
nor U3527 (N_3527,N_1759,N_1632);
nand U3528 (N_3528,N_1657,N_1589);
nand U3529 (N_3529,N_2121,N_1574);
nor U3530 (N_3530,N_2369,N_2726);
nand U3531 (N_3531,N_2698,N_2321);
and U3532 (N_3532,N_2865,N_2138);
xnor U3533 (N_3533,N_2006,N_1947);
nand U3534 (N_3534,N_2334,N_2174);
and U3535 (N_3535,N_2762,N_2128);
or U3536 (N_3536,N_2637,N_2226);
nand U3537 (N_3537,N_1727,N_2985);
nand U3538 (N_3538,N_2844,N_2135);
nand U3539 (N_3539,N_2644,N_1836);
or U3540 (N_3540,N_1815,N_2218);
nor U3541 (N_3541,N_1904,N_2733);
or U3542 (N_3542,N_2020,N_1831);
or U3543 (N_3543,N_2094,N_1893);
nand U3544 (N_3544,N_1571,N_2292);
and U3545 (N_3545,N_1504,N_1984);
and U3546 (N_3546,N_1513,N_2642);
or U3547 (N_3547,N_2054,N_2196);
and U3548 (N_3548,N_1783,N_1613);
nor U3549 (N_3549,N_2659,N_2866);
nor U3550 (N_3550,N_2306,N_2241);
or U3551 (N_3551,N_2266,N_2386);
or U3552 (N_3552,N_2828,N_1590);
or U3553 (N_3553,N_2172,N_2695);
and U3554 (N_3554,N_2771,N_1566);
or U3555 (N_3555,N_1583,N_1582);
or U3556 (N_3556,N_1656,N_2142);
xor U3557 (N_3557,N_2109,N_1740);
nand U3558 (N_3558,N_2947,N_1720);
nor U3559 (N_3559,N_1989,N_2931);
or U3560 (N_3560,N_2519,N_2191);
and U3561 (N_3561,N_1802,N_1512);
nand U3562 (N_3562,N_2260,N_2330);
or U3563 (N_3563,N_2148,N_2414);
nand U3564 (N_3564,N_2843,N_2383);
or U3565 (N_3565,N_2424,N_2337);
and U3566 (N_3566,N_2518,N_2106);
and U3567 (N_3567,N_2704,N_2356);
nor U3568 (N_3568,N_1937,N_2105);
nor U3569 (N_3569,N_2078,N_2144);
and U3570 (N_3570,N_2708,N_1554);
nor U3571 (N_3571,N_1733,N_2211);
and U3572 (N_3572,N_2520,N_2175);
and U3573 (N_3573,N_2663,N_2460);
nand U3574 (N_3574,N_2042,N_2227);
nand U3575 (N_3575,N_2576,N_2895);
nand U3576 (N_3576,N_2165,N_2953);
nand U3577 (N_3577,N_1933,N_2048);
xor U3578 (N_3578,N_2508,N_2548);
and U3579 (N_3579,N_1776,N_1941);
nor U3580 (N_3580,N_2529,N_2304);
nor U3581 (N_3581,N_2737,N_2404);
or U3582 (N_3582,N_2013,N_1942);
xnor U3583 (N_3583,N_2030,N_2021);
and U3584 (N_3584,N_2996,N_1818);
or U3585 (N_3585,N_2249,N_2894);
and U3586 (N_3586,N_1888,N_2965);
nor U3587 (N_3587,N_2715,N_1931);
nor U3588 (N_3588,N_2905,N_2069);
nand U3589 (N_3589,N_2275,N_1932);
nand U3590 (N_3590,N_2314,N_2063);
nand U3591 (N_3591,N_1854,N_2736);
nand U3592 (N_3592,N_2711,N_2792);
or U3593 (N_3593,N_2551,N_2245);
or U3594 (N_3594,N_2429,N_2203);
nand U3595 (N_3595,N_1839,N_2841);
nor U3596 (N_3596,N_1591,N_2178);
nand U3597 (N_3597,N_1756,N_2055);
nor U3598 (N_3598,N_2122,N_2775);
or U3599 (N_3599,N_2550,N_1864);
nor U3600 (N_3600,N_2879,N_2910);
or U3601 (N_3601,N_2269,N_2976);
xnor U3602 (N_3602,N_1680,N_2597);
and U3603 (N_3603,N_2370,N_2847);
or U3604 (N_3604,N_2564,N_1615);
nor U3605 (N_3605,N_2774,N_2329);
and U3606 (N_3606,N_1675,N_2415);
nor U3607 (N_3607,N_1687,N_1855);
and U3608 (N_3608,N_2788,N_2036);
or U3609 (N_3609,N_2977,N_1983);
nand U3610 (N_3610,N_2005,N_2072);
or U3611 (N_3611,N_1794,N_2377);
or U3612 (N_3612,N_2026,N_2907);
and U3613 (N_3613,N_1604,N_2748);
or U3614 (N_3614,N_2159,N_1568);
or U3615 (N_3615,N_2236,N_2133);
nor U3616 (N_3616,N_2777,N_2700);
nand U3617 (N_3617,N_1509,N_2590);
and U3618 (N_3618,N_1880,N_2009);
or U3619 (N_3619,N_1663,N_2354);
xnor U3620 (N_3620,N_1748,N_2493);
nand U3621 (N_3621,N_2734,N_1503);
nand U3622 (N_3622,N_2791,N_2222);
and U3623 (N_3623,N_2274,N_2084);
nand U3624 (N_3624,N_1884,N_1705);
nor U3625 (N_3625,N_1979,N_2994);
or U3626 (N_3626,N_2856,N_2755);
or U3627 (N_3627,N_2035,N_2261);
nor U3628 (N_3628,N_2485,N_1572);
nand U3629 (N_3629,N_1672,N_1648);
or U3630 (N_3630,N_1575,N_2139);
nor U3631 (N_3631,N_2694,N_1620);
or U3632 (N_3632,N_2641,N_1634);
nor U3633 (N_3633,N_1551,N_1779);
and U3634 (N_3634,N_2185,N_2852);
nor U3635 (N_3635,N_2225,N_2145);
or U3636 (N_3636,N_2604,N_2615);
or U3637 (N_3637,N_2382,N_1974);
nand U3638 (N_3638,N_2080,N_1946);
or U3639 (N_3639,N_1900,N_2656);
or U3640 (N_3640,N_2399,N_2566);
nor U3641 (N_3641,N_2332,N_2010);
nor U3642 (N_3642,N_1532,N_1919);
nand U3643 (N_3643,N_2492,N_1935);
nor U3644 (N_3644,N_2851,N_2658);
or U3645 (N_3645,N_2177,N_1543);
and U3646 (N_3646,N_2473,N_2024);
nand U3647 (N_3647,N_2449,N_2436);
or U3648 (N_3648,N_1997,N_2452);
nand U3649 (N_3649,N_1986,N_2541);
nand U3650 (N_3650,N_2933,N_2724);
and U3651 (N_3651,N_1650,N_2033);
and U3652 (N_3652,N_1789,N_2614);
and U3653 (N_3653,N_2149,N_2666);
nand U3654 (N_3654,N_2691,N_2620);
and U3655 (N_3655,N_2201,N_2246);
nand U3656 (N_3656,N_2333,N_1677);
or U3657 (N_3657,N_1982,N_2158);
nand U3658 (N_3658,N_2209,N_2110);
xnor U3659 (N_3659,N_2898,N_2675);
nand U3660 (N_3660,N_1528,N_2540);
nand U3661 (N_3661,N_1726,N_1834);
or U3662 (N_3662,N_2862,N_1577);
or U3663 (N_3663,N_2458,N_2723);
nor U3664 (N_3664,N_2230,N_1658);
or U3665 (N_3665,N_1948,N_2311);
nor U3666 (N_3666,N_1561,N_1928);
and U3667 (N_3667,N_2441,N_2526);
xor U3668 (N_3668,N_1624,N_2859);
xnor U3669 (N_3669,N_2141,N_2357);
and U3670 (N_3670,N_2767,N_1920);
nor U3671 (N_3671,N_2661,N_1697);
nand U3672 (N_3672,N_1682,N_2390);
nor U3673 (N_3673,N_2112,N_2465);
and U3674 (N_3674,N_2770,N_2884);
or U3675 (N_3675,N_2632,N_1712);
nor U3676 (N_3676,N_2967,N_2721);
or U3677 (N_3677,N_2565,N_2443);
or U3678 (N_3678,N_2206,N_2757);
or U3679 (N_3679,N_2004,N_2926);
nand U3680 (N_3680,N_2720,N_1596);
and U3681 (N_3681,N_1971,N_2647);
and U3682 (N_3682,N_2279,N_2842);
or U3683 (N_3683,N_2428,N_2100);
nand U3684 (N_3684,N_2189,N_2912);
and U3685 (N_3685,N_1903,N_2456);
or U3686 (N_3686,N_2327,N_1610);
nand U3687 (N_3687,N_2214,N_1763);
nor U3688 (N_3688,N_2280,N_1644);
nor U3689 (N_3689,N_2855,N_1685);
nor U3690 (N_3690,N_2411,N_2730);
or U3691 (N_3691,N_2412,N_2180);
nand U3692 (N_3692,N_2151,N_2499);
and U3693 (N_3693,N_2649,N_2968);
xnor U3694 (N_3694,N_2516,N_2003);
and U3695 (N_3695,N_2114,N_1950);
xor U3696 (N_3696,N_2039,N_1844);
nand U3697 (N_3697,N_1872,N_1736);
nor U3698 (N_3698,N_1876,N_1570);
nor U3699 (N_3699,N_2442,N_2962);
nand U3700 (N_3700,N_1508,N_2232);
and U3701 (N_3701,N_2381,N_2338);
and U3702 (N_3702,N_1981,N_2008);
and U3703 (N_3703,N_2389,N_2502);
nand U3704 (N_3704,N_2824,N_2331);
nand U3705 (N_3705,N_2235,N_1923);
and U3706 (N_3706,N_2887,N_2117);
or U3707 (N_3707,N_2062,N_1957);
or U3708 (N_3708,N_2812,N_1993);
nand U3709 (N_3709,N_1717,N_2626);
nand U3710 (N_3710,N_1780,N_2018);
or U3711 (N_3711,N_2490,N_1873);
nand U3712 (N_3712,N_2425,N_1781);
or U3713 (N_3713,N_2744,N_2582);
or U3714 (N_3714,N_2302,N_1871);
or U3715 (N_3715,N_2677,N_2975);
or U3716 (N_3716,N_1912,N_2047);
nand U3717 (N_3717,N_1832,N_2612);
and U3718 (N_3718,N_2633,N_1881);
or U3719 (N_3719,N_2794,N_1917);
or U3720 (N_3720,N_2041,N_2902);
nand U3721 (N_3721,N_2350,N_1714);
nand U3722 (N_3722,N_2630,N_2776);
and U3723 (N_3723,N_2839,N_1868);
nor U3724 (N_3724,N_2223,N_1799);
and U3725 (N_3725,N_2524,N_2915);
or U3726 (N_3726,N_1695,N_2296);
or U3727 (N_3727,N_1926,N_2707);
nor U3728 (N_3728,N_2545,N_2293);
or U3729 (N_3729,N_2217,N_2231);
nand U3730 (N_3730,N_1761,N_1706);
nor U3731 (N_3731,N_2081,N_2440);
nor U3732 (N_3732,N_1812,N_2556);
nor U3733 (N_3733,N_2507,N_2313);
and U3734 (N_3734,N_2539,N_1824);
nor U3735 (N_3735,N_1627,N_2779);
or U3736 (N_3736,N_1790,N_1580);
nor U3737 (N_3737,N_1749,N_2107);
and U3738 (N_3738,N_2134,N_2444);
or U3739 (N_3739,N_2999,N_2076);
nand U3740 (N_3740,N_2993,N_2239);
nand U3741 (N_3741,N_1899,N_2380);
xor U3742 (N_3742,N_2631,N_1576);
or U3743 (N_3743,N_2012,N_2375);
nand U3744 (N_3744,N_2092,N_1713);
and U3745 (N_3745,N_2417,N_1681);
nor U3746 (N_3746,N_1730,N_2578);
nor U3747 (N_3747,N_1762,N_2157);
nor U3748 (N_3748,N_2146,N_1896);
nand U3749 (N_3749,N_2923,N_2749);
and U3750 (N_3750,N_2640,N_2636);
or U3751 (N_3751,N_2331,N_2677);
or U3752 (N_3752,N_2319,N_2279);
and U3753 (N_3753,N_2979,N_2958);
or U3754 (N_3754,N_2170,N_2544);
and U3755 (N_3755,N_2901,N_2094);
nand U3756 (N_3756,N_2573,N_2627);
or U3757 (N_3757,N_1860,N_1574);
nand U3758 (N_3758,N_2967,N_2608);
or U3759 (N_3759,N_2542,N_2097);
nand U3760 (N_3760,N_1965,N_1735);
nor U3761 (N_3761,N_1842,N_2462);
nand U3762 (N_3762,N_2157,N_2272);
nor U3763 (N_3763,N_2707,N_2804);
and U3764 (N_3764,N_1766,N_2477);
or U3765 (N_3765,N_1802,N_2903);
nor U3766 (N_3766,N_1984,N_1822);
nor U3767 (N_3767,N_2319,N_2318);
and U3768 (N_3768,N_1558,N_2409);
nand U3769 (N_3769,N_1949,N_1928);
nand U3770 (N_3770,N_2404,N_2155);
xor U3771 (N_3771,N_1902,N_1947);
or U3772 (N_3772,N_2538,N_1981);
nor U3773 (N_3773,N_2061,N_2776);
or U3774 (N_3774,N_2355,N_2505);
xor U3775 (N_3775,N_2987,N_2126);
or U3776 (N_3776,N_2304,N_2444);
nor U3777 (N_3777,N_2731,N_2628);
nand U3778 (N_3778,N_1829,N_1639);
nor U3779 (N_3779,N_2310,N_1583);
xnor U3780 (N_3780,N_2207,N_2480);
nand U3781 (N_3781,N_2403,N_2982);
and U3782 (N_3782,N_2468,N_1522);
nor U3783 (N_3783,N_2376,N_1819);
xnor U3784 (N_3784,N_2835,N_2292);
nand U3785 (N_3785,N_1626,N_1879);
or U3786 (N_3786,N_2307,N_1643);
and U3787 (N_3787,N_2996,N_2128);
nand U3788 (N_3788,N_2754,N_2567);
and U3789 (N_3789,N_2098,N_2958);
nand U3790 (N_3790,N_2696,N_1755);
or U3791 (N_3791,N_2919,N_2568);
nor U3792 (N_3792,N_2523,N_2551);
nor U3793 (N_3793,N_2557,N_2848);
nor U3794 (N_3794,N_2627,N_1622);
xor U3795 (N_3795,N_2559,N_1928);
nand U3796 (N_3796,N_2788,N_1692);
nor U3797 (N_3797,N_2468,N_1777);
and U3798 (N_3798,N_1856,N_2608);
or U3799 (N_3799,N_2607,N_2990);
nor U3800 (N_3800,N_2671,N_2976);
or U3801 (N_3801,N_2065,N_2661);
and U3802 (N_3802,N_1767,N_2595);
and U3803 (N_3803,N_2216,N_2035);
xor U3804 (N_3804,N_1632,N_1668);
xnor U3805 (N_3805,N_2603,N_2032);
nand U3806 (N_3806,N_2164,N_1646);
xor U3807 (N_3807,N_2103,N_1972);
and U3808 (N_3808,N_1659,N_2249);
nor U3809 (N_3809,N_2673,N_2119);
xnor U3810 (N_3810,N_2572,N_1818);
xnor U3811 (N_3811,N_1955,N_2955);
or U3812 (N_3812,N_1764,N_1991);
and U3813 (N_3813,N_2167,N_2221);
nor U3814 (N_3814,N_2051,N_2469);
or U3815 (N_3815,N_2739,N_1951);
nand U3816 (N_3816,N_2716,N_2303);
nor U3817 (N_3817,N_2243,N_2901);
and U3818 (N_3818,N_2417,N_2718);
nor U3819 (N_3819,N_2586,N_2460);
nand U3820 (N_3820,N_1577,N_2473);
nand U3821 (N_3821,N_2542,N_1775);
xor U3822 (N_3822,N_2876,N_1589);
and U3823 (N_3823,N_1879,N_2934);
xnor U3824 (N_3824,N_2452,N_2333);
nor U3825 (N_3825,N_2485,N_2824);
xor U3826 (N_3826,N_1788,N_2531);
and U3827 (N_3827,N_1987,N_2594);
nand U3828 (N_3828,N_1798,N_2965);
or U3829 (N_3829,N_2467,N_2393);
or U3830 (N_3830,N_2233,N_2999);
and U3831 (N_3831,N_2392,N_2635);
or U3832 (N_3832,N_2074,N_2200);
nor U3833 (N_3833,N_2209,N_2026);
and U3834 (N_3834,N_1548,N_2659);
xnor U3835 (N_3835,N_1735,N_2311);
xnor U3836 (N_3836,N_2629,N_2067);
nor U3837 (N_3837,N_1872,N_2279);
nand U3838 (N_3838,N_2624,N_2321);
or U3839 (N_3839,N_2970,N_1715);
and U3840 (N_3840,N_1553,N_1741);
or U3841 (N_3841,N_1521,N_2585);
xor U3842 (N_3842,N_2348,N_2022);
and U3843 (N_3843,N_2646,N_2566);
or U3844 (N_3844,N_2217,N_2807);
nor U3845 (N_3845,N_2868,N_2441);
nor U3846 (N_3846,N_2070,N_1767);
nand U3847 (N_3847,N_2992,N_2323);
nand U3848 (N_3848,N_1721,N_2029);
xor U3849 (N_3849,N_2661,N_2854);
and U3850 (N_3850,N_2318,N_1585);
or U3851 (N_3851,N_2054,N_2520);
and U3852 (N_3852,N_2677,N_2282);
nor U3853 (N_3853,N_2839,N_2908);
xor U3854 (N_3854,N_1993,N_2103);
or U3855 (N_3855,N_1822,N_2004);
or U3856 (N_3856,N_1876,N_2143);
nor U3857 (N_3857,N_2360,N_1609);
nor U3858 (N_3858,N_2728,N_2601);
nor U3859 (N_3859,N_1692,N_1720);
and U3860 (N_3860,N_1995,N_2369);
nor U3861 (N_3861,N_1835,N_2207);
and U3862 (N_3862,N_2464,N_1500);
or U3863 (N_3863,N_2270,N_1721);
or U3864 (N_3864,N_2710,N_2554);
and U3865 (N_3865,N_2353,N_2452);
nand U3866 (N_3866,N_2265,N_2859);
and U3867 (N_3867,N_1815,N_1954);
or U3868 (N_3868,N_1688,N_1737);
and U3869 (N_3869,N_2495,N_1716);
or U3870 (N_3870,N_1681,N_1578);
nand U3871 (N_3871,N_1955,N_1660);
and U3872 (N_3872,N_2393,N_2532);
nor U3873 (N_3873,N_2994,N_2658);
xnor U3874 (N_3874,N_1931,N_2679);
and U3875 (N_3875,N_1569,N_2462);
or U3876 (N_3876,N_2509,N_2436);
or U3877 (N_3877,N_1822,N_2068);
xor U3878 (N_3878,N_2809,N_2984);
nand U3879 (N_3879,N_1538,N_2121);
and U3880 (N_3880,N_1754,N_2297);
nor U3881 (N_3881,N_2912,N_1756);
or U3882 (N_3882,N_2600,N_2041);
and U3883 (N_3883,N_2093,N_2306);
xnor U3884 (N_3884,N_2413,N_2803);
nand U3885 (N_3885,N_2596,N_1702);
or U3886 (N_3886,N_2143,N_1973);
nand U3887 (N_3887,N_2816,N_2148);
nor U3888 (N_3888,N_2284,N_2480);
xnor U3889 (N_3889,N_2452,N_2916);
nand U3890 (N_3890,N_2495,N_1960);
xor U3891 (N_3891,N_1956,N_2076);
or U3892 (N_3892,N_1686,N_2886);
nor U3893 (N_3893,N_2738,N_1954);
nand U3894 (N_3894,N_1509,N_1975);
and U3895 (N_3895,N_2171,N_2923);
or U3896 (N_3896,N_1626,N_2029);
and U3897 (N_3897,N_1946,N_2115);
or U3898 (N_3898,N_2340,N_2406);
and U3899 (N_3899,N_2361,N_2006);
and U3900 (N_3900,N_1573,N_2527);
and U3901 (N_3901,N_1905,N_1713);
or U3902 (N_3902,N_2583,N_1911);
or U3903 (N_3903,N_2633,N_1971);
nor U3904 (N_3904,N_2722,N_2077);
and U3905 (N_3905,N_2607,N_2103);
nor U3906 (N_3906,N_2615,N_1610);
or U3907 (N_3907,N_2542,N_1644);
nor U3908 (N_3908,N_2551,N_2133);
nand U3909 (N_3909,N_2608,N_1801);
or U3910 (N_3910,N_2675,N_2328);
xnor U3911 (N_3911,N_1768,N_2080);
or U3912 (N_3912,N_2235,N_1730);
and U3913 (N_3913,N_2807,N_2139);
xnor U3914 (N_3914,N_2507,N_2723);
and U3915 (N_3915,N_2733,N_2139);
and U3916 (N_3916,N_1688,N_1891);
or U3917 (N_3917,N_1607,N_2797);
nor U3918 (N_3918,N_1641,N_1853);
xor U3919 (N_3919,N_1683,N_2203);
nand U3920 (N_3920,N_1683,N_2679);
nor U3921 (N_3921,N_2725,N_1717);
nand U3922 (N_3922,N_2219,N_1873);
nor U3923 (N_3923,N_1882,N_2534);
nor U3924 (N_3924,N_1588,N_2742);
xnor U3925 (N_3925,N_2367,N_2765);
nor U3926 (N_3926,N_2427,N_2449);
nand U3927 (N_3927,N_2072,N_2762);
nor U3928 (N_3928,N_2119,N_1679);
nor U3929 (N_3929,N_2929,N_2498);
and U3930 (N_3930,N_1705,N_1504);
and U3931 (N_3931,N_2157,N_2840);
and U3932 (N_3932,N_2147,N_2922);
or U3933 (N_3933,N_2011,N_1990);
nand U3934 (N_3934,N_2745,N_2054);
xnor U3935 (N_3935,N_1599,N_1724);
and U3936 (N_3936,N_2200,N_1949);
and U3937 (N_3937,N_1987,N_2558);
or U3938 (N_3938,N_1643,N_2009);
or U3939 (N_3939,N_1920,N_2484);
nor U3940 (N_3940,N_2735,N_1866);
nand U3941 (N_3941,N_2837,N_1947);
and U3942 (N_3942,N_2001,N_2522);
and U3943 (N_3943,N_2685,N_2729);
and U3944 (N_3944,N_2338,N_2070);
and U3945 (N_3945,N_1580,N_2857);
nand U3946 (N_3946,N_2286,N_2379);
or U3947 (N_3947,N_2791,N_2449);
nand U3948 (N_3948,N_2386,N_1673);
nor U3949 (N_3949,N_2542,N_1980);
nor U3950 (N_3950,N_2488,N_1692);
nand U3951 (N_3951,N_2675,N_1768);
or U3952 (N_3952,N_1742,N_1682);
nor U3953 (N_3953,N_2175,N_2056);
nand U3954 (N_3954,N_2051,N_2311);
nor U3955 (N_3955,N_2712,N_2138);
nor U3956 (N_3956,N_2646,N_2402);
and U3957 (N_3957,N_2605,N_2243);
and U3958 (N_3958,N_2551,N_1619);
nor U3959 (N_3959,N_1786,N_1995);
nand U3960 (N_3960,N_2588,N_2798);
and U3961 (N_3961,N_2173,N_2188);
or U3962 (N_3962,N_2234,N_2625);
and U3963 (N_3963,N_1651,N_2366);
nor U3964 (N_3964,N_2354,N_2349);
and U3965 (N_3965,N_2970,N_1659);
and U3966 (N_3966,N_2790,N_2840);
or U3967 (N_3967,N_2056,N_2533);
and U3968 (N_3968,N_2101,N_2856);
or U3969 (N_3969,N_2466,N_2272);
and U3970 (N_3970,N_1846,N_2929);
nand U3971 (N_3971,N_2253,N_1549);
and U3972 (N_3972,N_2805,N_2871);
or U3973 (N_3973,N_1505,N_2706);
nand U3974 (N_3974,N_2042,N_1968);
and U3975 (N_3975,N_2987,N_2692);
or U3976 (N_3976,N_2942,N_1514);
and U3977 (N_3977,N_2130,N_2480);
xor U3978 (N_3978,N_1744,N_1694);
nand U3979 (N_3979,N_2176,N_1928);
and U3980 (N_3980,N_2817,N_2683);
and U3981 (N_3981,N_2084,N_2927);
nand U3982 (N_3982,N_2998,N_2692);
nand U3983 (N_3983,N_1860,N_2949);
and U3984 (N_3984,N_2125,N_2704);
and U3985 (N_3985,N_2939,N_2151);
and U3986 (N_3986,N_2656,N_2297);
or U3987 (N_3987,N_1656,N_2033);
or U3988 (N_3988,N_2224,N_2886);
nand U3989 (N_3989,N_2568,N_2569);
nand U3990 (N_3990,N_1791,N_1746);
nand U3991 (N_3991,N_1811,N_1576);
xor U3992 (N_3992,N_2418,N_1867);
nor U3993 (N_3993,N_1598,N_2550);
and U3994 (N_3994,N_2122,N_2582);
and U3995 (N_3995,N_2081,N_2048);
nand U3996 (N_3996,N_2195,N_1614);
nor U3997 (N_3997,N_2080,N_2507);
nand U3998 (N_3998,N_2697,N_2417);
and U3999 (N_3999,N_2217,N_1861);
nand U4000 (N_4000,N_2125,N_1821);
or U4001 (N_4001,N_1949,N_2284);
nor U4002 (N_4002,N_2985,N_1755);
xnor U4003 (N_4003,N_2147,N_1784);
xnor U4004 (N_4004,N_1505,N_2563);
nand U4005 (N_4005,N_2358,N_1556);
nand U4006 (N_4006,N_2965,N_2256);
and U4007 (N_4007,N_2764,N_1880);
and U4008 (N_4008,N_2115,N_2172);
and U4009 (N_4009,N_2627,N_2534);
nor U4010 (N_4010,N_1970,N_2468);
or U4011 (N_4011,N_2874,N_2237);
and U4012 (N_4012,N_2768,N_1979);
nor U4013 (N_4013,N_1832,N_2558);
and U4014 (N_4014,N_2231,N_2861);
and U4015 (N_4015,N_1749,N_2571);
or U4016 (N_4016,N_2085,N_1683);
nand U4017 (N_4017,N_2483,N_2641);
nor U4018 (N_4018,N_2380,N_2544);
and U4019 (N_4019,N_2907,N_1587);
or U4020 (N_4020,N_2065,N_2121);
xor U4021 (N_4021,N_2663,N_2338);
and U4022 (N_4022,N_2224,N_2664);
nor U4023 (N_4023,N_2835,N_2774);
nand U4024 (N_4024,N_2000,N_2678);
and U4025 (N_4025,N_2153,N_2885);
nor U4026 (N_4026,N_1734,N_2333);
or U4027 (N_4027,N_2425,N_2584);
nor U4028 (N_4028,N_2814,N_2562);
nand U4029 (N_4029,N_1626,N_2592);
xnor U4030 (N_4030,N_1537,N_2659);
and U4031 (N_4031,N_2621,N_2121);
nor U4032 (N_4032,N_1713,N_2718);
and U4033 (N_4033,N_1623,N_2614);
xor U4034 (N_4034,N_2007,N_2196);
nor U4035 (N_4035,N_1653,N_2338);
or U4036 (N_4036,N_2916,N_1871);
nand U4037 (N_4037,N_2478,N_2199);
and U4038 (N_4038,N_2047,N_2406);
nor U4039 (N_4039,N_1656,N_1960);
and U4040 (N_4040,N_1741,N_2082);
nor U4041 (N_4041,N_2231,N_2995);
nand U4042 (N_4042,N_2146,N_2989);
nand U4043 (N_4043,N_2260,N_2607);
nor U4044 (N_4044,N_1992,N_1869);
or U4045 (N_4045,N_1592,N_2336);
nand U4046 (N_4046,N_2848,N_2243);
or U4047 (N_4047,N_1947,N_2789);
nor U4048 (N_4048,N_2617,N_2065);
or U4049 (N_4049,N_1641,N_2263);
nor U4050 (N_4050,N_2790,N_1882);
or U4051 (N_4051,N_2254,N_2445);
and U4052 (N_4052,N_1515,N_2781);
nand U4053 (N_4053,N_2483,N_2560);
and U4054 (N_4054,N_2285,N_1990);
nor U4055 (N_4055,N_2928,N_2892);
or U4056 (N_4056,N_1750,N_2618);
or U4057 (N_4057,N_2487,N_1898);
or U4058 (N_4058,N_2484,N_1854);
or U4059 (N_4059,N_2825,N_2572);
nand U4060 (N_4060,N_2267,N_2268);
nand U4061 (N_4061,N_1745,N_2792);
nor U4062 (N_4062,N_2306,N_1582);
nand U4063 (N_4063,N_2651,N_1636);
nand U4064 (N_4064,N_2915,N_2330);
nand U4065 (N_4065,N_2598,N_2694);
xor U4066 (N_4066,N_2714,N_2221);
or U4067 (N_4067,N_2942,N_1862);
nor U4068 (N_4068,N_2094,N_2886);
nand U4069 (N_4069,N_2260,N_2545);
or U4070 (N_4070,N_2418,N_2843);
nor U4071 (N_4071,N_1978,N_1931);
nand U4072 (N_4072,N_1547,N_2319);
nand U4073 (N_4073,N_2748,N_2141);
and U4074 (N_4074,N_2528,N_2647);
nand U4075 (N_4075,N_1740,N_2398);
and U4076 (N_4076,N_1989,N_2165);
nand U4077 (N_4077,N_2547,N_1675);
and U4078 (N_4078,N_2370,N_1753);
nor U4079 (N_4079,N_2016,N_1620);
nand U4080 (N_4080,N_2294,N_2379);
nor U4081 (N_4081,N_2022,N_2080);
nand U4082 (N_4082,N_1884,N_2308);
nand U4083 (N_4083,N_1969,N_2382);
or U4084 (N_4084,N_2659,N_1946);
and U4085 (N_4085,N_1636,N_2806);
nor U4086 (N_4086,N_1696,N_2626);
or U4087 (N_4087,N_2772,N_2233);
or U4088 (N_4088,N_2416,N_2937);
or U4089 (N_4089,N_2623,N_2057);
or U4090 (N_4090,N_2323,N_2013);
or U4091 (N_4091,N_2754,N_1906);
nand U4092 (N_4092,N_2454,N_2882);
or U4093 (N_4093,N_2431,N_2784);
nor U4094 (N_4094,N_2816,N_2766);
and U4095 (N_4095,N_2336,N_2617);
nor U4096 (N_4096,N_2127,N_2960);
and U4097 (N_4097,N_2347,N_2187);
or U4098 (N_4098,N_2572,N_1916);
and U4099 (N_4099,N_2536,N_2910);
or U4100 (N_4100,N_2439,N_1839);
nor U4101 (N_4101,N_1792,N_1630);
xnor U4102 (N_4102,N_2481,N_2029);
or U4103 (N_4103,N_2339,N_1905);
and U4104 (N_4104,N_2210,N_2297);
and U4105 (N_4105,N_2806,N_1561);
or U4106 (N_4106,N_2582,N_1783);
or U4107 (N_4107,N_2231,N_2097);
or U4108 (N_4108,N_1618,N_2160);
nor U4109 (N_4109,N_2727,N_1711);
nor U4110 (N_4110,N_1822,N_2891);
nor U4111 (N_4111,N_2351,N_2797);
nor U4112 (N_4112,N_2337,N_2702);
nand U4113 (N_4113,N_1671,N_2487);
nand U4114 (N_4114,N_2610,N_1992);
nand U4115 (N_4115,N_1752,N_2854);
and U4116 (N_4116,N_2198,N_2260);
or U4117 (N_4117,N_1561,N_2374);
nor U4118 (N_4118,N_1527,N_2079);
xnor U4119 (N_4119,N_2243,N_2251);
nor U4120 (N_4120,N_1546,N_2971);
or U4121 (N_4121,N_2874,N_1589);
or U4122 (N_4122,N_2046,N_2684);
xor U4123 (N_4123,N_2435,N_1841);
nand U4124 (N_4124,N_2474,N_2039);
or U4125 (N_4125,N_2512,N_2074);
nand U4126 (N_4126,N_2846,N_2752);
and U4127 (N_4127,N_1945,N_1724);
nand U4128 (N_4128,N_1597,N_2271);
and U4129 (N_4129,N_2308,N_2521);
nand U4130 (N_4130,N_2498,N_1600);
or U4131 (N_4131,N_2351,N_2756);
nor U4132 (N_4132,N_2337,N_1742);
nand U4133 (N_4133,N_2411,N_2574);
xor U4134 (N_4134,N_1794,N_2600);
nand U4135 (N_4135,N_2285,N_1518);
nand U4136 (N_4136,N_1817,N_1585);
or U4137 (N_4137,N_2771,N_2494);
or U4138 (N_4138,N_2378,N_2932);
nand U4139 (N_4139,N_2666,N_1771);
and U4140 (N_4140,N_2164,N_1916);
or U4141 (N_4141,N_2384,N_2799);
nor U4142 (N_4142,N_1674,N_2291);
and U4143 (N_4143,N_2896,N_1572);
nand U4144 (N_4144,N_2809,N_1627);
nand U4145 (N_4145,N_1592,N_1624);
and U4146 (N_4146,N_1788,N_1523);
xnor U4147 (N_4147,N_2984,N_2968);
nor U4148 (N_4148,N_2794,N_2344);
or U4149 (N_4149,N_2344,N_2561);
nor U4150 (N_4150,N_2667,N_2218);
and U4151 (N_4151,N_2438,N_2581);
nor U4152 (N_4152,N_1612,N_1616);
and U4153 (N_4153,N_2904,N_1804);
nor U4154 (N_4154,N_2719,N_2341);
or U4155 (N_4155,N_2237,N_2697);
nor U4156 (N_4156,N_2962,N_2559);
nand U4157 (N_4157,N_2946,N_2125);
nand U4158 (N_4158,N_2308,N_2667);
and U4159 (N_4159,N_2113,N_2232);
nor U4160 (N_4160,N_2253,N_2769);
or U4161 (N_4161,N_2285,N_2598);
and U4162 (N_4162,N_2843,N_2105);
and U4163 (N_4163,N_2967,N_1516);
xor U4164 (N_4164,N_2933,N_1954);
nand U4165 (N_4165,N_2686,N_1972);
xnor U4166 (N_4166,N_2329,N_1892);
and U4167 (N_4167,N_1795,N_1906);
and U4168 (N_4168,N_2300,N_1587);
nand U4169 (N_4169,N_2400,N_1595);
and U4170 (N_4170,N_2848,N_2726);
xor U4171 (N_4171,N_2794,N_1719);
or U4172 (N_4172,N_2142,N_1706);
or U4173 (N_4173,N_1750,N_2857);
nand U4174 (N_4174,N_2544,N_2680);
or U4175 (N_4175,N_2789,N_2707);
and U4176 (N_4176,N_1855,N_2514);
nor U4177 (N_4177,N_1819,N_2465);
nand U4178 (N_4178,N_1609,N_1876);
or U4179 (N_4179,N_2235,N_2003);
nor U4180 (N_4180,N_2328,N_2234);
nand U4181 (N_4181,N_2665,N_1657);
and U4182 (N_4182,N_2176,N_1540);
xnor U4183 (N_4183,N_2915,N_1850);
nor U4184 (N_4184,N_2566,N_1567);
nand U4185 (N_4185,N_2842,N_2010);
or U4186 (N_4186,N_2612,N_2431);
xnor U4187 (N_4187,N_2236,N_1525);
xnor U4188 (N_4188,N_2972,N_2643);
nor U4189 (N_4189,N_2649,N_1939);
and U4190 (N_4190,N_1805,N_2777);
or U4191 (N_4191,N_1774,N_2279);
nor U4192 (N_4192,N_1934,N_1996);
nor U4193 (N_4193,N_1974,N_2443);
or U4194 (N_4194,N_1589,N_2120);
or U4195 (N_4195,N_1707,N_1721);
and U4196 (N_4196,N_1627,N_2846);
nand U4197 (N_4197,N_2493,N_1612);
nor U4198 (N_4198,N_2400,N_1712);
nand U4199 (N_4199,N_2581,N_2795);
nor U4200 (N_4200,N_2287,N_2474);
nand U4201 (N_4201,N_2503,N_2116);
xnor U4202 (N_4202,N_2269,N_1967);
and U4203 (N_4203,N_2246,N_1570);
nand U4204 (N_4204,N_1772,N_2414);
xnor U4205 (N_4205,N_1601,N_2858);
nor U4206 (N_4206,N_2326,N_1593);
nor U4207 (N_4207,N_2163,N_1850);
or U4208 (N_4208,N_1540,N_1753);
or U4209 (N_4209,N_2926,N_1734);
and U4210 (N_4210,N_2822,N_2763);
xor U4211 (N_4211,N_2046,N_2629);
xor U4212 (N_4212,N_1979,N_1734);
nand U4213 (N_4213,N_2049,N_2211);
and U4214 (N_4214,N_1721,N_2302);
and U4215 (N_4215,N_2738,N_2136);
and U4216 (N_4216,N_2070,N_2932);
nor U4217 (N_4217,N_2720,N_1844);
nor U4218 (N_4218,N_2889,N_2038);
xnor U4219 (N_4219,N_1504,N_2436);
nor U4220 (N_4220,N_2655,N_2503);
nand U4221 (N_4221,N_1762,N_1639);
nand U4222 (N_4222,N_2834,N_2229);
and U4223 (N_4223,N_1845,N_2952);
nor U4224 (N_4224,N_2294,N_1522);
nor U4225 (N_4225,N_2645,N_2125);
nor U4226 (N_4226,N_1914,N_1813);
nand U4227 (N_4227,N_1735,N_1550);
nand U4228 (N_4228,N_1712,N_1793);
xnor U4229 (N_4229,N_1506,N_2390);
nor U4230 (N_4230,N_2194,N_1872);
xnor U4231 (N_4231,N_2828,N_1833);
xor U4232 (N_4232,N_1521,N_1905);
nand U4233 (N_4233,N_2985,N_1724);
or U4234 (N_4234,N_1783,N_2804);
nor U4235 (N_4235,N_2129,N_2159);
nand U4236 (N_4236,N_2705,N_1694);
xnor U4237 (N_4237,N_2336,N_2415);
or U4238 (N_4238,N_1573,N_1692);
xor U4239 (N_4239,N_2499,N_2270);
or U4240 (N_4240,N_2414,N_2136);
nand U4241 (N_4241,N_2020,N_2751);
or U4242 (N_4242,N_2326,N_2332);
xnor U4243 (N_4243,N_1524,N_2545);
xor U4244 (N_4244,N_2282,N_1988);
and U4245 (N_4245,N_1670,N_1593);
nand U4246 (N_4246,N_1822,N_2073);
and U4247 (N_4247,N_2063,N_2765);
xnor U4248 (N_4248,N_1558,N_2439);
or U4249 (N_4249,N_2530,N_1708);
xnor U4250 (N_4250,N_2186,N_2442);
nor U4251 (N_4251,N_2488,N_2715);
or U4252 (N_4252,N_2893,N_1522);
or U4253 (N_4253,N_2897,N_2204);
xor U4254 (N_4254,N_1939,N_1696);
nor U4255 (N_4255,N_2401,N_2436);
or U4256 (N_4256,N_2673,N_2757);
or U4257 (N_4257,N_2444,N_2879);
and U4258 (N_4258,N_2946,N_2967);
nand U4259 (N_4259,N_2259,N_2860);
and U4260 (N_4260,N_2140,N_1948);
and U4261 (N_4261,N_1859,N_1654);
or U4262 (N_4262,N_1582,N_2810);
or U4263 (N_4263,N_1519,N_2626);
or U4264 (N_4264,N_2473,N_1849);
nand U4265 (N_4265,N_1805,N_2085);
or U4266 (N_4266,N_2064,N_1943);
xnor U4267 (N_4267,N_1816,N_1692);
xor U4268 (N_4268,N_2111,N_2078);
nor U4269 (N_4269,N_1946,N_1759);
nor U4270 (N_4270,N_2344,N_1602);
and U4271 (N_4271,N_1718,N_2357);
or U4272 (N_4272,N_1813,N_2224);
nand U4273 (N_4273,N_2087,N_1975);
or U4274 (N_4274,N_1571,N_2500);
or U4275 (N_4275,N_1978,N_1991);
nor U4276 (N_4276,N_2447,N_2902);
xor U4277 (N_4277,N_1959,N_2934);
nor U4278 (N_4278,N_2615,N_1878);
xnor U4279 (N_4279,N_2146,N_2235);
and U4280 (N_4280,N_2910,N_2706);
nand U4281 (N_4281,N_2200,N_1840);
nand U4282 (N_4282,N_1844,N_2656);
nor U4283 (N_4283,N_2135,N_1658);
nand U4284 (N_4284,N_1926,N_2071);
nor U4285 (N_4285,N_2577,N_1746);
or U4286 (N_4286,N_1908,N_2522);
or U4287 (N_4287,N_2446,N_2817);
nand U4288 (N_4288,N_2683,N_2273);
or U4289 (N_4289,N_2242,N_2783);
xnor U4290 (N_4290,N_2034,N_2395);
and U4291 (N_4291,N_1937,N_1874);
and U4292 (N_4292,N_2093,N_2299);
and U4293 (N_4293,N_1701,N_2051);
nor U4294 (N_4294,N_2469,N_1687);
nand U4295 (N_4295,N_1824,N_1633);
nand U4296 (N_4296,N_2681,N_2216);
nand U4297 (N_4297,N_1902,N_2785);
or U4298 (N_4298,N_2542,N_1666);
or U4299 (N_4299,N_2291,N_1828);
nand U4300 (N_4300,N_2726,N_1592);
nor U4301 (N_4301,N_2304,N_2757);
xor U4302 (N_4302,N_2748,N_2198);
or U4303 (N_4303,N_1968,N_1894);
nand U4304 (N_4304,N_1532,N_1784);
nor U4305 (N_4305,N_2917,N_2306);
or U4306 (N_4306,N_2070,N_2551);
nor U4307 (N_4307,N_2188,N_1638);
nor U4308 (N_4308,N_1696,N_1821);
xnor U4309 (N_4309,N_2424,N_1738);
xor U4310 (N_4310,N_2963,N_1590);
nand U4311 (N_4311,N_2708,N_1946);
nand U4312 (N_4312,N_2296,N_2993);
or U4313 (N_4313,N_1891,N_2224);
xor U4314 (N_4314,N_2321,N_2731);
or U4315 (N_4315,N_2195,N_2506);
and U4316 (N_4316,N_2966,N_1701);
and U4317 (N_4317,N_2696,N_2470);
nand U4318 (N_4318,N_2939,N_1563);
nand U4319 (N_4319,N_2535,N_2695);
and U4320 (N_4320,N_2946,N_2899);
or U4321 (N_4321,N_1556,N_2008);
and U4322 (N_4322,N_2383,N_1501);
and U4323 (N_4323,N_1883,N_1915);
nand U4324 (N_4324,N_1688,N_2326);
or U4325 (N_4325,N_2630,N_2904);
and U4326 (N_4326,N_2885,N_2040);
nor U4327 (N_4327,N_1820,N_1536);
nor U4328 (N_4328,N_2999,N_1569);
and U4329 (N_4329,N_1796,N_1736);
nor U4330 (N_4330,N_2973,N_1727);
nand U4331 (N_4331,N_1861,N_1806);
or U4332 (N_4332,N_1539,N_2692);
and U4333 (N_4333,N_2561,N_1615);
or U4334 (N_4334,N_1531,N_1825);
nand U4335 (N_4335,N_2058,N_2120);
and U4336 (N_4336,N_2654,N_2920);
nor U4337 (N_4337,N_2246,N_2003);
nand U4338 (N_4338,N_2988,N_2249);
or U4339 (N_4339,N_2168,N_2983);
and U4340 (N_4340,N_2978,N_2921);
or U4341 (N_4341,N_2896,N_2830);
or U4342 (N_4342,N_2073,N_2300);
and U4343 (N_4343,N_2669,N_2058);
or U4344 (N_4344,N_1754,N_2831);
xor U4345 (N_4345,N_2521,N_2759);
nand U4346 (N_4346,N_2109,N_2391);
nor U4347 (N_4347,N_1794,N_1639);
nand U4348 (N_4348,N_1743,N_1972);
and U4349 (N_4349,N_2310,N_2700);
and U4350 (N_4350,N_2573,N_2202);
nor U4351 (N_4351,N_2442,N_2481);
and U4352 (N_4352,N_2979,N_1871);
and U4353 (N_4353,N_2650,N_1683);
and U4354 (N_4354,N_2688,N_1980);
nand U4355 (N_4355,N_2599,N_2254);
nor U4356 (N_4356,N_1638,N_1630);
or U4357 (N_4357,N_1900,N_2353);
or U4358 (N_4358,N_2183,N_1727);
nand U4359 (N_4359,N_1692,N_2157);
nor U4360 (N_4360,N_1679,N_2979);
nor U4361 (N_4361,N_2441,N_2894);
nand U4362 (N_4362,N_2863,N_1533);
nand U4363 (N_4363,N_2981,N_2748);
or U4364 (N_4364,N_1614,N_2154);
nor U4365 (N_4365,N_1952,N_1958);
nand U4366 (N_4366,N_1921,N_2590);
and U4367 (N_4367,N_1583,N_2694);
and U4368 (N_4368,N_2074,N_2735);
nand U4369 (N_4369,N_1502,N_2850);
and U4370 (N_4370,N_2608,N_1866);
or U4371 (N_4371,N_2892,N_2962);
nand U4372 (N_4372,N_2631,N_2679);
xnor U4373 (N_4373,N_1828,N_2770);
nor U4374 (N_4374,N_1872,N_1549);
and U4375 (N_4375,N_1586,N_2706);
or U4376 (N_4376,N_1717,N_1720);
xnor U4377 (N_4377,N_1743,N_2904);
and U4378 (N_4378,N_2835,N_1543);
and U4379 (N_4379,N_2895,N_2575);
and U4380 (N_4380,N_1574,N_2974);
or U4381 (N_4381,N_2508,N_2664);
nor U4382 (N_4382,N_1850,N_2426);
nor U4383 (N_4383,N_1783,N_1838);
or U4384 (N_4384,N_2207,N_1528);
and U4385 (N_4385,N_2051,N_2420);
or U4386 (N_4386,N_2416,N_1985);
nor U4387 (N_4387,N_1648,N_2394);
and U4388 (N_4388,N_2157,N_2465);
and U4389 (N_4389,N_2907,N_2253);
nor U4390 (N_4390,N_1762,N_2744);
nand U4391 (N_4391,N_1942,N_2560);
and U4392 (N_4392,N_2040,N_1583);
or U4393 (N_4393,N_2196,N_2985);
or U4394 (N_4394,N_1746,N_1914);
and U4395 (N_4395,N_2136,N_2127);
nand U4396 (N_4396,N_2395,N_2064);
nor U4397 (N_4397,N_1890,N_2159);
or U4398 (N_4398,N_2947,N_2400);
and U4399 (N_4399,N_2780,N_2952);
xnor U4400 (N_4400,N_2185,N_2136);
xnor U4401 (N_4401,N_1806,N_1656);
or U4402 (N_4402,N_2754,N_2664);
and U4403 (N_4403,N_2891,N_1966);
nand U4404 (N_4404,N_2118,N_1582);
nand U4405 (N_4405,N_1982,N_1535);
nand U4406 (N_4406,N_2058,N_1963);
and U4407 (N_4407,N_2070,N_2889);
or U4408 (N_4408,N_2972,N_2376);
nand U4409 (N_4409,N_2929,N_1731);
or U4410 (N_4410,N_2592,N_1934);
nor U4411 (N_4411,N_2349,N_2534);
and U4412 (N_4412,N_2345,N_1670);
or U4413 (N_4413,N_2053,N_1727);
and U4414 (N_4414,N_1971,N_1529);
xnor U4415 (N_4415,N_2223,N_2146);
and U4416 (N_4416,N_1811,N_2736);
or U4417 (N_4417,N_2352,N_2538);
nand U4418 (N_4418,N_2660,N_2861);
xor U4419 (N_4419,N_2667,N_2287);
nand U4420 (N_4420,N_1873,N_2642);
nor U4421 (N_4421,N_2116,N_1929);
xnor U4422 (N_4422,N_1936,N_1720);
or U4423 (N_4423,N_2148,N_1527);
nor U4424 (N_4424,N_2781,N_2420);
nor U4425 (N_4425,N_1773,N_1963);
and U4426 (N_4426,N_2247,N_1737);
nand U4427 (N_4427,N_2208,N_2212);
or U4428 (N_4428,N_2681,N_1525);
nand U4429 (N_4429,N_2380,N_1580);
xnor U4430 (N_4430,N_2785,N_2300);
nand U4431 (N_4431,N_2060,N_1631);
or U4432 (N_4432,N_1636,N_2062);
and U4433 (N_4433,N_2415,N_2924);
xor U4434 (N_4434,N_2130,N_1981);
xor U4435 (N_4435,N_2617,N_2888);
or U4436 (N_4436,N_2351,N_1509);
and U4437 (N_4437,N_2633,N_2578);
and U4438 (N_4438,N_2332,N_1772);
nor U4439 (N_4439,N_2195,N_1965);
and U4440 (N_4440,N_2857,N_1618);
nand U4441 (N_4441,N_1573,N_2802);
nand U4442 (N_4442,N_2567,N_2397);
nor U4443 (N_4443,N_2740,N_2971);
and U4444 (N_4444,N_2046,N_2073);
nand U4445 (N_4445,N_2320,N_1653);
nand U4446 (N_4446,N_2009,N_1671);
and U4447 (N_4447,N_2830,N_2102);
and U4448 (N_4448,N_2991,N_1590);
or U4449 (N_4449,N_1758,N_2500);
or U4450 (N_4450,N_2104,N_2812);
or U4451 (N_4451,N_2327,N_1530);
and U4452 (N_4452,N_2088,N_1990);
nor U4453 (N_4453,N_1507,N_2731);
or U4454 (N_4454,N_1875,N_2690);
nand U4455 (N_4455,N_2153,N_1766);
and U4456 (N_4456,N_2504,N_2997);
nor U4457 (N_4457,N_2542,N_2905);
or U4458 (N_4458,N_2064,N_1980);
nand U4459 (N_4459,N_2791,N_2268);
xor U4460 (N_4460,N_2170,N_2112);
or U4461 (N_4461,N_1661,N_1581);
and U4462 (N_4462,N_2613,N_1737);
and U4463 (N_4463,N_2249,N_1800);
or U4464 (N_4464,N_1981,N_2381);
nor U4465 (N_4465,N_2767,N_1702);
or U4466 (N_4466,N_2213,N_2310);
or U4467 (N_4467,N_2657,N_2601);
nor U4468 (N_4468,N_2090,N_1687);
or U4469 (N_4469,N_2672,N_2688);
nor U4470 (N_4470,N_2771,N_2673);
nand U4471 (N_4471,N_1506,N_2045);
nand U4472 (N_4472,N_1739,N_2670);
or U4473 (N_4473,N_1890,N_2088);
xor U4474 (N_4474,N_2892,N_2439);
nand U4475 (N_4475,N_1619,N_1812);
nand U4476 (N_4476,N_1698,N_2494);
and U4477 (N_4477,N_2790,N_2859);
nor U4478 (N_4478,N_2452,N_1520);
nand U4479 (N_4479,N_2260,N_2560);
and U4480 (N_4480,N_2880,N_1778);
or U4481 (N_4481,N_2001,N_1831);
or U4482 (N_4482,N_2215,N_2930);
or U4483 (N_4483,N_1722,N_1854);
and U4484 (N_4484,N_1683,N_1814);
or U4485 (N_4485,N_2372,N_2757);
or U4486 (N_4486,N_1662,N_2296);
or U4487 (N_4487,N_2835,N_2793);
or U4488 (N_4488,N_2841,N_2895);
or U4489 (N_4489,N_1882,N_1790);
or U4490 (N_4490,N_1960,N_1833);
nand U4491 (N_4491,N_2299,N_2940);
or U4492 (N_4492,N_2688,N_2401);
nor U4493 (N_4493,N_1794,N_2966);
and U4494 (N_4494,N_2794,N_2091);
and U4495 (N_4495,N_2277,N_2050);
and U4496 (N_4496,N_2329,N_2953);
or U4497 (N_4497,N_2655,N_2302);
or U4498 (N_4498,N_2270,N_2051);
nand U4499 (N_4499,N_2366,N_2612);
and U4500 (N_4500,N_3440,N_4264);
nand U4501 (N_4501,N_4008,N_3928);
nand U4502 (N_4502,N_3313,N_3935);
or U4503 (N_4503,N_4203,N_4184);
or U4504 (N_4504,N_3645,N_3338);
or U4505 (N_4505,N_3770,N_3564);
or U4506 (N_4506,N_4132,N_4430);
or U4507 (N_4507,N_3450,N_3724);
and U4508 (N_4508,N_3815,N_4375);
xor U4509 (N_4509,N_4211,N_3876);
nor U4510 (N_4510,N_4340,N_3755);
nand U4511 (N_4511,N_4077,N_3942);
nor U4512 (N_4512,N_3048,N_3626);
nor U4513 (N_4513,N_3316,N_3256);
nor U4514 (N_4514,N_3831,N_3117);
or U4515 (N_4515,N_3054,N_3053);
or U4516 (N_4516,N_3192,N_3076);
or U4517 (N_4517,N_3540,N_3787);
nand U4518 (N_4518,N_4257,N_3668);
and U4519 (N_4519,N_4293,N_3152);
nand U4520 (N_4520,N_4178,N_3041);
nor U4521 (N_4521,N_4197,N_3940);
xor U4522 (N_4522,N_4338,N_3356);
nor U4523 (N_4523,N_4273,N_3701);
or U4524 (N_4524,N_4170,N_4139);
nor U4525 (N_4525,N_4045,N_4271);
or U4526 (N_4526,N_3678,N_4314);
nand U4527 (N_4527,N_3593,N_3308);
or U4528 (N_4528,N_3469,N_3527);
nand U4529 (N_4529,N_3186,N_4478);
nand U4530 (N_4530,N_4214,N_3400);
or U4531 (N_4531,N_3947,N_3491);
xnor U4532 (N_4532,N_3349,N_4252);
nor U4533 (N_4533,N_3382,N_3855);
and U4534 (N_4534,N_3269,N_3141);
and U4535 (N_4535,N_3811,N_3073);
and U4536 (N_4536,N_3500,N_4244);
nor U4537 (N_4537,N_4133,N_4243);
or U4538 (N_4538,N_3462,N_4018);
or U4539 (N_4539,N_3452,N_4124);
or U4540 (N_4540,N_3096,N_3871);
nor U4541 (N_4541,N_3489,N_4057);
and U4542 (N_4542,N_3771,N_4006);
nor U4543 (N_4543,N_3778,N_4023);
xnor U4544 (N_4544,N_3503,N_3359);
or U4545 (N_4545,N_3704,N_3923);
nor U4546 (N_4546,N_4072,N_3553);
nor U4547 (N_4547,N_3114,N_3348);
and U4548 (N_4548,N_3009,N_3063);
or U4549 (N_4549,N_3894,N_3859);
xnor U4550 (N_4550,N_3213,N_4476);
nand U4551 (N_4551,N_3666,N_3399);
nor U4552 (N_4552,N_4455,N_3994);
xnor U4553 (N_4553,N_4207,N_4377);
or U4554 (N_4554,N_3693,N_3608);
or U4555 (N_4555,N_3837,N_4277);
nand U4556 (N_4556,N_4356,N_4301);
and U4557 (N_4557,N_4471,N_3767);
or U4558 (N_4558,N_3458,N_3106);
nand U4559 (N_4559,N_3421,N_4318);
and U4560 (N_4560,N_4467,N_3765);
and U4561 (N_4561,N_4099,N_3436);
nor U4562 (N_4562,N_3074,N_3371);
nor U4563 (N_4563,N_4287,N_3333);
nor U4564 (N_4564,N_4482,N_4081);
or U4565 (N_4565,N_3861,N_3872);
and U4566 (N_4566,N_4158,N_4262);
and U4567 (N_4567,N_3546,N_3684);
or U4568 (N_4568,N_4283,N_3207);
or U4569 (N_4569,N_4216,N_4009);
nor U4570 (N_4570,N_4113,N_4186);
nor U4571 (N_4571,N_4369,N_3565);
nand U4572 (N_4572,N_3911,N_3146);
and U4573 (N_4573,N_3050,N_3892);
and U4574 (N_4574,N_3818,N_4382);
nand U4575 (N_4575,N_4343,N_3867);
or U4576 (N_4576,N_3548,N_3488);
or U4577 (N_4577,N_4483,N_4332);
or U4578 (N_4578,N_3325,N_3191);
xor U4579 (N_4579,N_3583,N_3844);
nor U4580 (N_4580,N_3560,N_3040);
nor U4581 (N_4581,N_3611,N_4342);
xnor U4582 (N_4582,N_3394,N_3429);
nor U4583 (N_4583,N_3632,N_3554);
and U4584 (N_4584,N_3951,N_3996);
or U4585 (N_4585,N_3949,N_3875);
and U4586 (N_4586,N_4017,N_3671);
nand U4587 (N_4587,N_4224,N_3194);
nand U4588 (N_4588,N_3707,N_4349);
and U4589 (N_4589,N_3957,N_4148);
and U4590 (N_4590,N_3840,N_4457);
nor U4591 (N_4591,N_4151,N_3142);
nand U4592 (N_4592,N_4385,N_3821);
nor U4593 (N_4593,N_3208,N_3024);
nor U4594 (N_4594,N_3910,N_4414);
xor U4595 (N_4595,N_4444,N_4289);
xor U4596 (N_4596,N_3428,N_3100);
or U4597 (N_4597,N_4226,N_3901);
nand U4598 (N_4598,N_3012,N_3884);
nand U4599 (N_4599,N_4095,N_3025);
nor U4600 (N_4600,N_3537,N_3315);
and U4601 (N_4601,N_3927,N_3365);
or U4602 (N_4602,N_4068,N_3786);
nand U4603 (N_4603,N_3902,N_3579);
xnor U4604 (N_4604,N_3918,N_3195);
nand U4605 (N_4605,N_3956,N_3280);
xnor U4606 (N_4606,N_4100,N_3013);
xnor U4607 (N_4607,N_4169,N_3703);
nor U4608 (N_4608,N_4119,N_4067);
nand U4609 (N_4609,N_4347,N_3014);
or U4610 (N_4610,N_3238,N_3418);
nor U4611 (N_4611,N_3022,N_3575);
nand U4612 (N_4612,N_3848,N_4215);
and U4613 (N_4613,N_4034,N_4461);
or U4614 (N_4614,N_3184,N_3622);
nor U4615 (N_4615,N_4429,N_4321);
or U4616 (N_4616,N_3110,N_3478);
and U4617 (N_4617,N_4128,N_4317);
and U4618 (N_4618,N_3895,N_3438);
or U4619 (N_4619,N_4161,N_4115);
and U4620 (N_4620,N_3835,N_4210);
and U4621 (N_4621,N_4070,N_4061);
nand U4622 (N_4622,N_3597,N_3705);
and U4623 (N_4623,N_3079,N_3206);
nand U4624 (N_4624,N_3634,N_3168);
and U4625 (N_4625,N_3392,N_4185);
nor U4626 (N_4626,N_4103,N_3943);
nand U4627 (N_4627,N_4396,N_3713);
nor U4628 (N_4628,N_3799,N_3427);
nor U4629 (N_4629,N_3497,N_4452);
nand U4630 (N_4630,N_3275,N_4263);
or U4631 (N_4631,N_3109,N_3710);
and U4632 (N_4632,N_3538,N_3714);
and U4633 (N_4633,N_3912,N_3588);
nand U4634 (N_4634,N_3619,N_3893);
nand U4635 (N_4635,N_3147,N_3341);
nor U4636 (N_4636,N_3766,N_3793);
or U4637 (N_4637,N_4033,N_3519);
and U4638 (N_4638,N_4098,N_4173);
or U4639 (N_4639,N_3490,N_3264);
and U4640 (N_4640,N_4005,N_4076);
or U4641 (N_4641,N_3285,N_4420);
nor U4642 (N_4642,N_3003,N_4378);
and U4643 (N_4643,N_4145,N_4047);
nor U4644 (N_4644,N_3924,N_3974);
nand U4645 (N_4645,N_4241,N_3986);
nand U4646 (N_4646,N_3143,N_3607);
nand U4647 (N_4647,N_3964,N_4162);
and U4648 (N_4648,N_3946,N_3290);
nand U4649 (N_4649,N_4495,N_4157);
or U4650 (N_4650,N_3144,N_3735);
and U4651 (N_4651,N_3753,N_3828);
or U4652 (N_4652,N_4167,N_4362);
or U4653 (N_4653,N_3993,N_4472);
or U4654 (N_4654,N_3202,N_4104);
nand U4655 (N_4655,N_4431,N_3788);
nand U4656 (N_4656,N_4065,N_3047);
nor U4657 (N_4657,N_3200,N_3153);
nand U4658 (N_4658,N_4451,N_4279);
or U4659 (N_4659,N_4160,N_3650);
and U4660 (N_4660,N_3448,N_3406);
nor U4661 (N_4661,N_3062,N_4330);
nor U4662 (N_4662,N_3921,N_3419);
xor U4663 (N_4663,N_3329,N_4380);
or U4664 (N_4664,N_3312,N_3915);
xor U4665 (N_4665,N_3457,N_3355);
nor U4666 (N_4666,N_3598,N_3283);
or U4667 (N_4667,N_3995,N_3535);
nand U4668 (N_4668,N_3610,N_4353);
and U4669 (N_4669,N_3485,N_3870);
nor U4670 (N_4670,N_4415,N_3299);
nor U4671 (N_4671,N_4080,N_3060);
or U4672 (N_4672,N_4155,N_4280);
or U4673 (N_4673,N_3865,N_4029);
or U4674 (N_4674,N_4274,N_4202);
nand U4675 (N_4675,N_3987,N_4335);
nand U4676 (N_4676,N_3220,N_4439);
xor U4677 (N_4677,N_4064,N_3412);
nand U4678 (N_4678,N_3107,N_3101);
or U4679 (N_4679,N_3730,N_3813);
or U4680 (N_4680,N_3112,N_3609);
and U4681 (N_4681,N_3732,N_3768);
nand U4682 (N_4682,N_3653,N_4046);
and U4683 (N_4683,N_3643,N_4013);
and U4684 (N_4684,N_3706,N_4464);
xnor U4685 (N_4685,N_3128,N_4019);
nand U4686 (N_4686,N_4110,N_3344);
nor U4687 (N_4687,N_4078,N_3629);
or U4688 (N_4688,N_3763,N_3690);
nor U4689 (N_4689,N_3027,N_3277);
xnor U4690 (N_4690,N_3644,N_3046);
or U4691 (N_4691,N_4101,N_4494);
nor U4692 (N_4692,N_3725,N_3375);
nor U4693 (N_4693,N_3646,N_3068);
and U4694 (N_4694,N_3850,N_3081);
nor U4695 (N_4695,N_4384,N_3601);
nor U4696 (N_4696,N_4003,N_4260);
nand U4697 (N_4697,N_3236,N_3196);
nor U4698 (N_4698,N_3467,N_4020);
and U4699 (N_4699,N_4350,N_3989);
xnor U4700 (N_4700,N_3403,N_3148);
nor U4701 (N_4701,N_4091,N_3094);
nor U4702 (N_4702,N_3878,N_3209);
and U4703 (N_4703,N_3245,N_3336);
and U4704 (N_4704,N_3664,N_4193);
nor U4705 (N_4705,N_4278,N_3604);
or U4706 (N_4706,N_3019,N_4305);
and U4707 (N_4707,N_3465,N_4038);
nand U4708 (N_4708,N_3669,N_3252);
nand U4709 (N_4709,N_3391,N_3139);
nand U4710 (N_4710,N_4194,N_4363);
nor U4711 (N_4711,N_3905,N_3098);
nor U4712 (N_4712,N_3332,N_3929);
nor U4713 (N_4713,N_4427,N_3323);
nor U4714 (N_4714,N_3971,N_3635);
xor U4715 (N_4715,N_4135,N_3441);
or U4716 (N_4716,N_3606,N_4147);
nor U4717 (N_4717,N_3775,N_4354);
and U4718 (N_4718,N_4176,N_3749);
or U4719 (N_4719,N_4021,N_4179);
nand U4720 (N_4720,N_3145,N_3791);
nor U4721 (N_4721,N_3476,N_4052);
nor U4722 (N_4722,N_3843,N_4223);
and U4723 (N_4723,N_4297,N_3164);
or U4724 (N_4724,N_4131,N_3108);
and U4725 (N_4725,N_3381,N_3086);
or U4726 (N_4726,N_4154,N_3018);
nor U4727 (N_4727,N_3237,N_3080);
and U4728 (N_4728,N_3230,N_3930);
and U4729 (N_4729,N_3259,N_3157);
nand U4730 (N_4730,N_3804,N_3590);
and U4731 (N_4731,N_3459,N_4242);
and U4732 (N_4732,N_3720,N_3033);
nor U4733 (N_4733,N_4355,N_3055);
and U4734 (N_4734,N_3756,N_3530);
nor U4735 (N_4735,N_3342,N_4367);
or U4736 (N_4736,N_4421,N_4360);
nor U4737 (N_4737,N_3827,N_3722);
nand U4738 (N_4738,N_3944,N_4393);
xnor U4739 (N_4739,N_4105,N_4090);
nand U4740 (N_4740,N_3816,N_3132);
and U4741 (N_4741,N_3834,N_3135);
xor U4742 (N_4742,N_3812,N_4399);
nor U4743 (N_4743,N_3558,N_4308);
or U4744 (N_4744,N_3838,N_3075);
and U4745 (N_4745,N_3008,N_3853);
and U4746 (N_4746,N_4097,N_3302);
nand U4747 (N_4747,N_3454,N_3512);
nor U4748 (N_4748,N_4372,N_4424);
nand U4749 (N_4749,N_3973,N_3176);
or U4750 (N_4750,N_3842,N_3574);
or U4751 (N_4751,N_3633,N_3303);
xor U4752 (N_4752,N_3326,N_3941);
and U4753 (N_4753,N_4007,N_3413);
nand U4754 (N_4754,N_3700,N_3197);
and U4755 (N_4755,N_4359,N_3493);
and U4756 (N_4756,N_4422,N_3455);
nand U4757 (N_4757,N_3000,N_3115);
nor U4758 (N_4758,N_3781,N_3832);
nor U4759 (N_4759,N_3387,N_4345);
nand U4760 (N_4760,N_3204,N_3199);
or U4761 (N_4761,N_3102,N_4298);
and U4762 (N_4762,N_3300,N_4351);
nor U4763 (N_4763,N_3695,N_3249);
and U4764 (N_4764,N_3233,N_3021);
or U4765 (N_4765,N_4171,N_3628);
and U4766 (N_4766,N_3092,N_4204);
nor U4767 (N_4767,N_4085,N_3950);
and U4768 (N_4768,N_4428,N_4096);
and U4769 (N_4769,N_3211,N_4475);
and U4770 (N_4770,N_3405,N_4190);
nor U4771 (N_4771,N_4329,N_3777);
or U4772 (N_4772,N_3226,N_4291);
nor U4773 (N_4773,N_4086,N_4470);
and U4774 (N_4774,N_3331,N_4499);
nor U4775 (N_4775,N_3396,N_4434);
or U4776 (N_4776,N_3594,N_3223);
nor U4777 (N_4777,N_4408,N_4391);
and U4778 (N_4778,N_3550,N_4447);
or U4779 (N_4779,N_4153,N_3502);
nor U4780 (N_4780,N_3566,N_3289);
nand U4781 (N_4781,N_3773,N_3327);
nand U4782 (N_4782,N_4348,N_4022);
xor U4783 (N_4783,N_3116,N_4395);
and U4784 (N_4784,N_4016,N_3402);
nor U4785 (N_4785,N_4480,N_3393);
xnor U4786 (N_4786,N_4358,N_3087);
or U4787 (N_4787,N_3728,N_3212);
or U4788 (N_4788,N_4460,N_4336);
or U4789 (N_4789,N_3011,N_3287);
nand U4790 (N_4790,N_4331,N_3415);
xor U4791 (N_4791,N_4235,N_3292);
and U4792 (N_4792,N_3711,N_3174);
nand U4793 (N_4793,N_3833,N_3939);
xnor U4794 (N_4794,N_4055,N_3802);
and U4795 (N_4795,N_4328,N_4056);
or U4796 (N_4796,N_4473,N_3625);
xnor U4797 (N_4797,N_3203,N_3061);
and U4798 (N_4798,N_4032,N_3888);
xor U4799 (N_4799,N_3661,N_3699);
nand U4800 (N_4800,N_3885,N_3297);
or U4801 (N_4801,N_3473,N_3555);
or U4802 (N_4802,N_4443,N_3506);
nor U4803 (N_4803,N_4163,N_3499);
and U4804 (N_4804,N_3999,N_4276);
or U4805 (N_4805,N_4387,N_3284);
or U4806 (N_4806,N_4191,N_3346);
nand U4807 (N_4807,N_3273,N_3260);
xor U4808 (N_4808,N_3907,N_3719);
nand U4809 (N_4809,N_4028,N_4140);
xnor U4810 (N_4810,N_4334,N_3983);
nor U4811 (N_4811,N_3547,N_4142);
or U4812 (N_4812,N_3004,N_3595);
and U4813 (N_4813,N_3568,N_4489);
nor U4814 (N_4814,N_3980,N_4322);
and U4815 (N_4815,N_3761,N_3914);
and U4816 (N_4816,N_3623,N_4364);
and U4817 (N_4817,N_3819,N_3696);
xnor U4818 (N_4818,N_4491,N_4165);
nor U4819 (N_4819,N_3352,N_3305);
and U4820 (N_4820,N_4062,N_3976);
nand U4821 (N_4821,N_3651,N_3536);
nand U4822 (N_4822,N_3288,N_4042);
or U4823 (N_4823,N_3686,N_3444);
or U4824 (N_4824,N_3747,N_4498);
or U4825 (N_4825,N_3077,N_3829);
nand U4826 (N_4826,N_3970,N_3361);
or U4827 (N_4827,N_3580,N_3680);
nand U4828 (N_4828,N_3962,N_4088);
nand U4829 (N_4829,N_3126,N_3582);
and U4830 (N_4830,N_3071,N_3961);
xnor U4831 (N_4831,N_3059,N_3231);
or U4832 (N_4832,N_4337,N_4462);
and U4833 (N_4833,N_3742,N_4406);
nand U4834 (N_4834,N_4156,N_3266);
nor U4835 (N_4835,N_3716,N_3453);
xor U4836 (N_4836,N_3800,N_3932);
nor U4837 (N_4837,N_3328,N_3420);
xor U4838 (N_4838,N_3909,N_4423);
nor U4839 (N_4839,N_4199,N_3692);
and U4840 (N_4840,N_4379,N_4180);
and U4841 (N_4841,N_4219,N_3304);
xor U4842 (N_4842,N_3374,N_3743);
nor U4843 (N_4843,N_3681,N_3534);
or U4844 (N_4844,N_4388,N_3529);
nor U4845 (N_4845,N_3250,N_3006);
nor U4846 (N_4846,N_3082,N_3868);
nand U4847 (N_4847,N_3267,N_3470);
or U4848 (N_4848,N_3464,N_3272);
and U4849 (N_4849,N_3521,N_3282);
xnor U4850 (N_4850,N_3841,N_3805);
nand U4851 (N_4851,N_4239,N_3298);
xor U4852 (N_4852,N_4383,N_3596);
xnor U4853 (N_4853,N_3642,N_3125);
and U4854 (N_4854,N_3442,N_3744);
xor U4855 (N_4855,N_3404,N_4466);
and U4856 (N_4856,N_3494,N_4270);
nor U4857 (N_4857,N_4325,N_3750);
nand U4858 (N_4858,N_3172,N_3072);
xor U4859 (N_4859,N_3005,N_4282);
or U4860 (N_4860,N_4401,N_4295);
or U4861 (N_4861,N_4411,N_3291);
or U4862 (N_4862,N_3789,N_4175);
and U4863 (N_4863,N_3416,N_4146);
nor U4864 (N_4864,N_3830,N_3443);
nand U4865 (N_4865,N_3067,N_3549);
xor U4866 (N_4866,N_3605,N_3158);
and U4867 (N_4867,N_3070,N_4053);
nand U4868 (N_4868,N_3010,N_3095);
or U4869 (N_4869,N_3599,N_4143);
or U4870 (N_4870,N_4370,N_3384);
nand U4871 (N_4871,N_4181,N_3614);
nor U4872 (N_4872,N_3702,N_3903);
and U4873 (N_4873,N_3543,N_3822);
or U4874 (N_4874,N_4392,N_3638);
or U4875 (N_4875,N_3592,N_4134);
and U4876 (N_4876,N_3603,N_3159);
nor U4877 (N_4877,N_3150,N_3891);
nand U4878 (N_4878,N_3665,N_3417);
nor U4879 (N_4879,N_3218,N_3089);
and U4880 (N_4880,N_3118,N_3475);
nor U4881 (N_4881,N_4413,N_4248);
nor U4882 (N_4882,N_4454,N_3562);
or U4883 (N_4883,N_4126,N_4082);
nor U4884 (N_4884,N_4094,N_3262);
or U4885 (N_4885,N_3044,N_3103);
nand U4886 (N_4886,N_4268,N_3339);
and U4887 (N_4887,N_4381,N_3990);
nand U4888 (N_4888,N_3477,N_4118);
or U4889 (N_4889,N_3487,N_3340);
and U4890 (N_4890,N_3439,N_3410);
xnor U4891 (N_4891,N_3078,N_3551);
nand U4892 (N_4892,N_3123,N_3613);
nor U4893 (N_4893,N_3065,N_4121);
nor U4894 (N_4894,N_4409,N_3655);
or U4895 (N_4895,N_3351,N_3869);
nand U4896 (N_4896,N_3296,N_3557);
nand U4897 (N_4897,N_3151,N_4299);
nor U4898 (N_4898,N_3414,N_4366);
and U4899 (N_4899,N_3461,N_3890);
or U4900 (N_4900,N_4002,N_3407);
nor U4901 (N_4901,N_3636,N_4405);
and U4902 (N_4902,N_3779,N_3317);
nand U4903 (N_4903,N_3149,N_3959);
nor U4904 (N_4904,N_3177,N_3463);
nand U4905 (N_4905,N_4357,N_3322);
nor U4906 (N_4906,N_3774,N_3481);
xor U4907 (N_4907,N_3227,N_3066);
nand U4908 (N_4908,N_3790,N_3193);
nor U4909 (N_4909,N_3175,N_3803);
and U4910 (N_4910,N_3105,N_3028);
and U4911 (N_4911,N_3225,N_3796);
nor U4912 (N_4912,N_3119,N_3166);
nor U4913 (N_4913,N_3247,N_4373);
or U4914 (N_4914,N_3372,N_4217);
or U4915 (N_4915,N_4228,N_3745);
or U4916 (N_4916,N_3764,N_4001);
nor U4917 (N_4917,N_3472,N_3657);
and U4918 (N_4918,N_3754,N_4221);
or U4919 (N_4919,N_3785,N_4326);
xor U4920 (N_4920,N_3577,N_3694);
nand U4921 (N_4921,N_3131,N_4416);
or U4922 (N_4922,N_3898,N_3882);
nor U4923 (N_4923,N_3663,N_3368);
and U4924 (N_4924,N_4041,N_3511);
or U4925 (N_4925,N_3165,N_4313);
xor U4926 (N_4926,N_4265,N_4106);
xnor U4927 (N_4927,N_3294,N_3656);
nor U4928 (N_4928,N_3992,N_3931);
nand U4929 (N_4929,N_3659,N_4039);
or U4930 (N_4930,N_4043,N_3385);
nor U4931 (N_4931,N_4316,N_4075);
nand U4932 (N_4932,N_4168,N_3293);
or U4933 (N_4933,N_3845,N_3170);
and U4934 (N_4934,N_3121,N_3255);
and U4935 (N_4935,N_4227,N_4344);
or U4936 (N_4936,N_3689,N_3520);
or U4937 (N_4937,N_3712,N_3569);
nor U4938 (N_4938,N_3883,N_3229);
or U4939 (N_4939,N_3591,N_4407);
xor U4940 (N_4940,N_3430,N_3997);
and U4941 (N_4941,N_4187,N_4024);
nand U4942 (N_4942,N_4398,N_3449);
xor U4943 (N_4943,N_4196,N_3030);
nor U4944 (N_4944,N_4333,N_3737);
xnor U4945 (N_4945,N_3683,N_3167);
nor U4946 (N_4946,N_3654,N_4102);
and U4947 (N_4947,N_4137,N_4084);
nand U4948 (N_4948,N_3134,N_3492);
nor U4949 (N_4949,N_4304,N_3254);
nor U4950 (N_4950,N_3451,N_4069);
and U4951 (N_4951,N_3278,N_4208);
nor U4952 (N_4952,N_3542,N_3357);
nor U4953 (N_4953,N_3007,N_3858);
and U4954 (N_4954,N_3045,N_4481);
nand U4955 (N_4955,N_4138,N_3064);
nand U4956 (N_4956,N_3408,N_3090);
and U4957 (N_4957,N_4025,N_3274);
and U4958 (N_4958,N_3846,N_3740);
and U4959 (N_4959,N_3515,N_3647);
nand U4960 (N_4960,N_3688,N_3034);
and U4961 (N_4961,N_3508,N_3482);
and U4962 (N_4962,N_3977,N_4073);
nor U4963 (N_4963,N_4292,N_3241);
and U4964 (N_4964,N_3938,N_3866);
nor U4965 (N_4965,N_3364,N_4129);
and U4966 (N_4966,N_4486,N_3251);
and U4967 (N_4967,N_3504,N_3897);
nand U4968 (N_4968,N_4339,N_3736);
nand U4969 (N_4969,N_3434,N_4266);
xor U4970 (N_4970,N_4015,N_4250);
and U4971 (N_4971,N_4122,N_3792);
nor U4972 (N_4972,N_3585,N_3026);
or U4973 (N_4973,N_3906,N_3801);
or U4974 (N_4974,N_4000,N_4327);
nor U4975 (N_4975,N_3425,N_4259);
nand U4976 (N_4976,N_3752,N_3637);
xnor U4977 (N_4977,N_3401,N_3358);
or U4978 (N_4978,N_3602,N_3670);
nand U4979 (N_4979,N_4492,N_3154);
or U4980 (N_4980,N_4164,N_3432);
or U4981 (N_4981,N_3780,N_4272);
nor U4982 (N_4982,N_3916,N_3017);
or U4983 (N_4983,N_3757,N_3038);
nor U4984 (N_4984,N_3738,N_4352);
nand U4985 (N_4985,N_4432,N_3232);
or U4986 (N_4986,N_3035,N_3390);
nand U4987 (N_4987,N_4437,N_3161);
nand U4988 (N_4988,N_4141,N_3945);
nand U4989 (N_4989,N_4425,N_4083);
and U4990 (N_4990,N_4400,N_3222);
xnor U4991 (N_4991,N_3395,N_3919);
or U4992 (N_4992,N_4111,N_3137);
and U4993 (N_4993,N_4306,N_3854);
nor U4994 (N_4994,N_3741,N_3426);
or U4995 (N_4995,N_3509,N_3133);
and U4996 (N_4996,N_3483,N_3171);
nand U4997 (N_4997,N_3963,N_4296);
nand U4998 (N_4998,N_3960,N_4284);
nand U4999 (N_4999,N_3968,N_4037);
nor U5000 (N_5000,N_4403,N_3772);
nor U5001 (N_5001,N_3486,N_3474);
or U5002 (N_5002,N_3198,N_3660);
nand U5003 (N_5003,N_4275,N_3379);
and U5004 (N_5004,N_3917,N_4249);
nand U5005 (N_5005,N_3263,N_3571);
and U5006 (N_5006,N_3958,N_3836);
or U5007 (N_5007,N_3388,N_4130);
nand U5008 (N_5008,N_3985,N_4397);
nor U5009 (N_5009,N_3039,N_4440);
nand U5010 (N_5010,N_3518,N_3697);
nand U5011 (N_5011,N_3015,N_3691);
nor U5012 (N_5012,N_3334,N_3268);
or U5013 (N_5013,N_4234,N_3445);
xnor U5014 (N_5014,N_3839,N_3934);
nor U5015 (N_5015,N_4426,N_3373);
or U5016 (N_5016,N_4035,N_4433);
xor U5017 (N_5017,N_4256,N_4004);
nor U5018 (N_5018,N_3221,N_4307);
and U5019 (N_5019,N_3526,N_3016);
nor U5020 (N_5020,N_3517,N_3466);
nor U5021 (N_5021,N_3219,N_3514);
or U5022 (N_5022,N_4449,N_3649);
xnor U5023 (N_5023,N_4269,N_3362);
nand U5024 (N_5024,N_3496,N_3672);
and U5025 (N_5025,N_4490,N_3925);
and U5026 (N_5026,N_3877,N_4183);
nand U5027 (N_5027,N_3814,N_3573);
nand U5028 (N_5028,N_3718,N_4189);
or U5029 (N_5029,N_3169,N_3544);
and U5030 (N_5030,N_3784,N_3782);
nor U5031 (N_5031,N_3320,N_3817);
and U5032 (N_5032,N_3952,N_3138);
nor U5033 (N_5033,N_4198,N_4152);
nor U5034 (N_5034,N_3337,N_3377);
or U5035 (N_5035,N_3510,N_4365);
and U5036 (N_5036,N_3658,N_3431);
nand U5037 (N_5037,N_3798,N_3258);
and U5038 (N_5038,N_3127,N_4442);
nand U5039 (N_5039,N_4071,N_3424);
nor U5040 (N_5040,N_3933,N_3129);
nand U5041 (N_5041,N_3624,N_4232);
xnor U5042 (N_5042,N_4031,N_4112);
nand U5043 (N_5043,N_3343,N_3920);
xnor U5044 (N_5044,N_3318,N_3052);
or U5045 (N_5045,N_3099,N_3495);
or U5046 (N_5046,N_4496,N_3386);
or U5047 (N_5047,N_4310,N_3776);
nor U5048 (N_5048,N_3279,N_3366);
nor U5049 (N_5049,N_3746,N_3242);
xor U5050 (N_5050,N_4441,N_3324);
and U5051 (N_5051,N_3335,N_4485);
nor U5052 (N_5052,N_4222,N_3246);
nand U5053 (N_5053,N_4311,N_4201);
or U5054 (N_5054,N_4346,N_4240);
nor U5055 (N_5055,N_4477,N_4127);
or U5056 (N_5056,N_3345,N_4074);
or U5057 (N_5057,N_4488,N_4066);
nand U5058 (N_5058,N_3797,N_3029);
or U5059 (N_5059,N_3734,N_3201);
or U5060 (N_5060,N_3908,N_3130);
nor U5061 (N_5061,N_3097,N_3541);
and U5062 (N_5062,N_3215,N_4079);
nor U5063 (N_5063,N_4469,N_3111);
nor U5064 (N_5064,N_3570,N_3600);
nor U5065 (N_5065,N_3572,N_4254);
nor U5066 (N_5066,N_3618,N_4300);
xnor U5067 (N_5067,N_3966,N_3760);
or U5068 (N_5068,N_4238,N_3446);
and U5069 (N_5069,N_3673,N_3674);
xor U5070 (N_5070,N_4247,N_3295);
nand U5071 (N_5071,N_3433,N_3378);
or U5072 (N_5072,N_4309,N_3733);
nor U5073 (N_5073,N_3620,N_3723);
nor U5074 (N_5074,N_3809,N_3460);
and U5075 (N_5075,N_3667,N_3383);
nand U5076 (N_5076,N_3376,N_3860);
nor U5077 (N_5077,N_3874,N_4174);
and U5078 (N_5078,N_4063,N_3709);
nor U5079 (N_5079,N_3857,N_4150);
or U5080 (N_5080,N_3042,N_3234);
xnor U5081 (N_5081,N_3528,N_3567);
and U5082 (N_5082,N_3679,N_3310);
and U5083 (N_5083,N_3615,N_3001);
nor U5084 (N_5084,N_3422,N_4177);
nor U5085 (N_5085,N_3759,N_3120);
and U5086 (N_5086,N_4195,N_4220);
or U5087 (N_5087,N_3978,N_4446);
nor U5088 (N_5088,N_3975,N_4484);
or U5089 (N_5089,N_3825,N_4450);
and U5090 (N_5090,N_4059,N_3584);
and U5091 (N_5091,N_3479,N_3367);
and U5092 (N_5092,N_4054,N_4012);
nand U5093 (N_5093,N_3953,N_4014);
or U5094 (N_5094,N_3253,N_3826);
and U5095 (N_5095,N_3214,N_3794);
or U5096 (N_5096,N_4109,N_3397);
nor U5097 (N_5097,N_3456,N_4117);
and U5098 (N_5098,N_4120,N_3281);
and U5099 (N_5099,N_3676,N_4246);
nor U5100 (N_5100,N_4051,N_4465);
or U5101 (N_5101,N_3155,N_4026);
nor U5102 (N_5102,N_4319,N_3190);
nand U5103 (N_5103,N_3437,N_4192);
or U5104 (N_5104,N_3612,N_4285);
and U5105 (N_5105,N_3271,N_3988);
nand U5106 (N_5106,N_3899,N_3856);
xor U5107 (N_5107,N_4458,N_4182);
nand U5108 (N_5108,N_3887,N_3363);
nand U5109 (N_5109,N_3900,N_3484);
and U5110 (N_5110,N_4114,N_3758);
or U5111 (N_5111,N_3187,N_4323);
or U5112 (N_5112,N_3808,N_4493);
xor U5113 (N_5113,N_3423,N_3183);
nand U5114 (N_5114,N_4412,N_4011);
and U5115 (N_5115,N_4136,N_4368);
or U5116 (N_5116,N_3981,N_3880);
and U5117 (N_5117,N_4027,N_3820);
or U5118 (N_5118,N_3717,N_4233);
and U5119 (N_5119,N_4361,N_3370);
nand U5120 (N_5120,N_4225,N_3049);
and U5121 (N_5121,N_3217,N_3389);
nand U5122 (N_5122,N_3954,N_3889);
nor U5123 (N_5123,N_4230,N_3104);
and U5124 (N_5124,N_4116,N_3851);
and U5125 (N_5125,N_3330,N_4288);
nand U5126 (N_5126,N_3156,N_3522);
nand U5127 (N_5127,N_3863,N_3685);
xnor U5128 (N_5128,N_3698,N_3913);
or U5129 (N_5129,N_3721,N_4213);
nand U5130 (N_5130,N_4468,N_3056);
xnor U5131 (N_5131,N_3824,N_3524);
and U5132 (N_5132,N_3037,N_3180);
or U5133 (N_5133,N_4341,N_3085);
nand U5134 (N_5134,N_4402,N_3307);
nand U5135 (N_5135,N_3556,N_3057);
or U5136 (N_5136,N_4404,N_3984);
nand U5137 (N_5137,N_3471,N_3552);
nor U5138 (N_5138,N_4459,N_3354);
xnor U5139 (N_5139,N_3682,N_3023);
and U5140 (N_5140,N_3729,N_3586);
and U5141 (N_5141,N_4302,N_3523);
nand U5142 (N_5142,N_3675,N_3727);
and U5143 (N_5143,N_3380,N_4389);
nor U5144 (N_5144,N_3687,N_3173);
or U5145 (N_5145,N_3587,N_4453);
xor U5146 (N_5146,N_3178,N_3873);
or U5147 (N_5147,N_3309,N_3228);
xnor U5148 (N_5148,N_4417,N_3998);
and U5149 (N_5149,N_3480,N_3864);
nor U5150 (N_5150,N_3043,N_4089);
nor U5151 (N_5151,N_3533,N_3020);
or U5152 (N_5152,N_3113,N_3648);
nor U5153 (N_5153,N_3937,N_3265);
or U5154 (N_5154,N_4060,N_4324);
or U5155 (N_5155,N_4386,N_3616);
nand U5156 (N_5156,N_3181,N_3058);
nand U5157 (N_5157,N_3160,N_3353);
nor U5158 (N_5158,N_3576,N_3969);
nor U5159 (N_5159,N_4231,N_3806);
nand U5160 (N_5160,N_4087,N_3091);
or U5161 (N_5161,N_4144,N_3505);
nor U5162 (N_5162,N_4281,N_3581);
nand U5163 (N_5163,N_3239,N_3276);
nand U5164 (N_5164,N_3715,N_3398);
nand U5165 (N_5165,N_3731,N_3748);
nor U5166 (N_5166,N_4236,N_3036);
nor U5167 (N_5167,N_3224,N_3631);
xnor U5168 (N_5168,N_3306,N_3140);
or U5169 (N_5169,N_3002,N_4229);
nand U5170 (N_5170,N_4479,N_4205);
nand U5171 (N_5171,N_4371,N_3124);
nor U5172 (N_5172,N_3189,N_3862);
nor U5173 (N_5173,N_3849,N_4294);
nand U5174 (N_5174,N_3350,N_4108);
and U5175 (N_5175,N_4487,N_3621);
nor U5176 (N_5176,N_3216,N_3409);
nor U5177 (N_5177,N_3726,N_3708);
nand U5178 (N_5178,N_4058,N_3769);
and U5179 (N_5179,N_3617,N_4092);
xnor U5180 (N_5180,N_3922,N_3301);
xnor U5181 (N_5181,N_4286,N_4315);
nand U5182 (N_5182,N_4463,N_3563);
nand U5183 (N_5183,N_3051,N_3852);
or U5184 (N_5184,N_3513,N_4188);
xor U5185 (N_5185,N_3369,N_4376);
nor U5186 (N_5186,N_4445,N_3032);
xnor U5187 (N_5187,N_3321,N_4125);
nor U5188 (N_5188,N_3501,N_3532);
or U5189 (N_5189,N_4049,N_3311);
xor U5190 (N_5190,N_3179,N_3795);
nand U5191 (N_5191,N_3347,N_4390);
or U5192 (N_5192,N_3240,N_3539);
nor U5193 (N_5193,N_3411,N_3188);
nor U5194 (N_5194,N_4253,N_3243);
nor U5195 (N_5195,N_3991,N_3069);
xnor U5196 (N_5196,N_4107,N_3435);
or U5197 (N_5197,N_3677,N_3589);
nor U5198 (N_5198,N_3525,N_3088);
and U5199 (N_5199,N_3639,N_4267);
nand U5200 (N_5200,N_3531,N_3641);
nor U5201 (N_5201,N_4435,N_3904);
and U5202 (N_5202,N_3972,N_3210);
xnor U5203 (N_5203,N_4374,N_3662);
and U5204 (N_5204,N_3948,N_3965);
nor U5205 (N_5205,N_4251,N_4209);
or U5206 (N_5206,N_4212,N_4200);
nor U5207 (N_5207,N_4172,N_4438);
or U5208 (N_5208,N_3652,N_4448);
and U5209 (N_5209,N_4312,N_3979);
or U5210 (N_5210,N_3468,N_3561);
nor U5211 (N_5211,N_3084,N_3936);
or U5212 (N_5212,N_4436,N_3270);
or U5213 (N_5213,N_3762,N_3447);
or U5214 (N_5214,N_3185,N_3360);
or U5215 (N_5215,N_3926,N_3205);
nor U5216 (N_5216,N_3516,N_3982);
and U5217 (N_5217,N_3498,N_4456);
nand U5218 (N_5218,N_3955,N_4474);
or U5219 (N_5219,N_3627,N_3881);
nor U5220 (N_5220,N_3640,N_3244);
nand U5221 (N_5221,N_3182,N_4255);
xor U5222 (N_5222,N_4258,N_3031);
nor U5223 (N_5223,N_4320,N_4497);
nand U5224 (N_5224,N_4410,N_4030);
or U5225 (N_5225,N_3823,N_3559);
nor U5226 (N_5226,N_3286,N_4149);
nand U5227 (N_5227,N_3879,N_3578);
and U5228 (N_5228,N_4010,N_4093);
and U5229 (N_5229,N_3545,N_4237);
nor U5230 (N_5230,N_4303,N_3122);
or U5231 (N_5231,N_4218,N_3319);
nand U5232 (N_5232,N_4206,N_4048);
or U5233 (N_5233,N_4166,N_3136);
or U5234 (N_5234,N_4123,N_4044);
and U5235 (N_5235,N_4245,N_4036);
and U5236 (N_5236,N_3967,N_4040);
nand U5237 (N_5237,N_3810,N_4159);
and U5238 (N_5238,N_3507,N_4050);
and U5239 (N_5239,N_3739,N_3314);
or U5240 (N_5240,N_3630,N_3886);
or U5241 (N_5241,N_3083,N_3257);
and U5242 (N_5242,N_3847,N_3896);
nand U5243 (N_5243,N_4394,N_4419);
nor U5244 (N_5244,N_3751,N_3162);
nand U5245 (N_5245,N_4261,N_3783);
nor U5246 (N_5246,N_4418,N_3093);
and U5247 (N_5247,N_3261,N_3235);
and U5248 (N_5248,N_3163,N_3248);
or U5249 (N_5249,N_4290,N_3807);
nor U5250 (N_5250,N_4347,N_3287);
nor U5251 (N_5251,N_3501,N_3592);
or U5252 (N_5252,N_4498,N_3036);
nand U5253 (N_5253,N_4327,N_4271);
nand U5254 (N_5254,N_3690,N_3555);
and U5255 (N_5255,N_3662,N_4435);
and U5256 (N_5256,N_3928,N_3709);
nor U5257 (N_5257,N_4350,N_3711);
or U5258 (N_5258,N_4185,N_3994);
or U5259 (N_5259,N_3300,N_4474);
and U5260 (N_5260,N_3673,N_3496);
and U5261 (N_5261,N_3000,N_3518);
nor U5262 (N_5262,N_3433,N_3516);
and U5263 (N_5263,N_3931,N_3377);
nand U5264 (N_5264,N_3134,N_3887);
nor U5265 (N_5265,N_3390,N_3221);
or U5266 (N_5266,N_4247,N_3697);
nor U5267 (N_5267,N_3193,N_4333);
nand U5268 (N_5268,N_3469,N_3515);
and U5269 (N_5269,N_3183,N_3874);
nand U5270 (N_5270,N_3875,N_4452);
nand U5271 (N_5271,N_4495,N_3503);
or U5272 (N_5272,N_3511,N_4385);
nor U5273 (N_5273,N_3943,N_4226);
or U5274 (N_5274,N_3354,N_4273);
or U5275 (N_5275,N_3511,N_4446);
nor U5276 (N_5276,N_3400,N_3413);
nand U5277 (N_5277,N_4345,N_4047);
or U5278 (N_5278,N_3129,N_3130);
nor U5279 (N_5279,N_4188,N_3974);
or U5280 (N_5280,N_3627,N_3283);
and U5281 (N_5281,N_4177,N_4309);
nor U5282 (N_5282,N_3375,N_3098);
and U5283 (N_5283,N_3452,N_3986);
and U5284 (N_5284,N_3078,N_3339);
nor U5285 (N_5285,N_3052,N_3669);
xnor U5286 (N_5286,N_4360,N_3355);
nand U5287 (N_5287,N_3261,N_3830);
xor U5288 (N_5288,N_3211,N_3916);
nor U5289 (N_5289,N_3624,N_3538);
or U5290 (N_5290,N_4146,N_3863);
or U5291 (N_5291,N_3421,N_3132);
and U5292 (N_5292,N_3819,N_3981);
nor U5293 (N_5293,N_3769,N_4118);
nor U5294 (N_5294,N_3115,N_3622);
nor U5295 (N_5295,N_3357,N_3563);
nand U5296 (N_5296,N_4389,N_4421);
nand U5297 (N_5297,N_3227,N_3635);
nor U5298 (N_5298,N_3660,N_3845);
nand U5299 (N_5299,N_3536,N_3952);
and U5300 (N_5300,N_3215,N_3870);
or U5301 (N_5301,N_4162,N_4124);
nand U5302 (N_5302,N_3103,N_3902);
nand U5303 (N_5303,N_3929,N_4327);
nor U5304 (N_5304,N_4085,N_4226);
and U5305 (N_5305,N_3766,N_3871);
or U5306 (N_5306,N_3580,N_3239);
nand U5307 (N_5307,N_3705,N_4078);
nand U5308 (N_5308,N_4317,N_3978);
nor U5309 (N_5309,N_3238,N_3780);
nor U5310 (N_5310,N_3871,N_4312);
and U5311 (N_5311,N_3842,N_3196);
xnor U5312 (N_5312,N_4297,N_3122);
or U5313 (N_5313,N_3649,N_4104);
nor U5314 (N_5314,N_3151,N_3557);
or U5315 (N_5315,N_3009,N_3523);
nor U5316 (N_5316,N_4408,N_3753);
or U5317 (N_5317,N_3205,N_4039);
nand U5318 (N_5318,N_3440,N_4341);
nor U5319 (N_5319,N_3360,N_3689);
and U5320 (N_5320,N_3356,N_3141);
nand U5321 (N_5321,N_4167,N_4356);
or U5322 (N_5322,N_3127,N_3645);
and U5323 (N_5323,N_4347,N_4251);
and U5324 (N_5324,N_4412,N_3903);
or U5325 (N_5325,N_3253,N_3100);
nor U5326 (N_5326,N_3681,N_3802);
and U5327 (N_5327,N_4185,N_3554);
nand U5328 (N_5328,N_4116,N_3731);
and U5329 (N_5329,N_4260,N_4417);
and U5330 (N_5330,N_4322,N_4472);
and U5331 (N_5331,N_3830,N_3589);
xor U5332 (N_5332,N_3740,N_3595);
xor U5333 (N_5333,N_4149,N_3110);
or U5334 (N_5334,N_3410,N_3917);
and U5335 (N_5335,N_3751,N_3192);
or U5336 (N_5336,N_4423,N_3231);
nand U5337 (N_5337,N_3228,N_3022);
and U5338 (N_5338,N_3138,N_3171);
nand U5339 (N_5339,N_3573,N_3719);
nand U5340 (N_5340,N_4011,N_3820);
nor U5341 (N_5341,N_3852,N_4182);
or U5342 (N_5342,N_3577,N_3962);
nor U5343 (N_5343,N_3686,N_4216);
nand U5344 (N_5344,N_3509,N_3728);
nand U5345 (N_5345,N_4274,N_4150);
nor U5346 (N_5346,N_3322,N_3076);
or U5347 (N_5347,N_4341,N_3850);
nor U5348 (N_5348,N_3306,N_4396);
and U5349 (N_5349,N_3449,N_4499);
nand U5350 (N_5350,N_3320,N_3556);
nand U5351 (N_5351,N_4055,N_4151);
or U5352 (N_5352,N_3428,N_4117);
nand U5353 (N_5353,N_3824,N_3313);
or U5354 (N_5354,N_4185,N_3449);
or U5355 (N_5355,N_3903,N_3173);
or U5356 (N_5356,N_3302,N_3708);
nand U5357 (N_5357,N_3277,N_3216);
or U5358 (N_5358,N_4189,N_4484);
xor U5359 (N_5359,N_4318,N_3614);
or U5360 (N_5360,N_4080,N_4019);
or U5361 (N_5361,N_3413,N_3339);
nor U5362 (N_5362,N_3963,N_3168);
and U5363 (N_5363,N_3373,N_4079);
nor U5364 (N_5364,N_3217,N_3494);
or U5365 (N_5365,N_3887,N_3779);
nor U5366 (N_5366,N_3888,N_3059);
and U5367 (N_5367,N_4239,N_4307);
nor U5368 (N_5368,N_3704,N_3904);
and U5369 (N_5369,N_3286,N_4102);
nor U5370 (N_5370,N_3750,N_4414);
xor U5371 (N_5371,N_3671,N_3590);
nor U5372 (N_5372,N_4341,N_3107);
and U5373 (N_5373,N_4152,N_3003);
or U5374 (N_5374,N_3589,N_3629);
and U5375 (N_5375,N_3894,N_4040);
and U5376 (N_5376,N_3494,N_3604);
nand U5377 (N_5377,N_3284,N_3424);
and U5378 (N_5378,N_3381,N_4073);
nand U5379 (N_5379,N_3047,N_3973);
or U5380 (N_5380,N_3144,N_4285);
and U5381 (N_5381,N_3403,N_4464);
and U5382 (N_5382,N_3886,N_3284);
nor U5383 (N_5383,N_3768,N_3336);
and U5384 (N_5384,N_3307,N_3098);
nand U5385 (N_5385,N_3817,N_3173);
nor U5386 (N_5386,N_3557,N_3847);
nor U5387 (N_5387,N_4260,N_4399);
or U5388 (N_5388,N_3270,N_4385);
or U5389 (N_5389,N_4380,N_3341);
and U5390 (N_5390,N_3216,N_3313);
or U5391 (N_5391,N_3486,N_4264);
xnor U5392 (N_5392,N_3816,N_3504);
nor U5393 (N_5393,N_3837,N_4420);
nand U5394 (N_5394,N_4465,N_3229);
and U5395 (N_5395,N_4423,N_3671);
and U5396 (N_5396,N_3003,N_3569);
nand U5397 (N_5397,N_4196,N_4320);
nor U5398 (N_5398,N_3002,N_4017);
nand U5399 (N_5399,N_4407,N_3622);
xnor U5400 (N_5400,N_4155,N_4481);
nand U5401 (N_5401,N_3457,N_4328);
nand U5402 (N_5402,N_3565,N_3895);
and U5403 (N_5403,N_3912,N_3725);
and U5404 (N_5404,N_3541,N_4277);
or U5405 (N_5405,N_3683,N_4403);
xnor U5406 (N_5406,N_3382,N_3837);
xnor U5407 (N_5407,N_3574,N_3054);
nor U5408 (N_5408,N_3232,N_3437);
or U5409 (N_5409,N_3797,N_3906);
nor U5410 (N_5410,N_3743,N_3449);
nor U5411 (N_5411,N_3627,N_3067);
nand U5412 (N_5412,N_3367,N_4298);
nand U5413 (N_5413,N_3547,N_3197);
nand U5414 (N_5414,N_4198,N_4179);
nand U5415 (N_5415,N_4018,N_3079);
and U5416 (N_5416,N_4101,N_3585);
xnor U5417 (N_5417,N_3703,N_3405);
xnor U5418 (N_5418,N_3307,N_4256);
or U5419 (N_5419,N_4118,N_3522);
and U5420 (N_5420,N_3166,N_3717);
and U5421 (N_5421,N_3414,N_3940);
nand U5422 (N_5422,N_3249,N_4487);
nand U5423 (N_5423,N_4499,N_3546);
xnor U5424 (N_5424,N_3307,N_3325);
or U5425 (N_5425,N_4061,N_3363);
nand U5426 (N_5426,N_3961,N_4026);
nand U5427 (N_5427,N_3168,N_3744);
nand U5428 (N_5428,N_3706,N_4448);
or U5429 (N_5429,N_4402,N_3841);
or U5430 (N_5430,N_3530,N_4338);
or U5431 (N_5431,N_4164,N_4096);
and U5432 (N_5432,N_3274,N_4053);
and U5433 (N_5433,N_3806,N_3298);
nor U5434 (N_5434,N_4175,N_3297);
or U5435 (N_5435,N_3359,N_3234);
or U5436 (N_5436,N_4408,N_4246);
and U5437 (N_5437,N_3345,N_3797);
and U5438 (N_5438,N_3174,N_3791);
nand U5439 (N_5439,N_3345,N_3304);
nor U5440 (N_5440,N_4262,N_4456);
nor U5441 (N_5441,N_3841,N_3282);
nand U5442 (N_5442,N_3019,N_3471);
or U5443 (N_5443,N_4219,N_3653);
nand U5444 (N_5444,N_4123,N_3318);
nand U5445 (N_5445,N_4182,N_3477);
and U5446 (N_5446,N_3873,N_3188);
xnor U5447 (N_5447,N_4361,N_3562);
and U5448 (N_5448,N_3818,N_3713);
or U5449 (N_5449,N_3293,N_3558);
nor U5450 (N_5450,N_3900,N_3481);
xor U5451 (N_5451,N_3290,N_4402);
nor U5452 (N_5452,N_3265,N_3656);
and U5453 (N_5453,N_3835,N_4239);
nor U5454 (N_5454,N_3670,N_3317);
or U5455 (N_5455,N_3172,N_3480);
nor U5456 (N_5456,N_3921,N_3073);
nor U5457 (N_5457,N_4284,N_3987);
nor U5458 (N_5458,N_4461,N_3491);
nor U5459 (N_5459,N_4126,N_4375);
and U5460 (N_5460,N_3013,N_4454);
xnor U5461 (N_5461,N_4416,N_4151);
and U5462 (N_5462,N_4309,N_3820);
or U5463 (N_5463,N_4183,N_4196);
and U5464 (N_5464,N_4425,N_4472);
and U5465 (N_5465,N_3218,N_3461);
nor U5466 (N_5466,N_3758,N_3715);
nand U5467 (N_5467,N_3845,N_3689);
nor U5468 (N_5468,N_3856,N_3927);
or U5469 (N_5469,N_3267,N_4225);
and U5470 (N_5470,N_4150,N_3326);
nor U5471 (N_5471,N_4361,N_3905);
nor U5472 (N_5472,N_3394,N_3178);
nand U5473 (N_5473,N_3410,N_3043);
nor U5474 (N_5474,N_4120,N_3417);
nand U5475 (N_5475,N_4485,N_4353);
and U5476 (N_5476,N_3798,N_3793);
nor U5477 (N_5477,N_3493,N_3036);
and U5478 (N_5478,N_3449,N_4405);
or U5479 (N_5479,N_4005,N_3348);
or U5480 (N_5480,N_3222,N_3200);
nand U5481 (N_5481,N_4376,N_3680);
and U5482 (N_5482,N_3703,N_3377);
nand U5483 (N_5483,N_3865,N_3802);
and U5484 (N_5484,N_3321,N_4356);
or U5485 (N_5485,N_4459,N_3304);
xnor U5486 (N_5486,N_3402,N_3732);
or U5487 (N_5487,N_3448,N_3546);
and U5488 (N_5488,N_4302,N_4278);
or U5489 (N_5489,N_3136,N_4040);
nand U5490 (N_5490,N_4162,N_3780);
nor U5491 (N_5491,N_4353,N_3376);
or U5492 (N_5492,N_3288,N_3945);
nor U5493 (N_5493,N_4487,N_3779);
and U5494 (N_5494,N_3295,N_4265);
or U5495 (N_5495,N_3795,N_3768);
or U5496 (N_5496,N_3197,N_3615);
or U5497 (N_5497,N_3707,N_4106);
xor U5498 (N_5498,N_3261,N_3717);
and U5499 (N_5499,N_3229,N_3908);
nand U5500 (N_5500,N_3730,N_4042);
xnor U5501 (N_5501,N_3618,N_4044);
nor U5502 (N_5502,N_3116,N_3471);
nand U5503 (N_5503,N_3555,N_4322);
and U5504 (N_5504,N_3521,N_3245);
nor U5505 (N_5505,N_3670,N_4150);
xnor U5506 (N_5506,N_3279,N_4195);
and U5507 (N_5507,N_3141,N_3406);
nor U5508 (N_5508,N_3987,N_3109);
or U5509 (N_5509,N_3901,N_3688);
nor U5510 (N_5510,N_3184,N_4158);
nand U5511 (N_5511,N_3556,N_3379);
and U5512 (N_5512,N_4467,N_4463);
xnor U5513 (N_5513,N_3200,N_3831);
and U5514 (N_5514,N_3611,N_3651);
or U5515 (N_5515,N_4187,N_4176);
nand U5516 (N_5516,N_4150,N_3629);
nand U5517 (N_5517,N_3031,N_4143);
nor U5518 (N_5518,N_3181,N_3414);
or U5519 (N_5519,N_3268,N_3040);
or U5520 (N_5520,N_4485,N_3796);
and U5521 (N_5521,N_3292,N_3565);
nand U5522 (N_5522,N_3189,N_3375);
nor U5523 (N_5523,N_3679,N_3080);
nor U5524 (N_5524,N_4213,N_4190);
nand U5525 (N_5525,N_3608,N_3492);
and U5526 (N_5526,N_3853,N_4435);
and U5527 (N_5527,N_4124,N_4263);
or U5528 (N_5528,N_3897,N_4413);
and U5529 (N_5529,N_3222,N_3449);
and U5530 (N_5530,N_3635,N_3219);
or U5531 (N_5531,N_4178,N_4391);
nor U5532 (N_5532,N_3687,N_3727);
nand U5533 (N_5533,N_3967,N_3208);
nor U5534 (N_5534,N_3476,N_3466);
and U5535 (N_5535,N_4459,N_4101);
or U5536 (N_5536,N_3938,N_4090);
xnor U5537 (N_5537,N_3552,N_3031);
and U5538 (N_5538,N_3641,N_4135);
and U5539 (N_5539,N_3875,N_4025);
nand U5540 (N_5540,N_3984,N_3313);
nand U5541 (N_5541,N_3407,N_3163);
nor U5542 (N_5542,N_4106,N_4331);
nand U5543 (N_5543,N_3797,N_4086);
or U5544 (N_5544,N_4423,N_3844);
nor U5545 (N_5545,N_3122,N_3940);
nor U5546 (N_5546,N_3717,N_3590);
xnor U5547 (N_5547,N_3286,N_4159);
nand U5548 (N_5548,N_3909,N_3137);
or U5549 (N_5549,N_3941,N_4052);
nand U5550 (N_5550,N_3725,N_3717);
nor U5551 (N_5551,N_3994,N_3181);
nand U5552 (N_5552,N_4404,N_3115);
or U5553 (N_5553,N_4152,N_3092);
and U5554 (N_5554,N_4337,N_3696);
nand U5555 (N_5555,N_3250,N_3217);
nor U5556 (N_5556,N_4263,N_3243);
nor U5557 (N_5557,N_3060,N_3471);
xor U5558 (N_5558,N_3221,N_4444);
or U5559 (N_5559,N_3145,N_3593);
nor U5560 (N_5560,N_3727,N_3435);
nand U5561 (N_5561,N_3325,N_4257);
and U5562 (N_5562,N_4268,N_4060);
and U5563 (N_5563,N_3363,N_3336);
or U5564 (N_5564,N_3646,N_3979);
and U5565 (N_5565,N_3941,N_3343);
nand U5566 (N_5566,N_4284,N_3520);
and U5567 (N_5567,N_3207,N_3782);
or U5568 (N_5568,N_4078,N_3288);
nand U5569 (N_5569,N_3911,N_4277);
nand U5570 (N_5570,N_3613,N_4045);
or U5571 (N_5571,N_4218,N_3509);
nor U5572 (N_5572,N_3218,N_3308);
and U5573 (N_5573,N_3361,N_4194);
xor U5574 (N_5574,N_4023,N_3874);
nand U5575 (N_5575,N_3611,N_3657);
and U5576 (N_5576,N_3431,N_4088);
or U5577 (N_5577,N_3467,N_3910);
and U5578 (N_5578,N_3338,N_3545);
and U5579 (N_5579,N_4485,N_4482);
or U5580 (N_5580,N_3019,N_3140);
nand U5581 (N_5581,N_4114,N_3052);
or U5582 (N_5582,N_3542,N_3677);
nand U5583 (N_5583,N_3874,N_3254);
and U5584 (N_5584,N_3694,N_3525);
and U5585 (N_5585,N_3623,N_3355);
and U5586 (N_5586,N_3126,N_3986);
nand U5587 (N_5587,N_3891,N_3464);
or U5588 (N_5588,N_3040,N_3926);
or U5589 (N_5589,N_3707,N_4479);
xnor U5590 (N_5590,N_3886,N_3193);
and U5591 (N_5591,N_3828,N_3469);
and U5592 (N_5592,N_3114,N_3263);
xnor U5593 (N_5593,N_3289,N_4339);
or U5594 (N_5594,N_4292,N_3235);
or U5595 (N_5595,N_3836,N_3941);
xor U5596 (N_5596,N_3989,N_3359);
and U5597 (N_5597,N_4087,N_4261);
or U5598 (N_5598,N_3204,N_3142);
nand U5599 (N_5599,N_3150,N_3299);
nor U5600 (N_5600,N_3086,N_3652);
nor U5601 (N_5601,N_3450,N_4499);
xnor U5602 (N_5602,N_4262,N_3526);
or U5603 (N_5603,N_3921,N_4219);
nor U5604 (N_5604,N_4269,N_3834);
nor U5605 (N_5605,N_3260,N_3445);
nand U5606 (N_5606,N_4189,N_3348);
xor U5607 (N_5607,N_4476,N_4412);
or U5608 (N_5608,N_4416,N_4158);
or U5609 (N_5609,N_3283,N_3028);
or U5610 (N_5610,N_3608,N_3315);
nand U5611 (N_5611,N_4095,N_3539);
xor U5612 (N_5612,N_3988,N_3128);
nand U5613 (N_5613,N_4354,N_3347);
nor U5614 (N_5614,N_4122,N_3038);
xnor U5615 (N_5615,N_4205,N_3099);
nand U5616 (N_5616,N_3617,N_3230);
or U5617 (N_5617,N_3609,N_4375);
or U5618 (N_5618,N_4392,N_3612);
xor U5619 (N_5619,N_3703,N_3596);
and U5620 (N_5620,N_3748,N_3490);
nor U5621 (N_5621,N_3866,N_4220);
and U5622 (N_5622,N_3832,N_3314);
nor U5623 (N_5623,N_4177,N_3838);
nand U5624 (N_5624,N_3266,N_3548);
nand U5625 (N_5625,N_3475,N_4419);
or U5626 (N_5626,N_3361,N_3200);
xor U5627 (N_5627,N_3473,N_3871);
xnor U5628 (N_5628,N_4133,N_3821);
nor U5629 (N_5629,N_4452,N_3890);
or U5630 (N_5630,N_3748,N_3426);
or U5631 (N_5631,N_3311,N_3379);
nand U5632 (N_5632,N_3714,N_3009);
and U5633 (N_5633,N_4308,N_3760);
nand U5634 (N_5634,N_3490,N_3897);
and U5635 (N_5635,N_3852,N_4241);
nand U5636 (N_5636,N_4149,N_3746);
nand U5637 (N_5637,N_4100,N_3609);
nor U5638 (N_5638,N_3352,N_3149);
nand U5639 (N_5639,N_3029,N_4106);
and U5640 (N_5640,N_4495,N_3956);
and U5641 (N_5641,N_3088,N_3215);
nand U5642 (N_5642,N_4003,N_4420);
nand U5643 (N_5643,N_3074,N_4328);
nand U5644 (N_5644,N_3505,N_3713);
nor U5645 (N_5645,N_4241,N_3603);
xor U5646 (N_5646,N_4180,N_3835);
or U5647 (N_5647,N_3977,N_4385);
or U5648 (N_5648,N_4050,N_4026);
and U5649 (N_5649,N_4226,N_3969);
nor U5650 (N_5650,N_3563,N_3379);
nor U5651 (N_5651,N_4351,N_4065);
and U5652 (N_5652,N_3850,N_3411);
or U5653 (N_5653,N_3166,N_4025);
nor U5654 (N_5654,N_3305,N_3770);
nand U5655 (N_5655,N_3692,N_4377);
xnor U5656 (N_5656,N_3382,N_3290);
nand U5657 (N_5657,N_3336,N_4234);
nor U5658 (N_5658,N_3619,N_3073);
nand U5659 (N_5659,N_3070,N_4248);
or U5660 (N_5660,N_3671,N_3795);
nor U5661 (N_5661,N_4020,N_4407);
nor U5662 (N_5662,N_3936,N_3383);
nand U5663 (N_5663,N_4401,N_3510);
nor U5664 (N_5664,N_4062,N_3382);
nor U5665 (N_5665,N_4253,N_3747);
xnor U5666 (N_5666,N_3758,N_4100);
and U5667 (N_5667,N_3887,N_4216);
nor U5668 (N_5668,N_3499,N_3157);
or U5669 (N_5669,N_4391,N_3018);
and U5670 (N_5670,N_4454,N_3628);
nand U5671 (N_5671,N_4251,N_4288);
or U5672 (N_5672,N_3817,N_4342);
or U5673 (N_5673,N_3360,N_3078);
and U5674 (N_5674,N_4014,N_4482);
or U5675 (N_5675,N_4466,N_3274);
xnor U5676 (N_5676,N_4236,N_4362);
or U5677 (N_5677,N_3735,N_4409);
and U5678 (N_5678,N_3687,N_3311);
or U5679 (N_5679,N_3037,N_4031);
nand U5680 (N_5680,N_3450,N_3900);
nor U5681 (N_5681,N_3386,N_4478);
nand U5682 (N_5682,N_4329,N_4188);
nor U5683 (N_5683,N_3239,N_4172);
xnor U5684 (N_5684,N_3465,N_4133);
and U5685 (N_5685,N_4102,N_3842);
nor U5686 (N_5686,N_3903,N_4222);
or U5687 (N_5687,N_3126,N_3172);
nand U5688 (N_5688,N_3715,N_3371);
xnor U5689 (N_5689,N_4154,N_3812);
or U5690 (N_5690,N_3010,N_3053);
and U5691 (N_5691,N_4314,N_4383);
nand U5692 (N_5692,N_4419,N_3632);
nand U5693 (N_5693,N_3389,N_3283);
or U5694 (N_5694,N_3867,N_4055);
nand U5695 (N_5695,N_3896,N_3743);
or U5696 (N_5696,N_4145,N_3499);
and U5697 (N_5697,N_4483,N_4167);
nand U5698 (N_5698,N_3345,N_3694);
or U5699 (N_5699,N_3527,N_3752);
and U5700 (N_5700,N_3053,N_3931);
nand U5701 (N_5701,N_4081,N_3751);
nor U5702 (N_5702,N_3769,N_3577);
or U5703 (N_5703,N_4022,N_3350);
or U5704 (N_5704,N_3047,N_3201);
nor U5705 (N_5705,N_3592,N_3849);
and U5706 (N_5706,N_4363,N_4144);
and U5707 (N_5707,N_4319,N_3917);
xnor U5708 (N_5708,N_3821,N_4239);
and U5709 (N_5709,N_3192,N_3983);
nand U5710 (N_5710,N_3573,N_4094);
and U5711 (N_5711,N_3627,N_4235);
nor U5712 (N_5712,N_3627,N_4204);
nand U5713 (N_5713,N_3331,N_3005);
nor U5714 (N_5714,N_4163,N_4025);
nor U5715 (N_5715,N_3592,N_3132);
nor U5716 (N_5716,N_3974,N_3328);
nor U5717 (N_5717,N_3138,N_4234);
or U5718 (N_5718,N_3368,N_3798);
or U5719 (N_5719,N_3557,N_3185);
or U5720 (N_5720,N_3347,N_4236);
nor U5721 (N_5721,N_4371,N_3931);
nor U5722 (N_5722,N_3111,N_3517);
xor U5723 (N_5723,N_4374,N_3452);
nand U5724 (N_5724,N_3878,N_4106);
nor U5725 (N_5725,N_4120,N_3476);
and U5726 (N_5726,N_4068,N_3876);
or U5727 (N_5727,N_4205,N_3570);
or U5728 (N_5728,N_3815,N_3772);
and U5729 (N_5729,N_4460,N_3150);
nor U5730 (N_5730,N_3015,N_3745);
nor U5731 (N_5731,N_3616,N_3527);
and U5732 (N_5732,N_3547,N_4134);
nor U5733 (N_5733,N_3620,N_4485);
nand U5734 (N_5734,N_3437,N_3939);
xor U5735 (N_5735,N_4464,N_3080);
or U5736 (N_5736,N_3152,N_4218);
and U5737 (N_5737,N_3766,N_3595);
nor U5738 (N_5738,N_3152,N_4439);
nor U5739 (N_5739,N_3094,N_3951);
and U5740 (N_5740,N_4436,N_4064);
xor U5741 (N_5741,N_4201,N_4425);
nand U5742 (N_5742,N_4429,N_3298);
nor U5743 (N_5743,N_3066,N_3660);
or U5744 (N_5744,N_3197,N_3458);
or U5745 (N_5745,N_3527,N_3735);
xor U5746 (N_5746,N_3087,N_3324);
or U5747 (N_5747,N_4190,N_3090);
nor U5748 (N_5748,N_4337,N_3563);
nor U5749 (N_5749,N_4134,N_3848);
and U5750 (N_5750,N_3518,N_3727);
or U5751 (N_5751,N_3960,N_3314);
nand U5752 (N_5752,N_4307,N_3175);
nor U5753 (N_5753,N_4084,N_3159);
and U5754 (N_5754,N_3103,N_4039);
and U5755 (N_5755,N_3681,N_4339);
nand U5756 (N_5756,N_4242,N_4229);
and U5757 (N_5757,N_4362,N_3372);
nor U5758 (N_5758,N_4286,N_3758);
xnor U5759 (N_5759,N_3358,N_3885);
and U5760 (N_5760,N_3358,N_3629);
nor U5761 (N_5761,N_3156,N_4094);
or U5762 (N_5762,N_3553,N_3947);
and U5763 (N_5763,N_3656,N_4162);
and U5764 (N_5764,N_3173,N_4499);
and U5765 (N_5765,N_3898,N_3278);
and U5766 (N_5766,N_3842,N_3141);
or U5767 (N_5767,N_4287,N_3569);
xnor U5768 (N_5768,N_4259,N_3244);
and U5769 (N_5769,N_3480,N_3383);
xor U5770 (N_5770,N_3351,N_3771);
xnor U5771 (N_5771,N_3926,N_3888);
nor U5772 (N_5772,N_3663,N_4163);
xor U5773 (N_5773,N_3483,N_4038);
nand U5774 (N_5774,N_3333,N_3903);
nor U5775 (N_5775,N_3012,N_3960);
and U5776 (N_5776,N_3747,N_3142);
nor U5777 (N_5777,N_3811,N_3901);
nor U5778 (N_5778,N_3567,N_3079);
nand U5779 (N_5779,N_3298,N_4400);
nor U5780 (N_5780,N_4046,N_3233);
and U5781 (N_5781,N_4119,N_4092);
nor U5782 (N_5782,N_4402,N_3580);
and U5783 (N_5783,N_3636,N_3037);
or U5784 (N_5784,N_4005,N_3322);
nor U5785 (N_5785,N_4439,N_3413);
nor U5786 (N_5786,N_3355,N_3820);
nor U5787 (N_5787,N_3314,N_4405);
xor U5788 (N_5788,N_4024,N_3293);
nor U5789 (N_5789,N_4223,N_3281);
and U5790 (N_5790,N_3277,N_4417);
nor U5791 (N_5791,N_3562,N_3479);
and U5792 (N_5792,N_3159,N_3832);
nand U5793 (N_5793,N_3411,N_4062);
nor U5794 (N_5794,N_3142,N_4263);
nor U5795 (N_5795,N_3168,N_3745);
or U5796 (N_5796,N_4437,N_4266);
nor U5797 (N_5797,N_3748,N_4259);
or U5798 (N_5798,N_3845,N_3104);
nor U5799 (N_5799,N_4338,N_3323);
or U5800 (N_5800,N_3090,N_3791);
or U5801 (N_5801,N_3796,N_4274);
and U5802 (N_5802,N_4030,N_3204);
or U5803 (N_5803,N_3994,N_3454);
and U5804 (N_5804,N_3910,N_3054);
nor U5805 (N_5805,N_4230,N_4334);
and U5806 (N_5806,N_4191,N_4456);
nand U5807 (N_5807,N_3811,N_3181);
and U5808 (N_5808,N_3414,N_3111);
or U5809 (N_5809,N_3092,N_3390);
and U5810 (N_5810,N_4214,N_4305);
and U5811 (N_5811,N_4137,N_3060);
nand U5812 (N_5812,N_4216,N_4288);
or U5813 (N_5813,N_3072,N_3337);
nor U5814 (N_5814,N_4368,N_3045);
or U5815 (N_5815,N_3651,N_3103);
xnor U5816 (N_5816,N_4133,N_3341);
or U5817 (N_5817,N_3698,N_3449);
or U5818 (N_5818,N_3072,N_3708);
and U5819 (N_5819,N_4145,N_4364);
or U5820 (N_5820,N_3375,N_3314);
and U5821 (N_5821,N_3554,N_3370);
xnor U5822 (N_5822,N_3118,N_3961);
nand U5823 (N_5823,N_3143,N_3257);
nor U5824 (N_5824,N_3069,N_3844);
nor U5825 (N_5825,N_3389,N_4268);
nor U5826 (N_5826,N_3052,N_3688);
and U5827 (N_5827,N_4361,N_3211);
or U5828 (N_5828,N_3803,N_4145);
or U5829 (N_5829,N_3154,N_3816);
nand U5830 (N_5830,N_3114,N_3661);
or U5831 (N_5831,N_4167,N_3843);
nor U5832 (N_5832,N_3640,N_3975);
nand U5833 (N_5833,N_4115,N_3532);
or U5834 (N_5834,N_3080,N_3178);
and U5835 (N_5835,N_3501,N_4158);
xnor U5836 (N_5836,N_3296,N_4489);
xnor U5837 (N_5837,N_3589,N_4144);
nand U5838 (N_5838,N_3619,N_4156);
nand U5839 (N_5839,N_4040,N_3768);
xor U5840 (N_5840,N_4005,N_3323);
and U5841 (N_5841,N_3537,N_4331);
nand U5842 (N_5842,N_4017,N_3223);
or U5843 (N_5843,N_3437,N_3054);
nand U5844 (N_5844,N_3037,N_3159);
or U5845 (N_5845,N_4251,N_3874);
nor U5846 (N_5846,N_4436,N_4359);
or U5847 (N_5847,N_3998,N_3513);
or U5848 (N_5848,N_3072,N_3358);
nand U5849 (N_5849,N_3060,N_4158);
and U5850 (N_5850,N_3947,N_4320);
or U5851 (N_5851,N_4405,N_3903);
and U5852 (N_5852,N_3510,N_4050);
nor U5853 (N_5853,N_4173,N_3260);
or U5854 (N_5854,N_4236,N_3292);
xnor U5855 (N_5855,N_3056,N_3447);
nand U5856 (N_5856,N_3611,N_4449);
or U5857 (N_5857,N_3822,N_3387);
nor U5858 (N_5858,N_3359,N_4040);
or U5859 (N_5859,N_4050,N_4410);
or U5860 (N_5860,N_4171,N_4023);
and U5861 (N_5861,N_3135,N_3861);
and U5862 (N_5862,N_3247,N_3330);
nor U5863 (N_5863,N_3393,N_4254);
nand U5864 (N_5864,N_3654,N_3846);
and U5865 (N_5865,N_3041,N_3638);
nand U5866 (N_5866,N_4198,N_3427);
nand U5867 (N_5867,N_3953,N_4027);
nor U5868 (N_5868,N_3073,N_3855);
nor U5869 (N_5869,N_3083,N_3603);
nor U5870 (N_5870,N_3626,N_4126);
nor U5871 (N_5871,N_4440,N_3227);
nor U5872 (N_5872,N_4393,N_4453);
or U5873 (N_5873,N_4097,N_4343);
nor U5874 (N_5874,N_4489,N_3070);
or U5875 (N_5875,N_3926,N_3214);
nand U5876 (N_5876,N_3958,N_3465);
xnor U5877 (N_5877,N_4027,N_4052);
nand U5878 (N_5878,N_3846,N_3938);
nand U5879 (N_5879,N_3252,N_3535);
nand U5880 (N_5880,N_3734,N_3202);
or U5881 (N_5881,N_3606,N_4389);
nor U5882 (N_5882,N_4062,N_3306);
nor U5883 (N_5883,N_3451,N_3368);
nor U5884 (N_5884,N_3748,N_3297);
or U5885 (N_5885,N_3192,N_4037);
and U5886 (N_5886,N_3733,N_4289);
nand U5887 (N_5887,N_3492,N_4030);
nor U5888 (N_5888,N_3548,N_3681);
or U5889 (N_5889,N_3852,N_3705);
xor U5890 (N_5890,N_3031,N_3737);
and U5891 (N_5891,N_3760,N_3603);
nand U5892 (N_5892,N_3039,N_3715);
and U5893 (N_5893,N_3259,N_4018);
nand U5894 (N_5894,N_3925,N_3018);
nand U5895 (N_5895,N_4369,N_3805);
nand U5896 (N_5896,N_4220,N_4065);
nor U5897 (N_5897,N_4029,N_3504);
nor U5898 (N_5898,N_3180,N_3292);
nor U5899 (N_5899,N_4172,N_3212);
nand U5900 (N_5900,N_3467,N_3776);
nand U5901 (N_5901,N_3541,N_3115);
nand U5902 (N_5902,N_3274,N_3846);
xnor U5903 (N_5903,N_4478,N_3035);
or U5904 (N_5904,N_4024,N_3706);
nand U5905 (N_5905,N_4109,N_3540);
or U5906 (N_5906,N_3220,N_3796);
xor U5907 (N_5907,N_4340,N_3044);
and U5908 (N_5908,N_4084,N_4452);
nor U5909 (N_5909,N_3385,N_4348);
nor U5910 (N_5910,N_3706,N_3330);
xnor U5911 (N_5911,N_4395,N_3904);
xor U5912 (N_5912,N_3544,N_3007);
or U5913 (N_5913,N_3717,N_3136);
nor U5914 (N_5914,N_3322,N_3812);
nand U5915 (N_5915,N_3076,N_4004);
or U5916 (N_5916,N_3342,N_4450);
nand U5917 (N_5917,N_4410,N_3312);
nand U5918 (N_5918,N_3381,N_4048);
xnor U5919 (N_5919,N_3225,N_3213);
and U5920 (N_5920,N_3590,N_4155);
or U5921 (N_5921,N_3932,N_3069);
nor U5922 (N_5922,N_3954,N_3963);
and U5923 (N_5923,N_3764,N_3196);
nor U5924 (N_5924,N_3505,N_4447);
and U5925 (N_5925,N_4351,N_4160);
and U5926 (N_5926,N_4482,N_3309);
and U5927 (N_5927,N_3151,N_3721);
nor U5928 (N_5928,N_3318,N_4091);
xnor U5929 (N_5929,N_3999,N_4110);
and U5930 (N_5930,N_3495,N_3921);
nand U5931 (N_5931,N_3966,N_4043);
and U5932 (N_5932,N_3300,N_3153);
and U5933 (N_5933,N_3404,N_3724);
or U5934 (N_5934,N_4181,N_4353);
nor U5935 (N_5935,N_3860,N_3794);
nand U5936 (N_5936,N_3539,N_3370);
nand U5937 (N_5937,N_3313,N_4143);
and U5938 (N_5938,N_4429,N_3116);
nor U5939 (N_5939,N_3007,N_3270);
nor U5940 (N_5940,N_3695,N_3428);
nor U5941 (N_5941,N_3049,N_4385);
or U5942 (N_5942,N_3046,N_3641);
nor U5943 (N_5943,N_3121,N_3231);
nand U5944 (N_5944,N_3976,N_3187);
nand U5945 (N_5945,N_3523,N_3265);
and U5946 (N_5946,N_3677,N_3074);
and U5947 (N_5947,N_4197,N_3542);
xnor U5948 (N_5948,N_3703,N_4198);
nand U5949 (N_5949,N_3934,N_4072);
or U5950 (N_5950,N_4329,N_4125);
nor U5951 (N_5951,N_3255,N_4093);
nor U5952 (N_5952,N_3874,N_4416);
and U5953 (N_5953,N_3568,N_4419);
and U5954 (N_5954,N_3409,N_3207);
or U5955 (N_5955,N_3534,N_3782);
or U5956 (N_5956,N_4008,N_3680);
nand U5957 (N_5957,N_3012,N_3239);
and U5958 (N_5958,N_3969,N_3162);
nor U5959 (N_5959,N_3509,N_3703);
nor U5960 (N_5960,N_3449,N_4307);
or U5961 (N_5961,N_3331,N_3502);
nor U5962 (N_5962,N_3503,N_3006);
nand U5963 (N_5963,N_3657,N_3155);
nor U5964 (N_5964,N_3316,N_3087);
nand U5965 (N_5965,N_3902,N_3040);
or U5966 (N_5966,N_4020,N_3694);
or U5967 (N_5967,N_3697,N_3297);
nand U5968 (N_5968,N_3891,N_3592);
and U5969 (N_5969,N_3706,N_3732);
or U5970 (N_5970,N_3706,N_3681);
nand U5971 (N_5971,N_3223,N_3029);
nor U5972 (N_5972,N_3237,N_3882);
nand U5973 (N_5973,N_3327,N_3563);
and U5974 (N_5974,N_3713,N_3899);
nor U5975 (N_5975,N_3506,N_4215);
nand U5976 (N_5976,N_3258,N_3311);
xnor U5977 (N_5977,N_3898,N_3488);
or U5978 (N_5978,N_3149,N_3670);
nand U5979 (N_5979,N_3926,N_4186);
xor U5980 (N_5980,N_4471,N_3189);
nor U5981 (N_5981,N_3844,N_4119);
and U5982 (N_5982,N_3352,N_4453);
and U5983 (N_5983,N_4309,N_4306);
or U5984 (N_5984,N_4275,N_4111);
nor U5985 (N_5985,N_3463,N_3791);
or U5986 (N_5986,N_3897,N_3078);
and U5987 (N_5987,N_4089,N_3424);
nor U5988 (N_5988,N_4138,N_3626);
nor U5989 (N_5989,N_3478,N_4481);
nor U5990 (N_5990,N_4130,N_3545);
xor U5991 (N_5991,N_3388,N_3886);
xor U5992 (N_5992,N_3145,N_4097);
nand U5993 (N_5993,N_3287,N_3585);
and U5994 (N_5994,N_3732,N_3576);
or U5995 (N_5995,N_3399,N_3091);
nor U5996 (N_5996,N_3561,N_4151);
and U5997 (N_5997,N_4324,N_4336);
nor U5998 (N_5998,N_4009,N_3415);
and U5999 (N_5999,N_3106,N_3397);
nor U6000 (N_6000,N_5446,N_5417);
or U6001 (N_6001,N_5030,N_4686);
nor U6002 (N_6002,N_5097,N_4973);
or U6003 (N_6003,N_5774,N_5922);
or U6004 (N_6004,N_5309,N_5914);
or U6005 (N_6005,N_5144,N_5258);
or U6006 (N_6006,N_4911,N_5749);
or U6007 (N_6007,N_5761,N_4868);
or U6008 (N_6008,N_5004,N_5586);
or U6009 (N_6009,N_5845,N_4965);
nor U6010 (N_6010,N_5305,N_4711);
or U6011 (N_6011,N_5946,N_5911);
nand U6012 (N_6012,N_4914,N_5278);
nand U6013 (N_6013,N_5671,N_5201);
nand U6014 (N_6014,N_5154,N_4756);
or U6015 (N_6015,N_4987,N_5053);
and U6016 (N_6016,N_5530,N_5992);
nor U6017 (N_6017,N_5033,N_5527);
xnor U6018 (N_6018,N_5467,N_5908);
and U6019 (N_6019,N_5390,N_4865);
nand U6020 (N_6020,N_5287,N_4579);
and U6021 (N_6021,N_5851,N_4584);
nand U6022 (N_6022,N_5898,N_5477);
nand U6023 (N_6023,N_4628,N_5624);
nand U6024 (N_6024,N_5596,N_5580);
nor U6025 (N_6025,N_5393,N_5869);
and U6026 (N_6026,N_5866,N_5308);
nor U6027 (N_6027,N_4891,N_4881);
or U6028 (N_6028,N_5065,N_5516);
or U6029 (N_6029,N_5823,N_5272);
nor U6030 (N_6030,N_4734,N_5350);
nand U6031 (N_6031,N_5369,N_4998);
and U6032 (N_6032,N_4918,N_5450);
nand U6033 (N_6033,N_4852,N_5737);
nand U6034 (N_6034,N_5262,N_5300);
nor U6035 (N_6035,N_5036,N_4720);
and U6036 (N_6036,N_5786,N_5564);
nand U6037 (N_6037,N_4989,N_4775);
nor U6038 (N_6038,N_5407,N_5005);
and U6039 (N_6039,N_5844,N_4971);
nand U6040 (N_6040,N_4674,N_5008);
xnor U6041 (N_6041,N_4599,N_5022);
or U6042 (N_6042,N_5076,N_5971);
and U6043 (N_6043,N_5158,N_4814);
nor U6044 (N_6044,N_5981,N_4548);
and U6045 (N_6045,N_4899,N_4532);
xor U6046 (N_6046,N_5521,N_4933);
or U6047 (N_6047,N_5820,N_5080);
nand U6048 (N_6048,N_5687,N_4692);
nand U6049 (N_6049,N_5345,N_5323);
and U6050 (N_6050,N_4701,N_5479);
or U6051 (N_6051,N_4633,N_4691);
nand U6052 (N_6052,N_5481,N_5608);
and U6053 (N_6053,N_5909,N_4901);
or U6054 (N_6054,N_4926,N_5821);
nor U6055 (N_6055,N_5319,N_5332);
xnor U6056 (N_6056,N_5705,N_4882);
xor U6057 (N_6057,N_5602,N_4920);
or U6058 (N_6058,N_5797,N_5701);
nand U6059 (N_6059,N_4854,N_5386);
nor U6060 (N_6060,N_5641,N_4554);
or U6061 (N_6061,N_5406,N_5493);
or U6062 (N_6062,N_5796,N_5807);
or U6063 (N_6063,N_4706,N_4813);
nor U6064 (N_6064,N_4904,N_5341);
and U6065 (N_6065,N_4763,N_5415);
nor U6066 (N_6066,N_4846,N_5181);
or U6067 (N_6067,N_5333,N_5413);
or U6068 (N_6068,N_4552,N_4961);
or U6069 (N_6069,N_5441,N_4540);
or U6070 (N_6070,N_4947,N_5924);
nand U6071 (N_6071,N_5685,N_5187);
nand U6072 (N_6072,N_5092,N_5681);
nand U6073 (N_6073,N_4767,N_5140);
nor U6074 (N_6074,N_5003,N_5155);
and U6075 (N_6075,N_4507,N_5280);
nor U6076 (N_6076,N_4531,N_4976);
nand U6077 (N_6077,N_5791,N_5253);
nor U6078 (N_6078,N_5546,N_4956);
and U6079 (N_6079,N_5178,N_5955);
nor U6080 (N_6080,N_4707,N_4716);
or U6081 (N_6081,N_4663,N_4627);
nand U6082 (N_6082,N_5795,N_5666);
and U6083 (N_6083,N_5805,N_5794);
and U6084 (N_6084,N_5301,N_5950);
nor U6085 (N_6085,N_5182,N_5104);
or U6086 (N_6086,N_5164,N_5355);
and U6087 (N_6087,N_5398,N_4796);
nor U6088 (N_6088,N_5524,N_5549);
or U6089 (N_6089,N_4872,N_4553);
nand U6090 (N_6090,N_5224,N_5903);
nand U6091 (N_6091,N_4644,N_5730);
xor U6092 (N_6092,N_5125,N_4656);
nor U6093 (N_6093,N_5512,N_4819);
nand U6094 (N_6094,N_5382,N_5622);
xor U6095 (N_6095,N_4608,N_4909);
and U6096 (N_6096,N_5281,N_4870);
xor U6097 (N_6097,N_4858,N_5090);
nor U6098 (N_6098,N_5001,N_5311);
nand U6099 (N_6099,N_4793,N_4855);
nand U6100 (N_6100,N_5352,N_5475);
nand U6101 (N_6101,N_4517,N_4768);
and U6102 (N_6102,N_4725,N_5228);
or U6103 (N_6103,N_5019,N_4839);
xor U6104 (N_6104,N_4984,N_5139);
nand U6105 (N_6105,N_5704,N_5128);
xnor U6106 (N_6106,N_5800,N_5348);
and U6107 (N_6107,N_5274,N_4685);
or U6108 (N_6108,N_5112,N_4774);
or U6109 (N_6109,N_5552,N_5566);
and U6110 (N_6110,N_5168,N_4829);
and U6111 (N_6111,N_4563,N_4510);
or U6112 (N_6112,N_4835,N_5130);
nor U6113 (N_6113,N_4542,N_5260);
nor U6114 (N_6114,N_5317,N_5222);
nand U6115 (N_6115,N_5978,N_5115);
xor U6116 (N_6116,N_5255,N_5659);
or U6117 (N_6117,N_4797,N_4986);
or U6118 (N_6118,N_4703,N_4903);
or U6119 (N_6119,N_5011,N_4597);
nand U6120 (N_6120,N_4958,N_5663);
nand U6121 (N_6121,N_5472,N_5344);
and U6122 (N_6122,N_5453,N_5949);
nor U6123 (N_6123,N_5536,N_5361);
and U6124 (N_6124,N_4577,N_5848);
or U6125 (N_6125,N_5623,N_4980);
nor U6126 (N_6126,N_4805,N_5331);
or U6127 (N_6127,N_5969,N_5604);
xnor U6128 (N_6128,N_4724,N_5018);
nor U6129 (N_6129,N_5902,N_4623);
or U6130 (N_6130,N_4880,N_5172);
nand U6131 (N_6131,N_4755,N_4772);
nand U6132 (N_6132,N_4594,N_5451);
xor U6133 (N_6133,N_5715,N_5392);
nand U6134 (N_6134,N_4782,N_5804);
and U6135 (N_6135,N_5123,N_4739);
and U6136 (N_6136,N_5121,N_5034);
and U6137 (N_6137,N_5551,N_4516);
nand U6138 (N_6138,N_4970,N_5970);
and U6139 (N_6139,N_5405,N_4940);
and U6140 (N_6140,N_5427,N_4524);
nor U6141 (N_6141,N_5174,N_4567);
nor U6142 (N_6142,N_4837,N_5058);
or U6143 (N_6143,N_5209,N_4543);
or U6144 (N_6144,N_5347,N_4727);
nand U6145 (N_6145,N_4888,N_5738);
or U6146 (N_6146,N_5818,N_5487);
and U6147 (N_6147,N_5132,N_5974);
nor U6148 (N_6148,N_5322,N_5967);
and U6149 (N_6149,N_4983,N_5858);
and U6150 (N_6150,N_5070,N_5489);
nor U6151 (N_6151,N_5229,N_5577);
and U6152 (N_6152,N_5147,N_5100);
nor U6153 (N_6153,N_5072,N_5270);
nand U6154 (N_6154,N_5779,N_4562);
nor U6155 (N_6155,N_4698,N_5134);
or U6156 (N_6156,N_4893,N_5513);
and U6157 (N_6157,N_4718,N_5921);
and U6158 (N_6158,N_5885,N_4972);
nor U6159 (N_6159,N_4683,N_5269);
nor U6160 (N_6160,N_5062,N_5627);
nand U6161 (N_6161,N_4700,N_4745);
nor U6162 (N_6162,N_5015,N_4557);
and U6163 (N_6163,N_5199,N_5785);
nor U6164 (N_6164,N_5867,N_5443);
nand U6165 (N_6165,N_4515,N_4907);
nor U6166 (N_6166,N_5116,N_5445);
nor U6167 (N_6167,N_4662,N_5849);
nor U6168 (N_6168,N_5051,N_4578);
or U6169 (N_6169,N_5086,N_5833);
or U6170 (N_6170,N_5888,N_5197);
or U6171 (N_6171,N_4821,N_4536);
xnor U6172 (N_6172,N_4714,N_4787);
or U6173 (N_6173,N_5702,N_5814);
or U6174 (N_6174,N_4635,N_5648);
nor U6175 (N_6175,N_4581,N_4619);
or U6176 (N_6176,N_5784,N_5929);
nor U6177 (N_6177,N_5223,N_4539);
nor U6178 (N_6178,N_5754,N_4664);
or U6179 (N_6179,N_4693,N_5872);
nor U6180 (N_6180,N_4896,N_5576);
or U6181 (N_6181,N_4670,N_5762);
and U6182 (N_6182,N_4849,N_4929);
nand U6183 (N_6183,N_4944,N_5395);
nand U6184 (N_6184,N_5662,N_4530);
or U6185 (N_6185,N_5620,N_5822);
nor U6186 (N_6186,N_4886,N_5161);
nand U6187 (N_6187,N_4570,N_5057);
nor U6188 (N_6188,N_5462,N_4509);
nor U6189 (N_6189,N_4967,N_4760);
and U6190 (N_6190,N_5440,N_4648);
nand U6191 (N_6191,N_5052,N_5141);
nor U6192 (N_6192,N_5593,N_5235);
nor U6193 (N_6193,N_4687,N_5327);
and U6194 (N_6194,N_5096,N_4874);
and U6195 (N_6195,N_4750,N_5965);
nand U6196 (N_6196,N_4501,N_4733);
nand U6197 (N_6197,N_5679,N_5519);
and U6198 (N_6198,N_5334,N_5084);
and U6199 (N_6199,N_4576,N_5979);
xor U6200 (N_6200,N_5460,N_5799);
nand U6201 (N_6201,N_5013,N_4786);
nor U6202 (N_6202,N_4746,N_5202);
nor U6203 (N_6203,N_5046,N_5753);
xor U6204 (N_6204,N_4593,N_5543);
and U6205 (N_6205,N_4943,N_5189);
nor U6206 (N_6206,N_5429,N_4521);
or U6207 (N_6207,N_5610,N_5863);
and U6208 (N_6208,N_5126,N_5721);
and U6209 (N_6209,N_5066,N_4777);
xnor U6210 (N_6210,N_4559,N_4595);
nand U6211 (N_6211,N_5289,N_5634);
nand U6212 (N_6212,N_5342,N_5220);
nand U6213 (N_6213,N_5233,N_5242);
and U6214 (N_6214,N_5094,N_5490);
nand U6215 (N_6215,N_5887,N_4761);
xor U6216 (N_6216,N_5259,N_4988);
nor U6217 (N_6217,N_5673,N_5617);
and U6218 (N_6218,N_5569,N_4827);
xnor U6219 (N_6219,N_5548,N_5353);
nor U6220 (N_6220,N_4678,N_5442);
nand U6221 (N_6221,N_5991,N_4556);
and U6222 (N_6222,N_5195,N_4938);
xnor U6223 (N_6223,N_5600,N_5205);
and U6224 (N_6224,N_5607,N_5166);
or U6225 (N_6225,N_4946,N_5938);
or U6226 (N_6226,N_4978,N_5896);
nand U6227 (N_6227,N_5919,N_4551);
xor U6228 (N_6228,N_5956,N_5783);
nor U6229 (N_6229,N_4916,N_5964);
nand U6230 (N_6230,N_5570,N_4728);
or U6231 (N_6231,N_5063,N_5905);
nand U6232 (N_6232,N_4751,N_5295);
xor U6233 (N_6233,N_5547,N_4915);
or U6234 (N_6234,N_5159,N_5684);
and U6235 (N_6235,N_4520,N_4999);
and U6236 (N_6236,N_5539,N_5145);
and U6237 (N_6237,N_5711,N_4809);
nor U6238 (N_6238,N_5320,N_4618);
and U6239 (N_6239,N_5410,N_5175);
nand U6240 (N_6240,N_5455,N_5689);
or U6241 (N_6241,N_5787,N_5364);
or U6242 (N_6242,N_5952,N_5012);
nand U6243 (N_6243,N_5709,N_5581);
xnor U6244 (N_6244,N_5691,N_5230);
and U6245 (N_6245,N_5582,N_5328);
nand U6246 (N_6246,N_5138,N_5387);
and U6247 (N_6247,N_4705,N_5501);
nor U6248 (N_6248,N_5492,N_4866);
nand U6249 (N_6249,N_4784,N_5384);
and U6250 (N_6250,N_4921,N_5719);
nand U6251 (N_6251,N_5628,N_5817);
and U6252 (N_6252,N_4922,N_4522);
or U6253 (N_6253,N_5024,N_5575);
or U6254 (N_6254,N_5926,N_5894);
nor U6255 (N_6255,N_5373,N_5183);
nand U6256 (N_6256,N_5559,N_5767);
nand U6257 (N_6257,N_5706,N_5854);
and U6258 (N_6258,N_5114,N_5944);
or U6259 (N_6259,N_5284,N_4824);
nand U6260 (N_6260,N_5133,N_5734);
or U6261 (N_6261,N_5621,N_5841);
nor U6262 (N_6262,N_5766,N_5626);
nand U6263 (N_6263,N_4964,N_5553);
nand U6264 (N_6264,N_5304,N_4651);
xnor U6265 (N_6265,N_5237,N_4936);
or U6266 (N_6266,N_4877,N_5870);
or U6267 (N_6267,N_5777,N_5054);
and U6268 (N_6268,N_5389,N_5639);
and U6269 (N_6269,N_5152,N_4995);
and U6270 (N_6270,N_5035,N_5079);
nand U6271 (N_6271,N_4785,N_4833);
nand U6272 (N_6272,N_5862,N_5474);
and U6273 (N_6273,N_5840,N_5055);
or U6274 (N_6274,N_5560,N_5645);
or U6275 (N_6275,N_5716,N_4639);
xor U6276 (N_6276,N_4723,N_5680);
or U6277 (N_6277,N_4658,N_5307);
or U6278 (N_6278,N_4607,N_5647);
and U6279 (N_6279,N_5297,N_5438);
nor U6280 (N_6280,N_5509,N_5023);
nand U6281 (N_6281,N_5942,N_5400);
or U6282 (N_6282,N_5574,N_5021);
nor U6283 (N_6283,N_4857,N_5589);
nor U6284 (N_6284,N_5940,N_5105);
or U6285 (N_6285,N_5402,N_4752);
or U6286 (N_6286,N_4677,N_4979);
and U6287 (N_6287,N_5976,N_5945);
nand U6288 (N_6288,N_5338,N_5835);
nand U6289 (N_6289,N_5522,N_5157);
or U6290 (N_6290,N_5765,N_5414);
and U6291 (N_6291,N_4759,N_4744);
or U6292 (N_6292,N_5782,N_5918);
and U6293 (N_6293,N_4631,N_4884);
xnor U6294 (N_6294,N_5408,N_5637);
nand U6295 (N_6295,N_5044,N_5473);
nor U6296 (N_6296,N_5668,N_5325);
nor U6297 (N_6297,N_4708,N_4569);
or U6298 (N_6298,N_5708,N_5912);
xor U6299 (N_6299,N_4828,N_4661);
or U6300 (N_6300,N_5456,N_5351);
nand U6301 (N_6301,N_4695,N_5310);
nor U6302 (N_6302,N_4737,N_5354);
or U6303 (N_6303,N_5561,N_5798);
xor U6304 (N_6304,N_4900,N_4905);
nor U6305 (N_6305,N_5091,N_4616);
nand U6306 (N_6306,N_4721,N_5215);
or U6307 (N_6307,N_4790,N_5266);
nand U6308 (N_6308,N_5583,N_4541);
nand U6309 (N_6309,N_5421,N_5367);
and U6310 (N_6310,N_5712,N_4859);
nand U6311 (N_6311,N_5953,N_4729);
nor U6312 (N_6312,N_5409,N_5993);
or U6313 (N_6313,N_4764,N_4694);
xor U6314 (N_6314,N_5847,N_5459);
xnor U6315 (N_6315,N_5486,N_5207);
xnor U6316 (N_6316,N_5119,N_4808);
nand U6317 (N_6317,N_5632,N_5435);
nand U6318 (N_6318,N_5741,N_4630);
and U6319 (N_6319,N_4843,N_5240);
or U6320 (N_6320,N_5430,N_5770);
nand U6321 (N_6321,N_4932,N_5177);
nor U6322 (N_6322,N_4713,N_5986);
and U6323 (N_6323,N_5692,N_5554);
nor U6324 (N_6324,N_5261,N_5020);
and U6325 (N_6325,N_5951,N_4625);
and U6326 (N_6326,N_5625,N_4959);
and U6327 (N_6327,N_4602,N_5745);
and U6328 (N_6328,N_5082,N_5667);
or U6329 (N_6329,N_4601,N_5191);
and U6330 (N_6330,N_5838,N_4996);
nor U6331 (N_6331,N_5349,N_4546);
nand U6332 (N_6332,N_5039,N_4732);
nor U6333 (N_6333,N_5049,N_4848);
or U6334 (N_6334,N_5683,N_5180);
xnor U6335 (N_6335,N_5935,N_5934);
or U6336 (N_6336,N_5127,N_5603);
nand U6337 (N_6337,N_4957,N_5428);
nor U6338 (N_6338,N_5907,N_5694);
and U6339 (N_6339,N_5495,N_4939);
nor U6340 (N_6340,N_4962,N_5366);
or U6341 (N_6341,N_5433,N_5592);
and U6342 (N_6342,N_5041,N_4640);
nand U6343 (N_6343,N_5775,N_5426);
nor U6344 (N_6344,N_5267,N_5131);
nor U6345 (N_6345,N_5980,N_4969);
nand U6346 (N_6346,N_4681,N_5025);
or U6347 (N_6347,N_4645,N_5078);
xnor U6348 (N_6348,N_4679,N_5109);
xor U6349 (N_6349,N_5383,N_5920);
nand U6350 (N_6350,N_5422,N_5707);
and U6351 (N_6351,N_5803,N_5163);
nor U6352 (N_6352,N_5448,N_5615);
nand U6353 (N_6353,N_5482,N_5497);
or U6354 (N_6354,N_4585,N_4842);
and U6355 (N_6355,N_5009,N_5954);
nor U6356 (N_6356,N_4758,N_5286);
nand U6357 (N_6357,N_4804,N_5491);
or U6358 (N_6358,N_5572,N_4527);
nand U6359 (N_6359,N_4950,N_5606);
or U6360 (N_6360,N_5032,N_5293);
xor U6361 (N_6361,N_5478,N_5578);
and U6362 (N_6362,N_5296,N_5654);
nand U6363 (N_6363,N_5876,N_4596);
and U6364 (N_6364,N_4652,N_5816);
nor U6365 (N_6365,N_5111,N_5312);
and U6366 (N_6366,N_5404,N_5585);
nor U6367 (N_6367,N_4642,N_4610);
nand U6368 (N_6368,N_5703,N_5877);
nor U6369 (N_6369,N_5802,N_4898);
nand U6370 (N_6370,N_5743,N_4773);
and U6371 (N_6371,N_4948,N_4781);
nor U6372 (N_6372,N_4923,N_4757);
xnor U6373 (N_6373,N_4794,N_4655);
nor U6374 (N_6374,N_5873,N_5045);
and U6375 (N_6375,N_4941,N_4803);
or U6376 (N_6376,N_5511,N_5047);
and U6377 (N_6377,N_5612,N_5732);
or U6378 (N_6378,N_4586,N_4518);
nand U6379 (N_6379,N_5378,N_5579);
or U6380 (N_6380,N_4966,N_4743);
or U6381 (N_6381,N_5672,N_4770);
or U6382 (N_6382,N_5864,N_4826);
xor U6383 (N_6383,N_5488,N_5326);
nand U6384 (N_6384,N_5218,N_5103);
nor U6385 (N_6385,N_5861,N_5239);
and U6386 (N_6386,N_5038,N_5542);
and U6387 (N_6387,N_5584,N_5498);
or U6388 (N_6388,N_4688,N_5941);
or U6389 (N_6389,N_4665,N_4798);
nand U6390 (N_6390,N_5609,N_4788);
nand U6391 (N_6391,N_4816,N_5678);
nor U6392 (N_6392,N_5660,N_5416);
nor U6393 (N_6393,N_4555,N_5273);
nand U6394 (N_6394,N_5891,N_5102);
nand U6395 (N_6395,N_5081,N_4748);
or U6396 (N_6396,N_5343,N_5257);
nand U6397 (N_6397,N_5882,N_5748);
or U6398 (N_6398,N_4573,N_5664);
nand U6399 (N_6399,N_5360,N_4825);
and U6400 (N_6400,N_5238,N_4762);
xnor U6401 (N_6401,N_4889,N_5359);
nor U6402 (N_6402,N_5670,N_5372);
nand U6403 (N_6403,N_4547,N_5120);
and U6404 (N_6404,N_5727,N_5613);
nand U6405 (N_6405,N_5346,N_4935);
and U6406 (N_6406,N_5243,N_5083);
nor U6407 (N_6407,N_4847,N_5595);
nand U6408 (N_6408,N_5532,N_4913);
or U6409 (N_6409,N_5983,N_5494);
nor U6410 (N_6410,N_5910,N_4831);
or U6411 (N_6411,N_5827,N_4609);
or U6412 (N_6412,N_4800,N_5151);
nand U6413 (N_6413,N_4869,N_5614);
nand U6414 (N_6414,N_5886,N_4666);
nor U6415 (N_6415,N_5788,N_5757);
nand U6416 (N_6416,N_5605,N_5675);
or U6417 (N_6417,N_5533,N_4657);
nor U6418 (N_6418,N_5436,N_5562);
nor U6419 (N_6419,N_5982,N_4840);
nand U6420 (N_6420,N_4856,N_5165);
and U6421 (N_6421,N_4985,N_4690);
nand U6422 (N_6422,N_5002,N_5074);
nand U6423 (N_6423,N_5192,N_5856);
and U6424 (N_6424,N_4942,N_5778);
nand U6425 (N_6425,N_5290,N_5150);
xor U6426 (N_6426,N_5837,N_5040);
nor U6427 (N_6427,N_4712,N_5294);
xnor U6428 (N_6428,N_4887,N_5529);
nor U6429 (N_6429,N_5813,N_4885);
xor U6430 (N_6430,N_4953,N_5206);
nand U6431 (N_6431,N_5998,N_5892);
and U6432 (N_6432,N_4931,N_5806);
or U6433 (N_6433,N_5618,N_5832);
and U6434 (N_6434,N_5283,N_5733);
xor U6435 (N_6435,N_5458,N_4955);
or U6436 (N_6436,N_4680,N_4912);
nor U6437 (N_6437,N_5231,N_4626);
nor U6438 (N_6438,N_4765,N_5850);
xor U6439 (N_6439,N_4861,N_4671);
xor U6440 (N_6440,N_5792,N_5819);
nor U6441 (N_6441,N_5194,N_5135);
nand U6442 (N_6442,N_4994,N_5517);
and U6443 (N_6443,N_4675,N_4769);
nand U6444 (N_6444,N_5972,N_5597);
and U6445 (N_6445,N_5504,N_5061);
and U6446 (N_6446,N_4937,N_5629);
xnor U6447 (N_6447,N_5789,N_4583);
nand U6448 (N_6448,N_5153,N_5682);
and U6449 (N_6449,N_5060,N_5056);
nand U6450 (N_6450,N_4673,N_5917);
nor U6451 (N_6451,N_5321,N_5977);
and U6452 (N_6452,N_5391,N_5931);
nand U6453 (N_6453,N_5298,N_4830);
and U6454 (N_6454,N_5381,N_5726);
nand U6455 (N_6455,N_5557,N_4776);
or U6456 (N_6456,N_5966,N_4799);
and U6457 (N_6457,N_4867,N_5809);
or U6458 (N_6458,N_5339,N_4982);
nand U6459 (N_6459,N_4974,N_5540);
or U6460 (N_6460,N_5196,N_5535);
nor U6461 (N_6461,N_5656,N_5865);
or U6462 (N_6462,N_5635,N_5520);
and U6463 (N_6463,N_4545,N_4871);
nand U6464 (N_6464,N_5468,N_5996);
nand U6465 (N_6465,N_5810,N_5943);
nand U6466 (N_6466,N_4611,N_5947);
nand U6467 (N_6467,N_4574,N_5507);
and U6468 (N_6468,N_5496,N_5883);
nand U6469 (N_6469,N_5176,N_5718);
and U6470 (N_6470,N_5484,N_4954);
nand U6471 (N_6471,N_5510,N_4636);
and U6472 (N_6472,N_5676,N_5285);
and U6473 (N_6473,N_5143,N_5000);
nor U6474 (N_6474,N_5210,N_5316);
or U6475 (N_6475,N_4910,N_4560);
xnor U6476 (N_6476,N_5480,N_5059);
or U6477 (N_6477,N_5544,N_5700);
nand U6478 (N_6478,N_5225,N_5633);
and U6479 (N_6479,N_5879,N_4836);
or U6480 (N_6480,N_5118,N_5252);
or U6481 (N_6481,N_4513,N_5302);
nor U6482 (N_6482,N_4612,N_4766);
or U6483 (N_6483,N_5631,N_5449);
nand U6484 (N_6484,N_5471,N_4704);
xnor U6485 (N_6485,N_5219,N_4702);
and U6486 (N_6486,N_5014,N_5279);
and U6487 (N_6487,N_4863,N_4778);
or U6488 (N_6488,N_5122,N_4741);
and U6489 (N_6489,N_5999,N_5423);
or U6490 (N_6490,N_4811,N_4506);
nor U6491 (N_6491,N_5336,N_5432);
nor U6492 (N_6492,N_5254,N_5193);
nor U6493 (N_6493,N_5071,N_4927);
nand U6494 (N_6494,N_5531,N_5973);
and U6495 (N_6495,N_4851,N_4591);
and U6496 (N_6496,N_5649,N_5661);
and U6497 (N_6497,N_5651,N_5825);
xnor U6498 (N_6498,N_4806,N_5688);
xnor U6499 (N_6499,N_4643,N_4802);
and U6500 (N_6500,N_4754,N_5048);
and U6501 (N_6501,N_5397,N_4544);
nand U6502 (N_6502,N_5098,N_5095);
or U6503 (N_6503,N_4845,N_5075);
or U6504 (N_6504,N_5503,N_5031);
nand U6505 (N_6505,N_5419,N_5265);
or U6506 (N_6506,N_4902,N_5650);
and U6507 (N_6507,N_4660,N_5485);
and U6508 (N_6508,N_5411,N_5108);
nand U6509 (N_6509,N_5901,N_4511);
or U6510 (N_6510,N_4620,N_5318);
or U6511 (N_6511,N_4622,N_4654);
and U6512 (N_6512,N_5171,N_5525);
nand U6513 (N_6513,N_4928,N_5958);
and U6514 (N_6514,N_5545,N_5099);
nand U6515 (N_6515,N_5747,N_5142);
nor U6516 (N_6516,N_5968,N_4590);
nor U6517 (N_6517,N_4977,N_5506);
nand U6518 (N_6518,N_5959,N_5288);
xnor U6519 (N_6519,N_5263,N_5502);
nand U6520 (N_6520,N_5363,N_5880);
and U6521 (N_6521,N_5466,N_5731);
nand U6522 (N_6522,N_5412,N_5368);
xnor U6523 (N_6523,N_5216,N_4710);
xor U6524 (N_6524,N_5042,N_4740);
and U6525 (N_6525,N_5994,N_5598);
xnor U6526 (N_6526,N_5167,N_4925);
xnor U6527 (N_6527,N_4722,N_4504);
nor U6528 (N_6528,N_5424,N_5227);
nand U6529 (N_6529,N_4792,N_5275);
or U6530 (N_6530,N_5722,N_4637);
nor U6531 (N_6531,N_5928,N_5010);
nor U6532 (N_6532,N_4862,N_4791);
or U6533 (N_6533,N_5751,N_5315);
or U6534 (N_6534,N_5808,N_4952);
xor U6535 (N_6535,N_5793,N_4917);
nand U6536 (N_6536,N_4629,N_5695);
nor U6537 (N_6537,N_5699,N_5790);
nor U6538 (N_6538,N_5812,N_5772);
nand U6539 (N_6539,N_5107,N_5616);
and U6540 (N_6540,N_5874,N_4589);
or U6541 (N_6541,N_5454,N_5160);
nand U6542 (N_6542,N_5370,N_4505);
or U6543 (N_6543,N_5420,N_4566);
nand U6544 (N_6544,N_5725,N_5246);
and U6545 (N_6545,N_5871,N_5069);
or U6546 (N_6546,N_5728,N_4614);
nor U6547 (N_6547,N_5884,N_4580);
nor U6548 (N_6548,N_5463,N_5906);
nor U6549 (N_6549,N_4876,N_5729);
and U6550 (N_6550,N_5232,N_5567);
nand U6551 (N_6551,N_5852,N_4731);
xor U6552 (N_6552,N_4508,N_5735);
and U6553 (N_6553,N_5717,N_4738);
and U6554 (N_6554,N_5764,N_5961);
or U6555 (N_6555,N_4834,N_4815);
or U6556 (N_6556,N_5388,N_4981);
nand U6557 (N_6557,N_5425,N_4844);
or U6558 (N_6558,N_4537,N_5444);
nand U6559 (N_6559,N_5271,N_5759);
or U6560 (N_6560,N_5169,N_5101);
or U6561 (N_6561,N_5198,N_4853);
nor U6562 (N_6562,N_4818,N_5299);
nand U6563 (N_6563,N_4747,N_5248);
nor U6564 (N_6564,N_5829,N_4565);
and U6565 (N_6565,N_5526,N_5895);
nor U6566 (N_6566,N_5889,N_4502);
nor U6567 (N_6567,N_5282,N_4615);
or U6568 (N_6568,N_5591,N_5439);
nor U6569 (N_6569,N_4951,N_4906);
or U6570 (N_6570,N_4575,N_5136);
nand U6571 (N_6571,N_4592,N_4650);
nand U6572 (N_6572,N_5916,N_5936);
nor U6573 (N_6573,N_4550,N_5358);
xnor U6574 (N_6574,N_5990,N_5093);
or U6575 (N_6575,N_5842,N_5106);
xor U6576 (N_6576,N_5362,N_5534);
nand U6577 (N_6577,N_5113,N_5619);
or U6578 (N_6578,N_5830,N_5963);
nand U6579 (N_6579,N_5244,N_5203);
or U6580 (N_6580,N_5881,N_5758);
nand U6581 (N_6581,N_5587,N_4822);
nand U6582 (N_6582,N_5962,N_5937);
or U6583 (N_6583,N_5465,N_5050);
nor U6584 (N_6584,N_5655,N_4993);
nand U6585 (N_6585,N_5697,N_4649);
xor U6586 (N_6586,N_5590,N_5418);
nand U6587 (N_6587,N_4699,N_4668);
and U6588 (N_6588,N_5173,N_5669);
or U6589 (N_6589,N_4696,N_5644);
nor U6590 (N_6590,N_5927,N_4512);
or U6591 (N_6591,N_5568,N_5630);
and U6592 (N_6592,N_5188,N_4503);
nor U6593 (N_6593,N_5213,N_5073);
nor U6594 (N_6594,N_4820,N_5904);
nand U6595 (N_6595,N_5646,N_4653);
nor U6596 (N_6596,N_4624,N_5768);
nand U6597 (N_6597,N_5515,N_5357);
nor U6598 (N_6598,N_5989,N_5211);
or U6599 (N_6599,N_4735,N_4715);
nand U6600 (N_6600,N_5826,N_5828);
or U6601 (N_6601,N_5129,N_4789);
and U6602 (N_6602,N_5016,N_5571);
and U6603 (N_6603,N_5162,N_5376);
or U6604 (N_6604,N_5760,N_4968);
and U6605 (N_6605,N_4807,N_5556);
nor U6606 (N_6606,N_4641,N_5356);
and U6607 (N_6607,N_5756,N_5170);
nand U6608 (N_6608,N_4990,N_4736);
nand U6609 (N_6609,N_5893,N_5746);
nand U6610 (N_6610,N_5179,N_4895);
nor U6611 (N_6611,N_5401,N_5464);
nor U6612 (N_6612,N_5736,N_4617);
or U6613 (N_6613,N_5755,N_5781);
nor U6614 (N_6614,N_4634,N_5500);
or U6615 (N_6615,N_4535,N_5988);
nor U6616 (N_6616,N_4838,N_5380);
nand U6617 (N_6617,N_5313,N_4526);
nor U6618 (N_6618,N_5868,N_5930);
nand U6619 (N_6619,N_5537,N_5200);
xor U6620 (N_6620,N_4883,N_5740);
nor U6621 (N_6621,N_4742,N_5599);
and U6622 (N_6622,N_4753,N_5693);
or U6623 (N_6623,N_4682,N_4908);
xor U6624 (N_6624,N_5452,N_4647);
or U6625 (N_6625,N_5037,N_5508);
or U6626 (N_6626,N_4646,N_4783);
and U6627 (N_6627,N_4684,N_5514);
or U6628 (N_6628,N_5523,N_5017);
or U6629 (N_6629,N_5714,N_5447);
nor U6630 (N_6630,N_5379,N_5696);
and U6631 (N_6631,N_4894,N_4672);
or U6632 (N_6632,N_4621,N_5241);
and U6633 (N_6633,N_5403,N_4689);
or U6634 (N_6634,N_5470,N_4749);
nor U6635 (N_6635,N_5247,N_4864);
or U6636 (N_6636,N_5505,N_5214);
or U6637 (N_6637,N_4605,N_5636);
and U6638 (N_6638,N_5149,N_5834);
nor U6639 (N_6639,N_5853,N_5337);
or U6640 (N_6640,N_5611,N_4500);
nand U6641 (N_6641,N_4523,N_4606);
and U6642 (N_6642,N_4558,N_5457);
or U6643 (N_6643,N_5763,N_5026);
and U6644 (N_6644,N_5801,N_5291);
nand U6645 (N_6645,N_4717,N_5713);
or U6646 (N_6646,N_4812,N_5839);
nand U6647 (N_6647,N_4588,N_5190);
nand U6648 (N_6648,N_5306,N_5997);
or U6649 (N_6649,N_5212,N_5750);
and U6650 (N_6650,N_4878,N_5890);
nand U6651 (N_6651,N_4582,N_5900);
nor U6652 (N_6652,N_5185,N_4945);
and U6653 (N_6653,N_5156,N_5780);
and U6654 (N_6654,N_4659,N_5277);
and U6655 (N_6655,N_4841,N_4801);
nor U6656 (N_6656,N_5565,N_4992);
nand U6657 (N_6657,N_5186,N_4533);
nor U6658 (N_6658,N_5377,N_5984);
and U6659 (N_6659,N_4525,N_5857);
xor U6660 (N_6660,N_5365,N_5957);
nor U6661 (N_6661,N_5913,N_5836);
or U6662 (N_6662,N_5690,N_5292);
or U6663 (N_6663,N_5742,N_5723);
or U6664 (N_6664,N_5824,N_5563);
xor U6665 (N_6665,N_4860,N_5434);
or U6666 (N_6666,N_5371,N_4963);
or U6667 (N_6667,N_5875,N_4529);
or U6668 (N_6668,N_5226,N_5249);
and U6669 (N_6669,N_5739,N_5588);
nand U6670 (N_6670,N_4991,N_5330);
nand U6671 (N_6671,N_4697,N_5276);
xor U6672 (N_6672,N_5939,N_5932);
nor U6673 (N_6673,N_4771,N_5686);
nor U6674 (N_6674,N_5665,N_5815);
or U6675 (N_6675,N_5773,N_4850);
nor U6676 (N_6676,N_4676,N_5985);
nand U6677 (N_6677,N_5217,N_5394);
and U6678 (N_6678,N_4528,N_5385);
nand U6679 (N_6679,N_5043,N_5028);
nand U6680 (N_6680,N_5710,N_4780);
xor U6681 (N_6681,N_5085,N_4779);
nand U6682 (N_6682,N_5483,N_5550);
nor U6683 (N_6683,N_4519,N_5831);
or U6684 (N_6684,N_5975,N_5329);
nor U6685 (N_6685,N_5064,N_5399);
and U6686 (N_6686,N_5769,N_4919);
nor U6687 (N_6687,N_4897,N_5221);
and U6688 (N_6688,N_4873,N_5846);
or U6689 (N_6689,N_5236,N_5340);
nand U6690 (N_6690,N_4890,N_4613);
and U6691 (N_6691,N_4638,N_5007);
or U6692 (N_6692,N_5776,N_4534);
nor U6693 (N_6693,N_4817,N_5860);
nand U6694 (N_6694,N_5897,N_4960);
or U6695 (N_6695,N_5724,N_5657);
nand U6696 (N_6696,N_4571,N_5987);
or U6697 (N_6697,N_5068,N_5771);
nor U6698 (N_6698,N_4572,N_5915);
nand U6699 (N_6699,N_5925,N_5461);
nand U6700 (N_6700,N_5184,N_5640);
nand U6701 (N_6701,N_5643,N_5933);
or U6702 (N_6702,N_5245,N_4667);
nor U6703 (N_6703,N_5324,N_4603);
and U6704 (N_6704,N_5878,N_5264);
or U6705 (N_6705,N_5087,N_5006);
nor U6706 (N_6706,N_4875,N_5431);
and U6707 (N_6707,N_4514,N_5960);
and U6708 (N_6708,N_5811,N_5251);
nor U6709 (N_6709,N_5555,N_4997);
nand U6710 (N_6710,N_5476,N_5843);
nand U6711 (N_6711,N_5601,N_5256);
nor U6712 (N_6712,N_4924,N_5995);
nand U6713 (N_6713,N_5652,N_5234);
or U6714 (N_6714,N_4564,N_5744);
or U6715 (N_6715,N_4719,N_4709);
nand U6716 (N_6716,N_5948,N_5117);
and U6717 (N_6717,N_4832,N_5396);
and U6718 (N_6718,N_5499,N_4538);
nand U6719 (N_6719,N_4879,N_4892);
nand U6720 (N_6720,N_4600,N_4604);
nor U6721 (N_6721,N_5752,N_5638);
nand U6722 (N_6722,N_5594,N_5653);
nand U6723 (N_6723,N_4823,N_4726);
xnor U6724 (N_6724,N_5642,N_5067);
and U6725 (N_6725,N_5268,N_4730);
nor U6726 (N_6726,N_5538,N_5541);
nor U6727 (N_6727,N_5528,N_5137);
nand U6728 (N_6728,N_4549,N_5658);
xnor U6729 (N_6729,N_4975,N_4810);
nand U6730 (N_6730,N_5698,N_4598);
and U6731 (N_6731,N_5027,N_5250);
nand U6732 (N_6732,N_4669,N_5077);
xnor U6733 (N_6733,N_5859,N_5375);
xnor U6734 (N_6734,N_5124,N_5089);
nand U6735 (N_6735,N_5303,N_4795);
and U6736 (N_6736,N_4587,N_5146);
nor U6737 (N_6737,N_5314,N_4949);
nand U6738 (N_6738,N_5677,N_5088);
nand U6739 (N_6739,N_5558,N_5437);
nand U6740 (N_6740,N_5573,N_5855);
nand U6741 (N_6741,N_5720,N_5029);
xnor U6742 (N_6742,N_5374,N_5518);
nand U6743 (N_6743,N_5204,N_5335);
and U6744 (N_6744,N_4561,N_5208);
xnor U6745 (N_6745,N_5923,N_5110);
or U6746 (N_6746,N_5899,N_5469);
nor U6747 (N_6747,N_4632,N_4934);
nor U6748 (N_6748,N_4930,N_5148);
or U6749 (N_6749,N_5674,N_4568);
xnor U6750 (N_6750,N_5854,N_4796);
or U6751 (N_6751,N_4777,N_4900);
nor U6752 (N_6752,N_4575,N_4724);
nand U6753 (N_6753,N_5388,N_5644);
nand U6754 (N_6754,N_4517,N_4849);
and U6755 (N_6755,N_4793,N_5824);
and U6756 (N_6756,N_5287,N_5927);
xnor U6757 (N_6757,N_4861,N_4819);
xnor U6758 (N_6758,N_4860,N_5857);
and U6759 (N_6759,N_5259,N_5303);
nand U6760 (N_6760,N_4735,N_4557);
nand U6761 (N_6761,N_4845,N_4913);
nor U6762 (N_6762,N_5693,N_5186);
or U6763 (N_6763,N_5005,N_4519);
xnor U6764 (N_6764,N_4957,N_5986);
nor U6765 (N_6765,N_5844,N_4776);
nor U6766 (N_6766,N_5354,N_4870);
and U6767 (N_6767,N_4986,N_5478);
and U6768 (N_6768,N_4556,N_5974);
or U6769 (N_6769,N_5794,N_5502);
or U6770 (N_6770,N_4587,N_5301);
xnor U6771 (N_6771,N_5419,N_5341);
nand U6772 (N_6772,N_5229,N_5524);
nor U6773 (N_6773,N_4749,N_5666);
nand U6774 (N_6774,N_5027,N_5062);
xor U6775 (N_6775,N_5123,N_4757);
or U6776 (N_6776,N_4947,N_5834);
and U6777 (N_6777,N_5394,N_4574);
nor U6778 (N_6778,N_4639,N_5159);
nor U6779 (N_6779,N_4693,N_5660);
nand U6780 (N_6780,N_4897,N_5293);
or U6781 (N_6781,N_5771,N_5006);
nor U6782 (N_6782,N_4782,N_5445);
and U6783 (N_6783,N_5421,N_4725);
nand U6784 (N_6784,N_5887,N_5879);
nand U6785 (N_6785,N_5151,N_5790);
or U6786 (N_6786,N_5892,N_5312);
and U6787 (N_6787,N_5618,N_5979);
or U6788 (N_6788,N_4600,N_5123);
or U6789 (N_6789,N_4635,N_4989);
or U6790 (N_6790,N_4973,N_5861);
nand U6791 (N_6791,N_5810,N_5743);
nand U6792 (N_6792,N_5632,N_5043);
nor U6793 (N_6793,N_5780,N_4808);
and U6794 (N_6794,N_4587,N_4663);
nand U6795 (N_6795,N_5197,N_5137);
or U6796 (N_6796,N_4819,N_5630);
nor U6797 (N_6797,N_4887,N_5672);
or U6798 (N_6798,N_5670,N_5153);
nand U6799 (N_6799,N_5187,N_4706);
nand U6800 (N_6800,N_5202,N_5316);
and U6801 (N_6801,N_5552,N_5498);
nand U6802 (N_6802,N_5607,N_5592);
and U6803 (N_6803,N_5120,N_5563);
nor U6804 (N_6804,N_5775,N_4747);
nor U6805 (N_6805,N_5595,N_5770);
or U6806 (N_6806,N_5210,N_5150);
or U6807 (N_6807,N_5406,N_5602);
nand U6808 (N_6808,N_5197,N_5505);
nor U6809 (N_6809,N_5966,N_4562);
nand U6810 (N_6810,N_4831,N_5226);
nand U6811 (N_6811,N_5311,N_5299);
nor U6812 (N_6812,N_5329,N_5359);
nand U6813 (N_6813,N_5866,N_4507);
nor U6814 (N_6814,N_5718,N_5151);
and U6815 (N_6815,N_5647,N_4999);
nand U6816 (N_6816,N_5305,N_4718);
and U6817 (N_6817,N_5347,N_5074);
nor U6818 (N_6818,N_4928,N_4570);
and U6819 (N_6819,N_5616,N_5625);
xnor U6820 (N_6820,N_5883,N_5189);
nor U6821 (N_6821,N_4949,N_5171);
or U6822 (N_6822,N_5290,N_5902);
nand U6823 (N_6823,N_4969,N_5389);
nand U6824 (N_6824,N_5909,N_4580);
nor U6825 (N_6825,N_5323,N_5929);
or U6826 (N_6826,N_5738,N_5997);
and U6827 (N_6827,N_5361,N_5865);
and U6828 (N_6828,N_4866,N_4911);
nor U6829 (N_6829,N_5683,N_5990);
or U6830 (N_6830,N_4914,N_5662);
nor U6831 (N_6831,N_5889,N_4963);
or U6832 (N_6832,N_5215,N_5682);
and U6833 (N_6833,N_4800,N_5723);
and U6834 (N_6834,N_4542,N_5696);
and U6835 (N_6835,N_5013,N_5658);
nor U6836 (N_6836,N_5716,N_4917);
and U6837 (N_6837,N_4818,N_4560);
or U6838 (N_6838,N_5551,N_4892);
nor U6839 (N_6839,N_5185,N_5165);
or U6840 (N_6840,N_5269,N_4945);
nand U6841 (N_6841,N_5132,N_5257);
nor U6842 (N_6842,N_5724,N_4554);
and U6843 (N_6843,N_4565,N_4500);
xnor U6844 (N_6844,N_5512,N_5608);
nor U6845 (N_6845,N_5348,N_5904);
xnor U6846 (N_6846,N_5076,N_4637);
or U6847 (N_6847,N_5558,N_4823);
or U6848 (N_6848,N_5239,N_5918);
nand U6849 (N_6849,N_5416,N_5436);
xor U6850 (N_6850,N_4783,N_4777);
xnor U6851 (N_6851,N_4656,N_4821);
nand U6852 (N_6852,N_5507,N_5669);
nor U6853 (N_6853,N_5119,N_4873);
and U6854 (N_6854,N_5802,N_5258);
or U6855 (N_6855,N_4572,N_4944);
nand U6856 (N_6856,N_5758,N_5347);
and U6857 (N_6857,N_5767,N_5215);
nand U6858 (N_6858,N_5837,N_4577);
or U6859 (N_6859,N_5126,N_5325);
or U6860 (N_6860,N_5336,N_4870);
nand U6861 (N_6861,N_5132,N_5175);
nor U6862 (N_6862,N_4759,N_5749);
and U6863 (N_6863,N_5586,N_5426);
nor U6864 (N_6864,N_4705,N_5543);
and U6865 (N_6865,N_5404,N_4809);
xnor U6866 (N_6866,N_5731,N_4513);
nand U6867 (N_6867,N_4715,N_5667);
nor U6868 (N_6868,N_4552,N_4874);
nor U6869 (N_6869,N_5477,N_5698);
xnor U6870 (N_6870,N_5172,N_4574);
nand U6871 (N_6871,N_4808,N_5121);
and U6872 (N_6872,N_4752,N_5197);
or U6873 (N_6873,N_4830,N_4671);
nand U6874 (N_6874,N_5277,N_4512);
and U6875 (N_6875,N_5720,N_5314);
or U6876 (N_6876,N_5516,N_4937);
nor U6877 (N_6877,N_5727,N_5851);
and U6878 (N_6878,N_5048,N_5447);
and U6879 (N_6879,N_5826,N_5996);
and U6880 (N_6880,N_4543,N_4644);
nand U6881 (N_6881,N_5642,N_4634);
or U6882 (N_6882,N_5695,N_5761);
nand U6883 (N_6883,N_4700,N_5702);
or U6884 (N_6884,N_5511,N_5967);
nand U6885 (N_6885,N_4839,N_4809);
nand U6886 (N_6886,N_4671,N_5018);
nor U6887 (N_6887,N_4524,N_4948);
and U6888 (N_6888,N_4549,N_4865);
or U6889 (N_6889,N_4899,N_5118);
and U6890 (N_6890,N_4676,N_5456);
nor U6891 (N_6891,N_4961,N_4925);
or U6892 (N_6892,N_5676,N_4757);
and U6893 (N_6893,N_5337,N_4723);
or U6894 (N_6894,N_5062,N_5513);
nor U6895 (N_6895,N_4503,N_4944);
nand U6896 (N_6896,N_5779,N_4806);
nor U6897 (N_6897,N_5364,N_5014);
and U6898 (N_6898,N_5435,N_5047);
nand U6899 (N_6899,N_5925,N_4690);
nand U6900 (N_6900,N_5727,N_5329);
nor U6901 (N_6901,N_5649,N_5914);
nor U6902 (N_6902,N_4506,N_5428);
and U6903 (N_6903,N_5046,N_5539);
nor U6904 (N_6904,N_5132,N_5383);
nand U6905 (N_6905,N_5965,N_4567);
nand U6906 (N_6906,N_4819,N_5766);
and U6907 (N_6907,N_5517,N_4925);
nor U6908 (N_6908,N_5641,N_4501);
or U6909 (N_6909,N_5820,N_5503);
or U6910 (N_6910,N_5799,N_5382);
nand U6911 (N_6911,N_5516,N_5244);
or U6912 (N_6912,N_5315,N_5784);
or U6913 (N_6913,N_4857,N_5628);
and U6914 (N_6914,N_5854,N_5379);
nand U6915 (N_6915,N_4724,N_5091);
nand U6916 (N_6916,N_5019,N_5480);
or U6917 (N_6917,N_5610,N_5731);
and U6918 (N_6918,N_4550,N_4519);
or U6919 (N_6919,N_5123,N_5355);
nor U6920 (N_6920,N_5517,N_4622);
and U6921 (N_6921,N_4986,N_5738);
nor U6922 (N_6922,N_5238,N_5183);
or U6923 (N_6923,N_4640,N_4646);
nor U6924 (N_6924,N_4555,N_5803);
or U6925 (N_6925,N_4844,N_5656);
and U6926 (N_6926,N_5438,N_5761);
or U6927 (N_6927,N_4841,N_4799);
and U6928 (N_6928,N_4922,N_5568);
nor U6929 (N_6929,N_5806,N_5058);
and U6930 (N_6930,N_4545,N_5957);
nand U6931 (N_6931,N_5662,N_5260);
nor U6932 (N_6932,N_5637,N_5986);
nor U6933 (N_6933,N_5493,N_5731);
or U6934 (N_6934,N_5684,N_5374);
and U6935 (N_6935,N_5535,N_4842);
xor U6936 (N_6936,N_5762,N_5961);
and U6937 (N_6937,N_5221,N_5192);
and U6938 (N_6938,N_5925,N_5685);
and U6939 (N_6939,N_5483,N_5568);
or U6940 (N_6940,N_4617,N_4809);
nor U6941 (N_6941,N_5497,N_5961);
xor U6942 (N_6942,N_5866,N_4698);
or U6943 (N_6943,N_4806,N_5363);
or U6944 (N_6944,N_4737,N_4927);
nor U6945 (N_6945,N_4899,N_5777);
xor U6946 (N_6946,N_5859,N_5870);
nor U6947 (N_6947,N_5094,N_5281);
nand U6948 (N_6948,N_5121,N_5885);
or U6949 (N_6949,N_5347,N_4828);
or U6950 (N_6950,N_5880,N_4776);
or U6951 (N_6951,N_5800,N_4529);
nor U6952 (N_6952,N_4647,N_4936);
or U6953 (N_6953,N_5968,N_5680);
nor U6954 (N_6954,N_5553,N_4646);
or U6955 (N_6955,N_5295,N_4755);
xnor U6956 (N_6956,N_5927,N_5510);
or U6957 (N_6957,N_4602,N_5639);
nor U6958 (N_6958,N_4786,N_5458);
nor U6959 (N_6959,N_4903,N_5578);
nand U6960 (N_6960,N_4953,N_5005);
xor U6961 (N_6961,N_4917,N_5723);
and U6962 (N_6962,N_5274,N_5094);
or U6963 (N_6963,N_5272,N_5190);
xor U6964 (N_6964,N_4569,N_5646);
and U6965 (N_6965,N_4618,N_5179);
xnor U6966 (N_6966,N_5779,N_5038);
xnor U6967 (N_6967,N_4585,N_4689);
and U6968 (N_6968,N_5440,N_5034);
nor U6969 (N_6969,N_5438,N_5270);
or U6970 (N_6970,N_4910,N_4741);
or U6971 (N_6971,N_4574,N_4860);
and U6972 (N_6972,N_5529,N_5256);
xnor U6973 (N_6973,N_5398,N_4949);
nand U6974 (N_6974,N_5474,N_4749);
nand U6975 (N_6975,N_5402,N_4735);
nand U6976 (N_6976,N_4857,N_5255);
nor U6977 (N_6977,N_5066,N_5211);
nor U6978 (N_6978,N_5540,N_5469);
or U6979 (N_6979,N_4531,N_5269);
or U6980 (N_6980,N_5088,N_5054);
xnor U6981 (N_6981,N_5863,N_5703);
or U6982 (N_6982,N_5535,N_5695);
nor U6983 (N_6983,N_5982,N_5314);
and U6984 (N_6984,N_5324,N_4524);
and U6985 (N_6985,N_5503,N_4771);
and U6986 (N_6986,N_5793,N_4778);
nor U6987 (N_6987,N_4531,N_5653);
or U6988 (N_6988,N_4749,N_5908);
nor U6989 (N_6989,N_5878,N_4605);
xor U6990 (N_6990,N_4999,N_5838);
nand U6991 (N_6991,N_5102,N_5268);
nor U6992 (N_6992,N_5515,N_5022);
nand U6993 (N_6993,N_5008,N_4953);
nor U6994 (N_6994,N_4539,N_5850);
xnor U6995 (N_6995,N_4893,N_5654);
nor U6996 (N_6996,N_5552,N_4853);
nand U6997 (N_6997,N_5954,N_5261);
xor U6998 (N_6998,N_4649,N_4539);
and U6999 (N_6999,N_5421,N_5648);
or U7000 (N_7000,N_4804,N_5645);
xnor U7001 (N_7001,N_5546,N_4921);
and U7002 (N_7002,N_5656,N_4916);
nor U7003 (N_7003,N_5397,N_4773);
or U7004 (N_7004,N_5688,N_5095);
nor U7005 (N_7005,N_4923,N_5152);
nor U7006 (N_7006,N_5902,N_5471);
or U7007 (N_7007,N_5556,N_5895);
xor U7008 (N_7008,N_5544,N_4722);
nor U7009 (N_7009,N_5236,N_4752);
or U7010 (N_7010,N_4825,N_5519);
and U7011 (N_7011,N_4838,N_4773);
nand U7012 (N_7012,N_4806,N_5035);
nor U7013 (N_7013,N_4641,N_5470);
or U7014 (N_7014,N_4821,N_5860);
or U7015 (N_7015,N_5519,N_5970);
nor U7016 (N_7016,N_4835,N_5824);
and U7017 (N_7017,N_5850,N_5353);
and U7018 (N_7018,N_5146,N_4563);
or U7019 (N_7019,N_5293,N_4958);
nor U7020 (N_7020,N_5323,N_5482);
and U7021 (N_7021,N_5465,N_4697);
nor U7022 (N_7022,N_5143,N_4601);
nand U7023 (N_7023,N_5373,N_5311);
nand U7024 (N_7024,N_5735,N_4747);
and U7025 (N_7025,N_4714,N_4864);
nand U7026 (N_7026,N_4653,N_5480);
or U7027 (N_7027,N_5899,N_5486);
or U7028 (N_7028,N_4782,N_5194);
nor U7029 (N_7029,N_5273,N_4878);
and U7030 (N_7030,N_5261,N_5622);
xnor U7031 (N_7031,N_4873,N_5955);
and U7032 (N_7032,N_4843,N_5040);
nor U7033 (N_7033,N_4916,N_4573);
nor U7034 (N_7034,N_5736,N_4552);
or U7035 (N_7035,N_4799,N_4937);
nand U7036 (N_7036,N_5265,N_5889);
nor U7037 (N_7037,N_5951,N_4970);
and U7038 (N_7038,N_5868,N_4752);
or U7039 (N_7039,N_5304,N_5932);
nor U7040 (N_7040,N_5770,N_4528);
nor U7041 (N_7041,N_5187,N_4636);
nor U7042 (N_7042,N_5441,N_4909);
nand U7043 (N_7043,N_5208,N_4952);
nand U7044 (N_7044,N_5289,N_5668);
or U7045 (N_7045,N_5614,N_5883);
nand U7046 (N_7046,N_5695,N_5393);
xor U7047 (N_7047,N_4839,N_5248);
and U7048 (N_7048,N_5749,N_5768);
nor U7049 (N_7049,N_5769,N_4615);
and U7050 (N_7050,N_4916,N_4508);
nor U7051 (N_7051,N_5825,N_4578);
nor U7052 (N_7052,N_5532,N_5928);
nor U7053 (N_7053,N_5183,N_5018);
nand U7054 (N_7054,N_5905,N_5537);
and U7055 (N_7055,N_4671,N_5109);
nor U7056 (N_7056,N_5936,N_5077);
xor U7057 (N_7057,N_5760,N_5250);
nor U7058 (N_7058,N_5610,N_5383);
and U7059 (N_7059,N_4977,N_4812);
nor U7060 (N_7060,N_5576,N_4985);
nand U7061 (N_7061,N_5940,N_5580);
and U7062 (N_7062,N_5409,N_4819);
nor U7063 (N_7063,N_4549,N_5037);
nor U7064 (N_7064,N_4709,N_5596);
nand U7065 (N_7065,N_5177,N_5387);
and U7066 (N_7066,N_5766,N_5872);
and U7067 (N_7067,N_4793,N_5227);
nor U7068 (N_7068,N_4647,N_5139);
and U7069 (N_7069,N_5197,N_4699);
and U7070 (N_7070,N_5849,N_5510);
nor U7071 (N_7071,N_5776,N_5856);
nor U7072 (N_7072,N_4768,N_5191);
and U7073 (N_7073,N_4875,N_5908);
xnor U7074 (N_7074,N_5645,N_4859);
or U7075 (N_7075,N_5606,N_5489);
and U7076 (N_7076,N_5882,N_5179);
nor U7077 (N_7077,N_5355,N_5705);
nand U7078 (N_7078,N_5968,N_4514);
nor U7079 (N_7079,N_4725,N_5055);
nand U7080 (N_7080,N_4934,N_5606);
or U7081 (N_7081,N_4924,N_5139);
and U7082 (N_7082,N_5407,N_5104);
nand U7083 (N_7083,N_5983,N_5528);
nor U7084 (N_7084,N_5815,N_5473);
and U7085 (N_7085,N_4676,N_5580);
and U7086 (N_7086,N_5453,N_5851);
or U7087 (N_7087,N_4971,N_5047);
and U7088 (N_7088,N_4502,N_5688);
nand U7089 (N_7089,N_5683,N_5593);
and U7090 (N_7090,N_4880,N_4960);
or U7091 (N_7091,N_4828,N_5786);
or U7092 (N_7092,N_4845,N_4653);
nor U7093 (N_7093,N_5911,N_5840);
nand U7094 (N_7094,N_4543,N_5598);
and U7095 (N_7095,N_5168,N_4682);
and U7096 (N_7096,N_5532,N_5266);
nand U7097 (N_7097,N_4703,N_4809);
and U7098 (N_7098,N_4692,N_5510);
xor U7099 (N_7099,N_5669,N_5188);
and U7100 (N_7100,N_5832,N_5736);
nor U7101 (N_7101,N_5639,N_5012);
and U7102 (N_7102,N_5503,N_5575);
or U7103 (N_7103,N_5929,N_4958);
nor U7104 (N_7104,N_5616,N_5963);
and U7105 (N_7105,N_5854,N_5378);
nand U7106 (N_7106,N_5908,N_5510);
or U7107 (N_7107,N_4660,N_5844);
xnor U7108 (N_7108,N_5773,N_5953);
and U7109 (N_7109,N_5626,N_5374);
nor U7110 (N_7110,N_5215,N_5297);
or U7111 (N_7111,N_5311,N_5860);
or U7112 (N_7112,N_4614,N_5267);
and U7113 (N_7113,N_5608,N_4600);
and U7114 (N_7114,N_4760,N_4562);
nand U7115 (N_7115,N_4673,N_5186);
nor U7116 (N_7116,N_5510,N_5519);
and U7117 (N_7117,N_5569,N_5102);
or U7118 (N_7118,N_5307,N_4824);
or U7119 (N_7119,N_5625,N_4524);
or U7120 (N_7120,N_4996,N_5546);
nor U7121 (N_7121,N_5281,N_5604);
and U7122 (N_7122,N_5275,N_5025);
nand U7123 (N_7123,N_5870,N_5988);
nand U7124 (N_7124,N_5578,N_5491);
nor U7125 (N_7125,N_5570,N_5092);
nor U7126 (N_7126,N_4899,N_5405);
nor U7127 (N_7127,N_4524,N_5836);
nand U7128 (N_7128,N_4792,N_5564);
nor U7129 (N_7129,N_4675,N_5421);
or U7130 (N_7130,N_4609,N_5094);
nand U7131 (N_7131,N_4555,N_5217);
nand U7132 (N_7132,N_5323,N_5144);
and U7133 (N_7133,N_4610,N_4690);
nand U7134 (N_7134,N_5240,N_5220);
and U7135 (N_7135,N_4732,N_5589);
nor U7136 (N_7136,N_5059,N_4993);
or U7137 (N_7137,N_4737,N_5873);
and U7138 (N_7138,N_5317,N_4970);
nor U7139 (N_7139,N_5495,N_5595);
or U7140 (N_7140,N_5978,N_4613);
or U7141 (N_7141,N_4648,N_5450);
nand U7142 (N_7142,N_5065,N_5994);
nand U7143 (N_7143,N_4979,N_5259);
and U7144 (N_7144,N_4590,N_5079);
and U7145 (N_7145,N_5778,N_4854);
xnor U7146 (N_7146,N_5974,N_5688);
xor U7147 (N_7147,N_5847,N_4855);
nand U7148 (N_7148,N_5997,N_5854);
nand U7149 (N_7149,N_5351,N_4951);
or U7150 (N_7150,N_5731,N_5506);
or U7151 (N_7151,N_5084,N_5188);
nand U7152 (N_7152,N_4743,N_4863);
or U7153 (N_7153,N_5645,N_5113);
nand U7154 (N_7154,N_4544,N_5341);
and U7155 (N_7155,N_4870,N_5372);
nand U7156 (N_7156,N_4537,N_4521);
nand U7157 (N_7157,N_5641,N_5798);
nor U7158 (N_7158,N_4708,N_5048);
nor U7159 (N_7159,N_5122,N_5918);
nor U7160 (N_7160,N_5603,N_5676);
nor U7161 (N_7161,N_5505,N_5739);
and U7162 (N_7162,N_4995,N_5165);
or U7163 (N_7163,N_4701,N_5804);
nand U7164 (N_7164,N_4718,N_5141);
nand U7165 (N_7165,N_4502,N_5476);
nor U7166 (N_7166,N_5651,N_4831);
nor U7167 (N_7167,N_5069,N_4660);
nand U7168 (N_7168,N_5571,N_5742);
nor U7169 (N_7169,N_5296,N_4969);
nor U7170 (N_7170,N_5003,N_4976);
or U7171 (N_7171,N_4985,N_5845);
and U7172 (N_7172,N_5217,N_5695);
nor U7173 (N_7173,N_5897,N_4930);
or U7174 (N_7174,N_5147,N_4738);
nor U7175 (N_7175,N_4515,N_4625);
and U7176 (N_7176,N_5505,N_4754);
nor U7177 (N_7177,N_4934,N_5780);
nand U7178 (N_7178,N_5940,N_5275);
or U7179 (N_7179,N_4991,N_5777);
nor U7180 (N_7180,N_4934,N_4993);
or U7181 (N_7181,N_5026,N_5148);
xor U7182 (N_7182,N_4925,N_5318);
or U7183 (N_7183,N_5047,N_5565);
nor U7184 (N_7184,N_5790,N_5595);
nor U7185 (N_7185,N_5257,N_4760);
xor U7186 (N_7186,N_4889,N_5435);
xnor U7187 (N_7187,N_5849,N_4978);
nand U7188 (N_7188,N_4867,N_5001);
or U7189 (N_7189,N_4646,N_5014);
xor U7190 (N_7190,N_5213,N_5832);
and U7191 (N_7191,N_4812,N_4927);
and U7192 (N_7192,N_5507,N_5994);
or U7193 (N_7193,N_4883,N_5613);
nor U7194 (N_7194,N_4675,N_5063);
nand U7195 (N_7195,N_5165,N_5015);
nor U7196 (N_7196,N_5917,N_4635);
nor U7197 (N_7197,N_4677,N_5012);
nand U7198 (N_7198,N_5473,N_4657);
nand U7199 (N_7199,N_4750,N_5504);
and U7200 (N_7200,N_4955,N_4670);
or U7201 (N_7201,N_5467,N_4914);
nor U7202 (N_7202,N_5611,N_5417);
and U7203 (N_7203,N_4583,N_4841);
nor U7204 (N_7204,N_5259,N_5865);
nor U7205 (N_7205,N_5248,N_4577);
and U7206 (N_7206,N_5349,N_4766);
nand U7207 (N_7207,N_5731,N_4724);
nor U7208 (N_7208,N_5272,N_5560);
or U7209 (N_7209,N_5883,N_5439);
nand U7210 (N_7210,N_4963,N_5291);
or U7211 (N_7211,N_4510,N_5543);
nor U7212 (N_7212,N_4962,N_4532);
and U7213 (N_7213,N_5738,N_5656);
nand U7214 (N_7214,N_5643,N_4550);
and U7215 (N_7215,N_5833,N_4529);
and U7216 (N_7216,N_5787,N_5022);
xnor U7217 (N_7217,N_4818,N_5626);
nand U7218 (N_7218,N_5727,N_4772);
or U7219 (N_7219,N_5154,N_5554);
nand U7220 (N_7220,N_5148,N_5330);
nor U7221 (N_7221,N_5794,N_4868);
nor U7222 (N_7222,N_5567,N_5881);
nor U7223 (N_7223,N_5222,N_5087);
and U7224 (N_7224,N_5806,N_5034);
or U7225 (N_7225,N_5142,N_5357);
and U7226 (N_7226,N_5260,N_4823);
nor U7227 (N_7227,N_5712,N_5143);
or U7228 (N_7228,N_5939,N_4503);
nand U7229 (N_7229,N_5697,N_5134);
or U7230 (N_7230,N_4542,N_4667);
xnor U7231 (N_7231,N_5016,N_5674);
nor U7232 (N_7232,N_4561,N_5633);
nand U7233 (N_7233,N_4705,N_4736);
nor U7234 (N_7234,N_4945,N_5910);
nand U7235 (N_7235,N_4951,N_5070);
nor U7236 (N_7236,N_4865,N_4687);
nor U7237 (N_7237,N_5917,N_5481);
or U7238 (N_7238,N_5453,N_5893);
or U7239 (N_7239,N_4679,N_5514);
and U7240 (N_7240,N_5208,N_5157);
nand U7241 (N_7241,N_5654,N_4903);
xor U7242 (N_7242,N_4974,N_5825);
and U7243 (N_7243,N_5176,N_5635);
and U7244 (N_7244,N_5771,N_5811);
or U7245 (N_7245,N_5826,N_5777);
xnor U7246 (N_7246,N_4558,N_5674);
and U7247 (N_7247,N_4955,N_4880);
or U7248 (N_7248,N_4831,N_5702);
and U7249 (N_7249,N_5448,N_5169);
xor U7250 (N_7250,N_4778,N_5930);
and U7251 (N_7251,N_5321,N_5344);
and U7252 (N_7252,N_5739,N_5718);
or U7253 (N_7253,N_5259,N_5516);
nor U7254 (N_7254,N_5957,N_5540);
and U7255 (N_7255,N_4866,N_5240);
nor U7256 (N_7256,N_4885,N_5215);
or U7257 (N_7257,N_5762,N_5136);
and U7258 (N_7258,N_5766,N_5862);
and U7259 (N_7259,N_5615,N_5869);
nand U7260 (N_7260,N_4949,N_5613);
xor U7261 (N_7261,N_4976,N_5428);
nand U7262 (N_7262,N_4839,N_5033);
nor U7263 (N_7263,N_4942,N_4595);
or U7264 (N_7264,N_5858,N_5717);
or U7265 (N_7265,N_4919,N_5550);
and U7266 (N_7266,N_5014,N_5314);
nor U7267 (N_7267,N_5551,N_5122);
and U7268 (N_7268,N_5832,N_4695);
and U7269 (N_7269,N_4760,N_4617);
nand U7270 (N_7270,N_5091,N_5893);
nor U7271 (N_7271,N_5785,N_5477);
xor U7272 (N_7272,N_4563,N_4837);
and U7273 (N_7273,N_5882,N_5983);
nor U7274 (N_7274,N_4902,N_5876);
or U7275 (N_7275,N_5524,N_5547);
nand U7276 (N_7276,N_4745,N_5487);
and U7277 (N_7277,N_5846,N_4811);
nor U7278 (N_7278,N_5954,N_4623);
or U7279 (N_7279,N_5899,N_5622);
or U7280 (N_7280,N_4749,N_4529);
nor U7281 (N_7281,N_5284,N_4737);
xnor U7282 (N_7282,N_5033,N_4885);
and U7283 (N_7283,N_5781,N_5895);
nand U7284 (N_7284,N_4755,N_4525);
nand U7285 (N_7285,N_4760,N_5246);
or U7286 (N_7286,N_4779,N_5984);
nor U7287 (N_7287,N_5160,N_5710);
nand U7288 (N_7288,N_5589,N_4523);
nor U7289 (N_7289,N_4516,N_5512);
or U7290 (N_7290,N_5665,N_5679);
nand U7291 (N_7291,N_5789,N_4654);
nor U7292 (N_7292,N_5601,N_5575);
nand U7293 (N_7293,N_4553,N_5089);
or U7294 (N_7294,N_5522,N_5626);
nor U7295 (N_7295,N_4561,N_5820);
or U7296 (N_7296,N_5200,N_5210);
or U7297 (N_7297,N_4611,N_4928);
nand U7298 (N_7298,N_5830,N_5435);
or U7299 (N_7299,N_5802,N_5854);
nor U7300 (N_7300,N_4768,N_4963);
xor U7301 (N_7301,N_4799,N_4535);
or U7302 (N_7302,N_5915,N_5776);
xor U7303 (N_7303,N_5695,N_5138);
nand U7304 (N_7304,N_4620,N_4736);
nor U7305 (N_7305,N_5894,N_5668);
or U7306 (N_7306,N_4897,N_5053);
nand U7307 (N_7307,N_5786,N_5030);
and U7308 (N_7308,N_5390,N_5814);
nand U7309 (N_7309,N_5967,N_5787);
or U7310 (N_7310,N_5326,N_5710);
and U7311 (N_7311,N_5191,N_4757);
and U7312 (N_7312,N_5056,N_5403);
and U7313 (N_7313,N_5391,N_4739);
nand U7314 (N_7314,N_5054,N_5515);
nand U7315 (N_7315,N_5754,N_5070);
nand U7316 (N_7316,N_5875,N_5026);
or U7317 (N_7317,N_5059,N_5975);
nand U7318 (N_7318,N_4768,N_4750);
or U7319 (N_7319,N_5067,N_4598);
or U7320 (N_7320,N_5289,N_5344);
nor U7321 (N_7321,N_4945,N_4534);
or U7322 (N_7322,N_5542,N_4573);
and U7323 (N_7323,N_4900,N_5394);
nand U7324 (N_7324,N_5850,N_5580);
nand U7325 (N_7325,N_4677,N_4584);
and U7326 (N_7326,N_4581,N_5957);
nand U7327 (N_7327,N_5948,N_5438);
xnor U7328 (N_7328,N_5082,N_5385);
nand U7329 (N_7329,N_5771,N_5787);
nor U7330 (N_7330,N_5403,N_5745);
or U7331 (N_7331,N_5377,N_5551);
or U7332 (N_7332,N_5066,N_5408);
or U7333 (N_7333,N_5251,N_5700);
nor U7334 (N_7334,N_5663,N_4910);
or U7335 (N_7335,N_5026,N_5430);
and U7336 (N_7336,N_4799,N_5029);
nor U7337 (N_7337,N_5986,N_5210);
nand U7338 (N_7338,N_4796,N_4578);
xnor U7339 (N_7339,N_4660,N_5123);
nand U7340 (N_7340,N_5238,N_5783);
and U7341 (N_7341,N_5355,N_4971);
nand U7342 (N_7342,N_5291,N_5313);
nor U7343 (N_7343,N_5760,N_5793);
or U7344 (N_7344,N_4894,N_5687);
and U7345 (N_7345,N_5938,N_5483);
nand U7346 (N_7346,N_4598,N_4796);
nand U7347 (N_7347,N_5382,N_4791);
nand U7348 (N_7348,N_5278,N_5031);
or U7349 (N_7349,N_5348,N_5119);
nand U7350 (N_7350,N_5967,N_4648);
and U7351 (N_7351,N_4792,N_5429);
nor U7352 (N_7352,N_5951,N_4981);
xor U7353 (N_7353,N_4942,N_4751);
nor U7354 (N_7354,N_4685,N_5967);
or U7355 (N_7355,N_5879,N_5842);
nor U7356 (N_7356,N_5498,N_4822);
or U7357 (N_7357,N_4552,N_5772);
or U7358 (N_7358,N_4697,N_5380);
nor U7359 (N_7359,N_5327,N_5182);
xnor U7360 (N_7360,N_4763,N_5899);
or U7361 (N_7361,N_5680,N_4772);
nor U7362 (N_7362,N_5914,N_5972);
and U7363 (N_7363,N_5073,N_5119);
or U7364 (N_7364,N_5627,N_5973);
xnor U7365 (N_7365,N_5975,N_4893);
or U7366 (N_7366,N_5380,N_5832);
nand U7367 (N_7367,N_4994,N_5423);
nor U7368 (N_7368,N_5812,N_5051);
nor U7369 (N_7369,N_5185,N_5183);
or U7370 (N_7370,N_5904,N_4511);
nand U7371 (N_7371,N_5101,N_5900);
or U7372 (N_7372,N_5560,N_4784);
nor U7373 (N_7373,N_5318,N_5954);
nand U7374 (N_7374,N_4809,N_5962);
nor U7375 (N_7375,N_5923,N_5229);
nand U7376 (N_7376,N_5037,N_5963);
nand U7377 (N_7377,N_4759,N_5209);
nor U7378 (N_7378,N_4982,N_5317);
nor U7379 (N_7379,N_5440,N_5950);
and U7380 (N_7380,N_5074,N_4673);
nand U7381 (N_7381,N_5508,N_4628);
or U7382 (N_7382,N_5999,N_5686);
nand U7383 (N_7383,N_5223,N_5153);
nand U7384 (N_7384,N_4914,N_4531);
nand U7385 (N_7385,N_5756,N_5129);
xnor U7386 (N_7386,N_4776,N_4705);
nor U7387 (N_7387,N_4581,N_5097);
and U7388 (N_7388,N_5219,N_5056);
or U7389 (N_7389,N_5279,N_4561);
or U7390 (N_7390,N_5330,N_4858);
or U7391 (N_7391,N_4511,N_4645);
nor U7392 (N_7392,N_5922,N_4539);
nor U7393 (N_7393,N_5747,N_5341);
and U7394 (N_7394,N_5811,N_4704);
or U7395 (N_7395,N_4980,N_4748);
nand U7396 (N_7396,N_4910,N_5146);
nor U7397 (N_7397,N_4906,N_5682);
or U7398 (N_7398,N_5821,N_5858);
nand U7399 (N_7399,N_5272,N_5794);
nor U7400 (N_7400,N_4888,N_4683);
nand U7401 (N_7401,N_5717,N_4658);
nand U7402 (N_7402,N_5296,N_5179);
nor U7403 (N_7403,N_5222,N_4596);
nor U7404 (N_7404,N_4837,N_5531);
nor U7405 (N_7405,N_5227,N_4889);
or U7406 (N_7406,N_4516,N_5132);
or U7407 (N_7407,N_5876,N_5057);
xor U7408 (N_7408,N_4802,N_4799);
and U7409 (N_7409,N_5406,N_4977);
nand U7410 (N_7410,N_5088,N_5639);
nor U7411 (N_7411,N_5724,N_4562);
nor U7412 (N_7412,N_5401,N_4911);
nand U7413 (N_7413,N_4720,N_5130);
nor U7414 (N_7414,N_5785,N_5554);
nor U7415 (N_7415,N_4900,N_5422);
xor U7416 (N_7416,N_5281,N_4639);
and U7417 (N_7417,N_5359,N_4607);
nand U7418 (N_7418,N_4814,N_5999);
xor U7419 (N_7419,N_4832,N_4982);
nand U7420 (N_7420,N_4729,N_5698);
nor U7421 (N_7421,N_5279,N_5631);
nor U7422 (N_7422,N_5537,N_4971);
nor U7423 (N_7423,N_5772,N_5744);
nand U7424 (N_7424,N_4843,N_5504);
and U7425 (N_7425,N_5902,N_5873);
or U7426 (N_7426,N_5410,N_5921);
or U7427 (N_7427,N_4721,N_4513);
or U7428 (N_7428,N_5079,N_4666);
xnor U7429 (N_7429,N_5340,N_5945);
nand U7430 (N_7430,N_5617,N_5568);
nand U7431 (N_7431,N_4645,N_5034);
and U7432 (N_7432,N_4729,N_4540);
or U7433 (N_7433,N_4508,N_5100);
nor U7434 (N_7434,N_5842,N_5246);
xor U7435 (N_7435,N_4778,N_5935);
nand U7436 (N_7436,N_4715,N_5203);
or U7437 (N_7437,N_4968,N_4842);
nand U7438 (N_7438,N_5228,N_5235);
nor U7439 (N_7439,N_4618,N_5543);
or U7440 (N_7440,N_5239,N_4681);
or U7441 (N_7441,N_5189,N_5524);
nand U7442 (N_7442,N_5997,N_5447);
nor U7443 (N_7443,N_5994,N_5132);
xnor U7444 (N_7444,N_5712,N_5580);
and U7445 (N_7445,N_5306,N_5205);
xor U7446 (N_7446,N_4937,N_5598);
nor U7447 (N_7447,N_5777,N_5520);
nand U7448 (N_7448,N_5986,N_5716);
xnor U7449 (N_7449,N_5985,N_5222);
xnor U7450 (N_7450,N_4935,N_5385);
nand U7451 (N_7451,N_5349,N_4988);
and U7452 (N_7452,N_5849,N_5938);
or U7453 (N_7453,N_5015,N_4617);
nor U7454 (N_7454,N_5852,N_4963);
nand U7455 (N_7455,N_4555,N_5181);
or U7456 (N_7456,N_5727,N_5391);
or U7457 (N_7457,N_5935,N_5760);
and U7458 (N_7458,N_4719,N_4905);
nand U7459 (N_7459,N_5786,N_5387);
and U7460 (N_7460,N_5991,N_5322);
and U7461 (N_7461,N_5432,N_4924);
nor U7462 (N_7462,N_4990,N_5971);
or U7463 (N_7463,N_5483,N_4695);
nor U7464 (N_7464,N_5477,N_4927);
or U7465 (N_7465,N_5650,N_5240);
xnor U7466 (N_7466,N_4798,N_4595);
and U7467 (N_7467,N_5566,N_5110);
nor U7468 (N_7468,N_4600,N_5017);
or U7469 (N_7469,N_5746,N_4941);
xor U7470 (N_7470,N_5236,N_4716);
or U7471 (N_7471,N_5494,N_4966);
and U7472 (N_7472,N_4813,N_4642);
nor U7473 (N_7473,N_5652,N_4677);
and U7474 (N_7474,N_5241,N_5628);
nor U7475 (N_7475,N_5493,N_5019);
or U7476 (N_7476,N_5363,N_5196);
nand U7477 (N_7477,N_5089,N_5280);
or U7478 (N_7478,N_5587,N_5298);
or U7479 (N_7479,N_5145,N_5723);
or U7480 (N_7480,N_5597,N_5960);
or U7481 (N_7481,N_4909,N_5396);
xnor U7482 (N_7482,N_4877,N_5257);
nor U7483 (N_7483,N_4744,N_5354);
and U7484 (N_7484,N_5939,N_4669);
or U7485 (N_7485,N_5921,N_5178);
or U7486 (N_7486,N_4881,N_4523);
xor U7487 (N_7487,N_5369,N_4687);
xor U7488 (N_7488,N_5109,N_5146);
or U7489 (N_7489,N_5319,N_5439);
nor U7490 (N_7490,N_4969,N_4612);
or U7491 (N_7491,N_4776,N_5030);
nor U7492 (N_7492,N_5404,N_5196);
nand U7493 (N_7493,N_4679,N_4995);
and U7494 (N_7494,N_5631,N_5785);
or U7495 (N_7495,N_4941,N_5600);
xor U7496 (N_7496,N_5968,N_4858);
nor U7497 (N_7497,N_5433,N_4518);
nor U7498 (N_7498,N_5503,N_5007);
and U7499 (N_7499,N_4612,N_4923);
nand U7500 (N_7500,N_6901,N_6462);
and U7501 (N_7501,N_7174,N_6861);
or U7502 (N_7502,N_6488,N_7270);
or U7503 (N_7503,N_6438,N_6599);
xnor U7504 (N_7504,N_7463,N_7362);
nand U7505 (N_7505,N_6848,N_6294);
or U7506 (N_7506,N_6543,N_7244);
nor U7507 (N_7507,N_7494,N_7460);
or U7508 (N_7508,N_6273,N_6692);
nand U7509 (N_7509,N_6963,N_6023);
nor U7510 (N_7510,N_7208,N_7262);
xnor U7511 (N_7511,N_6349,N_7311);
nand U7512 (N_7512,N_6869,N_6034);
nand U7513 (N_7513,N_6914,N_7221);
nand U7514 (N_7514,N_6479,N_7060);
or U7515 (N_7515,N_6474,N_6899);
xnor U7516 (N_7516,N_6766,N_6918);
and U7517 (N_7517,N_6062,N_6633);
and U7518 (N_7518,N_6293,N_7128);
and U7519 (N_7519,N_7374,N_6335);
or U7520 (N_7520,N_7031,N_6376);
nor U7521 (N_7521,N_6594,N_7384);
nand U7522 (N_7522,N_6454,N_6206);
nor U7523 (N_7523,N_6443,N_7442);
or U7524 (N_7524,N_6384,N_6976);
nand U7525 (N_7525,N_7102,N_7258);
and U7526 (N_7526,N_6211,N_6290);
and U7527 (N_7527,N_6671,N_6910);
and U7528 (N_7528,N_7488,N_6398);
xnor U7529 (N_7529,N_7487,N_6656);
or U7530 (N_7530,N_6455,N_6031);
nand U7531 (N_7531,N_6683,N_7201);
nand U7532 (N_7532,N_7429,N_6318);
xor U7533 (N_7533,N_6202,N_6077);
nand U7534 (N_7534,N_7329,N_7180);
and U7535 (N_7535,N_6597,N_7295);
or U7536 (N_7536,N_6020,N_6321);
and U7537 (N_7537,N_6965,N_6761);
nor U7538 (N_7538,N_6055,N_7004);
and U7539 (N_7539,N_6471,N_7432);
or U7540 (N_7540,N_6285,N_7039);
nand U7541 (N_7541,N_6138,N_6934);
nor U7542 (N_7542,N_6612,N_6307);
nand U7543 (N_7543,N_6857,N_6151);
and U7544 (N_7544,N_7300,N_6801);
nor U7545 (N_7545,N_7294,N_7019);
and U7546 (N_7546,N_7451,N_6047);
nor U7547 (N_7547,N_6448,N_7088);
or U7548 (N_7548,N_6267,N_6340);
or U7549 (N_7549,N_6859,N_6281);
nor U7550 (N_7550,N_6542,N_7469);
and U7551 (N_7551,N_7217,N_6070);
or U7552 (N_7552,N_6547,N_7117);
or U7553 (N_7553,N_7145,N_6263);
xnor U7554 (N_7554,N_6684,N_6163);
xnor U7555 (N_7555,N_6064,N_6527);
nor U7556 (N_7556,N_6170,N_6200);
nand U7557 (N_7557,N_7379,N_7148);
or U7558 (N_7558,N_6514,N_6646);
or U7559 (N_7559,N_6977,N_6484);
nand U7560 (N_7560,N_7055,N_6229);
nand U7561 (N_7561,N_7395,N_6639);
nand U7562 (N_7562,N_6722,N_7257);
nand U7563 (N_7563,N_6103,N_6213);
nand U7564 (N_7564,N_6305,N_6887);
or U7565 (N_7565,N_6003,N_7333);
nand U7566 (N_7566,N_6939,N_6092);
xnor U7567 (N_7567,N_7144,N_7116);
nor U7568 (N_7568,N_6112,N_6751);
xor U7569 (N_7569,N_6670,N_6736);
nand U7570 (N_7570,N_6541,N_6711);
nand U7571 (N_7571,N_6350,N_6578);
and U7572 (N_7572,N_6951,N_7169);
nand U7573 (N_7573,N_6571,N_7010);
nand U7574 (N_7574,N_6357,N_6962);
and U7575 (N_7575,N_7302,N_6396);
and U7576 (N_7576,N_6348,N_7313);
xnor U7577 (N_7577,N_6014,N_6109);
nand U7578 (N_7578,N_7438,N_7465);
or U7579 (N_7579,N_6368,N_6703);
nor U7580 (N_7580,N_7413,N_6416);
nand U7581 (N_7581,N_7236,N_6157);
or U7582 (N_7582,N_6605,N_7296);
or U7583 (N_7583,N_7334,N_7297);
or U7584 (N_7584,N_6695,N_7479);
nand U7585 (N_7585,N_6576,N_6071);
and U7586 (N_7586,N_7011,N_6943);
nand U7587 (N_7587,N_6940,N_6386);
nand U7588 (N_7588,N_6372,N_6166);
and U7589 (N_7589,N_6775,N_6572);
nand U7590 (N_7590,N_6570,N_6135);
and U7591 (N_7591,N_6422,N_6993);
and U7592 (N_7592,N_6247,N_6622);
or U7593 (N_7593,N_6126,N_7445);
nand U7594 (N_7594,N_7209,N_7133);
nor U7595 (N_7595,N_6179,N_6816);
and U7596 (N_7596,N_7285,N_7471);
nand U7597 (N_7597,N_6378,N_7301);
xor U7598 (N_7598,N_6959,N_6352);
or U7599 (N_7599,N_7363,N_6851);
nor U7600 (N_7600,N_6090,N_6041);
nor U7601 (N_7601,N_7357,N_7498);
nand U7602 (N_7602,N_7415,N_6905);
or U7603 (N_7603,N_6193,N_6391);
nand U7604 (N_7604,N_6926,N_7430);
nand U7605 (N_7605,N_6012,N_6282);
nor U7606 (N_7606,N_7085,N_6043);
or U7607 (N_7607,N_6536,N_7020);
nand U7608 (N_7608,N_7271,N_7204);
and U7609 (N_7609,N_7153,N_6116);
and U7610 (N_7610,N_6088,N_6158);
and U7611 (N_7611,N_6850,N_7084);
nor U7612 (N_7612,N_7110,N_6026);
and U7613 (N_7613,N_7380,N_7326);
or U7614 (N_7614,N_6203,N_6098);
nand U7615 (N_7615,N_7407,N_7224);
xor U7616 (N_7616,N_6945,N_6727);
nand U7617 (N_7617,N_7017,N_6145);
nor U7618 (N_7618,N_6373,N_6768);
or U7619 (N_7619,N_6207,N_7072);
and U7620 (N_7620,N_6436,N_7260);
nor U7621 (N_7621,N_6573,N_6925);
or U7622 (N_7622,N_6363,N_7067);
nor U7623 (N_7623,N_6440,N_6936);
or U7624 (N_7624,N_7437,N_7276);
or U7625 (N_7625,N_6171,N_6081);
and U7626 (N_7626,N_7192,N_7477);
and U7627 (N_7627,N_6555,N_6245);
nor U7628 (N_7628,N_6383,N_6623);
or U7629 (N_7629,N_6688,N_6666);
or U7630 (N_7630,N_6819,N_6029);
xor U7631 (N_7631,N_6094,N_7279);
nor U7632 (N_7632,N_7472,N_6676);
nor U7633 (N_7633,N_6678,N_6338);
or U7634 (N_7634,N_6968,N_7023);
nand U7635 (N_7635,N_6655,N_6627);
nor U7636 (N_7636,N_6818,N_7486);
xor U7637 (N_7637,N_6878,N_6563);
nor U7638 (N_7638,N_7495,N_6526);
xnor U7639 (N_7639,N_6565,N_6843);
nand U7640 (N_7640,N_6365,N_6786);
and U7641 (N_7641,N_6824,N_6217);
nor U7642 (N_7642,N_7417,N_6325);
nand U7643 (N_7643,N_7228,N_7408);
nor U7644 (N_7644,N_7149,N_6564);
xnor U7645 (N_7645,N_6212,N_6304);
or U7646 (N_7646,N_6482,N_6492);
nand U7647 (N_7647,N_6913,N_7125);
or U7648 (N_7648,N_6520,N_6517);
nor U7649 (N_7649,N_7012,N_7254);
nand U7650 (N_7650,N_6615,N_6499);
or U7651 (N_7651,N_6010,N_6310);
nor U7652 (N_7652,N_6328,N_6035);
or U7653 (N_7653,N_7284,N_6250);
nand U7654 (N_7654,N_6449,N_6429);
or U7655 (N_7655,N_7016,N_6297);
and U7656 (N_7656,N_6353,N_6214);
and U7657 (N_7657,N_7150,N_7218);
or U7658 (N_7658,N_7058,N_6370);
or U7659 (N_7659,N_6574,N_6985);
and U7660 (N_7660,N_6510,N_6280);
nor U7661 (N_7661,N_6792,N_6377);
nand U7662 (N_7662,N_7062,N_7327);
nand U7663 (N_7663,N_6235,N_6039);
or U7664 (N_7664,N_6518,N_7075);
and U7665 (N_7665,N_7410,N_6485);
and U7666 (N_7666,N_7111,N_6425);
or U7667 (N_7667,N_7159,N_7354);
and U7668 (N_7668,N_6345,N_7216);
or U7669 (N_7669,N_6466,N_7426);
nand U7670 (N_7670,N_6292,N_6960);
and U7671 (N_7671,N_7389,N_6949);
nand U7672 (N_7672,N_7423,N_6053);
and U7673 (N_7673,N_7307,N_6967);
and U7674 (N_7674,N_6649,N_7483);
or U7675 (N_7675,N_7127,N_6681);
and U7676 (N_7676,N_7248,N_7092);
and U7677 (N_7677,N_6698,N_6731);
nor U7678 (N_7678,N_7286,N_6794);
and U7679 (N_7679,N_6065,N_6424);
xnor U7680 (N_7680,N_7086,N_7446);
and U7681 (N_7681,N_6826,N_6236);
and U7682 (N_7682,N_7398,N_7227);
nor U7683 (N_7683,N_7237,N_7203);
nand U7684 (N_7684,N_7319,N_6874);
nor U7685 (N_7685,N_6266,N_6067);
or U7686 (N_7686,N_6314,N_6008);
nor U7687 (N_7687,N_6210,N_6154);
or U7688 (N_7688,N_7443,N_6674);
and U7689 (N_7689,N_7142,N_6856);
and U7690 (N_7690,N_6537,N_6323);
nor U7691 (N_7691,N_6840,N_7391);
or U7692 (N_7692,N_6531,N_6833);
and U7693 (N_7693,N_6603,N_6707);
nand U7694 (N_7694,N_6994,N_7360);
nand U7695 (N_7695,N_7120,N_6456);
nand U7696 (N_7696,N_6439,N_6152);
or U7697 (N_7697,N_6495,N_6757);
nor U7698 (N_7698,N_7403,N_7259);
nand U7699 (N_7699,N_6734,N_6589);
and U7700 (N_7700,N_6891,N_6596);
nand U7701 (N_7701,N_6930,N_6693);
and U7702 (N_7702,N_6991,N_6453);
nor U7703 (N_7703,N_6789,N_7310);
or U7704 (N_7704,N_6287,N_6033);
or U7705 (N_7705,N_6477,N_6886);
or U7706 (N_7706,N_7318,N_7137);
nor U7707 (N_7707,N_7378,N_6300);
xor U7708 (N_7708,N_6953,N_6700);
or U7709 (N_7709,N_6701,N_6421);
nor U7710 (N_7710,N_7015,N_6607);
or U7711 (N_7711,N_7467,N_7045);
nand U7712 (N_7712,N_7404,N_7365);
and U7713 (N_7713,N_6276,N_6868);
nand U7714 (N_7714,N_6097,N_6919);
and U7715 (N_7715,N_6972,N_6224);
xnor U7716 (N_7716,N_6189,N_6739);
and U7717 (N_7717,N_6941,N_7230);
nand U7718 (N_7718,N_6123,N_7104);
nand U7719 (N_7719,N_6955,N_7372);
nand U7720 (N_7720,N_6557,N_6277);
nand U7721 (N_7721,N_7298,N_6264);
or U7722 (N_7722,N_7397,N_6144);
and U7723 (N_7723,N_6710,N_7195);
or U7724 (N_7724,N_7275,N_7118);
nand U7725 (N_7725,N_6028,N_6269);
or U7726 (N_7726,N_6044,N_7419);
and U7727 (N_7727,N_6491,N_7197);
nor U7728 (N_7728,N_6654,N_7478);
nand U7729 (N_7729,N_7177,N_6301);
or U7730 (N_7730,N_6246,N_6476);
nand U7731 (N_7731,N_6938,N_6446);
nand U7732 (N_7732,N_6602,N_6842);
nor U7733 (N_7733,N_6942,N_6162);
or U7734 (N_7734,N_6244,N_7210);
and U7735 (N_7735,N_7124,N_6347);
nand U7736 (N_7736,N_6590,N_7416);
nor U7737 (N_7737,N_6503,N_7324);
or U7738 (N_7738,N_6897,N_6129);
or U7739 (N_7739,N_6497,N_7079);
xor U7740 (N_7740,N_6430,N_7074);
nand U7741 (N_7741,N_6853,N_6120);
and U7742 (N_7742,N_6782,N_7350);
nor U7743 (N_7743,N_6445,N_6185);
or U7744 (N_7744,N_6278,N_7029);
or U7745 (N_7745,N_6176,N_6830);
nor U7746 (N_7746,N_6755,N_7038);
nor U7747 (N_7747,N_6355,N_6558);
nand U7748 (N_7748,N_7049,N_6645);
nor U7749 (N_7749,N_6005,N_6876);
and U7750 (N_7750,N_6303,N_6101);
nand U7751 (N_7751,N_7033,N_6146);
xnor U7752 (N_7752,N_7249,N_7400);
and U7753 (N_7753,N_6772,N_6275);
nor U7754 (N_7754,N_6399,N_6360);
nand U7755 (N_7755,N_7123,N_7164);
or U7756 (N_7756,N_6356,N_6880);
or U7757 (N_7757,N_6545,N_6911);
nand U7758 (N_7758,N_6450,N_6616);
and U7759 (N_7759,N_6296,N_6270);
nand U7760 (N_7760,N_6773,N_6132);
nand U7761 (N_7761,N_7129,N_7476);
nand U7762 (N_7762,N_6327,N_6004);
nand U7763 (N_7763,N_6872,N_7273);
nor U7764 (N_7764,N_6617,N_7185);
nand U7765 (N_7765,N_7348,N_6877);
nand U7766 (N_7766,N_6444,N_6999);
and U7767 (N_7767,N_6342,N_7421);
xnor U7768 (N_7768,N_6408,N_7027);
or U7769 (N_7769,N_6458,N_7394);
nand U7770 (N_7770,N_6756,N_6242);
nand U7771 (N_7771,N_7042,N_7063);
xor U7772 (N_7772,N_6660,N_6435);
nor U7773 (N_7773,N_6253,N_7261);
xor U7774 (N_7774,N_6316,N_7005);
nor U7775 (N_7775,N_6778,N_7156);
xnor U7776 (N_7776,N_6511,N_6637);
nand U7777 (N_7777,N_6460,N_6420);
nor U7778 (N_7778,N_6080,N_6733);
and U7779 (N_7779,N_6036,N_6330);
nand U7780 (N_7780,N_6845,N_6587);
nor U7781 (N_7781,N_7482,N_7346);
or U7782 (N_7782,N_6410,N_7194);
and U7783 (N_7783,N_6238,N_6986);
and U7784 (N_7784,N_6762,N_6401);
nor U7785 (N_7785,N_7061,N_6837);
and U7786 (N_7786,N_7337,N_6337);
nor U7787 (N_7787,N_6898,N_7414);
and U7788 (N_7788,N_7096,N_7205);
nor U7789 (N_7789,N_6659,N_6793);
nor U7790 (N_7790,N_6204,N_6920);
and U7791 (N_7791,N_6192,N_7200);
or U7792 (N_7792,N_7351,N_6172);
and U7793 (N_7793,N_6021,N_6716);
or U7794 (N_7794,N_6174,N_6873);
or U7795 (N_7795,N_6298,N_7054);
xnor U7796 (N_7796,N_6932,N_7453);
and U7797 (N_7797,N_6480,N_6746);
and U7798 (N_7798,N_7048,N_6073);
and U7799 (N_7799,N_6165,N_6630);
nand U7800 (N_7800,N_7490,N_6744);
or U7801 (N_7801,N_6251,N_7047);
and U7802 (N_7802,N_6268,N_7225);
nor U7803 (N_7803,N_7368,N_6205);
nand U7804 (N_7804,N_6539,N_6506);
xor U7805 (N_7805,N_6709,N_7383);
and U7806 (N_7806,N_7293,N_7462);
nand U7807 (N_7807,N_6863,N_6087);
nor U7808 (N_7808,N_6767,N_6486);
nand U7809 (N_7809,N_7080,N_6608);
or U7810 (N_7810,N_6001,N_6127);
nand U7811 (N_7811,N_6504,N_6980);
or U7812 (N_7812,N_6956,N_7401);
nor U7813 (N_7813,N_7024,N_6075);
and U7814 (N_7814,N_7190,N_6704);
or U7815 (N_7815,N_6423,N_6817);
or U7816 (N_7816,N_6626,N_6802);
nor U7817 (N_7817,N_7214,N_6069);
nor U7818 (N_7818,N_6351,N_6361);
nand U7819 (N_7819,N_6631,N_6760);
nand U7820 (N_7820,N_7154,N_7459);
xnor U7821 (N_7821,N_7040,N_7412);
nand U7822 (N_7822,N_6946,N_6125);
nor U7823 (N_7823,N_6289,N_6395);
nand U7824 (N_7824,N_6196,N_6796);
nand U7825 (N_7825,N_6218,N_6969);
nor U7826 (N_7826,N_6379,N_6291);
or U7827 (N_7827,N_6983,N_7436);
nand U7828 (N_7828,N_6359,N_6550);
and U7829 (N_7829,N_6326,N_6821);
nor U7830 (N_7830,N_6839,N_6992);
and U7831 (N_7831,N_7339,N_7331);
and U7832 (N_7832,N_6134,N_7375);
or U7833 (N_7833,N_6647,N_6180);
or U7834 (N_7834,N_6343,N_7497);
nor U7835 (N_7835,N_6588,N_7424);
and U7836 (N_7836,N_7114,N_6417);
and U7837 (N_7837,N_6642,N_6534);
nand U7838 (N_7838,N_6388,N_6459);
and U7839 (N_7839,N_6513,N_7255);
nand U7840 (N_7840,N_6686,N_6791);
nor U7841 (N_7841,N_7172,N_7247);
nand U7842 (N_7842,N_7441,N_7387);
and U7843 (N_7843,N_6387,N_6078);
xor U7844 (N_7844,N_7392,N_6650);
nor U7845 (N_7845,N_7252,N_6159);
or U7846 (N_7846,N_6825,N_6182);
or U7847 (N_7847,N_7002,N_6810);
xnor U7848 (N_7848,N_7312,N_6827);
and U7849 (N_7849,N_6128,N_7233);
or U7850 (N_7850,N_6283,N_7468);
and U7851 (N_7851,N_6974,N_7157);
or U7852 (N_7852,N_6795,N_6059);
nor U7853 (N_7853,N_6519,N_6334);
or U7854 (N_7854,N_6544,N_7347);
nor U7855 (N_7855,N_6765,N_6705);
or U7856 (N_7856,N_6183,N_6262);
and U7857 (N_7857,N_7323,N_6600);
and U7858 (N_7858,N_7458,N_6892);
and U7859 (N_7859,N_6759,N_7034);
nor U7860 (N_7860,N_6917,N_6089);
nand U7861 (N_7861,N_6066,N_7282);
and U7862 (N_7862,N_6699,N_6105);
nand U7863 (N_7863,N_6742,N_6528);
nand U7864 (N_7864,N_6916,N_6111);
nor U7865 (N_7865,N_7189,N_6494);
and U7866 (N_7866,N_6288,N_6255);
or U7867 (N_7867,N_6011,N_7399);
nor U7868 (N_7868,N_6346,N_7030);
xor U7869 (N_7869,N_7455,N_7178);
or U7870 (N_7870,N_6516,N_7130);
xor U7871 (N_7871,N_6774,N_6753);
nor U7872 (N_7872,N_6988,N_6809);
nor U7873 (N_7873,N_6621,N_6836);
xnor U7874 (N_7874,N_7376,N_6852);
and U7875 (N_7875,N_7349,N_6052);
nor U7876 (N_7876,N_6997,N_6451);
or U7877 (N_7877,N_6694,N_6952);
nand U7878 (N_7878,N_7448,N_6770);
and U7879 (N_7879,N_6643,N_6331);
and U7880 (N_7880,N_7167,N_6858);
nor U7881 (N_7881,N_7435,N_6849);
nor U7882 (N_7882,N_6725,N_7449);
and U7883 (N_7883,N_6136,N_6981);
nand U7884 (N_7884,N_6382,N_6585);
and U7885 (N_7885,N_6505,N_6258);
nand U7886 (N_7886,N_6726,N_6815);
nand U7887 (N_7887,N_6016,N_6640);
nor U7888 (N_7888,N_7263,N_6056);
or U7889 (N_7889,N_6048,N_6613);
and U7890 (N_7890,N_7143,N_7340);
or U7891 (N_7891,N_6119,N_7089);
or U7892 (N_7892,N_6632,N_6045);
xor U7893 (N_7893,N_6604,N_6978);
nor U7894 (N_7894,N_7095,N_7053);
nor U7895 (N_7895,N_6906,N_6117);
or U7896 (N_7896,N_7121,N_7277);
and U7897 (N_7897,N_7139,N_6593);
and U7898 (N_7898,N_7485,N_6635);
nor U7899 (N_7899,N_7068,N_7489);
nand U7900 (N_7900,N_6114,N_7115);
or U7901 (N_7901,N_6478,N_7160);
nand U7902 (N_7902,N_6783,N_6764);
and U7903 (N_7903,N_7094,N_6142);
and U7904 (N_7904,N_7059,N_6822);
nor U7905 (N_7905,N_6405,N_6175);
and U7906 (N_7906,N_7343,N_6864);
nor U7907 (N_7907,N_7266,N_7454);
nand U7908 (N_7908,N_6489,N_6261);
or U7909 (N_7909,N_6583,N_6788);
and U7910 (N_7910,N_7132,N_7251);
nand U7911 (N_7911,N_6611,N_6638);
nand U7912 (N_7912,N_7099,N_7168);
nand U7913 (N_7913,N_7207,N_6561);
or U7914 (N_7914,N_6274,N_6402);
and U7915 (N_7915,N_6560,N_7256);
nand U7916 (N_7916,N_6222,N_6051);
nand U7917 (N_7917,N_6260,N_7308);
nor U7918 (N_7918,N_6618,N_6083);
nor U7919 (N_7919,N_6535,N_6890);
nor U7920 (N_7920,N_6173,N_7288);
or U7921 (N_7921,N_6644,N_7272);
nor U7922 (N_7922,N_6835,N_6271);
nor U7923 (N_7923,N_6964,N_6149);
nand U7924 (N_7924,N_6970,N_6664);
and U7925 (N_7925,N_6341,N_7182);
xor U7926 (N_7926,N_6893,N_6721);
nor U7927 (N_7927,N_7355,N_6168);
and U7928 (N_7928,N_6496,N_6812);
nor U7929 (N_7929,N_6050,N_7161);
xor U7930 (N_7930,N_6332,N_6061);
nand U7931 (N_7931,N_7014,N_7332);
xnor U7932 (N_7932,N_6362,N_7141);
nor U7933 (N_7933,N_7364,N_6808);
nand U7934 (N_7934,N_6322,N_7071);
nand U7935 (N_7935,N_6225,N_6257);
and U7936 (N_7936,N_7371,N_6024);
or U7937 (N_7937,N_6641,N_6820);
or U7938 (N_7938,N_6995,N_6829);
and U7939 (N_7939,N_6216,N_7215);
or U7940 (N_7940,N_7396,N_6201);
and U7941 (N_7941,N_6115,N_6164);
and U7942 (N_7942,N_6883,N_6404);
and U7943 (N_7943,N_7165,N_6702);
nand U7944 (N_7944,N_7037,N_6312);
nor U7945 (N_7945,N_6961,N_7474);
xnor U7946 (N_7946,N_6745,N_7166);
or U7947 (N_7947,N_7290,N_6191);
or U7948 (N_7948,N_7425,N_6614);
nor U7949 (N_7949,N_6344,N_7191);
nand U7950 (N_7950,N_7352,N_7051);
nand U7951 (N_7951,N_6018,N_7325);
nand U7952 (N_7952,N_7105,N_6254);
nand U7953 (N_7953,N_7093,N_6530);
xnor U7954 (N_7954,N_6900,N_7280);
nor U7955 (N_7955,N_7283,N_6668);
nand U7956 (N_7956,N_6975,N_6195);
xnor U7957 (N_7957,N_6592,N_6091);
nand U7958 (N_7958,N_6524,N_7341);
or U7959 (N_7959,N_7292,N_6186);
nand U7960 (N_7960,N_6426,N_6881);
and U7961 (N_7961,N_6380,N_6996);
or U7962 (N_7962,N_6990,N_7220);
nand U7963 (N_7963,N_7078,N_7278);
or U7964 (N_7964,N_7381,N_6629);
nor U7965 (N_7965,N_6928,N_6501);
nor U7966 (N_7966,N_6823,N_6375);
and U7967 (N_7967,N_6885,N_6190);
nand U7968 (N_7968,N_7119,N_6777);
nor U7969 (N_7969,N_6256,N_6844);
and U7970 (N_7970,N_6769,N_6807);
nor U7971 (N_7971,N_7480,N_6625);
or U7972 (N_7972,N_7028,N_6009);
xnor U7973 (N_7973,N_7193,N_7299);
or U7974 (N_7974,N_7101,N_6237);
and U7975 (N_7975,N_6086,N_6776);
nand U7976 (N_7976,N_6228,N_6966);
or U7977 (N_7977,N_6030,N_6971);
nand U7978 (N_7978,N_6933,N_6669);
nor U7979 (N_7979,N_6118,N_6636);
and U7980 (N_7980,N_6813,N_6317);
nor U7981 (N_7981,N_7083,N_6884);
and U7982 (N_7982,N_7036,N_6427);
nor U7983 (N_7983,N_6130,N_7253);
nor U7984 (N_7984,N_7183,N_7131);
or U7985 (N_7985,N_6329,N_6046);
and U7986 (N_7986,N_6441,N_7065);
nor U7987 (N_7987,N_6133,N_6309);
or U7988 (N_7988,N_6469,N_7493);
xnor U7989 (N_7989,N_7171,N_6598);
nand U7990 (N_7990,N_6921,N_7238);
or U7991 (N_7991,N_7491,N_6806);
xor U7992 (N_7992,N_7428,N_6232);
nor U7993 (N_7993,N_6832,N_6279);
nor U7994 (N_7994,N_6060,N_6935);
or U7995 (N_7995,N_6706,N_6568);
and U7996 (N_7996,N_6068,N_7212);
or U7997 (N_7997,N_6099,N_6582);
nor U7998 (N_7998,N_7473,N_6467);
and U7999 (N_7999,N_6548,N_6306);
or U8000 (N_8000,N_7450,N_6140);
nand U8001 (N_8001,N_7229,N_7082);
and U8002 (N_8002,N_6866,N_7440);
nor U8003 (N_8003,N_6392,N_7064);
or U8004 (N_8004,N_6634,N_6006);
nand U8005 (N_8005,N_6139,N_7052);
or U8006 (N_8006,N_6367,N_7335);
xor U8007 (N_8007,N_6673,N_6400);
nor U8008 (N_8008,N_6790,N_6025);
nor U8009 (N_8009,N_6998,N_6481);
nor U8010 (N_8010,N_6834,N_7175);
and U8011 (N_8011,N_6187,N_6743);
and U8012 (N_8012,N_6708,N_6085);
or U8013 (N_8013,N_6336,N_6754);
or U8014 (N_8014,N_7385,N_7187);
nor U8015 (N_8015,N_7211,N_6084);
nor U8016 (N_8016,N_6687,N_7402);
xor U8017 (N_8017,N_6908,N_6562);
and U8018 (N_8018,N_6882,N_6740);
nor U8019 (N_8019,N_6803,N_6723);
and U8020 (N_8020,N_6389,N_7136);
nor U8021 (N_8021,N_6575,N_7098);
nand U8022 (N_8022,N_7321,N_6780);
or U8023 (N_8023,N_6272,N_7070);
or U8024 (N_8024,N_7274,N_7170);
or U8025 (N_8025,N_6896,N_6680);
nor U8026 (N_8026,N_6160,N_6567);
and U8027 (N_8027,N_6601,N_7241);
xor U8028 (N_8028,N_6093,N_7044);
nand U8029 (N_8029,N_6369,N_6371);
and U8030 (N_8030,N_6197,N_6374);
nand U8031 (N_8031,N_7289,N_7000);
nand U8032 (N_8032,N_7138,N_7032);
and U8033 (N_8033,N_7222,N_6779);
or U8034 (N_8034,N_6784,N_7370);
or U8035 (N_8035,N_6063,N_6464);
nor U8036 (N_8036,N_6434,N_7135);
or U8037 (N_8037,N_6177,N_6735);
nor U8038 (N_8038,N_7305,N_6624);
or U8039 (N_8039,N_6320,N_6027);
or U8040 (N_8040,N_6937,N_6239);
or U8041 (N_8041,N_6233,N_6958);
nand U8042 (N_8042,N_6082,N_7345);
nand U8043 (N_8043,N_7091,N_6651);
and U8044 (N_8044,N_6414,N_7240);
xor U8045 (N_8045,N_7317,N_6929);
or U8046 (N_8046,N_6652,N_6865);
nand U8047 (N_8047,N_6227,N_6220);
or U8048 (N_8048,N_6619,N_6483);
xnor U8049 (N_8049,N_7366,N_6606);
and U8050 (N_8050,N_7434,N_6691);
nand U8051 (N_8051,N_6781,N_6302);
and U8052 (N_8052,N_6552,N_6493);
xnor U8053 (N_8053,N_7353,N_7390);
nand U8054 (N_8054,N_6717,N_6797);
nand U8055 (N_8055,N_6209,N_6104);
nor U8056 (N_8056,N_6465,N_6319);
or U8057 (N_8057,N_7322,N_7418);
nor U8058 (N_8058,N_7179,N_7219);
and U8059 (N_8059,N_6428,N_6749);
and U8060 (N_8060,N_6143,N_7202);
nand U8061 (N_8061,N_6591,N_7134);
xnor U8062 (N_8062,N_6131,N_7320);
nand U8063 (N_8063,N_6032,N_6903);
or U8064 (N_8064,N_6313,N_7267);
and U8065 (N_8065,N_6931,N_6248);
and U8066 (N_8066,N_6831,N_7050);
nand U8067 (N_8067,N_7043,N_7231);
and U8068 (N_8068,N_6973,N_6199);
and U8069 (N_8069,N_6719,N_7361);
nor U8070 (N_8070,N_6049,N_6713);
nor U8071 (N_8071,N_6000,N_7268);
and U8072 (N_8072,N_7126,N_6141);
nand U8073 (N_8073,N_7386,N_7213);
and U8074 (N_8074,N_7106,N_6690);
nand U8075 (N_8075,N_6533,N_6390);
nor U8076 (N_8076,N_6580,N_6894);
xnor U8077 (N_8077,N_7492,N_6787);
and U8078 (N_8078,N_6718,N_6512);
and U8079 (N_8079,N_6912,N_6595);
and U8080 (N_8080,N_7367,N_6240);
and U8081 (N_8081,N_6226,N_6546);
nor U8082 (N_8082,N_7007,N_7470);
xor U8083 (N_8083,N_6286,N_7081);
or U8084 (N_8084,N_6667,N_6752);
or U8085 (N_8085,N_6947,N_7496);
or U8086 (N_8086,N_6811,N_6663);
xor U8087 (N_8087,N_7265,N_6747);
nor U8088 (N_8088,N_6989,N_7336);
nand U8089 (N_8089,N_6521,N_7109);
nand U8090 (N_8090,N_6750,N_6665);
nand U8091 (N_8091,N_6072,N_7181);
xnor U8092 (N_8092,N_6184,N_7239);
nand U8093 (N_8093,N_6074,N_6463);
nand U8094 (N_8094,N_6771,N_6532);
and U8095 (N_8095,N_6411,N_7411);
or U8096 (N_8096,N_7427,N_6231);
nor U8097 (N_8097,N_6540,N_6737);
xnor U8098 (N_8098,N_6662,N_6556);
or U8099 (N_8099,N_7108,N_6358);
nor U8100 (N_8100,N_6879,N_6037);
and U8101 (N_8101,N_6208,N_6161);
or U8102 (N_8102,N_7309,N_6040);
or U8103 (N_8103,N_7306,N_6324);
or U8104 (N_8104,N_6846,N_6798);
nor U8105 (N_8105,N_6509,N_6311);
and U8106 (N_8106,N_6847,N_6418);
and U8107 (N_8107,N_6549,N_6895);
nor U8108 (N_8108,N_6019,N_6498);
nand U8109 (N_8109,N_6923,N_6814);
and U8110 (N_8110,N_6113,N_6354);
nor U8111 (N_8111,N_6017,N_6672);
or U8112 (N_8112,N_6508,N_6522);
xor U8113 (N_8113,N_7420,N_6147);
nor U8114 (N_8114,N_6339,N_6473);
nand U8115 (N_8115,N_7338,N_7382);
or U8116 (N_8116,N_6732,N_6584);
nand U8117 (N_8117,N_7146,N_6433);
nand U8118 (N_8118,N_6538,N_6393);
nor U8119 (N_8119,N_7107,N_6038);
nand U8120 (N_8120,N_7235,N_6106);
or U8121 (N_8121,N_6121,N_7499);
and U8122 (N_8122,N_7439,N_7393);
nor U8123 (N_8123,N_6295,N_6366);
nand U8124 (N_8124,N_6076,N_7484);
and U8125 (N_8125,N_6107,N_7147);
and U8126 (N_8126,N_7199,N_6249);
and U8127 (N_8127,N_6551,N_6153);
and U8128 (N_8128,N_7069,N_7155);
nand U8129 (N_8129,N_6241,N_7008);
and U8130 (N_8130,N_7316,N_6577);
or U8131 (N_8131,N_6252,N_6730);
nor U8132 (N_8132,N_6490,N_6927);
nand U8133 (N_8133,N_6299,N_7206);
or U8134 (N_8134,N_7073,N_7328);
nor U8135 (N_8135,N_7163,N_6167);
or U8136 (N_8136,N_7006,N_6862);
and U8137 (N_8137,N_6394,N_7461);
nor U8138 (N_8138,N_6397,N_6658);
xnor U8139 (N_8139,N_6738,N_6432);
nand U8140 (N_8140,N_6515,N_7388);
and U8141 (N_8141,N_7475,N_6875);
nor U8142 (N_8142,N_6137,N_6169);
and U8143 (N_8143,N_7291,N_6715);
nor U8144 (N_8144,N_6675,N_6696);
and U8145 (N_8145,N_6922,N_7264);
nor U8146 (N_8146,N_7287,N_7003);
xor U8147 (N_8147,N_6419,N_7444);
or U8148 (N_8148,N_6315,N_7377);
nand U8149 (N_8149,N_7242,N_6855);
nor U8150 (N_8150,N_6265,N_7041);
or U8151 (N_8151,N_7025,N_6924);
nand U8152 (N_8152,N_6333,N_6661);
or U8153 (N_8153,N_6569,N_6219);
or U8154 (N_8154,N_6215,N_6785);
nand U8155 (N_8155,N_6472,N_6487);
nor U8156 (N_8156,N_6697,N_6867);
and U8157 (N_8157,N_7406,N_6712);
and U8158 (N_8158,N_6554,N_6415);
xor U8159 (N_8159,N_7481,N_6407);
xor U8160 (N_8160,N_7369,N_6799);
nor U8161 (N_8161,N_7358,N_7184);
nand U8162 (N_8162,N_7122,N_6648);
nand U8163 (N_8163,N_7176,N_6860);
nor U8164 (N_8164,N_6741,N_6800);
and U8165 (N_8165,N_7113,N_7359);
nand U8166 (N_8166,N_7356,N_7269);
nor U8167 (N_8167,N_6308,N_6452);
nand U8168 (N_8168,N_6188,N_7303);
nor U8169 (N_8169,N_7022,N_7330);
or U8170 (N_8170,N_6724,N_7188);
nor U8171 (N_8171,N_7100,N_6944);
and U8172 (N_8172,N_6553,N_7246);
nand U8173 (N_8173,N_6748,N_6838);
nor U8174 (N_8174,N_6412,N_6096);
xor U8175 (N_8175,N_6230,N_7464);
nand U8176 (N_8176,N_7243,N_6653);
or U8177 (N_8177,N_7373,N_6364);
or U8178 (N_8178,N_7281,N_6610);
nand U8179 (N_8179,N_6628,N_7077);
and U8180 (N_8180,N_6181,N_7151);
nor U8181 (N_8181,N_6902,N_6502);
or U8182 (N_8182,N_6057,N_6156);
or U8183 (N_8183,N_7452,N_7342);
nor U8184 (N_8184,N_6682,N_6102);
nor U8185 (N_8185,N_6728,N_6679);
and U8186 (N_8186,N_6950,N_6108);
nand U8187 (N_8187,N_6870,N_7056);
nor U8188 (N_8188,N_6042,N_7066);
nand U8189 (N_8189,N_6403,N_7103);
xor U8190 (N_8190,N_6470,N_6178);
nor U8191 (N_8191,N_6475,N_6007);
and U8192 (N_8192,N_7405,N_6054);
or U8193 (N_8193,N_6854,N_6525);
nor U8194 (N_8194,N_6110,N_7431);
and U8195 (N_8195,N_6620,N_7009);
and U8196 (N_8196,N_7250,N_7422);
nand U8197 (N_8197,N_6948,N_6150);
nand U8198 (N_8198,N_7021,N_6058);
nand U8199 (N_8199,N_6442,N_6889);
nor U8200 (N_8200,N_6909,N_6579);
and U8201 (N_8201,N_6431,N_7026);
xnor U8202 (N_8202,N_6013,N_6984);
and U8203 (N_8203,N_6957,N_6406);
xnor U8204 (N_8204,N_6500,N_6915);
xor U8205 (N_8205,N_6015,N_7140);
nor U8206 (N_8206,N_6729,N_6888);
or U8207 (N_8207,N_7447,N_7226);
xnor U8208 (N_8208,N_6223,N_6804);
or U8209 (N_8209,N_7198,N_7001);
or U8210 (N_8210,N_7158,N_6982);
xor U8211 (N_8211,N_6409,N_6904);
or U8212 (N_8212,N_6689,N_7304);
xor U8213 (N_8213,N_7018,N_6720);
and U8214 (N_8214,N_6461,N_7173);
nor U8215 (N_8215,N_6507,N_7035);
nand U8216 (N_8216,N_6979,N_6437);
and U8217 (N_8217,N_7466,N_6657);
nor U8218 (N_8218,N_7456,N_7152);
or U8219 (N_8219,N_6566,N_6457);
nor U8220 (N_8220,N_6609,N_6841);
or U8221 (N_8221,N_6234,N_7013);
and U8222 (N_8222,N_7234,N_7087);
nand U8223 (N_8223,N_6259,N_6198);
or U8224 (N_8224,N_6221,N_6022);
nor U8225 (N_8225,N_6907,N_6581);
xnor U8226 (N_8226,N_6385,N_6559);
nor U8227 (N_8227,N_6523,N_6122);
and U8228 (N_8228,N_6758,N_6284);
and U8229 (N_8229,N_6381,N_7315);
nor U8230 (N_8230,N_7196,N_6468);
xor U8231 (N_8231,N_6805,N_7112);
nand U8232 (N_8232,N_7314,N_7046);
and U8233 (N_8233,N_6447,N_6685);
or U8234 (N_8234,N_7186,N_6714);
nor U8235 (N_8235,N_6828,N_7457);
nand U8236 (N_8236,N_6194,N_7223);
nor U8237 (N_8237,N_6155,N_6124);
nor U8238 (N_8238,N_7245,N_6079);
xnor U8239 (N_8239,N_6002,N_6954);
and U8240 (N_8240,N_7162,N_6100);
nand U8241 (N_8241,N_7097,N_7409);
nand U8242 (N_8242,N_6677,N_7433);
and U8243 (N_8243,N_6243,N_7232);
nand U8244 (N_8244,N_7076,N_6987);
xor U8245 (N_8245,N_6529,N_7090);
nand U8246 (N_8246,N_6413,N_6095);
or U8247 (N_8247,N_7057,N_6586);
nand U8248 (N_8248,N_7344,N_6148);
nand U8249 (N_8249,N_6763,N_6871);
and U8250 (N_8250,N_6515,N_6472);
nor U8251 (N_8251,N_6099,N_6872);
and U8252 (N_8252,N_6582,N_6318);
or U8253 (N_8253,N_7262,N_6068);
and U8254 (N_8254,N_6380,N_6649);
and U8255 (N_8255,N_7245,N_6437);
nand U8256 (N_8256,N_6150,N_6190);
and U8257 (N_8257,N_6535,N_7020);
or U8258 (N_8258,N_6483,N_6292);
or U8259 (N_8259,N_6138,N_7147);
or U8260 (N_8260,N_6512,N_7297);
nand U8261 (N_8261,N_7114,N_6671);
nor U8262 (N_8262,N_7270,N_6695);
nor U8263 (N_8263,N_6985,N_6154);
xnor U8264 (N_8264,N_7267,N_7212);
nand U8265 (N_8265,N_6126,N_6418);
nand U8266 (N_8266,N_6425,N_7405);
xor U8267 (N_8267,N_6486,N_6634);
xnor U8268 (N_8268,N_6461,N_6709);
nor U8269 (N_8269,N_7092,N_7093);
and U8270 (N_8270,N_6190,N_6620);
nor U8271 (N_8271,N_6103,N_7222);
nor U8272 (N_8272,N_6749,N_6448);
and U8273 (N_8273,N_6518,N_6913);
or U8274 (N_8274,N_6632,N_6602);
nand U8275 (N_8275,N_7371,N_6366);
nor U8276 (N_8276,N_7416,N_7011);
or U8277 (N_8277,N_6919,N_7491);
nand U8278 (N_8278,N_6880,N_6103);
and U8279 (N_8279,N_6474,N_7418);
nand U8280 (N_8280,N_6708,N_7131);
nand U8281 (N_8281,N_6728,N_6027);
nor U8282 (N_8282,N_6974,N_6098);
and U8283 (N_8283,N_7463,N_6938);
nand U8284 (N_8284,N_6332,N_6807);
or U8285 (N_8285,N_7106,N_7047);
and U8286 (N_8286,N_7245,N_6779);
nor U8287 (N_8287,N_6868,N_7052);
nor U8288 (N_8288,N_7369,N_6388);
nor U8289 (N_8289,N_6256,N_6549);
or U8290 (N_8290,N_7100,N_6964);
nand U8291 (N_8291,N_7140,N_6981);
and U8292 (N_8292,N_6968,N_6815);
nor U8293 (N_8293,N_6892,N_7385);
xnor U8294 (N_8294,N_7135,N_6503);
and U8295 (N_8295,N_6944,N_6806);
and U8296 (N_8296,N_6050,N_6765);
nor U8297 (N_8297,N_7448,N_6276);
xor U8298 (N_8298,N_6973,N_7257);
nor U8299 (N_8299,N_7423,N_6939);
nand U8300 (N_8300,N_6691,N_7272);
and U8301 (N_8301,N_7404,N_7132);
nand U8302 (N_8302,N_6859,N_6817);
or U8303 (N_8303,N_7138,N_7422);
or U8304 (N_8304,N_6503,N_6174);
nand U8305 (N_8305,N_6981,N_7378);
and U8306 (N_8306,N_6744,N_6098);
nor U8307 (N_8307,N_6194,N_6270);
or U8308 (N_8308,N_6471,N_6155);
nand U8309 (N_8309,N_6677,N_6125);
or U8310 (N_8310,N_6178,N_6919);
xor U8311 (N_8311,N_6309,N_6664);
nand U8312 (N_8312,N_6286,N_6852);
and U8313 (N_8313,N_6556,N_7390);
and U8314 (N_8314,N_6889,N_6381);
nand U8315 (N_8315,N_6077,N_6017);
or U8316 (N_8316,N_7227,N_7423);
nand U8317 (N_8317,N_6941,N_6523);
or U8318 (N_8318,N_6683,N_6732);
and U8319 (N_8319,N_6023,N_7424);
nand U8320 (N_8320,N_6890,N_6121);
or U8321 (N_8321,N_7253,N_7047);
nand U8322 (N_8322,N_7455,N_7291);
and U8323 (N_8323,N_7412,N_7365);
nand U8324 (N_8324,N_7163,N_7303);
and U8325 (N_8325,N_6916,N_6460);
nor U8326 (N_8326,N_6622,N_6784);
or U8327 (N_8327,N_6643,N_6946);
nand U8328 (N_8328,N_6890,N_6072);
nand U8329 (N_8329,N_6475,N_6945);
nor U8330 (N_8330,N_6095,N_6024);
nor U8331 (N_8331,N_6149,N_6516);
nand U8332 (N_8332,N_6775,N_6574);
or U8333 (N_8333,N_7283,N_6745);
xnor U8334 (N_8334,N_7315,N_6817);
or U8335 (N_8335,N_7475,N_7154);
or U8336 (N_8336,N_7320,N_6610);
and U8337 (N_8337,N_6206,N_6959);
and U8338 (N_8338,N_7278,N_6714);
or U8339 (N_8339,N_7019,N_7142);
nor U8340 (N_8340,N_7326,N_7351);
and U8341 (N_8341,N_7345,N_7399);
or U8342 (N_8342,N_7226,N_6500);
and U8343 (N_8343,N_6696,N_6687);
or U8344 (N_8344,N_6725,N_6206);
nand U8345 (N_8345,N_6893,N_6110);
nand U8346 (N_8346,N_6500,N_6130);
nor U8347 (N_8347,N_7455,N_6763);
nand U8348 (N_8348,N_7450,N_7359);
nand U8349 (N_8349,N_6052,N_7042);
nor U8350 (N_8350,N_6061,N_6721);
nor U8351 (N_8351,N_6347,N_6147);
or U8352 (N_8352,N_6180,N_6336);
nand U8353 (N_8353,N_7136,N_6261);
or U8354 (N_8354,N_7009,N_6378);
nor U8355 (N_8355,N_7467,N_7449);
nor U8356 (N_8356,N_7312,N_6464);
nand U8357 (N_8357,N_6508,N_7416);
and U8358 (N_8358,N_7344,N_6699);
nor U8359 (N_8359,N_6726,N_6076);
and U8360 (N_8360,N_6980,N_6222);
or U8361 (N_8361,N_6026,N_7192);
nand U8362 (N_8362,N_6177,N_7318);
or U8363 (N_8363,N_7348,N_6180);
and U8364 (N_8364,N_7113,N_6889);
xor U8365 (N_8365,N_7017,N_6680);
nand U8366 (N_8366,N_6258,N_6852);
nor U8367 (N_8367,N_6319,N_7362);
and U8368 (N_8368,N_6256,N_6886);
and U8369 (N_8369,N_6304,N_6256);
nor U8370 (N_8370,N_6792,N_6102);
nand U8371 (N_8371,N_7395,N_6439);
xor U8372 (N_8372,N_6032,N_7316);
nor U8373 (N_8373,N_7225,N_7009);
and U8374 (N_8374,N_7051,N_6421);
nand U8375 (N_8375,N_7172,N_6216);
nand U8376 (N_8376,N_7251,N_7306);
or U8377 (N_8377,N_7228,N_6096);
nand U8378 (N_8378,N_7091,N_7245);
nor U8379 (N_8379,N_6995,N_6910);
and U8380 (N_8380,N_6000,N_6050);
nand U8381 (N_8381,N_6093,N_6782);
or U8382 (N_8382,N_6107,N_7119);
nor U8383 (N_8383,N_6039,N_6254);
and U8384 (N_8384,N_6559,N_6835);
or U8385 (N_8385,N_6945,N_7417);
and U8386 (N_8386,N_7389,N_6304);
and U8387 (N_8387,N_7185,N_7327);
or U8388 (N_8388,N_7160,N_6447);
and U8389 (N_8389,N_7111,N_6131);
nand U8390 (N_8390,N_6820,N_6381);
or U8391 (N_8391,N_7060,N_7033);
nor U8392 (N_8392,N_6887,N_6116);
or U8393 (N_8393,N_6238,N_6245);
or U8394 (N_8394,N_6133,N_6776);
and U8395 (N_8395,N_6802,N_6870);
or U8396 (N_8396,N_6361,N_6748);
nor U8397 (N_8397,N_7034,N_6164);
and U8398 (N_8398,N_6456,N_6175);
and U8399 (N_8399,N_7499,N_7439);
or U8400 (N_8400,N_7069,N_7408);
nand U8401 (N_8401,N_7368,N_7172);
xor U8402 (N_8402,N_7360,N_6442);
or U8403 (N_8403,N_6748,N_6933);
and U8404 (N_8404,N_6746,N_6149);
nand U8405 (N_8405,N_6717,N_6570);
nand U8406 (N_8406,N_6329,N_6557);
nor U8407 (N_8407,N_7032,N_6438);
or U8408 (N_8408,N_6380,N_7145);
xnor U8409 (N_8409,N_7080,N_7467);
or U8410 (N_8410,N_7199,N_6939);
and U8411 (N_8411,N_7130,N_7388);
or U8412 (N_8412,N_7126,N_7401);
nand U8413 (N_8413,N_7208,N_6949);
nand U8414 (N_8414,N_6554,N_7440);
and U8415 (N_8415,N_6183,N_6608);
nor U8416 (N_8416,N_6463,N_7353);
nand U8417 (N_8417,N_6664,N_6442);
nor U8418 (N_8418,N_6733,N_7359);
and U8419 (N_8419,N_6237,N_7216);
xnor U8420 (N_8420,N_6140,N_6809);
and U8421 (N_8421,N_6010,N_6546);
or U8422 (N_8422,N_7069,N_6088);
nor U8423 (N_8423,N_6180,N_6935);
nand U8424 (N_8424,N_6978,N_6550);
nand U8425 (N_8425,N_7454,N_7092);
nor U8426 (N_8426,N_6144,N_6719);
xnor U8427 (N_8427,N_6277,N_6031);
or U8428 (N_8428,N_6659,N_6866);
nand U8429 (N_8429,N_7086,N_7148);
or U8430 (N_8430,N_6784,N_7498);
xnor U8431 (N_8431,N_6778,N_6408);
nand U8432 (N_8432,N_7172,N_6791);
and U8433 (N_8433,N_6590,N_7376);
nand U8434 (N_8434,N_7211,N_7410);
and U8435 (N_8435,N_7099,N_7304);
nor U8436 (N_8436,N_6043,N_7052);
or U8437 (N_8437,N_7334,N_6820);
or U8438 (N_8438,N_7016,N_7481);
nor U8439 (N_8439,N_7311,N_7333);
nor U8440 (N_8440,N_6470,N_7398);
and U8441 (N_8441,N_6856,N_6863);
or U8442 (N_8442,N_7412,N_7323);
or U8443 (N_8443,N_7184,N_6682);
or U8444 (N_8444,N_7211,N_6093);
and U8445 (N_8445,N_7411,N_6795);
nand U8446 (N_8446,N_6997,N_7466);
or U8447 (N_8447,N_6887,N_6439);
and U8448 (N_8448,N_7310,N_7303);
nor U8449 (N_8449,N_7425,N_7101);
nor U8450 (N_8450,N_7189,N_6214);
and U8451 (N_8451,N_6415,N_7307);
nor U8452 (N_8452,N_6730,N_7155);
or U8453 (N_8453,N_6885,N_6183);
nand U8454 (N_8454,N_6198,N_7272);
or U8455 (N_8455,N_6801,N_6099);
and U8456 (N_8456,N_7477,N_6957);
xor U8457 (N_8457,N_7200,N_6545);
or U8458 (N_8458,N_7099,N_6085);
nand U8459 (N_8459,N_6046,N_7485);
or U8460 (N_8460,N_6477,N_6315);
nor U8461 (N_8461,N_6393,N_6955);
nor U8462 (N_8462,N_6725,N_7245);
nor U8463 (N_8463,N_7280,N_6814);
and U8464 (N_8464,N_7279,N_7145);
nand U8465 (N_8465,N_6097,N_7007);
or U8466 (N_8466,N_7452,N_7188);
or U8467 (N_8467,N_7424,N_6090);
or U8468 (N_8468,N_7317,N_6742);
or U8469 (N_8469,N_7054,N_6985);
and U8470 (N_8470,N_7082,N_7348);
nor U8471 (N_8471,N_6502,N_6556);
nand U8472 (N_8472,N_6624,N_6141);
nand U8473 (N_8473,N_6176,N_6907);
or U8474 (N_8474,N_6846,N_7137);
and U8475 (N_8475,N_6905,N_7323);
nand U8476 (N_8476,N_7482,N_6271);
and U8477 (N_8477,N_6391,N_6390);
and U8478 (N_8478,N_7375,N_6728);
xnor U8479 (N_8479,N_6149,N_6447);
nand U8480 (N_8480,N_6863,N_6638);
nand U8481 (N_8481,N_7210,N_7215);
nor U8482 (N_8482,N_6240,N_6444);
nor U8483 (N_8483,N_6086,N_7032);
or U8484 (N_8484,N_7001,N_6390);
or U8485 (N_8485,N_6689,N_6649);
nor U8486 (N_8486,N_6239,N_6549);
xor U8487 (N_8487,N_7460,N_7042);
or U8488 (N_8488,N_7438,N_6165);
nor U8489 (N_8489,N_6206,N_7258);
nor U8490 (N_8490,N_7335,N_7201);
or U8491 (N_8491,N_6030,N_6534);
nor U8492 (N_8492,N_6410,N_6609);
nand U8493 (N_8493,N_6276,N_7237);
or U8494 (N_8494,N_6410,N_6634);
and U8495 (N_8495,N_6782,N_6356);
and U8496 (N_8496,N_6537,N_7216);
and U8497 (N_8497,N_6559,N_6796);
nand U8498 (N_8498,N_6933,N_6605);
or U8499 (N_8499,N_7048,N_7107);
nand U8500 (N_8500,N_6956,N_6032);
or U8501 (N_8501,N_6413,N_6147);
nor U8502 (N_8502,N_7282,N_6377);
or U8503 (N_8503,N_6933,N_7451);
and U8504 (N_8504,N_6807,N_7286);
or U8505 (N_8505,N_6410,N_7448);
nand U8506 (N_8506,N_6108,N_7089);
or U8507 (N_8507,N_6078,N_7261);
and U8508 (N_8508,N_6095,N_7177);
nand U8509 (N_8509,N_7082,N_6077);
nor U8510 (N_8510,N_6830,N_6591);
xor U8511 (N_8511,N_6050,N_7089);
nor U8512 (N_8512,N_7393,N_7416);
and U8513 (N_8513,N_6381,N_6866);
and U8514 (N_8514,N_6701,N_6560);
nor U8515 (N_8515,N_7267,N_7292);
or U8516 (N_8516,N_6201,N_6794);
nor U8517 (N_8517,N_6669,N_7136);
nor U8518 (N_8518,N_6856,N_6755);
or U8519 (N_8519,N_6585,N_6501);
nand U8520 (N_8520,N_6438,N_7378);
and U8521 (N_8521,N_6936,N_7457);
or U8522 (N_8522,N_6280,N_6754);
nand U8523 (N_8523,N_6899,N_6329);
or U8524 (N_8524,N_6682,N_6137);
nor U8525 (N_8525,N_6538,N_6133);
nor U8526 (N_8526,N_7192,N_6578);
nand U8527 (N_8527,N_6093,N_7462);
and U8528 (N_8528,N_6380,N_6543);
or U8529 (N_8529,N_6953,N_6962);
xor U8530 (N_8530,N_7189,N_6085);
xor U8531 (N_8531,N_6597,N_6701);
nand U8532 (N_8532,N_6421,N_7158);
or U8533 (N_8533,N_6754,N_7254);
nand U8534 (N_8534,N_6934,N_6196);
or U8535 (N_8535,N_6569,N_6292);
nand U8536 (N_8536,N_7164,N_6133);
nand U8537 (N_8537,N_6971,N_7343);
and U8538 (N_8538,N_6878,N_6883);
nor U8539 (N_8539,N_7001,N_7340);
nor U8540 (N_8540,N_7150,N_7049);
or U8541 (N_8541,N_6814,N_6326);
nor U8542 (N_8542,N_6126,N_6711);
nand U8543 (N_8543,N_7308,N_6632);
nor U8544 (N_8544,N_6124,N_7396);
nor U8545 (N_8545,N_7230,N_7031);
nand U8546 (N_8546,N_6330,N_6660);
nor U8547 (N_8547,N_7395,N_6890);
xnor U8548 (N_8548,N_6100,N_6771);
and U8549 (N_8549,N_6278,N_6760);
xor U8550 (N_8550,N_6881,N_6083);
or U8551 (N_8551,N_6098,N_6601);
or U8552 (N_8552,N_7338,N_6484);
and U8553 (N_8553,N_6321,N_6426);
nand U8554 (N_8554,N_6387,N_6731);
nor U8555 (N_8555,N_7479,N_6399);
nor U8556 (N_8556,N_6431,N_7481);
nand U8557 (N_8557,N_6286,N_7186);
nand U8558 (N_8558,N_7429,N_7044);
or U8559 (N_8559,N_7241,N_7465);
and U8560 (N_8560,N_6608,N_6976);
nand U8561 (N_8561,N_6405,N_7247);
xnor U8562 (N_8562,N_7498,N_7238);
nor U8563 (N_8563,N_6272,N_6620);
nand U8564 (N_8564,N_7305,N_6120);
nor U8565 (N_8565,N_6304,N_6625);
or U8566 (N_8566,N_6837,N_6958);
nor U8567 (N_8567,N_6886,N_7407);
nand U8568 (N_8568,N_6330,N_6112);
nor U8569 (N_8569,N_6414,N_7436);
nand U8570 (N_8570,N_6607,N_7209);
nand U8571 (N_8571,N_6403,N_6223);
nand U8572 (N_8572,N_6552,N_6183);
nor U8573 (N_8573,N_6074,N_6420);
and U8574 (N_8574,N_6200,N_7321);
and U8575 (N_8575,N_6069,N_6021);
or U8576 (N_8576,N_6667,N_6486);
and U8577 (N_8577,N_7009,N_7345);
nor U8578 (N_8578,N_7202,N_7371);
xnor U8579 (N_8579,N_7172,N_6059);
nand U8580 (N_8580,N_6003,N_6945);
nor U8581 (N_8581,N_7177,N_7146);
or U8582 (N_8582,N_6793,N_6026);
or U8583 (N_8583,N_7473,N_6962);
and U8584 (N_8584,N_7308,N_7079);
and U8585 (N_8585,N_6070,N_7376);
and U8586 (N_8586,N_7364,N_7030);
nand U8587 (N_8587,N_6307,N_6709);
or U8588 (N_8588,N_6515,N_6526);
or U8589 (N_8589,N_6098,N_6725);
and U8590 (N_8590,N_6219,N_6757);
and U8591 (N_8591,N_7169,N_6636);
nor U8592 (N_8592,N_6297,N_7258);
and U8593 (N_8593,N_7006,N_7025);
and U8594 (N_8594,N_6833,N_7295);
and U8595 (N_8595,N_7128,N_6240);
nand U8596 (N_8596,N_7256,N_7341);
and U8597 (N_8597,N_6864,N_6297);
and U8598 (N_8598,N_6872,N_6603);
nor U8599 (N_8599,N_6105,N_6900);
and U8600 (N_8600,N_7075,N_7495);
nor U8601 (N_8601,N_7008,N_6802);
xor U8602 (N_8602,N_7055,N_6513);
nor U8603 (N_8603,N_6780,N_7445);
and U8604 (N_8604,N_6394,N_6960);
nor U8605 (N_8605,N_7212,N_6484);
nand U8606 (N_8606,N_6575,N_6405);
or U8607 (N_8607,N_6866,N_7124);
or U8608 (N_8608,N_6512,N_6500);
nor U8609 (N_8609,N_6866,N_6967);
and U8610 (N_8610,N_6334,N_7192);
or U8611 (N_8611,N_6518,N_7023);
nand U8612 (N_8612,N_7059,N_7144);
or U8613 (N_8613,N_6895,N_7026);
nand U8614 (N_8614,N_6362,N_6896);
and U8615 (N_8615,N_6528,N_6803);
xor U8616 (N_8616,N_6752,N_6071);
xnor U8617 (N_8617,N_6306,N_6677);
nand U8618 (N_8618,N_6220,N_6686);
nand U8619 (N_8619,N_6501,N_7371);
nor U8620 (N_8620,N_6925,N_7035);
or U8621 (N_8621,N_6286,N_7107);
xor U8622 (N_8622,N_6228,N_6638);
or U8623 (N_8623,N_6773,N_6147);
and U8624 (N_8624,N_6835,N_6907);
and U8625 (N_8625,N_6554,N_7445);
nand U8626 (N_8626,N_6511,N_6620);
or U8627 (N_8627,N_6189,N_6008);
nand U8628 (N_8628,N_6962,N_7223);
nand U8629 (N_8629,N_6431,N_6245);
nand U8630 (N_8630,N_6199,N_6069);
and U8631 (N_8631,N_7335,N_6093);
nor U8632 (N_8632,N_7491,N_6111);
and U8633 (N_8633,N_6125,N_7483);
nor U8634 (N_8634,N_7301,N_7349);
nand U8635 (N_8635,N_7187,N_6264);
nand U8636 (N_8636,N_6216,N_7442);
and U8637 (N_8637,N_6458,N_6466);
or U8638 (N_8638,N_7126,N_6590);
and U8639 (N_8639,N_7451,N_6337);
xor U8640 (N_8640,N_7496,N_7123);
or U8641 (N_8641,N_7344,N_6195);
and U8642 (N_8642,N_7074,N_6018);
nand U8643 (N_8643,N_7207,N_7022);
nand U8644 (N_8644,N_6502,N_7098);
xor U8645 (N_8645,N_6019,N_7091);
and U8646 (N_8646,N_6020,N_6758);
or U8647 (N_8647,N_6208,N_6903);
nor U8648 (N_8648,N_6369,N_7351);
and U8649 (N_8649,N_6063,N_6537);
xor U8650 (N_8650,N_7166,N_6926);
and U8651 (N_8651,N_7145,N_6260);
nand U8652 (N_8652,N_7347,N_7413);
nor U8653 (N_8653,N_6989,N_6045);
nor U8654 (N_8654,N_6315,N_7176);
nor U8655 (N_8655,N_6958,N_6790);
nor U8656 (N_8656,N_6712,N_6554);
and U8657 (N_8657,N_7254,N_7469);
and U8658 (N_8658,N_6242,N_6700);
nand U8659 (N_8659,N_7178,N_6318);
or U8660 (N_8660,N_6494,N_7341);
and U8661 (N_8661,N_6160,N_7385);
and U8662 (N_8662,N_7309,N_6180);
or U8663 (N_8663,N_7240,N_7178);
nor U8664 (N_8664,N_6412,N_6687);
or U8665 (N_8665,N_6629,N_6224);
or U8666 (N_8666,N_7166,N_7300);
or U8667 (N_8667,N_6599,N_7063);
xor U8668 (N_8668,N_7376,N_6815);
xnor U8669 (N_8669,N_6350,N_6351);
and U8670 (N_8670,N_6691,N_6507);
and U8671 (N_8671,N_6215,N_7446);
nor U8672 (N_8672,N_6454,N_6830);
and U8673 (N_8673,N_6905,N_7058);
or U8674 (N_8674,N_7245,N_6750);
nor U8675 (N_8675,N_6782,N_6941);
or U8676 (N_8676,N_7155,N_6954);
nor U8677 (N_8677,N_6209,N_6237);
and U8678 (N_8678,N_6879,N_7428);
xor U8679 (N_8679,N_7175,N_7377);
and U8680 (N_8680,N_6664,N_6412);
and U8681 (N_8681,N_7007,N_6883);
nor U8682 (N_8682,N_6825,N_7473);
and U8683 (N_8683,N_6002,N_6157);
or U8684 (N_8684,N_6797,N_6589);
and U8685 (N_8685,N_6739,N_6039);
nor U8686 (N_8686,N_6715,N_6207);
and U8687 (N_8687,N_6202,N_6755);
or U8688 (N_8688,N_6093,N_6190);
nor U8689 (N_8689,N_6369,N_7059);
nand U8690 (N_8690,N_7005,N_7031);
or U8691 (N_8691,N_7485,N_6880);
nand U8692 (N_8692,N_7302,N_7187);
and U8693 (N_8693,N_7034,N_6034);
nor U8694 (N_8694,N_6337,N_6718);
or U8695 (N_8695,N_7046,N_6388);
nor U8696 (N_8696,N_6607,N_7498);
or U8697 (N_8697,N_6891,N_6892);
and U8698 (N_8698,N_6717,N_7039);
nand U8699 (N_8699,N_6830,N_7115);
or U8700 (N_8700,N_6826,N_6533);
xnor U8701 (N_8701,N_6118,N_6545);
or U8702 (N_8702,N_6997,N_6254);
xor U8703 (N_8703,N_6730,N_6902);
or U8704 (N_8704,N_6441,N_7454);
and U8705 (N_8705,N_7431,N_6091);
nand U8706 (N_8706,N_6921,N_6962);
nand U8707 (N_8707,N_6015,N_6278);
nor U8708 (N_8708,N_6704,N_6047);
and U8709 (N_8709,N_7260,N_6615);
or U8710 (N_8710,N_7100,N_6236);
and U8711 (N_8711,N_6813,N_6900);
xnor U8712 (N_8712,N_6759,N_7112);
or U8713 (N_8713,N_7178,N_6165);
and U8714 (N_8714,N_7436,N_6710);
or U8715 (N_8715,N_6237,N_6387);
nand U8716 (N_8716,N_6871,N_7386);
or U8717 (N_8717,N_7454,N_7498);
nand U8718 (N_8718,N_6805,N_6494);
nor U8719 (N_8719,N_7141,N_6708);
nand U8720 (N_8720,N_6746,N_6953);
or U8721 (N_8721,N_7038,N_6347);
xor U8722 (N_8722,N_7222,N_7165);
and U8723 (N_8723,N_6123,N_6906);
xor U8724 (N_8724,N_6319,N_6942);
nor U8725 (N_8725,N_6154,N_6763);
and U8726 (N_8726,N_6221,N_7095);
and U8727 (N_8727,N_7295,N_6763);
xor U8728 (N_8728,N_6148,N_6906);
or U8729 (N_8729,N_7312,N_6097);
or U8730 (N_8730,N_6152,N_6518);
and U8731 (N_8731,N_6301,N_6907);
or U8732 (N_8732,N_6956,N_7126);
nand U8733 (N_8733,N_6477,N_6404);
and U8734 (N_8734,N_6365,N_6247);
and U8735 (N_8735,N_6765,N_7027);
or U8736 (N_8736,N_6116,N_7228);
nor U8737 (N_8737,N_7469,N_7498);
nor U8738 (N_8738,N_6324,N_6578);
nor U8739 (N_8739,N_6868,N_6165);
xor U8740 (N_8740,N_7393,N_6814);
or U8741 (N_8741,N_6462,N_6793);
and U8742 (N_8742,N_6131,N_7471);
or U8743 (N_8743,N_7314,N_6749);
nor U8744 (N_8744,N_6569,N_6813);
or U8745 (N_8745,N_7369,N_6995);
or U8746 (N_8746,N_7164,N_6918);
nand U8747 (N_8747,N_6079,N_7454);
or U8748 (N_8748,N_7148,N_7135);
nor U8749 (N_8749,N_6265,N_7264);
or U8750 (N_8750,N_7230,N_7144);
nor U8751 (N_8751,N_6241,N_6282);
and U8752 (N_8752,N_6880,N_6603);
and U8753 (N_8753,N_6421,N_6327);
xor U8754 (N_8754,N_6534,N_7254);
xor U8755 (N_8755,N_6810,N_7303);
and U8756 (N_8756,N_7498,N_7406);
or U8757 (N_8757,N_6913,N_7412);
xor U8758 (N_8758,N_6383,N_7330);
or U8759 (N_8759,N_6655,N_7028);
nand U8760 (N_8760,N_7358,N_6855);
or U8761 (N_8761,N_6009,N_7196);
nand U8762 (N_8762,N_6751,N_6705);
nand U8763 (N_8763,N_6414,N_6920);
nand U8764 (N_8764,N_7241,N_6830);
nand U8765 (N_8765,N_6294,N_6074);
nor U8766 (N_8766,N_7351,N_6909);
xor U8767 (N_8767,N_6854,N_6551);
nor U8768 (N_8768,N_6086,N_7303);
and U8769 (N_8769,N_6544,N_7205);
nor U8770 (N_8770,N_6001,N_6768);
xor U8771 (N_8771,N_6219,N_6424);
nand U8772 (N_8772,N_7280,N_6147);
or U8773 (N_8773,N_6971,N_6319);
and U8774 (N_8774,N_7178,N_7270);
and U8775 (N_8775,N_7477,N_7342);
and U8776 (N_8776,N_6608,N_6953);
or U8777 (N_8777,N_6826,N_6539);
or U8778 (N_8778,N_6142,N_6851);
xnor U8779 (N_8779,N_6353,N_6576);
nand U8780 (N_8780,N_7185,N_6217);
and U8781 (N_8781,N_6169,N_7213);
and U8782 (N_8782,N_6790,N_7396);
and U8783 (N_8783,N_6312,N_6581);
nor U8784 (N_8784,N_6052,N_7069);
or U8785 (N_8785,N_6180,N_6296);
nand U8786 (N_8786,N_6453,N_6393);
nand U8787 (N_8787,N_6681,N_6646);
nor U8788 (N_8788,N_6545,N_6816);
and U8789 (N_8789,N_6233,N_6219);
nor U8790 (N_8790,N_6618,N_7410);
and U8791 (N_8791,N_6223,N_7229);
or U8792 (N_8792,N_6942,N_6126);
and U8793 (N_8793,N_7030,N_6595);
nand U8794 (N_8794,N_6441,N_6811);
or U8795 (N_8795,N_6594,N_6814);
nor U8796 (N_8796,N_6591,N_6405);
nor U8797 (N_8797,N_7060,N_6914);
nor U8798 (N_8798,N_6506,N_7085);
nor U8799 (N_8799,N_7301,N_6885);
xnor U8800 (N_8800,N_6768,N_6721);
and U8801 (N_8801,N_6774,N_6595);
nand U8802 (N_8802,N_7365,N_6665);
nand U8803 (N_8803,N_6714,N_6758);
and U8804 (N_8804,N_6076,N_6826);
nand U8805 (N_8805,N_7249,N_6774);
and U8806 (N_8806,N_6737,N_7182);
and U8807 (N_8807,N_6375,N_6782);
nand U8808 (N_8808,N_7448,N_7291);
nand U8809 (N_8809,N_6554,N_7474);
nand U8810 (N_8810,N_6949,N_7239);
and U8811 (N_8811,N_6471,N_6782);
nor U8812 (N_8812,N_7392,N_6596);
nand U8813 (N_8813,N_6222,N_6324);
nand U8814 (N_8814,N_7005,N_7486);
xor U8815 (N_8815,N_6198,N_6210);
xnor U8816 (N_8816,N_6885,N_7013);
nor U8817 (N_8817,N_6194,N_6325);
nor U8818 (N_8818,N_6004,N_6187);
nand U8819 (N_8819,N_6104,N_6870);
nor U8820 (N_8820,N_7154,N_6694);
nor U8821 (N_8821,N_6978,N_6255);
xor U8822 (N_8822,N_6002,N_6756);
nor U8823 (N_8823,N_6741,N_7110);
or U8824 (N_8824,N_7000,N_6218);
xnor U8825 (N_8825,N_6567,N_6939);
nor U8826 (N_8826,N_7456,N_7211);
or U8827 (N_8827,N_6148,N_6234);
nor U8828 (N_8828,N_6389,N_6543);
nand U8829 (N_8829,N_6648,N_6033);
or U8830 (N_8830,N_6546,N_6875);
and U8831 (N_8831,N_6475,N_6919);
nor U8832 (N_8832,N_6026,N_6081);
nand U8833 (N_8833,N_6072,N_7381);
nor U8834 (N_8834,N_6997,N_6580);
and U8835 (N_8835,N_7238,N_6692);
nand U8836 (N_8836,N_6646,N_6359);
or U8837 (N_8837,N_6097,N_6325);
or U8838 (N_8838,N_6855,N_6858);
nand U8839 (N_8839,N_7413,N_6774);
xor U8840 (N_8840,N_6779,N_6913);
or U8841 (N_8841,N_6461,N_6754);
nand U8842 (N_8842,N_7272,N_6103);
nor U8843 (N_8843,N_6076,N_6230);
xor U8844 (N_8844,N_6711,N_6637);
and U8845 (N_8845,N_7435,N_6312);
or U8846 (N_8846,N_6464,N_6577);
or U8847 (N_8847,N_7017,N_7263);
and U8848 (N_8848,N_7376,N_6569);
nand U8849 (N_8849,N_6862,N_7226);
nand U8850 (N_8850,N_6354,N_6337);
or U8851 (N_8851,N_6253,N_7419);
or U8852 (N_8852,N_6541,N_7404);
xor U8853 (N_8853,N_6198,N_7238);
nor U8854 (N_8854,N_6791,N_6844);
or U8855 (N_8855,N_7140,N_7190);
xnor U8856 (N_8856,N_6284,N_6050);
nor U8857 (N_8857,N_6182,N_6055);
or U8858 (N_8858,N_6277,N_7121);
xor U8859 (N_8859,N_6003,N_6753);
nand U8860 (N_8860,N_7450,N_7092);
and U8861 (N_8861,N_7000,N_6585);
nor U8862 (N_8862,N_6172,N_6013);
nand U8863 (N_8863,N_6046,N_7147);
xnor U8864 (N_8864,N_7111,N_7498);
and U8865 (N_8865,N_6189,N_6154);
nor U8866 (N_8866,N_7025,N_6638);
nand U8867 (N_8867,N_7389,N_7443);
nor U8868 (N_8868,N_6719,N_6060);
and U8869 (N_8869,N_7211,N_6530);
nor U8870 (N_8870,N_7070,N_7242);
and U8871 (N_8871,N_6777,N_7227);
or U8872 (N_8872,N_6249,N_6149);
or U8873 (N_8873,N_6954,N_6585);
or U8874 (N_8874,N_6742,N_7487);
nand U8875 (N_8875,N_6360,N_6645);
nand U8876 (N_8876,N_6962,N_6654);
nor U8877 (N_8877,N_7497,N_7262);
nor U8878 (N_8878,N_7025,N_6155);
nor U8879 (N_8879,N_7246,N_7165);
or U8880 (N_8880,N_7249,N_6823);
or U8881 (N_8881,N_6901,N_7239);
or U8882 (N_8882,N_6644,N_7288);
nand U8883 (N_8883,N_6078,N_6014);
and U8884 (N_8884,N_6309,N_7464);
nand U8885 (N_8885,N_6819,N_6710);
and U8886 (N_8886,N_7079,N_7001);
or U8887 (N_8887,N_6471,N_6381);
and U8888 (N_8888,N_6956,N_6170);
or U8889 (N_8889,N_6652,N_7414);
or U8890 (N_8890,N_6954,N_7350);
nand U8891 (N_8891,N_6838,N_7422);
xor U8892 (N_8892,N_6817,N_6917);
xnor U8893 (N_8893,N_6544,N_6438);
or U8894 (N_8894,N_7264,N_7445);
or U8895 (N_8895,N_6370,N_6233);
nor U8896 (N_8896,N_6247,N_7065);
and U8897 (N_8897,N_6856,N_6274);
nand U8898 (N_8898,N_7096,N_7415);
nand U8899 (N_8899,N_6823,N_7074);
and U8900 (N_8900,N_7108,N_6945);
nand U8901 (N_8901,N_6574,N_7079);
nand U8902 (N_8902,N_7133,N_6548);
and U8903 (N_8903,N_6748,N_6378);
or U8904 (N_8904,N_7459,N_6068);
or U8905 (N_8905,N_6371,N_6687);
or U8906 (N_8906,N_6297,N_6880);
or U8907 (N_8907,N_6666,N_7102);
nand U8908 (N_8908,N_7109,N_7006);
nand U8909 (N_8909,N_6081,N_7498);
nor U8910 (N_8910,N_6450,N_7370);
nor U8911 (N_8911,N_6647,N_6912);
nor U8912 (N_8912,N_6806,N_7458);
nor U8913 (N_8913,N_6541,N_7345);
xnor U8914 (N_8914,N_6926,N_7114);
and U8915 (N_8915,N_7110,N_6841);
nand U8916 (N_8916,N_6282,N_7374);
and U8917 (N_8917,N_6193,N_7079);
or U8918 (N_8918,N_7120,N_6084);
nand U8919 (N_8919,N_7249,N_6737);
nand U8920 (N_8920,N_6770,N_7392);
and U8921 (N_8921,N_6914,N_7004);
nor U8922 (N_8922,N_6014,N_6603);
or U8923 (N_8923,N_7160,N_6699);
nand U8924 (N_8924,N_6941,N_6612);
and U8925 (N_8925,N_6246,N_7356);
nor U8926 (N_8926,N_6613,N_6748);
nor U8927 (N_8927,N_6946,N_6642);
nand U8928 (N_8928,N_6471,N_6892);
nor U8929 (N_8929,N_6322,N_6332);
nand U8930 (N_8930,N_6498,N_7251);
nor U8931 (N_8931,N_7179,N_7431);
and U8932 (N_8932,N_6740,N_6152);
or U8933 (N_8933,N_6333,N_7476);
nor U8934 (N_8934,N_6889,N_7039);
nor U8935 (N_8935,N_6079,N_6173);
or U8936 (N_8936,N_7208,N_6944);
nand U8937 (N_8937,N_6477,N_6191);
and U8938 (N_8938,N_6048,N_6432);
and U8939 (N_8939,N_7222,N_6639);
xnor U8940 (N_8940,N_7356,N_6407);
or U8941 (N_8941,N_6577,N_6396);
nor U8942 (N_8942,N_6994,N_7079);
nor U8943 (N_8943,N_6534,N_7004);
nor U8944 (N_8944,N_6478,N_6520);
nand U8945 (N_8945,N_7079,N_7432);
or U8946 (N_8946,N_6716,N_7232);
or U8947 (N_8947,N_6690,N_6290);
and U8948 (N_8948,N_6707,N_6956);
and U8949 (N_8949,N_7258,N_7415);
or U8950 (N_8950,N_7344,N_7290);
or U8951 (N_8951,N_7055,N_7108);
or U8952 (N_8952,N_6680,N_6894);
or U8953 (N_8953,N_7308,N_6095);
nand U8954 (N_8954,N_6946,N_7283);
nand U8955 (N_8955,N_6657,N_7160);
nor U8956 (N_8956,N_6403,N_6898);
and U8957 (N_8957,N_7126,N_6024);
nand U8958 (N_8958,N_6983,N_6008);
and U8959 (N_8959,N_7358,N_6400);
nand U8960 (N_8960,N_6873,N_6719);
nor U8961 (N_8961,N_7268,N_6343);
and U8962 (N_8962,N_6956,N_6330);
nor U8963 (N_8963,N_7311,N_7013);
nor U8964 (N_8964,N_6583,N_6905);
and U8965 (N_8965,N_6926,N_6588);
or U8966 (N_8966,N_7279,N_7328);
or U8967 (N_8967,N_6962,N_6252);
nor U8968 (N_8968,N_6210,N_7061);
nor U8969 (N_8969,N_6838,N_7149);
nor U8970 (N_8970,N_7335,N_7169);
xor U8971 (N_8971,N_6854,N_6567);
nand U8972 (N_8972,N_7097,N_6927);
nor U8973 (N_8973,N_6382,N_6094);
and U8974 (N_8974,N_7043,N_6697);
nor U8975 (N_8975,N_6119,N_6683);
or U8976 (N_8976,N_6514,N_6323);
nand U8977 (N_8977,N_7408,N_7399);
nor U8978 (N_8978,N_6317,N_6340);
or U8979 (N_8979,N_6979,N_6610);
and U8980 (N_8980,N_7478,N_6551);
xnor U8981 (N_8981,N_6340,N_6087);
nor U8982 (N_8982,N_7397,N_6976);
or U8983 (N_8983,N_6221,N_7410);
and U8984 (N_8984,N_6426,N_7308);
or U8985 (N_8985,N_6601,N_6683);
or U8986 (N_8986,N_6133,N_7046);
and U8987 (N_8987,N_7339,N_6762);
xnor U8988 (N_8988,N_6546,N_7261);
nor U8989 (N_8989,N_7021,N_7257);
or U8990 (N_8990,N_6634,N_7223);
nand U8991 (N_8991,N_6184,N_6304);
xor U8992 (N_8992,N_6516,N_6829);
or U8993 (N_8993,N_7115,N_7433);
nand U8994 (N_8994,N_6826,N_7031);
or U8995 (N_8995,N_7478,N_6320);
or U8996 (N_8996,N_6524,N_6663);
nand U8997 (N_8997,N_6584,N_7312);
nand U8998 (N_8998,N_6371,N_7367);
xor U8999 (N_8999,N_7471,N_6556);
or U9000 (N_9000,N_8892,N_8985);
and U9001 (N_9001,N_8915,N_7982);
and U9002 (N_9002,N_8431,N_7636);
nor U9003 (N_9003,N_8815,N_8636);
and U9004 (N_9004,N_7954,N_8576);
and U9005 (N_9005,N_8963,N_8343);
xnor U9006 (N_9006,N_8353,N_7588);
nor U9007 (N_9007,N_8301,N_8617);
xnor U9008 (N_9008,N_7738,N_8467);
xnor U9009 (N_9009,N_7745,N_7553);
and U9010 (N_9010,N_8344,N_8639);
nand U9011 (N_9011,N_8604,N_8479);
and U9012 (N_9012,N_8950,N_8690);
nand U9013 (N_9013,N_7810,N_8633);
xnor U9014 (N_9014,N_7609,N_8172);
xnor U9015 (N_9015,N_7619,N_7763);
or U9016 (N_9016,N_7956,N_8265);
or U9017 (N_9017,N_8833,N_8644);
nor U9018 (N_9018,N_8623,N_8119);
nor U9019 (N_9019,N_7526,N_8981);
or U9020 (N_9020,N_8387,N_8895);
nand U9021 (N_9021,N_7963,N_7626);
xor U9022 (N_9022,N_8808,N_8851);
xnor U9023 (N_9023,N_7688,N_7727);
nand U9024 (N_9024,N_8540,N_8563);
and U9025 (N_9025,N_8316,N_8331);
nand U9026 (N_9026,N_8884,N_7864);
nor U9027 (N_9027,N_8830,N_8294);
xor U9028 (N_9028,N_8889,N_7530);
xor U9029 (N_9029,N_7991,N_8156);
xnor U9030 (N_9030,N_7573,N_8772);
xor U9031 (N_9031,N_7603,N_8930);
nor U9032 (N_9032,N_8153,N_7884);
nor U9033 (N_9033,N_8429,N_7611);
or U9034 (N_9034,N_7517,N_7572);
nor U9035 (N_9035,N_8448,N_8613);
and U9036 (N_9036,N_7950,N_8986);
and U9037 (N_9037,N_7882,N_7726);
or U9038 (N_9038,N_8380,N_7842);
or U9039 (N_9039,N_8136,N_7943);
nor U9040 (N_9040,N_7989,N_8253);
nor U9041 (N_9041,N_8532,N_8512);
nor U9042 (N_9042,N_8840,N_8612);
nand U9043 (N_9043,N_8242,N_7541);
nand U9044 (N_9044,N_7642,N_8568);
nor U9045 (N_9045,N_8192,N_7955);
nand U9046 (N_9046,N_7962,N_8785);
nor U9047 (N_9047,N_8250,N_7586);
or U9048 (N_9048,N_7694,N_7761);
or U9049 (N_9049,N_8761,N_8687);
nor U9050 (N_9050,N_7787,N_7511);
nand U9051 (N_9051,N_7545,N_7781);
nand U9052 (N_9052,N_8960,N_8675);
and U9053 (N_9053,N_7925,N_7786);
nand U9054 (N_9054,N_7812,N_8480);
nor U9055 (N_9055,N_8686,N_7702);
and U9056 (N_9056,N_8984,N_8476);
nand U9057 (N_9057,N_8740,N_7585);
nor U9058 (N_9058,N_8013,N_8206);
or U9059 (N_9059,N_8920,N_8086);
or U9060 (N_9060,N_8152,N_8526);
xnor U9061 (N_9061,N_7622,N_8426);
or U9062 (N_9062,N_8261,N_8183);
nand U9063 (N_9063,N_8088,N_8566);
and U9064 (N_9064,N_8271,N_8262);
or U9065 (N_9065,N_7684,N_8135);
and U9066 (N_9066,N_8908,N_7987);
nand U9067 (N_9067,N_8050,N_8988);
xor U9068 (N_9068,N_8427,N_8520);
or U9069 (N_9069,N_8412,N_8861);
nand U9070 (N_9070,N_8436,N_7880);
and U9071 (N_9071,N_8787,N_8441);
or U9072 (N_9072,N_7900,N_8043);
nor U9073 (N_9073,N_8051,N_8514);
and U9074 (N_9074,N_7858,N_7504);
or U9075 (N_9075,N_8508,N_8545);
and U9076 (N_9076,N_8795,N_8462);
xor U9077 (N_9077,N_8975,N_7779);
nor U9078 (N_9078,N_7932,N_7914);
or U9079 (N_9079,N_8789,N_8974);
and U9080 (N_9080,N_8866,N_8989);
or U9081 (N_9081,N_8034,N_8862);
and U9082 (N_9082,N_7853,N_7693);
and U9083 (N_9083,N_8956,N_7951);
and U9084 (N_9084,N_8729,N_8001);
and U9085 (N_9085,N_7966,N_8674);
or U9086 (N_9086,N_8921,N_8300);
nand U9087 (N_9087,N_8899,N_8324);
or U9088 (N_9088,N_8969,N_8857);
nand U9089 (N_9089,N_8798,N_8147);
nor U9090 (N_9090,N_7968,N_8337);
nand U9091 (N_9091,N_8796,N_8475);
and U9092 (N_9092,N_8310,N_8291);
xnor U9093 (N_9093,N_7592,N_8414);
nand U9094 (N_9094,N_7658,N_7927);
and U9095 (N_9095,N_7898,N_7773);
xor U9096 (N_9096,N_8537,N_8037);
xor U9097 (N_9097,N_8099,N_8205);
or U9098 (N_9098,N_7793,N_7581);
nor U9099 (N_9099,N_8834,N_7699);
or U9100 (N_9100,N_8401,N_7621);
or U9101 (N_9101,N_8155,N_8621);
nand U9102 (N_9102,N_8564,N_7679);
nand U9103 (N_9103,N_8408,N_8492);
or U9104 (N_9104,N_8252,N_8138);
nand U9105 (N_9105,N_7698,N_8757);
xnor U9106 (N_9106,N_8870,N_7670);
or U9107 (N_9107,N_8330,N_7835);
nand U9108 (N_9108,N_8054,N_8713);
nor U9109 (N_9109,N_8111,N_8482);
nor U9110 (N_9110,N_8752,N_8045);
nor U9111 (N_9111,N_8284,N_8768);
nor U9112 (N_9112,N_7969,N_8784);
or U9113 (N_9113,N_8854,N_7705);
nand U9114 (N_9114,N_8075,N_8125);
nor U9115 (N_9115,N_8531,N_8407);
nor U9116 (N_9116,N_8214,N_8556);
and U9117 (N_9117,N_8031,N_8006);
nor U9118 (N_9118,N_7796,N_7507);
and U9119 (N_9119,N_7997,N_8485);
xor U9120 (N_9120,N_8342,N_7529);
or U9121 (N_9121,N_8444,N_8428);
nand U9122 (N_9122,N_8906,N_8179);
and U9123 (N_9123,N_7790,N_8249);
xor U9124 (N_9124,N_8945,N_8498);
xor U9125 (N_9125,N_7683,N_8158);
and U9126 (N_9126,N_8773,N_7938);
and U9127 (N_9127,N_7614,N_8823);
and U9128 (N_9128,N_8523,N_8501);
and U9129 (N_9129,N_8048,N_8680);
and U9130 (N_9130,N_8517,N_8145);
nor U9131 (N_9131,N_8762,N_7605);
or U9132 (N_9132,N_7990,N_8141);
nor U9133 (N_9133,N_7704,N_8968);
nand U9134 (N_9134,N_8356,N_7729);
and U9135 (N_9135,N_8842,N_8766);
xor U9136 (N_9136,N_7865,N_7985);
or U9137 (N_9137,N_8868,N_8572);
and U9138 (N_9138,N_8229,N_8388);
or U9139 (N_9139,N_8259,N_8062);
nand U9140 (N_9140,N_8373,N_8581);
nor U9141 (N_9141,N_8635,N_8358);
or U9142 (N_9142,N_8519,N_7596);
and U9143 (N_9143,N_8392,N_7607);
nor U9144 (N_9144,N_8858,N_8064);
or U9145 (N_9145,N_8494,N_8570);
and U9146 (N_9146,N_8871,N_7533);
and U9147 (N_9147,N_8404,N_8187);
and U9148 (N_9148,N_7502,N_7947);
or U9149 (N_9149,N_7567,N_7744);
nand U9150 (N_9150,N_8692,N_8122);
and U9151 (N_9151,N_8257,N_8220);
and U9152 (N_9152,N_8308,N_8090);
and U9153 (N_9153,N_7595,N_8092);
or U9154 (N_9154,N_8694,N_7735);
or U9155 (N_9155,N_8233,N_8402);
xor U9156 (N_9156,N_8365,N_7833);
nand U9157 (N_9157,N_7849,N_8319);
and U9158 (N_9158,N_7893,N_8323);
nor U9159 (N_9159,N_8422,N_8182);
and U9160 (N_9160,N_8947,N_8491);
and U9161 (N_9161,N_8267,N_8790);
nand U9162 (N_9162,N_7952,N_8234);
or U9163 (N_9163,N_8421,N_8615);
nor U9164 (N_9164,N_8844,N_7756);
and U9165 (N_9165,N_8838,N_7570);
and U9166 (N_9166,N_7576,N_8406);
nor U9167 (N_9167,N_7762,N_7769);
nand U9168 (N_9168,N_7776,N_8811);
or U9169 (N_9169,N_8451,N_7945);
nand U9170 (N_9170,N_7571,N_8799);
or U9171 (N_9171,N_7926,N_8877);
or U9172 (N_9172,N_8195,N_7889);
or U9173 (N_9173,N_8129,N_8078);
nand U9174 (N_9174,N_7976,N_7960);
nor U9175 (N_9175,N_8726,N_8029);
and U9176 (N_9176,N_8541,N_7659);
xnor U9177 (N_9177,N_8595,N_8468);
nor U9178 (N_9178,N_7784,N_8228);
nor U9179 (N_9179,N_8438,N_7828);
nor U9180 (N_9180,N_8994,N_8363);
or U9181 (N_9181,N_8722,N_7528);
nand U9182 (N_9182,N_8927,N_8728);
and U9183 (N_9183,N_8416,N_8218);
xnor U9184 (N_9184,N_8652,N_8702);
or U9185 (N_9185,N_8669,N_8600);
nor U9186 (N_9186,N_8575,N_7964);
and U9187 (N_9187,N_8466,N_8569);
xor U9188 (N_9188,N_8212,N_8000);
xnor U9189 (N_9189,N_8277,N_7871);
xor U9190 (N_9190,N_8828,N_7905);
or U9191 (N_9191,N_8203,N_8350);
nor U9192 (N_9192,N_8712,N_8236);
nand U9193 (N_9193,N_8019,N_8032);
nand U9194 (N_9194,N_7675,N_8951);
nand U9195 (N_9195,N_7753,N_7998);
nor U9196 (N_9196,N_8351,N_7717);
nor U9197 (N_9197,N_8859,N_8139);
or U9198 (N_9198,N_7823,N_7593);
nand U9199 (N_9199,N_7718,N_7838);
nand U9200 (N_9200,N_8924,N_8176);
nand U9201 (N_9201,N_7637,N_8240);
nor U9202 (N_9202,N_7977,N_8530);
nor U9203 (N_9203,N_8737,N_8550);
and U9204 (N_9204,N_8609,N_8825);
or U9205 (N_9205,N_7760,N_8553);
nand U9206 (N_9206,N_8433,N_7851);
or U9207 (N_9207,N_8215,N_8150);
or U9208 (N_9208,N_8298,N_8080);
nor U9209 (N_9209,N_7805,N_8711);
and U9210 (N_9210,N_7886,N_8646);
nand U9211 (N_9211,N_7825,N_7712);
and U9212 (N_9212,N_8606,N_8368);
or U9213 (N_9213,N_8457,N_8489);
nand U9214 (N_9214,N_8852,N_8174);
xnor U9215 (N_9215,N_7808,N_7515);
and U9216 (N_9216,N_7821,N_7829);
nor U9217 (N_9217,N_8269,N_8593);
xnor U9218 (N_9218,N_8549,N_8608);
nor U9219 (N_9219,N_7663,N_8241);
or U9220 (N_9220,N_8446,N_7711);
nand U9221 (N_9221,N_8913,N_7701);
nand U9222 (N_9222,N_8898,N_8684);
or U9223 (N_9223,N_8177,N_8039);
nand U9224 (N_9224,N_8839,N_7980);
and U9225 (N_9225,N_8025,N_7696);
xor U9226 (N_9226,N_8528,N_8455);
nor U9227 (N_9227,N_8274,N_8382);
xor U9228 (N_9228,N_8848,N_8982);
nand U9229 (N_9229,N_7700,N_8202);
nand U9230 (N_9230,N_8474,N_8500);
nor U9231 (N_9231,N_7866,N_8698);
nor U9232 (N_9232,N_8797,N_8673);
and U9233 (N_9233,N_8181,N_7631);
and U9234 (N_9234,N_7872,N_8126);
nor U9235 (N_9235,N_8246,N_7780);
nand U9236 (N_9236,N_7503,N_7629);
nor U9237 (N_9237,N_8326,N_8546);
and U9238 (N_9238,N_8396,N_8562);
or U9239 (N_9239,N_8561,N_8081);
nor U9240 (N_9240,N_8118,N_8818);
and U9241 (N_9241,N_8629,N_8094);
nand U9242 (N_9242,N_7817,N_7692);
nand U9243 (N_9243,N_8026,N_7623);
nor U9244 (N_9244,N_8695,N_7691);
nor U9245 (N_9245,N_8809,N_7782);
or U9246 (N_9246,N_8021,N_8285);
and U9247 (N_9247,N_8666,N_8079);
nor U9248 (N_9248,N_8544,N_8535);
nor U9249 (N_9249,N_7772,N_7804);
and U9250 (N_9250,N_8354,N_8603);
and U9251 (N_9251,N_7830,N_8996);
nor U9252 (N_9252,N_7747,N_8023);
nand U9253 (N_9253,N_8810,N_8596);
and U9254 (N_9254,N_8946,N_8276);
nor U9255 (N_9255,N_8167,N_8410);
and U9256 (N_9256,N_8340,N_8584);
xnor U9257 (N_9257,N_7539,N_7818);
or U9258 (N_9258,N_8302,N_8391);
nor U9259 (N_9259,N_8164,N_8703);
nand U9260 (N_9260,N_8278,N_8149);
nand U9261 (N_9261,N_8620,N_7885);
or U9262 (N_9262,N_8447,N_8853);
nor U9263 (N_9263,N_8245,N_7999);
nor U9264 (N_9264,N_7709,N_8933);
or U9265 (N_9265,N_7937,N_7794);
nand U9266 (N_9266,N_8386,N_7819);
or U9267 (N_9267,N_7800,N_8266);
nor U9268 (N_9268,N_7640,N_8102);
and U9269 (N_9269,N_8338,N_7920);
nand U9270 (N_9270,N_8296,N_8357);
or U9271 (N_9271,N_7995,N_7618);
nand U9272 (N_9272,N_8471,N_8286);
xnor U9273 (N_9273,N_7903,N_7930);
and U9274 (N_9274,N_7560,N_8197);
and U9275 (N_9275,N_8835,N_7909);
or U9276 (N_9276,N_7754,N_8255);
or U9277 (N_9277,N_8688,N_8315);
and U9278 (N_9278,N_8030,N_8487);
and U9279 (N_9279,N_8018,N_8781);
and U9280 (N_9280,N_7648,N_8914);
xnor U9281 (N_9281,N_7854,N_8677);
xnor U9282 (N_9282,N_8040,N_8288);
nand U9283 (N_9283,N_8359,N_7890);
nor U9284 (N_9284,N_8622,N_7635);
nor U9285 (N_9285,N_7604,N_8097);
nand U9286 (N_9286,N_8105,N_8725);
nand U9287 (N_9287,N_7958,N_7510);
or U9288 (N_9288,N_8361,N_8939);
nand U9289 (N_9289,N_7506,N_8015);
xor U9290 (N_9290,N_8303,N_7577);
nand U9291 (N_9291,N_8979,N_8873);
and U9292 (N_9292,N_8515,N_8732);
or U9293 (N_9293,N_8837,N_8109);
xor U9294 (N_9294,N_8311,N_8157);
or U9295 (N_9295,N_8630,N_8901);
or U9296 (N_9296,N_8934,N_8536);
or U9297 (N_9297,N_8910,N_8509);
nand U9298 (N_9298,N_7583,N_8610);
or U9299 (N_9299,N_8033,N_7563);
nor U9300 (N_9300,N_8867,N_7759);
nand U9301 (N_9301,N_8325,N_8314);
and U9302 (N_9302,N_8628,N_8592);
nor U9303 (N_9303,N_8372,N_7894);
or U9304 (N_9304,N_8641,N_8788);
xnor U9305 (N_9305,N_8769,N_7775);
nand U9306 (N_9306,N_8778,N_8959);
nor U9307 (N_9307,N_7514,N_8896);
nand U9308 (N_9308,N_8685,N_8133);
or U9309 (N_9309,N_7877,N_7522);
xnor U9310 (N_9310,N_7959,N_8339);
or U9311 (N_9311,N_7612,N_8627);
and U9312 (N_9312,N_8887,N_8393);
xor U9313 (N_9313,N_8121,N_8578);
and U9314 (N_9314,N_7831,N_8559);
nand U9315 (N_9315,N_8763,N_8587);
nand U9316 (N_9316,N_7521,N_8112);
nand U9317 (N_9317,N_8998,N_8662);
xor U9318 (N_9318,N_7697,N_7500);
and U9319 (N_9319,N_8069,N_8120);
nand U9320 (N_9320,N_8124,N_7869);
xnor U9321 (N_9321,N_8367,N_7739);
or U9322 (N_9322,N_7624,N_7874);
or U9323 (N_9323,N_8411,N_8750);
nor U9324 (N_9324,N_7574,N_8189);
xor U9325 (N_9325,N_8072,N_7850);
xor U9326 (N_9326,N_8089,N_8502);
or U9327 (N_9327,N_8279,N_8897);
nor U9328 (N_9328,N_8589,N_7685);
nand U9329 (N_9329,N_8558,N_8087);
nor U9330 (N_9330,N_8771,N_8618);
and U9331 (N_9331,N_7806,N_8821);
nor U9332 (N_9332,N_7837,N_7501);
xnor U9333 (N_9333,N_7993,N_8071);
or U9334 (N_9334,N_8292,N_8199);
nand U9335 (N_9335,N_8847,N_8371);
nand U9336 (N_9336,N_7743,N_8070);
and U9337 (N_9337,N_8990,N_8272);
nand U9338 (N_9338,N_8547,N_8524);
nor U9339 (N_9339,N_7546,N_8642);
or U9340 (N_9340,N_8440,N_7979);
nor U9341 (N_9341,N_7752,N_8905);
nand U9342 (N_9342,N_8035,N_8850);
or U9343 (N_9343,N_7540,N_7771);
xor U9344 (N_9344,N_8170,N_8496);
or U9345 (N_9345,N_7557,N_8972);
nand U9346 (N_9346,N_7988,N_8076);
nor U9347 (N_9347,N_8225,N_8162);
and U9348 (N_9348,N_8191,N_8683);
and U9349 (N_9349,N_7633,N_8663);
and U9350 (N_9350,N_8281,N_7919);
nand U9351 (N_9351,N_8188,N_8534);
and U9352 (N_9352,N_7940,N_8970);
or U9353 (N_9353,N_8525,N_7834);
or U9354 (N_9354,N_7907,N_8417);
or U9355 (N_9355,N_8583,N_8495);
and U9356 (N_9356,N_7627,N_8116);
or U9357 (N_9357,N_8424,N_7597);
and U9358 (N_9358,N_8803,N_7941);
nand U9359 (N_9359,N_7836,N_8473);
or U9360 (N_9360,N_7895,N_8704);
and U9361 (N_9361,N_8949,N_8165);
nor U9362 (N_9362,N_7632,N_8879);
or U9363 (N_9363,N_7789,N_7839);
and U9364 (N_9364,N_8731,N_7878);
xor U9365 (N_9365,N_8060,N_7897);
and U9366 (N_9366,N_7733,N_8654);
nand U9367 (N_9367,N_8507,N_7513);
or U9368 (N_9368,N_8758,N_8755);
or U9369 (N_9369,N_8486,N_7931);
or U9370 (N_9370,N_7606,N_7899);
xnor U9371 (N_9371,N_7672,N_7859);
and U9372 (N_9372,N_8957,N_7928);
and U9373 (N_9373,N_7788,N_8754);
and U9374 (N_9374,N_8510,N_8012);
nand U9375 (N_9375,N_7911,N_8458);
xnor U9376 (N_9376,N_8634,N_7508);
and U9377 (N_9377,N_8816,N_8395);
nand U9378 (N_9378,N_8883,N_8379);
or U9379 (N_9379,N_8123,N_8591);
or U9380 (N_9380,N_8743,N_7534);
nor U9381 (N_9381,N_8938,N_7791);
or U9382 (N_9382,N_8506,N_8115);
and U9383 (N_9383,N_8332,N_7594);
nand U9384 (N_9384,N_7638,N_8942);
nand U9385 (N_9385,N_8130,N_8221);
nor U9386 (N_9386,N_7730,N_8701);
or U9387 (N_9387,N_8082,N_7795);
and U9388 (N_9388,N_8777,N_8464);
and U9389 (N_9389,N_8890,N_8527);
and U9390 (N_9390,N_8439,N_7918);
nor U9391 (N_9391,N_8742,N_8096);
nand U9392 (N_9392,N_7970,N_8909);
or U9393 (N_9393,N_8052,N_7863);
xnor U9394 (N_9394,N_8567,N_8976);
or U9395 (N_9395,N_7535,N_7856);
nand U9396 (N_9396,N_8375,N_7896);
or U9397 (N_9397,N_8201,N_7868);
or U9398 (N_9398,N_8953,N_7876);
nand U9399 (N_9399,N_8437,N_8585);
or U9400 (N_9400,N_8955,N_8280);
or U9401 (N_9401,N_7660,N_8318);
and U9402 (N_9402,N_8672,N_7974);
xor U9403 (N_9403,N_8727,N_8876);
xnor U9404 (N_9404,N_8103,N_7714);
nor U9405 (N_9405,N_8493,N_8399);
nand U9406 (N_9406,N_8046,N_8222);
nor U9407 (N_9407,N_8926,N_8813);
xnor U9408 (N_9408,N_7548,N_8571);
nor U9409 (N_9409,N_8794,N_7720);
xnor U9410 (N_9410,N_8144,N_8248);
or U9411 (N_9411,N_8260,N_8804);
nand U9412 (N_9412,N_8538,N_7537);
nor U9413 (N_9413,N_8865,N_7891);
or U9414 (N_9414,N_7848,N_7532);
xor U9415 (N_9415,N_8605,N_7860);
nor U9416 (N_9416,N_7750,N_7873);
or U9417 (N_9417,N_8024,N_8289);
and U9418 (N_9418,N_8465,N_8007);
xor U9419 (N_9419,N_7628,N_8003);
nand U9420 (N_9420,N_8329,N_7644);
or U9421 (N_9421,N_8577,N_7881);
and U9422 (N_9422,N_8614,N_7827);
nor U9423 (N_9423,N_8954,N_8805);
xnor U9424 (N_9424,N_7687,N_8738);
and U9425 (N_9425,N_8263,N_7680);
nand U9426 (N_9426,N_8709,N_8961);
nor U9427 (N_9427,N_8902,N_7942);
or U9428 (N_9428,N_7867,N_8208);
or U9429 (N_9429,N_8231,N_8084);
or U9430 (N_9430,N_8352,N_7814);
or U9431 (N_9431,N_8894,N_8327);
nand U9432 (N_9432,N_7575,N_7973);
nand U9433 (N_9433,N_7556,N_7620);
nand U9434 (N_9434,N_8626,N_8503);
or U9435 (N_9435,N_8829,N_7590);
and U9436 (N_9436,N_8590,N_7716);
nor U9437 (N_9437,N_7971,N_7666);
or U9438 (N_9438,N_7767,N_7566);
and U9439 (N_9439,N_8461,N_7758);
or U9440 (N_9440,N_8378,N_8819);
xor U9441 (N_9441,N_8376,N_8657);
nor U9442 (N_9442,N_8529,N_7965);
and U9443 (N_9443,N_8760,N_8597);
xor U9444 (N_9444,N_8283,N_8028);
nand U9445 (N_9445,N_7674,N_8321);
nor U9446 (N_9446,N_7667,N_8113);
or U9447 (N_9447,N_7676,N_8059);
or U9448 (N_9448,N_8987,N_7832);
nand U9449 (N_9449,N_8083,N_8940);
or U9450 (N_9450,N_8748,N_7820);
and U9451 (N_9451,N_7561,N_8782);
nand U9452 (N_9452,N_8077,N_7957);
nand U9453 (N_9453,N_8293,N_8708);
nand U9454 (N_9454,N_7870,N_8235);
or U9455 (N_9455,N_7742,N_7923);
nor U9456 (N_9456,N_7519,N_8042);
or U9457 (N_9457,N_7559,N_8312);
and U9458 (N_9458,N_8916,N_7652);
nand U9459 (N_9459,N_7887,N_7996);
nor U9460 (N_9460,N_8721,N_7843);
or U9461 (N_9461,N_7732,N_8611);
nand U9462 (N_9462,N_8952,N_8864);
and U9463 (N_9463,N_8607,N_7531);
or U9464 (N_9464,N_7783,N_8377);
nand U9465 (N_9465,N_8875,N_8131);
nand U9466 (N_9466,N_7706,N_8730);
nor U9467 (N_9467,N_7906,N_8390);
and U9468 (N_9468,N_7662,N_7654);
nor U9469 (N_9469,N_8911,N_7728);
nor U9470 (N_9470,N_7845,N_7936);
or U9471 (N_9471,N_8999,N_8888);
nand U9472 (N_9472,N_8161,N_8557);
and U9473 (N_9473,N_8710,N_8186);
and U9474 (N_9474,N_7669,N_7749);
or U9475 (N_9475,N_8980,N_8100);
nor U9476 (N_9476,N_8063,N_8200);
and U9477 (N_9477,N_8290,N_8925);
or U9478 (N_9478,N_8917,N_7523);
nand U9479 (N_9479,N_8705,N_8226);
nand U9480 (N_9480,N_8010,N_8793);
nand U9481 (N_9481,N_8127,N_7852);
and U9482 (N_9482,N_7785,N_8305);
and U9483 (N_9483,N_7948,N_8670);
nor U9484 (N_9484,N_7857,N_8454);
nand U9485 (N_9485,N_8159,N_7792);
and U9486 (N_9486,N_7554,N_7582);
nor U9487 (N_9487,N_8425,N_7643);
or U9488 (N_9488,N_8309,N_7578);
or U9489 (N_9489,N_8227,N_8484);
and U9490 (N_9490,N_8780,N_8700);
and U9491 (N_9491,N_8676,N_8659);
or U9492 (N_9492,N_7516,N_8400);
or U9493 (N_9493,N_8238,N_8775);
or U9494 (N_9494,N_8744,N_8055);
nand U9495 (N_9495,N_8160,N_8759);
or U9496 (N_9496,N_8085,N_8747);
or U9497 (N_9497,N_8997,N_8991);
nand U9498 (N_9498,N_8068,N_8282);
nand U9499 (N_9499,N_8004,N_8366);
nand U9500 (N_9500,N_8671,N_8586);
or U9501 (N_9501,N_7992,N_8247);
or U9502 (N_9502,N_7922,N_8995);
nor U9503 (N_9503,N_8008,N_7944);
nand U9504 (N_9504,N_7768,N_8746);
and U9505 (N_9505,N_8560,N_8180);
and U9506 (N_9506,N_7809,N_8574);
nor U9507 (N_9507,N_8107,N_8812);
xnor U9508 (N_9508,N_8814,N_8716);
and U9509 (N_9509,N_8114,N_8678);
or U9510 (N_9510,N_8983,N_8460);
or U9511 (N_9511,N_7844,N_8445);
xor U9512 (N_9512,N_8706,N_7765);
or U9513 (N_9513,N_8638,N_8009);
nor U9514 (N_9514,N_8194,N_8900);
nor U9515 (N_9515,N_7653,N_8154);
and U9516 (N_9516,N_7562,N_8313);
nand U9517 (N_9517,N_7751,N_8335);
nor U9518 (N_9518,N_7855,N_8516);
xor U9519 (N_9519,N_7840,N_7686);
nor U9520 (N_9520,N_7713,N_8625);
or U9521 (N_9521,N_8881,N_8217);
nand U9522 (N_9522,N_8432,N_7565);
and U9523 (N_9523,N_7984,N_7737);
nand U9524 (N_9524,N_8932,N_8903);
nor U9525 (N_9525,N_7549,N_7847);
nor U9526 (N_9526,N_7655,N_8661);
nor U9527 (N_9527,N_8885,N_8251);
nor U9528 (N_9528,N_8478,N_8355);
or U9529 (N_9529,N_8106,N_8011);
or U9530 (N_9530,N_7664,N_8173);
nor U9531 (N_9531,N_7509,N_7661);
nor U9532 (N_9532,N_8936,N_8792);
and U9533 (N_9533,N_8993,N_8216);
nand U9534 (N_9534,N_8565,N_8207);
or U9535 (N_9535,N_8397,N_7657);
or U9536 (N_9536,N_8863,N_8364);
or U9537 (N_9537,N_8967,N_8333);
nand U9538 (N_9538,N_8846,N_7746);
xor U9539 (N_9539,N_8832,N_7740);
or U9540 (N_9540,N_8268,N_8632);
nor U9541 (N_9541,N_8598,N_8715);
and U9542 (N_9542,N_7723,N_7719);
or U9543 (N_9543,N_8764,N_8341);
xnor U9544 (N_9544,N_8893,N_8542);
xor U9545 (N_9545,N_8017,N_8459);
xnor U9546 (N_9546,N_8962,N_7524);
xor U9547 (N_9547,N_8224,N_8923);
nand U9548 (N_9548,N_8770,N_8717);
nor U9549 (N_9549,N_7778,N_8091);
nor U9550 (N_9550,N_8822,N_8827);
nor U9551 (N_9551,N_7589,N_7921);
nor U9552 (N_9552,N_8650,N_8806);
nand U9553 (N_9553,N_8398,N_7678);
or U9554 (N_9554,N_8944,N_7912);
and U9555 (N_9555,N_7724,N_7813);
nand U9556 (N_9556,N_8415,N_8655);
or U9557 (N_9557,N_7981,N_7862);
and U9558 (N_9558,N_8204,N_8637);
and U9559 (N_9559,N_8649,N_8552);
nand U9560 (N_9560,N_8679,N_7797);
and U9561 (N_9561,N_8275,N_7888);
xor U9562 (N_9562,N_8579,N_8134);
xor U9563 (N_9563,N_7822,N_8992);
xnor U9564 (N_9564,N_8456,N_8418);
xnor U9565 (N_9565,N_8230,N_7580);
nor U9566 (N_9566,N_8067,N_8749);
nor U9567 (N_9567,N_8522,N_8168);
xnor U9568 (N_9568,N_8551,N_7967);
or U9569 (N_9569,N_7703,N_8370);
or U9570 (N_9570,N_7901,N_7766);
or U9571 (N_9571,N_8682,N_8449);
nand U9572 (N_9572,N_8306,N_8117);
xor U9573 (N_9573,N_7544,N_8714);
nand U9574 (N_9574,N_7879,N_8322);
nand U9575 (N_9575,N_7904,N_8582);
and U9576 (N_9576,N_8723,N_8718);
nor U9577 (N_9577,N_8140,N_8101);
nor U9578 (N_9578,N_8210,N_7978);
nor U9579 (N_9579,N_7721,N_7731);
and U9580 (N_9580,N_8619,N_8499);
nand U9581 (N_9581,N_8964,N_8175);
nor U9582 (N_9582,N_7639,N_8328);
or U9583 (N_9583,N_7710,N_7681);
nor U9584 (N_9584,N_8691,N_8831);
xnor U9585 (N_9585,N_7599,N_7861);
and U9586 (N_9586,N_8504,N_8347);
nor U9587 (N_9587,N_8602,N_7949);
and U9588 (N_9588,N_7646,N_8041);
xor U9589 (N_9589,N_8490,N_8741);
and U9590 (N_9590,N_7630,N_8707);
and U9591 (N_9591,N_8074,N_8668);
or U9592 (N_9592,N_8874,N_8518);
nand U9593 (N_9593,N_8511,N_8966);
nand U9594 (N_9594,N_8624,N_8057);
or U9595 (N_9595,N_8488,N_8151);
or U9596 (N_9596,N_8334,N_8573);
nor U9597 (N_9597,N_8845,N_7677);
xnor U9598 (N_9598,N_8450,N_8880);
nand U9599 (N_9599,N_8651,N_8211);
nor U9600 (N_9600,N_7520,N_7641);
nand U9601 (N_9601,N_8066,N_8689);
nand U9602 (N_9602,N_8855,N_7916);
xnor U9603 (N_9603,N_8481,N_8435);
and U9604 (N_9604,N_7799,N_8349);
xnor U9605 (N_9605,N_8497,N_8434);
and U9606 (N_9606,N_7707,N_7826);
nor U9607 (N_9607,N_8038,N_8720);
nand U9608 (N_9608,N_7933,N_8643);
and U9609 (N_9609,N_8307,N_8904);
nor U9610 (N_9610,N_8640,N_8779);
nand U9611 (N_9611,N_8184,N_7598);
or U9612 (N_9612,N_8886,N_8270);
nand U9613 (N_9613,N_8384,N_8907);
and U9614 (N_9614,N_8463,N_8256);
and U9615 (N_9615,N_8430,N_8776);
or U9616 (N_9616,N_8696,N_7708);
and U9617 (N_9617,N_8002,N_7913);
and U9618 (N_9618,N_7649,N_8791);
nor U9619 (N_9619,N_8369,N_8753);
and U9620 (N_9620,N_8601,N_8543);
nor U9621 (N_9621,N_8016,N_7682);
nand U9622 (N_9622,N_8783,N_8767);
nor U9623 (N_9623,N_8093,N_8110);
nand U9624 (N_9624,N_8965,N_8548);
and U9625 (N_9625,N_8420,N_8719);
nor U9626 (N_9626,N_8027,N_8580);
or U9627 (N_9627,N_7656,N_8166);
and U9628 (N_9628,N_8053,N_7892);
xor U9629 (N_9629,N_8403,N_8681);
nand U9630 (N_9630,N_7616,N_8273);
and U9631 (N_9631,N_8736,N_8143);
and U9632 (N_9632,N_8505,N_8442);
nor U9633 (N_9633,N_7801,N_8599);
and U9634 (N_9634,N_8693,N_8653);
nor U9635 (N_9635,N_8196,N_8047);
xor U9636 (N_9636,N_7695,N_7986);
xor U9637 (N_9637,N_7807,N_7846);
xnor U9638 (N_9638,N_7587,N_8800);
nor U9639 (N_9639,N_8836,N_7725);
or U9640 (N_9640,N_7841,N_8345);
and U9641 (N_9641,N_8616,N_8137);
nand U9642 (N_9642,N_8383,N_8647);
or U9643 (N_9643,N_8697,N_7591);
nor U9644 (N_9644,N_8860,N_8443);
and U9645 (N_9645,N_8244,N_8756);
or U9646 (N_9646,N_8631,N_8922);
and U9647 (N_9647,N_8469,N_7690);
and U9648 (N_9648,N_8699,N_7645);
and U9649 (N_9649,N_7601,N_7736);
or U9650 (N_9650,N_7983,N_8849);
nor U9651 (N_9651,N_8095,N_7610);
nand U9652 (N_9652,N_8190,N_8973);
and U9653 (N_9653,N_8588,N_7815);
nand U9654 (N_9654,N_7505,N_7543);
or U9655 (N_9655,N_8142,N_8304);
xnor U9656 (N_9656,N_8385,N_8128);
nand U9657 (N_9657,N_8237,N_8477);
nor U9658 (N_9658,N_7741,N_7798);
or U9659 (N_9659,N_8919,N_8470);
and U9660 (N_9660,N_8193,N_8943);
nor U9661 (N_9661,N_8036,N_8521);
nor U9662 (N_9662,N_7917,N_7908);
nor U9663 (N_9663,N_8841,N_8409);
xor U9664 (N_9664,N_8374,N_8648);
or U9665 (N_9665,N_8452,N_8824);
nor U9666 (N_9666,N_8098,N_8941);
nor U9667 (N_9667,N_7803,N_8665);
nand U9668 (N_9668,N_7734,N_8073);
xor U9669 (N_9669,N_7961,N_8745);
nor U9670 (N_9670,N_7934,N_8058);
and U9671 (N_9671,N_7665,N_8419);
nand U9672 (N_9672,N_8317,N_7994);
or U9673 (N_9673,N_7689,N_7552);
nor U9674 (N_9674,N_8882,N_8872);
xnor U9675 (N_9675,N_8163,N_8348);
nand U9676 (N_9676,N_8483,N_7634);
nand U9677 (N_9677,N_8453,N_7816);
nand U9678 (N_9678,N_7647,N_7824);
or U9679 (N_9679,N_8169,N_8978);
and U9680 (N_9680,N_8594,N_8014);
and U9681 (N_9681,N_7608,N_7613);
nor U9682 (N_9682,N_7525,N_8724);
or U9683 (N_9683,N_7935,N_8807);
and U9684 (N_9684,N_8132,N_8658);
or U9685 (N_9685,N_8295,N_8394);
nand U9686 (N_9686,N_8912,N_8533);
and U9687 (N_9687,N_8878,N_8209);
or U9688 (N_9688,N_8786,N_7518);
nor U9689 (N_9689,N_7512,N_7579);
nor U9690 (N_9690,N_7910,N_7569);
and U9691 (N_9691,N_8299,N_7558);
nand U9692 (N_9692,N_8664,N_7584);
and U9693 (N_9693,N_8774,N_7875);
or U9694 (N_9694,N_8146,N_8287);
nor U9695 (N_9695,N_8243,N_7774);
or U9696 (N_9696,N_7617,N_7568);
or U9697 (N_9697,N_7883,N_7972);
or U9698 (N_9698,N_8049,N_8958);
or U9699 (N_9699,N_8336,N_7902);
and U9700 (N_9700,N_8044,N_7668);
nand U9701 (N_9701,N_7757,N_8826);
nor U9702 (N_9702,N_8801,N_8423);
nand U9703 (N_9703,N_8232,N_8891);
nor U9704 (N_9704,N_8320,N_8554);
nand U9705 (N_9705,N_7650,N_8405);
and U9706 (N_9706,N_8061,N_7602);
and U9707 (N_9707,N_8297,N_8381);
nand U9708 (N_9708,N_7811,N_7924);
and U9709 (N_9709,N_8977,N_8178);
and U9710 (N_9710,N_8022,N_8667);
nor U9711 (N_9711,N_7550,N_7777);
and U9712 (N_9712,N_7764,N_7542);
or U9713 (N_9713,N_7770,N_8765);
nand U9714 (N_9714,N_8928,N_8751);
or U9715 (N_9715,N_8513,N_8555);
nand U9716 (N_9716,N_8360,N_7547);
nand U9717 (N_9717,N_7722,N_8258);
or U9718 (N_9718,N_8660,N_8005);
nand U9719 (N_9719,N_8856,N_8948);
nor U9720 (N_9720,N_8148,N_7755);
or U9721 (N_9721,N_8171,N_8735);
nand U9722 (N_9722,N_7538,N_8020);
xnor U9723 (N_9723,N_8213,N_8843);
and U9724 (N_9724,N_7555,N_8656);
or U9725 (N_9725,N_7929,N_7673);
and U9726 (N_9726,N_7615,N_7975);
or U9727 (N_9727,N_7946,N_8065);
nand U9728 (N_9728,N_8472,N_7536);
and U9729 (N_9729,N_8346,N_7564);
nor U9730 (N_9730,N_8539,N_7651);
or U9731 (N_9731,N_8104,N_8056);
or U9732 (N_9732,N_7715,N_8239);
or U9733 (N_9733,N_8645,N_7527);
or U9734 (N_9734,N_8413,N_7748);
xor U9735 (N_9735,N_8929,N_8108);
nor U9736 (N_9736,N_8937,N_8817);
nand U9737 (N_9737,N_7671,N_8971);
or U9738 (N_9738,N_7600,N_8185);
and U9739 (N_9739,N_7551,N_8931);
nor U9740 (N_9740,N_8734,N_8802);
nor U9741 (N_9741,N_8918,N_8739);
and U9742 (N_9742,N_8198,N_8219);
nand U9743 (N_9743,N_7915,N_7802);
nand U9744 (N_9744,N_8254,N_7625);
nor U9745 (N_9745,N_8264,N_8733);
nand U9746 (N_9746,N_8362,N_8389);
or U9747 (N_9747,N_8935,N_7953);
nand U9748 (N_9748,N_7939,N_8820);
or U9749 (N_9749,N_8869,N_8223);
or U9750 (N_9750,N_7885,N_7909);
nand U9751 (N_9751,N_8916,N_7738);
or U9752 (N_9752,N_8390,N_8911);
and U9753 (N_9753,N_7645,N_8658);
xnor U9754 (N_9754,N_7652,N_8194);
or U9755 (N_9755,N_7833,N_7732);
or U9756 (N_9756,N_8858,N_8919);
nand U9757 (N_9757,N_8678,N_7813);
nor U9758 (N_9758,N_8940,N_8741);
nand U9759 (N_9759,N_7979,N_7972);
nor U9760 (N_9760,N_8715,N_8260);
nand U9761 (N_9761,N_7763,N_8794);
nor U9762 (N_9762,N_7860,N_8752);
or U9763 (N_9763,N_7932,N_8406);
nand U9764 (N_9764,N_7574,N_7628);
xor U9765 (N_9765,N_8283,N_7841);
and U9766 (N_9766,N_8381,N_8937);
or U9767 (N_9767,N_7966,N_8335);
nand U9768 (N_9768,N_8730,N_8476);
nor U9769 (N_9769,N_7932,N_7972);
nor U9770 (N_9770,N_8540,N_8296);
xnor U9771 (N_9771,N_8248,N_8800);
nand U9772 (N_9772,N_7577,N_7874);
or U9773 (N_9773,N_7533,N_7686);
nor U9774 (N_9774,N_8992,N_7538);
nor U9775 (N_9775,N_8395,N_7604);
or U9776 (N_9776,N_8137,N_8399);
nor U9777 (N_9777,N_8551,N_8869);
or U9778 (N_9778,N_8429,N_8048);
nor U9779 (N_9779,N_8978,N_8321);
nor U9780 (N_9780,N_7840,N_8240);
and U9781 (N_9781,N_8600,N_8061);
nand U9782 (N_9782,N_8052,N_8883);
nor U9783 (N_9783,N_8515,N_8695);
and U9784 (N_9784,N_7820,N_7513);
or U9785 (N_9785,N_7715,N_7512);
nand U9786 (N_9786,N_7604,N_8084);
xor U9787 (N_9787,N_8905,N_8671);
nand U9788 (N_9788,N_7980,N_8756);
nand U9789 (N_9789,N_7768,N_7890);
nor U9790 (N_9790,N_8411,N_8796);
and U9791 (N_9791,N_8359,N_8335);
xor U9792 (N_9792,N_8530,N_8044);
nor U9793 (N_9793,N_8548,N_8559);
nor U9794 (N_9794,N_8312,N_7651);
xnor U9795 (N_9795,N_8315,N_8720);
nand U9796 (N_9796,N_7736,N_7858);
nand U9797 (N_9797,N_7737,N_8850);
and U9798 (N_9798,N_7934,N_7968);
nor U9799 (N_9799,N_8503,N_8513);
xnor U9800 (N_9800,N_7923,N_8501);
nor U9801 (N_9801,N_7586,N_8878);
nor U9802 (N_9802,N_8743,N_7828);
nor U9803 (N_9803,N_8010,N_8696);
nor U9804 (N_9804,N_8175,N_7832);
nor U9805 (N_9805,N_7944,N_7680);
nor U9806 (N_9806,N_7509,N_7971);
nor U9807 (N_9807,N_7591,N_7908);
and U9808 (N_9808,N_7969,N_8577);
nand U9809 (N_9809,N_8263,N_8887);
nor U9810 (N_9810,N_7851,N_7800);
nor U9811 (N_9811,N_8438,N_8626);
nor U9812 (N_9812,N_8191,N_8975);
or U9813 (N_9813,N_7512,N_7772);
nor U9814 (N_9814,N_8022,N_8402);
nor U9815 (N_9815,N_8874,N_8741);
nor U9816 (N_9816,N_8871,N_7734);
xor U9817 (N_9817,N_7946,N_8387);
and U9818 (N_9818,N_8637,N_8346);
nand U9819 (N_9819,N_8030,N_8803);
xnor U9820 (N_9820,N_8459,N_7685);
nand U9821 (N_9821,N_8957,N_8047);
nor U9822 (N_9822,N_8232,N_8306);
and U9823 (N_9823,N_7511,N_8499);
xor U9824 (N_9824,N_8318,N_7689);
nand U9825 (N_9825,N_8149,N_8657);
xnor U9826 (N_9826,N_8853,N_8410);
nor U9827 (N_9827,N_8913,N_7838);
or U9828 (N_9828,N_8615,N_8017);
and U9829 (N_9829,N_8279,N_7992);
nand U9830 (N_9830,N_8845,N_7809);
and U9831 (N_9831,N_8476,N_8967);
nor U9832 (N_9832,N_7803,N_8624);
and U9833 (N_9833,N_8947,N_8294);
and U9834 (N_9834,N_7923,N_8409);
and U9835 (N_9835,N_8271,N_8298);
and U9836 (N_9836,N_8305,N_8287);
and U9837 (N_9837,N_7648,N_8589);
xnor U9838 (N_9838,N_7818,N_7777);
or U9839 (N_9839,N_8394,N_8509);
or U9840 (N_9840,N_7538,N_8124);
and U9841 (N_9841,N_8351,N_7793);
nand U9842 (N_9842,N_8434,N_8023);
nand U9843 (N_9843,N_8736,N_8132);
and U9844 (N_9844,N_8482,N_8720);
or U9845 (N_9845,N_8522,N_7971);
nor U9846 (N_9846,N_8438,N_7813);
nor U9847 (N_9847,N_8281,N_7777);
nand U9848 (N_9848,N_7938,N_8751);
xnor U9849 (N_9849,N_8067,N_7705);
nor U9850 (N_9850,N_8236,N_7745);
and U9851 (N_9851,N_8393,N_8826);
nor U9852 (N_9852,N_8149,N_8685);
or U9853 (N_9853,N_8878,N_8311);
or U9854 (N_9854,N_8158,N_8771);
nand U9855 (N_9855,N_8126,N_8424);
xnor U9856 (N_9856,N_7922,N_8619);
or U9857 (N_9857,N_8133,N_8512);
nand U9858 (N_9858,N_7665,N_7932);
nand U9859 (N_9859,N_8716,N_8384);
nor U9860 (N_9860,N_7615,N_7800);
xor U9861 (N_9861,N_7541,N_8163);
and U9862 (N_9862,N_8143,N_8186);
nor U9863 (N_9863,N_8030,N_8483);
nor U9864 (N_9864,N_7688,N_7848);
and U9865 (N_9865,N_8201,N_7551);
nand U9866 (N_9866,N_8393,N_7812);
and U9867 (N_9867,N_8663,N_7608);
or U9868 (N_9868,N_8506,N_8687);
and U9869 (N_9869,N_8103,N_8687);
and U9870 (N_9870,N_7892,N_7538);
nor U9871 (N_9871,N_8853,N_8108);
nor U9872 (N_9872,N_8744,N_8303);
and U9873 (N_9873,N_7814,N_7581);
or U9874 (N_9874,N_8610,N_7943);
xor U9875 (N_9875,N_8226,N_8742);
nor U9876 (N_9876,N_7862,N_8009);
xor U9877 (N_9877,N_8481,N_8188);
nand U9878 (N_9878,N_8735,N_8149);
nand U9879 (N_9879,N_7564,N_8127);
nor U9880 (N_9880,N_8657,N_8967);
nor U9881 (N_9881,N_7633,N_7650);
or U9882 (N_9882,N_7513,N_8777);
nand U9883 (N_9883,N_7798,N_7606);
nand U9884 (N_9884,N_8424,N_8684);
nand U9885 (N_9885,N_7810,N_7534);
nor U9886 (N_9886,N_8358,N_8768);
nand U9887 (N_9887,N_8359,N_8234);
or U9888 (N_9888,N_8474,N_8020);
xnor U9889 (N_9889,N_7813,N_8072);
nand U9890 (N_9890,N_8749,N_7643);
or U9891 (N_9891,N_8702,N_7913);
or U9892 (N_9892,N_8058,N_8010);
and U9893 (N_9893,N_8042,N_8132);
or U9894 (N_9894,N_7764,N_8988);
nand U9895 (N_9895,N_8033,N_8976);
nor U9896 (N_9896,N_7519,N_8177);
nand U9897 (N_9897,N_8535,N_8196);
nand U9898 (N_9898,N_8327,N_8482);
nand U9899 (N_9899,N_7568,N_8239);
nor U9900 (N_9900,N_7650,N_7618);
nand U9901 (N_9901,N_7978,N_8191);
or U9902 (N_9902,N_8129,N_8311);
and U9903 (N_9903,N_8633,N_8494);
and U9904 (N_9904,N_8373,N_8263);
and U9905 (N_9905,N_8731,N_7942);
or U9906 (N_9906,N_8372,N_8699);
and U9907 (N_9907,N_8190,N_8099);
nor U9908 (N_9908,N_8885,N_7851);
or U9909 (N_9909,N_8123,N_7634);
nor U9910 (N_9910,N_7851,N_8082);
or U9911 (N_9911,N_8668,N_7998);
or U9912 (N_9912,N_8860,N_8815);
nor U9913 (N_9913,N_7694,N_8748);
or U9914 (N_9914,N_8190,N_7808);
and U9915 (N_9915,N_8325,N_8373);
or U9916 (N_9916,N_7523,N_8753);
nor U9917 (N_9917,N_8109,N_7783);
or U9918 (N_9918,N_8635,N_8564);
nor U9919 (N_9919,N_7945,N_8650);
or U9920 (N_9920,N_8073,N_8451);
nand U9921 (N_9921,N_8623,N_8797);
and U9922 (N_9922,N_8013,N_8778);
nor U9923 (N_9923,N_8647,N_7846);
xnor U9924 (N_9924,N_8267,N_8614);
xor U9925 (N_9925,N_7964,N_7584);
nor U9926 (N_9926,N_8365,N_8496);
nor U9927 (N_9927,N_7701,N_7963);
or U9928 (N_9928,N_8639,N_7987);
nand U9929 (N_9929,N_8152,N_8324);
or U9930 (N_9930,N_8472,N_8632);
nor U9931 (N_9931,N_7705,N_7506);
nor U9932 (N_9932,N_7502,N_8749);
and U9933 (N_9933,N_7678,N_8680);
nor U9934 (N_9934,N_8909,N_8442);
nand U9935 (N_9935,N_8361,N_8534);
nand U9936 (N_9936,N_7647,N_8311);
and U9937 (N_9937,N_7846,N_8974);
and U9938 (N_9938,N_8609,N_7716);
or U9939 (N_9939,N_8921,N_8394);
nor U9940 (N_9940,N_8632,N_8492);
nand U9941 (N_9941,N_8786,N_7543);
xnor U9942 (N_9942,N_7979,N_7869);
nand U9943 (N_9943,N_8719,N_8187);
nand U9944 (N_9944,N_7955,N_8680);
or U9945 (N_9945,N_8683,N_7557);
or U9946 (N_9946,N_8179,N_7596);
or U9947 (N_9947,N_8842,N_8136);
or U9948 (N_9948,N_8828,N_8691);
or U9949 (N_9949,N_8900,N_8951);
nand U9950 (N_9950,N_8166,N_8007);
nor U9951 (N_9951,N_7940,N_8596);
nor U9952 (N_9952,N_7734,N_7873);
nand U9953 (N_9953,N_7536,N_7848);
or U9954 (N_9954,N_8874,N_7924);
nor U9955 (N_9955,N_8415,N_7834);
nand U9956 (N_9956,N_7797,N_8497);
or U9957 (N_9957,N_7981,N_8312);
and U9958 (N_9958,N_7907,N_8815);
and U9959 (N_9959,N_8164,N_8100);
and U9960 (N_9960,N_7566,N_8026);
nand U9961 (N_9961,N_7989,N_7659);
nand U9962 (N_9962,N_8473,N_8103);
and U9963 (N_9963,N_7791,N_7597);
and U9964 (N_9964,N_8121,N_7795);
and U9965 (N_9965,N_8091,N_7947);
xnor U9966 (N_9966,N_8546,N_8574);
xor U9967 (N_9967,N_7936,N_8138);
and U9968 (N_9968,N_8375,N_8148);
nor U9969 (N_9969,N_8916,N_8663);
nor U9970 (N_9970,N_8734,N_8884);
xor U9971 (N_9971,N_8527,N_7501);
nor U9972 (N_9972,N_8084,N_8812);
xnor U9973 (N_9973,N_8677,N_8430);
xnor U9974 (N_9974,N_8989,N_7604);
and U9975 (N_9975,N_8203,N_8966);
nor U9976 (N_9976,N_8108,N_8113);
nand U9977 (N_9977,N_7895,N_8609);
or U9978 (N_9978,N_8245,N_8702);
and U9979 (N_9979,N_8784,N_8130);
nor U9980 (N_9980,N_8193,N_8043);
or U9981 (N_9981,N_8013,N_8927);
or U9982 (N_9982,N_8054,N_8601);
or U9983 (N_9983,N_8769,N_7683);
nand U9984 (N_9984,N_8334,N_8402);
nor U9985 (N_9985,N_7894,N_8158);
nand U9986 (N_9986,N_8063,N_8606);
and U9987 (N_9987,N_8519,N_8406);
nand U9988 (N_9988,N_7851,N_7750);
or U9989 (N_9989,N_8802,N_7935);
nor U9990 (N_9990,N_7650,N_8587);
nor U9991 (N_9991,N_8202,N_7757);
nand U9992 (N_9992,N_8853,N_8044);
or U9993 (N_9993,N_8998,N_8895);
nand U9994 (N_9994,N_8292,N_8077);
or U9995 (N_9995,N_8449,N_7719);
and U9996 (N_9996,N_8449,N_8900);
or U9997 (N_9997,N_8626,N_8435);
nor U9998 (N_9998,N_8448,N_8737);
or U9999 (N_9999,N_8197,N_8935);
nor U10000 (N_10000,N_8108,N_8573);
and U10001 (N_10001,N_8583,N_8784);
nor U10002 (N_10002,N_8227,N_8311);
or U10003 (N_10003,N_8996,N_8920);
and U10004 (N_10004,N_8617,N_8058);
nand U10005 (N_10005,N_8332,N_7767);
nand U10006 (N_10006,N_8687,N_8429);
nor U10007 (N_10007,N_7873,N_8174);
or U10008 (N_10008,N_7706,N_8538);
nor U10009 (N_10009,N_8749,N_8922);
and U10010 (N_10010,N_7998,N_8431);
or U10011 (N_10011,N_8135,N_8567);
and U10012 (N_10012,N_8453,N_8965);
or U10013 (N_10013,N_8768,N_8668);
and U10014 (N_10014,N_7781,N_7883);
nand U10015 (N_10015,N_8452,N_8381);
and U10016 (N_10016,N_8013,N_8035);
nand U10017 (N_10017,N_8469,N_8071);
nand U10018 (N_10018,N_8109,N_8713);
and U10019 (N_10019,N_8420,N_8182);
and U10020 (N_10020,N_7671,N_7729);
and U10021 (N_10021,N_8335,N_8904);
nor U10022 (N_10022,N_8691,N_8998);
or U10023 (N_10023,N_8931,N_8519);
or U10024 (N_10024,N_8719,N_8592);
or U10025 (N_10025,N_7879,N_7963);
nand U10026 (N_10026,N_7616,N_7569);
or U10027 (N_10027,N_8146,N_8956);
nand U10028 (N_10028,N_7543,N_8570);
and U10029 (N_10029,N_8223,N_8605);
nand U10030 (N_10030,N_7538,N_8361);
nand U10031 (N_10031,N_8389,N_8931);
or U10032 (N_10032,N_7985,N_8817);
nor U10033 (N_10033,N_8370,N_7927);
and U10034 (N_10034,N_7762,N_8993);
or U10035 (N_10035,N_8120,N_8240);
xnor U10036 (N_10036,N_7547,N_7949);
nor U10037 (N_10037,N_8141,N_8553);
or U10038 (N_10038,N_8032,N_8889);
nor U10039 (N_10039,N_8181,N_7834);
nand U10040 (N_10040,N_7803,N_8096);
nor U10041 (N_10041,N_8676,N_8333);
nand U10042 (N_10042,N_8868,N_8398);
or U10043 (N_10043,N_8069,N_8671);
or U10044 (N_10044,N_8641,N_8785);
and U10045 (N_10045,N_8376,N_7609);
nor U10046 (N_10046,N_8913,N_8749);
nand U10047 (N_10047,N_8492,N_8337);
nor U10048 (N_10048,N_8979,N_8009);
or U10049 (N_10049,N_7616,N_8622);
and U10050 (N_10050,N_8784,N_7779);
or U10051 (N_10051,N_8880,N_8030);
or U10052 (N_10052,N_8736,N_7966);
nor U10053 (N_10053,N_8288,N_8744);
nor U10054 (N_10054,N_8478,N_7504);
nand U10055 (N_10055,N_8305,N_8320);
nor U10056 (N_10056,N_8146,N_8070);
and U10057 (N_10057,N_8539,N_8726);
or U10058 (N_10058,N_8105,N_8167);
nand U10059 (N_10059,N_8763,N_8759);
or U10060 (N_10060,N_7820,N_8232);
xor U10061 (N_10061,N_8098,N_7749);
or U10062 (N_10062,N_8391,N_8819);
nor U10063 (N_10063,N_8587,N_7779);
and U10064 (N_10064,N_7857,N_7827);
nand U10065 (N_10065,N_8450,N_8425);
or U10066 (N_10066,N_8071,N_7524);
and U10067 (N_10067,N_7563,N_7582);
and U10068 (N_10068,N_7840,N_7636);
nand U10069 (N_10069,N_8181,N_8062);
nor U10070 (N_10070,N_7569,N_7628);
or U10071 (N_10071,N_8580,N_7970);
xnor U10072 (N_10072,N_8316,N_7601);
and U10073 (N_10073,N_8028,N_8341);
nor U10074 (N_10074,N_8953,N_8226);
and U10075 (N_10075,N_8208,N_8700);
nor U10076 (N_10076,N_7930,N_8610);
nand U10077 (N_10077,N_8540,N_8779);
nor U10078 (N_10078,N_8004,N_8771);
nor U10079 (N_10079,N_7798,N_8156);
or U10080 (N_10080,N_7594,N_8241);
nand U10081 (N_10081,N_8117,N_8469);
and U10082 (N_10082,N_8831,N_8067);
nor U10083 (N_10083,N_7757,N_8142);
and U10084 (N_10084,N_8870,N_8599);
nand U10085 (N_10085,N_7810,N_7948);
or U10086 (N_10086,N_8704,N_8367);
nor U10087 (N_10087,N_7657,N_8327);
and U10088 (N_10088,N_8493,N_8264);
nor U10089 (N_10089,N_7635,N_8969);
nand U10090 (N_10090,N_8515,N_8265);
nor U10091 (N_10091,N_8942,N_8410);
and U10092 (N_10092,N_8286,N_8752);
and U10093 (N_10093,N_7569,N_7947);
or U10094 (N_10094,N_7523,N_8642);
nor U10095 (N_10095,N_8560,N_8026);
nand U10096 (N_10096,N_8666,N_7998);
nand U10097 (N_10097,N_8261,N_7580);
or U10098 (N_10098,N_8881,N_8431);
nor U10099 (N_10099,N_8968,N_8999);
nand U10100 (N_10100,N_8220,N_8721);
or U10101 (N_10101,N_7956,N_8137);
and U10102 (N_10102,N_8677,N_8964);
nand U10103 (N_10103,N_8524,N_8502);
and U10104 (N_10104,N_7503,N_8222);
nand U10105 (N_10105,N_8549,N_7695);
nor U10106 (N_10106,N_8123,N_7753);
nor U10107 (N_10107,N_8703,N_8982);
nor U10108 (N_10108,N_8479,N_8666);
nor U10109 (N_10109,N_7712,N_8030);
and U10110 (N_10110,N_8528,N_8746);
or U10111 (N_10111,N_7524,N_8444);
or U10112 (N_10112,N_8827,N_8006);
or U10113 (N_10113,N_8405,N_8856);
xor U10114 (N_10114,N_8829,N_7788);
nand U10115 (N_10115,N_8920,N_8298);
and U10116 (N_10116,N_7643,N_8792);
and U10117 (N_10117,N_8850,N_7556);
and U10118 (N_10118,N_7999,N_8490);
or U10119 (N_10119,N_8712,N_8656);
nor U10120 (N_10120,N_7626,N_8355);
nor U10121 (N_10121,N_8155,N_8936);
nor U10122 (N_10122,N_8907,N_7958);
or U10123 (N_10123,N_8257,N_8140);
or U10124 (N_10124,N_8358,N_7629);
xor U10125 (N_10125,N_8167,N_8366);
and U10126 (N_10126,N_8807,N_8659);
nand U10127 (N_10127,N_8644,N_8910);
nor U10128 (N_10128,N_8450,N_8476);
and U10129 (N_10129,N_7533,N_8240);
nand U10130 (N_10130,N_8108,N_7697);
nor U10131 (N_10131,N_8648,N_8136);
and U10132 (N_10132,N_8658,N_8500);
nor U10133 (N_10133,N_7642,N_8694);
nor U10134 (N_10134,N_8988,N_8674);
nor U10135 (N_10135,N_8417,N_8730);
and U10136 (N_10136,N_7798,N_8253);
xnor U10137 (N_10137,N_8253,N_7631);
nor U10138 (N_10138,N_8374,N_8963);
or U10139 (N_10139,N_8020,N_7840);
or U10140 (N_10140,N_8710,N_8935);
xnor U10141 (N_10141,N_8567,N_8941);
xor U10142 (N_10142,N_8593,N_8084);
xnor U10143 (N_10143,N_8320,N_7684);
or U10144 (N_10144,N_8319,N_8972);
nor U10145 (N_10145,N_8087,N_7684);
xnor U10146 (N_10146,N_8840,N_8037);
and U10147 (N_10147,N_7880,N_8491);
or U10148 (N_10148,N_8462,N_8728);
nor U10149 (N_10149,N_8947,N_8695);
or U10150 (N_10150,N_8812,N_7919);
nand U10151 (N_10151,N_8435,N_8340);
or U10152 (N_10152,N_8221,N_8729);
nand U10153 (N_10153,N_8847,N_8682);
nor U10154 (N_10154,N_7955,N_8654);
and U10155 (N_10155,N_7696,N_8895);
or U10156 (N_10156,N_7870,N_8257);
or U10157 (N_10157,N_7830,N_8775);
nor U10158 (N_10158,N_7891,N_8175);
or U10159 (N_10159,N_8571,N_7706);
nor U10160 (N_10160,N_8689,N_8711);
or U10161 (N_10161,N_8101,N_8127);
nand U10162 (N_10162,N_7555,N_8388);
xnor U10163 (N_10163,N_7900,N_8477);
nor U10164 (N_10164,N_8243,N_8620);
nand U10165 (N_10165,N_8717,N_7644);
nand U10166 (N_10166,N_8997,N_8816);
or U10167 (N_10167,N_8254,N_7560);
or U10168 (N_10168,N_7758,N_7827);
and U10169 (N_10169,N_7671,N_8404);
nand U10170 (N_10170,N_7565,N_7764);
or U10171 (N_10171,N_8118,N_8235);
nand U10172 (N_10172,N_8547,N_7704);
nor U10173 (N_10173,N_8946,N_8927);
nand U10174 (N_10174,N_8064,N_7974);
xnor U10175 (N_10175,N_8399,N_8314);
xnor U10176 (N_10176,N_7595,N_7874);
nor U10177 (N_10177,N_7842,N_7703);
or U10178 (N_10178,N_8737,N_8862);
or U10179 (N_10179,N_8385,N_7949);
nor U10180 (N_10180,N_8532,N_8497);
and U10181 (N_10181,N_7515,N_7757);
nand U10182 (N_10182,N_7642,N_8021);
nor U10183 (N_10183,N_7557,N_8175);
nor U10184 (N_10184,N_7645,N_8568);
or U10185 (N_10185,N_8997,N_8346);
nor U10186 (N_10186,N_7528,N_8009);
nor U10187 (N_10187,N_7819,N_8339);
or U10188 (N_10188,N_8052,N_8259);
xnor U10189 (N_10189,N_8030,N_8318);
xnor U10190 (N_10190,N_8976,N_8344);
nor U10191 (N_10191,N_7638,N_7782);
and U10192 (N_10192,N_8159,N_8837);
and U10193 (N_10193,N_7518,N_8363);
or U10194 (N_10194,N_8952,N_7940);
and U10195 (N_10195,N_8297,N_8467);
xnor U10196 (N_10196,N_8789,N_8805);
or U10197 (N_10197,N_8680,N_8581);
xor U10198 (N_10198,N_8088,N_8288);
nand U10199 (N_10199,N_8867,N_8022);
xor U10200 (N_10200,N_8727,N_7508);
nor U10201 (N_10201,N_8583,N_8865);
nor U10202 (N_10202,N_7849,N_8996);
and U10203 (N_10203,N_7612,N_8956);
and U10204 (N_10204,N_7711,N_8615);
nand U10205 (N_10205,N_8716,N_8435);
or U10206 (N_10206,N_7928,N_8357);
nand U10207 (N_10207,N_7651,N_7650);
xnor U10208 (N_10208,N_8525,N_8413);
nor U10209 (N_10209,N_7916,N_8620);
and U10210 (N_10210,N_8593,N_7987);
xnor U10211 (N_10211,N_8799,N_7726);
xnor U10212 (N_10212,N_8627,N_8891);
and U10213 (N_10213,N_8269,N_8509);
nor U10214 (N_10214,N_7571,N_7906);
nand U10215 (N_10215,N_8577,N_8158);
nor U10216 (N_10216,N_7687,N_7563);
or U10217 (N_10217,N_7838,N_8235);
nand U10218 (N_10218,N_8667,N_8358);
nand U10219 (N_10219,N_8070,N_8952);
and U10220 (N_10220,N_7871,N_8347);
and U10221 (N_10221,N_8427,N_8780);
nand U10222 (N_10222,N_7621,N_8537);
nor U10223 (N_10223,N_7599,N_8311);
and U10224 (N_10224,N_8712,N_8819);
nand U10225 (N_10225,N_7744,N_8408);
and U10226 (N_10226,N_8825,N_8599);
and U10227 (N_10227,N_8575,N_8194);
or U10228 (N_10228,N_8503,N_8230);
or U10229 (N_10229,N_8872,N_7800);
and U10230 (N_10230,N_8759,N_8943);
or U10231 (N_10231,N_8734,N_8688);
or U10232 (N_10232,N_7844,N_8926);
or U10233 (N_10233,N_7537,N_7904);
xor U10234 (N_10234,N_8151,N_7934);
nand U10235 (N_10235,N_8280,N_8403);
and U10236 (N_10236,N_8653,N_8261);
and U10237 (N_10237,N_8673,N_8554);
nor U10238 (N_10238,N_8582,N_8050);
or U10239 (N_10239,N_8026,N_8153);
xor U10240 (N_10240,N_8623,N_8629);
nand U10241 (N_10241,N_8383,N_8783);
nand U10242 (N_10242,N_8396,N_8198);
nor U10243 (N_10243,N_8366,N_8605);
or U10244 (N_10244,N_8716,N_8076);
nor U10245 (N_10245,N_8095,N_8815);
nor U10246 (N_10246,N_7810,N_8141);
nand U10247 (N_10247,N_8365,N_8117);
or U10248 (N_10248,N_8925,N_7974);
or U10249 (N_10249,N_7785,N_8488);
or U10250 (N_10250,N_7681,N_7655);
nor U10251 (N_10251,N_8455,N_8194);
nor U10252 (N_10252,N_7900,N_8337);
and U10253 (N_10253,N_7863,N_8125);
and U10254 (N_10254,N_7918,N_7649);
or U10255 (N_10255,N_8196,N_8989);
nor U10256 (N_10256,N_7991,N_8363);
nor U10257 (N_10257,N_8096,N_7966);
nor U10258 (N_10258,N_8179,N_8336);
nand U10259 (N_10259,N_8893,N_7810);
xor U10260 (N_10260,N_8509,N_7674);
xor U10261 (N_10261,N_7848,N_8115);
and U10262 (N_10262,N_8360,N_8150);
or U10263 (N_10263,N_8645,N_7688);
or U10264 (N_10264,N_7987,N_8531);
nor U10265 (N_10265,N_8863,N_7917);
xnor U10266 (N_10266,N_8745,N_7553);
and U10267 (N_10267,N_7589,N_8513);
nand U10268 (N_10268,N_8602,N_7975);
nand U10269 (N_10269,N_8345,N_7771);
or U10270 (N_10270,N_7838,N_8018);
and U10271 (N_10271,N_8499,N_8948);
and U10272 (N_10272,N_7671,N_7886);
xor U10273 (N_10273,N_8318,N_8249);
or U10274 (N_10274,N_7614,N_8879);
and U10275 (N_10275,N_8229,N_8271);
and U10276 (N_10276,N_8382,N_8736);
xor U10277 (N_10277,N_8978,N_8877);
or U10278 (N_10278,N_7939,N_8046);
nor U10279 (N_10279,N_8403,N_8812);
nor U10280 (N_10280,N_8092,N_8592);
nor U10281 (N_10281,N_8721,N_8920);
or U10282 (N_10282,N_8269,N_7993);
xor U10283 (N_10283,N_8676,N_7829);
nand U10284 (N_10284,N_8697,N_8375);
and U10285 (N_10285,N_8010,N_8121);
nand U10286 (N_10286,N_8762,N_8697);
or U10287 (N_10287,N_8094,N_7819);
nand U10288 (N_10288,N_8766,N_8753);
or U10289 (N_10289,N_8253,N_7771);
nand U10290 (N_10290,N_7557,N_8874);
and U10291 (N_10291,N_8450,N_8108);
or U10292 (N_10292,N_8717,N_8364);
nor U10293 (N_10293,N_8068,N_8540);
xnor U10294 (N_10294,N_8848,N_8650);
or U10295 (N_10295,N_7575,N_8855);
nand U10296 (N_10296,N_8628,N_8576);
xnor U10297 (N_10297,N_8169,N_8795);
and U10298 (N_10298,N_8240,N_8713);
nand U10299 (N_10299,N_7595,N_7714);
nor U10300 (N_10300,N_8180,N_7692);
nor U10301 (N_10301,N_8724,N_8739);
and U10302 (N_10302,N_8025,N_8254);
or U10303 (N_10303,N_7933,N_8521);
nand U10304 (N_10304,N_8645,N_8963);
and U10305 (N_10305,N_7654,N_8869);
or U10306 (N_10306,N_7897,N_8382);
and U10307 (N_10307,N_8395,N_8391);
or U10308 (N_10308,N_8575,N_8161);
nor U10309 (N_10309,N_8285,N_7810);
and U10310 (N_10310,N_8055,N_8697);
or U10311 (N_10311,N_8283,N_8731);
or U10312 (N_10312,N_8047,N_7889);
nand U10313 (N_10313,N_8235,N_8485);
and U10314 (N_10314,N_7874,N_8295);
nor U10315 (N_10315,N_7528,N_8284);
and U10316 (N_10316,N_7806,N_8716);
and U10317 (N_10317,N_8760,N_8342);
and U10318 (N_10318,N_8042,N_7952);
nor U10319 (N_10319,N_8278,N_8184);
and U10320 (N_10320,N_8851,N_8751);
nor U10321 (N_10321,N_8285,N_8039);
or U10322 (N_10322,N_7774,N_7962);
nor U10323 (N_10323,N_8027,N_7793);
xor U10324 (N_10324,N_8872,N_8068);
and U10325 (N_10325,N_8840,N_7733);
nand U10326 (N_10326,N_7615,N_8840);
and U10327 (N_10327,N_8045,N_8571);
and U10328 (N_10328,N_8204,N_7553);
or U10329 (N_10329,N_7861,N_8537);
nor U10330 (N_10330,N_8772,N_7821);
and U10331 (N_10331,N_8927,N_7753);
or U10332 (N_10332,N_8065,N_8586);
nor U10333 (N_10333,N_8207,N_7956);
nor U10334 (N_10334,N_7829,N_7717);
and U10335 (N_10335,N_8507,N_8667);
nor U10336 (N_10336,N_8123,N_8192);
nand U10337 (N_10337,N_7839,N_7628);
nand U10338 (N_10338,N_7853,N_8282);
nor U10339 (N_10339,N_8842,N_7653);
nand U10340 (N_10340,N_7526,N_7549);
nor U10341 (N_10341,N_7580,N_7681);
and U10342 (N_10342,N_7893,N_7732);
xor U10343 (N_10343,N_7530,N_7541);
nor U10344 (N_10344,N_7855,N_8114);
or U10345 (N_10345,N_7959,N_7693);
and U10346 (N_10346,N_7999,N_8376);
and U10347 (N_10347,N_8185,N_8554);
nor U10348 (N_10348,N_8265,N_8316);
nand U10349 (N_10349,N_8917,N_8497);
nand U10350 (N_10350,N_7983,N_7686);
and U10351 (N_10351,N_7623,N_8149);
nand U10352 (N_10352,N_8477,N_8721);
or U10353 (N_10353,N_8876,N_8049);
or U10354 (N_10354,N_8868,N_8128);
and U10355 (N_10355,N_8255,N_7640);
nand U10356 (N_10356,N_8654,N_8588);
nor U10357 (N_10357,N_8501,N_8351);
and U10358 (N_10358,N_8972,N_7605);
nand U10359 (N_10359,N_7933,N_8850);
and U10360 (N_10360,N_7699,N_7662);
nor U10361 (N_10361,N_7947,N_8023);
or U10362 (N_10362,N_8629,N_8351);
nand U10363 (N_10363,N_8708,N_8460);
and U10364 (N_10364,N_7971,N_8617);
nand U10365 (N_10365,N_7501,N_8975);
xor U10366 (N_10366,N_8575,N_7603);
nand U10367 (N_10367,N_8185,N_8214);
nor U10368 (N_10368,N_8415,N_7981);
or U10369 (N_10369,N_8622,N_8712);
or U10370 (N_10370,N_8729,N_8356);
nand U10371 (N_10371,N_8365,N_7783);
or U10372 (N_10372,N_8882,N_7694);
or U10373 (N_10373,N_8326,N_7605);
or U10374 (N_10374,N_8038,N_7514);
or U10375 (N_10375,N_8520,N_8835);
nor U10376 (N_10376,N_8360,N_8154);
xor U10377 (N_10377,N_8185,N_8990);
or U10378 (N_10378,N_7543,N_8683);
and U10379 (N_10379,N_8229,N_8237);
or U10380 (N_10380,N_8904,N_8275);
nand U10381 (N_10381,N_8489,N_7523);
nor U10382 (N_10382,N_8399,N_8318);
nor U10383 (N_10383,N_8525,N_7531);
nor U10384 (N_10384,N_7589,N_8062);
nand U10385 (N_10385,N_7646,N_7915);
or U10386 (N_10386,N_7767,N_8104);
nand U10387 (N_10387,N_7857,N_8879);
and U10388 (N_10388,N_8081,N_8735);
or U10389 (N_10389,N_7959,N_7731);
nand U10390 (N_10390,N_8879,N_8967);
nor U10391 (N_10391,N_7650,N_8681);
and U10392 (N_10392,N_8685,N_8360);
xor U10393 (N_10393,N_7844,N_8897);
and U10394 (N_10394,N_8746,N_8686);
nand U10395 (N_10395,N_7662,N_7848);
and U10396 (N_10396,N_8476,N_8687);
xnor U10397 (N_10397,N_8030,N_8981);
and U10398 (N_10398,N_7501,N_7563);
and U10399 (N_10399,N_7651,N_7547);
nor U10400 (N_10400,N_8444,N_8788);
and U10401 (N_10401,N_7816,N_8231);
or U10402 (N_10402,N_7704,N_8678);
or U10403 (N_10403,N_7971,N_8169);
xor U10404 (N_10404,N_8133,N_8758);
nor U10405 (N_10405,N_8448,N_8717);
nor U10406 (N_10406,N_7708,N_8236);
or U10407 (N_10407,N_7769,N_8564);
or U10408 (N_10408,N_7872,N_8080);
nor U10409 (N_10409,N_8393,N_8071);
or U10410 (N_10410,N_8700,N_7757);
and U10411 (N_10411,N_7888,N_8838);
and U10412 (N_10412,N_7592,N_8571);
nor U10413 (N_10413,N_8574,N_8173);
or U10414 (N_10414,N_7879,N_7689);
nand U10415 (N_10415,N_8173,N_7811);
or U10416 (N_10416,N_8697,N_8172);
nor U10417 (N_10417,N_8723,N_8696);
and U10418 (N_10418,N_7956,N_7768);
nor U10419 (N_10419,N_8912,N_8596);
nand U10420 (N_10420,N_8602,N_8419);
nand U10421 (N_10421,N_7519,N_7715);
or U10422 (N_10422,N_8575,N_8938);
nor U10423 (N_10423,N_8592,N_8951);
nand U10424 (N_10424,N_7929,N_8064);
or U10425 (N_10425,N_8724,N_8776);
nand U10426 (N_10426,N_7824,N_8010);
and U10427 (N_10427,N_8786,N_7794);
and U10428 (N_10428,N_7886,N_7935);
or U10429 (N_10429,N_7778,N_8329);
xor U10430 (N_10430,N_8523,N_8195);
nor U10431 (N_10431,N_8443,N_8927);
nor U10432 (N_10432,N_7574,N_7612);
nand U10433 (N_10433,N_8658,N_7714);
and U10434 (N_10434,N_8042,N_8059);
nor U10435 (N_10435,N_7836,N_8134);
nand U10436 (N_10436,N_8710,N_7857);
nand U10437 (N_10437,N_8390,N_8486);
and U10438 (N_10438,N_7661,N_8653);
and U10439 (N_10439,N_8293,N_8395);
nor U10440 (N_10440,N_8707,N_8367);
xnor U10441 (N_10441,N_8969,N_7505);
nor U10442 (N_10442,N_8092,N_7600);
xor U10443 (N_10443,N_8091,N_8432);
nor U10444 (N_10444,N_8447,N_8416);
and U10445 (N_10445,N_8999,N_7545);
nor U10446 (N_10446,N_7613,N_7958);
or U10447 (N_10447,N_7518,N_7909);
or U10448 (N_10448,N_8542,N_8805);
nand U10449 (N_10449,N_7958,N_8452);
nor U10450 (N_10450,N_8234,N_8760);
nand U10451 (N_10451,N_8865,N_8722);
nand U10452 (N_10452,N_7573,N_8860);
nand U10453 (N_10453,N_8417,N_8491);
nor U10454 (N_10454,N_7884,N_7858);
or U10455 (N_10455,N_7873,N_7831);
nand U10456 (N_10456,N_8784,N_7909);
nor U10457 (N_10457,N_7850,N_8870);
nand U10458 (N_10458,N_7516,N_8081);
and U10459 (N_10459,N_8237,N_8034);
xnor U10460 (N_10460,N_8721,N_7944);
xor U10461 (N_10461,N_8214,N_8493);
xnor U10462 (N_10462,N_8752,N_7837);
or U10463 (N_10463,N_7884,N_8141);
nor U10464 (N_10464,N_7776,N_8293);
nand U10465 (N_10465,N_8742,N_8608);
nand U10466 (N_10466,N_7772,N_7849);
and U10467 (N_10467,N_7740,N_7602);
nand U10468 (N_10468,N_7614,N_7576);
nor U10469 (N_10469,N_8521,N_8730);
or U10470 (N_10470,N_7685,N_8640);
nand U10471 (N_10471,N_7566,N_8633);
nand U10472 (N_10472,N_7811,N_8899);
and U10473 (N_10473,N_8650,N_8540);
or U10474 (N_10474,N_8200,N_7913);
nand U10475 (N_10475,N_8799,N_8790);
xor U10476 (N_10476,N_8956,N_7800);
and U10477 (N_10477,N_8452,N_8063);
nand U10478 (N_10478,N_7932,N_7595);
and U10479 (N_10479,N_8199,N_7794);
nor U10480 (N_10480,N_8244,N_8904);
or U10481 (N_10481,N_7722,N_8119);
nor U10482 (N_10482,N_8373,N_8593);
and U10483 (N_10483,N_8865,N_8920);
and U10484 (N_10484,N_7718,N_8999);
xnor U10485 (N_10485,N_8278,N_8759);
or U10486 (N_10486,N_7854,N_8930);
and U10487 (N_10487,N_7606,N_8890);
or U10488 (N_10488,N_8006,N_7630);
xor U10489 (N_10489,N_8826,N_8846);
nand U10490 (N_10490,N_8140,N_8330);
nor U10491 (N_10491,N_7537,N_8190);
xor U10492 (N_10492,N_7916,N_7552);
nand U10493 (N_10493,N_7632,N_7645);
nor U10494 (N_10494,N_7813,N_8724);
nor U10495 (N_10495,N_8189,N_8629);
or U10496 (N_10496,N_7594,N_8876);
or U10497 (N_10497,N_8585,N_8728);
nand U10498 (N_10498,N_8524,N_7933);
nand U10499 (N_10499,N_8413,N_8151);
or U10500 (N_10500,N_9066,N_10451);
nor U10501 (N_10501,N_9991,N_10061);
xor U10502 (N_10502,N_9732,N_10133);
or U10503 (N_10503,N_10317,N_9765);
and U10504 (N_10504,N_9290,N_10208);
or U10505 (N_10505,N_9615,N_9703);
nor U10506 (N_10506,N_9087,N_9639);
nor U10507 (N_10507,N_9630,N_9638);
and U10508 (N_10508,N_9436,N_9936);
xor U10509 (N_10509,N_9728,N_10494);
nor U10510 (N_10510,N_9879,N_9642);
nor U10511 (N_10511,N_9123,N_10254);
and U10512 (N_10512,N_10441,N_9182);
nor U10513 (N_10513,N_10038,N_10427);
nor U10514 (N_10514,N_9247,N_9328);
and U10515 (N_10515,N_9627,N_9214);
or U10516 (N_10516,N_9572,N_9095);
nor U10517 (N_10517,N_10414,N_9990);
nor U10518 (N_10518,N_10306,N_9121);
xnor U10519 (N_10519,N_9604,N_9992);
nor U10520 (N_10520,N_10042,N_9553);
and U10521 (N_10521,N_10300,N_9145);
or U10522 (N_10522,N_9249,N_10380);
and U10523 (N_10523,N_9804,N_9813);
and U10524 (N_10524,N_10394,N_9499);
nand U10525 (N_10525,N_10333,N_9834);
nor U10526 (N_10526,N_9281,N_9006);
nand U10527 (N_10527,N_9403,N_10008);
or U10528 (N_10528,N_9124,N_9125);
nand U10529 (N_10529,N_9374,N_9002);
xor U10530 (N_10530,N_9028,N_9402);
nand U10531 (N_10531,N_10175,N_9306);
and U10532 (N_10532,N_9942,N_9746);
nor U10533 (N_10533,N_9021,N_9581);
nor U10534 (N_10534,N_10288,N_9138);
and U10535 (N_10535,N_9391,N_9201);
nand U10536 (N_10536,N_9322,N_9544);
nand U10537 (N_10537,N_10043,N_10097);
and U10538 (N_10538,N_9756,N_9856);
and U10539 (N_10539,N_10383,N_9761);
nor U10540 (N_10540,N_9419,N_9174);
or U10541 (N_10541,N_9954,N_10379);
or U10542 (N_10542,N_9415,N_9038);
and U10543 (N_10543,N_10396,N_9375);
nand U10544 (N_10544,N_9131,N_9845);
nor U10545 (N_10545,N_9350,N_9571);
or U10546 (N_10546,N_9452,N_10103);
or U10547 (N_10547,N_9672,N_9521);
or U10548 (N_10548,N_10140,N_9458);
nand U10549 (N_10549,N_9790,N_10395);
or U10550 (N_10550,N_9674,N_10011);
and U10551 (N_10551,N_10471,N_9248);
or U10552 (N_10552,N_9673,N_9871);
nand U10553 (N_10553,N_9805,N_10044);
and U10554 (N_10554,N_10204,N_10415);
nand U10555 (N_10555,N_9044,N_9163);
nand U10556 (N_10556,N_10195,N_9475);
or U10557 (N_10557,N_10192,N_10174);
and U10558 (N_10558,N_9963,N_9652);
nor U10559 (N_10559,N_10230,N_9139);
and U10560 (N_10560,N_10100,N_9166);
or U10561 (N_10561,N_9893,N_9218);
nor U10562 (N_10562,N_9558,N_9720);
nand U10563 (N_10563,N_9680,N_9435);
xnor U10564 (N_10564,N_9294,N_9037);
xor U10565 (N_10565,N_10385,N_9794);
nand U10566 (N_10566,N_9657,N_9046);
or U10567 (N_10567,N_9230,N_9598);
and U10568 (N_10568,N_9244,N_9269);
and U10569 (N_10569,N_9068,N_10036);
and U10570 (N_10570,N_10473,N_9196);
or U10571 (N_10571,N_10191,N_9461);
nor U10572 (N_10572,N_9377,N_9821);
or U10573 (N_10573,N_10322,N_9513);
nor U10574 (N_10574,N_10054,N_10163);
nand U10575 (N_10575,N_9624,N_10002);
xor U10576 (N_10576,N_9355,N_10072);
xor U10577 (N_10577,N_9008,N_9841);
and U10578 (N_10578,N_9034,N_10299);
nand U10579 (N_10579,N_10261,N_9707);
and U10580 (N_10580,N_9913,N_9874);
and U10581 (N_10581,N_9787,N_9986);
or U10582 (N_10582,N_9384,N_9326);
nor U10583 (N_10583,N_9187,N_9042);
and U10584 (N_10584,N_9511,N_9001);
nand U10585 (N_10585,N_10423,N_10474);
and U10586 (N_10586,N_9519,N_10210);
and U10587 (N_10587,N_9906,N_9440);
nor U10588 (N_10588,N_10183,N_9227);
nand U10589 (N_10589,N_9449,N_9243);
and U10590 (N_10590,N_9751,N_9752);
and U10591 (N_10591,N_9870,N_9482);
xor U10592 (N_10592,N_10050,N_9955);
and U10593 (N_10593,N_9520,N_10089);
or U10594 (N_10594,N_9601,N_9516);
or U10595 (N_10595,N_9303,N_9261);
and U10596 (N_10596,N_10307,N_9047);
and U10597 (N_10597,N_9378,N_9550);
or U10598 (N_10598,N_9983,N_9147);
and U10599 (N_10599,N_9089,N_9929);
or U10600 (N_10600,N_10200,N_10264);
nand U10601 (N_10601,N_9600,N_10040);
or U10602 (N_10602,N_10284,N_10001);
or U10603 (N_10603,N_10392,N_9305);
and U10604 (N_10604,N_9842,N_9860);
or U10605 (N_10605,N_10095,N_10127);
or U10606 (N_10606,N_9070,N_10013);
nand U10607 (N_10607,N_9867,N_10320);
or U10608 (N_10608,N_9545,N_10374);
or U10609 (N_10609,N_9722,N_9744);
nand U10610 (N_10610,N_9573,N_9013);
nor U10611 (N_10611,N_9775,N_9512);
xnor U10612 (N_10612,N_9921,N_10298);
or U10613 (N_10613,N_9351,N_9721);
or U10614 (N_10614,N_9809,N_10165);
or U10615 (N_10615,N_10170,N_9503);
and U10616 (N_10616,N_9067,N_9768);
nand U10617 (N_10617,N_9058,N_9956);
or U10618 (N_10618,N_10067,N_10367);
nand U10619 (N_10619,N_9644,N_9670);
and U10620 (N_10620,N_10278,N_10139);
nand U10621 (N_10621,N_9240,N_9446);
or U10622 (N_10622,N_10227,N_10371);
and U10623 (N_10623,N_10430,N_9223);
nor U10624 (N_10624,N_9190,N_10289);
xor U10625 (N_10625,N_9122,N_9018);
or U10626 (N_10626,N_10041,N_10128);
or U10627 (N_10627,N_9059,N_9362);
nand U10628 (N_10628,N_9549,N_10022);
nand U10629 (N_10629,N_9372,N_9035);
and U10630 (N_10630,N_10272,N_9233);
nor U10631 (N_10631,N_10481,N_9143);
nand U10632 (N_10632,N_9608,N_9200);
or U10633 (N_10633,N_9743,N_10434);
and U10634 (N_10634,N_9431,N_9160);
or U10635 (N_10635,N_10108,N_9114);
nand U10636 (N_10636,N_9137,N_10418);
nand U10637 (N_10637,N_10166,N_10142);
nand U10638 (N_10638,N_10122,N_9840);
nand U10639 (N_10639,N_9057,N_9537);
and U10640 (N_10640,N_9812,N_9994);
nor U10641 (N_10641,N_9696,N_10478);
xnor U10642 (N_10642,N_9607,N_9335);
nor U10643 (N_10643,N_10487,N_9547);
xnor U10644 (N_10644,N_10292,N_9882);
nand U10645 (N_10645,N_10270,N_10260);
and U10646 (N_10646,N_9525,N_9847);
nand U10647 (N_10647,N_9949,N_9327);
and U10648 (N_10648,N_10068,N_9040);
and U10649 (N_10649,N_9154,N_9857);
or U10650 (N_10650,N_9151,N_9665);
or U10651 (N_10651,N_9896,N_9694);
nand U10652 (N_10652,N_10426,N_10386);
xnor U10653 (N_10653,N_10455,N_9268);
nand U10654 (N_10654,N_10123,N_9141);
and U10655 (N_10655,N_9486,N_9394);
and U10656 (N_10656,N_10151,N_9974);
nor U10657 (N_10657,N_9731,N_9366);
or U10658 (N_10658,N_9967,N_9282);
and U10659 (N_10659,N_9623,N_9155);
nor U10660 (N_10660,N_10156,N_10410);
and U10661 (N_10661,N_9144,N_10063);
nor U10662 (N_10662,N_9039,N_9259);
or U10663 (N_10663,N_9389,N_9915);
nand U10664 (N_10664,N_9510,N_9031);
or U10665 (N_10665,N_10448,N_9060);
nor U10666 (N_10666,N_10257,N_10342);
or U10667 (N_10667,N_9307,N_9146);
and U10668 (N_10668,N_10463,N_9656);
or U10669 (N_10669,N_9472,N_9448);
nand U10670 (N_10670,N_10345,N_10185);
nor U10671 (N_10671,N_10469,N_9023);
or U10672 (N_10672,N_9304,N_9689);
nor U10673 (N_10673,N_9235,N_9245);
nor U10674 (N_10674,N_9169,N_9487);
nand U10675 (N_10675,N_10472,N_9236);
and U10676 (N_10676,N_10433,N_9667);
nor U10677 (N_10677,N_9186,N_9183);
or U10678 (N_10678,N_10492,N_9853);
or U10679 (N_10679,N_10475,N_9276);
nor U10680 (N_10680,N_9800,N_10496);
nand U10681 (N_10681,N_9589,N_9334);
nor U10682 (N_10682,N_9944,N_9602);
and U10683 (N_10683,N_10028,N_9376);
nor U10684 (N_10684,N_9858,N_10483);
xnor U10685 (N_10685,N_9718,N_9302);
xor U10686 (N_10686,N_9171,N_10118);
nand U10687 (N_10687,N_9109,N_9202);
and U10688 (N_10688,N_10154,N_9907);
or U10689 (N_10689,N_9234,N_9381);
nand U10690 (N_10690,N_9273,N_9748);
or U10691 (N_10691,N_9153,N_9692);
or U10692 (N_10692,N_9798,N_10422);
nor U10693 (N_10693,N_9951,N_10450);
nand U10694 (N_10694,N_9285,N_9246);
nand U10695 (N_10695,N_10023,N_10334);
nor U10696 (N_10696,N_9317,N_9099);
or U10697 (N_10697,N_10032,N_9876);
nor U10698 (N_10698,N_9833,N_9816);
or U10699 (N_10699,N_9881,N_9941);
or U10700 (N_10700,N_9112,N_10150);
xor U10701 (N_10701,N_9632,N_9465);
nor U10702 (N_10702,N_10184,N_9479);
or U10703 (N_10703,N_9168,N_9727);
nand U10704 (N_10704,N_10031,N_9167);
xor U10705 (N_10705,N_10027,N_10484);
nand U10706 (N_10706,N_10148,N_10060);
or U10707 (N_10707,N_9074,N_10256);
and U10708 (N_10708,N_9204,N_9613);
nor U10709 (N_10709,N_9725,N_10355);
and U10710 (N_10710,N_10222,N_10255);
nand U10711 (N_10711,N_9651,N_9393);
and U10712 (N_10712,N_9687,N_9705);
and U10713 (N_10713,N_10213,N_10155);
xor U10714 (N_10714,N_9940,N_10235);
nand U10715 (N_10715,N_9184,N_9353);
or U10716 (N_10716,N_9164,N_9451);
and U10717 (N_10717,N_10246,N_9136);
nand U10718 (N_10718,N_9988,N_10413);
nor U10719 (N_10719,N_10194,N_9467);
nand U10720 (N_10720,N_9669,N_9385);
nand U10721 (N_10721,N_10079,N_9769);
and U10722 (N_10722,N_9864,N_10018);
nand U10723 (N_10723,N_9062,N_9129);
or U10724 (N_10724,N_9736,N_9635);
or U10725 (N_10725,N_9219,N_9312);
nor U10726 (N_10726,N_9016,N_9421);
nand U10727 (N_10727,N_9408,N_10078);
and U10728 (N_10728,N_9869,N_10399);
or U10729 (N_10729,N_9178,N_9948);
nor U10730 (N_10730,N_10297,N_9577);
and U10731 (N_10731,N_10188,N_9000);
xnor U10732 (N_10732,N_9661,N_10171);
nor U10733 (N_10733,N_9119,N_9428);
nand U10734 (N_10734,N_10065,N_9814);
and U10735 (N_10735,N_9701,N_9773);
nand U10736 (N_10736,N_9959,N_9026);
nand U10737 (N_10737,N_10326,N_9097);
nand U10738 (N_10738,N_9082,N_10055);
and U10739 (N_10739,N_10069,N_9646);
nor U10740 (N_10740,N_9104,N_9005);
nand U10741 (N_10741,N_9298,N_9270);
and U10742 (N_10742,N_9274,N_9284);
or U10743 (N_10743,N_9556,N_9532);
nand U10744 (N_10744,N_10083,N_9213);
and U10745 (N_10745,N_9785,N_9817);
nand U10746 (N_10746,N_9457,N_10117);
or U10747 (N_10747,N_9085,N_9898);
or U10748 (N_10748,N_10488,N_10304);
and U10749 (N_10749,N_9232,N_9799);
or U10750 (N_10750,N_9390,N_9496);
nor U10751 (N_10751,N_9173,N_10181);
or U10752 (N_10752,N_9872,N_9596);
and U10753 (N_10753,N_10274,N_10335);
and U10754 (N_10754,N_10003,N_9237);
or U10755 (N_10755,N_10231,N_9383);
xnor U10756 (N_10756,N_9760,N_10111);
and U10757 (N_10757,N_9420,N_9517);
or U10758 (N_10758,N_10164,N_10405);
nand U10759 (N_10759,N_9352,N_9917);
and U10760 (N_10760,N_9560,N_10080);
xnor U10761 (N_10761,N_9622,N_10332);
and U10762 (N_10762,N_9172,N_9386);
and U10763 (N_10763,N_9012,N_10015);
and U10764 (N_10764,N_9019,N_9704);
or U10765 (N_10765,N_9260,N_9478);
nor U10766 (N_10766,N_9469,N_9685);
nand U10767 (N_10767,N_10412,N_9837);
nor U10768 (N_10768,N_10263,N_9032);
nor U10769 (N_10769,N_9181,N_10404);
nand U10770 (N_10770,N_9552,N_9413);
or U10771 (N_10771,N_9215,N_9810);
xor U10772 (N_10772,N_10269,N_9682);
and U10773 (N_10773,N_9092,N_9447);
or U10774 (N_10774,N_10301,N_10305);
or U10775 (N_10775,N_10406,N_10341);
or U10776 (N_10776,N_9149,N_10039);
and U10777 (N_10777,N_9111,N_9286);
and U10778 (N_10778,N_9597,N_9781);
and U10779 (N_10779,N_9321,N_10336);
nand U10780 (N_10780,N_10282,N_9830);
nand U10781 (N_10781,N_9797,N_9340);
and U10782 (N_10782,N_9148,N_10358);
nor U10783 (N_10783,N_10313,N_10102);
xor U10784 (N_10784,N_9690,N_9093);
and U10785 (N_10785,N_9877,N_9433);
nor U10786 (N_10786,N_9371,N_9014);
nand U10787 (N_10787,N_9654,N_9636);
xor U10788 (N_10788,N_9029,N_10037);
and U10789 (N_10789,N_10145,N_10338);
nand U10790 (N_10790,N_10279,N_9476);
and U10791 (N_10791,N_10408,N_9369);
or U10792 (N_10792,N_9387,N_9806);
nor U10793 (N_10793,N_9889,N_9464);
nor U10794 (N_10794,N_10081,N_9717);
or U10795 (N_10795,N_9649,N_10271);
nand U10796 (N_10796,N_9256,N_9106);
nand U10797 (N_10797,N_10168,N_10076);
nor U10798 (N_10798,N_10224,N_9128);
nor U10799 (N_10799,N_10024,N_10169);
nor U10800 (N_10800,N_10093,N_10071);
nor U10801 (N_10801,N_9702,N_10053);
or U10802 (N_10802,N_9928,N_10343);
nand U10803 (N_10803,N_10310,N_9481);
nand U10804 (N_10804,N_9116,N_10048);
and U10805 (N_10805,N_10215,N_10131);
nor U10806 (N_10806,N_9699,N_10370);
nand U10807 (N_10807,N_9901,N_9902);
or U10808 (N_10808,N_9922,N_9653);
nand U10809 (N_10809,N_9784,N_9466);
nand U10810 (N_10810,N_9554,N_10092);
or U10811 (N_10811,N_10137,N_9076);
nor U10812 (N_10812,N_9590,N_9414);
or U10813 (N_10813,N_9484,N_10085);
nand U10814 (N_10814,N_10232,N_10357);
nor U10815 (N_10815,N_10363,N_9135);
nor U10816 (N_10816,N_9003,N_9884);
nand U10817 (N_10817,N_10075,N_9619);
nand U10818 (N_10818,N_9659,N_9706);
xor U10819 (N_10819,N_9947,N_10315);
and U10820 (N_10820,N_10115,N_9753);
or U10821 (N_10821,N_9398,N_9418);
and U10822 (N_10822,N_10021,N_9679);
nand U10823 (N_10823,N_10025,N_10107);
and U10824 (N_10824,N_9348,N_9684);
or U10825 (N_10825,N_10203,N_9015);
nor U10826 (N_10826,N_9480,N_10465);
and U10827 (N_10827,N_10331,N_9987);
nor U10828 (N_10828,N_9966,N_9443);
nand U10829 (N_10829,N_9908,N_9337);
nand U10830 (N_10830,N_9497,N_9559);
or U10831 (N_10831,N_10016,N_9495);
and U10832 (N_10832,N_9820,N_10147);
nor U10833 (N_10833,N_10321,N_10311);
and U10834 (N_10834,N_9439,N_9786);
and U10835 (N_10835,N_10344,N_9952);
nand U10836 (N_10836,N_9265,N_9441);
and U10837 (N_10837,N_9868,N_9207);
nand U10838 (N_10838,N_10220,N_10152);
nand U10839 (N_10839,N_9631,N_10202);
nor U10840 (N_10840,N_9177,N_9041);
xor U10841 (N_10841,N_9888,N_9264);
nor U10842 (N_10842,N_9427,N_9514);
nand U10843 (N_10843,N_10398,N_9828);
and U10844 (N_10844,N_9330,N_10466);
and U10845 (N_10845,N_9980,N_9189);
or U10846 (N_10846,N_10134,N_9894);
nand U10847 (N_10847,N_9075,N_9849);
and U10848 (N_10848,N_10328,N_9742);
or U10849 (N_10849,N_10411,N_9634);
and U10850 (N_10850,N_10239,N_10449);
nand U10851 (N_10851,N_9320,N_10218);
and U10852 (N_10852,N_9055,N_9660);
and U10853 (N_10853,N_10062,N_10497);
nand U10854 (N_10854,N_10206,N_9628);
xor U10855 (N_10855,N_9540,N_9257);
nor U10856 (N_10856,N_9783,N_9228);
nor U10857 (N_10857,N_9338,N_10340);
nor U10858 (N_10858,N_9932,N_10431);
nor U10859 (N_10859,N_10476,N_9360);
xor U10860 (N_10860,N_10082,N_9771);
and U10861 (N_10861,N_10366,N_9493);
nor U10862 (N_10862,N_9846,N_10401);
or U10863 (N_10863,N_9645,N_9142);
nand U10864 (N_10864,N_9729,N_10113);
nor U10865 (N_10865,N_9671,N_9905);
and U10866 (N_10866,N_9359,N_9970);
nand U10867 (N_10867,N_9530,N_9417);
or U10868 (N_10868,N_9848,N_9020);
and U10869 (N_10869,N_10126,N_9803);
or U10870 (N_10870,N_10086,N_9100);
xor U10871 (N_10871,N_10325,N_9217);
or U10872 (N_10872,N_9332,N_10236);
nor U10873 (N_10873,N_9555,N_9110);
or U10874 (N_10874,N_9221,N_9161);
or U10875 (N_10875,N_9678,N_9438);
nand U10876 (N_10876,N_9222,N_10327);
or U10877 (N_10877,N_9585,N_9925);
nand U10878 (N_10878,N_9299,N_10295);
or U10879 (N_10879,N_9755,N_10425);
nand U10880 (N_10880,N_10432,N_9064);
or U10881 (N_10881,N_10262,N_9823);
and U10882 (N_10882,N_9934,N_10144);
and U10883 (N_10883,N_10324,N_9593);
nor U10884 (N_10884,N_9017,N_10479);
nand U10885 (N_10885,N_10377,N_9176);
nor U10886 (N_10886,N_9788,N_9777);
and U10887 (N_10887,N_9763,N_9548);
nor U10888 (N_10888,N_9808,N_10136);
nor U10889 (N_10889,N_10084,N_9538);
nor U10890 (N_10890,N_10167,N_10189);
nor U10891 (N_10891,N_10012,N_10209);
and U10892 (N_10892,N_9293,N_10064);
nor U10893 (N_10893,N_9984,N_9209);
xor U10894 (N_10894,N_9568,N_9115);
xnor U10895 (N_10895,N_9982,N_9561);
nor U10896 (N_10896,N_9741,N_10467);
nand U10897 (N_10897,N_9133,N_9036);
nor U10898 (N_10898,N_9523,N_9407);
nand U10899 (N_10899,N_9778,N_9489);
or U10900 (N_10900,N_9250,N_9838);
or U10901 (N_10901,N_9007,N_9367);
nand U10902 (N_10902,N_9911,N_10098);
nor U10903 (N_10903,N_9267,N_9724);
nand U10904 (N_10904,N_10182,N_9958);
nand U10905 (N_10905,N_9919,N_9924);
and U10906 (N_10906,N_9357,N_10444);
and U10907 (N_10907,N_10252,N_9198);
and U10908 (N_10908,N_10490,N_9968);
or U10909 (N_10909,N_9676,N_9165);
nand U10910 (N_10910,N_9818,N_9570);
nor U10911 (N_10911,N_9090,N_10006);
nor U10912 (N_10912,N_9754,N_10233);
xor U10913 (N_10913,N_9890,N_9895);
or U10914 (N_10914,N_10382,N_9611);
and U10915 (N_10915,N_9971,N_9410);
or U10916 (N_10916,N_9580,N_9749);
nand U10917 (N_10917,N_9998,N_9594);
or U10918 (N_10918,N_10017,N_9683);
and U10919 (N_10919,N_9295,N_10266);
or U10920 (N_10920,N_9185,N_9188);
and U10921 (N_10921,N_9278,N_9050);
xnor U10922 (N_10922,N_9048,N_9363);
nor U10923 (N_10923,N_9080,N_10217);
and U10924 (N_10924,N_9474,N_9750);
and U10925 (N_10925,N_9695,N_9536);
and U10926 (N_10926,N_10049,N_10088);
nor U10927 (N_10927,N_9107,N_10409);
and U10928 (N_10928,N_9253,N_10201);
nand U10929 (N_10929,N_9101,N_9210);
and U10930 (N_10930,N_10241,N_9931);
and U10931 (N_10931,N_9972,N_9344);
or U10932 (N_10932,N_9677,N_9807);
nand U10933 (N_10933,N_9609,N_9300);
and U10934 (N_10934,N_10400,N_10424);
or U10935 (N_10935,N_10364,N_9319);
or U10936 (N_10936,N_9345,N_9488);
nor U10937 (N_10937,N_10353,N_9875);
or U10938 (N_10938,N_9258,N_9734);
and U10939 (N_10939,N_10309,N_9526);
xnor U10940 (N_10940,N_9324,N_10458);
nor U10941 (N_10941,N_9450,N_10187);
or U10942 (N_10942,N_10197,N_10318);
and U10943 (N_10943,N_10229,N_10214);
xor U10944 (N_10944,N_9975,N_9272);
or U10945 (N_10945,N_9897,N_9616);
and U10946 (N_10946,N_10014,N_10468);
and U10947 (N_10947,N_10244,N_9675);
nor U10948 (N_10948,N_9380,N_10438);
or U10949 (N_10949,N_9126,N_9522);
or U10950 (N_10950,N_9113,N_9061);
nand U10951 (N_10951,N_9506,N_9557);
nand U10952 (N_10952,N_10141,N_9518);
nor U10953 (N_10953,N_9132,N_9708);
nor U10954 (N_10954,N_9004,N_10009);
or U10955 (N_10955,N_9108,N_10005);
or U10956 (N_10956,N_9159,N_10099);
or U10957 (N_10957,N_9156,N_10339);
nand U10958 (N_10958,N_9291,N_9152);
or U10959 (N_10959,N_10238,N_10275);
nor U10960 (N_10960,N_9425,N_9899);
or U10961 (N_10961,N_9205,N_9698);
nand U10962 (N_10962,N_9117,N_10407);
nand U10963 (N_10963,N_9621,N_9565);
and U10964 (N_10964,N_10453,N_9996);
nand U10965 (N_10965,N_9444,N_9575);
nor U10966 (N_10966,N_9501,N_9423);
and U10967 (N_10967,N_10273,N_9158);
nand U10968 (N_10968,N_10459,N_10178);
nor U10969 (N_10969,N_10234,N_9505);
or U10970 (N_10970,N_9331,N_9633);
and U10971 (N_10971,N_9595,N_10372);
nand U10972 (N_10972,N_10077,N_10205);
or U10973 (N_10973,N_10314,N_10250);
nor U10974 (N_10974,N_9292,N_9605);
nand U10975 (N_10975,N_10109,N_9714);
or U10976 (N_10976,N_9979,N_10158);
or U10977 (N_10977,N_9733,N_10489);
or U10978 (N_10978,N_10291,N_9873);
or U10979 (N_10979,N_9162,N_9551);
nor U10980 (N_10980,N_9587,N_9999);
and U10981 (N_10981,N_9666,N_9831);
and U10982 (N_10982,N_9892,N_9863);
or U10983 (N_10983,N_10116,N_10190);
or U10984 (N_10984,N_9065,N_9625);
xor U10985 (N_10985,N_9102,N_9078);
nand U10986 (N_10986,N_10135,N_9658);
and U10987 (N_10987,N_9206,N_9280);
and U10988 (N_10988,N_9491,N_9802);
nor U10989 (N_10989,N_9854,N_9766);
and U10990 (N_10990,N_9758,N_10143);
nor U10991 (N_10991,N_10251,N_9342);
or U10992 (N_10992,N_10337,N_9715);
nand U10993 (N_10993,N_9747,N_10051);
nor U10994 (N_10994,N_9574,N_10237);
xor U10995 (N_10995,N_9325,N_9309);
and U10996 (N_10996,N_10198,N_9719);
or U10997 (N_10997,N_9477,N_9964);
nand U10998 (N_10998,N_9194,N_9978);
or U10999 (N_10999,N_9356,N_9997);
nor U11000 (N_11000,N_10114,N_9515);
and U11001 (N_11001,N_9829,N_9529);
nand U11002 (N_11002,N_9697,N_10435);
and U11003 (N_11003,N_9664,N_9399);
or U11004 (N_11004,N_9681,N_9382);
and U11005 (N_11005,N_9826,N_10352);
nand U11006 (N_11006,N_9211,N_9069);
nand U11007 (N_11007,N_9938,N_9195);
and U11008 (N_11008,N_9916,N_10429);
or U11009 (N_11009,N_10493,N_9539);
or U11010 (N_11010,N_9716,N_10359);
and U11011 (N_11011,N_9103,N_10428);
nor U11012 (N_11012,N_10420,N_9546);
nor U11013 (N_11013,N_9175,N_10119);
or U11014 (N_11014,N_9365,N_9442);
xor U11015 (N_11015,N_10452,N_9416);
nand U11016 (N_11016,N_10074,N_9401);
xnor U11017 (N_11017,N_10348,N_9266);
nor U11018 (N_11018,N_9468,N_10312);
or U11019 (N_11019,N_9969,N_9531);
nor U11020 (N_11020,N_10457,N_9379);
nor U11021 (N_11021,N_9445,N_9225);
or U11022 (N_11022,N_9835,N_10265);
and U11023 (N_11023,N_9400,N_9426);
and U11024 (N_11024,N_9471,N_9203);
xor U11025 (N_11025,N_10057,N_10351);
nand U11026 (N_11026,N_9617,N_9308);
or U11027 (N_11027,N_9700,N_9584);
and U11028 (N_11028,N_9212,N_9086);
or U11029 (N_11029,N_9976,N_9543);
or U11030 (N_11030,N_10347,N_9880);
or U11031 (N_11031,N_9098,N_10035);
nor U11032 (N_11032,N_9852,N_10101);
or U11033 (N_11033,N_9010,N_9460);
nor U11034 (N_11034,N_9603,N_9789);
xor U11035 (N_11035,N_9022,N_9454);
nand U11036 (N_11036,N_9030,N_9396);
nand U11037 (N_11037,N_10361,N_9346);
xnor U11038 (N_11038,N_10482,N_9134);
nand U11039 (N_11039,N_9735,N_9640);
nand U11040 (N_11040,N_10296,N_9843);
or U11041 (N_11041,N_9463,N_9850);
nor U11042 (N_11042,N_9462,N_10007);
or U11043 (N_11043,N_9025,N_9767);
nand U11044 (N_11044,N_10267,N_9774);
nor U11045 (N_11045,N_10302,N_9535);
nand U11046 (N_11046,N_10160,N_9822);
nand U11047 (N_11047,N_10381,N_9437);
xor U11048 (N_11048,N_9470,N_10393);
or U11049 (N_11049,N_10059,N_10096);
or U11050 (N_11050,N_10004,N_9509);
and U11051 (N_11051,N_9839,N_9582);
nor U11052 (N_11052,N_10177,N_9796);
nand U11053 (N_11053,N_9981,N_9686);
nand U11054 (N_11054,N_9933,N_9579);
and U11055 (N_11055,N_9251,N_10290);
or U11056 (N_11056,N_10248,N_9693);
nor U11057 (N_11057,N_10362,N_9712);
and U11058 (N_11058,N_10121,N_10391);
or U11059 (N_11059,N_10045,N_9844);
or U11060 (N_11060,N_9855,N_10480);
xnor U11061 (N_11061,N_10470,N_9937);
nor U11062 (N_11062,N_9541,N_9373);
and U11063 (N_11063,N_9626,N_10354);
nor U11064 (N_11064,N_10056,N_9866);
nand U11065 (N_11065,N_9564,N_9170);
or U11066 (N_11066,N_9887,N_9323);
and U11067 (N_11067,N_10268,N_9197);
xor U11068 (N_11068,N_10477,N_10286);
nor U11069 (N_11069,N_9710,N_10416);
nor U11070 (N_11070,N_10456,N_9358);
and U11071 (N_11071,N_10010,N_9943);
nand U11072 (N_11072,N_9648,N_9819);
and U11073 (N_11073,N_9226,N_9578);
nand U11074 (N_11074,N_9606,N_10442);
nor U11075 (N_11075,N_9492,N_10106);
nand U11076 (N_11076,N_10019,N_9388);
nor U11077 (N_11077,N_9024,N_9930);
or U11078 (N_11078,N_9759,N_10173);
nand U11079 (N_11079,N_9610,N_10130);
and U11080 (N_11080,N_10125,N_10437);
or U11081 (N_11081,N_9662,N_9878);
nand U11082 (N_11082,N_9923,N_9563);
nor U11083 (N_11083,N_9524,N_10447);
or U11084 (N_11084,N_10421,N_10058);
or U11085 (N_11085,N_9527,N_10073);
nand U11086 (N_11086,N_9953,N_9770);
and U11087 (N_11087,N_9562,N_9637);
nand U11088 (N_11088,N_9430,N_9063);
and U11089 (N_11089,N_9668,N_10294);
and U11090 (N_11090,N_9453,N_9739);
or U11091 (N_11091,N_9072,N_9081);
and U11092 (N_11092,N_9220,N_9157);
nand U11093 (N_11093,N_9824,N_9832);
nor U11094 (N_11094,N_10159,N_9150);
nor U11095 (N_11095,N_9946,N_10249);
nor U11096 (N_11096,N_9782,N_9009);
or U11097 (N_11097,N_10287,N_9027);
or U11098 (N_11098,N_9051,N_9229);
nand U11099 (N_11099,N_10196,N_10157);
nor U11100 (N_11100,N_9629,N_9792);
nor U11101 (N_11101,N_9392,N_9909);
and U11102 (N_11102,N_10199,N_10094);
xnor U11103 (N_11103,N_9566,N_10216);
xnor U11104 (N_11104,N_9711,N_9455);
and U11105 (N_11105,N_10323,N_9056);
nor U11106 (N_11106,N_9508,N_9130);
or U11107 (N_11107,N_9071,N_10461);
or U11108 (N_11108,N_10066,N_9912);
and U11109 (N_11109,N_9354,N_10223);
and U11110 (N_11110,N_10402,N_10030);
nand U11111 (N_11111,N_9612,N_10120);
nor U11112 (N_11112,N_9494,N_10486);
nand U11113 (N_11113,N_9973,N_10211);
and U11114 (N_11114,N_10498,N_9301);
and U11115 (N_11115,N_10228,N_10091);
nor U11116 (N_11116,N_10462,N_9737);
and U11117 (N_11117,N_9199,N_9275);
nand U11118 (N_11118,N_10046,N_10247);
or U11119 (N_11119,N_9935,N_10360);
xnor U11120 (N_11120,N_9411,N_10403);
xnor U11121 (N_11121,N_10285,N_10436);
nand U11122 (N_11122,N_9641,N_9569);
xor U11123 (N_11123,N_10446,N_9730);
nor U11124 (N_11124,N_9588,N_10464);
or U11125 (N_11125,N_9179,N_9094);
and U11126 (N_11126,N_9723,N_10389);
or U11127 (N_11127,N_10240,N_9297);
nor U11128 (N_11128,N_9088,N_9242);
xnor U11129 (N_11129,N_9483,N_9333);
or U11130 (N_11130,N_10445,N_9096);
and U11131 (N_11131,N_9740,N_9409);
or U11132 (N_11132,N_10242,N_10226);
xnor U11133 (N_11133,N_10225,N_9045);
xnor U11134 (N_11134,N_10138,N_9655);
nor U11135 (N_11135,N_9314,N_9528);
and U11136 (N_11136,N_9618,N_9918);
and U11137 (N_11137,N_10153,N_9504);
nor U11138 (N_11138,N_9962,N_9791);
nor U11139 (N_11139,N_9271,N_9647);
and U11140 (N_11140,N_9339,N_9811);
xor U11141 (N_11141,N_9825,N_10090);
nand U11142 (N_11142,N_9395,N_9336);
xnor U11143 (N_11143,N_9757,N_9283);
nand U11144 (N_11144,N_9995,N_9311);
nand U11145 (N_11145,N_10276,N_9591);
or U11146 (N_11146,N_9764,N_9180);
nand U11147 (N_11147,N_10207,N_10047);
or U11148 (N_11148,N_10180,N_9950);
xor U11149 (N_11149,N_10052,N_10350);
nor U11150 (N_11150,N_10293,N_9650);
or U11151 (N_11151,N_9091,N_9485);
or U11152 (N_11152,N_9910,N_9405);
or U11153 (N_11153,N_10245,N_10000);
nor U11154 (N_11154,N_10329,N_10132);
and U11155 (N_11155,N_9780,N_9347);
nor U11156 (N_11156,N_10349,N_9957);
and U11157 (N_11157,N_9079,N_9208);
nor U11158 (N_11158,N_10186,N_10346);
and U11159 (N_11159,N_9432,N_10308);
nor U11160 (N_11160,N_9989,N_9502);
nor U11161 (N_11161,N_9434,N_9105);
xnor U11162 (N_11162,N_9490,N_10365);
xor U11163 (N_11163,N_10319,N_10417);
nor U11164 (N_11164,N_9795,N_9533);
nand U11165 (N_11165,N_9914,N_9576);
nand U11166 (N_11166,N_9263,N_9851);
nor U11167 (N_11167,N_10259,N_10029);
and U11168 (N_11168,N_9279,N_9713);
nand U11169 (N_11169,N_9836,N_9620);
nor U11170 (N_11170,N_9745,N_10277);
nor U11171 (N_11171,N_10179,N_10258);
nor U11172 (N_11172,N_9567,N_10439);
nand U11173 (N_11173,N_9329,N_9586);
nor U11174 (N_11174,N_10316,N_9429);
and U11175 (N_11175,N_9793,N_10375);
nor U11176 (N_11176,N_9900,N_9191);
and U11177 (N_11177,N_9216,N_9779);
nor U11178 (N_11178,N_9961,N_9599);
nor U11179 (N_11179,N_9772,N_9313);
or U11180 (N_11180,N_9288,N_9691);
nand U11181 (N_11181,N_9891,N_9343);
nand U11182 (N_11182,N_10104,N_10330);
and U11183 (N_11183,N_9507,N_10162);
nor U11184 (N_11184,N_9404,N_9456);
and U11185 (N_11185,N_10460,N_10176);
xor U11186 (N_11186,N_9643,N_9316);
nor U11187 (N_11187,N_9052,N_10387);
or U11188 (N_11188,N_9084,N_9663);
xor U11189 (N_11189,N_10087,N_9287);
nand U11190 (N_11190,N_10105,N_9885);
or U11191 (N_11191,N_9310,N_10281);
or U11192 (N_11192,N_9224,N_9920);
nor U11193 (N_11193,N_9709,N_9127);
nand U11194 (N_11194,N_10440,N_9827);
and U11195 (N_11195,N_9801,N_10443);
nor U11196 (N_11196,N_9583,N_10419);
or U11197 (N_11197,N_10388,N_10161);
nor U11198 (N_11198,N_10368,N_10212);
or U11199 (N_11199,N_9239,N_9960);
nand U11200 (N_11200,N_9927,N_9542);
or U11201 (N_11201,N_9776,N_9977);
nand U11202 (N_11202,N_10280,N_9262);
or U11203 (N_11203,N_10283,N_10146);
and U11204 (N_11204,N_10129,N_10397);
nor U11205 (N_11205,N_9500,N_9592);
xnor U11206 (N_11206,N_9862,N_10491);
nand U11207 (N_11207,N_10499,N_10172);
nor U11208 (N_11208,N_9859,N_9762);
nand U11209 (N_11209,N_9118,N_9993);
or U11210 (N_11210,N_10124,N_10219);
nand U11211 (N_11211,N_10485,N_10454);
nand U11212 (N_11212,N_10112,N_9945);
nor U11213 (N_11213,N_10033,N_9083);
nor U11214 (N_11214,N_9349,N_10378);
xor U11215 (N_11215,N_9054,N_9193);
xor U11216 (N_11216,N_10356,N_10221);
and U11217 (N_11217,N_10495,N_9865);
or U11218 (N_11218,N_10193,N_9883);
and U11219 (N_11219,N_9985,N_10026);
nor U11220 (N_11220,N_9473,N_9815);
xnor U11221 (N_11221,N_9368,N_10390);
nor U11222 (N_11222,N_9049,N_9296);
and U11223 (N_11223,N_9926,N_9241);
nor U11224 (N_11224,N_9688,N_9033);
nor U11225 (N_11225,N_9424,N_9614);
and U11226 (N_11226,N_9120,N_10253);
or U11227 (N_11227,N_9043,N_9315);
and U11228 (N_11228,N_10384,N_9231);
or U11229 (N_11229,N_9534,N_10110);
or U11230 (N_11230,N_9459,N_9341);
nor U11231 (N_11231,N_10369,N_9238);
xor U11232 (N_11232,N_9140,N_9738);
and U11233 (N_11233,N_9053,N_9498);
xnor U11234 (N_11234,N_10070,N_9318);
nor U11235 (N_11235,N_9412,N_9073);
nor U11236 (N_11236,N_9886,N_9726);
nand U11237 (N_11237,N_10034,N_9422);
and U11238 (N_11238,N_9011,N_10149);
and U11239 (N_11239,N_9406,N_9361);
or U11240 (N_11240,N_9965,N_9289);
or U11241 (N_11241,N_10243,N_10303);
and U11242 (N_11242,N_10376,N_10373);
and U11243 (N_11243,N_9939,N_10020);
and U11244 (N_11244,N_9904,N_9192);
xor U11245 (N_11245,N_9397,N_9364);
nand U11246 (N_11246,N_9370,N_9077);
and U11247 (N_11247,N_9255,N_9254);
xor U11248 (N_11248,N_9861,N_9903);
nor U11249 (N_11249,N_9252,N_9277);
nand U11250 (N_11250,N_9936,N_9727);
nand U11251 (N_11251,N_9379,N_10106);
or U11252 (N_11252,N_9638,N_9387);
xor U11253 (N_11253,N_9000,N_10455);
or U11254 (N_11254,N_9095,N_9118);
nor U11255 (N_11255,N_10462,N_10113);
and U11256 (N_11256,N_10354,N_10496);
and U11257 (N_11257,N_9218,N_9086);
and U11258 (N_11258,N_9293,N_9002);
and U11259 (N_11259,N_9891,N_9306);
or U11260 (N_11260,N_9838,N_9830);
nor U11261 (N_11261,N_10000,N_9289);
xor U11262 (N_11262,N_9335,N_9796);
nand U11263 (N_11263,N_10234,N_9199);
and U11264 (N_11264,N_9157,N_9185);
or U11265 (N_11265,N_9846,N_9658);
nand U11266 (N_11266,N_10141,N_9370);
and U11267 (N_11267,N_9881,N_9676);
nand U11268 (N_11268,N_9187,N_9382);
or U11269 (N_11269,N_9767,N_9161);
and U11270 (N_11270,N_10088,N_10216);
and U11271 (N_11271,N_9183,N_9500);
and U11272 (N_11272,N_9947,N_9465);
or U11273 (N_11273,N_9867,N_9396);
and U11274 (N_11274,N_9654,N_9432);
nor U11275 (N_11275,N_10037,N_9158);
nor U11276 (N_11276,N_9361,N_9009);
or U11277 (N_11277,N_10451,N_9399);
nand U11278 (N_11278,N_9484,N_9245);
nor U11279 (N_11279,N_9228,N_9100);
and U11280 (N_11280,N_9682,N_9324);
and U11281 (N_11281,N_9913,N_9029);
or U11282 (N_11282,N_9525,N_9227);
or U11283 (N_11283,N_9817,N_9728);
and U11284 (N_11284,N_9349,N_9815);
nor U11285 (N_11285,N_9625,N_10156);
or U11286 (N_11286,N_10317,N_9086);
nand U11287 (N_11287,N_9035,N_9875);
nor U11288 (N_11288,N_9566,N_9117);
and U11289 (N_11289,N_9526,N_9829);
and U11290 (N_11290,N_10455,N_10496);
or U11291 (N_11291,N_9803,N_10117);
or U11292 (N_11292,N_9498,N_10348);
and U11293 (N_11293,N_10029,N_10446);
nor U11294 (N_11294,N_9784,N_9419);
xnor U11295 (N_11295,N_9765,N_10233);
and U11296 (N_11296,N_10371,N_9659);
and U11297 (N_11297,N_10222,N_9015);
nor U11298 (N_11298,N_9574,N_9573);
or U11299 (N_11299,N_9595,N_10427);
nand U11300 (N_11300,N_9877,N_9918);
or U11301 (N_11301,N_10266,N_9422);
xor U11302 (N_11302,N_9602,N_10300);
and U11303 (N_11303,N_10105,N_9508);
nand U11304 (N_11304,N_9964,N_10111);
and U11305 (N_11305,N_9893,N_9641);
or U11306 (N_11306,N_9907,N_9026);
and U11307 (N_11307,N_9816,N_9660);
and U11308 (N_11308,N_10169,N_9020);
xor U11309 (N_11309,N_10081,N_10031);
nor U11310 (N_11310,N_10046,N_9301);
nor U11311 (N_11311,N_9441,N_9376);
nor U11312 (N_11312,N_10376,N_9690);
nor U11313 (N_11313,N_9104,N_9308);
nor U11314 (N_11314,N_9318,N_10321);
and U11315 (N_11315,N_9204,N_10149);
nand U11316 (N_11316,N_9819,N_9880);
nor U11317 (N_11317,N_9651,N_10124);
nor U11318 (N_11318,N_10005,N_9906);
nor U11319 (N_11319,N_9858,N_10209);
nor U11320 (N_11320,N_9504,N_9384);
nand U11321 (N_11321,N_9299,N_10130);
nand U11322 (N_11322,N_9276,N_10356);
and U11323 (N_11323,N_9517,N_9080);
and U11324 (N_11324,N_9667,N_10069);
nor U11325 (N_11325,N_10045,N_9220);
or U11326 (N_11326,N_10056,N_9428);
and U11327 (N_11327,N_9344,N_9476);
or U11328 (N_11328,N_10186,N_10135);
nor U11329 (N_11329,N_9156,N_10009);
and U11330 (N_11330,N_9666,N_10163);
nand U11331 (N_11331,N_10244,N_9479);
or U11332 (N_11332,N_10060,N_9870);
or U11333 (N_11333,N_10031,N_9531);
or U11334 (N_11334,N_9278,N_10342);
nand U11335 (N_11335,N_9651,N_9924);
or U11336 (N_11336,N_10112,N_9407);
nand U11337 (N_11337,N_9515,N_10015);
nand U11338 (N_11338,N_9342,N_9576);
nor U11339 (N_11339,N_9510,N_9386);
or U11340 (N_11340,N_10137,N_9662);
and U11341 (N_11341,N_9791,N_10009);
and U11342 (N_11342,N_9612,N_9622);
nor U11343 (N_11343,N_9466,N_9075);
and U11344 (N_11344,N_9273,N_9603);
xor U11345 (N_11345,N_9325,N_9120);
nor U11346 (N_11346,N_10124,N_10371);
and U11347 (N_11347,N_9039,N_10187);
nor U11348 (N_11348,N_9368,N_10201);
nand U11349 (N_11349,N_9818,N_9097);
and U11350 (N_11350,N_9261,N_9206);
or U11351 (N_11351,N_9650,N_10312);
and U11352 (N_11352,N_9078,N_9815);
or U11353 (N_11353,N_9344,N_9020);
or U11354 (N_11354,N_9066,N_10389);
nand U11355 (N_11355,N_9095,N_9073);
nor U11356 (N_11356,N_9501,N_10406);
nor U11357 (N_11357,N_9603,N_9121);
and U11358 (N_11358,N_10074,N_10203);
and U11359 (N_11359,N_9747,N_9626);
and U11360 (N_11360,N_9796,N_9958);
nand U11361 (N_11361,N_9993,N_10359);
nand U11362 (N_11362,N_9821,N_9764);
nand U11363 (N_11363,N_10260,N_9397);
xnor U11364 (N_11364,N_9965,N_9110);
and U11365 (N_11365,N_9942,N_9764);
or U11366 (N_11366,N_10363,N_9694);
nor U11367 (N_11367,N_9809,N_10467);
and U11368 (N_11368,N_10135,N_9089);
or U11369 (N_11369,N_10487,N_9188);
xor U11370 (N_11370,N_10340,N_10217);
or U11371 (N_11371,N_10110,N_9281);
or U11372 (N_11372,N_9058,N_9017);
xor U11373 (N_11373,N_9011,N_9964);
nand U11374 (N_11374,N_9952,N_9614);
nor U11375 (N_11375,N_10052,N_9475);
and U11376 (N_11376,N_10257,N_10326);
or U11377 (N_11377,N_9651,N_9591);
nor U11378 (N_11378,N_9105,N_9694);
nand U11379 (N_11379,N_9427,N_9922);
xor U11380 (N_11380,N_9169,N_10259);
nand U11381 (N_11381,N_10272,N_10080);
nand U11382 (N_11382,N_9277,N_9881);
nor U11383 (N_11383,N_10055,N_10450);
nand U11384 (N_11384,N_10466,N_10047);
nand U11385 (N_11385,N_9200,N_10156);
nand U11386 (N_11386,N_9923,N_9604);
and U11387 (N_11387,N_9609,N_9132);
nand U11388 (N_11388,N_9818,N_10455);
xor U11389 (N_11389,N_9855,N_9560);
nor U11390 (N_11390,N_10248,N_9598);
nor U11391 (N_11391,N_9332,N_9581);
nand U11392 (N_11392,N_10483,N_9329);
or U11393 (N_11393,N_9846,N_9515);
and U11394 (N_11394,N_9962,N_10333);
nor U11395 (N_11395,N_10330,N_9523);
nand U11396 (N_11396,N_10474,N_10245);
nand U11397 (N_11397,N_10067,N_10251);
nand U11398 (N_11398,N_9961,N_10457);
nor U11399 (N_11399,N_10051,N_10272);
and U11400 (N_11400,N_9776,N_10490);
and U11401 (N_11401,N_9501,N_9493);
and U11402 (N_11402,N_9003,N_9757);
and U11403 (N_11403,N_9920,N_9292);
or U11404 (N_11404,N_9655,N_10169);
and U11405 (N_11405,N_9557,N_10172);
or U11406 (N_11406,N_10308,N_10033);
xor U11407 (N_11407,N_10492,N_9590);
and U11408 (N_11408,N_9554,N_9951);
or U11409 (N_11409,N_9614,N_9051);
xnor U11410 (N_11410,N_10207,N_10390);
nand U11411 (N_11411,N_9369,N_9972);
xnor U11412 (N_11412,N_9598,N_9683);
or U11413 (N_11413,N_9705,N_10382);
nand U11414 (N_11414,N_9520,N_10130);
and U11415 (N_11415,N_9739,N_9112);
and U11416 (N_11416,N_9609,N_9447);
and U11417 (N_11417,N_9074,N_9487);
and U11418 (N_11418,N_9972,N_9057);
nand U11419 (N_11419,N_9204,N_10217);
and U11420 (N_11420,N_10492,N_10403);
or U11421 (N_11421,N_9973,N_10414);
nor U11422 (N_11422,N_10097,N_9325);
or U11423 (N_11423,N_9601,N_9619);
and U11424 (N_11424,N_10033,N_9501);
or U11425 (N_11425,N_10174,N_9769);
nand U11426 (N_11426,N_9787,N_9158);
nand U11427 (N_11427,N_9328,N_9508);
xor U11428 (N_11428,N_9264,N_9522);
and U11429 (N_11429,N_10272,N_9946);
and U11430 (N_11430,N_10163,N_9867);
nor U11431 (N_11431,N_9955,N_9751);
nor U11432 (N_11432,N_10041,N_9930);
and U11433 (N_11433,N_10113,N_9747);
nor U11434 (N_11434,N_9004,N_9521);
and U11435 (N_11435,N_9605,N_10088);
nand U11436 (N_11436,N_9319,N_10384);
and U11437 (N_11437,N_10474,N_10074);
xor U11438 (N_11438,N_9465,N_9766);
nor U11439 (N_11439,N_9788,N_9321);
nor U11440 (N_11440,N_10014,N_10340);
or U11441 (N_11441,N_10241,N_10450);
nand U11442 (N_11442,N_10032,N_9413);
nand U11443 (N_11443,N_10323,N_9757);
or U11444 (N_11444,N_9314,N_9895);
and U11445 (N_11445,N_10133,N_9549);
nand U11446 (N_11446,N_9695,N_9478);
and U11447 (N_11447,N_9581,N_9913);
nor U11448 (N_11448,N_9460,N_9518);
and U11449 (N_11449,N_9459,N_10487);
nor U11450 (N_11450,N_9337,N_9697);
nand U11451 (N_11451,N_9282,N_9733);
xnor U11452 (N_11452,N_9183,N_9841);
nand U11453 (N_11453,N_10389,N_10291);
nand U11454 (N_11454,N_9790,N_9287);
and U11455 (N_11455,N_9613,N_10034);
nor U11456 (N_11456,N_9942,N_10151);
nand U11457 (N_11457,N_10268,N_9475);
nand U11458 (N_11458,N_9180,N_9517);
and U11459 (N_11459,N_10400,N_9957);
nand U11460 (N_11460,N_9717,N_10416);
and U11461 (N_11461,N_10458,N_9201);
nand U11462 (N_11462,N_10008,N_9404);
nand U11463 (N_11463,N_9245,N_10323);
and U11464 (N_11464,N_10278,N_10338);
nor U11465 (N_11465,N_10095,N_9077);
nand U11466 (N_11466,N_9759,N_9284);
and U11467 (N_11467,N_9766,N_9011);
nand U11468 (N_11468,N_10363,N_9993);
nand U11469 (N_11469,N_9858,N_9959);
or U11470 (N_11470,N_10316,N_10189);
nor U11471 (N_11471,N_9288,N_9311);
or U11472 (N_11472,N_10480,N_9597);
or U11473 (N_11473,N_10375,N_9222);
nand U11474 (N_11474,N_9090,N_9136);
or U11475 (N_11475,N_9103,N_9584);
nand U11476 (N_11476,N_9934,N_9083);
nand U11477 (N_11477,N_9903,N_9722);
nor U11478 (N_11478,N_9171,N_9861);
nor U11479 (N_11479,N_10085,N_9979);
nor U11480 (N_11480,N_9732,N_9393);
and U11481 (N_11481,N_9824,N_9815);
or U11482 (N_11482,N_9651,N_9471);
nor U11483 (N_11483,N_9928,N_10102);
nand U11484 (N_11484,N_10356,N_9790);
and U11485 (N_11485,N_9476,N_9209);
nand U11486 (N_11486,N_9537,N_10336);
nand U11487 (N_11487,N_9048,N_9310);
and U11488 (N_11488,N_10112,N_9891);
nand U11489 (N_11489,N_9270,N_9529);
and U11490 (N_11490,N_9131,N_10275);
and U11491 (N_11491,N_9581,N_9146);
or U11492 (N_11492,N_9443,N_10280);
xnor U11493 (N_11493,N_10212,N_9387);
nor U11494 (N_11494,N_9382,N_9064);
nand U11495 (N_11495,N_9848,N_9580);
or U11496 (N_11496,N_9441,N_9969);
nor U11497 (N_11497,N_9560,N_10429);
nor U11498 (N_11498,N_10129,N_10453);
nor U11499 (N_11499,N_9824,N_9201);
nand U11500 (N_11500,N_9939,N_9890);
and U11501 (N_11501,N_9446,N_9889);
nand U11502 (N_11502,N_10443,N_9313);
nor U11503 (N_11503,N_10302,N_9737);
nor U11504 (N_11504,N_10246,N_10289);
or U11505 (N_11505,N_9896,N_9645);
and U11506 (N_11506,N_9352,N_9096);
nor U11507 (N_11507,N_10466,N_9982);
or U11508 (N_11508,N_9139,N_9684);
nor U11509 (N_11509,N_10439,N_9986);
xnor U11510 (N_11510,N_10410,N_9769);
xnor U11511 (N_11511,N_9485,N_10091);
nor U11512 (N_11512,N_9472,N_9069);
or U11513 (N_11513,N_9184,N_9039);
nor U11514 (N_11514,N_9876,N_9748);
nor U11515 (N_11515,N_9827,N_10380);
or U11516 (N_11516,N_9756,N_10408);
xnor U11517 (N_11517,N_10144,N_10368);
and U11518 (N_11518,N_9546,N_10335);
nor U11519 (N_11519,N_9141,N_9643);
nor U11520 (N_11520,N_9822,N_9713);
or U11521 (N_11521,N_10354,N_10494);
nor U11522 (N_11522,N_10304,N_9959);
or U11523 (N_11523,N_9584,N_9900);
nor U11524 (N_11524,N_9120,N_10245);
and U11525 (N_11525,N_9583,N_9306);
nand U11526 (N_11526,N_9089,N_9375);
or U11527 (N_11527,N_9614,N_10245);
nand U11528 (N_11528,N_10064,N_10420);
xnor U11529 (N_11529,N_9591,N_10008);
and U11530 (N_11530,N_9104,N_10430);
or U11531 (N_11531,N_9988,N_10377);
xnor U11532 (N_11532,N_9034,N_9487);
and U11533 (N_11533,N_10115,N_9739);
or U11534 (N_11534,N_10498,N_9832);
or U11535 (N_11535,N_10228,N_9642);
xnor U11536 (N_11536,N_9879,N_10356);
nor U11537 (N_11537,N_9343,N_10153);
or U11538 (N_11538,N_10495,N_10477);
and U11539 (N_11539,N_10311,N_9032);
or U11540 (N_11540,N_9908,N_9740);
nor U11541 (N_11541,N_10303,N_9714);
or U11542 (N_11542,N_10039,N_9778);
and U11543 (N_11543,N_9498,N_9329);
and U11544 (N_11544,N_9879,N_9148);
and U11545 (N_11545,N_9209,N_9097);
or U11546 (N_11546,N_9683,N_9455);
xnor U11547 (N_11547,N_9402,N_9378);
or U11548 (N_11548,N_9534,N_9803);
or U11549 (N_11549,N_9377,N_9302);
or U11550 (N_11550,N_9065,N_9358);
nand U11551 (N_11551,N_9245,N_9411);
xnor U11552 (N_11552,N_10034,N_9073);
or U11553 (N_11553,N_10492,N_9962);
nor U11554 (N_11554,N_9303,N_10141);
nand U11555 (N_11555,N_10455,N_9255);
or U11556 (N_11556,N_9914,N_9438);
xor U11557 (N_11557,N_9735,N_9376);
and U11558 (N_11558,N_9273,N_10378);
nor U11559 (N_11559,N_10400,N_10083);
or U11560 (N_11560,N_9790,N_9294);
and U11561 (N_11561,N_9643,N_9086);
and U11562 (N_11562,N_9242,N_9453);
or U11563 (N_11563,N_10273,N_9032);
nor U11564 (N_11564,N_10353,N_9994);
nor U11565 (N_11565,N_9989,N_9731);
and U11566 (N_11566,N_9683,N_9671);
or U11567 (N_11567,N_9250,N_10010);
nand U11568 (N_11568,N_9638,N_9025);
and U11569 (N_11569,N_10418,N_9464);
nand U11570 (N_11570,N_9280,N_9637);
and U11571 (N_11571,N_10458,N_9362);
or U11572 (N_11572,N_10193,N_9974);
and U11573 (N_11573,N_9846,N_9427);
and U11574 (N_11574,N_9408,N_9336);
or U11575 (N_11575,N_9729,N_9446);
nor U11576 (N_11576,N_9028,N_10144);
nor U11577 (N_11577,N_10341,N_9977);
nor U11578 (N_11578,N_9867,N_9286);
nor U11579 (N_11579,N_10159,N_10392);
nor U11580 (N_11580,N_10295,N_10204);
or U11581 (N_11581,N_9344,N_9831);
or U11582 (N_11582,N_9142,N_10027);
nor U11583 (N_11583,N_9722,N_9351);
xor U11584 (N_11584,N_10219,N_10408);
or U11585 (N_11585,N_9552,N_9324);
nand U11586 (N_11586,N_9868,N_10288);
and U11587 (N_11587,N_10390,N_9269);
nor U11588 (N_11588,N_10204,N_9642);
and U11589 (N_11589,N_9813,N_9537);
xor U11590 (N_11590,N_9732,N_9561);
nand U11591 (N_11591,N_9565,N_10038);
nand U11592 (N_11592,N_9249,N_9838);
or U11593 (N_11593,N_9786,N_9192);
nor U11594 (N_11594,N_10234,N_9382);
or U11595 (N_11595,N_9643,N_9416);
nor U11596 (N_11596,N_9192,N_9942);
and U11597 (N_11597,N_9254,N_9778);
and U11598 (N_11598,N_10424,N_9351);
nor U11599 (N_11599,N_10122,N_9062);
and U11600 (N_11600,N_10062,N_10341);
nand U11601 (N_11601,N_9318,N_10281);
and U11602 (N_11602,N_9368,N_10435);
xnor U11603 (N_11603,N_9124,N_9074);
nand U11604 (N_11604,N_10038,N_10422);
or U11605 (N_11605,N_9136,N_9176);
and U11606 (N_11606,N_9678,N_9214);
or U11607 (N_11607,N_9010,N_9483);
or U11608 (N_11608,N_9044,N_10053);
nor U11609 (N_11609,N_10482,N_10202);
nand U11610 (N_11610,N_10186,N_9904);
and U11611 (N_11611,N_9070,N_9128);
xnor U11612 (N_11612,N_10188,N_9355);
nor U11613 (N_11613,N_9797,N_9367);
nor U11614 (N_11614,N_9161,N_9589);
or U11615 (N_11615,N_9380,N_10183);
xnor U11616 (N_11616,N_9529,N_10041);
nand U11617 (N_11617,N_10120,N_10357);
and U11618 (N_11618,N_10121,N_10060);
and U11619 (N_11619,N_9666,N_9447);
and U11620 (N_11620,N_10101,N_9163);
or U11621 (N_11621,N_10385,N_9648);
and U11622 (N_11622,N_10212,N_9001);
nor U11623 (N_11623,N_10046,N_9553);
and U11624 (N_11624,N_9607,N_9793);
xor U11625 (N_11625,N_9539,N_10300);
or U11626 (N_11626,N_9447,N_9335);
nand U11627 (N_11627,N_9350,N_9252);
nand U11628 (N_11628,N_9906,N_10308);
and U11629 (N_11629,N_9464,N_9172);
nand U11630 (N_11630,N_9638,N_10090);
nor U11631 (N_11631,N_9293,N_9057);
or U11632 (N_11632,N_9523,N_9831);
nor U11633 (N_11633,N_10316,N_9701);
nand U11634 (N_11634,N_9404,N_9723);
or U11635 (N_11635,N_9498,N_9397);
or U11636 (N_11636,N_10194,N_9515);
xnor U11637 (N_11637,N_9282,N_9820);
or U11638 (N_11638,N_10189,N_9521);
nor U11639 (N_11639,N_10335,N_9085);
nand U11640 (N_11640,N_10454,N_10449);
nand U11641 (N_11641,N_9316,N_10253);
nor U11642 (N_11642,N_9674,N_10391);
and U11643 (N_11643,N_9534,N_9005);
or U11644 (N_11644,N_10330,N_9061);
nand U11645 (N_11645,N_9596,N_9209);
and U11646 (N_11646,N_10101,N_10315);
nor U11647 (N_11647,N_9058,N_9686);
nor U11648 (N_11648,N_9159,N_9324);
nand U11649 (N_11649,N_9440,N_10419);
or U11650 (N_11650,N_10036,N_9245);
and U11651 (N_11651,N_9747,N_9353);
and U11652 (N_11652,N_9568,N_10427);
or U11653 (N_11653,N_9235,N_9015);
nand U11654 (N_11654,N_9448,N_9204);
nand U11655 (N_11655,N_9384,N_9643);
nor U11656 (N_11656,N_10195,N_9434);
nand U11657 (N_11657,N_9862,N_9655);
and U11658 (N_11658,N_9880,N_10183);
or U11659 (N_11659,N_10161,N_9371);
and U11660 (N_11660,N_9830,N_10074);
or U11661 (N_11661,N_9024,N_9358);
nand U11662 (N_11662,N_9234,N_10290);
nor U11663 (N_11663,N_9594,N_9347);
and U11664 (N_11664,N_10337,N_9021);
or U11665 (N_11665,N_9341,N_9395);
and U11666 (N_11666,N_9435,N_9503);
or U11667 (N_11667,N_9540,N_9951);
or U11668 (N_11668,N_9034,N_9770);
nand U11669 (N_11669,N_9335,N_9327);
or U11670 (N_11670,N_9627,N_9320);
or U11671 (N_11671,N_10328,N_10343);
and U11672 (N_11672,N_9586,N_10321);
and U11673 (N_11673,N_9919,N_10262);
nand U11674 (N_11674,N_9825,N_9548);
nor U11675 (N_11675,N_10204,N_9462);
xnor U11676 (N_11676,N_10300,N_10348);
nand U11677 (N_11677,N_9941,N_9351);
and U11678 (N_11678,N_9944,N_10077);
nor U11679 (N_11679,N_9248,N_9765);
or U11680 (N_11680,N_9577,N_9822);
nor U11681 (N_11681,N_9719,N_9275);
and U11682 (N_11682,N_9655,N_9984);
and U11683 (N_11683,N_9900,N_10443);
nand U11684 (N_11684,N_9330,N_9053);
nand U11685 (N_11685,N_10097,N_10256);
nand U11686 (N_11686,N_10071,N_9764);
xnor U11687 (N_11687,N_10097,N_10226);
and U11688 (N_11688,N_9364,N_10220);
or U11689 (N_11689,N_10408,N_9008);
nor U11690 (N_11690,N_10202,N_9452);
and U11691 (N_11691,N_9909,N_10107);
nand U11692 (N_11692,N_10011,N_9341);
and U11693 (N_11693,N_10301,N_9931);
nand U11694 (N_11694,N_10408,N_9314);
nor U11695 (N_11695,N_9401,N_9427);
nor U11696 (N_11696,N_9317,N_10108);
or U11697 (N_11697,N_9410,N_10409);
nand U11698 (N_11698,N_10098,N_9300);
nand U11699 (N_11699,N_10182,N_9179);
and U11700 (N_11700,N_9107,N_10017);
nor U11701 (N_11701,N_9484,N_9930);
or U11702 (N_11702,N_9759,N_10039);
nand U11703 (N_11703,N_9894,N_9435);
and U11704 (N_11704,N_9117,N_9268);
or U11705 (N_11705,N_9021,N_10308);
nor U11706 (N_11706,N_9555,N_9699);
and U11707 (N_11707,N_10357,N_10062);
or U11708 (N_11708,N_9579,N_9043);
or U11709 (N_11709,N_9597,N_10368);
xor U11710 (N_11710,N_9236,N_10287);
or U11711 (N_11711,N_9946,N_10409);
or U11712 (N_11712,N_9585,N_10252);
or U11713 (N_11713,N_10464,N_9687);
nand U11714 (N_11714,N_9242,N_10357);
nor U11715 (N_11715,N_9771,N_10090);
and U11716 (N_11716,N_9568,N_9262);
and U11717 (N_11717,N_9494,N_9655);
nor U11718 (N_11718,N_9341,N_9489);
and U11719 (N_11719,N_9127,N_9689);
and U11720 (N_11720,N_10310,N_9675);
and U11721 (N_11721,N_9846,N_10037);
and U11722 (N_11722,N_10028,N_9902);
nand U11723 (N_11723,N_9529,N_10245);
or U11724 (N_11724,N_9996,N_9911);
nor U11725 (N_11725,N_9645,N_9597);
nor U11726 (N_11726,N_9302,N_9828);
nor U11727 (N_11727,N_10297,N_10030);
nor U11728 (N_11728,N_9262,N_10396);
nor U11729 (N_11729,N_9823,N_9419);
nor U11730 (N_11730,N_10195,N_9342);
nand U11731 (N_11731,N_9352,N_10036);
xnor U11732 (N_11732,N_9057,N_10268);
nand U11733 (N_11733,N_10405,N_9989);
nand U11734 (N_11734,N_10476,N_9041);
and U11735 (N_11735,N_9107,N_10159);
nor U11736 (N_11736,N_10132,N_9418);
nand U11737 (N_11737,N_9636,N_9846);
or U11738 (N_11738,N_9396,N_9475);
and U11739 (N_11739,N_10428,N_9373);
nor U11740 (N_11740,N_9437,N_10343);
nand U11741 (N_11741,N_9163,N_9837);
or U11742 (N_11742,N_9643,N_10458);
nand U11743 (N_11743,N_9959,N_9811);
or U11744 (N_11744,N_10156,N_10406);
or U11745 (N_11745,N_9201,N_9761);
or U11746 (N_11746,N_9659,N_9239);
nor U11747 (N_11747,N_9607,N_10320);
or U11748 (N_11748,N_10198,N_10111);
nand U11749 (N_11749,N_9883,N_9268);
xor U11750 (N_11750,N_9488,N_9476);
or U11751 (N_11751,N_9211,N_10460);
or U11752 (N_11752,N_10088,N_9046);
nand U11753 (N_11753,N_9910,N_10366);
nor U11754 (N_11754,N_9056,N_9794);
nand U11755 (N_11755,N_9876,N_10077);
and U11756 (N_11756,N_10231,N_9056);
xnor U11757 (N_11757,N_9443,N_10336);
xor U11758 (N_11758,N_10302,N_9244);
and U11759 (N_11759,N_9528,N_10057);
and U11760 (N_11760,N_9345,N_10014);
and U11761 (N_11761,N_10275,N_9955);
nand U11762 (N_11762,N_10483,N_10448);
xnor U11763 (N_11763,N_9608,N_10116);
or U11764 (N_11764,N_9409,N_9233);
nand U11765 (N_11765,N_10143,N_9305);
xnor U11766 (N_11766,N_10146,N_9355);
nand U11767 (N_11767,N_9935,N_10083);
and U11768 (N_11768,N_10001,N_9767);
nor U11769 (N_11769,N_9959,N_9146);
nor U11770 (N_11770,N_10128,N_9359);
nand U11771 (N_11771,N_9236,N_9773);
or U11772 (N_11772,N_9145,N_9836);
nor U11773 (N_11773,N_9782,N_9551);
or U11774 (N_11774,N_10499,N_9879);
and U11775 (N_11775,N_10261,N_9414);
and U11776 (N_11776,N_10070,N_10494);
and U11777 (N_11777,N_9528,N_10116);
xor U11778 (N_11778,N_9918,N_10168);
or U11779 (N_11779,N_9250,N_9624);
nand U11780 (N_11780,N_9825,N_9068);
nor U11781 (N_11781,N_9555,N_9171);
nor U11782 (N_11782,N_10233,N_9825);
nand U11783 (N_11783,N_9104,N_9672);
nand U11784 (N_11784,N_9036,N_9668);
xor U11785 (N_11785,N_9622,N_9866);
or U11786 (N_11786,N_9569,N_9801);
nand U11787 (N_11787,N_9621,N_10108);
or U11788 (N_11788,N_9740,N_9316);
nand U11789 (N_11789,N_10373,N_9299);
nand U11790 (N_11790,N_9681,N_9455);
nor U11791 (N_11791,N_9274,N_9444);
nand U11792 (N_11792,N_10202,N_9411);
or U11793 (N_11793,N_10204,N_10197);
and U11794 (N_11794,N_10274,N_10155);
nand U11795 (N_11795,N_9550,N_10358);
xnor U11796 (N_11796,N_9476,N_9494);
nand U11797 (N_11797,N_10022,N_10496);
nand U11798 (N_11798,N_9696,N_9841);
or U11799 (N_11799,N_9735,N_9843);
nor U11800 (N_11800,N_10064,N_9365);
xor U11801 (N_11801,N_10434,N_9354);
or U11802 (N_11802,N_9849,N_9334);
nand U11803 (N_11803,N_9592,N_9667);
nor U11804 (N_11804,N_10275,N_10032);
or U11805 (N_11805,N_9281,N_10204);
or U11806 (N_11806,N_9193,N_9191);
nor U11807 (N_11807,N_9942,N_10212);
nand U11808 (N_11808,N_9083,N_9752);
or U11809 (N_11809,N_9477,N_10131);
and U11810 (N_11810,N_9704,N_9792);
nor U11811 (N_11811,N_9948,N_9973);
or U11812 (N_11812,N_9169,N_9942);
nand U11813 (N_11813,N_10346,N_9491);
and U11814 (N_11814,N_10285,N_9531);
nand U11815 (N_11815,N_10388,N_10081);
or U11816 (N_11816,N_9069,N_9635);
or U11817 (N_11817,N_9984,N_9672);
or U11818 (N_11818,N_9173,N_10011);
nand U11819 (N_11819,N_10009,N_10341);
or U11820 (N_11820,N_9756,N_10237);
and U11821 (N_11821,N_9960,N_9535);
or U11822 (N_11822,N_9504,N_10159);
and U11823 (N_11823,N_9629,N_9900);
or U11824 (N_11824,N_10245,N_9670);
nand U11825 (N_11825,N_10462,N_9372);
nand U11826 (N_11826,N_10364,N_9201);
nand U11827 (N_11827,N_9827,N_10460);
or U11828 (N_11828,N_9503,N_9722);
and U11829 (N_11829,N_9861,N_9335);
nand U11830 (N_11830,N_10172,N_10289);
nor U11831 (N_11831,N_10360,N_9004);
nor U11832 (N_11832,N_9525,N_9791);
or U11833 (N_11833,N_9619,N_9676);
and U11834 (N_11834,N_9095,N_9473);
or U11835 (N_11835,N_9392,N_10139);
nor U11836 (N_11836,N_10154,N_10006);
nand U11837 (N_11837,N_10470,N_9150);
nor U11838 (N_11838,N_10277,N_9072);
and U11839 (N_11839,N_10210,N_10397);
and U11840 (N_11840,N_9823,N_10345);
nor U11841 (N_11841,N_9618,N_9669);
and U11842 (N_11842,N_9907,N_9848);
or U11843 (N_11843,N_9768,N_9347);
nor U11844 (N_11844,N_9096,N_9294);
nor U11845 (N_11845,N_9309,N_10489);
nor U11846 (N_11846,N_10076,N_9774);
nor U11847 (N_11847,N_9522,N_9368);
nand U11848 (N_11848,N_10413,N_9027);
or U11849 (N_11849,N_9477,N_9478);
nand U11850 (N_11850,N_10489,N_9183);
nor U11851 (N_11851,N_9526,N_9141);
nand U11852 (N_11852,N_9781,N_9074);
and U11853 (N_11853,N_10467,N_9899);
or U11854 (N_11854,N_9449,N_10088);
and U11855 (N_11855,N_9915,N_10057);
xor U11856 (N_11856,N_9783,N_9311);
nand U11857 (N_11857,N_9778,N_9129);
nor U11858 (N_11858,N_9949,N_10372);
xor U11859 (N_11859,N_10330,N_9460);
nand U11860 (N_11860,N_9437,N_9519);
and U11861 (N_11861,N_9673,N_9862);
and U11862 (N_11862,N_9660,N_9983);
nand U11863 (N_11863,N_9183,N_9163);
or U11864 (N_11864,N_9442,N_9329);
nand U11865 (N_11865,N_9493,N_9360);
nor U11866 (N_11866,N_10413,N_9555);
nand U11867 (N_11867,N_9187,N_10035);
nor U11868 (N_11868,N_9481,N_9826);
and U11869 (N_11869,N_10300,N_9341);
nand U11870 (N_11870,N_9424,N_10381);
or U11871 (N_11871,N_9712,N_9738);
and U11872 (N_11872,N_9598,N_9738);
or U11873 (N_11873,N_9435,N_9504);
and U11874 (N_11874,N_9261,N_9633);
and U11875 (N_11875,N_9794,N_9768);
nand U11876 (N_11876,N_9052,N_10078);
and U11877 (N_11877,N_10099,N_10304);
nor U11878 (N_11878,N_9411,N_9068);
or U11879 (N_11879,N_10163,N_9305);
nand U11880 (N_11880,N_10315,N_9465);
or U11881 (N_11881,N_10033,N_9611);
xnor U11882 (N_11882,N_9278,N_9971);
or U11883 (N_11883,N_9811,N_9697);
nor U11884 (N_11884,N_9969,N_10287);
nor U11885 (N_11885,N_9694,N_10406);
or U11886 (N_11886,N_9967,N_10032);
or U11887 (N_11887,N_10396,N_10479);
or U11888 (N_11888,N_9533,N_9984);
nor U11889 (N_11889,N_10081,N_9866);
or U11890 (N_11890,N_9477,N_9540);
nor U11891 (N_11891,N_10053,N_10090);
and U11892 (N_11892,N_9989,N_9644);
nand U11893 (N_11893,N_10088,N_9767);
nor U11894 (N_11894,N_10029,N_9676);
nor U11895 (N_11895,N_9371,N_9842);
nor U11896 (N_11896,N_10383,N_9869);
xnor U11897 (N_11897,N_10231,N_9914);
nor U11898 (N_11898,N_10257,N_9147);
and U11899 (N_11899,N_10110,N_9652);
or U11900 (N_11900,N_9884,N_9252);
nand U11901 (N_11901,N_9808,N_9172);
or U11902 (N_11902,N_9262,N_9396);
nor U11903 (N_11903,N_10142,N_9070);
nor U11904 (N_11904,N_10198,N_9301);
and U11905 (N_11905,N_9863,N_10344);
nand U11906 (N_11906,N_9912,N_10089);
nor U11907 (N_11907,N_9322,N_9676);
nor U11908 (N_11908,N_9122,N_9633);
and U11909 (N_11909,N_9046,N_9498);
and U11910 (N_11910,N_9993,N_9069);
and U11911 (N_11911,N_9943,N_9093);
and U11912 (N_11912,N_10292,N_9577);
nor U11913 (N_11913,N_10306,N_9103);
and U11914 (N_11914,N_10346,N_9565);
and U11915 (N_11915,N_9586,N_10107);
or U11916 (N_11916,N_9518,N_10447);
nand U11917 (N_11917,N_9454,N_9848);
or U11918 (N_11918,N_9523,N_10290);
and U11919 (N_11919,N_10127,N_9009);
nor U11920 (N_11920,N_9866,N_10494);
nor U11921 (N_11921,N_9570,N_10042);
nor U11922 (N_11922,N_9313,N_9168);
nand U11923 (N_11923,N_9447,N_10072);
or U11924 (N_11924,N_9577,N_9707);
nor U11925 (N_11925,N_10293,N_9594);
nand U11926 (N_11926,N_9506,N_9355);
or U11927 (N_11927,N_10480,N_10207);
xnor U11928 (N_11928,N_9588,N_9917);
nand U11929 (N_11929,N_9003,N_9509);
nor U11930 (N_11930,N_9436,N_9898);
and U11931 (N_11931,N_9906,N_9963);
nand U11932 (N_11932,N_9156,N_10310);
xnor U11933 (N_11933,N_9357,N_10370);
and U11934 (N_11934,N_10162,N_9575);
or U11935 (N_11935,N_9736,N_9807);
and U11936 (N_11936,N_9989,N_10085);
or U11937 (N_11937,N_10462,N_10129);
nand U11938 (N_11938,N_9036,N_9938);
nor U11939 (N_11939,N_9754,N_10179);
and U11940 (N_11940,N_9282,N_10450);
and U11941 (N_11941,N_9278,N_9566);
or U11942 (N_11942,N_9043,N_9328);
nor U11943 (N_11943,N_9252,N_10146);
and U11944 (N_11944,N_10412,N_9276);
and U11945 (N_11945,N_9106,N_10184);
nor U11946 (N_11946,N_9417,N_9393);
nand U11947 (N_11947,N_9779,N_9558);
or U11948 (N_11948,N_9305,N_9228);
xor U11949 (N_11949,N_9150,N_9382);
nor U11950 (N_11950,N_9119,N_9398);
or U11951 (N_11951,N_9814,N_9637);
xor U11952 (N_11952,N_9913,N_10472);
nand U11953 (N_11953,N_9177,N_10120);
or U11954 (N_11954,N_9299,N_10490);
nand U11955 (N_11955,N_10448,N_9892);
or U11956 (N_11956,N_10317,N_10196);
xnor U11957 (N_11957,N_9942,N_9307);
and U11958 (N_11958,N_10283,N_10123);
nor U11959 (N_11959,N_9923,N_9932);
nand U11960 (N_11960,N_10275,N_9271);
nand U11961 (N_11961,N_9244,N_9483);
and U11962 (N_11962,N_9223,N_9593);
or U11963 (N_11963,N_9787,N_9832);
nand U11964 (N_11964,N_10234,N_10211);
nand U11965 (N_11965,N_9460,N_9393);
nand U11966 (N_11966,N_9470,N_9852);
and U11967 (N_11967,N_9616,N_9388);
nand U11968 (N_11968,N_10082,N_9513);
nor U11969 (N_11969,N_9514,N_10466);
nor U11970 (N_11970,N_10031,N_9331);
and U11971 (N_11971,N_10280,N_9936);
or U11972 (N_11972,N_9114,N_10391);
nor U11973 (N_11973,N_9934,N_9859);
or U11974 (N_11974,N_9940,N_9514);
xnor U11975 (N_11975,N_10178,N_10190);
nand U11976 (N_11976,N_9328,N_9175);
nand U11977 (N_11977,N_10124,N_10092);
or U11978 (N_11978,N_9906,N_10119);
xnor U11979 (N_11979,N_10285,N_10343);
or U11980 (N_11980,N_9374,N_9261);
and U11981 (N_11981,N_10467,N_9523);
or U11982 (N_11982,N_10181,N_10400);
and U11983 (N_11983,N_9429,N_9063);
xor U11984 (N_11984,N_9446,N_9799);
xnor U11985 (N_11985,N_9965,N_10022);
xor U11986 (N_11986,N_9337,N_10406);
and U11987 (N_11987,N_10073,N_10107);
nand U11988 (N_11988,N_9826,N_9087);
xnor U11989 (N_11989,N_9330,N_10241);
and U11990 (N_11990,N_10156,N_10423);
nand U11991 (N_11991,N_9186,N_10436);
or U11992 (N_11992,N_9055,N_10239);
nand U11993 (N_11993,N_9026,N_10143);
or U11994 (N_11994,N_10254,N_9377);
nand U11995 (N_11995,N_10247,N_10042);
or U11996 (N_11996,N_9960,N_9216);
nor U11997 (N_11997,N_9252,N_9954);
and U11998 (N_11998,N_10034,N_10474);
nor U11999 (N_11999,N_9738,N_9528);
xnor U12000 (N_12000,N_11537,N_11693);
or U12001 (N_12001,N_10679,N_11869);
and U12002 (N_12002,N_11302,N_11007);
nand U12003 (N_12003,N_11996,N_11492);
or U12004 (N_12004,N_10634,N_10862);
nor U12005 (N_12005,N_10536,N_11541);
nor U12006 (N_12006,N_11001,N_10906);
or U12007 (N_12007,N_11150,N_10603);
nor U12008 (N_12008,N_11810,N_10855);
xnor U12009 (N_12009,N_11061,N_11047);
nor U12010 (N_12010,N_10509,N_11963);
or U12011 (N_12011,N_10578,N_10973);
and U12012 (N_12012,N_11742,N_11057);
and U12013 (N_12013,N_10954,N_11507);
or U12014 (N_12014,N_10826,N_11257);
or U12015 (N_12015,N_11465,N_11657);
and U12016 (N_12016,N_11813,N_11382);
or U12017 (N_12017,N_11448,N_11484);
and U12018 (N_12018,N_11571,N_11972);
xnor U12019 (N_12019,N_10733,N_10922);
and U12020 (N_12020,N_11032,N_11591);
nor U12021 (N_12021,N_10763,N_11982);
and U12022 (N_12022,N_11539,N_11493);
and U12023 (N_12023,N_11974,N_11727);
nand U12024 (N_12024,N_11383,N_11169);
xor U12025 (N_12025,N_10622,N_11654);
nand U12026 (N_12026,N_11311,N_11845);
and U12027 (N_12027,N_11512,N_11253);
nand U12028 (N_12028,N_11337,N_11165);
nor U12029 (N_12029,N_10769,N_10527);
nor U12030 (N_12030,N_11538,N_11917);
nand U12031 (N_12031,N_11044,N_11503);
nand U12032 (N_12032,N_11937,N_11413);
nand U12033 (N_12033,N_11981,N_10682);
nor U12034 (N_12034,N_11264,N_11475);
nor U12035 (N_12035,N_11569,N_10939);
nor U12036 (N_12036,N_11714,N_11216);
and U12037 (N_12037,N_11901,N_10550);
nor U12038 (N_12038,N_10932,N_11780);
nand U12039 (N_12039,N_10976,N_10827);
nor U12040 (N_12040,N_10684,N_10705);
or U12041 (N_12041,N_11035,N_11928);
nand U12042 (N_12042,N_11091,N_11243);
and U12043 (N_12043,N_11862,N_11325);
nor U12044 (N_12044,N_11868,N_11580);
nor U12045 (N_12045,N_11707,N_11694);
and U12046 (N_12046,N_11348,N_10978);
or U12047 (N_12047,N_10800,N_10895);
nand U12048 (N_12048,N_11902,N_10598);
nand U12049 (N_12049,N_10689,N_11432);
xor U12050 (N_12050,N_10723,N_11685);
or U12051 (N_12051,N_10729,N_10822);
nand U12052 (N_12052,N_10866,N_11676);
and U12053 (N_12053,N_10890,N_11523);
nor U12054 (N_12054,N_10852,N_11343);
xnor U12055 (N_12055,N_11418,N_10905);
nor U12056 (N_12056,N_11596,N_11369);
nor U12057 (N_12057,N_11883,N_11679);
nor U12058 (N_12058,N_11396,N_11684);
nand U12059 (N_12059,N_10628,N_11565);
nand U12060 (N_12060,N_11765,N_11556);
xnor U12061 (N_12061,N_10882,N_11345);
nor U12062 (N_12062,N_10874,N_11313);
or U12063 (N_12063,N_11612,N_11763);
nor U12064 (N_12064,N_10853,N_10685);
nor U12065 (N_12065,N_11147,N_11158);
nand U12066 (N_12066,N_10668,N_11162);
nand U12067 (N_12067,N_11808,N_11701);
or U12068 (N_12068,N_10728,N_11255);
and U12069 (N_12069,N_10957,N_10662);
nand U12070 (N_12070,N_11796,N_11910);
or U12071 (N_12071,N_11244,N_10879);
or U12072 (N_12072,N_10665,N_11856);
nand U12073 (N_12073,N_11398,N_11823);
and U12074 (N_12074,N_11951,N_10540);
or U12075 (N_12075,N_10572,N_10519);
and U12076 (N_12076,N_11485,N_10580);
nor U12077 (N_12077,N_11745,N_10927);
nor U12078 (N_12078,N_11127,N_11985);
nor U12079 (N_12079,N_11578,N_11043);
and U12080 (N_12080,N_10907,N_10664);
and U12081 (N_12081,N_11460,N_11561);
and U12082 (N_12082,N_11277,N_10865);
nor U12083 (N_12083,N_10696,N_10570);
nand U12084 (N_12084,N_11399,N_10576);
nor U12085 (N_12085,N_11378,N_11582);
xor U12086 (N_12086,N_11852,N_11599);
and U12087 (N_12087,N_11752,N_11078);
or U12088 (N_12088,N_10507,N_11124);
and U12089 (N_12089,N_10913,N_11833);
nand U12090 (N_12090,N_11254,N_11074);
and U12091 (N_12091,N_10697,N_11611);
xnor U12092 (N_12092,N_10500,N_11024);
nand U12093 (N_12093,N_11228,N_11093);
and U12094 (N_12094,N_11584,N_10633);
nand U12095 (N_12095,N_11370,N_11342);
nand U12096 (N_12096,N_10746,N_11853);
nand U12097 (N_12097,N_10611,N_10673);
xnor U12098 (N_12098,N_10641,N_11719);
nor U12099 (N_12099,N_10702,N_11242);
and U12100 (N_12100,N_11712,N_11510);
nor U12101 (N_12101,N_11638,N_10864);
xnor U12102 (N_12102,N_10991,N_10845);
nand U12103 (N_12103,N_10715,N_10678);
nand U12104 (N_12104,N_10716,N_10885);
or U12105 (N_12105,N_10686,N_10860);
xnor U12106 (N_12106,N_11774,N_11529);
nor U12107 (N_12107,N_10695,N_10876);
or U12108 (N_12108,N_11881,N_10599);
or U12109 (N_12109,N_11675,N_10902);
nand U12110 (N_12110,N_10815,N_11106);
nand U12111 (N_12111,N_11291,N_11923);
and U12112 (N_12112,N_11112,N_11490);
and U12113 (N_12113,N_10887,N_10900);
nor U12114 (N_12114,N_11543,N_11049);
nor U12115 (N_12115,N_11177,N_10960);
nor U12116 (N_12116,N_11632,N_11247);
nand U12117 (N_12117,N_11394,N_11802);
and U12118 (N_12118,N_11170,N_10805);
and U12119 (N_12119,N_11986,N_11117);
xor U12120 (N_12120,N_11748,N_11933);
or U12121 (N_12121,N_10501,N_11831);
and U12122 (N_12122,N_10640,N_11705);
nor U12123 (N_12123,N_11240,N_11308);
nand U12124 (N_12124,N_11773,N_11161);
and U12125 (N_12125,N_10972,N_11900);
nor U12126 (N_12126,N_10787,N_11027);
nor U12127 (N_12127,N_11740,N_10595);
nor U12128 (N_12128,N_10713,N_11518);
and U12129 (N_12129,N_11155,N_11878);
or U12130 (N_12130,N_11843,N_11662);
nor U12131 (N_12131,N_11689,N_11948);
nor U12132 (N_12132,N_11906,N_10796);
and U12133 (N_12133,N_11703,N_10940);
or U12134 (N_12134,N_11559,N_11055);
nor U12135 (N_12135,N_11410,N_11022);
and U12136 (N_12136,N_11659,N_10581);
or U12137 (N_12137,N_11011,N_11272);
nand U12138 (N_12138,N_10765,N_11767);
xnor U12139 (N_12139,N_11588,N_11251);
nor U12140 (N_12140,N_11889,N_11809);
or U12141 (N_12141,N_11952,N_11961);
xnor U12142 (N_12142,N_11290,N_10745);
nor U12143 (N_12143,N_11445,N_10571);
and U12144 (N_12144,N_10961,N_11614);
nor U12145 (N_12145,N_11229,N_11674);
and U12146 (N_12146,N_11141,N_11506);
and U12147 (N_12147,N_10620,N_10680);
xor U12148 (N_12148,N_11927,N_11930);
and U12149 (N_12149,N_11099,N_10828);
nand U12150 (N_12150,N_11704,N_10893);
and U12151 (N_12151,N_11971,N_11605);
and U12152 (N_12152,N_11407,N_10513);
and U12153 (N_12153,N_11286,N_11877);
nand U12154 (N_12154,N_11871,N_11083);
nand U12155 (N_12155,N_10968,N_10937);
xnor U12156 (N_12156,N_11756,N_11620);
or U12157 (N_12157,N_11395,N_10647);
nor U12158 (N_12158,N_10766,N_11747);
or U12159 (N_12159,N_10962,N_11608);
xnor U12160 (N_12160,N_10761,N_10969);
and U12161 (N_12161,N_10677,N_11594);
or U12162 (N_12162,N_11235,N_10943);
and U12163 (N_12163,N_11603,N_11534);
nand U12164 (N_12164,N_11459,N_11371);
nand U12165 (N_12165,N_10808,N_11281);
or U12166 (N_12166,N_10514,N_11716);
nor U12167 (N_12167,N_11696,N_11664);
or U12168 (N_12168,N_10672,N_11860);
and U12169 (N_12169,N_11002,N_10614);
and U12170 (N_12170,N_11838,N_11331);
and U12171 (N_12171,N_10639,N_11914);
xor U12172 (N_12172,N_10706,N_11230);
or U12173 (N_12173,N_11820,N_10574);
and U12174 (N_12174,N_11516,N_11895);
or U12175 (N_12175,N_11783,N_11922);
and U12176 (N_12176,N_10825,N_11225);
and U12177 (N_12177,N_11393,N_11785);
and U12178 (N_12178,N_10789,N_11304);
nor U12179 (N_12179,N_11129,N_11320);
or U12180 (N_12180,N_11790,N_11275);
nor U12181 (N_12181,N_11893,N_11289);
nor U12182 (N_12182,N_10583,N_11522);
nand U12183 (N_12183,N_11202,N_11573);
nor U12184 (N_12184,N_10607,N_10989);
nor U12185 (N_12185,N_10594,N_11096);
nand U12186 (N_12186,N_11233,N_10621);
nand U12187 (N_12187,N_11652,N_10916);
and U12188 (N_12188,N_11646,N_11904);
nand U12189 (N_12189,N_10503,N_10608);
xnor U12190 (N_12190,N_10924,N_10644);
or U12191 (N_12191,N_11265,N_11363);
nand U12192 (N_12192,N_10707,N_11958);
nand U12193 (N_12193,N_10901,N_10833);
or U12194 (N_12194,N_11786,N_11212);
or U12195 (N_12195,N_10563,N_10667);
xnor U12196 (N_12196,N_11000,N_11444);
nor U12197 (N_12197,N_11322,N_10749);
nand U12198 (N_12198,N_10836,N_11208);
or U12199 (N_12199,N_11306,N_10824);
xor U12200 (N_12200,N_11550,N_11113);
or U12201 (N_12201,N_10688,N_10889);
or U12202 (N_12202,N_11065,N_11944);
xnor U12203 (N_12203,N_11069,N_11172);
and U12204 (N_12204,N_11143,N_10784);
nand U12205 (N_12205,N_10711,N_10632);
or U12206 (N_12206,N_10791,N_11200);
and U12207 (N_12207,N_10588,N_11915);
or U12208 (N_12208,N_10929,N_10502);
nor U12209 (N_12209,N_11692,N_11521);
or U12210 (N_12210,N_11419,N_11181);
nand U12211 (N_12211,N_11204,N_10987);
nor U12212 (N_12212,N_11339,N_11688);
nand U12213 (N_12213,N_10870,N_11734);
nand U12214 (N_12214,N_11495,N_11451);
or U12215 (N_12215,N_11458,N_11126);
and U12216 (N_12216,N_11417,N_11630);
nor U12217 (N_12217,N_11139,N_10859);
nand U12218 (N_12218,N_11649,N_10670);
and U12219 (N_12219,N_11333,N_10949);
nor U12220 (N_12220,N_11103,N_11332);
nor U12221 (N_12221,N_11054,N_10575);
or U12222 (N_12222,N_11666,N_10528);
nand U12223 (N_12223,N_11822,N_11837);
nand U12224 (N_12224,N_10760,N_10935);
xnor U12225 (N_12225,N_10966,N_10704);
and U12226 (N_12226,N_11669,N_10835);
and U12227 (N_12227,N_11248,N_10963);
nor U12228 (N_12228,N_11353,N_11759);
or U12229 (N_12229,N_10510,N_11939);
and U12230 (N_12230,N_11108,N_10653);
and U12231 (N_12231,N_11135,N_11076);
and U12232 (N_12232,N_11387,N_10521);
nor U12233 (N_12233,N_11344,N_11048);
or U12234 (N_12234,N_10810,N_11803);
nand U12235 (N_12235,N_11520,N_10964);
and U12236 (N_12236,N_10854,N_10892);
and U12237 (N_12237,N_11564,N_11287);
xnor U12238 (N_12238,N_11077,N_11566);
nand U12239 (N_12239,N_10559,N_10910);
nand U12240 (N_12240,N_10525,N_11633);
and U12241 (N_12241,N_11142,N_11373);
and U12242 (N_12242,N_11995,N_11016);
nor U12243 (N_12243,N_11372,N_10798);
and U12244 (N_12244,N_10947,N_11595);
or U12245 (N_12245,N_11245,N_10736);
xnor U12246 (N_12246,N_10617,N_11966);
nor U12247 (N_12247,N_11825,N_11136);
and U12248 (N_12248,N_10631,N_10731);
nand U12249 (N_12249,N_11408,N_11454);
xnor U12250 (N_12250,N_10857,N_11514);
xnor U12251 (N_12251,N_11766,N_11532);
nand U12252 (N_12252,N_10856,N_10681);
nand U12253 (N_12253,N_10817,N_10524);
nand U12254 (N_12254,N_10867,N_11979);
nor U12255 (N_12255,N_10593,N_11690);
nand U12256 (N_12256,N_10983,N_11658);
and U12257 (N_12257,N_10561,N_10586);
or U12258 (N_12258,N_10752,N_11660);
nor U12259 (N_12259,N_10814,N_10661);
and U12260 (N_12260,N_11513,N_11872);
nor U12261 (N_12261,N_11366,N_11384);
nand U12262 (N_12262,N_11184,N_10714);
nor U12263 (N_12263,N_11997,N_10584);
nor U12264 (N_12264,N_10650,N_11056);
or U12265 (N_12265,N_11653,N_11462);
nand U12266 (N_12266,N_11051,N_10657);
or U12267 (N_12267,N_11029,N_11897);
nand U12268 (N_12268,N_11480,N_11467);
xnor U12269 (N_12269,N_11310,N_11730);
nand U12270 (N_12270,N_11975,N_11307);
nor U12271 (N_12271,N_11101,N_11953);
nand U12272 (N_12272,N_10930,N_11179);
nand U12273 (N_12273,N_11583,N_10786);
xnor U12274 (N_12274,N_11806,N_10975);
or U12275 (N_12275,N_10844,N_10724);
xor U12276 (N_12276,N_10693,N_11683);
nor U12277 (N_12277,N_11945,N_10602);
or U12278 (N_12278,N_11214,N_11597);
and U12279 (N_12279,N_11270,N_11918);
and U12280 (N_12280,N_11711,N_10629);
nor U12281 (N_12281,N_10651,N_11764);
nand U12282 (N_12282,N_10819,N_11138);
xor U12283 (N_12283,N_11315,N_11435);
or U12284 (N_12284,N_10720,N_11992);
or U12285 (N_12285,N_11262,N_11062);
nor U12286 (N_12286,N_11585,N_11284);
nand U12287 (N_12287,N_10881,N_10535);
nor U12288 (N_12288,N_11028,N_11779);
nor U12289 (N_12289,N_11505,N_11560);
nand U12290 (N_12290,N_10549,N_11276);
nor U12291 (N_12291,N_11601,N_11402);
and U12292 (N_12292,N_11196,N_11053);
xnor U12293 (N_12293,N_11544,N_11386);
nand U12294 (N_12294,N_11776,N_11104);
or U12295 (N_12295,N_11227,N_11328);
nor U12296 (N_12296,N_11224,N_11496);
nor U12297 (N_12297,N_11125,N_10750);
and U12298 (N_12298,N_11105,N_11645);
nor U12299 (N_12299,N_10532,N_11610);
or U12300 (N_12300,N_11964,N_11088);
and U12301 (N_12301,N_10625,N_10596);
nand U12302 (N_12302,N_10872,N_11526);
xnor U12303 (N_12303,N_11536,N_11535);
nand U12304 (N_12304,N_11613,N_10839);
nand U12305 (N_12305,N_10911,N_10623);
or U12306 (N_12306,N_11941,N_10624);
nand U12307 (N_12307,N_10795,N_11206);
nor U12308 (N_12308,N_11469,N_11215);
and U12309 (N_12309,N_10908,N_11401);
or U12310 (N_12310,N_11361,N_11625);
nand U12311 (N_12311,N_11163,N_10952);
nand U12312 (N_12312,N_11167,N_10708);
nor U12313 (N_12313,N_11892,N_11587);
nand U12314 (N_12314,N_11487,N_11725);
nor U12315 (N_12315,N_10547,N_10558);
or U12316 (N_12316,N_10601,N_10831);
nand U12317 (N_12317,N_11033,N_11626);
or U12318 (N_12318,N_11152,N_11699);
and U12319 (N_12319,N_11807,N_11440);
nand U12320 (N_12320,N_11661,N_11183);
or U12321 (N_12321,N_11651,N_10508);
and U12322 (N_12322,N_11846,N_10888);
and U12323 (N_12323,N_11221,N_11994);
nor U12324 (N_12324,N_10884,N_11470);
nand U12325 (N_12325,N_10850,N_10703);
nand U12326 (N_12326,N_11477,N_10829);
xnor U12327 (N_12327,N_11488,N_11947);
xor U12328 (N_12328,N_11874,N_10871);
or U12329 (N_12329,N_11085,N_11118);
nand U12330 (N_12330,N_10959,N_10544);
xor U12331 (N_12331,N_11644,N_11086);
nand U12332 (N_12332,N_11187,N_10868);
or U12333 (N_12333,N_11935,N_11882);
or U12334 (N_12334,N_10951,N_10912);
nor U12335 (N_12335,N_10861,N_11973);
or U12336 (N_12336,N_10812,N_10515);
nand U12337 (N_12337,N_11362,N_11607);
xor U12338 (N_12338,N_11801,N_11358);
xor U12339 (N_12339,N_11301,N_11347);
nor U12340 (N_12340,N_11884,N_11282);
or U12341 (N_12341,N_11864,N_10757);
nor U12342 (N_12342,N_10873,N_11030);
nor U12343 (N_12343,N_10880,N_10582);
or U12344 (N_12344,N_11025,N_10569);
or U12345 (N_12345,N_10565,N_11412);
or U12346 (N_12346,N_11377,N_11060);
and U12347 (N_12347,N_11319,N_10663);
nor U12348 (N_12348,N_11406,N_11102);
or U12349 (N_12349,N_11524,N_11197);
and U12350 (N_12350,N_11473,N_11530);
and U12351 (N_12351,N_11075,N_10683);
and U12352 (N_12352,N_10774,N_11844);
nor U12353 (N_12353,N_10919,N_10666);
nand U12354 (N_12354,N_10698,N_11346);
and U12355 (N_12355,N_10701,N_11068);
and U12356 (N_12356,N_10654,N_11762);
nor U12357 (N_12357,N_11008,N_11794);
nand U12358 (N_12358,N_11489,N_11283);
nor U12359 (N_12359,N_10778,N_11017);
and U12360 (N_12360,N_11443,N_11671);
nor U12361 (N_12361,N_11191,N_10807);
or U12362 (N_12362,N_11080,N_10899);
and U12363 (N_12363,N_11154,N_11219);
and U12364 (N_12364,N_11005,N_10556);
and U12365 (N_12365,N_11134,N_10655);
xnor U12366 (N_12366,N_11555,N_11799);
nand U12367 (N_12367,N_11702,N_11781);
nand U12368 (N_12368,N_11950,N_11157);
and U12369 (N_12369,N_10981,N_11640);
nand U12370 (N_12370,N_11380,N_11122);
xnor U12371 (N_12371,N_10504,N_10838);
nor U12372 (N_12372,N_10539,N_10938);
and U12373 (N_12373,N_11226,N_10554);
and U12374 (N_12374,N_11405,N_11317);
nand U12375 (N_12375,N_11411,N_11357);
xor U12376 (N_12376,N_11873,N_11217);
or U12377 (N_12377,N_11772,N_10587);
nor U12378 (N_12378,N_10591,N_11929);
nor U12379 (N_12379,N_11153,N_10782);
nand U12380 (N_12380,N_11903,N_11334);
nor U12381 (N_12381,N_11811,N_11542);
nand U12382 (N_12382,N_10771,N_11617);
nand U12383 (N_12383,N_11084,N_11720);
nand U12384 (N_12384,N_11115,N_11335);
xor U12385 (N_12385,N_10636,N_11144);
or U12386 (N_12386,N_11107,N_10643);
nor U12387 (N_12387,N_11563,N_11977);
xor U12388 (N_12388,N_11241,N_11842);
nand U12389 (N_12389,N_10725,N_10883);
nand U12390 (N_12390,N_11857,N_11744);
or U12391 (N_12391,N_10649,N_10538);
nor U12392 (N_12392,N_11549,N_11800);
nand U12393 (N_12393,N_11554,N_11887);
and U12394 (N_12394,N_11476,N_10573);
or U12395 (N_12395,N_11851,N_11092);
nor U12396 (N_12396,N_10646,N_11305);
and U12397 (N_12397,N_10506,N_11274);
or U12398 (N_12398,N_11111,N_11920);
xor U12399 (N_12399,N_10970,N_11483);
nor U12400 (N_12400,N_10917,N_11285);
and U12401 (N_12401,N_10553,N_10523);
and U12402 (N_12402,N_11379,N_10891);
or U12403 (N_12403,N_11899,N_10762);
nor U12404 (N_12404,N_11680,N_11618);
xor U12405 (N_12405,N_11097,N_11604);
nand U12406 (N_12406,N_10710,N_11968);
or U12407 (N_12407,N_10546,N_11193);
nor U12408 (N_12408,N_11998,N_11294);
nor U12409 (N_12409,N_10904,N_11804);
nor U12410 (N_12410,N_11830,N_10590);
nand U12411 (N_12411,N_11231,N_10609);
nand U12412 (N_12412,N_11098,N_11623);
xnor U12413 (N_12413,N_11858,N_10942);
or U12414 (N_12414,N_11050,N_11976);
nand U12415 (N_12415,N_10718,N_11354);
nand U12416 (N_12416,N_11461,N_11970);
or U12417 (N_12417,N_11014,N_10747);
nor U12418 (N_12418,N_11246,N_11066);
xnor U12419 (N_12419,N_10877,N_11237);
nand U12420 (N_12420,N_10744,N_11898);
nand U12421 (N_12421,N_10985,N_10896);
and U12422 (N_12422,N_10635,N_11643);
nor U12423 (N_12423,N_11441,N_11558);
xor U12424 (N_12424,N_11295,N_11736);
xnor U12425 (N_12425,N_11905,N_11203);
or U12426 (N_12426,N_11672,N_11751);
nor U12427 (N_12427,N_11722,N_11156);
or U12428 (N_12428,N_10903,N_10886);
or U12429 (N_12429,N_10564,N_10505);
and U12430 (N_12430,N_10548,N_11501);
nand U12431 (N_12431,N_11464,N_10996);
and U12432 (N_12432,N_11252,N_11504);
and U12433 (N_12433,N_11389,N_11708);
or U12434 (N_12434,N_11743,N_11637);
nor U12435 (N_12435,N_11416,N_11567);
and U12436 (N_12436,N_11700,N_10699);
and U12437 (N_12437,N_11999,N_11223);
nand U12438 (N_12438,N_11816,N_11656);
nor U12439 (N_12439,N_11040,N_11616);
and U12440 (N_12440,N_11349,N_11123);
xnor U12441 (N_12441,N_11186,N_11168);
xnor U12442 (N_12442,N_10648,N_11983);
nand U12443 (N_12443,N_11450,N_10980);
and U12444 (N_12444,N_11797,N_10770);
xnor U12445 (N_12445,N_10915,N_11052);
and U12446 (N_12446,N_11886,N_11201);
nand U12447 (N_12447,N_11385,N_11499);
or U12448 (N_12448,N_11481,N_11414);
nor U12449 (N_12449,N_11042,N_11758);
nand U12450 (N_12450,N_11374,N_11434);
or U12451 (N_12451,N_10619,N_11913);
or U12452 (N_12452,N_11258,N_11427);
or U12453 (N_12453,N_10530,N_11222);
and U12454 (N_12454,N_11525,N_10560);
and U12455 (N_12455,N_11280,N_11479);
or U12456 (N_12456,N_10792,N_11815);
or U12457 (N_12457,N_10990,N_10753);
nand U12458 (N_12458,N_10848,N_11073);
nand U12459 (N_12459,N_11909,N_11321);
nor U12460 (N_12460,N_11238,N_11236);
nand U12461 (N_12461,N_11261,N_11159);
and U12462 (N_12462,N_10933,N_10537);
nand U12463 (N_12463,N_11148,N_11404);
and U12464 (N_12464,N_11207,N_11557);
or U12465 (N_12465,N_11424,N_11463);
or U12466 (N_12466,N_11628,N_11859);
or U12467 (N_12467,N_10652,N_10567);
nand U12468 (N_12468,N_11121,N_10982);
or U12469 (N_12469,N_11409,N_11494);
nor U12470 (N_12470,N_10818,N_10984);
or U12471 (N_12471,N_10656,N_11515);
xnor U12472 (N_12472,N_11826,N_11647);
and U12473 (N_12473,N_11213,N_11593);
and U12474 (N_12474,N_11400,N_10604);
and U12475 (N_12475,N_10790,N_11021);
or U12476 (N_12476,N_10743,N_11425);
nor U12477 (N_12477,N_10605,N_10944);
or U12478 (N_12478,N_10722,N_11063);
nand U12479 (N_12479,N_11698,N_11619);
xnor U12480 (N_12480,N_11205,N_11581);
or U12481 (N_12481,N_10734,N_10803);
nor U12482 (N_12482,N_10977,N_11891);
and U12483 (N_12483,N_11792,N_10780);
nor U12484 (N_12484,N_10909,N_10717);
nor U12485 (N_12485,N_10645,N_10566);
or U12486 (N_12486,N_11273,N_11256);
nand U12487 (N_12487,N_10709,N_10858);
nand U12488 (N_12488,N_11771,N_11834);
or U12489 (N_12489,N_11749,N_11218);
xor U12490 (N_12490,N_10785,N_11015);
nand U12491 (N_12491,N_11486,N_11472);
and U12492 (N_12492,N_11729,N_10783);
and U12493 (N_12493,N_11634,N_11220);
and U12494 (N_12494,N_11036,N_10687);
or U12495 (N_12495,N_11038,N_11828);
nor U12496 (N_12496,N_10869,N_11880);
and U12497 (N_12497,N_11896,N_10941);
nor U12498 (N_12498,N_11491,N_11376);
nand U12499 (N_12499,N_11735,N_11519);
xor U12500 (N_12500,N_10920,N_11166);
and U12501 (N_12501,N_10511,N_10998);
nand U12502 (N_12502,N_10759,N_11131);
nor U12503 (N_12503,N_11706,N_11436);
nor U12504 (N_12504,N_10742,N_11787);
nor U12505 (N_12505,N_11314,N_11188);
or U12506 (N_12506,N_11171,N_11137);
nor U12507 (N_12507,N_10799,N_11990);
and U12508 (N_12508,N_11840,N_10545);
and U12509 (N_12509,N_10950,N_11733);
and U12510 (N_12510,N_10526,N_11368);
xnor U12511 (N_12511,N_10543,N_10847);
and U12512 (N_12512,N_10552,N_11836);
nor U12513 (N_12513,N_11962,N_10531);
nand U12514 (N_12514,N_10764,N_11854);
or U12515 (N_12515,N_11266,N_11020);
xor U12516 (N_12516,N_11791,N_11439);
or U12517 (N_12517,N_11279,N_11867);
nor U12518 (N_12518,N_11728,N_11079);
nand U12519 (N_12519,N_10712,N_11814);
nor U12520 (N_12520,N_11110,N_10613);
nor U12521 (N_12521,N_11827,N_10863);
xnor U12522 (N_12522,N_10809,N_11012);
nor U12523 (N_12523,N_11013,N_11303);
and U12524 (N_12524,N_11081,N_11919);
nand U12525 (N_12525,N_11004,N_11509);
and U12526 (N_12526,N_11798,N_10627);
and U12527 (N_12527,N_10562,N_10926);
or U12528 (N_12528,N_10557,N_11648);
nand U12529 (N_12529,N_11232,N_11789);
nor U12530 (N_12530,N_10995,N_11039);
nor U12531 (N_12531,N_11821,N_11949);
or U12532 (N_12532,N_11466,N_11936);
and U12533 (N_12533,N_11397,N_11782);
nor U12534 (N_12534,N_11511,N_10658);
nor U12535 (N_12535,N_11760,N_11849);
nand U12536 (N_12536,N_11009,N_10755);
and U12537 (N_12537,N_11269,N_10737);
nor U12538 (N_12538,N_10914,N_11297);
or U12539 (N_12539,N_11352,N_11655);
and U12540 (N_12540,N_11540,N_11456);
or U12541 (N_12541,N_11978,N_11433);
xnor U12542 (N_12542,N_11932,N_10974);
and U12543 (N_12543,N_11602,N_10691);
and U12544 (N_12544,N_11090,N_11145);
or U12545 (N_12545,N_11064,N_11442);
nand U12546 (N_12546,N_11931,N_11318);
nor U12547 (N_12547,N_11691,N_10842);
or U12548 (N_12548,N_10597,N_11180);
nand U12549 (N_12549,N_10776,N_10732);
or U12550 (N_12550,N_11635,N_11908);
and U12551 (N_12551,N_10637,N_11775);
xnor U12552 (N_12552,N_11114,N_11641);
xnor U12553 (N_12553,N_11551,N_10801);
and U12554 (N_12554,N_11817,N_11754);
and U12555 (N_12555,N_11907,N_10659);
and U12556 (N_12556,N_11839,N_11336);
nor U12557 (N_12557,N_11575,N_10956);
or U12558 (N_12558,N_11642,N_11446);
or U12559 (N_12559,N_10541,N_11210);
or U12560 (N_12560,N_11673,N_11316);
nand U12561 (N_12561,N_11431,N_11682);
and U12562 (N_12562,N_10754,N_11453);
or U12563 (N_12563,N_11726,N_10946);
and U12564 (N_12564,N_11631,N_11710);
nor U12565 (N_12565,N_11323,N_11130);
nor U12566 (N_12566,N_11173,N_11967);
nand U12567 (N_12567,N_10965,N_11709);
nor U12568 (N_12568,N_10520,N_10804);
or U12569 (N_12569,N_10630,N_11579);
nor U12570 (N_12570,N_10577,N_11500);
or U12571 (N_12571,N_11006,N_11211);
nand U12572 (N_12572,N_11375,N_11023);
and U12573 (N_12573,N_10832,N_11681);
nor U12574 (N_12574,N_10788,N_11422);
nand U12575 (N_12575,N_10589,N_11421);
or U12576 (N_12576,N_11959,N_11003);
or U12577 (N_12577,N_10739,N_10726);
nand U12578 (N_12578,N_10758,N_11768);
or U12579 (N_12579,N_11070,N_11769);
nor U12580 (N_12580,N_11082,N_10542);
nand U12581 (N_12581,N_11697,N_11570);
nor U12582 (N_12582,N_10606,N_11732);
nand U12583 (N_12583,N_11824,N_11589);
and U12584 (N_12584,N_10875,N_10534);
xnor U12585 (N_12585,N_10529,N_11890);
or U12586 (N_12586,N_10994,N_11474);
xor U12587 (N_12587,N_11943,N_11568);
and U12588 (N_12588,N_11478,N_11058);
nor U12589 (N_12589,N_11312,N_11546);
nand U12590 (N_12590,N_11761,N_10721);
or U12591 (N_12591,N_10928,N_11875);
or U12592 (N_12592,N_11132,N_10768);
nor U12593 (N_12593,N_11946,N_11819);
or U12594 (N_12594,N_10740,N_11133);
nand U12595 (N_12595,N_11338,N_10843);
nand U12596 (N_12596,N_11415,N_11598);
or U12597 (N_12597,N_11753,N_11686);
nor U12598 (N_12598,N_10675,N_11452);
nor U12599 (N_12599,N_11750,N_10841);
or U12600 (N_12600,N_11071,N_10730);
xor U12601 (N_12601,N_11468,N_10616);
xnor U12602 (N_12602,N_10999,N_11299);
nand U12603 (N_12603,N_10971,N_11687);
and U12604 (N_12604,N_11508,N_10793);
nor U12605 (N_12605,N_11606,N_11778);
or U12606 (N_12606,N_11739,N_11615);
or U12607 (N_12607,N_11146,N_11100);
and U12608 (N_12608,N_11757,N_11234);
nand U12609 (N_12609,N_11987,N_11502);
nor U12610 (N_12610,N_10615,N_11777);
nand U12611 (N_12611,N_10958,N_10806);
nand U12612 (N_12612,N_11094,N_10551);
xor U12613 (N_12613,N_10516,N_10518);
or U12614 (N_12614,N_11151,N_10773);
or U12615 (N_12615,N_11866,N_11288);
nor U12616 (N_12616,N_10979,N_11423);
and U12617 (N_12617,N_11109,N_11695);
nor U12618 (N_12618,N_11087,N_11046);
nand U12619 (N_12619,N_11420,N_11341);
xnor U12620 (N_12620,N_11911,N_11259);
nand U12621 (N_12621,N_10802,N_10997);
nand U12622 (N_12622,N_11527,N_11190);
nor U12623 (N_12623,N_10600,N_11293);
and U12624 (N_12624,N_11531,N_11267);
nor U12625 (N_12625,N_11388,N_11260);
nand U12626 (N_12626,N_11517,N_11176);
or U12627 (N_12627,N_11574,N_10813);
nor U12628 (N_12628,N_11984,N_10953);
nor U12629 (N_12629,N_11182,N_11365);
nor U12630 (N_12630,N_11164,N_10955);
or U12631 (N_12631,N_10692,N_11533);
or U12632 (N_12632,N_11940,N_11178);
and U12633 (N_12633,N_11865,N_11116);
and U12634 (N_12634,N_10821,N_11805);
and U12635 (N_12635,N_10638,N_11942);
or U12636 (N_12636,N_11832,N_10756);
and U12637 (N_12637,N_11592,N_10897);
or U12638 (N_12638,N_11359,N_11876);
nor U12639 (N_12639,N_11969,N_10837);
and U12640 (N_12640,N_11924,N_11916);
xor U12641 (N_12641,N_11552,N_10986);
or U12642 (N_12642,N_11189,N_11993);
and U12643 (N_12643,N_11249,N_11912);
xnor U12644 (N_12644,N_10700,N_11741);
or U12645 (N_12645,N_11980,N_11650);
nand U12646 (N_12646,N_10735,N_11149);
or U12647 (N_12647,N_11037,N_11770);
and U12648 (N_12648,N_10512,N_11989);
nand U12649 (N_12649,N_10820,N_11829);
or U12650 (N_12650,N_11329,N_11367);
or U12651 (N_12651,N_11841,N_11818);
nor U12652 (N_12652,N_11128,N_11089);
or U12653 (N_12653,N_11430,N_10694);
nand U12654 (N_12654,N_11621,N_10775);
and U12655 (N_12655,N_10878,N_11271);
nand U12656 (N_12656,N_11713,N_11784);
nor U12657 (N_12657,N_11350,N_11848);
nand U12658 (N_12658,N_11471,N_11600);
and U12659 (N_12659,N_11576,N_11296);
or U12660 (N_12660,N_10610,N_11715);
nand U12661 (N_12661,N_11010,N_11925);
nand U12662 (N_12662,N_11723,N_11586);
or U12663 (N_12663,N_11175,N_11390);
nor U12664 (N_12664,N_11545,N_11629);
or U12665 (N_12665,N_11622,N_11300);
and U12666 (N_12666,N_11309,N_11326);
xor U12667 (N_12667,N_11938,N_11018);
nor U12668 (N_12668,N_10931,N_11327);
or U12669 (N_12669,N_11528,N_11059);
nand U12670 (N_12670,N_11879,N_11250);
nand U12671 (N_12671,N_10671,N_11746);
nand U12672 (N_12672,N_11360,N_11160);
nor U12673 (N_12673,N_11340,N_11562);
or U12674 (N_12674,N_10992,N_11934);
or U12675 (N_12675,N_11731,N_10748);
and U12676 (N_12676,N_10719,N_10727);
nand U12677 (N_12677,N_11678,N_10967);
nand U12678 (N_12678,N_11381,N_10988);
nor U12679 (N_12679,N_10816,N_10921);
and U12680 (N_12680,N_11668,N_11263);
or U12681 (N_12681,N_10894,N_10517);
nand U12682 (N_12682,N_11438,N_10948);
nor U12683 (N_12683,N_11268,N_11355);
and U12684 (N_12684,N_11447,N_11639);
and U12685 (N_12685,N_11026,N_10936);
nor U12686 (N_12686,N_11194,N_11855);
nand U12687 (N_12687,N_11185,N_11174);
nand U12688 (N_12688,N_10751,N_11965);
or U12689 (N_12689,N_11199,N_11737);
nor U12690 (N_12690,N_11437,N_11861);
nor U12691 (N_12691,N_10918,N_11847);
and U12692 (N_12692,N_11278,N_11324);
nand U12693 (N_12693,N_11956,N_11835);
or U12694 (N_12694,N_11717,N_10840);
and U12695 (N_12695,N_11870,N_10579);
and U12696 (N_12696,N_11991,N_11239);
nor U12697 (N_12697,N_11624,N_11590);
nor U12698 (N_12698,N_10993,N_11364);
or U12699 (N_12699,N_10522,N_11954);
nor U12700 (N_12700,N_11392,N_10618);
and U12701 (N_12701,N_11894,N_10925);
or U12702 (N_12702,N_10823,N_11356);
and U12703 (N_12703,N_11482,N_10612);
nor U12704 (N_12704,N_10797,N_11095);
nor U12705 (N_12705,N_11636,N_11497);
xnor U12706 (N_12706,N_11921,N_11455);
nand U12707 (N_12707,N_11960,N_11195);
and U12708 (N_12708,N_11041,N_10642);
nand U12709 (N_12709,N_11738,N_11547);
xnor U12710 (N_12710,N_11888,N_10794);
or U12711 (N_12711,N_11677,N_11457);
and U12712 (N_12712,N_10738,N_10533);
and U12713 (N_12713,N_11426,N_10779);
and U12714 (N_12714,N_10676,N_11031);
or U12715 (N_12715,N_11140,N_11755);
or U12716 (N_12716,N_11609,N_11988);
nor U12717 (N_12717,N_11667,N_11330);
and U12718 (N_12718,N_10669,N_11391);
and U12719 (N_12719,N_11957,N_11627);
xor U12720 (N_12720,N_10777,N_11192);
and U12721 (N_12721,N_11351,N_10934);
and U12722 (N_12722,N_11034,N_11572);
nand U12723 (N_12723,N_11793,N_11665);
nand U12724 (N_12724,N_11863,N_11724);
and U12725 (N_12725,N_10811,N_11119);
or U12726 (N_12726,N_10846,N_11019);
and U12727 (N_12727,N_10592,N_10945);
nand U12728 (N_12728,N_10830,N_11449);
nor U12729 (N_12729,N_11067,N_11812);
or U12730 (N_12730,N_11209,N_11548);
nor U12731 (N_12731,N_11428,N_10660);
or U12732 (N_12732,N_11926,N_10674);
nor U12733 (N_12733,N_10585,N_10767);
xnor U12734 (N_12734,N_11577,N_11850);
nor U12735 (N_12735,N_11670,N_11498);
nand U12736 (N_12736,N_10781,N_11955);
or U12737 (N_12737,N_10626,N_10898);
nand U12738 (N_12738,N_10568,N_10741);
or U12739 (N_12739,N_11045,N_11298);
nand U12740 (N_12740,N_10772,N_11403);
nand U12741 (N_12741,N_11120,N_11718);
or U12742 (N_12742,N_11292,N_11721);
nor U12743 (N_12743,N_11429,N_11663);
and U12744 (N_12744,N_11795,N_11885);
nand U12745 (N_12745,N_10690,N_11198);
and U12746 (N_12746,N_11553,N_10849);
nor U12747 (N_12747,N_10851,N_11788);
and U12748 (N_12748,N_10834,N_10923);
and U12749 (N_12749,N_10555,N_11072);
or U12750 (N_12750,N_11683,N_10853);
or U12751 (N_12751,N_11896,N_11985);
xor U12752 (N_12752,N_11675,N_11256);
nand U12753 (N_12753,N_10864,N_10861);
or U12754 (N_12754,N_10840,N_11226);
or U12755 (N_12755,N_11137,N_10840);
and U12756 (N_12756,N_10929,N_10692);
and U12757 (N_12757,N_11303,N_11478);
nand U12758 (N_12758,N_11771,N_10612);
or U12759 (N_12759,N_11458,N_11205);
nor U12760 (N_12760,N_11351,N_11008);
nand U12761 (N_12761,N_10533,N_11324);
and U12762 (N_12762,N_10930,N_11637);
nand U12763 (N_12763,N_10752,N_11724);
nand U12764 (N_12764,N_11209,N_11214);
or U12765 (N_12765,N_11889,N_10736);
and U12766 (N_12766,N_10519,N_11348);
nor U12767 (N_12767,N_11495,N_11920);
nand U12768 (N_12768,N_11921,N_11518);
nand U12769 (N_12769,N_11937,N_11970);
and U12770 (N_12770,N_11994,N_11774);
and U12771 (N_12771,N_10971,N_10834);
nand U12772 (N_12772,N_10975,N_10690);
nor U12773 (N_12773,N_11035,N_11687);
nor U12774 (N_12774,N_11465,N_11015);
nand U12775 (N_12775,N_10708,N_11660);
xnor U12776 (N_12776,N_10870,N_11137);
or U12777 (N_12777,N_10896,N_11606);
or U12778 (N_12778,N_11509,N_11922);
nor U12779 (N_12779,N_11022,N_10568);
or U12780 (N_12780,N_10714,N_11419);
and U12781 (N_12781,N_11758,N_10653);
nand U12782 (N_12782,N_11481,N_11466);
xnor U12783 (N_12783,N_10773,N_10590);
and U12784 (N_12784,N_11475,N_11341);
and U12785 (N_12785,N_10588,N_11255);
xor U12786 (N_12786,N_11273,N_11470);
nand U12787 (N_12787,N_10801,N_11652);
nand U12788 (N_12788,N_11701,N_11106);
or U12789 (N_12789,N_11881,N_11006);
nand U12790 (N_12790,N_10737,N_10703);
nor U12791 (N_12791,N_11327,N_11926);
or U12792 (N_12792,N_11410,N_11025);
nand U12793 (N_12793,N_11610,N_11499);
xor U12794 (N_12794,N_10735,N_10666);
nand U12795 (N_12795,N_11682,N_11132);
or U12796 (N_12796,N_10501,N_11623);
xor U12797 (N_12797,N_10890,N_11812);
xnor U12798 (N_12798,N_10600,N_11145);
nand U12799 (N_12799,N_10643,N_10585);
nand U12800 (N_12800,N_11514,N_10950);
nor U12801 (N_12801,N_11885,N_11573);
and U12802 (N_12802,N_11970,N_10921);
or U12803 (N_12803,N_11258,N_10820);
nand U12804 (N_12804,N_11145,N_11874);
nand U12805 (N_12805,N_11547,N_11287);
nand U12806 (N_12806,N_11444,N_11187);
xnor U12807 (N_12807,N_11513,N_11997);
nand U12808 (N_12808,N_10624,N_11681);
nand U12809 (N_12809,N_10776,N_10579);
nand U12810 (N_12810,N_11329,N_10752);
nor U12811 (N_12811,N_11138,N_11924);
or U12812 (N_12812,N_11218,N_11975);
and U12813 (N_12813,N_11583,N_10753);
nand U12814 (N_12814,N_10729,N_11974);
xnor U12815 (N_12815,N_10917,N_11310);
or U12816 (N_12816,N_11909,N_10888);
nand U12817 (N_12817,N_10502,N_11269);
and U12818 (N_12818,N_10883,N_11084);
nand U12819 (N_12819,N_11086,N_11690);
and U12820 (N_12820,N_11720,N_11827);
or U12821 (N_12821,N_10643,N_11826);
nand U12822 (N_12822,N_10694,N_11567);
and U12823 (N_12823,N_11843,N_11045);
nor U12824 (N_12824,N_11727,N_11076);
nor U12825 (N_12825,N_11594,N_11645);
or U12826 (N_12826,N_11472,N_11745);
and U12827 (N_12827,N_11057,N_11938);
and U12828 (N_12828,N_11140,N_11541);
and U12829 (N_12829,N_11536,N_11477);
nor U12830 (N_12830,N_11932,N_10646);
and U12831 (N_12831,N_11226,N_11656);
nor U12832 (N_12832,N_10672,N_10580);
nand U12833 (N_12833,N_10753,N_11272);
or U12834 (N_12834,N_11407,N_11099);
or U12835 (N_12835,N_10985,N_11177);
nand U12836 (N_12836,N_10700,N_11161);
nor U12837 (N_12837,N_11103,N_11449);
nor U12838 (N_12838,N_11667,N_11416);
or U12839 (N_12839,N_10515,N_10739);
nor U12840 (N_12840,N_11179,N_11799);
and U12841 (N_12841,N_10800,N_10726);
nand U12842 (N_12842,N_11065,N_10523);
nand U12843 (N_12843,N_10954,N_10605);
nor U12844 (N_12844,N_10590,N_11543);
nand U12845 (N_12845,N_11224,N_10670);
nand U12846 (N_12846,N_10657,N_11183);
and U12847 (N_12847,N_11178,N_10628);
nand U12848 (N_12848,N_11959,N_10592);
or U12849 (N_12849,N_11931,N_11021);
and U12850 (N_12850,N_10732,N_11326);
nand U12851 (N_12851,N_10842,N_10953);
or U12852 (N_12852,N_11950,N_11875);
nor U12853 (N_12853,N_11435,N_11942);
nand U12854 (N_12854,N_10832,N_10871);
xor U12855 (N_12855,N_10895,N_11004);
nand U12856 (N_12856,N_10729,N_11356);
nand U12857 (N_12857,N_11880,N_10587);
nor U12858 (N_12858,N_10856,N_11717);
nor U12859 (N_12859,N_10993,N_10826);
nand U12860 (N_12860,N_10517,N_11761);
and U12861 (N_12861,N_11316,N_11908);
or U12862 (N_12862,N_10797,N_10916);
nand U12863 (N_12863,N_11308,N_11827);
nand U12864 (N_12864,N_10615,N_11110);
and U12865 (N_12865,N_11119,N_11670);
xnor U12866 (N_12866,N_11053,N_11502);
and U12867 (N_12867,N_11718,N_10848);
and U12868 (N_12868,N_10719,N_10924);
nand U12869 (N_12869,N_11456,N_10950);
and U12870 (N_12870,N_11799,N_10913);
nand U12871 (N_12871,N_10714,N_11314);
nor U12872 (N_12872,N_11482,N_11852);
nand U12873 (N_12873,N_11270,N_10743);
nand U12874 (N_12874,N_10969,N_11674);
nor U12875 (N_12875,N_10850,N_11199);
or U12876 (N_12876,N_10919,N_10602);
nor U12877 (N_12877,N_10953,N_11436);
nor U12878 (N_12878,N_11207,N_11719);
nand U12879 (N_12879,N_11837,N_11173);
nand U12880 (N_12880,N_10838,N_11751);
xor U12881 (N_12881,N_11799,N_10744);
or U12882 (N_12882,N_11048,N_11087);
xor U12883 (N_12883,N_11037,N_11524);
or U12884 (N_12884,N_10941,N_11928);
nand U12885 (N_12885,N_11588,N_10632);
nor U12886 (N_12886,N_11259,N_11202);
and U12887 (N_12887,N_11887,N_10939);
and U12888 (N_12888,N_11139,N_10731);
or U12889 (N_12889,N_11062,N_11430);
xnor U12890 (N_12890,N_10508,N_11915);
nor U12891 (N_12891,N_11283,N_10987);
and U12892 (N_12892,N_11254,N_11156);
and U12893 (N_12893,N_10519,N_11989);
nor U12894 (N_12894,N_10525,N_11510);
or U12895 (N_12895,N_10591,N_10744);
nand U12896 (N_12896,N_11402,N_11979);
and U12897 (N_12897,N_10941,N_11875);
nand U12898 (N_12898,N_10707,N_11035);
nor U12899 (N_12899,N_11703,N_10810);
and U12900 (N_12900,N_11815,N_10718);
nor U12901 (N_12901,N_10906,N_11705);
nor U12902 (N_12902,N_10663,N_10898);
nor U12903 (N_12903,N_10571,N_11651);
or U12904 (N_12904,N_11948,N_11919);
nor U12905 (N_12905,N_10769,N_11005);
nand U12906 (N_12906,N_11402,N_10828);
nor U12907 (N_12907,N_11877,N_11745);
nand U12908 (N_12908,N_11929,N_11583);
nand U12909 (N_12909,N_11974,N_11924);
or U12910 (N_12910,N_10770,N_11933);
nand U12911 (N_12911,N_11779,N_11503);
and U12912 (N_12912,N_10932,N_10828);
or U12913 (N_12913,N_11902,N_11624);
xnor U12914 (N_12914,N_11881,N_11149);
nor U12915 (N_12915,N_11757,N_11918);
nand U12916 (N_12916,N_11385,N_10800);
nor U12917 (N_12917,N_11998,N_10519);
or U12918 (N_12918,N_11202,N_10680);
and U12919 (N_12919,N_11349,N_10887);
nor U12920 (N_12920,N_11346,N_10703);
and U12921 (N_12921,N_11958,N_11756);
xor U12922 (N_12922,N_11095,N_11806);
xnor U12923 (N_12923,N_11089,N_11001);
or U12924 (N_12924,N_10617,N_10599);
nand U12925 (N_12925,N_11339,N_10841);
nor U12926 (N_12926,N_10786,N_10873);
nor U12927 (N_12927,N_11285,N_10635);
nand U12928 (N_12928,N_11980,N_11798);
nor U12929 (N_12929,N_10507,N_11714);
and U12930 (N_12930,N_10690,N_10978);
nand U12931 (N_12931,N_10834,N_11026);
xor U12932 (N_12932,N_11714,N_11217);
nand U12933 (N_12933,N_11717,N_10708);
and U12934 (N_12934,N_10763,N_11492);
nor U12935 (N_12935,N_10857,N_10966);
nor U12936 (N_12936,N_11264,N_10677);
and U12937 (N_12937,N_11614,N_11305);
nor U12938 (N_12938,N_11261,N_10753);
nor U12939 (N_12939,N_10779,N_11869);
nor U12940 (N_12940,N_11834,N_10830);
or U12941 (N_12941,N_11876,N_11701);
xnor U12942 (N_12942,N_11719,N_10812);
nor U12943 (N_12943,N_11828,N_11739);
and U12944 (N_12944,N_11864,N_11849);
and U12945 (N_12945,N_11256,N_10878);
nor U12946 (N_12946,N_11181,N_11284);
and U12947 (N_12947,N_11298,N_11771);
or U12948 (N_12948,N_10833,N_11126);
nor U12949 (N_12949,N_11851,N_11167);
nand U12950 (N_12950,N_11072,N_11005);
nand U12951 (N_12951,N_11971,N_11681);
nor U12952 (N_12952,N_11394,N_11012);
and U12953 (N_12953,N_11187,N_11572);
xor U12954 (N_12954,N_11718,N_11212);
or U12955 (N_12955,N_11617,N_11604);
nor U12956 (N_12956,N_10563,N_11614);
xnor U12957 (N_12957,N_11507,N_11680);
nand U12958 (N_12958,N_11710,N_11588);
nor U12959 (N_12959,N_11076,N_11875);
and U12960 (N_12960,N_10707,N_11154);
nor U12961 (N_12961,N_11013,N_10631);
nand U12962 (N_12962,N_11311,N_11668);
nor U12963 (N_12963,N_10709,N_11584);
and U12964 (N_12964,N_11668,N_10769);
xor U12965 (N_12965,N_11740,N_10634);
nand U12966 (N_12966,N_11450,N_11757);
xor U12967 (N_12967,N_11683,N_10680);
or U12968 (N_12968,N_11737,N_11154);
nor U12969 (N_12969,N_10656,N_10638);
and U12970 (N_12970,N_10781,N_10623);
nor U12971 (N_12971,N_10960,N_11738);
and U12972 (N_12972,N_11110,N_11685);
xnor U12973 (N_12973,N_11037,N_11528);
nor U12974 (N_12974,N_11834,N_10799);
nand U12975 (N_12975,N_10801,N_11605);
nand U12976 (N_12976,N_11348,N_11752);
xor U12977 (N_12977,N_11734,N_11958);
nor U12978 (N_12978,N_11221,N_10926);
xnor U12979 (N_12979,N_10862,N_10848);
nor U12980 (N_12980,N_11015,N_11027);
or U12981 (N_12981,N_11267,N_10529);
nor U12982 (N_12982,N_11271,N_11877);
nor U12983 (N_12983,N_11556,N_11461);
nand U12984 (N_12984,N_10999,N_10625);
nand U12985 (N_12985,N_11705,N_10825);
nor U12986 (N_12986,N_10876,N_11926);
nor U12987 (N_12987,N_10822,N_11899);
or U12988 (N_12988,N_10673,N_11403);
or U12989 (N_12989,N_10728,N_11392);
nand U12990 (N_12990,N_10569,N_11389);
and U12991 (N_12991,N_11454,N_11446);
nor U12992 (N_12992,N_10678,N_11911);
and U12993 (N_12993,N_10667,N_11597);
nor U12994 (N_12994,N_10769,N_10823);
or U12995 (N_12995,N_11633,N_11785);
and U12996 (N_12996,N_10824,N_10813);
and U12997 (N_12997,N_11134,N_11896);
or U12998 (N_12998,N_11692,N_10805);
or U12999 (N_12999,N_10520,N_11559);
nor U13000 (N_13000,N_11706,N_11562);
nor U13001 (N_13001,N_11364,N_11924);
and U13002 (N_13002,N_11477,N_10926);
nand U13003 (N_13003,N_11171,N_11369);
nor U13004 (N_13004,N_11593,N_10979);
nor U13005 (N_13005,N_10969,N_11211);
nand U13006 (N_13006,N_11809,N_10562);
and U13007 (N_13007,N_11865,N_11814);
and U13008 (N_13008,N_11102,N_10685);
and U13009 (N_13009,N_10975,N_11237);
nand U13010 (N_13010,N_11811,N_11903);
nand U13011 (N_13011,N_11851,N_11586);
xor U13012 (N_13012,N_11723,N_10561);
or U13013 (N_13013,N_11181,N_11085);
nand U13014 (N_13014,N_10561,N_11372);
nand U13015 (N_13015,N_11460,N_11446);
nand U13016 (N_13016,N_11903,N_11858);
or U13017 (N_13017,N_10991,N_10771);
or U13018 (N_13018,N_11546,N_11559);
nor U13019 (N_13019,N_11526,N_10526);
and U13020 (N_13020,N_11112,N_10882);
nand U13021 (N_13021,N_11078,N_11330);
xnor U13022 (N_13022,N_11389,N_11369);
nor U13023 (N_13023,N_11342,N_10643);
nor U13024 (N_13024,N_11040,N_10949);
nand U13025 (N_13025,N_11567,N_10711);
and U13026 (N_13026,N_10819,N_11008);
nand U13027 (N_13027,N_11487,N_10892);
nor U13028 (N_13028,N_11415,N_10544);
xnor U13029 (N_13029,N_10909,N_10532);
nand U13030 (N_13030,N_11692,N_11679);
xnor U13031 (N_13031,N_11884,N_10953);
or U13032 (N_13032,N_11291,N_11641);
nor U13033 (N_13033,N_10814,N_11286);
and U13034 (N_13034,N_11813,N_11623);
nand U13035 (N_13035,N_11507,N_11399);
or U13036 (N_13036,N_10880,N_11901);
or U13037 (N_13037,N_11813,N_11398);
and U13038 (N_13038,N_11803,N_11785);
and U13039 (N_13039,N_10747,N_11298);
xor U13040 (N_13040,N_10520,N_11371);
and U13041 (N_13041,N_10568,N_11249);
nor U13042 (N_13042,N_10596,N_10599);
nand U13043 (N_13043,N_11752,N_11372);
or U13044 (N_13044,N_11560,N_11989);
and U13045 (N_13045,N_11290,N_11190);
nor U13046 (N_13046,N_11611,N_11207);
or U13047 (N_13047,N_10854,N_11410);
nor U13048 (N_13048,N_10524,N_11212);
nand U13049 (N_13049,N_11567,N_11340);
nor U13050 (N_13050,N_11531,N_10632);
nand U13051 (N_13051,N_11357,N_11630);
xor U13052 (N_13052,N_11581,N_11852);
and U13053 (N_13053,N_11581,N_10910);
xnor U13054 (N_13054,N_11990,N_10677);
nand U13055 (N_13055,N_10543,N_10813);
nor U13056 (N_13056,N_10827,N_11345);
nor U13057 (N_13057,N_10904,N_11219);
and U13058 (N_13058,N_11739,N_11913);
or U13059 (N_13059,N_11194,N_11851);
or U13060 (N_13060,N_10614,N_11053);
or U13061 (N_13061,N_11835,N_11780);
nor U13062 (N_13062,N_11152,N_11338);
or U13063 (N_13063,N_10997,N_10590);
xor U13064 (N_13064,N_11623,N_10802);
nand U13065 (N_13065,N_10955,N_11725);
nor U13066 (N_13066,N_10965,N_10972);
nand U13067 (N_13067,N_10570,N_10898);
nand U13068 (N_13068,N_11518,N_10597);
and U13069 (N_13069,N_11721,N_10628);
and U13070 (N_13070,N_11004,N_10931);
and U13071 (N_13071,N_10537,N_11127);
and U13072 (N_13072,N_11758,N_10810);
nand U13073 (N_13073,N_11236,N_10766);
nand U13074 (N_13074,N_11951,N_10613);
and U13075 (N_13075,N_11842,N_10747);
and U13076 (N_13076,N_10565,N_10714);
nor U13077 (N_13077,N_10648,N_10920);
and U13078 (N_13078,N_10896,N_11348);
nand U13079 (N_13079,N_11729,N_10766);
nor U13080 (N_13080,N_11592,N_10872);
nor U13081 (N_13081,N_11950,N_11945);
or U13082 (N_13082,N_11627,N_11348);
nor U13083 (N_13083,N_11069,N_10636);
nand U13084 (N_13084,N_11609,N_10740);
and U13085 (N_13085,N_11866,N_11683);
nand U13086 (N_13086,N_11562,N_11955);
nor U13087 (N_13087,N_10572,N_11657);
or U13088 (N_13088,N_11751,N_10681);
or U13089 (N_13089,N_11619,N_10593);
nand U13090 (N_13090,N_11914,N_10723);
and U13091 (N_13091,N_10842,N_11311);
nor U13092 (N_13092,N_10983,N_11937);
xnor U13093 (N_13093,N_11729,N_10756);
and U13094 (N_13094,N_11923,N_10911);
or U13095 (N_13095,N_11576,N_10909);
or U13096 (N_13096,N_10797,N_10831);
nand U13097 (N_13097,N_11406,N_10583);
xnor U13098 (N_13098,N_11638,N_10693);
xnor U13099 (N_13099,N_10811,N_11215);
nand U13100 (N_13100,N_11110,N_10663);
nor U13101 (N_13101,N_10804,N_10826);
and U13102 (N_13102,N_11034,N_11011);
or U13103 (N_13103,N_11128,N_10603);
nor U13104 (N_13104,N_11415,N_11541);
or U13105 (N_13105,N_11953,N_11119);
and U13106 (N_13106,N_10546,N_11780);
nor U13107 (N_13107,N_11302,N_11655);
nand U13108 (N_13108,N_10547,N_11094);
or U13109 (N_13109,N_10909,N_11639);
or U13110 (N_13110,N_11229,N_10858);
and U13111 (N_13111,N_11441,N_11035);
and U13112 (N_13112,N_11872,N_10961);
or U13113 (N_13113,N_10912,N_11565);
nand U13114 (N_13114,N_11064,N_11770);
and U13115 (N_13115,N_11343,N_11548);
and U13116 (N_13116,N_11880,N_11062);
or U13117 (N_13117,N_11032,N_10524);
and U13118 (N_13118,N_10511,N_11908);
or U13119 (N_13119,N_11133,N_10856);
nor U13120 (N_13120,N_10798,N_11169);
or U13121 (N_13121,N_11742,N_11822);
and U13122 (N_13122,N_10707,N_10895);
nor U13123 (N_13123,N_11768,N_10608);
and U13124 (N_13124,N_11277,N_11735);
and U13125 (N_13125,N_11441,N_11763);
and U13126 (N_13126,N_11889,N_10857);
or U13127 (N_13127,N_10735,N_11826);
nor U13128 (N_13128,N_11025,N_11246);
and U13129 (N_13129,N_11537,N_10655);
nor U13130 (N_13130,N_11360,N_10991);
nor U13131 (N_13131,N_11422,N_10807);
nor U13132 (N_13132,N_10507,N_11532);
nand U13133 (N_13133,N_11019,N_10905);
nor U13134 (N_13134,N_10817,N_11564);
and U13135 (N_13135,N_10724,N_11746);
or U13136 (N_13136,N_11936,N_11430);
nand U13137 (N_13137,N_11080,N_11750);
nor U13138 (N_13138,N_11189,N_10658);
nand U13139 (N_13139,N_11735,N_11896);
xnor U13140 (N_13140,N_11134,N_11675);
or U13141 (N_13141,N_10699,N_11181);
nand U13142 (N_13142,N_11628,N_10851);
and U13143 (N_13143,N_10595,N_10658);
or U13144 (N_13144,N_10823,N_11864);
and U13145 (N_13145,N_11483,N_11182);
nand U13146 (N_13146,N_10737,N_11092);
or U13147 (N_13147,N_11734,N_11679);
xnor U13148 (N_13148,N_10573,N_11210);
and U13149 (N_13149,N_10795,N_11010);
and U13150 (N_13150,N_11523,N_11032);
nor U13151 (N_13151,N_11362,N_11848);
xor U13152 (N_13152,N_11041,N_10674);
and U13153 (N_13153,N_11067,N_11510);
and U13154 (N_13154,N_11481,N_11456);
nand U13155 (N_13155,N_11123,N_11557);
and U13156 (N_13156,N_11996,N_11581);
and U13157 (N_13157,N_11131,N_11212);
and U13158 (N_13158,N_11310,N_10608);
and U13159 (N_13159,N_11363,N_10579);
nor U13160 (N_13160,N_11932,N_10926);
nand U13161 (N_13161,N_10976,N_11343);
nand U13162 (N_13162,N_10935,N_11314);
nand U13163 (N_13163,N_10896,N_11073);
xnor U13164 (N_13164,N_11774,N_11172);
or U13165 (N_13165,N_11484,N_11474);
and U13166 (N_13166,N_11129,N_10691);
and U13167 (N_13167,N_11100,N_11150);
or U13168 (N_13168,N_10745,N_10687);
nand U13169 (N_13169,N_11834,N_10570);
or U13170 (N_13170,N_11637,N_10946);
nand U13171 (N_13171,N_11660,N_10698);
or U13172 (N_13172,N_11084,N_11164);
nand U13173 (N_13173,N_11523,N_11633);
nor U13174 (N_13174,N_11727,N_10573);
nor U13175 (N_13175,N_11366,N_11003);
or U13176 (N_13176,N_11847,N_11632);
or U13177 (N_13177,N_10895,N_11078);
nand U13178 (N_13178,N_11588,N_11595);
or U13179 (N_13179,N_11741,N_11342);
or U13180 (N_13180,N_11196,N_10522);
nor U13181 (N_13181,N_11874,N_10842);
nand U13182 (N_13182,N_11609,N_11334);
xnor U13183 (N_13183,N_10982,N_11386);
nand U13184 (N_13184,N_11558,N_11072);
and U13185 (N_13185,N_11108,N_10935);
nand U13186 (N_13186,N_11875,N_11116);
and U13187 (N_13187,N_11659,N_10938);
nand U13188 (N_13188,N_10825,N_11388);
nor U13189 (N_13189,N_11510,N_11313);
nand U13190 (N_13190,N_11037,N_11748);
and U13191 (N_13191,N_10535,N_10521);
nand U13192 (N_13192,N_11984,N_10708);
and U13193 (N_13193,N_10619,N_11725);
xnor U13194 (N_13194,N_10787,N_11440);
or U13195 (N_13195,N_10943,N_11597);
xor U13196 (N_13196,N_10596,N_10527);
nor U13197 (N_13197,N_10807,N_10535);
nor U13198 (N_13198,N_11525,N_11157);
nor U13199 (N_13199,N_11727,N_10748);
or U13200 (N_13200,N_11967,N_11688);
nand U13201 (N_13201,N_10716,N_10801);
xnor U13202 (N_13202,N_10651,N_11386);
or U13203 (N_13203,N_11499,N_10896);
or U13204 (N_13204,N_11086,N_11541);
or U13205 (N_13205,N_11098,N_10744);
or U13206 (N_13206,N_10582,N_11583);
nand U13207 (N_13207,N_11343,N_10652);
nor U13208 (N_13208,N_11100,N_10589);
and U13209 (N_13209,N_10936,N_11932);
or U13210 (N_13210,N_11002,N_11283);
or U13211 (N_13211,N_11671,N_10793);
nor U13212 (N_13212,N_11738,N_11060);
nand U13213 (N_13213,N_11697,N_11461);
nand U13214 (N_13214,N_11734,N_11294);
nor U13215 (N_13215,N_11108,N_10613);
xnor U13216 (N_13216,N_11948,N_10605);
and U13217 (N_13217,N_10698,N_11291);
and U13218 (N_13218,N_10603,N_11803);
nor U13219 (N_13219,N_10566,N_10917);
and U13220 (N_13220,N_11091,N_10884);
nand U13221 (N_13221,N_10890,N_10645);
nor U13222 (N_13222,N_10950,N_11203);
or U13223 (N_13223,N_10705,N_10914);
nand U13224 (N_13224,N_11408,N_11948);
xor U13225 (N_13225,N_11164,N_10913);
nor U13226 (N_13226,N_11018,N_11027);
nor U13227 (N_13227,N_10806,N_10914);
xnor U13228 (N_13228,N_10709,N_10894);
or U13229 (N_13229,N_10865,N_10862);
nor U13230 (N_13230,N_11440,N_11452);
or U13231 (N_13231,N_11883,N_11156);
nand U13232 (N_13232,N_11109,N_10886);
nand U13233 (N_13233,N_11213,N_11561);
and U13234 (N_13234,N_11849,N_10923);
or U13235 (N_13235,N_11897,N_11277);
nand U13236 (N_13236,N_11084,N_10873);
nor U13237 (N_13237,N_11895,N_11572);
nand U13238 (N_13238,N_11781,N_11124);
and U13239 (N_13239,N_11462,N_11345);
or U13240 (N_13240,N_11859,N_10618);
and U13241 (N_13241,N_11584,N_11480);
and U13242 (N_13242,N_10789,N_11145);
nand U13243 (N_13243,N_10977,N_11967);
or U13244 (N_13244,N_11330,N_10914);
or U13245 (N_13245,N_11005,N_11687);
or U13246 (N_13246,N_11570,N_11138);
nand U13247 (N_13247,N_11687,N_10712);
nand U13248 (N_13248,N_11793,N_11271);
nor U13249 (N_13249,N_11724,N_10821);
or U13250 (N_13250,N_11561,N_10684);
and U13251 (N_13251,N_11729,N_11470);
and U13252 (N_13252,N_11342,N_11326);
and U13253 (N_13253,N_11168,N_11887);
and U13254 (N_13254,N_11287,N_11000);
nor U13255 (N_13255,N_10679,N_11385);
and U13256 (N_13256,N_10599,N_11174);
nor U13257 (N_13257,N_10909,N_10694);
nor U13258 (N_13258,N_11656,N_10923);
or U13259 (N_13259,N_11371,N_11948);
and U13260 (N_13260,N_11910,N_11839);
nand U13261 (N_13261,N_11347,N_11861);
and U13262 (N_13262,N_11578,N_10884);
or U13263 (N_13263,N_11359,N_10653);
or U13264 (N_13264,N_10882,N_11613);
or U13265 (N_13265,N_10563,N_11243);
xor U13266 (N_13266,N_11585,N_10917);
nand U13267 (N_13267,N_10564,N_11285);
nand U13268 (N_13268,N_11830,N_11890);
and U13269 (N_13269,N_10840,N_11166);
xnor U13270 (N_13270,N_11562,N_10598);
and U13271 (N_13271,N_11692,N_11213);
and U13272 (N_13272,N_11373,N_10977);
xnor U13273 (N_13273,N_11301,N_11075);
nor U13274 (N_13274,N_10949,N_11197);
nand U13275 (N_13275,N_10965,N_10582);
or U13276 (N_13276,N_10598,N_11383);
and U13277 (N_13277,N_10915,N_10972);
and U13278 (N_13278,N_10652,N_10892);
or U13279 (N_13279,N_11548,N_11200);
nand U13280 (N_13280,N_11714,N_11314);
nor U13281 (N_13281,N_10590,N_10952);
or U13282 (N_13282,N_11081,N_10772);
xor U13283 (N_13283,N_11771,N_11945);
nor U13284 (N_13284,N_11087,N_11215);
and U13285 (N_13285,N_10787,N_11978);
or U13286 (N_13286,N_11588,N_10994);
nand U13287 (N_13287,N_10508,N_11289);
and U13288 (N_13288,N_11160,N_11321);
or U13289 (N_13289,N_10784,N_11368);
or U13290 (N_13290,N_11996,N_11815);
nor U13291 (N_13291,N_10722,N_11287);
nor U13292 (N_13292,N_10556,N_11998);
nand U13293 (N_13293,N_11042,N_11783);
nand U13294 (N_13294,N_10994,N_11601);
nor U13295 (N_13295,N_11908,N_10802);
or U13296 (N_13296,N_10925,N_11876);
and U13297 (N_13297,N_10902,N_11595);
nor U13298 (N_13298,N_11367,N_11044);
and U13299 (N_13299,N_11903,N_11899);
nor U13300 (N_13300,N_11594,N_10948);
or U13301 (N_13301,N_11146,N_11132);
and U13302 (N_13302,N_10961,N_11105);
or U13303 (N_13303,N_10617,N_11306);
xnor U13304 (N_13304,N_11936,N_10927);
or U13305 (N_13305,N_11524,N_10608);
and U13306 (N_13306,N_11351,N_10735);
nor U13307 (N_13307,N_11025,N_10530);
and U13308 (N_13308,N_11935,N_10607);
nand U13309 (N_13309,N_10687,N_11440);
or U13310 (N_13310,N_11639,N_11410);
nand U13311 (N_13311,N_11914,N_10534);
or U13312 (N_13312,N_10652,N_11326);
nand U13313 (N_13313,N_11014,N_11077);
nand U13314 (N_13314,N_10636,N_11563);
and U13315 (N_13315,N_11764,N_11884);
and U13316 (N_13316,N_11391,N_11012);
xor U13317 (N_13317,N_10777,N_11938);
nor U13318 (N_13318,N_11622,N_10752);
or U13319 (N_13319,N_10568,N_11628);
nand U13320 (N_13320,N_10794,N_11617);
nor U13321 (N_13321,N_10587,N_11545);
xnor U13322 (N_13322,N_11570,N_11752);
nor U13323 (N_13323,N_11773,N_11404);
nand U13324 (N_13324,N_11103,N_11161);
and U13325 (N_13325,N_10962,N_11205);
nor U13326 (N_13326,N_11373,N_10963);
and U13327 (N_13327,N_11534,N_10894);
or U13328 (N_13328,N_11575,N_11442);
nor U13329 (N_13329,N_10661,N_11406);
xnor U13330 (N_13330,N_11270,N_11217);
nor U13331 (N_13331,N_11369,N_11921);
and U13332 (N_13332,N_10602,N_10722);
nand U13333 (N_13333,N_11336,N_11057);
xor U13334 (N_13334,N_11304,N_11307);
nand U13335 (N_13335,N_11538,N_11143);
nor U13336 (N_13336,N_11448,N_11441);
nand U13337 (N_13337,N_10729,N_11339);
and U13338 (N_13338,N_11007,N_11696);
nand U13339 (N_13339,N_11666,N_11691);
nor U13340 (N_13340,N_11165,N_11972);
nor U13341 (N_13341,N_11735,N_11367);
nand U13342 (N_13342,N_11567,N_11529);
or U13343 (N_13343,N_11624,N_11340);
and U13344 (N_13344,N_10747,N_10959);
and U13345 (N_13345,N_11304,N_11327);
xnor U13346 (N_13346,N_11136,N_11617);
nor U13347 (N_13347,N_10630,N_11993);
xnor U13348 (N_13348,N_11992,N_11850);
nand U13349 (N_13349,N_11000,N_11819);
nand U13350 (N_13350,N_10670,N_11615);
nand U13351 (N_13351,N_10888,N_11651);
and U13352 (N_13352,N_11513,N_11316);
and U13353 (N_13353,N_10534,N_11074);
xor U13354 (N_13354,N_11359,N_11037);
nor U13355 (N_13355,N_11573,N_10699);
or U13356 (N_13356,N_11118,N_11834);
or U13357 (N_13357,N_11944,N_11337);
nor U13358 (N_13358,N_10646,N_11336);
or U13359 (N_13359,N_11133,N_11469);
nor U13360 (N_13360,N_11660,N_10645);
or U13361 (N_13361,N_10958,N_11625);
and U13362 (N_13362,N_10963,N_11422);
or U13363 (N_13363,N_11629,N_10812);
xor U13364 (N_13364,N_11830,N_11068);
nor U13365 (N_13365,N_11174,N_11613);
nand U13366 (N_13366,N_10684,N_10816);
or U13367 (N_13367,N_11688,N_11568);
nor U13368 (N_13368,N_11653,N_11454);
and U13369 (N_13369,N_10514,N_11961);
nand U13370 (N_13370,N_10836,N_10654);
or U13371 (N_13371,N_10730,N_11414);
and U13372 (N_13372,N_10741,N_11385);
xor U13373 (N_13373,N_10837,N_10934);
nor U13374 (N_13374,N_10744,N_10921);
or U13375 (N_13375,N_11647,N_11740);
nand U13376 (N_13376,N_11601,N_11524);
nand U13377 (N_13377,N_11184,N_11994);
nand U13378 (N_13378,N_11303,N_11621);
and U13379 (N_13379,N_10638,N_11431);
xnor U13380 (N_13380,N_11151,N_11938);
or U13381 (N_13381,N_11379,N_10848);
or U13382 (N_13382,N_11792,N_11195);
xnor U13383 (N_13383,N_11183,N_11442);
nor U13384 (N_13384,N_11341,N_10662);
xor U13385 (N_13385,N_11550,N_11093);
nor U13386 (N_13386,N_11379,N_11440);
and U13387 (N_13387,N_10999,N_11337);
nor U13388 (N_13388,N_11197,N_11251);
and U13389 (N_13389,N_10529,N_10856);
xor U13390 (N_13390,N_10801,N_11379);
nor U13391 (N_13391,N_11216,N_11398);
and U13392 (N_13392,N_11121,N_11133);
nand U13393 (N_13393,N_11366,N_11395);
nand U13394 (N_13394,N_11718,N_11277);
nor U13395 (N_13395,N_11774,N_11256);
or U13396 (N_13396,N_11547,N_11560);
or U13397 (N_13397,N_11282,N_11501);
nor U13398 (N_13398,N_10955,N_10873);
xnor U13399 (N_13399,N_11026,N_10654);
nand U13400 (N_13400,N_11113,N_11332);
xnor U13401 (N_13401,N_11382,N_11883);
and U13402 (N_13402,N_10832,N_11523);
or U13403 (N_13403,N_11441,N_10812);
nand U13404 (N_13404,N_11364,N_11164);
or U13405 (N_13405,N_10868,N_11205);
or U13406 (N_13406,N_11392,N_10713);
nand U13407 (N_13407,N_11020,N_11066);
or U13408 (N_13408,N_11208,N_11957);
nor U13409 (N_13409,N_11732,N_11538);
nor U13410 (N_13410,N_10845,N_11268);
nand U13411 (N_13411,N_11509,N_11982);
nand U13412 (N_13412,N_11971,N_11975);
or U13413 (N_13413,N_11769,N_11764);
nor U13414 (N_13414,N_11573,N_11773);
nor U13415 (N_13415,N_10512,N_11326);
xor U13416 (N_13416,N_10751,N_11829);
or U13417 (N_13417,N_10572,N_10637);
nand U13418 (N_13418,N_11775,N_10763);
nor U13419 (N_13419,N_11773,N_11621);
nand U13420 (N_13420,N_10541,N_11870);
or U13421 (N_13421,N_11438,N_11304);
nor U13422 (N_13422,N_10866,N_10741);
nor U13423 (N_13423,N_11699,N_11514);
nor U13424 (N_13424,N_10824,N_11089);
nor U13425 (N_13425,N_11881,N_11260);
nand U13426 (N_13426,N_11654,N_10840);
nand U13427 (N_13427,N_11601,N_11041);
and U13428 (N_13428,N_11001,N_10903);
and U13429 (N_13429,N_10735,N_10868);
or U13430 (N_13430,N_10521,N_11476);
and U13431 (N_13431,N_11257,N_11982);
nand U13432 (N_13432,N_11174,N_10877);
and U13433 (N_13433,N_10812,N_11986);
and U13434 (N_13434,N_10669,N_10903);
nor U13435 (N_13435,N_10606,N_11861);
and U13436 (N_13436,N_11207,N_11258);
nor U13437 (N_13437,N_10541,N_11691);
nor U13438 (N_13438,N_10926,N_10754);
nand U13439 (N_13439,N_10777,N_11173);
or U13440 (N_13440,N_11110,N_11734);
xnor U13441 (N_13441,N_11166,N_11778);
or U13442 (N_13442,N_10921,N_10552);
or U13443 (N_13443,N_11841,N_11510);
nor U13444 (N_13444,N_11986,N_11099);
or U13445 (N_13445,N_10806,N_11361);
and U13446 (N_13446,N_10918,N_10994);
or U13447 (N_13447,N_10509,N_10980);
nor U13448 (N_13448,N_10945,N_11821);
nand U13449 (N_13449,N_11739,N_11170);
and U13450 (N_13450,N_10734,N_11284);
or U13451 (N_13451,N_11823,N_11475);
xnor U13452 (N_13452,N_10905,N_11293);
nor U13453 (N_13453,N_11138,N_10978);
nor U13454 (N_13454,N_11600,N_11182);
and U13455 (N_13455,N_11138,N_11744);
nand U13456 (N_13456,N_11586,N_10505);
nand U13457 (N_13457,N_10797,N_10622);
nand U13458 (N_13458,N_11034,N_11272);
xnor U13459 (N_13459,N_11080,N_11680);
xor U13460 (N_13460,N_11783,N_10949);
and U13461 (N_13461,N_11563,N_11247);
or U13462 (N_13462,N_11276,N_10918);
xor U13463 (N_13463,N_11955,N_11791);
and U13464 (N_13464,N_11052,N_11483);
nor U13465 (N_13465,N_10665,N_11886);
xnor U13466 (N_13466,N_10685,N_11435);
or U13467 (N_13467,N_11452,N_11866);
or U13468 (N_13468,N_10671,N_10958);
nor U13469 (N_13469,N_11360,N_11238);
and U13470 (N_13470,N_10509,N_11629);
or U13471 (N_13471,N_11554,N_11877);
nor U13472 (N_13472,N_11146,N_11452);
nand U13473 (N_13473,N_11203,N_11284);
nand U13474 (N_13474,N_11185,N_11116);
and U13475 (N_13475,N_11689,N_11693);
nand U13476 (N_13476,N_11612,N_11357);
nand U13477 (N_13477,N_11375,N_10724);
nand U13478 (N_13478,N_10621,N_10770);
and U13479 (N_13479,N_11252,N_11882);
nor U13480 (N_13480,N_11970,N_10577);
nand U13481 (N_13481,N_10536,N_10591);
and U13482 (N_13482,N_11530,N_10906);
nor U13483 (N_13483,N_10550,N_11628);
nand U13484 (N_13484,N_11620,N_11694);
and U13485 (N_13485,N_11454,N_10967);
nand U13486 (N_13486,N_11819,N_11438);
and U13487 (N_13487,N_11410,N_11655);
and U13488 (N_13488,N_11326,N_11770);
and U13489 (N_13489,N_10921,N_11917);
nand U13490 (N_13490,N_11247,N_11818);
xor U13491 (N_13491,N_10930,N_10939);
and U13492 (N_13492,N_11652,N_11668);
or U13493 (N_13493,N_10578,N_11353);
nor U13494 (N_13494,N_10878,N_11329);
nor U13495 (N_13495,N_10657,N_10553);
nor U13496 (N_13496,N_11356,N_11853);
xor U13497 (N_13497,N_11906,N_10946);
and U13498 (N_13498,N_11270,N_10654);
nand U13499 (N_13499,N_11573,N_11832);
and U13500 (N_13500,N_12164,N_12146);
nand U13501 (N_13501,N_12068,N_12256);
nor U13502 (N_13502,N_12231,N_13439);
nand U13503 (N_13503,N_12438,N_12924);
nor U13504 (N_13504,N_13048,N_12052);
nor U13505 (N_13505,N_12279,N_12436);
and U13506 (N_13506,N_12107,N_13478);
xnor U13507 (N_13507,N_13124,N_13071);
nand U13508 (N_13508,N_13097,N_12347);
and U13509 (N_13509,N_13093,N_12978);
nor U13510 (N_13510,N_13473,N_12062);
and U13511 (N_13511,N_12834,N_12562);
nand U13512 (N_13512,N_12717,N_12819);
xor U13513 (N_13513,N_13450,N_12796);
and U13514 (N_13514,N_12223,N_12678);
nor U13515 (N_13515,N_13249,N_12595);
or U13516 (N_13516,N_12518,N_12544);
nor U13517 (N_13517,N_13045,N_12890);
nand U13518 (N_13518,N_12989,N_12971);
or U13519 (N_13519,N_12214,N_12101);
or U13520 (N_13520,N_13369,N_12321);
or U13521 (N_13521,N_12616,N_12966);
and U13522 (N_13522,N_13156,N_12898);
nand U13523 (N_13523,N_13022,N_12694);
nand U13524 (N_13524,N_12975,N_12646);
and U13525 (N_13525,N_12071,N_13125);
or U13526 (N_13526,N_13354,N_13260);
nand U13527 (N_13527,N_12617,N_12284);
xor U13528 (N_13528,N_12198,N_13217);
or U13529 (N_13529,N_12155,N_12764);
nor U13530 (N_13530,N_12389,N_12761);
or U13531 (N_13531,N_13037,N_12602);
and U13532 (N_13532,N_12638,N_12470);
nor U13533 (N_13533,N_13286,N_12405);
or U13534 (N_13534,N_12201,N_12772);
or U13535 (N_13535,N_12365,N_13328);
and U13536 (N_13536,N_12152,N_12866);
xnor U13537 (N_13537,N_12639,N_12383);
and U13538 (N_13538,N_12105,N_13207);
nand U13539 (N_13539,N_12727,N_12681);
xnor U13540 (N_13540,N_12150,N_12973);
nand U13541 (N_13541,N_12426,N_12200);
xnor U13542 (N_13542,N_13176,N_12700);
and U13543 (N_13543,N_13279,N_13385);
or U13544 (N_13544,N_12098,N_12250);
xor U13545 (N_13545,N_13122,N_13219);
and U13546 (N_13546,N_12013,N_13179);
nand U13547 (N_13547,N_13213,N_12386);
nor U13548 (N_13548,N_12099,N_13497);
and U13549 (N_13549,N_13226,N_12521);
nor U13550 (N_13550,N_12525,N_12850);
nand U13551 (N_13551,N_12628,N_12604);
nor U13552 (N_13552,N_12444,N_12636);
nand U13553 (N_13553,N_12790,N_13418);
nor U13554 (N_13554,N_12449,N_13117);
or U13555 (N_13555,N_12260,N_12766);
and U13556 (N_13556,N_12016,N_12137);
xor U13557 (N_13557,N_12401,N_12596);
and U13558 (N_13558,N_12046,N_12882);
or U13559 (N_13559,N_12356,N_13277);
or U13560 (N_13560,N_12163,N_12781);
nor U13561 (N_13561,N_12059,N_12793);
nand U13562 (N_13562,N_12582,N_12945);
nand U13563 (N_13563,N_12268,N_12317);
and U13564 (N_13564,N_12339,N_12479);
nor U13565 (N_13565,N_12635,N_12075);
and U13566 (N_13566,N_13088,N_12912);
xnor U13567 (N_13567,N_13084,N_12650);
nand U13568 (N_13568,N_12782,N_12710);
or U13569 (N_13569,N_12111,N_12474);
nor U13570 (N_13570,N_12311,N_12952);
or U13571 (N_13571,N_12141,N_13101);
or U13572 (N_13572,N_12699,N_12172);
and U13573 (N_13573,N_13359,N_13333);
or U13574 (N_13574,N_13018,N_13379);
nand U13575 (N_13575,N_12011,N_12193);
and U13576 (N_13576,N_12630,N_12951);
or U13577 (N_13577,N_12759,N_12249);
nor U13578 (N_13578,N_13490,N_12457);
or U13579 (N_13579,N_12686,N_12149);
nor U13580 (N_13580,N_12734,N_13388);
or U13581 (N_13581,N_12601,N_13325);
nand U13582 (N_13582,N_13335,N_13167);
nand U13583 (N_13583,N_13066,N_12070);
and U13584 (N_13584,N_12891,N_12134);
or U13585 (N_13585,N_12599,N_12048);
nand U13586 (N_13586,N_12432,N_12925);
nand U13587 (N_13587,N_13400,N_12998);
nor U13588 (N_13588,N_13347,N_12001);
or U13589 (N_13589,N_13240,N_13063);
or U13590 (N_13590,N_12154,N_12283);
nor U13591 (N_13591,N_12454,N_12281);
or U13592 (N_13592,N_12004,N_13368);
nand U13593 (N_13593,N_12296,N_13484);
or U13594 (N_13594,N_12063,N_12698);
xor U13595 (N_13595,N_12008,N_12667);
or U13596 (N_13596,N_12445,N_12826);
xor U13597 (N_13597,N_12682,N_13153);
nor U13598 (N_13598,N_12888,N_12805);
nor U13599 (N_13599,N_13381,N_12655);
and U13600 (N_13600,N_12371,N_12707);
and U13601 (N_13601,N_13214,N_13134);
xnor U13602 (N_13602,N_13476,N_12919);
and U13603 (N_13603,N_12695,N_12609);
or U13604 (N_13604,N_13405,N_13040);
and U13605 (N_13605,N_12418,N_12468);
and U13606 (N_13606,N_13420,N_12329);
nor U13607 (N_13607,N_12563,N_12056);
nor U13608 (N_13608,N_13269,N_12206);
or U13609 (N_13609,N_12334,N_12920);
and U13610 (N_13610,N_12871,N_12132);
and U13611 (N_13611,N_12490,N_12645);
nand U13612 (N_13612,N_12160,N_12394);
and U13613 (N_13613,N_12133,N_12855);
nand U13614 (N_13614,N_13411,N_12519);
nor U13615 (N_13615,N_12026,N_13350);
nand U13616 (N_13616,N_12522,N_12683);
xor U13617 (N_13617,N_12566,N_12740);
nor U13618 (N_13618,N_13356,N_13460);
nand U13619 (N_13619,N_13376,N_13199);
xnor U13620 (N_13620,N_13262,N_13232);
nand U13621 (N_13621,N_12554,N_12974);
nand U13622 (N_13622,N_12170,N_12262);
nand U13623 (N_13623,N_13428,N_12584);
and U13624 (N_13624,N_12520,N_12195);
and U13625 (N_13625,N_13442,N_13268);
and U13626 (N_13626,N_12382,N_12091);
or U13627 (N_13627,N_12349,N_13218);
and U13628 (N_13628,N_12300,N_12439);
and U13629 (N_13629,N_13014,N_12400);
nand U13630 (N_13630,N_12019,N_12488);
or U13631 (N_13631,N_12908,N_12406);
nor U13632 (N_13632,N_12778,N_13235);
or U13633 (N_13633,N_13449,N_12224);
nor U13634 (N_13634,N_12838,N_13160);
xnor U13635 (N_13635,N_12320,N_13427);
or U13636 (N_13636,N_12969,N_13024);
and U13637 (N_13637,N_13041,N_13104);
nand U13638 (N_13638,N_13409,N_12940);
and U13639 (N_13639,N_12392,N_12553);
or U13640 (N_13640,N_12128,N_12081);
and U13641 (N_13641,N_13194,N_12665);
and U13642 (N_13642,N_12598,N_12823);
and U13643 (N_13643,N_12179,N_13245);
and U13644 (N_13644,N_12258,N_12552);
or U13645 (N_13645,N_12947,N_13119);
nor U13646 (N_13646,N_12374,N_13284);
or U13647 (N_13647,N_13304,N_13493);
and U13648 (N_13648,N_12275,N_12226);
nand U13649 (N_13649,N_12014,N_12192);
and U13650 (N_13650,N_12165,N_13023);
nor U13651 (N_13651,N_12950,N_12096);
or U13652 (N_13652,N_12247,N_13469);
or U13653 (N_13653,N_12034,N_13013);
nand U13654 (N_13654,N_12097,N_12411);
xnor U13655 (N_13655,N_12476,N_13086);
xor U13656 (N_13656,N_13181,N_12309);
xnor U13657 (N_13657,N_13187,N_12803);
or U13658 (N_13658,N_13070,N_13271);
or U13659 (N_13659,N_12791,N_13380);
xnor U13660 (N_13660,N_12147,N_12385);
or U13661 (N_13661,N_12093,N_12215);
and U13662 (N_13662,N_12197,N_12496);
xnor U13663 (N_13663,N_12835,N_13083);
xor U13664 (N_13664,N_12469,N_12357);
nand U13665 (N_13665,N_13128,N_12836);
xor U13666 (N_13666,N_12965,N_12103);
or U13667 (N_13667,N_12350,N_12372);
or U13668 (N_13668,N_13183,N_13108);
xnor U13669 (N_13669,N_12829,N_12581);
nor U13670 (N_13670,N_12183,N_12032);
nand U13671 (N_13671,N_12813,N_13374);
nor U13672 (N_13672,N_13270,N_12410);
nor U13673 (N_13673,N_12253,N_13052);
or U13674 (N_13674,N_12252,N_13384);
nand U13675 (N_13675,N_13263,N_13238);
nor U13676 (N_13676,N_12914,N_12378);
nor U13677 (N_13677,N_12775,N_12227);
and U13678 (N_13678,N_12728,N_12946);
or U13679 (N_13679,N_12876,N_13436);
xnor U13680 (N_13680,N_12025,N_12837);
or U13681 (N_13681,N_13025,N_12769);
nor U13682 (N_13682,N_13002,N_13005);
xor U13683 (N_13683,N_12851,N_12328);
and U13684 (N_13684,N_12038,N_12676);
and U13685 (N_13685,N_12027,N_12292);
nand U13686 (N_13686,N_12771,N_12348);
or U13687 (N_13687,N_12467,N_12987);
and U13688 (N_13688,N_12934,N_13211);
or U13689 (N_13689,N_13383,N_13246);
nand U13690 (N_13690,N_12961,N_12663);
nor U13691 (N_13691,N_12369,N_13060);
nor U13692 (N_13692,N_13390,N_12425);
nand U13693 (N_13693,N_13445,N_13349);
or U13694 (N_13694,N_12176,N_12084);
nand U13695 (N_13695,N_12868,N_12344);
xor U13696 (N_13696,N_13216,N_13301);
nand U13697 (N_13697,N_12561,N_12933);
nand U13698 (N_13698,N_12669,N_12941);
and U13699 (N_13699,N_12911,N_12618);
nor U13700 (N_13700,N_12118,N_13431);
or U13701 (N_13701,N_12758,N_12433);
or U13702 (N_13702,N_13254,N_12442);
or U13703 (N_13703,N_12472,N_13239);
or U13704 (N_13704,N_13393,N_12028);
nand U13705 (N_13705,N_12594,N_13244);
and U13706 (N_13706,N_12798,N_13107);
nand U13707 (N_13707,N_12583,N_13140);
nor U13708 (N_13708,N_13265,N_13452);
nand U13709 (N_13709,N_13371,N_12662);
and U13710 (N_13710,N_12722,N_13495);
or U13711 (N_13711,N_12576,N_13451);
nand U13712 (N_13712,N_12360,N_13441);
nand U13713 (N_13713,N_12640,N_13079);
nor U13714 (N_13714,N_12023,N_12712);
or U13715 (N_13715,N_12885,N_12342);
xnor U13716 (N_13716,N_12964,N_13064);
and U13717 (N_13717,N_12867,N_12687);
and U13718 (N_13718,N_12484,N_12354);
nor U13719 (N_13719,N_12963,N_13042);
or U13720 (N_13720,N_13186,N_12634);
nor U13721 (N_13721,N_12742,N_12313);
xnor U13722 (N_13722,N_12104,N_12615);
nor U13723 (N_13723,N_12304,N_12471);
and U13724 (N_13724,N_12731,N_12658);
or U13725 (N_13725,N_12962,N_12340);
and U13726 (N_13726,N_12930,N_13486);
nand U13727 (N_13727,N_12550,N_13250);
nand U13728 (N_13728,N_12029,N_12714);
xor U13729 (N_13729,N_12337,N_12232);
and U13730 (N_13730,N_12674,N_13321);
and U13731 (N_13731,N_13424,N_12863);
and U13732 (N_13732,N_12514,N_12512);
nand U13733 (N_13733,N_13141,N_12416);
and U13734 (N_13734,N_12996,N_12960);
nand U13735 (N_13735,N_12906,N_13166);
nor U13736 (N_13736,N_13402,N_13289);
nand U13737 (N_13737,N_12802,N_12915);
nand U13738 (N_13738,N_13471,N_12331);
xnor U13739 (N_13739,N_13099,N_13299);
nand U13740 (N_13740,N_13261,N_12039);
and U13741 (N_13741,N_12431,N_12959);
nor U13742 (N_13742,N_13419,N_12624);
nand U13743 (N_13743,N_13120,N_12985);
or U13744 (N_13744,N_12086,N_12187);
nand U13745 (N_13745,N_12532,N_13296);
nand U13746 (N_13746,N_13038,N_13200);
nand U13747 (N_13747,N_13466,N_12564);
nor U13748 (N_13748,N_12345,N_12589);
and U13749 (N_13749,N_12244,N_12642);
and U13750 (N_13750,N_13144,N_13098);
nor U13751 (N_13751,N_12185,N_12573);
nand U13752 (N_13752,N_12827,N_13027);
and U13753 (N_13753,N_12286,N_13282);
nor U13754 (N_13754,N_13090,N_12862);
nand U13755 (N_13755,N_13326,N_12546);
nor U13756 (N_13756,N_13248,N_12773);
nor U13757 (N_13757,N_12629,N_12899);
nor U13758 (N_13758,N_13154,N_12818);
xor U13759 (N_13759,N_12242,N_12012);
nor U13760 (N_13760,N_12363,N_13285);
and U13761 (N_13761,N_12462,N_12225);
xnor U13762 (N_13762,N_12089,N_12361);
and U13763 (N_13763,N_12233,N_12325);
nand U13764 (N_13764,N_12709,N_12451);
nor U13765 (N_13765,N_13338,N_13257);
nor U13766 (N_13766,N_12459,N_12897);
nor U13767 (N_13767,N_13480,N_13126);
and U13768 (N_13768,N_13075,N_12733);
nand U13769 (N_13769,N_12362,N_13165);
and U13770 (N_13770,N_12235,N_12095);
and U13771 (N_13771,N_12677,N_12419);
nand U13772 (N_13772,N_12659,N_12293);
nand U13773 (N_13773,N_12979,N_12353);
nand U13774 (N_13774,N_12917,N_12992);
or U13775 (N_13775,N_12237,N_12113);
nor U13776 (N_13776,N_12127,N_13100);
nand U13777 (N_13777,N_12626,N_12050);
xnor U13778 (N_13778,N_12794,N_13209);
nand U13779 (N_13779,N_12741,N_12205);
and U13780 (N_13780,N_13311,N_12637);
or U13781 (N_13781,N_12289,N_13482);
nand U13782 (N_13782,N_12312,N_12230);
xnor U13783 (N_13783,N_12783,N_12757);
or U13784 (N_13784,N_12865,N_12976);
nand U13785 (N_13785,N_13102,N_12305);
or U13786 (N_13786,N_12387,N_12831);
or U13787 (N_13787,N_12844,N_13342);
nand U13788 (N_13788,N_12124,N_13343);
nand U13789 (N_13789,N_12009,N_12861);
nor U13790 (N_13790,N_13173,N_12115);
or U13791 (N_13791,N_13177,N_12984);
nor U13792 (N_13792,N_12592,N_12716);
xnor U13793 (N_13793,N_12267,N_13274);
nand U13794 (N_13794,N_12777,N_12248);
and U13795 (N_13795,N_12399,N_13080);
nand U13796 (N_13796,N_12792,N_12801);
xor U13797 (N_13797,N_13170,N_12749);
and U13798 (N_13798,N_12136,N_12572);
or U13799 (N_13799,N_12222,N_12273);
and U13800 (N_13800,N_13044,N_13496);
nand U13801 (N_13801,N_13017,N_13172);
and U13802 (N_13802,N_12204,N_13307);
nand U13803 (N_13803,N_13346,N_13355);
or U13804 (N_13804,N_12180,N_12010);
nor U13805 (N_13805,N_13036,N_12833);
nand U13806 (N_13806,N_12822,N_12397);
nor U13807 (N_13807,N_13230,N_12623);
and U13808 (N_13808,N_13458,N_13111);
nand U13809 (N_13809,N_12458,N_13422);
and U13810 (N_13810,N_12555,N_12367);
nor U13811 (N_13811,N_13446,N_12720);
nor U13812 (N_13812,N_12290,N_13318);
xor U13813 (N_13813,N_12788,N_13208);
nor U13814 (N_13814,N_12527,N_12144);
and U13815 (N_13815,N_12213,N_12210);
or U13816 (N_13816,N_13327,N_13201);
or U13817 (N_13817,N_13395,N_13032);
and U13818 (N_13818,N_12184,N_13416);
and U13819 (N_13819,N_12619,N_12441);
nand U13820 (N_13820,N_12421,N_12053);
nor U13821 (N_13821,N_12005,N_12703);
nor U13822 (N_13822,N_12427,N_12509);
nor U13823 (N_13823,N_12724,N_12577);
nand U13824 (N_13824,N_13241,N_13396);
xnor U13825 (N_13825,N_12526,N_12219);
or U13826 (N_13826,N_12282,N_12756);
nand U13827 (N_13827,N_12003,N_12178);
and U13828 (N_13828,N_13309,N_13375);
and U13829 (N_13829,N_13468,N_13258);
and U13830 (N_13830,N_13443,N_12825);
and U13831 (N_13831,N_12108,N_13222);
nand U13832 (N_13832,N_13103,N_13292);
or U13833 (N_13833,N_12307,N_12540);
nor U13834 (N_13834,N_13212,N_12571);
nand U13835 (N_13835,N_13288,N_12366);
and U13836 (N_13836,N_12228,N_12768);
nor U13837 (N_13837,N_13168,N_13348);
or U13838 (N_13838,N_13358,N_12955);
nor U13839 (N_13839,N_12938,N_12907);
or U13840 (N_13840,N_13295,N_12671);
nand U13841 (N_13841,N_12483,N_13363);
nor U13842 (N_13842,N_12675,N_12335);
nand U13843 (N_13843,N_12785,N_12872);
and U13844 (N_13844,N_13164,N_12087);
or U13845 (N_13845,N_12368,N_12280);
nor U13846 (N_13846,N_12738,N_12739);
nor U13847 (N_13847,N_12511,N_12043);
nand U13848 (N_13848,N_12770,N_12294);
or U13849 (N_13849,N_12988,N_12860);
or U13850 (N_13850,N_12916,N_12121);
nand U13851 (N_13851,N_13115,N_13039);
and U13852 (N_13852,N_13357,N_13378);
nor U13853 (N_13853,N_12536,N_13372);
and U13854 (N_13854,N_12875,N_12024);
nor U13855 (N_13855,N_12776,N_13129);
nand U13856 (N_13856,N_13315,N_12905);
or U13857 (N_13857,N_12751,N_13123);
or U13858 (N_13858,N_13415,N_12495);
nor U13859 (N_13859,N_12549,N_12902);
nor U13860 (N_13860,N_12900,N_13314);
nand U13861 (N_13861,N_13132,N_12593);
nand U13862 (N_13862,N_12437,N_12171);
nand U13863 (N_13863,N_12539,N_12567);
or U13864 (N_13864,N_13407,N_12452);
and U13865 (N_13865,N_12689,N_12654);
or U13866 (N_13866,N_12719,N_12610);
nand U13867 (N_13867,N_12035,N_12697);
nand U13868 (N_13868,N_12688,N_12516);
and U13869 (N_13869,N_13303,N_12660);
xnor U13870 (N_13870,N_13077,N_13344);
and U13871 (N_13871,N_12278,N_13290);
nor U13872 (N_13872,N_12100,N_12332);
or U13873 (N_13873,N_12753,N_12748);
or U13874 (N_13874,N_12114,N_12664);
nor U13875 (N_13875,N_12621,N_13252);
or U13876 (N_13876,N_13043,N_13330);
nor U13877 (N_13877,N_12212,N_12373);
nor U13878 (N_13878,N_12398,N_12843);
and U13879 (N_13879,N_12575,N_12054);
and U13880 (N_13880,N_13397,N_12981);
nor U13881 (N_13881,N_13401,N_12261);
xor U13882 (N_13882,N_12591,N_12430);
nand U13883 (N_13883,N_13437,N_12896);
or U13884 (N_13884,N_12196,N_13494);
nor U13885 (N_13885,N_12505,N_12887);
and U13886 (N_13886,N_13293,N_13399);
nor U13887 (N_13887,N_13297,N_12523);
nand U13888 (N_13888,N_12859,N_12811);
xor U13889 (N_13889,N_12568,N_12088);
nand U13890 (N_13890,N_12893,N_12143);
and U13891 (N_13891,N_12608,N_12935);
nor U13892 (N_13892,N_13197,N_12560);
nor U13893 (N_13893,N_12795,N_12082);
or U13894 (N_13894,N_12894,N_13272);
and U13895 (N_13895,N_13015,N_12221);
and U13896 (N_13896,N_13391,N_13247);
and U13897 (N_13897,N_13137,N_13465);
and U13898 (N_13898,N_12856,N_13215);
xor U13899 (N_13899,N_13011,N_12102);
xor U13900 (N_13900,N_13332,N_12611);
and U13901 (N_13901,N_13387,N_12701);
nand U13902 (N_13902,N_12763,N_13377);
and U13903 (N_13903,N_13145,N_12497);
and U13904 (N_13904,N_12853,N_12306);
nand U13905 (N_13905,N_12883,N_13227);
nand U13906 (N_13906,N_13291,N_12450);
and U13907 (N_13907,N_12943,N_12447);
or U13908 (N_13908,N_12409,N_12972);
and U13909 (N_13909,N_12338,N_12420);
nor U13910 (N_13910,N_12182,N_13298);
nor U13911 (N_13911,N_13464,N_12545);
nand U13912 (N_13912,N_12644,N_12181);
or U13913 (N_13913,N_13434,N_12393);
and U13914 (N_13914,N_12648,N_13210);
and U13915 (N_13915,N_12083,N_13065);
or U13916 (N_13916,N_13202,N_12932);
and U13917 (N_13917,N_12080,N_13142);
nand U13918 (N_13918,N_12804,N_13281);
and U13919 (N_13919,N_13483,N_12928);
xor U13920 (N_13920,N_13035,N_12809);
nand U13921 (N_13921,N_13455,N_13074);
nand U13922 (N_13922,N_12218,N_12434);
nor U13923 (N_13923,N_13435,N_12852);
xnor U13924 (N_13924,N_12291,N_12060);
nand U13925 (N_13925,N_13193,N_12239);
or U13926 (N_13926,N_12276,N_12762);
and U13927 (N_13927,N_12018,N_13453);
nor U13928 (N_13928,N_12380,N_12995);
nor U13929 (N_13929,N_12310,N_12047);
xor U13930 (N_13930,N_12847,N_12322);
nand U13931 (N_13931,N_12417,N_12504);
nand U13932 (N_13932,N_13184,N_13205);
nor U13933 (N_13933,N_12569,N_13135);
nand U13934 (N_13934,N_12997,N_12491);
or U13935 (N_13935,N_13195,N_12333);
or U13936 (N_13936,N_13082,N_12424);
nand U13937 (N_13937,N_12375,N_12877);
xnor U13938 (N_13938,N_12040,N_12548);
or U13939 (N_13939,N_13109,N_12493);
nor U13940 (N_13940,N_13362,N_12355);
or U13941 (N_13941,N_13116,N_12255);
or U13942 (N_13942,N_12797,N_12492);
and U13943 (N_13943,N_12202,N_12874);
and U13944 (N_13944,N_12473,N_13055);
and U13945 (N_13945,N_13152,N_12407);
nor U13946 (N_13946,N_13146,N_12993);
or U13947 (N_13947,N_12841,N_12120);
nand U13948 (N_13948,N_12880,N_12041);
and U13949 (N_13949,N_12585,N_12298);
nand U13950 (N_13950,N_12500,N_12174);
or U13951 (N_13951,N_13429,N_13361);
and U13952 (N_13952,N_13106,N_13426);
xor U13953 (N_13953,N_13251,N_13178);
nor U13954 (N_13954,N_12020,N_13322);
or U13955 (N_13955,N_13457,N_13139);
xnor U13956 (N_13956,N_12641,N_13169);
or U13957 (N_13957,N_13339,N_12057);
nand U13958 (N_13958,N_12287,N_13481);
nand U13959 (N_13959,N_12774,N_12747);
nand U13960 (N_13960,N_13417,N_12986);
and U13961 (N_13961,N_12007,N_12435);
or U13962 (N_13962,N_12922,N_13294);
and U13963 (N_13963,N_12343,N_12161);
nand U13964 (N_13964,N_12314,N_12869);
nor U13965 (N_13965,N_12346,N_12092);
nor U13966 (N_13966,N_12944,N_13413);
and U13967 (N_13967,N_12543,N_12649);
and U13968 (N_13968,N_13021,N_12269);
nor U13969 (N_13969,N_13155,N_12999);
and U13970 (N_13970,N_12970,N_13305);
and U13971 (N_13971,N_13477,N_12746);
nand U13972 (N_13972,N_13470,N_12953);
nor U13973 (N_13973,N_12901,N_13054);
nand U13974 (N_13974,N_13050,N_12840);
nor U13975 (N_13975,N_12381,N_12415);
nor U13976 (N_13976,N_13461,N_13454);
or U13977 (N_13977,N_13408,N_12587);
xnor U13978 (N_13978,N_12551,N_12254);
or U13979 (N_13979,N_12752,N_12884);
nor U13980 (N_13980,N_13433,N_13488);
nor U13981 (N_13981,N_13456,N_12456);
xor U13982 (N_13982,N_12743,N_12849);
and U13983 (N_13983,N_13394,N_12209);
nand U13984 (N_13984,N_13459,N_13033);
nand U13985 (N_13985,N_12590,N_13280);
nor U13986 (N_13986,N_12072,N_12806);
nand U13987 (N_13987,N_12679,N_12693);
nor U13988 (N_13988,N_13192,N_12706);
nand U13989 (N_13989,N_13068,N_12502);
and U13990 (N_13990,N_12303,N_12112);
nor U13991 (N_13991,N_12440,N_12680);
and U13992 (N_13992,N_12513,N_12559);
nor U13993 (N_13993,N_12927,N_13283);
and U13994 (N_13994,N_12515,N_12251);
nor U13995 (N_13995,N_13138,N_13485);
and U13996 (N_13996,N_13421,N_13008);
nand U13997 (N_13997,N_12318,N_12745);
and U13998 (N_13998,N_12846,N_12002);
nor U13999 (N_13999,N_13130,N_13206);
and U14000 (N_14000,N_13061,N_12983);
nand U14001 (N_14001,N_12189,N_12428);
and U14002 (N_14002,N_12169,N_12191);
or U14003 (N_14003,N_12271,N_13105);
and U14004 (N_14004,N_12461,N_13414);
or U14005 (N_14005,N_12530,N_12323);
nand U14006 (N_14006,N_12816,N_12903);
nand U14007 (N_14007,N_12243,N_12157);
nor U14008 (N_14008,N_12274,N_13386);
nor U14009 (N_14009,N_12556,N_13204);
and U14010 (N_14010,N_12625,N_12607);
and U14011 (N_14011,N_13341,N_12824);
nor U14012 (N_14012,N_13058,N_12037);
and U14013 (N_14013,N_12463,N_12537);
nor U14014 (N_14014,N_12538,N_12295);
nor U14015 (N_14015,N_12481,N_12135);
or U14016 (N_14016,N_13007,N_12090);
nand U14017 (N_14017,N_13096,N_12064);
nand U14018 (N_14018,N_13034,N_13329);
nand U14019 (N_14019,N_12238,N_13233);
and U14020 (N_14020,N_12036,N_12580);
nand U14021 (N_14021,N_12460,N_12220);
and U14022 (N_14022,N_12787,N_12156);
nand U14023 (N_14023,N_12711,N_12379);
and U14024 (N_14024,N_12633,N_13029);
or U14025 (N_14025,N_12547,N_12475);
xor U14026 (N_14026,N_12670,N_13188);
nor U14027 (N_14027,N_12767,N_12684);
nor U14028 (N_14028,N_12503,N_12858);
nor U14029 (N_14029,N_12647,N_12388);
nand U14030 (N_14030,N_12718,N_12404);
and U14031 (N_14031,N_12288,N_12842);
or U14032 (N_14032,N_12507,N_12168);
or U14033 (N_14033,N_12051,N_12166);
or U14034 (N_14034,N_12129,N_12094);
nor U14035 (N_14035,N_12968,N_13078);
nand U14036 (N_14036,N_13028,N_13091);
nor U14037 (N_14037,N_12229,N_12958);
or U14038 (N_14038,N_13228,N_13440);
and U14039 (N_14039,N_12982,N_12316);
or U14040 (N_14040,N_12498,N_13475);
nand U14041 (N_14041,N_12848,N_12078);
nand U14042 (N_14042,N_12597,N_12487);
and U14043 (N_14043,N_12508,N_13073);
nand U14044 (N_14044,N_13320,N_12881);
xor U14045 (N_14045,N_13425,N_13081);
and U14046 (N_14046,N_12923,N_13162);
xnor U14047 (N_14047,N_12510,N_13031);
nor U14048 (N_14048,N_13069,N_12123);
nand U14049 (N_14049,N_12478,N_13059);
and U14050 (N_14050,N_13191,N_13300);
and U14051 (N_14051,N_12177,N_12603);
nor U14052 (N_14052,N_12186,N_13148);
nand U14053 (N_14053,N_12839,N_12814);
nor U14054 (N_14054,N_13175,N_12125);
and U14055 (N_14055,N_12854,N_12830);
nand U14056 (N_14056,N_13317,N_12980);
xor U14057 (N_14057,N_12175,N_12750);
and U14058 (N_14058,N_13462,N_13112);
or U14059 (N_14059,N_12297,N_12408);
xor U14060 (N_14060,N_12216,N_12726);
or U14061 (N_14061,N_12453,N_12142);
or U14062 (N_14062,N_13150,N_13259);
or U14063 (N_14063,N_13174,N_12692);
nand U14064 (N_14064,N_12528,N_13474);
nor U14065 (N_14065,N_13331,N_13382);
and U14066 (N_14066,N_13275,N_12886);
or U14067 (N_14067,N_13337,N_13182);
or U14068 (N_14068,N_12263,N_12448);
nor U14069 (N_14069,N_12464,N_12485);
and U14070 (N_14070,N_12030,N_13180);
nand U14071 (N_14071,N_12391,N_12574);
or U14072 (N_14072,N_13319,N_13302);
or U14073 (N_14073,N_12892,N_12390);
and U14074 (N_14074,N_12613,N_13020);
nand U14075 (N_14075,N_12870,N_12131);
or U14076 (N_14076,N_12126,N_12494);
or U14077 (N_14077,N_13310,N_12412);
and U14078 (N_14078,N_13345,N_12815);
xnor U14079 (N_14079,N_13432,N_12194);
or U14080 (N_14080,N_13278,N_13367);
or U14081 (N_14081,N_12612,N_13221);
or U14082 (N_14082,N_12116,N_13352);
and U14083 (N_14083,N_13273,N_13092);
nand U14084 (N_14084,N_12696,N_13364);
and U14085 (N_14085,N_13256,N_13203);
and U14086 (N_14086,N_12259,N_12359);
xnor U14087 (N_14087,N_12395,N_12810);
nor U14088 (N_14088,N_13373,N_13340);
nor U14089 (N_14089,N_12489,N_12302);
xor U14090 (N_14090,N_12049,N_13229);
nand U14091 (N_14091,N_12396,N_12167);
or U14092 (N_14092,N_12236,N_12913);
nor U14093 (N_14093,N_12954,N_12614);
nand U14094 (N_14094,N_12730,N_12140);
xor U14095 (N_14095,N_12370,N_12657);
xnor U14096 (N_14096,N_12106,N_12672);
nand U14097 (N_14097,N_12246,N_13127);
or U14098 (N_14098,N_13085,N_12257);
or U14099 (N_14099,N_12529,N_12588);
nand U14100 (N_14100,N_13151,N_12936);
nor U14101 (N_14101,N_12058,N_12967);
nand U14102 (N_14102,N_13467,N_12073);
nor U14103 (N_14103,N_12673,N_12151);
nand U14104 (N_14104,N_12931,N_13010);
or U14105 (N_14105,N_13487,N_12319);
nor U14106 (N_14106,N_12377,N_12578);
nand U14107 (N_14107,N_12352,N_12808);
nand U14108 (N_14108,N_12879,N_12055);
nor U14109 (N_14109,N_12817,N_12364);
nand U14110 (N_14110,N_12110,N_12949);
nand U14111 (N_14111,N_12145,N_12465);
and U14112 (N_14112,N_12760,N_12315);
nor U14113 (N_14113,N_13438,N_12918);
and U14114 (N_14114,N_12765,N_12755);
or U14115 (N_14115,N_12729,N_13267);
or U14116 (N_14116,N_13026,N_12721);
nand U14117 (N_14117,N_12606,N_13370);
or U14118 (N_14118,N_12651,N_13463);
nand U14119 (N_14119,N_12845,N_12017);
or U14120 (N_14120,N_13121,N_12942);
and U14121 (N_14121,N_12270,N_13051);
nor U14122 (N_14122,N_12725,N_12708);
and U14123 (N_14123,N_12266,N_12702);
or U14124 (N_14124,N_13198,N_12744);
and U14125 (N_14125,N_13049,N_12044);
and U14126 (N_14126,N_13062,N_12446);
nor U14127 (N_14127,N_12241,N_13133);
and U14128 (N_14128,N_12119,N_13136);
xnor U14129 (N_14129,N_13479,N_13056);
xnor U14130 (N_14130,N_12977,N_13447);
or U14131 (N_14131,N_12939,N_12937);
and U14132 (N_14132,N_12668,N_13323);
or U14133 (N_14133,N_13113,N_12486);
and U14134 (N_14134,N_13234,N_12627);
nand U14135 (N_14135,N_12413,N_13163);
nand U14136 (N_14136,N_12820,N_12807);
or U14137 (N_14137,N_12109,N_12812);
and U14138 (N_14138,N_13223,N_13114);
or U14139 (N_14139,N_12031,N_12524);
xnor U14140 (N_14140,N_13236,N_12138);
nand U14141 (N_14141,N_12789,N_12895);
and U14142 (N_14142,N_13110,N_12605);
nand U14143 (N_14143,N_12784,N_12889);
nor U14144 (N_14144,N_12117,N_12904);
and U14145 (N_14145,N_12455,N_13001);
or U14146 (N_14146,N_12956,N_12737);
nand U14147 (N_14147,N_12327,N_12557);
or U14148 (N_14148,N_12800,N_12130);
xnor U14149 (N_14149,N_13243,N_12074);
and U14150 (N_14150,N_12857,N_12285);
nand U14151 (N_14151,N_12301,N_13171);
xor U14152 (N_14152,N_13403,N_12277);
or U14153 (N_14153,N_12506,N_12517);
nand U14154 (N_14154,N_12066,N_12565);
or U14155 (N_14155,N_13313,N_13276);
nand U14156 (N_14156,N_12643,N_12873);
xnor U14157 (N_14157,N_13006,N_12085);
nor U14158 (N_14158,N_13094,N_13316);
nor U14159 (N_14159,N_12480,N_13161);
or U14160 (N_14160,N_12022,N_12653);
or U14161 (N_14161,N_12926,N_12376);
nand U14162 (N_14162,N_13143,N_12723);
or U14163 (N_14163,N_13336,N_13489);
and U14164 (N_14164,N_13423,N_13266);
and U14165 (N_14165,N_12234,N_13147);
nor U14166 (N_14166,N_12077,N_12754);
or U14167 (N_14167,N_12203,N_12579);
nor U14168 (N_14168,N_13053,N_12533);
and U14169 (N_14169,N_12990,N_12423);
nand U14170 (N_14170,N_12531,N_13365);
nand U14171 (N_14171,N_12909,N_12336);
nor U14172 (N_14172,N_12910,N_13448);
nor U14173 (N_14173,N_12190,N_13095);
or U14174 (N_14174,N_12878,N_12042);
nand U14175 (N_14175,N_12736,N_12821);
nor U14176 (N_14176,N_12994,N_13009);
nor U14177 (N_14177,N_13224,N_12240);
and U14178 (N_14178,N_12330,N_12620);
nand U14179 (N_14179,N_13159,N_12705);
or U14180 (N_14180,N_12570,N_12541);
or U14181 (N_14181,N_12265,N_12308);
nand U14182 (N_14182,N_12199,N_12122);
or U14183 (N_14183,N_12341,N_12600);
or U14184 (N_14184,N_12208,N_12076);
xnor U14185 (N_14185,N_13057,N_12158);
nand U14186 (N_14186,N_13231,N_12786);
xor U14187 (N_14187,N_12033,N_12631);
or U14188 (N_14188,N_12324,N_12652);
nand U14189 (N_14189,N_12173,N_12403);
or U14190 (N_14190,N_12351,N_12384);
or U14191 (N_14191,N_12006,N_12832);
nand U14192 (N_14192,N_12690,N_12466);
nand U14193 (N_14193,N_13016,N_13360);
or U14194 (N_14194,N_12780,N_13087);
or U14195 (N_14195,N_13157,N_13012);
nor U14196 (N_14196,N_13499,N_13004);
and U14197 (N_14197,N_12735,N_13149);
nand U14198 (N_14198,N_12402,N_12299);
or U14199 (N_14199,N_13410,N_12264);
nand U14200 (N_14200,N_12443,N_13047);
nand U14201 (N_14201,N_12217,N_13389);
or U14202 (N_14202,N_12991,N_12929);
and U14203 (N_14203,N_12704,N_12661);
xor U14204 (N_14204,N_12207,N_12148);
and U14205 (N_14205,N_12632,N_12779);
and U14206 (N_14206,N_13306,N_13131);
nor U14207 (N_14207,N_12429,N_12477);
nor U14208 (N_14208,N_13351,N_12828);
and U14209 (N_14209,N_13444,N_13190);
nand U14210 (N_14210,N_13308,N_13366);
and U14211 (N_14211,N_12622,N_12501);
and U14212 (N_14212,N_12656,N_13430);
nor U14213 (N_14213,N_12948,N_12159);
or U14214 (N_14214,N_13312,N_13067);
and U14215 (N_14215,N_13491,N_12732);
and U14216 (N_14216,N_12713,N_13046);
or U14217 (N_14217,N_12691,N_13404);
nand U14218 (N_14218,N_12069,N_12414);
or U14219 (N_14219,N_13003,N_13019);
xor U14220 (N_14220,N_13472,N_13498);
xor U14221 (N_14221,N_13030,N_12015);
nand U14222 (N_14222,N_13492,N_12021);
nand U14223 (N_14223,N_13287,N_13392);
and U14224 (N_14224,N_13118,N_12422);
xor U14225 (N_14225,N_12921,N_12499);
or U14226 (N_14226,N_12153,N_13076);
and U14227 (N_14227,N_12586,N_12045);
nor U14228 (N_14228,N_12139,N_13406);
nand U14229 (N_14229,N_12558,N_12162);
nor U14230 (N_14230,N_13242,N_12079);
nand U14231 (N_14231,N_12000,N_12864);
and U14232 (N_14232,N_12065,N_13196);
or U14233 (N_14233,N_12799,N_13237);
nor U14234 (N_14234,N_13398,N_12188);
xor U14235 (N_14235,N_12272,N_12542);
and U14236 (N_14236,N_12482,N_13089);
nand U14237 (N_14237,N_13264,N_13412);
or U14238 (N_14238,N_13253,N_12061);
xnor U14239 (N_14239,N_13158,N_13334);
nor U14240 (N_14240,N_12358,N_13220);
nand U14241 (N_14241,N_13353,N_13324);
nand U14242 (N_14242,N_13185,N_13072);
and U14243 (N_14243,N_13189,N_12957);
and U14244 (N_14244,N_12326,N_12715);
xnor U14245 (N_14245,N_12685,N_13255);
nor U14246 (N_14246,N_12211,N_12535);
xor U14247 (N_14247,N_13000,N_12534);
and U14248 (N_14248,N_13225,N_12666);
or U14249 (N_14249,N_12245,N_12067);
nor U14250 (N_14250,N_12915,N_12170);
nor U14251 (N_14251,N_13064,N_12846);
nor U14252 (N_14252,N_13238,N_12975);
nor U14253 (N_14253,N_12054,N_12165);
and U14254 (N_14254,N_13188,N_13384);
nor U14255 (N_14255,N_12433,N_12600);
nand U14256 (N_14256,N_12750,N_13140);
and U14257 (N_14257,N_12268,N_12103);
or U14258 (N_14258,N_13284,N_12912);
nand U14259 (N_14259,N_12813,N_13357);
nor U14260 (N_14260,N_13156,N_12608);
nor U14261 (N_14261,N_12014,N_12250);
or U14262 (N_14262,N_13323,N_12924);
nor U14263 (N_14263,N_12673,N_12737);
nand U14264 (N_14264,N_12158,N_12956);
nor U14265 (N_14265,N_12707,N_13158);
or U14266 (N_14266,N_12477,N_12099);
nand U14267 (N_14267,N_13163,N_12180);
nor U14268 (N_14268,N_12742,N_12091);
nand U14269 (N_14269,N_13037,N_13410);
or U14270 (N_14270,N_12673,N_13365);
and U14271 (N_14271,N_12992,N_13043);
and U14272 (N_14272,N_13024,N_12556);
or U14273 (N_14273,N_12954,N_12943);
or U14274 (N_14274,N_13489,N_13354);
or U14275 (N_14275,N_12646,N_12334);
nor U14276 (N_14276,N_12049,N_12953);
xor U14277 (N_14277,N_12558,N_12792);
xnor U14278 (N_14278,N_13388,N_13361);
or U14279 (N_14279,N_13402,N_13201);
nor U14280 (N_14280,N_12813,N_13140);
and U14281 (N_14281,N_12002,N_13354);
and U14282 (N_14282,N_12192,N_12151);
and U14283 (N_14283,N_13358,N_12425);
nor U14284 (N_14284,N_12490,N_13040);
nand U14285 (N_14285,N_12573,N_12042);
nor U14286 (N_14286,N_13397,N_12839);
and U14287 (N_14287,N_12822,N_13468);
nor U14288 (N_14288,N_12191,N_13171);
nor U14289 (N_14289,N_12403,N_12842);
and U14290 (N_14290,N_13392,N_12176);
or U14291 (N_14291,N_13158,N_13473);
and U14292 (N_14292,N_12097,N_13337);
nand U14293 (N_14293,N_12106,N_13196);
or U14294 (N_14294,N_12736,N_13016);
nand U14295 (N_14295,N_12626,N_12041);
nand U14296 (N_14296,N_13361,N_13049);
or U14297 (N_14297,N_13358,N_12330);
and U14298 (N_14298,N_13294,N_12507);
nand U14299 (N_14299,N_12112,N_12949);
nand U14300 (N_14300,N_12564,N_12588);
and U14301 (N_14301,N_12828,N_13439);
and U14302 (N_14302,N_12740,N_12797);
nor U14303 (N_14303,N_12942,N_12201);
and U14304 (N_14304,N_12942,N_12223);
nor U14305 (N_14305,N_12839,N_12375);
and U14306 (N_14306,N_12647,N_13340);
and U14307 (N_14307,N_12569,N_12458);
nand U14308 (N_14308,N_13210,N_12484);
nand U14309 (N_14309,N_13019,N_12059);
or U14310 (N_14310,N_12672,N_12537);
and U14311 (N_14311,N_13407,N_12916);
or U14312 (N_14312,N_12152,N_13349);
nand U14313 (N_14313,N_12484,N_12721);
or U14314 (N_14314,N_12079,N_12722);
nor U14315 (N_14315,N_12282,N_13028);
or U14316 (N_14316,N_12237,N_12122);
or U14317 (N_14317,N_13192,N_12629);
or U14318 (N_14318,N_12900,N_12227);
or U14319 (N_14319,N_12558,N_12414);
and U14320 (N_14320,N_12677,N_12129);
xnor U14321 (N_14321,N_12823,N_12805);
or U14322 (N_14322,N_12239,N_12463);
xor U14323 (N_14323,N_13237,N_13362);
and U14324 (N_14324,N_13252,N_13008);
or U14325 (N_14325,N_13364,N_12284);
nand U14326 (N_14326,N_13402,N_13364);
nand U14327 (N_14327,N_13256,N_12703);
xnor U14328 (N_14328,N_13200,N_12051);
or U14329 (N_14329,N_12455,N_12860);
nor U14330 (N_14330,N_12848,N_13393);
and U14331 (N_14331,N_12737,N_12403);
or U14332 (N_14332,N_12025,N_13356);
xnor U14333 (N_14333,N_12089,N_13035);
and U14334 (N_14334,N_12267,N_12525);
nor U14335 (N_14335,N_12994,N_12998);
and U14336 (N_14336,N_12731,N_12583);
nand U14337 (N_14337,N_12763,N_12157);
nor U14338 (N_14338,N_12078,N_13050);
and U14339 (N_14339,N_12733,N_12618);
and U14340 (N_14340,N_12844,N_13389);
nor U14341 (N_14341,N_13251,N_12540);
or U14342 (N_14342,N_12014,N_13274);
or U14343 (N_14343,N_12460,N_12018);
or U14344 (N_14344,N_12969,N_12647);
and U14345 (N_14345,N_12759,N_12669);
or U14346 (N_14346,N_12636,N_12541);
and U14347 (N_14347,N_12135,N_12063);
nor U14348 (N_14348,N_13220,N_12465);
nand U14349 (N_14349,N_13091,N_12375);
nor U14350 (N_14350,N_12116,N_13017);
and U14351 (N_14351,N_12892,N_13453);
and U14352 (N_14352,N_13341,N_12460);
nor U14353 (N_14353,N_12825,N_12001);
and U14354 (N_14354,N_12229,N_12792);
nand U14355 (N_14355,N_12780,N_12788);
or U14356 (N_14356,N_12703,N_13125);
and U14357 (N_14357,N_12733,N_12201);
xnor U14358 (N_14358,N_12552,N_12544);
nor U14359 (N_14359,N_12293,N_12840);
and U14360 (N_14360,N_13011,N_13261);
and U14361 (N_14361,N_12980,N_12412);
or U14362 (N_14362,N_12739,N_13439);
and U14363 (N_14363,N_13099,N_12068);
and U14364 (N_14364,N_12625,N_13408);
xor U14365 (N_14365,N_12623,N_12898);
nor U14366 (N_14366,N_13058,N_13438);
nand U14367 (N_14367,N_13414,N_12849);
or U14368 (N_14368,N_12141,N_12264);
and U14369 (N_14369,N_13408,N_12494);
nand U14370 (N_14370,N_12270,N_13114);
or U14371 (N_14371,N_13039,N_13260);
or U14372 (N_14372,N_12921,N_12616);
xnor U14373 (N_14373,N_12908,N_12456);
or U14374 (N_14374,N_13393,N_12529);
nor U14375 (N_14375,N_13360,N_12094);
or U14376 (N_14376,N_13482,N_12680);
nand U14377 (N_14377,N_12794,N_13285);
or U14378 (N_14378,N_13461,N_12306);
nand U14379 (N_14379,N_12247,N_12608);
or U14380 (N_14380,N_12894,N_12794);
nor U14381 (N_14381,N_13218,N_12717);
nor U14382 (N_14382,N_13346,N_12418);
nand U14383 (N_14383,N_12323,N_13471);
and U14384 (N_14384,N_13243,N_12336);
and U14385 (N_14385,N_12080,N_13158);
or U14386 (N_14386,N_12084,N_12357);
xor U14387 (N_14387,N_13153,N_12746);
and U14388 (N_14388,N_12583,N_12430);
and U14389 (N_14389,N_13423,N_12707);
nand U14390 (N_14390,N_12808,N_13109);
xor U14391 (N_14391,N_13283,N_12199);
nand U14392 (N_14392,N_12465,N_12100);
xor U14393 (N_14393,N_13279,N_12874);
nand U14394 (N_14394,N_12770,N_13301);
and U14395 (N_14395,N_12363,N_12977);
nand U14396 (N_14396,N_12032,N_12499);
nand U14397 (N_14397,N_12843,N_12630);
and U14398 (N_14398,N_12389,N_12367);
nor U14399 (N_14399,N_13426,N_12216);
and U14400 (N_14400,N_12689,N_12856);
or U14401 (N_14401,N_12861,N_12294);
nor U14402 (N_14402,N_12902,N_12832);
or U14403 (N_14403,N_12014,N_13488);
nand U14404 (N_14404,N_13262,N_12361);
nand U14405 (N_14405,N_12962,N_12616);
nor U14406 (N_14406,N_13403,N_12171);
nor U14407 (N_14407,N_13407,N_12913);
or U14408 (N_14408,N_12304,N_12248);
nor U14409 (N_14409,N_12581,N_12344);
nand U14410 (N_14410,N_13238,N_12729);
or U14411 (N_14411,N_13323,N_13280);
nand U14412 (N_14412,N_13435,N_12686);
nor U14413 (N_14413,N_12566,N_12483);
or U14414 (N_14414,N_12959,N_12626);
xor U14415 (N_14415,N_12989,N_12609);
or U14416 (N_14416,N_12265,N_12981);
nand U14417 (N_14417,N_12787,N_13050);
nor U14418 (N_14418,N_13180,N_12016);
or U14419 (N_14419,N_12216,N_12456);
nand U14420 (N_14420,N_12570,N_12762);
nor U14421 (N_14421,N_13152,N_13221);
nor U14422 (N_14422,N_12833,N_12126);
nand U14423 (N_14423,N_12125,N_12565);
or U14424 (N_14424,N_12829,N_12781);
or U14425 (N_14425,N_13033,N_12490);
nand U14426 (N_14426,N_13175,N_12692);
and U14427 (N_14427,N_12458,N_12055);
nor U14428 (N_14428,N_13379,N_12645);
or U14429 (N_14429,N_13340,N_13226);
nand U14430 (N_14430,N_12279,N_12158);
nor U14431 (N_14431,N_13207,N_12405);
nand U14432 (N_14432,N_13419,N_12347);
or U14433 (N_14433,N_13220,N_12052);
and U14434 (N_14434,N_13321,N_12889);
nor U14435 (N_14435,N_13093,N_13263);
xnor U14436 (N_14436,N_12712,N_12327);
nand U14437 (N_14437,N_13335,N_13258);
or U14438 (N_14438,N_12624,N_12515);
nand U14439 (N_14439,N_12244,N_13286);
nor U14440 (N_14440,N_12788,N_13306);
or U14441 (N_14441,N_12520,N_13075);
or U14442 (N_14442,N_12383,N_13403);
nor U14443 (N_14443,N_12478,N_12620);
or U14444 (N_14444,N_12053,N_12433);
nor U14445 (N_14445,N_12418,N_12478);
nand U14446 (N_14446,N_12185,N_12002);
xnor U14447 (N_14447,N_12458,N_12263);
and U14448 (N_14448,N_13242,N_13143);
or U14449 (N_14449,N_13432,N_12270);
and U14450 (N_14450,N_12461,N_13276);
and U14451 (N_14451,N_12004,N_12691);
xor U14452 (N_14452,N_13079,N_13406);
nor U14453 (N_14453,N_13013,N_12783);
or U14454 (N_14454,N_12486,N_12176);
nor U14455 (N_14455,N_13070,N_12341);
and U14456 (N_14456,N_13343,N_13297);
or U14457 (N_14457,N_12033,N_13197);
or U14458 (N_14458,N_12148,N_13437);
and U14459 (N_14459,N_13168,N_12398);
and U14460 (N_14460,N_12960,N_12858);
nor U14461 (N_14461,N_12825,N_12713);
or U14462 (N_14462,N_13063,N_12884);
nand U14463 (N_14463,N_12803,N_12934);
nor U14464 (N_14464,N_12531,N_12452);
or U14465 (N_14465,N_12988,N_13349);
nor U14466 (N_14466,N_13179,N_12435);
nand U14467 (N_14467,N_12355,N_12142);
and U14468 (N_14468,N_12301,N_12873);
or U14469 (N_14469,N_12658,N_12341);
and U14470 (N_14470,N_12664,N_13136);
or U14471 (N_14471,N_13127,N_12953);
nor U14472 (N_14472,N_12606,N_13157);
xor U14473 (N_14473,N_13091,N_12922);
xnor U14474 (N_14474,N_12868,N_13291);
and U14475 (N_14475,N_12029,N_12806);
nor U14476 (N_14476,N_12281,N_12684);
nor U14477 (N_14477,N_13128,N_12001);
nor U14478 (N_14478,N_13081,N_12947);
nand U14479 (N_14479,N_12406,N_12806);
nor U14480 (N_14480,N_12960,N_13100);
and U14481 (N_14481,N_12149,N_13377);
xor U14482 (N_14482,N_13421,N_12909);
nor U14483 (N_14483,N_13381,N_12041);
xnor U14484 (N_14484,N_12995,N_12958);
nor U14485 (N_14485,N_12434,N_12641);
or U14486 (N_14486,N_12475,N_12436);
and U14487 (N_14487,N_12569,N_12958);
nor U14488 (N_14488,N_12109,N_12851);
nand U14489 (N_14489,N_13291,N_12263);
nand U14490 (N_14490,N_12882,N_12508);
nand U14491 (N_14491,N_12627,N_13008);
and U14492 (N_14492,N_12392,N_12246);
nor U14493 (N_14493,N_13166,N_12881);
and U14494 (N_14494,N_12259,N_12204);
or U14495 (N_14495,N_12595,N_13403);
nand U14496 (N_14496,N_13002,N_12373);
nor U14497 (N_14497,N_12959,N_12325);
nor U14498 (N_14498,N_12058,N_12497);
and U14499 (N_14499,N_12615,N_12530);
and U14500 (N_14500,N_12474,N_12437);
and U14501 (N_14501,N_12632,N_12962);
and U14502 (N_14502,N_13373,N_13116);
nor U14503 (N_14503,N_12055,N_13436);
nor U14504 (N_14504,N_13243,N_12594);
and U14505 (N_14505,N_12461,N_13326);
or U14506 (N_14506,N_12980,N_12704);
and U14507 (N_14507,N_12973,N_13207);
nor U14508 (N_14508,N_13282,N_12083);
xnor U14509 (N_14509,N_12543,N_13195);
xor U14510 (N_14510,N_12465,N_12558);
nor U14511 (N_14511,N_12721,N_13397);
nand U14512 (N_14512,N_12975,N_12372);
nand U14513 (N_14513,N_12181,N_12209);
or U14514 (N_14514,N_13148,N_12885);
xnor U14515 (N_14515,N_12526,N_12108);
nor U14516 (N_14516,N_12873,N_12256);
nor U14517 (N_14517,N_12107,N_12292);
or U14518 (N_14518,N_12224,N_12622);
nand U14519 (N_14519,N_13413,N_13432);
and U14520 (N_14520,N_13278,N_13201);
and U14521 (N_14521,N_12741,N_12390);
nand U14522 (N_14522,N_13083,N_13000);
xnor U14523 (N_14523,N_12508,N_12980);
xnor U14524 (N_14524,N_12625,N_12562);
or U14525 (N_14525,N_13453,N_12495);
and U14526 (N_14526,N_13206,N_13166);
and U14527 (N_14527,N_13056,N_12663);
nand U14528 (N_14528,N_12419,N_12527);
nor U14529 (N_14529,N_12065,N_12756);
nor U14530 (N_14530,N_13461,N_13073);
or U14531 (N_14531,N_12606,N_13392);
nand U14532 (N_14532,N_12205,N_12752);
or U14533 (N_14533,N_12084,N_12589);
and U14534 (N_14534,N_13464,N_13034);
or U14535 (N_14535,N_12711,N_13160);
nand U14536 (N_14536,N_12297,N_13111);
and U14537 (N_14537,N_13264,N_12308);
nor U14538 (N_14538,N_12989,N_12535);
or U14539 (N_14539,N_13251,N_12361);
and U14540 (N_14540,N_12606,N_13292);
nor U14541 (N_14541,N_13273,N_12564);
and U14542 (N_14542,N_12435,N_12417);
nand U14543 (N_14543,N_12070,N_13260);
or U14544 (N_14544,N_13097,N_12625);
nor U14545 (N_14545,N_12919,N_12447);
or U14546 (N_14546,N_12183,N_12007);
nand U14547 (N_14547,N_13272,N_12984);
nand U14548 (N_14548,N_13052,N_12012);
nor U14549 (N_14549,N_12396,N_12828);
or U14550 (N_14550,N_12897,N_13314);
xnor U14551 (N_14551,N_13076,N_13316);
or U14552 (N_14552,N_12382,N_12601);
nor U14553 (N_14553,N_12510,N_12837);
or U14554 (N_14554,N_13272,N_12075);
or U14555 (N_14555,N_12959,N_13129);
xor U14556 (N_14556,N_12680,N_12540);
or U14557 (N_14557,N_12328,N_12149);
nor U14558 (N_14558,N_12183,N_13098);
or U14559 (N_14559,N_13475,N_12956);
nand U14560 (N_14560,N_13415,N_13350);
xor U14561 (N_14561,N_13382,N_13456);
nand U14562 (N_14562,N_13082,N_12691);
xor U14563 (N_14563,N_12807,N_13446);
nor U14564 (N_14564,N_13082,N_12933);
nand U14565 (N_14565,N_13170,N_12373);
or U14566 (N_14566,N_12420,N_12951);
and U14567 (N_14567,N_12153,N_12089);
nand U14568 (N_14568,N_12762,N_12842);
nand U14569 (N_14569,N_12459,N_13218);
and U14570 (N_14570,N_13426,N_12320);
nor U14571 (N_14571,N_12086,N_13270);
nor U14572 (N_14572,N_12853,N_12652);
nand U14573 (N_14573,N_12180,N_12012);
nand U14574 (N_14574,N_12118,N_13044);
or U14575 (N_14575,N_12166,N_12694);
and U14576 (N_14576,N_13487,N_12588);
nand U14577 (N_14577,N_13139,N_12602);
or U14578 (N_14578,N_12903,N_13102);
nand U14579 (N_14579,N_13471,N_13127);
nor U14580 (N_14580,N_12667,N_12774);
or U14581 (N_14581,N_13349,N_12679);
xor U14582 (N_14582,N_12330,N_12744);
nand U14583 (N_14583,N_13066,N_12506);
nor U14584 (N_14584,N_12879,N_12564);
and U14585 (N_14585,N_12384,N_12368);
or U14586 (N_14586,N_12485,N_12470);
nand U14587 (N_14587,N_12773,N_12472);
nor U14588 (N_14588,N_13151,N_12628);
nor U14589 (N_14589,N_12055,N_12361);
and U14590 (N_14590,N_12958,N_12584);
or U14591 (N_14591,N_13050,N_12760);
nand U14592 (N_14592,N_12295,N_12939);
nor U14593 (N_14593,N_12378,N_12411);
nor U14594 (N_14594,N_13318,N_12187);
or U14595 (N_14595,N_12378,N_12623);
nor U14596 (N_14596,N_13458,N_12984);
nand U14597 (N_14597,N_12646,N_12846);
nand U14598 (N_14598,N_12489,N_12154);
or U14599 (N_14599,N_12193,N_12088);
nand U14600 (N_14600,N_12570,N_12575);
xnor U14601 (N_14601,N_12512,N_12191);
or U14602 (N_14602,N_12205,N_13213);
nand U14603 (N_14603,N_12457,N_13171);
or U14604 (N_14604,N_13237,N_12198);
and U14605 (N_14605,N_13466,N_12732);
or U14606 (N_14606,N_12880,N_12980);
or U14607 (N_14607,N_13314,N_12652);
nand U14608 (N_14608,N_12949,N_12393);
or U14609 (N_14609,N_12698,N_13189);
nor U14610 (N_14610,N_12295,N_13353);
nor U14611 (N_14611,N_12348,N_13389);
or U14612 (N_14612,N_12798,N_12818);
and U14613 (N_14613,N_13254,N_12589);
nor U14614 (N_14614,N_13366,N_12557);
or U14615 (N_14615,N_12623,N_12023);
and U14616 (N_14616,N_12585,N_12068);
nor U14617 (N_14617,N_12896,N_12665);
nand U14618 (N_14618,N_12658,N_12500);
nand U14619 (N_14619,N_12705,N_12559);
nor U14620 (N_14620,N_12738,N_12576);
and U14621 (N_14621,N_12692,N_12593);
xor U14622 (N_14622,N_13291,N_13364);
and U14623 (N_14623,N_12270,N_13487);
and U14624 (N_14624,N_13466,N_12084);
xor U14625 (N_14625,N_13448,N_12380);
nor U14626 (N_14626,N_12393,N_12124);
nand U14627 (N_14627,N_12022,N_12167);
or U14628 (N_14628,N_12244,N_12173);
xnor U14629 (N_14629,N_12726,N_12593);
or U14630 (N_14630,N_12956,N_13073);
nor U14631 (N_14631,N_13219,N_12268);
and U14632 (N_14632,N_12536,N_12192);
nand U14633 (N_14633,N_12735,N_12109);
and U14634 (N_14634,N_13216,N_12369);
nor U14635 (N_14635,N_12734,N_13301);
xnor U14636 (N_14636,N_12521,N_12536);
nand U14637 (N_14637,N_12113,N_12849);
or U14638 (N_14638,N_12772,N_13327);
nand U14639 (N_14639,N_12110,N_13354);
nand U14640 (N_14640,N_12028,N_12033);
nor U14641 (N_14641,N_12192,N_13030);
nand U14642 (N_14642,N_13378,N_13460);
and U14643 (N_14643,N_12762,N_13486);
nor U14644 (N_14644,N_13326,N_12763);
and U14645 (N_14645,N_12566,N_12860);
or U14646 (N_14646,N_12491,N_13191);
nand U14647 (N_14647,N_12130,N_12043);
and U14648 (N_14648,N_13118,N_12958);
and U14649 (N_14649,N_12090,N_13274);
nand U14650 (N_14650,N_12272,N_13447);
xnor U14651 (N_14651,N_13420,N_13179);
and U14652 (N_14652,N_12469,N_12344);
nand U14653 (N_14653,N_12586,N_13381);
nor U14654 (N_14654,N_13366,N_13373);
and U14655 (N_14655,N_13137,N_13222);
nand U14656 (N_14656,N_12035,N_12496);
nand U14657 (N_14657,N_12484,N_12249);
or U14658 (N_14658,N_12223,N_13049);
nand U14659 (N_14659,N_12198,N_12235);
nor U14660 (N_14660,N_13018,N_13131);
or U14661 (N_14661,N_12335,N_12796);
nand U14662 (N_14662,N_12789,N_12976);
nor U14663 (N_14663,N_12823,N_13146);
nor U14664 (N_14664,N_12362,N_13091);
and U14665 (N_14665,N_13117,N_12471);
nand U14666 (N_14666,N_13025,N_12563);
or U14667 (N_14667,N_13240,N_12178);
or U14668 (N_14668,N_13439,N_12230);
and U14669 (N_14669,N_12350,N_13189);
and U14670 (N_14670,N_13440,N_12717);
xnor U14671 (N_14671,N_12325,N_12298);
xor U14672 (N_14672,N_13127,N_12935);
and U14673 (N_14673,N_12887,N_12525);
and U14674 (N_14674,N_12871,N_13353);
and U14675 (N_14675,N_12039,N_13118);
nor U14676 (N_14676,N_13194,N_12588);
and U14677 (N_14677,N_13391,N_12279);
or U14678 (N_14678,N_13007,N_13343);
or U14679 (N_14679,N_13114,N_12871);
nand U14680 (N_14680,N_12278,N_12803);
and U14681 (N_14681,N_12863,N_12997);
or U14682 (N_14682,N_12150,N_13475);
and U14683 (N_14683,N_12129,N_12039);
and U14684 (N_14684,N_12908,N_12330);
or U14685 (N_14685,N_12535,N_12813);
or U14686 (N_14686,N_12511,N_13440);
nor U14687 (N_14687,N_12177,N_13372);
and U14688 (N_14688,N_12609,N_12373);
nor U14689 (N_14689,N_13093,N_12643);
nor U14690 (N_14690,N_13375,N_12178);
and U14691 (N_14691,N_12042,N_13263);
and U14692 (N_14692,N_12472,N_13084);
xnor U14693 (N_14693,N_13260,N_12288);
nand U14694 (N_14694,N_12959,N_12101);
and U14695 (N_14695,N_12639,N_13442);
nand U14696 (N_14696,N_13492,N_12318);
and U14697 (N_14697,N_12673,N_12494);
or U14698 (N_14698,N_13123,N_12585);
or U14699 (N_14699,N_12316,N_12916);
xnor U14700 (N_14700,N_13237,N_13188);
and U14701 (N_14701,N_12423,N_12322);
and U14702 (N_14702,N_12974,N_13423);
xnor U14703 (N_14703,N_12122,N_13332);
nor U14704 (N_14704,N_13132,N_12677);
or U14705 (N_14705,N_13248,N_13351);
xnor U14706 (N_14706,N_12618,N_12020);
and U14707 (N_14707,N_13347,N_12043);
or U14708 (N_14708,N_12735,N_13380);
nand U14709 (N_14709,N_12750,N_12332);
nor U14710 (N_14710,N_12398,N_12422);
nand U14711 (N_14711,N_13091,N_12487);
nor U14712 (N_14712,N_12998,N_12923);
nor U14713 (N_14713,N_13233,N_13242);
or U14714 (N_14714,N_12018,N_12378);
or U14715 (N_14715,N_12599,N_13000);
xnor U14716 (N_14716,N_13058,N_13127);
and U14717 (N_14717,N_12596,N_13490);
nor U14718 (N_14718,N_13488,N_13206);
and U14719 (N_14719,N_13448,N_13457);
nand U14720 (N_14720,N_12059,N_12722);
or U14721 (N_14721,N_12041,N_12285);
nor U14722 (N_14722,N_13179,N_12639);
nor U14723 (N_14723,N_12934,N_13377);
or U14724 (N_14724,N_13430,N_12941);
xnor U14725 (N_14725,N_12800,N_12538);
nand U14726 (N_14726,N_12794,N_12591);
nor U14727 (N_14727,N_12673,N_13332);
nor U14728 (N_14728,N_13462,N_12871);
and U14729 (N_14729,N_13425,N_12013);
nor U14730 (N_14730,N_12808,N_12299);
and U14731 (N_14731,N_13296,N_12345);
or U14732 (N_14732,N_12837,N_13342);
nand U14733 (N_14733,N_12078,N_13288);
or U14734 (N_14734,N_12771,N_12362);
nor U14735 (N_14735,N_12678,N_12482);
nand U14736 (N_14736,N_12464,N_13356);
nor U14737 (N_14737,N_13223,N_12838);
or U14738 (N_14738,N_13470,N_13281);
and U14739 (N_14739,N_13010,N_12868);
nand U14740 (N_14740,N_12920,N_12888);
nor U14741 (N_14741,N_13032,N_12807);
xnor U14742 (N_14742,N_12820,N_12052);
and U14743 (N_14743,N_12852,N_12987);
xnor U14744 (N_14744,N_12998,N_12285);
or U14745 (N_14745,N_13474,N_12192);
nand U14746 (N_14746,N_12677,N_12305);
nor U14747 (N_14747,N_12615,N_12045);
xnor U14748 (N_14748,N_12984,N_12210);
and U14749 (N_14749,N_12629,N_12631);
xnor U14750 (N_14750,N_12703,N_12292);
nor U14751 (N_14751,N_12488,N_13305);
xnor U14752 (N_14752,N_12436,N_12078);
nand U14753 (N_14753,N_12972,N_13083);
nor U14754 (N_14754,N_12424,N_13221);
or U14755 (N_14755,N_13458,N_12486);
nor U14756 (N_14756,N_12761,N_13469);
nor U14757 (N_14757,N_13253,N_13175);
xnor U14758 (N_14758,N_12929,N_13018);
nor U14759 (N_14759,N_12392,N_12777);
nor U14760 (N_14760,N_13133,N_12016);
nand U14761 (N_14761,N_12988,N_12372);
nor U14762 (N_14762,N_12843,N_13056);
nor U14763 (N_14763,N_13342,N_12596);
nand U14764 (N_14764,N_13299,N_13417);
or U14765 (N_14765,N_13211,N_12743);
or U14766 (N_14766,N_12868,N_13151);
nor U14767 (N_14767,N_12511,N_13287);
nand U14768 (N_14768,N_12479,N_12173);
or U14769 (N_14769,N_12071,N_13155);
nor U14770 (N_14770,N_12678,N_12869);
nand U14771 (N_14771,N_12247,N_13136);
nor U14772 (N_14772,N_13323,N_13262);
nand U14773 (N_14773,N_12384,N_12602);
and U14774 (N_14774,N_12030,N_12292);
xor U14775 (N_14775,N_13175,N_12411);
nand U14776 (N_14776,N_12351,N_12675);
nand U14777 (N_14777,N_12135,N_12397);
nor U14778 (N_14778,N_12151,N_12686);
or U14779 (N_14779,N_13398,N_12723);
nor U14780 (N_14780,N_12125,N_13298);
nor U14781 (N_14781,N_12155,N_13252);
and U14782 (N_14782,N_13229,N_12689);
xor U14783 (N_14783,N_12602,N_12555);
nand U14784 (N_14784,N_13417,N_13359);
or U14785 (N_14785,N_13012,N_12258);
or U14786 (N_14786,N_13372,N_12349);
nor U14787 (N_14787,N_13356,N_12953);
or U14788 (N_14788,N_12540,N_13007);
nand U14789 (N_14789,N_12115,N_12312);
nor U14790 (N_14790,N_13366,N_12666);
nand U14791 (N_14791,N_12752,N_12277);
nand U14792 (N_14792,N_12578,N_12171);
or U14793 (N_14793,N_13109,N_13017);
nand U14794 (N_14794,N_13357,N_12050);
nand U14795 (N_14795,N_12987,N_12007);
nor U14796 (N_14796,N_13007,N_12645);
or U14797 (N_14797,N_12760,N_12194);
or U14798 (N_14798,N_12555,N_12521);
and U14799 (N_14799,N_13342,N_12597);
or U14800 (N_14800,N_13486,N_12597);
nor U14801 (N_14801,N_12552,N_12071);
or U14802 (N_14802,N_13407,N_13461);
nor U14803 (N_14803,N_13205,N_13485);
and U14804 (N_14804,N_12224,N_13232);
or U14805 (N_14805,N_12918,N_13330);
and U14806 (N_14806,N_12198,N_12519);
nand U14807 (N_14807,N_13226,N_12145);
nor U14808 (N_14808,N_12138,N_12814);
or U14809 (N_14809,N_12898,N_12674);
xor U14810 (N_14810,N_13489,N_12377);
or U14811 (N_14811,N_12084,N_13348);
and U14812 (N_14812,N_12269,N_12402);
and U14813 (N_14813,N_13069,N_12698);
or U14814 (N_14814,N_12605,N_12347);
nand U14815 (N_14815,N_12380,N_12976);
and U14816 (N_14816,N_13265,N_13239);
xor U14817 (N_14817,N_12301,N_12648);
and U14818 (N_14818,N_13366,N_13128);
and U14819 (N_14819,N_13220,N_12054);
or U14820 (N_14820,N_12760,N_12737);
and U14821 (N_14821,N_12502,N_12935);
xnor U14822 (N_14822,N_12512,N_12640);
nand U14823 (N_14823,N_12099,N_12094);
xor U14824 (N_14824,N_13237,N_12807);
xor U14825 (N_14825,N_13172,N_13240);
or U14826 (N_14826,N_13343,N_13374);
and U14827 (N_14827,N_12352,N_13484);
nand U14828 (N_14828,N_13018,N_12206);
nor U14829 (N_14829,N_12478,N_12101);
or U14830 (N_14830,N_12367,N_12182);
nand U14831 (N_14831,N_12239,N_12306);
nand U14832 (N_14832,N_13075,N_12932);
nor U14833 (N_14833,N_13492,N_12771);
nor U14834 (N_14834,N_12242,N_12059);
or U14835 (N_14835,N_12538,N_13328);
and U14836 (N_14836,N_12424,N_12537);
nand U14837 (N_14837,N_13310,N_12452);
nor U14838 (N_14838,N_12120,N_12836);
or U14839 (N_14839,N_12454,N_12633);
and U14840 (N_14840,N_12319,N_13144);
xnor U14841 (N_14841,N_12651,N_12392);
and U14842 (N_14842,N_12115,N_12666);
and U14843 (N_14843,N_12629,N_13172);
and U14844 (N_14844,N_13306,N_13248);
and U14845 (N_14845,N_12180,N_12621);
or U14846 (N_14846,N_12310,N_12134);
nand U14847 (N_14847,N_12896,N_12849);
nor U14848 (N_14848,N_12351,N_12980);
and U14849 (N_14849,N_12900,N_12464);
and U14850 (N_14850,N_12598,N_12882);
nor U14851 (N_14851,N_12443,N_13077);
nor U14852 (N_14852,N_13449,N_12935);
nor U14853 (N_14853,N_12156,N_13414);
nand U14854 (N_14854,N_12614,N_12608);
nor U14855 (N_14855,N_13297,N_12341);
nor U14856 (N_14856,N_12206,N_12998);
or U14857 (N_14857,N_12729,N_13059);
and U14858 (N_14858,N_12030,N_12862);
nand U14859 (N_14859,N_12208,N_12240);
nand U14860 (N_14860,N_13226,N_12468);
and U14861 (N_14861,N_12066,N_13047);
xor U14862 (N_14862,N_12026,N_12390);
or U14863 (N_14863,N_12852,N_12284);
or U14864 (N_14864,N_12313,N_12943);
or U14865 (N_14865,N_12510,N_13237);
or U14866 (N_14866,N_13067,N_13174);
xor U14867 (N_14867,N_12698,N_12826);
or U14868 (N_14868,N_12710,N_12832);
xor U14869 (N_14869,N_13449,N_12296);
nand U14870 (N_14870,N_12440,N_12098);
or U14871 (N_14871,N_12048,N_12505);
and U14872 (N_14872,N_12041,N_12179);
nor U14873 (N_14873,N_12630,N_12065);
or U14874 (N_14874,N_12035,N_13040);
or U14875 (N_14875,N_12186,N_13195);
and U14876 (N_14876,N_13354,N_12533);
nand U14877 (N_14877,N_13042,N_12109);
or U14878 (N_14878,N_13125,N_12538);
nor U14879 (N_14879,N_12252,N_13448);
nor U14880 (N_14880,N_12611,N_12766);
nor U14881 (N_14881,N_12437,N_12840);
and U14882 (N_14882,N_12091,N_12598);
nor U14883 (N_14883,N_12169,N_12374);
nor U14884 (N_14884,N_12342,N_12836);
nand U14885 (N_14885,N_13035,N_12521);
or U14886 (N_14886,N_12582,N_13320);
nor U14887 (N_14887,N_12525,N_12218);
and U14888 (N_14888,N_13036,N_12651);
nor U14889 (N_14889,N_12975,N_12185);
nand U14890 (N_14890,N_12089,N_12170);
nand U14891 (N_14891,N_13123,N_12432);
nand U14892 (N_14892,N_13413,N_13287);
and U14893 (N_14893,N_12885,N_12727);
xor U14894 (N_14894,N_13445,N_13122);
nand U14895 (N_14895,N_12481,N_12774);
and U14896 (N_14896,N_12225,N_12800);
nand U14897 (N_14897,N_12897,N_12542);
nor U14898 (N_14898,N_13178,N_12472);
nand U14899 (N_14899,N_12001,N_12639);
or U14900 (N_14900,N_12541,N_13088);
xor U14901 (N_14901,N_12116,N_12474);
nor U14902 (N_14902,N_12600,N_12220);
nor U14903 (N_14903,N_12586,N_13080);
and U14904 (N_14904,N_12407,N_12244);
nor U14905 (N_14905,N_12248,N_12355);
or U14906 (N_14906,N_12685,N_13060);
nor U14907 (N_14907,N_12526,N_12185);
or U14908 (N_14908,N_12348,N_13404);
and U14909 (N_14909,N_12618,N_12016);
and U14910 (N_14910,N_12284,N_12602);
nor U14911 (N_14911,N_12385,N_13181);
nand U14912 (N_14912,N_12817,N_12470);
nand U14913 (N_14913,N_12909,N_12497);
and U14914 (N_14914,N_13268,N_12653);
nand U14915 (N_14915,N_13403,N_13472);
or U14916 (N_14916,N_13092,N_12523);
nand U14917 (N_14917,N_12078,N_13474);
nand U14918 (N_14918,N_12470,N_12459);
and U14919 (N_14919,N_13032,N_12425);
nor U14920 (N_14920,N_12523,N_13050);
and U14921 (N_14921,N_12841,N_13491);
nor U14922 (N_14922,N_13019,N_12617);
and U14923 (N_14923,N_13264,N_12406);
xor U14924 (N_14924,N_12757,N_13115);
nand U14925 (N_14925,N_13022,N_12688);
and U14926 (N_14926,N_13080,N_12026);
nor U14927 (N_14927,N_12061,N_13080);
or U14928 (N_14928,N_12280,N_13130);
nand U14929 (N_14929,N_12350,N_12633);
or U14930 (N_14930,N_13314,N_13492);
nor U14931 (N_14931,N_12281,N_12119);
nand U14932 (N_14932,N_12225,N_13216);
xor U14933 (N_14933,N_12556,N_12996);
and U14934 (N_14934,N_12109,N_13246);
or U14935 (N_14935,N_13117,N_13402);
and U14936 (N_14936,N_13024,N_13063);
nor U14937 (N_14937,N_12265,N_12653);
and U14938 (N_14938,N_13043,N_12557);
or U14939 (N_14939,N_12715,N_12174);
nor U14940 (N_14940,N_13126,N_12056);
and U14941 (N_14941,N_12043,N_13136);
or U14942 (N_14942,N_12191,N_12314);
or U14943 (N_14943,N_12948,N_13444);
and U14944 (N_14944,N_12661,N_12884);
or U14945 (N_14945,N_13043,N_13350);
xnor U14946 (N_14946,N_13285,N_12583);
or U14947 (N_14947,N_12728,N_12546);
xnor U14948 (N_14948,N_12177,N_13122);
nand U14949 (N_14949,N_13055,N_12963);
and U14950 (N_14950,N_12273,N_13227);
nor U14951 (N_14951,N_13127,N_12578);
or U14952 (N_14952,N_12522,N_12441);
nand U14953 (N_14953,N_13362,N_12384);
nand U14954 (N_14954,N_12334,N_12210);
nor U14955 (N_14955,N_12977,N_13436);
or U14956 (N_14956,N_13059,N_13049);
nor U14957 (N_14957,N_12281,N_12003);
nand U14958 (N_14958,N_12341,N_13055);
or U14959 (N_14959,N_12519,N_12462);
or U14960 (N_14960,N_12378,N_12197);
and U14961 (N_14961,N_13106,N_12289);
nor U14962 (N_14962,N_12715,N_12079);
xor U14963 (N_14963,N_12484,N_13188);
or U14964 (N_14964,N_12338,N_12035);
nor U14965 (N_14965,N_12310,N_12391);
or U14966 (N_14966,N_12426,N_12904);
nand U14967 (N_14967,N_12449,N_12626);
nand U14968 (N_14968,N_12006,N_13015);
and U14969 (N_14969,N_12912,N_12458);
xnor U14970 (N_14970,N_13127,N_12577);
or U14971 (N_14971,N_12015,N_13372);
or U14972 (N_14972,N_12567,N_12356);
or U14973 (N_14973,N_12955,N_12740);
nand U14974 (N_14974,N_12299,N_12913);
nand U14975 (N_14975,N_12063,N_12171);
and U14976 (N_14976,N_12080,N_13364);
nor U14977 (N_14977,N_12904,N_12871);
nor U14978 (N_14978,N_13007,N_13119);
nor U14979 (N_14979,N_12397,N_12286);
nand U14980 (N_14980,N_12088,N_13099);
nor U14981 (N_14981,N_12729,N_12539);
and U14982 (N_14982,N_13153,N_12425);
xor U14983 (N_14983,N_12563,N_12586);
nand U14984 (N_14984,N_12818,N_12870);
nor U14985 (N_14985,N_13454,N_12385);
nand U14986 (N_14986,N_12683,N_12619);
xor U14987 (N_14987,N_12597,N_12561);
nand U14988 (N_14988,N_13257,N_12253);
nor U14989 (N_14989,N_12137,N_13101);
nand U14990 (N_14990,N_12302,N_13103);
nand U14991 (N_14991,N_12780,N_13113);
nor U14992 (N_14992,N_13045,N_12224);
nor U14993 (N_14993,N_12078,N_12118);
nor U14994 (N_14994,N_12596,N_12176);
and U14995 (N_14995,N_13052,N_13110);
nor U14996 (N_14996,N_12380,N_13241);
nor U14997 (N_14997,N_12910,N_12168);
xnor U14998 (N_14998,N_12201,N_13145);
and U14999 (N_14999,N_13369,N_12028);
nand UO_0 (O_0,N_14956,N_13599);
nor UO_1 (O_1,N_13735,N_14161);
nand UO_2 (O_2,N_13892,N_14055);
nand UO_3 (O_3,N_14301,N_14336);
or UO_4 (O_4,N_14367,N_14768);
or UO_5 (O_5,N_13527,N_13752);
and UO_6 (O_6,N_14230,N_14364);
nand UO_7 (O_7,N_14431,N_14528);
nor UO_8 (O_8,N_14943,N_14154);
xor UO_9 (O_9,N_14619,N_14734);
nor UO_10 (O_10,N_14084,N_14683);
nand UO_11 (O_11,N_13611,N_13720);
nor UO_12 (O_12,N_14485,N_14441);
and UO_13 (O_13,N_14899,N_14333);
and UO_14 (O_14,N_14326,N_14624);
and UO_15 (O_15,N_14184,N_14162);
or UO_16 (O_16,N_14742,N_14814);
nor UO_17 (O_17,N_14639,N_13588);
and UO_18 (O_18,N_14136,N_14110);
or UO_19 (O_19,N_14483,N_14242);
xor UO_20 (O_20,N_14179,N_13780);
or UO_21 (O_21,N_14349,N_14335);
nor UO_22 (O_22,N_14965,N_14362);
nand UO_23 (O_23,N_14173,N_14781);
or UO_24 (O_24,N_14744,N_13900);
nand UO_25 (O_25,N_13691,N_13754);
or UO_26 (O_26,N_14312,N_13681);
and UO_27 (O_27,N_14967,N_14477);
or UO_28 (O_28,N_13570,N_14822);
nand UO_29 (O_29,N_13859,N_14203);
nor UO_30 (O_30,N_13705,N_14709);
or UO_31 (O_31,N_14157,N_14352);
or UO_32 (O_32,N_13765,N_14314);
nand UO_33 (O_33,N_14823,N_14450);
or UO_34 (O_34,N_14239,N_14511);
and UO_35 (O_35,N_13614,N_13888);
nand UO_36 (O_36,N_14950,N_14491);
xnor UO_37 (O_37,N_13983,N_14394);
nor UO_38 (O_38,N_13761,N_14425);
or UO_39 (O_39,N_14539,N_14011);
or UO_40 (O_40,N_14338,N_14987);
or UO_41 (O_41,N_13822,N_14885);
and UO_42 (O_42,N_14196,N_14262);
or UO_43 (O_43,N_13805,N_14166);
or UO_44 (O_44,N_13824,N_13972);
and UO_45 (O_45,N_14070,N_14473);
xor UO_46 (O_46,N_14276,N_14663);
and UO_47 (O_47,N_13626,N_14628);
nand UO_48 (O_48,N_14192,N_14104);
or UO_49 (O_49,N_14007,N_13856);
and UO_50 (O_50,N_14339,N_14711);
xnor UO_51 (O_51,N_14507,N_13955);
xor UO_52 (O_52,N_14325,N_14625);
or UO_53 (O_53,N_14068,N_13910);
or UO_54 (O_54,N_14804,N_14465);
nand UO_55 (O_55,N_13948,N_14834);
and UO_56 (O_56,N_14486,N_14611);
nand UO_57 (O_57,N_14605,N_14034);
or UO_58 (O_58,N_14089,N_14656);
nand UO_59 (O_59,N_13810,N_14828);
nand UO_60 (O_60,N_13627,N_13865);
and UO_61 (O_61,N_13645,N_14937);
nand UO_62 (O_62,N_14005,N_14248);
nand UO_63 (O_63,N_13815,N_14988);
and UO_64 (O_64,N_13637,N_14889);
xnor UO_65 (O_65,N_14621,N_14134);
or UO_66 (O_66,N_14847,N_14298);
nand UO_67 (O_67,N_14016,N_14788);
or UO_68 (O_68,N_13869,N_14740);
nand UO_69 (O_69,N_14942,N_13990);
nor UO_70 (O_70,N_14668,N_14064);
nand UO_71 (O_71,N_14460,N_13795);
nor UO_72 (O_72,N_13619,N_13947);
or UO_73 (O_73,N_14585,N_14653);
and UO_74 (O_74,N_14532,N_14258);
nand UO_75 (O_75,N_14470,N_14216);
nor UO_76 (O_76,N_14295,N_13731);
nand UO_77 (O_77,N_13759,N_13580);
xor UO_78 (O_78,N_14054,N_14633);
or UO_79 (O_79,N_14447,N_14687);
nor UO_80 (O_80,N_13982,N_14344);
nor UO_81 (O_81,N_13531,N_14384);
or UO_82 (O_82,N_14593,N_14553);
nand UO_83 (O_83,N_14733,N_14693);
xnor UO_84 (O_84,N_14446,N_14210);
xnor UO_85 (O_85,N_14418,N_14776);
nor UO_86 (O_86,N_13564,N_14752);
nand UO_87 (O_87,N_14741,N_13678);
and UO_88 (O_88,N_14391,N_13624);
or UO_89 (O_89,N_13794,N_14358);
nor UO_90 (O_90,N_14481,N_14850);
nand UO_91 (O_91,N_13646,N_13673);
or UO_92 (O_92,N_14671,N_14724);
nand UO_93 (O_93,N_14267,N_14255);
nand UO_94 (O_94,N_14222,N_13834);
nand UO_95 (O_95,N_14601,N_14971);
nor UO_96 (O_96,N_14717,N_14591);
nand UO_97 (O_97,N_13844,N_14327);
nor UO_98 (O_98,N_14449,N_14835);
nand UO_99 (O_99,N_13617,N_13850);
nor UO_100 (O_100,N_13860,N_14434);
xnor UO_101 (O_101,N_13830,N_14798);
xor UO_102 (O_102,N_14562,N_14320);
or UO_103 (O_103,N_13781,N_14445);
nand UO_104 (O_104,N_14690,N_14898);
nor UO_105 (O_105,N_14574,N_13886);
and UO_106 (O_106,N_14403,N_14001);
nor UO_107 (O_107,N_14359,N_14266);
nand UO_108 (O_108,N_14341,N_14091);
nand UO_109 (O_109,N_13751,N_13921);
nand UO_110 (O_110,N_14947,N_13538);
and UO_111 (O_111,N_14815,N_14506);
nand UO_112 (O_112,N_14840,N_14722);
nor UO_113 (O_113,N_14848,N_14827);
or UO_114 (O_114,N_14309,N_14864);
or UO_115 (O_115,N_13808,N_14737);
nor UO_116 (O_116,N_13700,N_14223);
or UO_117 (O_117,N_13616,N_14921);
or UO_118 (O_118,N_13989,N_13738);
and UO_119 (O_119,N_14159,N_13845);
and UO_120 (O_120,N_14175,N_14609);
or UO_121 (O_121,N_13543,N_14202);
nand UO_122 (O_122,N_14908,N_14660);
nor UO_123 (O_123,N_14669,N_14891);
and UO_124 (O_124,N_14705,N_14517);
nor UO_125 (O_125,N_14342,N_13529);
nor UO_126 (O_126,N_14880,N_14354);
nand UO_127 (O_127,N_14316,N_14172);
nand UO_128 (O_128,N_14227,N_13858);
nor UO_129 (O_129,N_14137,N_13978);
nor UO_130 (O_130,N_14514,N_14785);
xor UO_131 (O_131,N_13942,N_14347);
and UO_132 (O_132,N_14385,N_13940);
and UO_133 (O_133,N_14148,N_14424);
nand UO_134 (O_134,N_13715,N_14030);
and UO_135 (O_135,N_13618,N_14778);
nor UO_136 (O_136,N_13994,N_14045);
nor UO_137 (O_137,N_14564,N_14754);
nand UO_138 (O_138,N_14402,N_13908);
nand UO_139 (O_139,N_13604,N_13927);
and UO_140 (O_140,N_14544,N_13505);
nor UO_141 (O_141,N_14576,N_14407);
nor UO_142 (O_142,N_14953,N_14875);
xor UO_143 (O_143,N_14925,N_14659);
nand UO_144 (O_144,N_14286,N_13551);
and UO_145 (O_145,N_14990,N_14968);
nand UO_146 (O_146,N_13728,N_14206);
nand UO_147 (O_147,N_14524,N_14608);
and UO_148 (O_148,N_13647,N_14432);
nand UO_149 (O_149,N_14600,N_14551);
nor UO_150 (O_150,N_13634,N_14760);
and UO_151 (O_151,N_13710,N_14069);
or UO_152 (O_152,N_14060,N_14302);
nand UO_153 (O_153,N_14887,N_14368);
xnor UO_154 (O_154,N_13699,N_13514);
nand UO_155 (O_155,N_14962,N_14904);
xor UO_156 (O_156,N_13807,N_13911);
nand UO_157 (O_157,N_14076,N_14801);
and UO_158 (O_158,N_13937,N_14080);
nor UO_159 (O_159,N_13756,N_14836);
nand UO_160 (O_160,N_13961,N_14476);
and UO_161 (O_161,N_13509,N_13852);
xnor UO_162 (O_162,N_13562,N_13660);
and UO_163 (O_163,N_13851,N_13920);
nand UO_164 (O_164,N_14926,N_14578);
and UO_165 (O_165,N_14749,N_14819);
nor UO_166 (O_166,N_14322,N_13550);
nand UO_167 (O_167,N_14996,N_14145);
xor UO_168 (O_168,N_14509,N_14504);
or UO_169 (O_169,N_14494,N_14598);
and UO_170 (O_170,N_13584,N_14582);
xnor UO_171 (O_171,N_14348,N_14259);
nand UO_172 (O_172,N_14405,N_14974);
xor UO_173 (O_173,N_13596,N_14146);
and UO_174 (O_174,N_14411,N_13512);
and UO_175 (O_175,N_13686,N_14000);
nand UO_176 (O_176,N_14584,N_14490);
nor UO_177 (O_177,N_14195,N_14073);
nand UO_178 (O_178,N_13557,N_14098);
and UO_179 (O_179,N_13758,N_14099);
nor UO_180 (O_180,N_14508,N_13750);
nand UO_181 (O_181,N_14153,N_13674);
nand UO_182 (O_182,N_13726,N_14896);
and UO_183 (O_183,N_14294,N_13517);
or UO_184 (O_184,N_13966,N_13802);
nor UO_185 (O_185,N_14397,N_13714);
nor UO_186 (O_186,N_14905,N_14868);
nor UO_187 (O_187,N_14805,N_14113);
xnor UO_188 (O_188,N_14300,N_14428);
or UO_189 (O_189,N_14330,N_13537);
nor UO_190 (O_190,N_13820,N_14277);
nand UO_191 (O_191,N_14332,N_13784);
or UO_192 (O_192,N_13901,N_14408);
nand UO_193 (O_193,N_13960,N_13721);
xnor UO_194 (O_194,N_14542,N_14592);
or UO_195 (O_195,N_14141,N_14061);
nand UO_196 (O_196,N_13930,N_14612);
nand UO_197 (O_197,N_14058,N_13546);
nor UO_198 (O_198,N_14699,N_14221);
nand UO_199 (O_199,N_14256,N_14127);
or UO_200 (O_200,N_13826,N_14537);
nand UO_201 (O_201,N_13526,N_14863);
and UO_202 (O_202,N_14251,N_13657);
nand UO_203 (O_203,N_13649,N_13642);
nand UO_204 (O_204,N_14328,N_14573);
or UO_205 (O_205,N_14096,N_14254);
and UO_206 (O_206,N_13722,N_14211);
or UO_207 (O_207,N_14019,N_14548);
nand UO_208 (O_208,N_14409,N_14991);
or UO_209 (O_209,N_14090,N_14082);
and UO_210 (O_210,N_14932,N_13747);
nor UO_211 (O_211,N_14351,N_14552);
nor UO_212 (O_212,N_13702,N_13522);
and UO_213 (O_213,N_14272,N_14201);
xnor UO_214 (O_214,N_14353,N_13589);
or UO_215 (O_215,N_13572,N_14097);
xnor UO_216 (O_216,N_14541,N_14510);
nand UO_217 (O_217,N_13866,N_14452);
or UO_218 (O_218,N_14273,N_13719);
or UO_219 (O_219,N_13501,N_13958);
or UO_220 (O_220,N_14743,N_13541);
and UO_221 (O_221,N_13988,N_13682);
nor UO_222 (O_222,N_14969,N_14185);
nand UO_223 (O_223,N_14042,N_13676);
nand UO_224 (O_224,N_14940,N_14252);
nand UO_225 (O_225,N_14916,N_14261);
nor UO_226 (O_226,N_13707,N_14149);
or UO_227 (O_227,N_14535,N_14174);
nand UO_228 (O_228,N_14720,N_14121);
and UO_229 (O_229,N_14519,N_14998);
and UO_230 (O_230,N_13629,N_14117);
nor UO_231 (O_231,N_13934,N_14412);
nand UO_232 (O_232,N_14033,N_13772);
or UO_233 (O_233,N_13950,N_13867);
nor UO_234 (O_234,N_14870,N_14571);
or UO_235 (O_235,N_13500,N_14038);
nor UO_236 (O_236,N_14500,N_14503);
or UO_237 (O_237,N_14062,N_13662);
nor UO_238 (O_238,N_14648,N_14867);
and UO_239 (O_239,N_13929,N_13668);
nor UO_240 (O_240,N_14824,N_14063);
xor UO_241 (O_241,N_14757,N_14997);
xor UO_242 (O_242,N_13612,N_13928);
or UO_243 (O_243,N_14212,N_14973);
nor UO_244 (O_244,N_13953,N_14696);
or UO_245 (O_245,N_13832,N_14310);
nand UO_246 (O_246,N_14949,N_13553);
and UO_247 (O_247,N_14453,N_14673);
and UO_248 (O_248,N_13503,N_14730);
or UO_249 (O_249,N_14726,N_14247);
nand UO_250 (O_250,N_14704,N_14946);
nand UO_251 (O_251,N_14417,N_14550);
nand UO_252 (O_252,N_13895,N_14182);
nand UO_253 (O_253,N_14959,N_14809);
nand UO_254 (O_254,N_14004,N_14280);
nand UO_255 (O_255,N_13661,N_14793);
xnor UO_256 (O_256,N_13963,N_14786);
or UO_257 (O_257,N_14093,N_14324);
or UO_258 (O_258,N_14290,N_14041);
nand UO_259 (O_259,N_14284,N_13643);
or UO_260 (O_260,N_14178,N_14457);
nor UO_261 (O_261,N_14627,N_13936);
or UO_262 (O_262,N_13943,N_14787);
nand UO_263 (O_263,N_14023,N_14115);
and UO_264 (O_264,N_14913,N_13783);
and UO_265 (O_265,N_14305,N_14479);
or UO_266 (O_266,N_14365,N_14855);
and UO_267 (O_267,N_14976,N_13849);
xor UO_268 (O_268,N_14219,N_14977);
nor UO_269 (O_269,N_14106,N_14533);
and UO_270 (O_270,N_14369,N_13919);
nor UO_271 (O_271,N_14516,N_14686);
nor UO_272 (O_272,N_14520,N_14777);
nor UO_273 (O_273,N_14646,N_14296);
nand UO_274 (O_274,N_14264,N_13945);
and UO_275 (O_275,N_13764,N_14455);
or UO_276 (O_276,N_14225,N_14945);
or UO_277 (O_277,N_13569,N_13737);
or UO_278 (O_278,N_13524,N_13644);
nor UO_279 (O_279,N_14811,N_14231);
and UO_280 (O_280,N_14773,N_13595);
nor UO_281 (O_281,N_14388,N_13633);
and UO_282 (O_282,N_14919,N_14638);
nand UO_283 (O_283,N_13991,N_14961);
nand UO_284 (O_284,N_14651,N_14872);
and UO_285 (O_285,N_14766,N_13977);
nor UO_286 (O_286,N_13975,N_13535);
nor UO_287 (O_287,N_14466,N_14924);
or UO_288 (O_288,N_14051,N_13656);
and UO_289 (O_289,N_13732,N_14176);
or UO_290 (O_290,N_14829,N_13609);
nand UO_291 (O_291,N_14390,N_14554);
xor UO_292 (O_292,N_14235,N_14072);
nor UO_293 (O_293,N_14436,N_14345);
or UO_294 (O_294,N_13981,N_13566);
xor UO_295 (O_295,N_14472,N_14763);
or UO_296 (O_296,N_14094,N_14401);
xor UO_297 (O_297,N_14637,N_14665);
and UO_298 (O_298,N_13749,N_13918);
nand UO_299 (O_299,N_14135,N_13677);
nor UO_300 (O_300,N_14088,N_14065);
nor UO_301 (O_301,N_13855,N_13944);
nand UO_302 (O_302,N_13812,N_14423);
nand UO_303 (O_303,N_13818,N_13969);
nor UO_304 (O_304,N_13763,N_14549);
nand UO_305 (O_305,N_13903,N_14536);
nand UO_306 (O_306,N_14204,N_14933);
or UO_307 (O_307,N_14451,N_13560);
nand UO_308 (O_308,N_14794,N_14732);
or UO_309 (O_309,N_14092,N_14167);
or UO_310 (O_310,N_14382,N_14198);
xor UO_311 (O_311,N_13979,N_13799);
or UO_312 (O_312,N_14691,N_14140);
nand UO_313 (O_313,N_14229,N_13797);
nor UO_314 (O_314,N_14642,N_14652);
nor UO_315 (O_315,N_14771,N_13974);
nand UO_316 (O_316,N_13711,N_14907);
and UO_317 (O_317,N_14556,N_13742);
nor UO_318 (O_318,N_14900,N_13829);
nor UO_319 (O_319,N_14143,N_13873);
or UO_320 (O_320,N_14496,N_14666);
nor UO_321 (O_321,N_13768,N_14200);
and UO_322 (O_322,N_14645,N_13891);
nand UO_323 (O_323,N_14077,N_14501);
or UO_324 (O_324,N_14939,N_13771);
nand UO_325 (O_325,N_14293,N_13793);
nor UO_326 (O_326,N_13938,N_14265);
or UO_327 (O_327,N_14240,N_14983);
and UO_328 (O_328,N_13843,N_13636);
and UO_329 (O_329,N_14782,N_13857);
or UO_330 (O_330,N_14631,N_14802);
xnor UO_331 (O_331,N_14437,N_13603);
nand UO_332 (O_332,N_14049,N_14614);
nor UO_333 (O_333,N_14795,N_14395);
xnor UO_334 (O_334,N_14253,N_13713);
nand UO_335 (O_335,N_14169,N_14980);
and UO_336 (O_336,N_13987,N_14731);
nand UO_337 (O_337,N_13907,N_13884);
or UO_338 (O_338,N_14199,N_14789);
or UO_339 (O_339,N_14715,N_14587);
nor UO_340 (O_340,N_14886,N_14912);
nand UO_341 (O_341,N_14037,N_14989);
and UO_342 (O_342,N_14181,N_14685);
and UO_343 (O_343,N_13821,N_14241);
nor UO_344 (O_344,N_13878,N_13916);
or UO_345 (O_345,N_13727,N_14321);
or UO_346 (O_346,N_13653,N_14853);
nor UO_347 (O_347,N_14689,N_13641);
xnor UO_348 (O_348,N_13698,N_14006);
nor UO_349 (O_349,N_14406,N_14799);
or UO_350 (O_350,N_14881,N_14878);
or UO_351 (O_351,N_14040,N_14599);
or UO_352 (O_352,N_14677,N_13534);
nor UO_353 (O_353,N_14420,N_14812);
nand UO_354 (O_354,N_14676,N_13868);
nand UO_355 (O_355,N_14337,N_14684);
and UO_356 (O_356,N_13757,N_13862);
xor UO_357 (O_357,N_13804,N_13610);
or UO_358 (O_358,N_13545,N_14170);
nand UO_359 (O_359,N_14057,N_14502);
xnor UO_360 (O_360,N_13544,N_14075);
and UO_361 (O_361,N_14606,N_14079);
or UO_362 (O_362,N_14360,N_14462);
or UO_363 (O_363,N_13659,N_13600);
xnor UO_364 (O_364,N_14540,N_13515);
or UO_365 (O_365,N_14066,N_14243);
nand UO_366 (O_366,N_14171,N_13760);
and UO_367 (O_367,N_13774,N_14414);
or UO_368 (O_368,N_13578,N_14716);
and UO_369 (O_369,N_14107,N_13847);
or UO_370 (O_370,N_14101,N_14753);
and UO_371 (O_371,N_13792,N_14616);
or UO_372 (O_372,N_13741,N_13879);
or UO_373 (O_373,N_13558,N_13898);
xnor UO_374 (O_374,N_14165,N_13554);
or UO_375 (O_375,N_14439,N_14910);
and UO_376 (O_376,N_14116,N_13816);
nor UO_377 (O_377,N_13716,N_13555);
or UO_378 (O_378,N_14422,N_14630);
nand UO_379 (O_379,N_14765,N_13739);
or UO_380 (O_380,N_13587,N_14702);
nor UO_381 (O_381,N_13952,N_14882);
xor UO_382 (O_382,N_14438,N_14100);
and UO_383 (O_383,N_14263,N_14529);
or UO_384 (O_384,N_13906,N_14972);
or UO_385 (O_385,N_13912,N_13909);
or UO_386 (O_386,N_14194,N_14433);
nor UO_387 (O_387,N_14215,N_13880);
xnor UO_388 (O_388,N_14489,N_14993);
nor UO_389 (O_389,N_14022,N_14806);
and UO_390 (O_390,N_13571,N_13788);
or UO_391 (O_391,N_14112,N_13746);
nand UO_392 (O_392,N_14634,N_13870);
or UO_393 (O_393,N_14700,N_13563);
or UO_394 (O_394,N_14197,N_13791);
xor UO_395 (O_395,N_14257,N_14934);
or UO_396 (O_396,N_14003,N_14487);
xor UO_397 (O_397,N_14865,N_14085);
nand UO_398 (O_398,N_13725,N_13670);
or UO_399 (O_399,N_14825,N_14071);
nor UO_400 (O_400,N_14727,N_14721);
nand UO_401 (O_401,N_13941,N_14189);
nor UO_402 (O_402,N_14586,N_13933);
or UO_403 (O_403,N_14285,N_14467);
xnor UO_404 (O_404,N_14657,N_13671);
nor UO_405 (O_405,N_14398,N_14128);
or UO_406 (O_406,N_14393,N_13896);
nor UO_407 (O_407,N_14565,N_14780);
nand UO_408 (O_408,N_13782,N_13736);
or UO_409 (O_409,N_14187,N_13689);
or UO_410 (O_410,N_13533,N_13775);
and UO_411 (O_411,N_13559,N_14783);
or UO_412 (O_412,N_14122,N_14762);
nand UO_413 (O_413,N_13598,N_13897);
or UO_414 (O_414,N_14315,N_13931);
nand UO_415 (O_415,N_14307,N_13523);
and UO_416 (O_416,N_14603,N_14118);
nor UO_417 (O_417,N_14563,N_14797);
or UO_418 (O_418,N_13790,N_14756);
nor UO_419 (O_419,N_13814,N_14607);
nor UO_420 (O_420,N_14083,N_14670);
nand UO_421 (O_421,N_13590,N_14658);
and UO_422 (O_422,N_14644,N_14888);
nor UO_423 (O_423,N_13513,N_14764);
nand UO_424 (O_424,N_14289,N_14713);
nor UO_425 (O_425,N_13828,N_13872);
nand UO_426 (O_426,N_14426,N_14897);
nand UO_427 (O_427,N_14817,N_14569);
nor UO_428 (O_428,N_13984,N_14957);
and UO_429 (O_429,N_14861,N_14796);
nand UO_430 (O_430,N_13980,N_14994);
nor UO_431 (O_431,N_14738,N_13753);
xnor UO_432 (O_432,N_13575,N_14530);
or UO_433 (O_433,N_14010,N_14859);
nor UO_434 (O_434,N_14791,N_14664);
or UO_435 (O_435,N_14274,N_14581);
nor UO_436 (O_436,N_14031,N_13766);
nor UO_437 (O_437,N_14761,N_14807);
and UO_438 (O_438,N_14936,N_14821);
nand UO_439 (O_439,N_14456,N_13997);
and UO_440 (O_440,N_14350,N_14613);
nand UO_441 (O_441,N_14133,N_13740);
and UO_442 (O_442,N_14356,N_14012);
xor UO_443 (O_443,N_14960,N_13785);
and UO_444 (O_444,N_13854,N_14234);
or UO_445 (O_445,N_13968,N_14813);
xnor UO_446 (O_446,N_14719,N_13992);
or UO_447 (O_447,N_14736,N_13679);
or UO_448 (O_448,N_14186,N_14238);
or UO_449 (O_449,N_13730,N_14674);
nor UO_450 (O_450,N_14020,N_14832);
xor UO_451 (O_451,N_14468,N_13876);
nor UO_452 (O_452,N_13519,N_13962);
nand UO_453 (O_453,N_13506,N_14319);
nand UO_454 (O_454,N_13620,N_14379);
and UO_455 (O_455,N_14226,N_14308);
nand UO_456 (O_456,N_14377,N_14361);
or UO_457 (O_457,N_14545,N_13813);
nand UO_458 (O_458,N_14838,N_14803);
nand UO_459 (O_459,N_14546,N_14014);
nand UO_460 (O_460,N_14728,N_14981);
or UO_461 (O_461,N_13631,N_14978);
nor UO_462 (O_462,N_13532,N_13885);
and UO_463 (O_463,N_14318,N_14281);
or UO_464 (O_464,N_14497,N_14790);
nor UO_465 (O_465,N_13536,N_14044);
and UO_466 (O_466,N_14109,N_13675);
nand UO_467 (O_467,N_14979,N_14930);
nor UO_468 (O_468,N_14518,N_13508);
and UO_469 (O_469,N_14846,N_14087);
or UO_470 (O_470,N_13615,N_13712);
or UO_471 (O_471,N_14124,N_13632);
nand UO_472 (O_472,N_14028,N_14842);
nand UO_473 (O_473,N_14002,N_14622);
nor UO_474 (O_474,N_13809,N_14357);
nor UO_475 (O_475,N_13796,N_14279);
or UO_476 (O_476,N_13577,N_13913);
or UO_477 (O_477,N_13755,N_14521);
nand UO_478 (O_478,N_13680,N_14052);
and UO_479 (O_479,N_14735,N_14929);
nand UO_480 (O_480,N_13623,N_14583);
or UO_481 (O_481,N_14680,N_13925);
or UO_482 (O_482,N_14081,N_14493);
xnor UO_483 (O_483,N_13574,N_14056);
nand UO_484 (O_484,N_14567,N_14268);
xor UO_485 (O_485,N_13717,N_13801);
nor UO_486 (O_486,N_14214,N_14986);
nand UO_487 (O_487,N_14059,N_14236);
and UO_488 (O_488,N_14024,N_13597);
and UO_489 (O_489,N_14323,N_14751);
or UO_490 (O_490,N_14590,N_13540);
or UO_491 (O_491,N_14523,N_13581);
nand UO_492 (O_492,N_14681,N_14952);
nand UO_493 (O_493,N_14635,N_13723);
nand UO_494 (O_494,N_14849,N_13967);
nand UO_495 (O_495,N_13579,N_14386);
nand UO_496 (O_496,N_13899,N_13767);
nor UO_497 (O_497,N_13548,N_13654);
nor UO_498 (O_498,N_14816,N_14901);
or UO_499 (O_499,N_14480,N_13696);
nand UO_500 (O_500,N_14538,N_14557);
and UO_501 (O_501,N_13743,N_13542);
nand UO_502 (O_502,N_14769,N_14931);
nor UO_503 (O_503,N_14958,N_13835);
nor UO_504 (O_504,N_13666,N_14770);
and UO_505 (O_505,N_13504,N_14095);
nor UO_506 (O_506,N_14954,N_14404);
nand UO_507 (O_507,N_14871,N_14566);
and UO_508 (O_508,N_14706,N_14224);
and UO_509 (O_509,N_14917,N_14561);
and UO_510 (O_510,N_14833,N_14050);
and UO_511 (O_511,N_14410,N_13964);
or UO_512 (O_512,N_14443,N_14679);
nor UO_513 (O_513,N_13704,N_14906);
xnor UO_514 (O_514,N_13510,N_14938);
nor UO_515 (O_515,N_14602,N_14775);
xor UO_516 (O_516,N_13965,N_14559);
and UO_517 (O_517,N_14013,N_13956);
nor UO_518 (O_518,N_13594,N_13745);
and UO_519 (O_519,N_13621,N_14800);
and UO_520 (O_520,N_14808,N_14421);
nor UO_521 (O_521,N_14026,N_14589);
xnor UO_522 (O_522,N_13871,N_13669);
nand UO_523 (O_523,N_14640,N_14304);
xor UO_524 (O_524,N_14374,N_14205);
and UO_525 (O_525,N_14278,N_13697);
nor UO_526 (O_526,N_13665,N_14555);
xnor UO_527 (O_527,N_13874,N_13638);
or UO_528 (O_528,N_14649,N_14662);
nand UO_529 (O_529,N_13923,N_14488);
xor UO_530 (O_530,N_13786,N_14188);
nand UO_531 (O_531,N_13561,N_14505);
and UO_532 (O_532,N_14866,N_14909);
and UO_533 (O_533,N_13762,N_14464);
nand UO_534 (O_534,N_14046,N_13976);
nor UO_535 (O_535,N_14697,N_13530);
xor UO_536 (O_536,N_14841,N_14282);
nor UO_537 (O_537,N_13839,N_13825);
nand UO_538 (O_538,N_14911,N_14883);
xor UO_539 (O_539,N_14854,N_13939);
nand UO_540 (O_540,N_14246,N_14130);
or UO_541 (O_541,N_13652,N_13708);
or UO_542 (O_542,N_13724,N_14220);
nand UO_543 (O_543,N_14249,N_13658);
nand UO_544 (O_544,N_13568,N_13733);
or UO_545 (O_545,N_14661,N_14484);
and UO_546 (O_546,N_14371,N_13650);
xnor UO_547 (O_547,N_14610,N_14725);
or UO_548 (O_548,N_13635,N_13863);
and UO_549 (O_549,N_14471,N_14672);
nor UO_550 (O_550,N_14454,N_14183);
nor UO_551 (O_551,N_14918,N_14655);
or UO_552 (O_552,N_14444,N_14707);
nor UO_553 (O_553,N_14982,N_13817);
nand UO_554 (O_554,N_14269,N_14710);
and UO_555 (O_555,N_14400,N_13890);
or UO_556 (O_556,N_14914,N_14475);
and UO_557 (O_557,N_14383,N_13718);
and UO_558 (O_558,N_13882,N_13777);
and UO_559 (O_559,N_14869,N_14543);
or UO_560 (O_560,N_13573,N_13881);
nor UO_561 (O_561,N_14568,N_14288);
xor UO_562 (O_562,N_14618,N_14144);
or UO_563 (O_563,N_13688,N_13511);
or UO_564 (O_564,N_14902,N_14739);
and UO_565 (O_565,N_13819,N_13685);
and UO_566 (O_566,N_13773,N_14570);
or UO_567 (O_567,N_13946,N_14851);
or UO_568 (O_568,N_14442,N_14572);
or UO_569 (O_569,N_14892,N_13779);
nor UO_570 (O_570,N_14857,N_13889);
xnor UO_571 (O_571,N_14125,N_14876);
and UO_572 (O_572,N_14132,N_14879);
and UO_573 (O_573,N_13769,N_14531);
xor UO_574 (O_574,N_14675,N_14074);
and UO_575 (O_575,N_13803,N_13576);
or UO_576 (O_576,N_14858,N_14250);
or UO_577 (O_577,N_14928,N_14966);
nor UO_578 (O_578,N_14209,N_14862);
nand UO_579 (O_579,N_14306,N_14440);
and UO_580 (O_580,N_14604,N_14376);
and UO_581 (O_581,N_14894,N_14355);
nor UO_582 (O_582,N_13973,N_13831);
nor UO_583 (O_583,N_14852,N_14158);
or UO_584 (O_584,N_14667,N_14283);
and UO_585 (O_585,N_14126,N_13602);
nand UO_586 (O_586,N_14047,N_13954);
nor UO_587 (O_587,N_13827,N_13525);
nor UO_588 (O_588,N_14513,N_13986);
and UO_589 (O_589,N_14032,N_14208);
and UO_590 (O_590,N_13593,N_14698);
nor UO_591 (O_591,N_14856,N_13864);
nand UO_592 (O_592,N_13917,N_13687);
and UO_593 (O_593,N_14948,N_13613);
nor UO_594 (O_594,N_13837,N_14837);
nand UO_595 (O_595,N_13922,N_14463);
nand UO_596 (O_596,N_14629,N_13556);
and UO_597 (O_597,N_14594,N_13672);
nand UO_598 (O_598,N_14723,N_13663);
nor UO_599 (O_599,N_14129,N_13823);
nand UO_600 (O_600,N_14228,N_14193);
nand UO_601 (O_601,N_14845,N_14703);
nor UO_602 (O_602,N_13787,N_14147);
and UO_603 (O_603,N_14180,N_13914);
or UO_604 (O_604,N_14123,N_14746);
nand UO_605 (O_605,N_14008,N_13776);
nor UO_606 (O_606,N_14313,N_13694);
nor UO_607 (O_607,N_14317,N_13630);
and UO_608 (O_608,N_14035,N_14413);
and UO_609 (O_609,N_13552,N_14922);
or UO_610 (O_610,N_14429,N_14650);
and UO_611 (O_611,N_14381,N_14784);
and UO_612 (O_612,N_14389,N_14139);
nor UO_613 (O_613,N_14415,N_13996);
nand UO_614 (O_614,N_13693,N_13887);
nor UO_615 (O_615,N_14340,N_13778);
nor UO_616 (O_616,N_13601,N_13846);
nor UO_617 (O_617,N_14498,N_13841);
or UO_618 (O_618,N_14903,N_13998);
and UO_619 (O_619,N_14748,N_13518);
nand UO_620 (O_620,N_14527,N_14142);
xor UO_621 (O_621,N_13875,N_14039);
or UO_622 (O_622,N_14620,N_13606);
nor UO_623 (O_623,N_14370,N_14131);
nand UO_624 (O_624,N_14964,N_14373);
nand UO_625 (O_625,N_14963,N_14469);
nor UO_626 (O_626,N_14820,N_14792);
or UO_627 (O_627,N_14164,N_14053);
or UO_628 (O_628,N_14779,N_13521);
xor UO_629 (O_629,N_14036,N_13894);
nor UO_630 (O_630,N_14708,N_13628);
and UO_631 (O_631,N_14334,N_14985);
and UO_632 (O_632,N_14311,N_14114);
and UO_633 (O_633,N_13648,N_14927);
nor UO_634 (O_634,N_13567,N_14515);
and UO_635 (O_635,N_14168,N_14156);
nand UO_636 (O_636,N_14435,N_13585);
nand UO_637 (O_637,N_14297,N_14120);
and UO_638 (O_638,N_13949,N_14392);
nor UO_639 (O_639,N_13692,N_14287);
xor UO_640 (O_640,N_14009,N_14207);
nand UO_641 (O_641,N_14772,N_14459);
nand UO_642 (O_642,N_14955,N_14458);
or UO_643 (O_643,N_13971,N_14138);
nor UO_644 (O_644,N_13592,N_14048);
nand UO_645 (O_645,N_14580,N_14579);
nand UO_646 (O_646,N_14999,N_14363);
and UO_647 (O_647,N_14152,N_14018);
and UO_648 (O_648,N_14299,N_13848);
nor UO_649 (O_649,N_14213,N_14067);
and UO_650 (O_650,N_14893,N_14758);
or UO_651 (O_651,N_13935,N_13995);
nor UO_652 (O_652,N_13549,N_13547);
xor UO_653 (O_653,N_14366,N_14818);
nor UO_654 (O_654,N_14682,N_13516);
nand UO_655 (O_655,N_14831,N_14755);
nand UO_656 (O_656,N_13605,N_13591);
or UO_657 (O_657,N_14163,N_14292);
nand UO_658 (O_658,N_13520,N_13683);
and UO_659 (O_659,N_14111,N_13893);
nor UO_660 (O_660,N_13706,N_14935);
nor UO_661 (O_661,N_14615,N_14522);
nand UO_662 (O_662,N_14915,N_13770);
nand UO_663 (O_663,N_14596,N_13951);
or UO_664 (O_664,N_14478,N_14078);
nor UO_665 (O_665,N_13798,N_14021);
and UO_666 (O_666,N_14448,N_14839);
or UO_667 (O_667,N_13842,N_14495);
or UO_668 (O_668,N_13748,N_14025);
and UO_669 (O_669,N_13502,N_13902);
nor UO_670 (O_670,N_13924,N_13664);
and UO_671 (O_671,N_14729,N_14043);
nand UO_672 (O_672,N_14396,N_14558);
nand UO_673 (O_673,N_13701,N_14105);
nor UO_674 (O_674,N_14547,N_13904);
and UO_675 (O_675,N_14944,N_14419);
nand UO_676 (O_676,N_14995,N_13565);
xor UO_677 (O_677,N_13690,N_14029);
or UO_678 (O_678,N_14430,N_14218);
and UO_679 (O_679,N_14577,N_14623);
and UO_680 (O_680,N_14492,N_14108);
or UO_681 (O_681,N_13999,N_13583);
or UO_682 (O_682,N_14160,N_13970);
xor UO_683 (O_683,N_14232,N_14474);
and UO_684 (O_684,N_14920,N_14923);
nor UO_685 (O_685,N_13622,N_14970);
nand UO_686 (O_686,N_14271,N_14830);
nand UO_687 (O_687,N_13607,N_14427);
nor UO_688 (O_688,N_14810,N_14086);
nor UO_689 (O_689,N_14695,N_13667);
xnor UO_690 (O_690,N_14873,N_14826);
nor UO_691 (O_691,N_13625,N_14688);
nand UO_692 (O_692,N_13840,N_14237);
nor UO_693 (O_693,N_14890,N_14595);
and UO_694 (O_694,N_14270,N_14015);
and UO_695 (O_695,N_14647,N_14102);
nand UO_696 (O_696,N_14244,N_14027);
and UO_697 (O_697,N_14745,N_14877);
nand UO_698 (O_698,N_14641,N_13582);
or UO_699 (O_699,N_14372,N_14375);
nor UO_700 (O_700,N_14701,N_14233);
nor UO_701 (O_701,N_13684,N_14692);
nand UO_702 (O_702,N_14759,N_14346);
and UO_703 (O_703,N_14941,N_14245);
and UO_704 (O_704,N_14378,N_13861);
nand UO_705 (O_705,N_14260,N_14190);
or UO_706 (O_706,N_14119,N_14387);
and UO_707 (O_707,N_14482,N_14844);
and UO_708 (O_708,N_14884,N_13836);
and UO_709 (O_709,N_14975,N_14747);
nand UO_710 (O_710,N_14416,N_14399);
nand UO_711 (O_711,N_14588,N_13744);
nor UO_712 (O_712,N_14774,N_14560);
or UO_713 (O_713,N_13703,N_13507);
and UO_714 (O_714,N_13811,N_13957);
nand UO_715 (O_715,N_14654,N_13608);
or UO_716 (O_716,N_14331,N_13993);
and UO_717 (O_717,N_14860,N_14678);
nor UO_718 (O_718,N_14767,N_13695);
nor UO_719 (O_719,N_13926,N_13915);
nor UO_720 (O_720,N_14843,N_13959);
and UO_721 (O_721,N_14177,N_14329);
nor UO_722 (O_722,N_13985,N_14617);
or UO_723 (O_723,N_14718,N_14499);
nand UO_724 (O_724,N_14017,N_14636);
or UO_725 (O_725,N_14712,N_13806);
nor UO_726 (O_726,N_14526,N_13651);
and UO_727 (O_727,N_13789,N_14714);
and UO_728 (O_728,N_14951,N_14191);
and UO_729 (O_729,N_14343,N_14626);
nor UO_730 (O_730,N_14694,N_13655);
nand UO_731 (O_731,N_14461,N_14103);
nor UO_732 (O_732,N_14575,N_13838);
and UO_733 (O_733,N_13883,N_14525);
or UO_734 (O_734,N_13734,N_14512);
nor UO_735 (O_735,N_14151,N_14534);
nor UO_736 (O_736,N_13853,N_14992);
or UO_737 (O_737,N_13800,N_14984);
nor UO_738 (O_738,N_13528,N_14275);
nand UO_739 (O_739,N_14750,N_13539);
and UO_740 (O_740,N_14643,N_14632);
nor UO_741 (O_741,N_14874,N_14597);
or UO_742 (O_742,N_13640,N_14303);
xnor UO_743 (O_743,N_14155,N_13639);
nand UO_744 (O_744,N_14150,N_13833);
nor UO_745 (O_745,N_13932,N_13729);
and UO_746 (O_746,N_13586,N_14217);
nand UO_747 (O_747,N_13877,N_14895);
nor UO_748 (O_748,N_13905,N_14291);
nand UO_749 (O_749,N_13709,N_14380);
nor UO_750 (O_750,N_13712,N_14017);
nand UO_751 (O_751,N_14648,N_14244);
and UO_752 (O_752,N_13835,N_14022);
or UO_753 (O_753,N_14935,N_14053);
nor UO_754 (O_754,N_14023,N_14635);
or UO_755 (O_755,N_14082,N_14302);
nor UO_756 (O_756,N_13955,N_13987);
or UO_757 (O_757,N_14495,N_14293);
and UO_758 (O_758,N_14269,N_14247);
xor UO_759 (O_759,N_14911,N_14447);
or UO_760 (O_760,N_13670,N_14682);
nor UO_761 (O_761,N_13844,N_14955);
or UO_762 (O_762,N_13509,N_14507);
nand UO_763 (O_763,N_14721,N_14916);
and UO_764 (O_764,N_14760,N_14164);
xnor UO_765 (O_765,N_14179,N_14976);
or UO_766 (O_766,N_14523,N_14046);
nand UO_767 (O_767,N_14652,N_14959);
or UO_768 (O_768,N_13976,N_14362);
nand UO_769 (O_769,N_13542,N_14142);
and UO_770 (O_770,N_13669,N_14786);
xnor UO_771 (O_771,N_14496,N_14469);
or UO_772 (O_772,N_14161,N_14961);
xnor UO_773 (O_773,N_13526,N_14746);
nor UO_774 (O_774,N_14814,N_14869);
xor UO_775 (O_775,N_14609,N_14714);
nor UO_776 (O_776,N_14961,N_13773);
and UO_777 (O_777,N_14792,N_13858);
or UO_778 (O_778,N_14653,N_14821);
nand UO_779 (O_779,N_14012,N_13526);
nor UO_780 (O_780,N_13892,N_14910);
and UO_781 (O_781,N_14448,N_14059);
and UO_782 (O_782,N_13582,N_13972);
nand UO_783 (O_783,N_13579,N_13593);
nand UO_784 (O_784,N_14969,N_14326);
and UO_785 (O_785,N_13853,N_14055);
and UO_786 (O_786,N_14278,N_14371);
or UO_787 (O_787,N_13722,N_13920);
and UO_788 (O_788,N_14571,N_13603);
and UO_789 (O_789,N_14080,N_13741);
or UO_790 (O_790,N_14890,N_14230);
or UO_791 (O_791,N_14048,N_14138);
xnor UO_792 (O_792,N_13601,N_14475);
or UO_793 (O_793,N_13549,N_14492);
nand UO_794 (O_794,N_13745,N_14993);
nor UO_795 (O_795,N_13748,N_14973);
or UO_796 (O_796,N_14158,N_14487);
and UO_797 (O_797,N_14706,N_13604);
nand UO_798 (O_798,N_14673,N_13771);
nand UO_799 (O_799,N_13687,N_14391);
or UO_800 (O_800,N_14754,N_13748);
nor UO_801 (O_801,N_14820,N_14723);
or UO_802 (O_802,N_13779,N_14909);
or UO_803 (O_803,N_13959,N_13788);
or UO_804 (O_804,N_13504,N_14644);
or UO_805 (O_805,N_13854,N_14959);
nand UO_806 (O_806,N_14153,N_14242);
nor UO_807 (O_807,N_14831,N_13807);
and UO_808 (O_808,N_14333,N_13929);
or UO_809 (O_809,N_14634,N_14564);
nor UO_810 (O_810,N_14150,N_14975);
or UO_811 (O_811,N_13996,N_14569);
or UO_812 (O_812,N_13948,N_13842);
or UO_813 (O_813,N_13824,N_13673);
or UO_814 (O_814,N_13819,N_14313);
nand UO_815 (O_815,N_14196,N_14198);
nand UO_816 (O_816,N_13911,N_14189);
or UO_817 (O_817,N_14591,N_13564);
nor UO_818 (O_818,N_14916,N_14847);
or UO_819 (O_819,N_14439,N_13565);
and UO_820 (O_820,N_14057,N_13653);
or UO_821 (O_821,N_14635,N_13695);
nor UO_822 (O_822,N_14546,N_13708);
or UO_823 (O_823,N_14879,N_13683);
nand UO_824 (O_824,N_14061,N_13867);
nor UO_825 (O_825,N_14922,N_13856);
and UO_826 (O_826,N_14254,N_14897);
nand UO_827 (O_827,N_14427,N_14033);
and UO_828 (O_828,N_14804,N_14064);
or UO_829 (O_829,N_14230,N_13851);
nand UO_830 (O_830,N_14672,N_14131);
nand UO_831 (O_831,N_14179,N_14616);
and UO_832 (O_832,N_14431,N_14506);
nand UO_833 (O_833,N_13555,N_14447);
or UO_834 (O_834,N_13550,N_13940);
nor UO_835 (O_835,N_14837,N_14408);
nor UO_836 (O_836,N_14596,N_14326);
or UO_837 (O_837,N_13885,N_14495);
nor UO_838 (O_838,N_14305,N_14304);
xor UO_839 (O_839,N_14214,N_14168);
nand UO_840 (O_840,N_14267,N_13672);
nand UO_841 (O_841,N_14381,N_13705);
and UO_842 (O_842,N_14473,N_14891);
and UO_843 (O_843,N_14456,N_14534);
nand UO_844 (O_844,N_13916,N_13525);
nand UO_845 (O_845,N_14747,N_14803);
and UO_846 (O_846,N_14895,N_14034);
nor UO_847 (O_847,N_14137,N_14487);
and UO_848 (O_848,N_14477,N_14320);
nor UO_849 (O_849,N_14490,N_14660);
or UO_850 (O_850,N_14805,N_14605);
nand UO_851 (O_851,N_13620,N_13664);
nor UO_852 (O_852,N_13512,N_14997);
nor UO_853 (O_853,N_14477,N_14705);
nand UO_854 (O_854,N_14482,N_14220);
xor UO_855 (O_855,N_13698,N_13564);
nor UO_856 (O_856,N_14165,N_14222);
nand UO_857 (O_857,N_14037,N_13613);
or UO_858 (O_858,N_14393,N_14001);
nand UO_859 (O_859,N_14415,N_14769);
and UO_860 (O_860,N_14801,N_13675);
xnor UO_861 (O_861,N_14278,N_13820);
nand UO_862 (O_862,N_14231,N_14491);
and UO_863 (O_863,N_13962,N_14365);
nand UO_864 (O_864,N_14226,N_14798);
nor UO_865 (O_865,N_14822,N_14929);
or UO_866 (O_866,N_14748,N_14948);
nand UO_867 (O_867,N_14954,N_14362);
or UO_868 (O_868,N_14451,N_14513);
or UO_869 (O_869,N_13706,N_14103);
and UO_870 (O_870,N_13505,N_14023);
or UO_871 (O_871,N_13536,N_14524);
and UO_872 (O_872,N_14686,N_14110);
xor UO_873 (O_873,N_13503,N_14957);
or UO_874 (O_874,N_14614,N_14394);
or UO_875 (O_875,N_13876,N_14746);
nand UO_876 (O_876,N_14943,N_14520);
and UO_877 (O_877,N_14991,N_14044);
and UO_878 (O_878,N_14194,N_14398);
or UO_879 (O_879,N_13777,N_13758);
nand UO_880 (O_880,N_14986,N_14906);
nand UO_881 (O_881,N_13634,N_14705);
nand UO_882 (O_882,N_14908,N_13930);
and UO_883 (O_883,N_14694,N_14862);
xor UO_884 (O_884,N_14533,N_14140);
nor UO_885 (O_885,N_14427,N_13958);
and UO_886 (O_886,N_13903,N_14556);
or UO_887 (O_887,N_14870,N_13803);
and UO_888 (O_888,N_14193,N_14972);
or UO_889 (O_889,N_14971,N_13967);
and UO_890 (O_890,N_13569,N_13709);
nor UO_891 (O_891,N_14780,N_14216);
xnor UO_892 (O_892,N_14975,N_14738);
nand UO_893 (O_893,N_14272,N_14834);
and UO_894 (O_894,N_14902,N_13581);
or UO_895 (O_895,N_14478,N_14879);
nand UO_896 (O_896,N_14884,N_14540);
nand UO_897 (O_897,N_13690,N_14834);
nand UO_898 (O_898,N_14989,N_14074);
and UO_899 (O_899,N_14730,N_14987);
nor UO_900 (O_900,N_14238,N_13938);
nand UO_901 (O_901,N_13701,N_14579);
nor UO_902 (O_902,N_14086,N_14841);
nand UO_903 (O_903,N_14743,N_14451);
nor UO_904 (O_904,N_14601,N_14129);
and UO_905 (O_905,N_14705,N_13662);
xnor UO_906 (O_906,N_13567,N_13719);
nand UO_907 (O_907,N_14356,N_14704);
or UO_908 (O_908,N_14751,N_13614);
or UO_909 (O_909,N_13650,N_13652);
and UO_910 (O_910,N_13688,N_14823);
xnor UO_911 (O_911,N_13925,N_14319);
and UO_912 (O_912,N_13906,N_13765);
and UO_913 (O_913,N_13803,N_13966);
nand UO_914 (O_914,N_14810,N_14973);
or UO_915 (O_915,N_14585,N_14581);
and UO_916 (O_916,N_14446,N_13695);
and UO_917 (O_917,N_14792,N_14672);
nor UO_918 (O_918,N_13595,N_13809);
or UO_919 (O_919,N_14359,N_14661);
and UO_920 (O_920,N_14905,N_14073);
nor UO_921 (O_921,N_14322,N_13968);
nand UO_922 (O_922,N_13529,N_14856);
nor UO_923 (O_923,N_13819,N_13993);
nor UO_924 (O_924,N_14527,N_14033);
nor UO_925 (O_925,N_14820,N_14651);
and UO_926 (O_926,N_13638,N_13891);
nand UO_927 (O_927,N_13993,N_14211);
nor UO_928 (O_928,N_14143,N_14504);
and UO_929 (O_929,N_14136,N_13718);
or UO_930 (O_930,N_13646,N_14183);
and UO_931 (O_931,N_14662,N_14829);
nor UO_932 (O_932,N_14098,N_13834);
nand UO_933 (O_933,N_14010,N_14068);
and UO_934 (O_934,N_14451,N_14760);
and UO_935 (O_935,N_13656,N_14751);
or UO_936 (O_936,N_14067,N_14027);
nand UO_937 (O_937,N_14018,N_14935);
and UO_938 (O_938,N_14702,N_14838);
xnor UO_939 (O_939,N_14541,N_14713);
and UO_940 (O_940,N_13860,N_14535);
or UO_941 (O_941,N_14435,N_13700);
nand UO_942 (O_942,N_14445,N_13561);
or UO_943 (O_943,N_14284,N_14358);
nand UO_944 (O_944,N_13598,N_14439);
and UO_945 (O_945,N_14827,N_14970);
nand UO_946 (O_946,N_14430,N_13856);
nand UO_947 (O_947,N_13679,N_14128);
nor UO_948 (O_948,N_13784,N_14247);
or UO_949 (O_949,N_13927,N_14956);
or UO_950 (O_950,N_13997,N_13577);
or UO_951 (O_951,N_14907,N_14887);
and UO_952 (O_952,N_14678,N_14252);
or UO_953 (O_953,N_13775,N_13941);
nand UO_954 (O_954,N_14010,N_13809);
and UO_955 (O_955,N_14040,N_13564);
or UO_956 (O_956,N_14034,N_13805);
xnor UO_957 (O_957,N_13679,N_13995);
xnor UO_958 (O_958,N_14607,N_13770);
nor UO_959 (O_959,N_14083,N_13572);
or UO_960 (O_960,N_14220,N_13542);
nand UO_961 (O_961,N_14397,N_14265);
nand UO_962 (O_962,N_13614,N_14588);
nand UO_963 (O_963,N_14596,N_14245);
and UO_964 (O_964,N_14005,N_14762);
xnor UO_965 (O_965,N_14384,N_14855);
nor UO_966 (O_966,N_13650,N_14025);
or UO_967 (O_967,N_14587,N_13938);
nand UO_968 (O_968,N_13974,N_14125);
nand UO_969 (O_969,N_13843,N_14814);
nand UO_970 (O_970,N_14759,N_14763);
and UO_971 (O_971,N_14186,N_14640);
nand UO_972 (O_972,N_13726,N_13920);
nand UO_973 (O_973,N_13996,N_14133);
nor UO_974 (O_974,N_13772,N_14131);
nor UO_975 (O_975,N_14983,N_14895);
nor UO_976 (O_976,N_13955,N_14553);
and UO_977 (O_977,N_14879,N_14963);
nor UO_978 (O_978,N_14584,N_14009);
xor UO_979 (O_979,N_14746,N_14542);
or UO_980 (O_980,N_13569,N_13513);
and UO_981 (O_981,N_14593,N_14968);
or UO_982 (O_982,N_14757,N_14732);
nand UO_983 (O_983,N_14894,N_14184);
nor UO_984 (O_984,N_13849,N_14861);
and UO_985 (O_985,N_14605,N_14085);
nand UO_986 (O_986,N_14208,N_14961);
and UO_987 (O_987,N_14912,N_13901);
nor UO_988 (O_988,N_14132,N_14582);
and UO_989 (O_989,N_14772,N_14599);
and UO_990 (O_990,N_14719,N_13784);
and UO_991 (O_991,N_14249,N_14813);
nor UO_992 (O_992,N_14907,N_14726);
or UO_993 (O_993,N_14410,N_14477);
xnor UO_994 (O_994,N_14048,N_14316);
and UO_995 (O_995,N_14513,N_14845);
or UO_996 (O_996,N_14355,N_14518);
nand UO_997 (O_997,N_14173,N_14812);
nor UO_998 (O_998,N_14350,N_13766);
and UO_999 (O_999,N_14133,N_14276);
nand UO_1000 (O_1000,N_14027,N_14177);
and UO_1001 (O_1001,N_13706,N_14682);
nor UO_1002 (O_1002,N_14053,N_14893);
nand UO_1003 (O_1003,N_13703,N_14296);
xor UO_1004 (O_1004,N_13836,N_13710);
or UO_1005 (O_1005,N_14445,N_14165);
nor UO_1006 (O_1006,N_13887,N_13683);
xnor UO_1007 (O_1007,N_13595,N_14292);
nand UO_1008 (O_1008,N_13947,N_13894);
and UO_1009 (O_1009,N_14881,N_13978);
or UO_1010 (O_1010,N_14035,N_14491);
nand UO_1011 (O_1011,N_13682,N_14480);
nor UO_1012 (O_1012,N_14048,N_13643);
nor UO_1013 (O_1013,N_13875,N_13748);
and UO_1014 (O_1014,N_14474,N_13606);
nor UO_1015 (O_1015,N_14236,N_13537);
and UO_1016 (O_1016,N_14031,N_13500);
nor UO_1017 (O_1017,N_14780,N_14739);
nand UO_1018 (O_1018,N_14420,N_13717);
and UO_1019 (O_1019,N_14308,N_14600);
and UO_1020 (O_1020,N_14643,N_13912);
nand UO_1021 (O_1021,N_13854,N_13645);
nand UO_1022 (O_1022,N_14519,N_14296);
xor UO_1023 (O_1023,N_14339,N_14883);
nor UO_1024 (O_1024,N_13698,N_13800);
nand UO_1025 (O_1025,N_13981,N_14384);
and UO_1026 (O_1026,N_13863,N_14509);
nand UO_1027 (O_1027,N_14712,N_14481);
nand UO_1028 (O_1028,N_14546,N_13583);
nand UO_1029 (O_1029,N_14742,N_14349);
nand UO_1030 (O_1030,N_13733,N_13715);
nor UO_1031 (O_1031,N_14497,N_13538);
nor UO_1032 (O_1032,N_13536,N_14783);
or UO_1033 (O_1033,N_14993,N_14341);
nor UO_1034 (O_1034,N_13656,N_13711);
nand UO_1035 (O_1035,N_14356,N_13885);
or UO_1036 (O_1036,N_14157,N_13991);
nor UO_1037 (O_1037,N_13751,N_13814);
nand UO_1038 (O_1038,N_13686,N_13591);
nor UO_1039 (O_1039,N_14926,N_14530);
and UO_1040 (O_1040,N_14636,N_13741);
nand UO_1041 (O_1041,N_14127,N_14716);
nand UO_1042 (O_1042,N_13654,N_14216);
and UO_1043 (O_1043,N_14917,N_14098);
nor UO_1044 (O_1044,N_14768,N_13682);
nor UO_1045 (O_1045,N_14755,N_14920);
nor UO_1046 (O_1046,N_13583,N_14519);
nor UO_1047 (O_1047,N_14437,N_13761);
and UO_1048 (O_1048,N_13736,N_14132);
or UO_1049 (O_1049,N_14861,N_13744);
or UO_1050 (O_1050,N_14905,N_14993);
or UO_1051 (O_1051,N_14285,N_14123);
xor UO_1052 (O_1052,N_14505,N_13847);
nand UO_1053 (O_1053,N_13821,N_14414);
nor UO_1054 (O_1054,N_14362,N_14542);
nand UO_1055 (O_1055,N_14632,N_13604);
or UO_1056 (O_1056,N_13904,N_14577);
or UO_1057 (O_1057,N_13735,N_13559);
or UO_1058 (O_1058,N_13735,N_14953);
nand UO_1059 (O_1059,N_14285,N_14081);
nor UO_1060 (O_1060,N_13918,N_13777);
and UO_1061 (O_1061,N_14720,N_14792);
nor UO_1062 (O_1062,N_14786,N_14406);
nand UO_1063 (O_1063,N_14883,N_14624);
or UO_1064 (O_1064,N_13588,N_13959);
nor UO_1065 (O_1065,N_14300,N_14387);
nand UO_1066 (O_1066,N_13823,N_14976);
nand UO_1067 (O_1067,N_13763,N_14809);
and UO_1068 (O_1068,N_14536,N_13984);
and UO_1069 (O_1069,N_14162,N_13916);
or UO_1070 (O_1070,N_14355,N_14703);
nor UO_1071 (O_1071,N_14852,N_14297);
and UO_1072 (O_1072,N_13990,N_14405);
or UO_1073 (O_1073,N_14572,N_14867);
or UO_1074 (O_1074,N_14168,N_14269);
nor UO_1075 (O_1075,N_13772,N_14085);
xnor UO_1076 (O_1076,N_14830,N_13999);
nand UO_1077 (O_1077,N_13655,N_13690);
nand UO_1078 (O_1078,N_14324,N_13984);
or UO_1079 (O_1079,N_14819,N_13831);
nand UO_1080 (O_1080,N_13715,N_14163);
or UO_1081 (O_1081,N_14468,N_13875);
nand UO_1082 (O_1082,N_13840,N_14515);
xnor UO_1083 (O_1083,N_13565,N_13581);
and UO_1084 (O_1084,N_13967,N_14694);
nand UO_1085 (O_1085,N_14768,N_13766);
and UO_1086 (O_1086,N_14067,N_14188);
and UO_1087 (O_1087,N_14993,N_14384);
or UO_1088 (O_1088,N_13905,N_14073);
and UO_1089 (O_1089,N_13529,N_14163);
and UO_1090 (O_1090,N_13598,N_14345);
nand UO_1091 (O_1091,N_14600,N_14614);
and UO_1092 (O_1092,N_13855,N_13933);
nor UO_1093 (O_1093,N_13915,N_14529);
nand UO_1094 (O_1094,N_13983,N_13501);
and UO_1095 (O_1095,N_13561,N_13740);
and UO_1096 (O_1096,N_14827,N_14133);
nand UO_1097 (O_1097,N_14599,N_13687);
nand UO_1098 (O_1098,N_13964,N_14238);
xnor UO_1099 (O_1099,N_13556,N_13565);
or UO_1100 (O_1100,N_13607,N_14529);
nand UO_1101 (O_1101,N_13582,N_14314);
xnor UO_1102 (O_1102,N_13624,N_14690);
or UO_1103 (O_1103,N_13702,N_14434);
nand UO_1104 (O_1104,N_14850,N_13937);
and UO_1105 (O_1105,N_14325,N_14152);
and UO_1106 (O_1106,N_14515,N_14404);
and UO_1107 (O_1107,N_14846,N_14520);
nand UO_1108 (O_1108,N_14071,N_14590);
nor UO_1109 (O_1109,N_14929,N_13812);
and UO_1110 (O_1110,N_13525,N_14854);
or UO_1111 (O_1111,N_14660,N_13553);
nor UO_1112 (O_1112,N_14227,N_14701);
or UO_1113 (O_1113,N_13920,N_14625);
or UO_1114 (O_1114,N_13748,N_13996);
and UO_1115 (O_1115,N_14805,N_13597);
nor UO_1116 (O_1116,N_14100,N_13784);
nand UO_1117 (O_1117,N_13795,N_14581);
nor UO_1118 (O_1118,N_14201,N_13827);
nand UO_1119 (O_1119,N_14121,N_14706);
or UO_1120 (O_1120,N_14224,N_14149);
nand UO_1121 (O_1121,N_14646,N_14693);
nand UO_1122 (O_1122,N_14388,N_14392);
nor UO_1123 (O_1123,N_14107,N_13991);
or UO_1124 (O_1124,N_13661,N_13600);
nand UO_1125 (O_1125,N_13692,N_14377);
and UO_1126 (O_1126,N_14992,N_14556);
and UO_1127 (O_1127,N_13713,N_13817);
or UO_1128 (O_1128,N_14456,N_13614);
and UO_1129 (O_1129,N_14732,N_14958);
and UO_1130 (O_1130,N_14391,N_14285);
xnor UO_1131 (O_1131,N_13913,N_14157);
nor UO_1132 (O_1132,N_13721,N_13623);
and UO_1133 (O_1133,N_13516,N_13502);
or UO_1134 (O_1134,N_14505,N_13677);
or UO_1135 (O_1135,N_14067,N_14704);
nor UO_1136 (O_1136,N_13521,N_14774);
and UO_1137 (O_1137,N_14092,N_14078);
nor UO_1138 (O_1138,N_14868,N_13670);
and UO_1139 (O_1139,N_14233,N_13939);
nor UO_1140 (O_1140,N_14390,N_14198);
xnor UO_1141 (O_1141,N_13829,N_13846);
and UO_1142 (O_1142,N_13516,N_13616);
and UO_1143 (O_1143,N_14266,N_14122);
or UO_1144 (O_1144,N_13871,N_14208);
nor UO_1145 (O_1145,N_14712,N_13987);
nand UO_1146 (O_1146,N_14630,N_13526);
or UO_1147 (O_1147,N_14699,N_13777);
xor UO_1148 (O_1148,N_13813,N_14751);
nand UO_1149 (O_1149,N_14645,N_14969);
or UO_1150 (O_1150,N_13585,N_14267);
nor UO_1151 (O_1151,N_13545,N_13514);
nand UO_1152 (O_1152,N_14576,N_13583);
nor UO_1153 (O_1153,N_14593,N_14112);
and UO_1154 (O_1154,N_14905,N_14456);
nor UO_1155 (O_1155,N_14488,N_14356);
nor UO_1156 (O_1156,N_13658,N_13776);
xor UO_1157 (O_1157,N_13674,N_14168);
nor UO_1158 (O_1158,N_13975,N_14122);
nand UO_1159 (O_1159,N_13563,N_14418);
nand UO_1160 (O_1160,N_13825,N_14187);
nand UO_1161 (O_1161,N_14593,N_14487);
nand UO_1162 (O_1162,N_13780,N_14349);
and UO_1163 (O_1163,N_13816,N_14789);
xor UO_1164 (O_1164,N_13829,N_13965);
or UO_1165 (O_1165,N_14411,N_14082);
or UO_1166 (O_1166,N_14035,N_14166);
and UO_1167 (O_1167,N_14420,N_13711);
nor UO_1168 (O_1168,N_14195,N_14386);
or UO_1169 (O_1169,N_14976,N_14910);
or UO_1170 (O_1170,N_13844,N_14000);
and UO_1171 (O_1171,N_14603,N_14315);
and UO_1172 (O_1172,N_14815,N_13853);
and UO_1173 (O_1173,N_14745,N_14273);
nand UO_1174 (O_1174,N_14395,N_14977);
and UO_1175 (O_1175,N_14913,N_13872);
nor UO_1176 (O_1176,N_14310,N_14948);
and UO_1177 (O_1177,N_13684,N_13888);
or UO_1178 (O_1178,N_14162,N_13587);
xor UO_1179 (O_1179,N_14448,N_14866);
or UO_1180 (O_1180,N_14161,N_14269);
and UO_1181 (O_1181,N_14310,N_14537);
nand UO_1182 (O_1182,N_14634,N_13983);
and UO_1183 (O_1183,N_14357,N_14127);
or UO_1184 (O_1184,N_14078,N_13592);
and UO_1185 (O_1185,N_13780,N_14075);
nand UO_1186 (O_1186,N_14542,N_14768);
and UO_1187 (O_1187,N_14610,N_14641);
nand UO_1188 (O_1188,N_14018,N_13547);
or UO_1189 (O_1189,N_14210,N_14550);
nand UO_1190 (O_1190,N_14016,N_14701);
nor UO_1191 (O_1191,N_13507,N_13634);
nor UO_1192 (O_1192,N_13835,N_14554);
or UO_1193 (O_1193,N_14524,N_14333);
nor UO_1194 (O_1194,N_13788,N_14956);
nor UO_1195 (O_1195,N_13505,N_14779);
nor UO_1196 (O_1196,N_14951,N_14081);
xnor UO_1197 (O_1197,N_13550,N_13564);
nor UO_1198 (O_1198,N_14473,N_13808);
xor UO_1199 (O_1199,N_13775,N_14338);
nor UO_1200 (O_1200,N_14295,N_13848);
or UO_1201 (O_1201,N_14150,N_14909);
nor UO_1202 (O_1202,N_14158,N_14098);
or UO_1203 (O_1203,N_14347,N_13510);
or UO_1204 (O_1204,N_14693,N_13601);
xnor UO_1205 (O_1205,N_13778,N_13861);
or UO_1206 (O_1206,N_14119,N_14741);
nor UO_1207 (O_1207,N_14978,N_14539);
and UO_1208 (O_1208,N_14269,N_14701);
xnor UO_1209 (O_1209,N_13639,N_13653);
and UO_1210 (O_1210,N_14996,N_13615);
nor UO_1211 (O_1211,N_14687,N_14289);
and UO_1212 (O_1212,N_14997,N_14595);
or UO_1213 (O_1213,N_13555,N_13868);
nor UO_1214 (O_1214,N_14435,N_13778);
nor UO_1215 (O_1215,N_13580,N_13696);
nand UO_1216 (O_1216,N_13505,N_13877);
and UO_1217 (O_1217,N_14083,N_14084);
nor UO_1218 (O_1218,N_14042,N_14556);
nand UO_1219 (O_1219,N_14253,N_13801);
or UO_1220 (O_1220,N_13860,N_14718);
nor UO_1221 (O_1221,N_13641,N_14494);
nand UO_1222 (O_1222,N_13733,N_14370);
nor UO_1223 (O_1223,N_14592,N_13895);
nor UO_1224 (O_1224,N_13627,N_14215);
or UO_1225 (O_1225,N_14071,N_14887);
nand UO_1226 (O_1226,N_14195,N_13804);
nor UO_1227 (O_1227,N_13515,N_14530);
nor UO_1228 (O_1228,N_14923,N_14596);
and UO_1229 (O_1229,N_14429,N_14272);
nor UO_1230 (O_1230,N_14339,N_13734);
nor UO_1231 (O_1231,N_14660,N_14579);
and UO_1232 (O_1232,N_13785,N_13876);
xor UO_1233 (O_1233,N_13572,N_14646);
nand UO_1234 (O_1234,N_14881,N_13590);
and UO_1235 (O_1235,N_14115,N_14495);
nand UO_1236 (O_1236,N_14495,N_14853);
and UO_1237 (O_1237,N_13978,N_14901);
nor UO_1238 (O_1238,N_14816,N_13923);
or UO_1239 (O_1239,N_13729,N_14574);
nor UO_1240 (O_1240,N_14958,N_14143);
nor UO_1241 (O_1241,N_13765,N_14162);
nor UO_1242 (O_1242,N_14916,N_13983);
or UO_1243 (O_1243,N_13958,N_14217);
nor UO_1244 (O_1244,N_14866,N_14617);
and UO_1245 (O_1245,N_14357,N_14289);
or UO_1246 (O_1246,N_13642,N_14826);
nand UO_1247 (O_1247,N_14676,N_13938);
nand UO_1248 (O_1248,N_14945,N_14231);
or UO_1249 (O_1249,N_14764,N_13982);
and UO_1250 (O_1250,N_14824,N_14763);
nand UO_1251 (O_1251,N_14672,N_14858);
and UO_1252 (O_1252,N_14386,N_14800);
and UO_1253 (O_1253,N_14281,N_13629);
and UO_1254 (O_1254,N_13524,N_14188);
or UO_1255 (O_1255,N_14384,N_14312);
or UO_1256 (O_1256,N_14218,N_13759);
and UO_1257 (O_1257,N_14230,N_14867);
or UO_1258 (O_1258,N_14310,N_14341);
xnor UO_1259 (O_1259,N_13763,N_13657);
and UO_1260 (O_1260,N_14563,N_14782);
and UO_1261 (O_1261,N_14115,N_13793);
xor UO_1262 (O_1262,N_14184,N_14396);
or UO_1263 (O_1263,N_13949,N_13951);
nand UO_1264 (O_1264,N_14213,N_14095);
nand UO_1265 (O_1265,N_14665,N_13959);
nor UO_1266 (O_1266,N_14054,N_13857);
nor UO_1267 (O_1267,N_13648,N_14475);
and UO_1268 (O_1268,N_14074,N_13897);
nor UO_1269 (O_1269,N_14249,N_14694);
or UO_1270 (O_1270,N_14179,N_14919);
xnor UO_1271 (O_1271,N_13702,N_14929);
nand UO_1272 (O_1272,N_14160,N_14480);
and UO_1273 (O_1273,N_13679,N_14748);
nand UO_1274 (O_1274,N_14857,N_13800);
nand UO_1275 (O_1275,N_14694,N_13787);
nor UO_1276 (O_1276,N_14926,N_13502);
or UO_1277 (O_1277,N_14477,N_14162);
and UO_1278 (O_1278,N_14658,N_13811);
nand UO_1279 (O_1279,N_14364,N_14994);
and UO_1280 (O_1280,N_13820,N_14412);
nor UO_1281 (O_1281,N_14770,N_13997);
and UO_1282 (O_1282,N_13656,N_13680);
and UO_1283 (O_1283,N_14365,N_13587);
nand UO_1284 (O_1284,N_14304,N_13510);
or UO_1285 (O_1285,N_14526,N_13550);
and UO_1286 (O_1286,N_13989,N_14514);
nand UO_1287 (O_1287,N_13999,N_14410);
nand UO_1288 (O_1288,N_14585,N_13886);
and UO_1289 (O_1289,N_14307,N_13945);
or UO_1290 (O_1290,N_14732,N_14727);
and UO_1291 (O_1291,N_14456,N_14794);
nand UO_1292 (O_1292,N_14160,N_14516);
nor UO_1293 (O_1293,N_14640,N_14103);
and UO_1294 (O_1294,N_14335,N_14511);
nor UO_1295 (O_1295,N_13699,N_13547);
xor UO_1296 (O_1296,N_14520,N_13744);
and UO_1297 (O_1297,N_14017,N_14102);
nand UO_1298 (O_1298,N_14246,N_14406);
or UO_1299 (O_1299,N_14514,N_13520);
nor UO_1300 (O_1300,N_14714,N_13886);
nor UO_1301 (O_1301,N_13842,N_14414);
nor UO_1302 (O_1302,N_14651,N_14695);
xnor UO_1303 (O_1303,N_14560,N_14687);
nor UO_1304 (O_1304,N_14823,N_14221);
nand UO_1305 (O_1305,N_14225,N_14345);
or UO_1306 (O_1306,N_14447,N_14740);
nor UO_1307 (O_1307,N_14714,N_13840);
and UO_1308 (O_1308,N_14718,N_13583);
xnor UO_1309 (O_1309,N_14665,N_13939);
or UO_1310 (O_1310,N_14877,N_14553);
or UO_1311 (O_1311,N_14454,N_13888);
or UO_1312 (O_1312,N_14763,N_14393);
nand UO_1313 (O_1313,N_14121,N_14796);
nand UO_1314 (O_1314,N_14605,N_13895);
nand UO_1315 (O_1315,N_14981,N_13971);
nand UO_1316 (O_1316,N_14470,N_13616);
nor UO_1317 (O_1317,N_13511,N_14420);
nand UO_1318 (O_1318,N_13738,N_13978);
or UO_1319 (O_1319,N_14749,N_14219);
or UO_1320 (O_1320,N_14520,N_14624);
or UO_1321 (O_1321,N_14004,N_13616);
nor UO_1322 (O_1322,N_13811,N_14410);
and UO_1323 (O_1323,N_13790,N_14173);
xor UO_1324 (O_1324,N_13815,N_13989);
nand UO_1325 (O_1325,N_13666,N_14983);
nand UO_1326 (O_1326,N_13700,N_14006);
or UO_1327 (O_1327,N_13781,N_14619);
or UO_1328 (O_1328,N_14962,N_14283);
xor UO_1329 (O_1329,N_13581,N_14116);
nor UO_1330 (O_1330,N_14248,N_14471);
and UO_1331 (O_1331,N_14079,N_14474);
or UO_1332 (O_1332,N_14601,N_14237);
or UO_1333 (O_1333,N_14562,N_14670);
and UO_1334 (O_1334,N_13925,N_14647);
or UO_1335 (O_1335,N_13529,N_14907);
nor UO_1336 (O_1336,N_14256,N_14204);
nand UO_1337 (O_1337,N_14645,N_14079);
or UO_1338 (O_1338,N_14484,N_14093);
xnor UO_1339 (O_1339,N_14255,N_14654);
and UO_1340 (O_1340,N_14218,N_14201);
or UO_1341 (O_1341,N_13599,N_14663);
nor UO_1342 (O_1342,N_14702,N_14849);
and UO_1343 (O_1343,N_13954,N_14214);
nand UO_1344 (O_1344,N_14529,N_14713);
nor UO_1345 (O_1345,N_14253,N_13945);
nor UO_1346 (O_1346,N_14652,N_13775);
and UO_1347 (O_1347,N_14283,N_14780);
nand UO_1348 (O_1348,N_13986,N_14539);
or UO_1349 (O_1349,N_14547,N_14762);
nand UO_1350 (O_1350,N_13999,N_13971);
or UO_1351 (O_1351,N_14263,N_14057);
nor UO_1352 (O_1352,N_13907,N_13677);
nand UO_1353 (O_1353,N_13833,N_14192);
and UO_1354 (O_1354,N_13862,N_14697);
or UO_1355 (O_1355,N_14390,N_13938);
nor UO_1356 (O_1356,N_14970,N_14041);
xnor UO_1357 (O_1357,N_14705,N_14351);
or UO_1358 (O_1358,N_14211,N_13641);
nor UO_1359 (O_1359,N_14341,N_14260);
and UO_1360 (O_1360,N_13583,N_14757);
or UO_1361 (O_1361,N_14139,N_13823);
or UO_1362 (O_1362,N_14873,N_13946);
xor UO_1363 (O_1363,N_13608,N_14804);
nand UO_1364 (O_1364,N_13546,N_14734);
nor UO_1365 (O_1365,N_14741,N_14983);
or UO_1366 (O_1366,N_14599,N_13562);
or UO_1367 (O_1367,N_14885,N_14553);
and UO_1368 (O_1368,N_14541,N_14607);
and UO_1369 (O_1369,N_14138,N_13987);
or UO_1370 (O_1370,N_13969,N_14592);
xor UO_1371 (O_1371,N_14863,N_14795);
nor UO_1372 (O_1372,N_14996,N_13791);
or UO_1373 (O_1373,N_14430,N_14186);
xor UO_1374 (O_1374,N_14328,N_13944);
xor UO_1375 (O_1375,N_13847,N_13700);
or UO_1376 (O_1376,N_13585,N_14590);
and UO_1377 (O_1377,N_13904,N_14228);
nor UO_1378 (O_1378,N_14440,N_14083);
nor UO_1379 (O_1379,N_14202,N_14953);
nor UO_1380 (O_1380,N_14441,N_14137);
and UO_1381 (O_1381,N_13898,N_13527);
nand UO_1382 (O_1382,N_14307,N_14525);
and UO_1383 (O_1383,N_14791,N_13665);
nand UO_1384 (O_1384,N_13828,N_14659);
or UO_1385 (O_1385,N_14601,N_14670);
nand UO_1386 (O_1386,N_13719,N_13976);
nand UO_1387 (O_1387,N_13983,N_14828);
nand UO_1388 (O_1388,N_14091,N_13652);
xor UO_1389 (O_1389,N_14397,N_14529);
and UO_1390 (O_1390,N_13659,N_14811);
nor UO_1391 (O_1391,N_14456,N_14740);
and UO_1392 (O_1392,N_14009,N_14416);
or UO_1393 (O_1393,N_14145,N_14265);
nor UO_1394 (O_1394,N_14679,N_14970);
and UO_1395 (O_1395,N_13906,N_14995);
or UO_1396 (O_1396,N_13736,N_14890);
or UO_1397 (O_1397,N_14606,N_14336);
or UO_1398 (O_1398,N_13660,N_14410);
or UO_1399 (O_1399,N_14195,N_14696);
and UO_1400 (O_1400,N_13505,N_14784);
and UO_1401 (O_1401,N_14804,N_13530);
and UO_1402 (O_1402,N_13918,N_14348);
xor UO_1403 (O_1403,N_14476,N_14781);
nor UO_1404 (O_1404,N_13547,N_14255);
nor UO_1405 (O_1405,N_14445,N_14908);
nand UO_1406 (O_1406,N_14599,N_14748);
nor UO_1407 (O_1407,N_13957,N_14138);
nand UO_1408 (O_1408,N_14820,N_14552);
nand UO_1409 (O_1409,N_13602,N_13998);
and UO_1410 (O_1410,N_14293,N_14144);
or UO_1411 (O_1411,N_14041,N_14962);
or UO_1412 (O_1412,N_14762,N_14706);
nand UO_1413 (O_1413,N_14246,N_14942);
xor UO_1414 (O_1414,N_14033,N_13848);
and UO_1415 (O_1415,N_14908,N_14275);
nor UO_1416 (O_1416,N_14928,N_13517);
nor UO_1417 (O_1417,N_14226,N_14073);
and UO_1418 (O_1418,N_14159,N_14600);
nor UO_1419 (O_1419,N_14922,N_13787);
nor UO_1420 (O_1420,N_13917,N_14692);
nor UO_1421 (O_1421,N_13825,N_13763);
nor UO_1422 (O_1422,N_14737,N_13871);
xor UO_1423 (O_1423,N_13761,N_14713);
nand UO_1424 (O_1424,N_13770,N_14163);
nand UO_1425 (O_1425,N_14233,N_13530);
nor UO_1426 (O_1426,N_14669,N_13601);
nand UO_1427 (O_1427,N_14766,N_14844);
nand UO_1428 (O_1428,N_14666,N_14342);
nand UO_1429 (O_1429,N_14440,N_13958);
nor UO_1430 (O_1430,N_14132,N_14897);
xor UO_1431 (O_1431,N_13553,N_14362);
and UO_1432 (O_1432,N_13667,N_13719);
and UO_1433 (O_1433,N_14922,N_14419);
nand UO_1434 (O_1434,N_14290,N_14006);
and UO_1435 (O_1435,N_13873,N_13775);
or UO_1436 (O_1436,N_14351,N_14671);
nand UO_1437 (O_1437,N_13789,N_14859);
nor UO_1438 (O_1438,N_14344,N_14612);
xor UO_1439 (O_1439,N_14168,N_14663);
nand UO_1440 (O_1440,N_14671,N_14486);
and UO_1441 (O_1441,N_13693,N_14556);
nand UO_1442 (O_1442,N_14764,N_14987);
and UO_1443 (O_1443,N_14977,N_14328);
nor UO_1444 (O_1444,N_13619,N_14392);
nor UO_1445 (O_1445,N_14429,N_13864);
and UO_1446 (O_1446,N_14387,N_14814);
nor UO_1447 (O_1447,N_14471,N_13799);
or UO_1448 (O_1448,N_14426,N_14295);
nor UO_1449 (O_1449,N_14581,N_13530);
or UO_1450 (O_1450,N_13792,N_13791);
and UO_1451 (O_1451,N_14574,N_13629);
xor UO_1452 (O_1452,N_14079,N_14497);
nor UO_1453 (O_1453,N_14602,N_13634);
nand UO_1454 (O_1454,N_14972,N_14720);
and UO_1455 (O_1455,N_14683,N_14705);
nand UO_1456 (O_1456,N_13908,N_13777);
nand UO_1457 (O_1457,N_14743,N_13640);
nand UO_1458 (O_1458,N_14778,N_14139);
nand UO_1459 (O_1459,N_13960,N_14592);
nand UO_1460 (O_1460,N_14445,N_13623);
and UO_1461 (O_1461,N_14560,N_13781);
xor UO_1462 (O_1462,N_14703,N_14509);
and UO_1463 (O_1463,N_14977,N_14855);
nand UO_1464 (O_1464,N_14354,N_14211);
xnor UO_1465 (O_1465,N_14296,N_14746);
nor UO_1466 (O_1466,N_14781,N_14027);
nand UO_1467 (O_1467,N_14733,N_14845);
and UO_1468 (O_1468,N_14149,N_14942);
or UO_1469 (O_1469,N_14956,N_14712);
or UO_1470 (O_1470,N_14907,N_13734);
and UO_1471 (O_1471,N_14711,N_13989);
or UO_1472 (O_1472,N_14014,N_14297);
and UO_1473 (O_1473,N_14257,N_14521);
or UO_1474 (O_1474,N_14005,N_13750);
or UO_1475 (O_1475,N_13932,N_13526);
and UO_1476 (O_1476,N_14113,N_14228);
nand UO_1477 (O_1477,N_13920,N_14719);
or UO_1478 (O_1478,N_14837,N_14523);
nand UO_1479 (O_1479,N_13539,N_13926);
nor UO_1480 (O_1480,N_14149,N_14074);
and UO_1481 (O_1481,N_13951,N_14246);
or UO_1482 (O_1482,N_13976,N_14311);
nand UO_1483 (O_1483,N_13556,N_13883);
or UO_1484 (O_1484,N_14414,N_13848);
and UO_1485 (O_1485,N_14362,N_13580);
nor UO_1486 (O_1486,N_13925,N_14366);
and UO_1487 (O_1487,N_13532,N_13750);
nand UO_1488 (O_1488,N_14840,N_13847);
or UO_1489 (O_1489,N_14433,N_14827);
nor UO_1490 (O_1490,N_14810,N_14301);
nand UO_1491 (O_1491,N_13877,N_14258);
and UO_1492 (O_1492,N_14909,N_14765);
nor UO_1493 (O_1493,N_14998,N_14792);
nor UO_1494 (O_1494,N_14657,N_13840);
nor UO_1495 (O_1495,N_13681,N_14059);
nor UO_1496 (O_1496,N_14569,N_13857);
or UO_1497 (O_1497,N_14494,N_14133);
nor UO_1498 (O_1498,N_14865,N_14702);
or UO_1499 (O_1499,N_14489,N_14713);
nand UO_1500 (O_1500,N_14649,N_13574);
nor UO_1501 (O_1501,N_14066,N_13970);
nand UO_1502 (O_1502,N_14841,N_13856);
xor UO_1503 (O_1503,N_13852,N_13986);
nand UO_1504 (O_1504,N_14597,N_14418);
or UO_1505 (O_1505,N_14708,N_14680);
nand UO_1506 (O_1506,N_14300,N_14043);
nand UO_1507 (O_1507,N_13994,N_14673);
or UO_1508 (O_1508,N_14553,N_14699);
and UO_1509 (O_1509,N_14946,N_14759);
and UO_1510 (O_1510,N_14296,N_14142);
or UO_1511 (O_1511,N_14862,N_14539);
nand UO_1512 (O_1512,N_14723,N_14913);
and UO_1513 (O_1513,N_13594,N_13668);
nand UO_1514 (O_1514,N_13985,N_14161);
nand UO_1515 (O_1515,N_14237,N_13603);
nand UO_1516 (O_1516,N_14659,N_14636);
or UO_1517 (O_1517,N_13875,N_14978);
and UO_1518 (O_1518,N_14919,N_14141);
and UO_1519 (O_1519,N_14742,N_14823);
or UO_1520 (O_1520,N_13782,N_14280);
nand UO_1521 (O_1521,N_14632,N_13801);
and UO_1522 (O_1522,N_14817,N_14049);
or UO_1523 (O_1523,N_14713,N_13639);
nand UO_1524 (O_1524,N_13712,N_14496);
or UO_1525 (O_1525,N_13752,N_14145);
nand UO_1526 (O_1526,N_14239,N_14825);
and UO_1527 (O_1527,N_14941,N_13573);
and UO_1528 (O_1528,N_13792,N_14090);
and UO_1529 (O_1529,N_14981,N_13561);
nor UO_1530 (O_1530,N_14793,N_13608);
and UO_1531 (O_1531,N_14265,N_14965);
nor UO_1532 (O_1532,N_14836,N_13658);
and UO_1533 (O_1533,N_13986,N_14083);
and UO_1534 (O_1534,N_14648,N_14393);
nand UO_1535 (O_1535,N_14326,N_14450);
and UO_1536 (O_1536,N_13767,N_14816);
nand UO_1537 (O_1537,N_14766,N_14840);
or UO_1538 (O_1538,N_13569,N_14275);
nand UO_1539 (O_1539,N_14682,N_13531);
nand UO_1540 (O_1540,N_14933,N_14790);
nor UO_1541 (O_1541,N_14333,N_13643);
and UO_1542 (O_1542,N_14857,N_14276);
xnor UO_1543 (O_1543,N_13916,N_14687);
or UO_1544 (O_1544,N_14380,N_14318);
nor UO_1545 (O_1545,N_14609,N_14014);
and UO_1546 (O_1546,N_14993,N_13949);
xor UO_1547 (O_1547,N_13805,N_13759);
and UO_1548 (O_1548,N_13983,N_14431);
or UO_1549 (O_1549,N_14525,N_14346);
nor UO_1550 (O_1550,N_14240,N_13976);
xnor UO_1551 (O_1551,N_14007,N_14298);
nand UO_1552 (O_1552,N_14103,N_13979);
nand UO_1553 (O_1553,N_14962,N_14477);
nand UO_1554 (O_1554,N_13522,N_14122);
xnor UO_1555 (O_1555,N_14518,N_13575);
and UO_1556 (O_1556,N_14805,N_13700);
nor UO_1557 (O_1557,N_14562,N_14283);
nand UO_1558 (O_1558,N_13658,N_14050);
and UO_1559 (O_1559,N_14868,N_13683);
and UO_1560 (O_1560,N_13952,N_14366);
nor UO_1561 (O_1561,N_14465,N_13692);
and UO_1562 (O_1562,N_14465,N_14950);
nor UO_1563 (O_1563,N_14728,N_14799);
and UO_1564 (O_1564,N_14009,N_14813);
and UO_1565 (O_1565,N_14860,N_14692);
xor UO_1566 (O_1566,N_14762,N_14614);
and UO_1567 (O_1567,N_13642,N_14340);
or UO_1568 (O_1568,N_14663,N_13588);
nand UO_1569 (O_1569,N_13846,N_14818);
and UO_1570 (O_1570,N_13674,N_14418);
nor UO_1571 (O_1571,N_14863,N_14647);
nand UO_1572 (O_1572,N_13609,N_14830);
nor UO_1573 (O_1573,N_14713,N_14306);
or UO_1574 (O_1574,N_14492,N_13853);
nor UO_1575 (O_1575,N_13840,N_14977);
nor UO_1576 (O_1576,N_14668,N_14541);
nand UO_1577 (O_1577,N_14612,N_14334);
nand UO_1578 (O_1578,N_13821,N_14256);
and UO_1579 (O_1579,N_13589,N_13997);
nand UO_1580 (O_1580,N_14618,N_14273);
nand UO_1581 (O_1581,N_13889,N_13658);
nand UO_1582 (O_1582,N_14114,N_14790);
and UO_1583 (O_1583,N_14051,N_14237);
nor UO_1584 (O_1584,N_14046,N_13536);
nor UO_1585 (O_1585,N_14868,N_14014);
nor UO_1586 (O_1586,N_14891,N_14235);
or UO_1587 (O_1587,N_14357,N_13623);
nand UO_1588 (O_1588,N_14784,N_14427);
or UO_1589 (O_1589,N_13879,N_13948);
nor UO_1590 (O_1590,N_14962,N_14147);
nor UO_1591 (O_1591,N_13673,N_13577);
and UO_1592 (O_1592,N_14937,N_13974);
xor UO_1593 (O_1593,N_13576,N_14370);
nor UO_1594 (O_1594,N_14061,N_14728);
xor UO_1595 (O_1595,N_14212,N_13594);
nor UO_1596 (O_1596,N_14849,N_13650);
nand UO_1597 (O_1597,N_13930,N_14881);
nor UO_1598 (O_1598,N_14377,N_13849);
nand UO_1599 (O_1599,N_13597,N_13529);
nor UO_1600 (O_1600,N_13901,N_14693);
xnor UO_1601 (O_1601,N_14843,N_13580);
or UO_1602 (O_1602,N_13754,N_13626);
xnor UO_1603 (O_1603,N_14664,N_14528);
nor UO_1604 (O_1604,N_13777,N_14447);
and UO_1605 (O_1605,N_14604,N_13631);
or UO_1606 (O_1606,N_13810,N_14514);
nor UO_1607 (O_1607,N_13922,N_14850);
or UO_1608 (O_1608,N_13942,N_14433);
or UO_1609 (O_1609,N_13619,N_13888);
nand UO_1610 (O_1610,N_14384,N_14054);
and UO_1611 (O_1611,N_14829,N_14623);
nor UO_1612 (O_1612,N_14077,N_14902);
nor UO_1613 (O_1613,N_14013,N_13591);
and UO_1614 (O_1614,N_13702,N_14406);
and UO_1615 (O_1615,N_13818,N_13849);
nand UO_1616 (O_1616,N_14754,N_13811);
nor UO_1617 (O_1617,N_14434,N_14775);
nand UO_1618 (O_1618,N_13710,N_14729);
xor UO_1619 (O_1619,N_13703,N_13803);
or UO_1620 (O_1620,N_14873,N_14550);
and UO_1621 (O_1621,N_14080,N_13656);
nand UO_1622 (O_1622,N_14013,N_14899);
or UO_1623 (O_1623,N_14611,N_14524);
nor UO_1624 (O_1624,N_14228,N_13649);
xor UO_1625 (O_1625,N_14466,N_14244);
or UO_1626 (O_1626,N_14928,N_13894);
nor UO_1627 (O_1627,N_14208,N_14006);
xor UO_1628 (O_1628,N_14148,N_14178);
nand UO_1629 (O_1629,N_14102,N_14705);
or UO_1630 (O_1630,N_14256,N_13712);
or UO_1631 (O_1631,N_14898,N_13749);
and UO_1632 (O_1632,N_14670,N_14266);
xor UO_1633 (O_1633,N_14331,N_14653);
nand UO_1634 (O_1634,N_14885,N_14126);
or UO_1635 (O_1635,N_14157,N_13981);
nor UO_1636 (O_1636,N_14788,N_14089);
nor UO_1637 (O_1637,N_14368,N_14033);
nor UO_1638 (O_1638,N_14969,N_14028);
nor UO_1639 (O_1639,N_14763,N_14965);
or UO_1640 (O_1640,N_14817,N_14519);
or UO_1641 (O_1641,N_13732,N_14834);
and UO_1642 (O_1642,N_14101,N_13878);
xnor UO_1643 (O_1643,N_14419,N_14583);
nor UO_1644 (O_1644,N_13511,N_14004);
xor UO_1645 (O_1645,N_14840,N_13894);
nand UO_1646 (O_1646,N_14459,N_14679);
nor UO_1647 (O_1647,N_14099,N_13663);
nor UO_1648 (O_1648,N_14754,N_14128);
or UO_1649 (O_1649,N_14032,N_14865);
and UO_1650 (O_1650,N_14444,N_13811);
and UO_1651 (O_1651,N_14287,N_14158);
nor UO_1652 (O_1652,N_14743,N_14879);
nand UO_1653 (O_1653,N_13744,N_13843);
nor UO_1654 (O_1654,N_13630,N_13700);
or UO_1655 (O_1655,N_13657,N_14198);
nand UO_1656 (O_1656,N_13585,N_14499);
nand UO_1657 (O_1657,N_14623,N_14133);
and UO_1658 (O_1658,N_13654,N_13979);
and UO_1659 (O_1659,N_14965,N_14783);
nor UO_1660 (O_1660,N_13879,N_14680);
nor UO_1661 (O_1661,N_13730,N_14533);
nand UO_1662 (O_1662,N_14749,N_14957);
nor UO_1663 (O_1663,N_14440,N_13768);
or UO_1664 (O_1664,N_13556,N_14818);
nand UO_1665 (O_1665,N_13500,N_13809);
nand UO_1666 (O_1666,N_14849,N_13578);
nand UO_1667 (O_1667,N_14194,N_14309);
nand UO_1668 (O_1668,N_14058,N_14651);
nor UO_1669 (O_1669,N_14449,N_14540);
or UO_1670 (O_1670,N_14045,N_14861);
nor UO_1671 (O_1671,N_14516,N_14520);
nor UO_1672 (O_1672,N_14742,N_14249);
or UO_1673 (O_1673,N_14103,N_14881);
and UO_1674 (O_1674,N_14273,N_13637);
or UO_1675 (O_1675,N_13938,N_13783);
nor UO_1676 (O_1676,N_13779,N_13659);
nor UO_1677 (O_1677,N_14096,N_14702);
or UO_1678 (O_1678,N_13758,N_14089);
or UO_1679 (O_1679,N_14655,N_14541);
or UO_1680 (O_1680,N_14443,N_14534);
or UO_1681 (O_1681,N_14244,N_14698);
nand UO_1682 (O_1682,N_14689,N_14089);
and UO_1683 (O_1683,N_14419,N_14938);
or UO_1684 (O_1684,N_13568,N_14184);
xor UO_1685 (O_1685,N_14638,N_14530);
nor UO_1686 (O_1686,N_14663,N_14820);
and UO_1687 (O_1687,N_13884,N_14156);
xnor UO_1688 (O_1688,N_13938,N_13852);
or UO_1689 (O_1689,N_13881,N_13864);
and UO_1690 (O_1690,N_13761,N_14787);
nand UO_1691 (O_1691,N_14121,N_14605);
nand UO_1692 (O_1692,N_14736,N_14339);
or UO_1693 (O_1693,N_14665,N_14519);
nand UO_1694 (O_1694,N_14119,N_13909);
and UO_1695 (O_1695,N_14097,N_13625);
nand UO_1696 (O_1696,N_14909,N_13771);
and UO_1697 (O_1697,N_13859,N_14909);
and UO_1698 (O_1698,N_14876,N_14237);
and UO_1699 (O_1699,N_13990,N_14694);
and UO_1700 (O_1700,N_13655,N_14792);
xor UO_1701 (O_1701,N_14959,N_13986);
or UO_1702 (O_1702,N_14388,N_14135);
and UO_1703 (O_1703,N_13973,N_14303);
xor UO_1704 (O_1704,N_14704,N_14689);
and UO_1705 (O_1705,N_14572,N_14763);
and UO_1706 (O_1706,N_13729,N_14714);
xor UO_1707 (O_1707,N_14867,N_14896);
and UO_1708 (O_1708,N_14286,N_14330);
and UO_1709 (O_1709,N_14892,N_14160);
or UO_1710 (O_1710,N_14464,N_14985);
xor UO_1711 (O_1711,N_13713,N_14234);
nor UO_1712 (O_1712,N_14927,N_13669);
or UO_1713 (O_1713,N_13914,N_13980);
and UO_1714 (O_1714,N_14236,N_14980);
or UO_1715 (O_1715,N_14114,N_14080);
or UO_1716 (O_1716,N_14373,N_14104);
nand UO_1717 (O_1717,N_13900,N_13793);
and UO_1718 (O_1718,N_13762,N_13719);
nand UO_1719 (O_1719,N_14419,N_13671);
and UO_1720 (O_1720,N_14732,N_13507);
or UO_1721 (O_1721,N_14843,N_14483);
and UO_1722 (O_1722,N_14970,N_14492);
or UO_1723 (O_1723,N_14859,N_14072);
nor UO_1724 (O_1724,N_13700,N_14785);
nand UO_1725 (O_1725,N_13816,N_14172);
and UO_1726 (O_1726,N_14390,N_14846);
xnor UO_1727 (O_1727,N_14881,N_13939);
nor UO_1728 (O_1728,N_14306,N_14712);
and UO_1729 (O_1729,N_13742,N_14176);
or UO_1730 (O_1730,N_14557,N_14508);
and UO_1731 (O_1731,N_14220,N_13742);
or UO_1732 (O_1732,N_13686,N_14859);
xnor UO_1733 (O_1733,N_14460,N_13868);
nor UO_1734 (O_1734,N_14052,N_14509);
and UO_1735 (O_1735,N_13894,N_13568);
and UO_1736 (O_1736,N_13987,N_14031);
nor UO_1737 (O_1737,N_14421,N_14198);
nand UO_1738 (O_1738,N_14209,N_13874);
and UO_1739 (O_1739,N_13516,N_14622);
and UO_1740 (O_1740,N_13503,N_13515);
or UO_1741 (O_1741,N_13623,N_13678);
or UO_1742 (O_1742,N_14000,N_14175);
nor UO_1743 (O_1743,N_13928,N_14501);
nand UO_1744 (O_1744,N_14482,N_13810);
nand UO_1745 (O_1745,N_14870,N_14210);
nor UO_1746 (O_1746,N_13562,N_14681);
nor UO_1747 (O_1747,N_14309,N_14726);
or UO_1748 (O_1748,N_14964,N_14929);
and UO_1749 (O_1749,N_13898,N_14724);
or UO_1750 (O_1750,N_14406,N_13540);
xor UO_1751 (O_1751,N_14195,N_13757);
nor UO_1752 (O_1752,N_13965,N_14998);
and UO_1753 (O_1753,N_14997,N_13552);
and UO_1754 (O_1754,N_14498,N_13784);
and UO_1755 (O_1755,N_13598,N_14333);
or UO_1756 (O_1756,N_13538,N_13779);
or UO_1757 (O_1757,N_14550,N_14229);
and UO_1758 (O_1758,N_14636,N_13686);
and UO_1759 (O_1759,N_14399,N_13793);
nor UO_1760 (O_1760,N_14815,N_14556);
xnor UO_1761 (O_1761,N_14748,N_14974);
or UO_1762 (O_1762,N_14036,N_14375);
nor UO_1763 (O_1763,N_14579,N_14317);
nand UO_1764 (O_1764,N_13810,N_14414);
nand UO_1765 (O_1765,N_13947,N_13852);
xor UO_1766 (O_1766,N_14298,N_14624);
nor UO_1767 (O_1767,N_14123,N_14582);
nor UO_1768 (O_1768,N_14565,N_13810);
nor UO_1769 (O_1769,N_14966,N_14287);
nand UO_1770 (O_1770,N_13672,N_14068);
nor UO_1771 (O_1771,N_13599,N_14718);
nor UO_1772 (O_1772,N_14276,N_13897);
or UO_1773 (O_1773,N_14460,N_13968);
xnor UO_1774 (O_1774,N_14642,N_14146);
nor UO_1775 (O_1775,N_14635,N_14631);
or UO_1776 (O_1776,N_14472,N_14518);
xor UO_1777 (O_1777,N_14939,N_13954);
nor UO_1778 (O_1778,N_14193,N_14988);
or UO_1779 (O_1779,N_13578,N_14652);
and UO_1780 (O_1780,N_14278,N_14309);
xnor UO_1781 (O_1781,N_14334,N_14303);
xnor UO_1782 (O_1782,N_14296,N_14414);
xor UO_1783 (O_1783,N_14701,N_14285);
nor UO_1784 (O_1784,N_14778,N_13501);
and UO_1785 (O_1785,N_14223,N_14037);
or UO_1786 (O_1786,N_14375,N_14198);
and UO_1787 (O_1787,N_14339,N_13973);
xor UO_1788 (O_1788,N_14455,N_14992);
nand UO_1789 (O_1789,N_13874,N_14917);
xor UO_1790 (O_1790,N_14360,N_14102);
nand UO_1791 (O_1791,N_14064,N_14024);
nor UO_1792 (O_1792,N_13848,N_14988);
or UO_1793 (O_1793,N_14292,N_14852);
or UO_1794 (O_1794,N_13857,N_13971);
nand UO_1795 (O_1795,N_14098,N_14188);
xor UO_1796 (O_1796,N_14861,N_14959);
nor UO_1797 (O_1797,N_13656,N_14170);
nor UO_1798 (O_1798,N_14781,N_14274);
or UO_1799 (O_1799,N_13741,N_14482);
and UO_1800 (O_1800,N_14392,N_14089);
or UO_1801 (O_1801,N_14626,N_13721);
nor UO_1802 (O_1802,N_14131,N_14532);
or UO_1803 (O_1803,N_14547,N_14414);
or UO_1804 (O_1804,N_13951,N_14817);
and UO_1805 (O_1805,N_13628,N_14738);
nor UO_1806 (O_1806,N_14685,N_14127);
xor UO_1807 (O_1807,N_14706,N_14193);
or UO_1808 (O_1808,N_14918,N_14971);
xor UO_1809 (O_1809,N_14211,N_14434);
nor UO_1810 (O_1810,N_13580,N_13654);
xor UO_1811 (O_1811,N_13813,N_14577);
nor UO_1812 (O_1812,N_13678,N_14124);
nand UO_1813 (O_1813,N_13563,N_14373);
nand UO_1814 (O_1814,N_14829,N_14270);
nand UO_1815 (O_1815,N_14955,N_14068);
and UO_1816 (O_1816,N_14486,N_14043);
or UO_1817 (O_1817,N_13633,N_13707);
and UO_1818 (O_1818,N_14036,N_14925);
nand UO_1819 (O_1819,N_14621,N_14829);
nor UO_1820 (O_1820,N_14167,N_14275);
or UO_1821 (O_1821,N_14908,N_13753);
nor UO_1822 (O_1822,N_13586,N_14455);
nor UO_1823 (O_1823,N_14039,N_14680);
nand UO_1824 (O_1824,N_14324,N_14247);
and UO_1825 (O_1825,N_13867,N_13530);
or UO_1826 (O_1826,N_14260,N_13894);
or UO_1827 (O_1827,N_14602,N_14621);
or UO_1828 (O_1828,N_14719,N_14622);
nand UO_1829 (O_1829,N_14473,N_14485);
nor UO_1830 (O_1830,N_13974,N_13901);
xor UO_1831 (O_1831,N_14422,N_14834);
or UO_1832 (O_1832,N_14949,N_13539);
nand UO_1833 (O_1833,N_14125,N_14769);
or UO_1834 (O_1834,N_14863,N_13647);
nor UO_1835 (O_1835,N_14027,N_14162);
and UO_1836 (O_1836,N_14067,N_14518);
nor UO_1837 (O_1837,N_14256,N_14374);
nor UO_1838 (O_1838,N_13564,N_14370);
nor UO_1839 (O_1839,N_13571,N_14576);
nand UO_1840 (O_1840,N_14127,N_14903);
or UO_1841 (O_1841,N_14421,N_13752);
or UO_1842 (O_1842,N_13540,N_14250);
and UO_1843 (O_1843,N_14564,N_14681);
or UO_1844 (O_1844,N_13905,N_13835);
and UO_1845 (O_1845,N_14155,N_13605);
nand UO_1846 (O_1846,N_14003,N_14377);
or UO_1847 (O_1847,N_14533,N_14327);
nor UO_1848 (O_1848,N_13728,N_14700);
and UO_1849 (O_1849,N_14771,N_14322);
nor UO_1850 (O_1850,N_14031,N_13637);
and UO_1851 (O_1851,N_14081,N_14219);
nand UO_1852 (O_1852,N_14287,N_14298);
and UO_1853 (O_1853,N_14788,N_13726);
nor UO_1854 (O_1854,N_13901,N_14760);
nand UO_1855 (O_1855,N_14064,N_14881);
xor UO_1856 (O_1856,N_13506,N_14004);
nor UO_1857 (O_1857,N_14129,N_14723);
or UO_1858 (O_1858,N_14071,N_14335);
or UO_1859 (O_1859,N_14314,N_14838);
nand UO_1860 (O_1860,N_14501,N_13933);
nor UO_1861 (O_1861,N_13584,N_14575);
nor UO_1862 (O_1862,N_14396,N_14922);
or UO_1863 (O_1863,N_14184,N_13683);
and UO_1864 (O_1864,N_14765,N_14516);
or UO_1865 (O_1865,N_13625,N_14306);
nand UO_1866 (O_1866,N_13632,N_14451);
xnor UO_1867 (O_1867,N_14095,N_14596);
nand UO_1868 (O_1868,N_14011,N_14237);
and UO_1869 (O_1869,N_14892,N_14601);
and UO_1870 (O_1870,N_13901,N_14670);
and UO_1871 (O_1871,N_13936,N_14609);
nand UO_1872 (O_1872,N_14684,N_14811);
nand UO_1873 (O_1873,N_14769,N_13738);
nor UO_1874 (O_1874,N_14296,N_14214);
and UO_1875 (O_1875,N_14132,N_14682);
nor UO_1876 (O_1876,N_13712,N_14243);
nand UO_1877 (O_1877,N_14337,N_13524);
nor UO_1878 (O_1878,N_14837,N_14198);
nand UO_1879 (O_1879,N_14487,N_13726);
and UO_1880 (O_1880,N_14008,N_13940);
and UO_1881 (O_1881,N_13605,N_14994);
nor UO_1882 (O_1882,N_14372,N_14063);
or UO_1883 (O_1883,N_14724,N_14436);
nor UO_1884 (O_1884,N_14914,N_13680);
xnor UO_1885 (O_1885,N_13666,N_13964);
and UO_1886 (O_1886,N_14057,N_13659);
and UO_1887 (O_1887,N_14895,N_14999);
nor UO_1888 (O_1888,N_14211,N_13706);
and UO_1889 (O_1889,N_14818,N_13761);
nand UO_1890 (O_1890,N_13733,N_13881);
or UO_1891 (O_1891,N_14588,N_14689);
xor UO_1892 (O_1892,N_14065,N_14865);
nor UO_1893 (O_1893,N_13603,N_14924);
or UO_1894 (O_1894,N_14503,N_14153);
nor UO_1895 (O_1895,N_14552,N_14290);
and UO_1896 (O_1896,N_13873,N_14583);
or UO_1897 (O_1897,N_13793,N_14819);
nor UO_1898 (O_1898,N_13797,N_14551);
nand UO_1899 (O_1899,N_14241,N_13837);
and UO_1900 (O_1900,N_14613,N_13548);
nor UO_1901 (O_1901,N_13593,N_14422);
or UO_1902 (O_1902,N_14422,N_13851);
or UO_1903 (O_1903,N_14224,N_14492);
or UO_1904 (O_1904,N_14200,N_13924);
nor UO_1905 (O_1905,N_14574,N_14174);
nand UO_1906 (O_1906,N_13578,N_14629);
nor UO_1907 (O_1907,N_14038,N_14919);
or UO_1908 (O_1908,N_14047,N_14457);
nand UO_1909 (O_1909,N_14021,N_14705);
nor UO_1910 (O_1910,N_13612,N_14606);
xor UO_1911 (O_1911,N_13542,N_13822);
xnor UO_1912 (O_1912,N_14592,N_14952);
and UO_1913 (O_1913,N_14903,N_13797);
nor UO_1914 (O_1914,N_13859,N_13996);
xnor UO_1915 (O_1915,N_13913,N_13709);
and UO_1916 (O_1916,N_14748,N_14653);
or UO_1917 (O_1917,N_13763,N_13952);
or UO_1918 (O_1918,N_13871,N_14101);
nand UO_1919 (O_1919,N_14567,N_13811);
and UO_1920 (O_1920,N_14293,N_14501);
and UO_1921 (O_1921,N_13789,N_14987);
and UO_1922 (O_1922,N_13718,N_14250);
and UO_1923 (O_1923,N_14225,N_14947);
nor UO_1924 (O_1924,N_14860,N_14485);
nand UO_1925 (O_1925,N_14007,N_14154);
and UO_1926 (O_1926,N_14254,N_14344);
or UO_1927 (O_1927,N_14594,N_14417);
nor UO_1928 (O_1928,N_13510,N_14545);
nand UO_1929 (O_1929,N_14531,N_14128);
xnor UO_1930 (O_1930,N_14867,N_13843);
and UO_1931 (O_1931,N_14213,N_13510);
nor UO_1932 (O_1932,N_14454,N_14421);
nor UO_1933 (O_1933,N_13617,N_13880);
or UO_1934 (O_1934,N_13526,N_13733);
nand UO_1935 (O_1935,N_14825,N_14066);
or UO_1936 (O_1936,N_14213,N_14904);
nor UO_1937 (O_1937,N_14751,N_14438);
nor UO_1938 (O_1938,N_14449,N_14542);
or UO_1939 (O_1939,N_14837,N_14653);
xor UO_1940 (O_1940,N_14469,N_13685);
and UO_1941 (O_1941,N_13848,N_14990);
xnor UO_1942 (O_1942,N_13694,N_14116);
xnor UO_1943 (O_1943,N_14194,N_14491);
and UO_1944 (O_1944,N_14267,N_13816);
or UO_1945 (O_1945,N_14159,N_13599);
and UO_1946 (O_1946,N_14117,N_14581);
and UO_1947 (O_1947,N_14212,N_13875);
nor UO_1948 (O_1948,N_14897,N_13729);
nor UO_1949 (O_1949,N_14905,N_13772);
or UO_1950 (O_1950,N_13773,N_14641);
nor UO_1951 (O_1951,N_14280,N_14922);
nand UO_1952 (O_1952,N_13534,N_14500);
nand UO_1953 (O_1953,N_14319,N_13998);
nand UO_1954 (O_1954,N_13552,N_13758);
or UO_1955 (O_1955,N_13681,N_14056);
and UO_1956 (O_1956,N_14577,N_14735);
or UO_1957 (O_1957,N_14042,N_14034);
or UO_1958 (O_1958,N_13591,N_14576);
nand UO_1959 (O_1959,N_14496,N_14421);
nand UO_1960 (O_1960,N_14882,N_13614);
nor UO_1961 (O_1961,N_13757,N_14751);
nor UO_1962 (O_1962,N_14587,N_14517);
or UO_1963 (O_1963,N_13823,N_14186);
or UO_1964 (O_1964,N_13604,N_13722);
or UO_1965 (O_1965,N_14899,N_14487);
and UO_1966 (O_1966,N_14094,N_13978);
xnor UO_1967 (O_1967,N_14836,N_14852);
xor UO_1968 (O_1968,N_14381,N_14762);
or UO_1969 (O_1969,N_13603,N_13539);
or UO_1970 (O_1970,N_13953,N_14843);
nand UO_1971 (O_1971,N_14737,N_14003);
or UO_1972 (O_1972,N_13775,N_14876);
xor UO_1973 (O_1973,N_13935,N_14120);
nor UO_1974 (O_1974,N_13776,N_14490);
or UO_1975 (O_1975,N_14053,N_14873);
nand UO_1976 (O_1976,N_14537,N_14411);
nor UO_1977 (O_1977,N_14941,N_13994);
nor UO_1978 (O_1978,N_14815,N_13824);
and UO_1979 (O_1979,N_14076,N_13811);
or UO_1980 (O_1980,N_14962,N_14835);
nand UO_1981 (O_1981,N_13746,N_14027);
nor UO_1982 (O_1982,N_14376,N_14466);
or UO_1983 (O_1983,N_14074,N_13678);
xnor UO_1984 (O_1984,N_14050,N_14609);
nor UO_1985 (O_1985,N_13945,N_14192);
or UO_1986 (O_1986,N_14578,N_14182);
or UO_1987 (O_1987,N_13579,N_14945);
xnor UO_1988 (O_1988,N_13718,N_13935);
nor UO_1989 (O_1989,N_13816,N_14388);
nor UO_1990 (O_1990,N_14239,N_13983);
and UO_1991 (O_1991,N_14675,N_13537);
nand UO_1992 (O_1992,N_13644,N_14458);
and UO_1993 (O_1993,N_13737,N_13574);
nor UO_1994 (O_1994,N_14900,N_14624);
nand UO_1995 (O_1995,N_14998,N_14445);
nor UO_1996 (O_1996,N_13719,N_14231);
or UO_1997 (O_1997,N_14312,N_14917);
nand UO_1998 (O_1998,N_14781,N_13731);
and UO_1999 (O_1999,N_14891,N_13684);
endmodule