module basic_1000_10000_1500_10_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_568,In_222);
or U1 (N_1,In_697,In_225);
xor U2 (N_2,In_48,In_761);
and U3 (N_3,In_352,In_724);
nand U4 (N_4,In_117,In_994);
and U5 (N_5,In_688,In_919);
or U6 (N_6,In_247,In_323);
or U7 (N_7,In_634,In_39);
or U8 (N_8,In_715,In_576);
or U9 (N_9,In_740,In_844);
nor U10 (N_10,In_194,In_252);
or U11 (N_11,In_760,In_596);
or U12 (N_12,In_971,In_89);
nand U13 (N_13,In_903,In_192);
or U14 (N_14,In_402,In_917);
nor U15 (N_15,In_977,In_446);
nand U16 (N_16,In_622,In_597);
and U17 (N_17,In_215,In_338);
nand U18 (N_18,In_613,In_214);
nand U19 (N_19,In_379,In_17);
and U20 (N_20,In_506,In_423);
and U21 (N_21,In_610,In_955);
and U22 (N_22,In_502,In_793);
nand U23 (N_23,In_242,In_435);
or U24 (N_24,In_546,In_282);
xnor U25 (N_25,In_186,In_53);
and U26 (N_26,In_381,In_751);
nand U27 (N_27,In_561,In_907);
nor U28 (N_28,In_40,In_463);
nor U29 (N_29,In_654,In_738);
nor U30 (N_30,In_968,In_881);
and U31 (N_31,In_636,In_816);
nor U32 (N_32,In_768,In_120);
nor U33 (N_33,In_615,In_23);
and U34 (N_34,In_393,In_839);
nand U35 (N_35,In_863,In_46);
nor U36 (N_36,In_771,In_900);
or U37 (N_37,In_341,In_467);
or U38 (N_38,In_468,In_679);
nor U39 (N_39,In_79,In_555);
or U40 (N_40,In_948,In_535);
nand U41 (N_41,In_623,In_21);
nor U42 (N_42,In_814,In_890);
nor U43 (N_43,In_50,In_44);
nand U44 (N_44,In_963,In_314);
nor U45 (N_45,In_197,In_587);
and U46 (N_46,In_95,In_429);
nor U47 (N_47,In_820,In_267);
and U48 (N_48,In_929,In_922);
nor U49 (N_49,In_982,In_200);
nand U50 (N_50,In_389,In_359);
and U51 (N_51,In_794,In_664);
and U52 (N_52,In_360,In_81);
or U53 (N_53,In_918,In_706);
nor U54 (N_54,In_933,In_873);
xnor U55 (N_55,In_43,In_415);
nor U56 (N_56,In_280,In_572);
nor U57 (N_57,In_908,In_265);
or U58 (N_58,In_791,In_744);
nand U59 (N_59,In_151,In_749);
nor U60 (N_60,In_297,In_251);
nor U61 (N_61,In_902,In_16);
and U62 (N_62,In_975,In_210);
nand U63 (N_63,In_951,In_727);
nor U64 (N_64,In_388,In_722);
or U65 (N_65,In_20,In_399);
nand U66 (N_66,In_512,In_603);
xnor U67 (N_67,In_403,In_625);
or U68 (N_68,In_148,In_6);
and U69 (N_69,In_520,In_133);
nand U70 (N_70,In_471,In_432);
and U71 (N_71,In_608,In_363);
nor U72 (N_72,In_111,In_51);
nand U73 (N_73,In_992,In_822);
and U74 (N_74,In_418,In_209);
nor U75 (N_75,In_556,In_583);
and U76 (N_76,In_894,In_702);
nor U77 (N_77,In_147,In_327);
or U78 (N_78,In_876,In_776);
xnor U79 (N_79,In_213,In_125);
and U80 (N_80,In_538,In_686);
and U81 (N_81,In_217,In_725);
nor U82 (N_82,In_377,In_859);
nand U83 (N_83,In_532,In_315);
nor U84 (N_84,In_369,In_368);
nand U85 (N_85,In_316,In_885);
or U86 (N_86,In_266,In_788);
and U87 (N_87,In_499,In_806);
nor U88 (N_88,In_159,In_362);
nor U89 (N_89,In_650,In_15);
nand U90 (N_90,In_443,In_481);
nor U91 (N_91,In_144,In_166);
nand U92 (N_92,In_414,In_237);
and U93 (N_93,In_705,In_105);
nor U94 (N_94,In_807,In_519);
nand U95 (N_95,In_272,In_123);
and U96 (N_96,In_748,In_921);
xor U97 (N_97,In_784,In_943);
xnor U98 (N_98,In_993,In_978);
nor U99 (N_99,In_387,In_726);
nor U100 (N_100,In_464,In_714);
nor U101 (N_101,In_590,In_938);
or U102 (N_102,In_313,In_182);
nand U103 (N_103,In_54,In_234);
or U104 (N_104,In_452,In_457);
nand U105 (N_105,In_884,In_490);
or U106 (N_106,In_841,In_243);
and U107 (N_107,In_823,In_661);
or U108 (N_108,In_757,In_137);
or U109 (N_109,In_756,In_284);
nor U110 (N_110,In_762,In_665);
nand U111 (N_111,In_212,In_495);
or U112 (N_112,In_719,In_301);
or U113 (N_113,In_484,In_766);
nor U114 (N_114,In_527,In_798);
xnor U115 (N_115,In_947,In_537);
nor U116 (N_116,In_472,In_515);
nand U117 (N_117,In_255,In_276);
and U118 (N_118,In_68,In_383);
nand U119 (N_119,In_351,In_801);
and U120 (N_120,In_828,In_101);
xor U121 (N_121,In_263,In_513);
or U122 (N_122,In_674,In_303);
and U123 (N_123,In_451,In_602);
and U124 (N_124,In_773,In_343);
nor U125 (N_125,In_775,In_239);
and U126 (N_126,In_398,In_504);
nand U127 (N_127,In_183,In_509);
nand U128 (N_128,In_616,In_617);
or U129 (N_129,In_819,In_106);
nand U130 (N_130,In_643,In_781);
and U131 (N_131,In_96,In_962);
and U132 (N_132,In_211,In_118);
nand U133 (N_133,In_928,In_796);
nor U134 (N_134,In_447,In_685);
nand U135 (N_135,In_420,In_638);
nor U136 (N_136,In_18,In_808);
or U137 (N_137,In_114,In_476);
and U138 (N_138,In_861,In_789);
xnor U139 (N_139,In_256,In_904);
or U140 (N_140,In_168,In_345);
and U141 (N_141,In_618,In_244);
or U142 (N_142,In_969,In_677);
or U143 (N_143,In_678,In_462);
nor U144 (N_144,In_895,In_75);
or U145 (N_145,In_205,In_246);
nand U146 (N_146,In_826,In_669);
nor U147 (N_147,In_136,In_708);
nand U148 (N_148,In_397,In_132);
xor U149 (N_149,In_530,In_245);
xnor U150 (N_150,In_812,In_455);
nor U151 (N_151,In_219,In_356);
nor U152 (N_152,In_914,In_346);
and U153 (N_153,In_645,In_827);
nor U154 (N_154,In_286,In_510);
nor U155 (N_155,In_162,In_175);
nand U156 (N_156,In_199,In_989);
nor U157 (N_157,In_391,In_845);
and U158 (N_158,In_439,In_64);
and U159 (N_159,In_26,In_283);
xor U160 (N_160,In_547,In_410);
and U161 (N_161,In_134,In_772);
or U162 (N_162,In_931,In_730);
or U163 (N_163,In_41,In_913);
nand U164 (N_164,In_795,In_121);
nor U165 (N_165,In_142,In_38);
or U166 (N_166,In_747,In_552);
or U167 (N_167,In_655,In_642);
nor U168 (N_168,In_87,In_325);
nor U169 (N_169,In_293,In_470);
nor U170 (N_170,In_573,In_474);
or U171 (N_171,In_701,In_396);
nand U172 (N_172,In_171,In_30);
nand U173 (N_173,In_713,In_690);
xor U174 (N_174,In_337,In_56);
nor U175 (N_175,In_249,In_326);
or U176 (N_176,In_201,In_566);
nand U177 (N_177,In_767,In_32);
and U178 (N_178,In_544,In_723);
nor U179 (N_179,In_563,In_191);
nor U180 (N_180,In_743,In_551);
or U181 (N_181,In_334,In_478);
xor U182 (N_182,In_940,In_459);
and U183 (N_183,In_187,In_868);
and U184 (N_184,In_763,In_196);
nand U185 (N_185,In_952,In_299);
nor U186 (N_186,In_970,In_324);
or U187 (N_187,In_640,In_503);
xnor U188 (N_188,In_434,In_296);
or U189 (N_189,In_840,In_516);
nand U190 (N_190,In_736,In_318);
nor U191 (N_191,In_739,In_250);
or U192 (N_192,In_945,In_545);
nand U193 (N_193,In_371,In_233);
nor U194 (N_194,In_90,In_8);
and U195 (N_195,In_311,In_534);
or U196 (N_196,In_208,In_291);
or U197 (N_197,In_69,In_995);
nor U198 (N_198,In_99,In_139);
or U199 (N_199,In_865,In_979);
and U200 (N_200,In_58,In_601);
and U201 (N_201,In_290,In_554);
nand U202 (N_202,In_92,In_699);
or U203 (N_203,In_711,In_73);
nand U204 (N_204,In_382,In_899);
xor U205 (N_205,In_526,In_817);
nor U206 (N_206,In_12,In_925);
nor U207 (N_207,In_855,In_731);
nor U208 (N_208,In_611,In_335);
or U209 (N_209,In_100,In_430);
nand U210 (N_210,In_492,In_891);
nor U211 (N_211,In_305,In_878);
and U212 (N_212,In_658,In_445);
and U213 (N_213,In_80,In_720);
xor U214 (N_214,In_689,In_501);
or U215 (N_215,In_486,In_864);
nor U216 (N_216,In_231,In_70);
nor U217 (N_217,In_366,In_539);
nand U218 (N_218,In_433,In_924);
or U219 (N_219,In_307,In_769);
nand U220 (N_220,In_941,In_949);
and U221 (N_221,In_164,In_442);
or U222 (N_222,In_787,In_646);
nor U223 (N_223,In_600,In_893);
nand U224 (N_224,In_564,In_167);
nor U225 (N_225,In_329,In_934);
nor U226 (N_226,In_858,In_72);
xor U227 (N_227,In_479,In_936);
nand U228 (N_228,In_440,In_27);
and U229 (N_229,In_660,In_112);
xor U230 (N_230,In_718,In_764);
nor U231 (N_231,In_851,In_47);
nor U232 (N_232,In_74,In_797);
nand U233 (N_233,In_274,In_942);
nor U234 (N_234,In_332,In_695);
or U235 (N_235,In_946,In_635);
and U236 (N_236,In_514,In_227);
nand U237 (N_237,In_422,In_392);
nor U238 (N_238,In_540,In_927);
or U239 (N_239,In_473,In_427);
nand U240 (N_240,In_444,In_224);
nand U241 (N_241,In_548,In_852);
and U242 (N_242,In_523,In_721);
or U243 (N_243,In_333,In_77);
and U244 (N_244,In_588,In_872);
xnor U245 (N_245,In_649,In_687);
nor U246 (N_246,In_803,In_61);
nand U247 (N_247,In_581,In_999);
or U248 (N_248,In_83,In_24);
and U249 (N_249,In_298,In_684);
or U250 (N_250,In_113,In_958);
or U251 (N_251,In_582,In_683);
nand U252 (N_252,In_939,In_277);
and U253 (N_253,In_657,In_521);
nor U254 (N_254,In_441,In_838);
or U255 (N_255,In_785,In_857);
and U256 (N_256,In_384,In_469);
or U257 (N_257,In_138,In_836);
nor U258 (N_258,In_579,In_831);
and U259 (N_259,In_889,In_169);
or U260 (N_260,In_179,In_742);
or U261 (N_261,In_408,In_577);
nor U262 (N_262,In_883,In_498);
and U263 (N_263,In_511,In_892);
nand U264 (N_264,In_854,In_569);
nand U265 (N_265,In_153,In_9);
xnor U266 (N_266,In_631,In_830);
or U267 (N_267,In_322,In_374);
nand U268 (N_268,In_52,In_825);
nor U269 (N_269,In_104,In_593);
nor U270 (N_270,In_604,In_198);
or U271 (N_271,In_524,In_10);
nand U272 (N_272,In_364,In_328);
or U273 (N_273,In_984,In_753);
or U274 (N_274,In_436,In_912);
and U275 (N_275,In_656,In_370);
nor U276 (N_276,In_570,In_230);
nand U277 (N_277,In_270,In_480);
and U278 (N_278,In_84,In_620);
nor U279 (N_279,In_732,In_957);
nor U280 (N_280,In_110,In_965);
and U281 (N_281,In_361,In_578);
or U282 (N_282,In_632,In_416);
nand U283 (N_283,In_652,In_3);
and U284 (N_284,In_140,In_254);
xnor U285 (N_285,In_754,In_562);
or U286 (N_286,In_536,In_188);
and U287 (N_287,In_639,In_347);
or U288 (N_288,In_853,In_671);
nand U289 (N_289,In_496,In_216);
nor U290 (N_290,In_97,In_1);
nor U291 (N_291,In_232,In_896);
nand U292 (N_292,In_517,In_240);
or U293 (N_293,In_765,In_960);
or U294 (N_294,In_413,In_189);
nand U295 (N_295,In_135,In_466);
xnor U296 (N_296,In_355,In_107);
and U297 (N_297,In_783,In_897);
nor U298 (N_298,In_983,In_707);
nand U299 (N_299,In_165,In_7);
or U300 (N_300,In_150,In_505);
nand U301 (N_301,In_614,In_867);
or U302 (N_302,In_82,In_609);
nor U303 (N_303,In_915,In_281);
and U304 (N_304,In_986,In_28);
nand U305 (N_305,In_241,In_580);
or U306 (N_306,In_882,In_847);
nand U307 (N_307,In_950,In_449);
nor U308 (N_308,In_595,In_228);
and U309 (N_309,In_628,In_287);
xnor U310 (N_310,In_585,In_629);
or U311 (N_311,In_354,In_586);
or U312 (N_312,In_717,In_170);
or U313 (N_313,In_821,In_86);
nand U314 (N_314,In_729,In_932);
nor U315 (N_315,In_62,In_380);
or U316 (N_316,In_833,In_849);
nand U317 (N_317,In_980,In_181);
nand U318 (N_318,In_497,In_437);
and U319 (N_319,In_626,In_734);
and U320 (N_320,In_592,In_676);
nor U321 (N_321,In_42,In_531);
and U322 (N_322,In_944,In_605);
and U323 (N_323,In_911,In_935);
nor U324 (N_324,In_888,In_152);
and U325 (N_325,In_786,In_115);
xor U326 (N_326,In_312,In_483);
xor U327 (N_327,In_220,In_348);
and U328 (N_328,In_195,In_782);
nor U329 (N_329,In_874,In_559);
xnor U330 (N_330,In_741,In_494);
nor U331 (N_331,In_320,In_996);
nand U332 (N_332,In_953,In_612);
nand U333 (N_333,In_647,In_458);
or U334 (N_334,In_920,In_594);
and U335 (N_335,In_964,In_353);
nand U336 (N_336,In_336,In_342);
or U337 (N_337,In_550,In_759);
and U338 (N_338,In_589,In_712);
nand U339 (N_339,In_367,In_755);
or U340 (N_340,In_160,In_302);
nor U341 (N_341,In_163,In_800);
nand U342 (N_342,In_930,In_257);
or U343 (N_343,In_675,In_223);
nand U344 (N_344,In_295,In_401);
or U345 (N_345,In_633,In_973);
and U346 (N_346,In_130,In_461);
nor U347 (N_347,In_651,In_76);
or U348 (N_348,In_818,In_119);
or U349 (N_349,In_906,In_704);
nand U350 (N_350,In_485,In_78);
nor U351 (N_351,In_155,In_176);
nand U352 (N_352,In_365,In_507);
nand U353 (N_353,In_268,In_644);
nand U354 (N_354,In_275,In_752);
nand U355 (N_355,In_967,In_571);
nor U356 (N_356,In_774,In_682);
nand U357 (N_357,In_238,In_35);
and U358 (N_358,In_630,In_694);
nor U359 (N_359,In_407,In_696);
or U360 (N_360,In_428,In_22);
nor U361 (N_361,In_584,In_394);
or U362 (N_362,In_288,In_832);
nand U363 (N_363,In_558,In_116);
and U364 (N_364,In_218,In_835);
nand U365 (N_365,In_131,In_278);
nor U366 (N_366,In_799,In_491);
nand U367 (N_367,In_66,In_508);
nor U368 (N_368,In_733,In_606);
and U369 (N_369,In_319,In_489);
nor U370 (N_370,In_438,In_770);
or U371 (N_371,In_203,In_465);
xor U372 (N_372,In_149,In_659);
or U373 (N_373,In_59,In_190);
nor U374 (N_374,In_412,In_745);
or U375 (N_375,In_4,In_681);
nand U376 (N_376,In_518,In_529);
and U377 (N_377,In_161,In_780);
or U378 (N_378,In_236,In_567);
xor U379 (N_379,In_488,In_691);
nand U380 (N_380,In_259,In_905);
xnor U381 (N_381,In_703,In_177);
and U382 (N_382,In_901,In_372);
and U383 (N_383,In_487,In_350);
nor U384 (N_384,In_271,In_395);
nor U385 (N_385,In_456,In_842);
nand U386 (N_386,In_289,In_937);
nand U387 (N_387,In_25,In_103);
nand U388 (N_388,In_339,In_321);
nor U389 (N_389,In_829,In_94);
nor U390 (N_390,In_627,In_49);
nand U391 (N_391,In_425,In_998);
nand U392 (N_392,In_98,In_709);
and U393 (N_393,In_248,In_11);
nor U394 (N_394,In_837,In_141);
and U395 (N_395,In_624,In_285);
nor U396 (N_396,In_304,In_431);
nand U397 (N_397,In_981,In_790);
or U398 (N_398,In_460,In_972);
nand U399 (N_399,In_127,In_405);
or U400 (N_400,In_746,In_5);
nor U401 (N_401,In_128,In_990);
nand U402 (N_402,In_693,In_376);
or U403 (N_403,In_331,In_813);
nor U404 (N_404,In_173,In_976);
nand U405 (N_405,In_373,In_330);
and U406 (N_406,In_65,In_31);
and U407 (N_407,In_777,In_923);
xor U408 (N_408,In_549,In_317);
nand U409 (N_409,In_543,In_154);
xor U410 (N_410,In_871,In_204);
nor U411 (N_411,In_804,In_126);
nor U412 (N_412,In_988,In_528);
nor U413 (N_413,In_260,In_802);
or U414 (N_414,In_680,In_88);
or U415 (N_415,In_273,In_178);
and U416 (N_416,In_560,In_557);
or U417 (N_417,In_124,In_292);
nand U418 (N_418,In_926,In_898);
nand U419 (N_419,In_641,In_673);
or U420 (N_420,In_700,In_426);
or U421 (N_421,In_565,In_843);
nand U422 (N_422,In_869,In_916);
nor U423 (N_423,In_668,In_985);
or U424 (N_424,In_834,In_279);
nor U425 (N_425,In_129,In_55);
or U426 (N_426,In_109,In_310);
nand U427 (N_427,In_146,In_991);
nand U428 (N_428,In_824,In_666);
and U429 (N_429,In_409,In_909);
or U430 (N_430,In_974,In_886);
nand U431 (N_431,In_60,In_598);
nor U432 (N_432,In_959,In_344);
nor U433 (N_433,In_987,In_961);
or U434 (N_434,In_728,In_454);
nor U435 (N_435,In_340,In_14);
and U436 (N_436,In_261,In_19);
nand U437 (N_437,In_758,In_648);
nor U438 (N_438,In_525,In_406);
nand U439 (N_439,In_357,In_663);
or U440 (N_440,In_156,In_294);
or U441 (N_441,In_621,In_37);
nor U442 (N_442,In_997,In_856);
nand U443 (N_443,In_180,In_493);
and U444 (N_444,In_93,In_235);
nand U445 (N_445,In_887,In_848);
and U446 (N_446,In_229,In_378);
and U447 (N_447,In_448,In_419);
and U448 (N_448,In_862,In_145);
or U449 (N_449,In_33,In_522);
or U450 (N_450,In_450,In_866);
and U451 (N_451,In_306,In_309);
nor U452 (N_452,In_750,In_108);
xor U453 (N_453,In_102,In_34);
and U454 (N_454,In_637,In_390);
nand U455 (N_455,In_846,In_36);
nand U456 (N_456,In_143,In_157);
nor U457 (N_457,In_475,In_850);
xor U458 (N_458,In_253,In_185);
nand U459 (N_459,In_533,In_349);
nor U460 (N_460,In_2,In_29);
or U461 (N_461,In_158,In_85);
or U462 (N_462,In_122,In_63);
nor U463 (N_463,In_477,In_956);
nand U464 (N_464,In_662,In_880);
nand U465 (N_465,In_716,In_910);
or U466 (N_466,In_174,In_778);
and U467 (N_467,In_400,In_553);
nand U468 (N_468,In_207,In_879);
nor U469 (N_469,In_453,In_184);
or U470 (N_470,In_667,In_67);
and U471 (N_471,In_591,In_811);
nand U472 (N_472,In_411,In_779);
nand U473 (N_473,In_206,In_308);
or U474 (N_474,In_877,In_172);
nand U475 (N_475,In_202,In_599);
and U476 (N_476,In_264,In_870);
and U477 (N_477,In_385,In_672);
or U478 (N_478,In_735,In_193);
and U479 (N_479,In_860,In_221);
or U480 (N_480,In_358,In_421);
nand U481 (N_481,In_424,In_875);
nor U482 (N_482,In_809,In_574);
or U483 (N_483,In_262,In_619);
or U484 (N_484,In_13,In_482);
and U485 (N_485,In_0,In_670);
and U486 (N_486,In_710,In_269);
or U487 (N_487,In_575,In_698);
and U488 (N_488,In_386,In_500);
xnor U489 (N_489,In_815,In_417);
nor U490 (N_490,In_404,In_91);
nand U491 (N_491,In_45,In_57);
and U492 (N_492,In_737,In_226);
nor U493 (N_493,In_541,In_966);
nand U494 (N_494,In_71,In_954);
or U495 (N_495,In_692,In_607);
nand U496 (N_496,In_792,In_258);
and U497 (N_497,In_300,In_653);
or U498 (N_498,In_542,In_805);
or U499 (N_499,In_810,In_375);
nand U500 (N_500,In_176,In_974);
and U501 (N_501,In_383,In_441);
nand U502 (N_502,In_380,In_478);
xor U503 (N_503,In_844,In_560);
nand U504 (N_504,In_65,In_481);
and U505 (N_505,In_923,In_45);
and U506 (N_506,In_779,In_574);
or U507 (N_507,In_474,In_425);
nor U508 (N_508,In_951,In_159);
nor U509 (N_509,In_462,In_986);
or U510 (N_510,In_360,In_671);
or U511 (N_511,In_5,In_744);
and U512 (N_512,In_509,In_444);
nor U513 (N_513,In_716,In_997);
and U514 (N_514,In_710,In_597);
and U515 (N_515,In_167,In_217);
or U516 (N_516,In_495,In_243);
nor U517 (N_517,In_717,In_129);
nor U518 (N_518,In_186,In_116);
xor U519 (N_519,In_778,In_607);
nand U520 (N_520,In_524,In_212);
nand U521 (N_521,In_346,In_577);
nand U522 (N_522,In_183,In_637);
xor U523 (N_523,In_782,In_344);
nor U524 (N_524,In_661,In_163);
or U525 (N_525,In_574,In_913);
or U526 (N_526,In_705,In_121);
and U527 (N_527,In_353,In_454);
nand U528 (N_528,In_124,In_62);
nand U529 (N_529,In_738,In_599);
nor U530 (N_530,In_662,In_132);
and U531 (N_531,In_918,In_593);
and U532 (N_532,In_838,In_978);
or U533 (N_533,In_354,In_536);
or U534 (N_534,In_158,In_460);
nand U535 (N_535,In_194,In_165);
nand U536 (N_536,In_421,In_266);
and U537 (N_537,In_31,In_143);
nor U538 (N_538,In_806,In_416);
or U539 (N_539,In_434,In_606);
nand U540 (N_540,In_774,In_58);
nand U541 (N_541,In_360,In_421);
nor U542 (N_542,In_597,In_843);
or U543 (N_543,In_465,In_898);
nor U544 (N_544,In_58,In_462);
nand U545 (N_545,In_814,In_60);
xnor U546 (N_546,In_812,In_552);
and U547 (N_547,In_983,In_951);
or U548 (N_548,In_201,In_269);
and U549 (N_549,In_746,In_136);
nand U550 (N_550,In_655,In_746);
nand U551 (N_551,In_356,In_484);
nand U552 (N_552,In_735,In_74);
or U553 (N_553,In_881,In_402);
or U554 (N_554,In_604,In_998);
or U555 (N_555,In_950,In_505);
or U556 (N_556,In_375,In_724);
xnor U557 (N_557,In_988,In_396);
and U558 (N_558,In_873,In_277);
nor U559 (N_559,In_4,In_65);
and U560 (N_560,In_107,In_624);
and U561 (N_561,In_559,In_111);
or U562 (N_562,In_327,In_200);
nor U563 (N_563,In_729,In_803);
nand U564 (N_564,In_720,In_360);
nor U565 (N_565,In_212,In_33);
nand U566 (N_566,In_509,In_904);
nor U567 (N_567,In_559,In_870);
or U568 (N_568,In_916,In_393);
or U569 (N_569,In_548,In_305);
and U570 (N_570,In_512,In_371);
or U571 (N_571,In_579,In_589);
nor U572 (N_572,In_462,In_663);
nand U573 (N_573,In_32,In_753);
nor U574 (N_574,In_229,In_524);
nor U575 (N_575,In_113,In_434);
nand U576 (N_576,In_254,In_582);
nor U577 (N_577,In_578,In_509);
nand U578 (N_578,In_216,In_678);
nand U579 (N_579,In_140,In_779);
and U580 (N_580,In_868,In_815);
or U581 (N_581,In_325,In_960);
nor U582 (N_582,In_363,In_419);
nand U583 (N_583,In_690,In_397);
and U584 (N_584,In_974,In_796);
or U585 (N_585,In_316,In_4);
nand U586 (N_586,In_109,In_510);
nand U587 (N_587,In_795,In_858);
nand U588 (N_588,In_390,In_712);
nand U589 (N_589,In_635,In_122);
nor U590 (N_590,In_287,In_178);
and U591 (N_591,In_303,In_38);
nor U592 (N_592,In_500,In_23);
nand U593 (N_593,In_244,In_25);
nor U594 (N_594,In_199,In_686);
nor U595 (N_595,In_953,In_908);
and U596 (N_596,In_455,In_267);
and U597 (N_597,In_343,In_769);
nand U598 (N_598,In_642,In_353);
xor U599 (N_599,In_398,In_522);
nand U600 (N_600,In_528,In_307);
nor U601 (N_601,In_552,In_18);
nand U602 (N_602,In_388,In_159);
or U603 (N_603,In_390,In_864);
or U604 (N_604,In_880,In_450);
nor U605 (N_605,In_236,In_561);
and U606 (N_606,In_867,In_793);
nand U607 (N_607,In_372,In_61);
or U608 (N_608,In_871,In_742);
and U609 (N_609,In_279,In_300);
xor U610 (N_610,In_561,In_862);
or U611 (N_611,In_397,In_944);
nor U612 (N_612,In_133,In_365);
and U613 (N_613,In_447,In_876);
and U614 (N_614,In_383,In_220);
or U615 (N_615,In_617,In_17);
nand U616 (N_616,In_203,In_347);
nor U617 (N_617,In_837,In_316);
xnor U618 (N_618,In_787,In_120);
or U619 (N_619,In_512,In_915);
or U620 (N_620,In_312,In_698);
and U621 (N_621,In_123,In_339);
nor U622 (N_622,In_221,In_849);
nor U623 (N_623,In_817,In_897);
xor U624 (N_624,In_653,In_46);
and U625 (N_625,In_275,In_596);
nand U626 (N_626,In_548,In_779);
xor U627 (N_627,In_585,In_86);
or U628 (N_628,In_588,In_658);
and U629 (N_629,In_631,In_35);
and U630 (N_630,In_915,In_982);
or U631 (N_631,In_801,In_995);
and U632 (N_632,In_698,In_221);
nand U633 (N_633,In_227,In_381);
xor U634 (N_634,In_410,In_143);
nand U635 (N_635,In_217,In_246);
nand U636 (N_636,In_44,In_401);
nand U637 (N_637,In_37,In_629);
nand U638 (N_638,In_538,In_522);
and U639 (N_639,In_337,In_55);
or U640 (N_640,In_812,In_243);
nor U641 (N_641,In_618,In_304);
nand U642 (N_642,In_35,In_440);
or U643 (N_643,In_22,In_769);
or U644 (N_644,In_852,In_570);
nand U645 (N_645,In_327,In_543);
nand U646 (N_646,In_842,In_914);
nor U647 (N_647,In_596,In_934);
nand U648 (N_648,In_239,In_704);
xnor U649 (N_649,In_453,In_470);
nor U650 (N_650,In_92,In_232);
or U651 (N_651,In_944,In_259);
nand U652 (N_652,In_859,In_821);
or U653 (N_653,In_366,In_321);
nand U654 (N_654,In_778,In_180);
nor U655 (N_655,In_35,In_158);
nand U656 (N_656,In_242,In_62);
xnor U657 (N_657,In_397,In_40);
and U658 (N_658,In_58,In_307);
nand U659 (N_659,In_817,In_756);
nand U660 (N_660,In_351,In_436);
or U661 (N_661,In_608,In_6);
or U662 (N_662,In_131,In_302);
nor U663 (N_663,In_422,In_293);
or U664 (N_664,In_181,In_339);
nor U665 (N_665,In_954,In_297);
nand U666 (N_666,In_969,In_420);
nand U667 (N_667,In_337,In_873);
or U668 (N_668,In_784,In_562);
or U669 (N_669,In_50,In_976);
xor U670 (N_670,In_522,In_4);
nand U671 (N_671,In_361,In_76);
or U672 (N_672,In_658,In_47);
nor U673 (N_673,In_726,In_599);
nand U674 (N_674,In_438,In_857);
and U675 (N_675,In_759,In_680);
and U676 (N_676,In_868,In_51);
nand U677 (N_677,In_695,In_102);
and U678 (N_678,In_49,In_286);
nor U679 (N_679,In_348,In_475);
nor U680 (N_680,In_378,In_308);
and U681 (N_681,In_889,In_566);
or U682 (N_682,In_75,In_186);
nor U683 (N_683,In_655,In_985);
and U684 (N_684,In_563,In_86);
nor U685 (N_685,In_133,In_557);
and U686 (N_686,In_160,In_471);
nand U687 (N_687,In_470,In_142);
nand U688 (N_688,In_847,In_149);
nor U689 (N_689,In_20,In_729);
xor U690 (N_690,In_711,In_701);
xor U691 (N_691,In_179,In_515);
nand U692 (N_692,In_608,In_507);
xnor U693 (N_693,In_875,In_666);
or U694 (N_694,In_447,In_326);
nor U695 (N_695,In_391,In_565);
or U696 (N_696,In_45,In_766);
and U697 (N_697,In_214,In_464);
nand U698 (N_698,In_141,In_618);
and U699 (N_699,In_380,In_282);
or U700 (N_700,In_333,In_742);
nor U701 (N_701,In_511,In_397);
or U702 (N_702,In_542,In_362);
xor U703 (N_703,In_488,In_985);
nand U704 (N_704,In_487,In_806);
nor U705 (N_705,In_325,In_451);
and U706 (N_706,In_646,In_119);
nand U707 (N_707,In_500,In_871);
and U708 (N_708,In_82,In_649);
or U709 (N_709,In_232,In_952);
nor U710 (N_710,In_385,In_461);
nand U711 (N_711,In_289,In_736);
nor U712 (N_712,In_11,In_66);
nor U713 (N_713,In_908,In_131);
nand U714 (N_714,In_71,In_47);
and U715 (N_715,In_79,In_638);
nand U716 (N_716,In_28,In_519);
and U717 (N_717,In_949,In_463);
nand U718 (N_718,In_793,In_72);
nand U719 (N_719,In_410,In_561);
and U720 (N_720,In_481,In_809);
and U721 (N_721,In_965,In_451);
nor U722 (N_722,In_130,In_908);
nor U723 (N_723,In_569,In_704);
nor U724 (N_724,In_403,In_351);
or U725 (N_725,In_407,In_48);
nand U726 (N_726,In_847,In_899);
xnor U727 (N_727,In_454,In_695);
or U728 (N_728,In_223,In_689);
nor U729 (N_729,In_352,In_935);
nand U730 (N_730,In_768,In_36);
or U731 (N_731,In_490,In_999);
or U732 (N_732,In_243,In_283);
and U733 (N_733,In_83,In_828);
or U734 (N_734,In_409,In_604);
xor U735 (N_735,In_45,In_487);
nor U736 (N_736,In_737,In_261);
and U737 (N_737,In_183,In_561);
nand U738 (N_738,In_15,In_888);
nand U739 (N_739,In_676,In_543);
or U740 (N_740,In_566,In_329);
nor U741 (N_741,In_833,In_88);
nor U742 (N_742,In_401,In_226);
nor U743 (N_743,In_663,In_264);
xnor U744 (N_744,In_306,In_904);
and U745 (N_745,In_513,In_914);
or U746 (N_746,In_146,In_495);
nand U747 (N_747,In_767,In_579);
nand U748 (N_748,In_233,In_865);
xnor U749 (N_749,In_885,In_367);
nand U750 (N_750,In_855,In_66);
nor U751 (N_751,In_222,In_106);
and U752 (N_752,In_366,In_531);
and U753 (N_753,In_435,In_905);
or U754 (N_754,In_838,In_257);
xnor U755 (N_755,In_712,In_70);
or U756 (N_756,In_839,In_652);
or U757 (N_757,In_794,In_690);
xor U758 (N_758,In_487,In_979);
and U759 (N_759,In_624,In_178);
xor U760 (N_760,In_813,In_841);
and U761 (N_761,In_524,In_980);
nor U762 (N_762,In_105,In_613);
nand U763 (N_763,In_681,In_442);
nand U764 (N_764,In_95,In_159);
and U765 (N_765,In_86,In_37);
xor U766 (N_766,In_181,In_389);
nand U767 (N_767,In_686,In_139);
nor U768 (N_768,In_860,In_700);
nor U769 (N_769,In_971,In_121);
nand U770 (N_770,In_221,In_987);
or U771 (N_771,In_624,In_665);
or U772 (N_772,In_172,In_134);
nand U773 (N_773,In_187,In_339);
and U774 (N_774,In_327,In_936);
and U775 (N_775,In_703,In_706);
and U776 (N_776,In_472,In_738);
nand U777 (N_777,In_719,In_407);
or U778 (N_778,In_314,In_309);
nand U779 (N_779,In_652,In_681);
and U780 (N_780,In_236,In_209);
nand U781 (N_781,In_969,In_406);
or U782 (N_782,In_964,In_436);
and U783 (N_783,In_526,In_401);
nor U784 (N_784,In_392,In_366);
nor U785 (N_785,In_347,In_843);
nor U786 (N_786,In_319,In_573);
nand U787 (N_787,In_590,In_802);
nand U788 (N_788,In_199,In_7);
nor U789 (N_789,In_43,In_633);
nor U790 (N_790,In_170,In_792);
nand U791 (N_791,In_796,In_865);
and U792 (N_792,In_792,In_681);
xnor U793 (N_793,In_483,In_381);
or U794 (N_794,In_699,In_405);
nand U795 (N_795,In_570,In_734);
nor U796 (N_796,In_201,In_649);
nor U797 (N_797,In_660,In_693);
and U798 (N_798,In_677,In_868);
and U799 (N_799,In_975,In_782);
or U800 (N_800,In_715,In_33);
or U801 (N_801,In_172,In_25);
nand U802 (N_802,In_899,In_410);
nor U803 (N_803,In_39,In_497);
nor U804 (N_804,In_895,In_205);
and U805 (N_805,In_717,In_194);
nand U806 (N_806,In_747,In_303);
or U807 (N_807,In_895,In_569);
xnor U808 (N_808,In_517,In_25);
and U809 (N_809,In_769,In_411);
or U810 (N_810,In_406,In_402);
or U811 (N_811,In_891,In_661);
nand U812 (N_812,In_573,In_170);
nand U813 (N_813,In_392,In_574);
or U814 (N_814,In_191,In_916);
and U815 (N_815,In_901,In_907);
or U816 (N_816,In_280,In_517);
and U817 (N_817,In_402,In_9);
nand U818 (N_818,In_633,In_396);
nor U819 (N_819,In_69,In_547);
or U820 (N_820,In_819,In_635);
or U821 (N_821,In_331,In_696);
or U822 (N_822,In_754,In_614);
nand U823 (N_823,In_376,In_429);
and U824 (N_824,In_984,In_563);
or U825 (N_825,In_477,In_468);
nor U826 (N_826,In_362,In_660);
or U827 (N_827,In_608,In_228);
nand U828 (N_828,In_197,In_606);
nand U829 (N_829,In_694,In_356);
or U830 (N_830,In_715,In_808);
nor U831 (N_831,In_64,In_897);
or U832 (N_832,In_156,In_522);
nor U833 (N_833,In_182,In_553);
nand U834 (N_834,In_435,In_419);
and U835 (N_835,In_8,In_192);
and U836 (N_836,In_74,In_623);
or U837 (N_837,In_846,In_897);
nand U838 (N_838,In_638,In_404);
nand U839 (N_839,In_942,In_627);
and U840 (N_840,In_158,In_775);
nor U841 (N_841,In_547,In_498);
xnor U842 (N_842,In_756,In_861);
nor U843 (N_843,In_340,In_297);
nand U844 (N_844,In_582,In_454);
and U845 (N_845,In_225,In_515);
nor U846 (N_846,In_14,In_405);
and U847 (N_847,In_163,In_754);
or U848 (N_848,In_167,In_423);
xnor U849 (N_849,In_876,In_886);
and U850 (N_850,In_121,In_133);
or U851 (N_851,In_501,In_505);
nor U852 (N_852,In_349,In_398);
or U853 (N_853,In_506,In_994);
or U854 (N_854,In_845,In_431);
nor U855 (N_855,In_898,In_23);
nand U856 (N_856,In_259,In_336);
and U857 (N_857,In_685,In_563);
xnor U858 (N_858,In_102,In_291);
and U859 (N_859,In_762,In_565);
and U860 (N_860,In_40,In_120);
and U861 (N_861,In_939,In_723);
nor U862 (N_862,In_132,In_961);
or U863 (N_863,In_787,In_256);
nand U864 (N_864,In_963,In_83);
xor U865 (N_865,In_244,In_872);
nand U866 (N_866,In_850,In_738);
nor U867 (N_867,In_920,In_182);
nor U868 (N_868,In_846,In_639);
or U869 (N_869,In_605,In_217);
or U870 (N_870,In_205,In_808);
nor U871 (N_871,In_521,In_630);
nor U872 (N_872,In_502,In_540);
nand U873 (N_873,In_513,In_908);
and U874 (N_874,In_601,In_754);
or U875 (N_875,In_541,In_38);
nor U876 (N_876,In_583,In_410);
nand U877 (N_877,In_892,In_977);
xnor U878 (N_878,In_351,In_36);
nand U879 (N_879,In_89,In_595);
nand U880 (N_880,In_482,In_576);
nor U881 (N_881,In_533,In_590);
or U882 (N_882,In_368,In_305);
nand U883 (N_883,In_648,In_713);
and U884 (N_884,In_334,In_265);
nor U885 (N_885,In_835,In_18);
and U886 (N_886,In_678,In_819);
nand U887 (N_887,In_571,In_602);
nand U888 (N_888,In_997,In_670);
nor U889 (N_889,In_276,In_378);
xor U890 (N_890,In_591,In_307);
nand U891 (N_891,In_902,In_716);
nor U892 (N_892,In_48,In_665);
or U893 (N_893,In_42,In_128);
nand U894 (N_894,In_637,In_646);
xor U895 (N_895,In_622,In_805);
xnor U896 (N_896,In_966,In_794);
or U897 (N_897,In_881,In_56);
and U898 (N_898,In_963,In_442);
or U899 (N_899,In_563,In_709);
or U900 (N_900,In_201,In_840);
or U901 (N_901,In_793,In_338);
and U902 (N_902,In_506,In_963);
nand U903 (N_903,In_943,In_989);
xnor U904 (N_904,In_584,In_197);
xnor U905 (N_905,In_811,In_370);
or U906 (N_906,In_313,In_70);
nand U907 (N_907,In_429,In_260);
nand U908 (N_908,In_269,In_118);
nor U909 (N_909,In_946,In_269);
or U910 (N_910,In_962,In_564);
and U911 (N_911,In_451,In_883);
and U912 (N_912,In_577,In_360);
nand U913 (N_913,In_525,In_429);
nand U914 (N_914,In_605,In_594);
or U915 (N_915,In_571,In_761);
nor U916 (N_916,In_47,In_571);
or U917 (N_917,In_45,In_414);
and U918 (N_918,In_949,In_540);
and U919 (N_919,In_364,In_704);
nand U920 (N_920,In_151,In_830);
nor U921 (N_921,In_726,In_282);
and U922 (N_922,In_468,In_864);
nor U923 (N_923,In_143,In_476);
nor U924 (N_924,In_438,In_811);
nor U925 (N_925,In_331,In_499);
nor U926 (N_926,In_352,In_58);
nand U927 (N_927,In_445,In_856);
nand U928 (N_928,In_250,In_118);
and U929 (N_929,In_404,In_412);
or U930 (N_930,In_734,In_987);
or U931 (N_931,In_173,In_495);
and U932 (N_932,In_817,In_442);
nor U933 (N_933,In_269,In_539);
nor U934 (N_934,In_578,In_617);
and U935 (N_935,In_618,In_190);
and U936 (N_936,In_131,In_273);
or U937 (N_937,In_914,In_650);
nand U938 (N_938,In_932,In_205);
or U939 (N_939,In_744,In_443);
and U940 (N_940,In_259,In_395);
xor U941 (N_941,In_114,In_900);
nor U942 (N_942,In_993,In_567);
or U943 (N_943,In_275,In_317);
and U944 (N_944,In_93,In_733);
or U945 (N_945,In_381,In_974);
xnor U946 (N_946,In_86,In_97);
or U947 (N_947,In_143,In_237);
nor U948 (N_948,In_809,In_752);
and U949 (N_949,In_216,In_419);
xor U950 (N_950,In_14,In_579);
nor U951 (N_951,In_949,In_185);
xor U952 (N_952,In_704,In_162);
nor U953 (N_953,In_886,In_994);
nor U954 (N_954,In_620,In_305);
xnor U955 (N_955,In_275,In_342);
or U956 (N_956,In_732,In_404);
and U957 (N_957,In_717,In_243);
and U958 (N_958,In_216,In_702);
nand U959 (N_959,In_856,In_71);
nand U960 (N_960,In_446,In_318);
nor U961 (N_961,In_810,In_661);
nand U962 (N_962,In_397,In_142);
nor U963 (N_963,In_494,In_890);
nor U964 (N_964,In_469,In_912);
and U965 (N_965,In_526,In_822);
xor U966 (N_966,In_866,In_190);
nor U967 (N_967,In_142,In_717);
nor U968 (N_968,In_890,In_334);
nand U969 (N_969,In_696,In_631);
nor U970 (N_970,In_254,In_239);
and U971 (N_971,In_597,In_955);
or U972 (N_972,In_994,In_261);
or U973 (N_973,In_339,In_291);
nand U974 (N_974,In_143,In_98);
xnor U975 (N_975,In_522,In_205);
or U976 (N_976,In_819,In_763);
or U977 (N_977,In_963,In_172);
nand U978 (N_978,In_62,In_757);
xor U979 (N_979,In_69,In_600);
nand U980 (N_980,In_345,In_164);
nor U981 (N_981,In_782,In_548);
nor U982 (N_982,In_544,In_812);
nor U983 (N_983,In_82,In_486);
or U984 (N_984,In_389,In_960);
nor U985 (N_985,In_287,In_539);
nand U986 (N_986,In_274,In_351);
and U987 (N_987,In_727,In_5);
or U988 (N_988,In_131,In_327);
or U989 (N_989,In_613,In_771);
and U990 (N_990,In_604,In_1);
or U991 (N_991,In_157,In_309);
nand U992 (N_992,In_996,In_233);
and U993 (N_993,In_161,In_792);
nand U994 (N_994,In_743,In_521);
nand U995 (N_995,In_733,In_374);
nand U996 (N_996,In_348,In_439);
xor U997 (N_997,In_924,In_478);
and U998 (N_998,In_431,In_454);
nand U999 (N_999,In_547,In_672);
nand U1000 (N_1000,N_67,N_19);
and U1001 (N_1001,N_362,N_882);
and U1002 (N_1002,N_546,N_545);
and U1003 (N_1003,N_473,N_62);
nor U1004 (N_1004,N_820,N_971);
nor U1005 (N_1005,N_942,N_678);
nor U1006 (N_1006,N_395,N_975);
nand U1007 (N_1007,N_755,N_339);
nor U1008 (N_1008,N_415,N_303);
nor U1009 (N_1009,N_736,N_624);
or U1010 (N_1010,N_246,N_80);
xnor U1011 (N_1011,N_326,N_850);
nor U1012 (N_1012,N_503,N_717);
nand U1013 (N_1013,N_720,N_286);
nand U1014 (N_1014,N_550,N_846);
nand U1015 (N_1015,N_579,N_306);
xnor U1016 (N_1016,N_281,N_895);
and U1017 (N_1017,N_636,N_158);
nor U1018 (N_1018,N_154,N_474);
nor U1019 (N_1019,N_94,N_176);
or U1020 (N_1020,N_481,N_144);
and U1021 (N_1021,N_581,N_741);
or U1022 (N_1022,N_276,N_22);
nand U1023 (N_1023,N_799,N_890);
nor U1024 (N_1024,N_431,N_310);
xor U1025 (N_1025,N_702,N_382);
and U1026 (N_1026,N_47,N_124);
and U1027 (N_1027,N_860,N_322);
nand U1028 (N_1028,N_355,N_617);
nand U1029 (N_1029,N_968,N_112);
or U1030 (N_1030,N_920,N_990);
nand U1031 (N_1031,N_252,N_423);
or U1032 (N_1032,N_663,N_771);
or U1033 (N_1033,N_48,N_831);
or U1034 (N_1034,N_390,N_806);
and U1035 (N_1035,N_6,N_951);
nand U1036 (N_1036,N_563,N_89);
nor U1037 (N_1037,N_294,N_120);
or U1038 (N_1038,N_236,N_163);
nor U1039 (N_1039,N_714,N_956);
and U1040 (N_1040,N_819,N_602);
nand U1041 (N_1041,N_227,N_599);
and U1042 (N_1042,N_607,N_271);
nand U1043 (N_1043,N_433,N_943);
and U1044 (N_1044,N_471,N_90);
or U1045 (N_1045,N_959,N_134);
and U1046 (N_1046,N_878,N_705);
xnor U1047 (N_1047,N_967,N_765);
or U1048 (N_1048,N_74,N_997);
and U1049 (N_1049,N_265,N_987);
xor U1050 (N_1050,N_369,N_643);
nand U1051 (N_1051,N_254,N_147);
or U1052 (N_1052,N_349,N_283);
or U1053 (N_1053,N_760,N_424);
or U1054 (N_1054,N_105,N_111);
nand U1055 (N_1055,N_278,N_569);
and U1056 (N_1056,N_786,N_743);
and U1057 (N_1057,N_325,N_425);
or U1058 (N_1058,N_148,N_564);
nor U1059 (N_1059,N_204,N_312);
or U1060 (N_1060,N_691,N_940);
nand U1061 (N_1061,N_353,N_331);
or U1062 (N_1062,N_186,N_722);
and U1063 (N_1063,N_950,N_202);
nor U1064 (N_1064,N_7,N_20);
and U1065 (N_1065,N_634,N_804);
nand U1066 (N_1066,N_296,N_522);
nor U1067 (N_1067,N_110,N_213);
or U1068 (N_1068,N_251,N_827);
nor U1069 (N_1069,N_776,N_696);
or U1070 (N_1070,N_73,N_809);
and U1071 (N_1071,N_243,N_169);
xor U1072 (N_1072,N_610,N_348);
nand U1073 (N_1073,N_58,N_407);
or U1074 (N_1074,N_554,N_674);
nor U1075 (N_1075,N_561,N_323);
and U1076 (N_1076,N_410,N_964);
nand U1077 (N_1077,N_963,N_397);
or U1078 (N_1078,N_12,N_157);
and U1079 (N_1079,N_883,N_291);
nand U1080 (N_1080,N_637,N_576);
nand U1081 (N_1081,N_64,N_716);
nor U1082 (N_1082,N_5,N_66);
or U1083 (N_1083,N_29,N_393);
nor U1084 (N_1084,N_396,N_700);
and U1085 (N_1085,N_909,N_256);
nor U1086 (N_1086,N_656,N_69);
and U1087 (N_1087,N_268,N_906);
nand U1088 (N_1088,N_233,N_181);
and U1089 (N_1089,N_289,N_752);
and U1090 (N_1090,N_869,N_224);
nor U1091 (N_1091,N_622,N_40);
nand U1092 (N_1092,N_866,N_653);
nand U1093 (N_1093,N_733,N_635);
or U1094 (N_1094,N_146,N_217);
and U1095 (N_1095,N_960,N_936);
and U1096 (N_1096,N_223,N_703);
nand U1097 (N_1097,N_807,N_982);
xor U1098 (N_1098,N_619,N_215);
nor U1099 (N_1099,N_125,N_896);
nor U1100 (N_1100,N_342,N_562);
or U1101 (N_1101,N_475,N_930);
xor U1102 (N_1102,N_17,N_992);
or U1103 (N_1103,N_195,N_293);
nand U1104 (N_1104,N_208,N_808);
or U1105 (N_1105,N_958,N_483);
nor U1106 (N_1106,N_308,N_498);
and U1107 (N_1107,N_317,N_924);
nand U1108 (N_1108,N_26,N_13);
or U1109 (N_1109,N_680,N_32);
and U1110 (N_1110,N_63,N_641);
nor U1111 (N_1111,N_220,N_790);
nand U1112 (N_1112,N_472,N_161);
nor U1113 (N_1113,N_182,N_302);
and U1114 (N_1114,N_46,N_83);
and U1115 (N_1115,N_3,N_870);
and U1116 (N_1116,N_626,N_152);
and U1117 (N_1117,N_409,N_568);
or U1118 (N_1118,N_451,N_638);
nand U1119 (N_1119,N_874,N_973);
nor U1120 (N_1120,N_615,N_439);
or U1121 (N_1121,N_847,N_668);
nand U1122 (N_1122,N_718,N_295);
and U1123 (N_1123,N_368,N_8);
nor U1124 (N_1124,N_976,N_868);
or U1125 (N_1125,N_872,N_487);
or U1126 (N_1126,N_694,N_701);
nor U1127 (N_1127,N_59,N_387);
nor U1128 (N_1128,N_121,N_623);
nor U1129 (N_1129,N_779,N_954);
and U1130 (N_1130,N_721,N_957);
xnor U1131 (N_1131,N_685,N_378);
nand U1132 (N_1132,N_84,N_570);
and U1133 (N_1133,N_572,N_458);
and U1134 (N_1134,N_854,N_681);
or U1135 (N_1135,N_240,N_404);
nor U1136 (N_1136,N_259,N_994);
and U1137 (N_1137,N_961,N_127);
and U1138 (N_1138,N_785,N_537);
nand U1139 (N_1139,N_797,N_732);
and U1140 (N_1140,N_379,N_504);
xnor U1141 (N_1141,N_632,N_174);
nor U1142 (N_1142,N_341,N_782);
and U1143 (N_1143,N_788,N_130);
and U1144 (N_1144,N_71,N_898);
or U1145 (N_1145,N_260,N_513);
or U1146 (N_1146,N_794,N_333);
or U1147 (N_1147,N_78,N_477);
xor U1148 (N_1148,N_2,N_507);
nand U1149 (N_1149,N_320,N_666);
and U1150 (N_1150,N_842,N_447);
nand U1151 (N_1151,N_995,N_298);
or U1152 (N_1152,N_363,N_115);
and U1153 (N_1153,N_500,N_993);
or U1154 (N_1154,N_783,N_170);
and U1155 (N_1155,N_996,N_177);
or U1156 (N_1156,N_324,N_597);
nor U1157 (N_1157,N_465,N_109);
nand U1158 (N_1158,N_81,N_955);
nor U1159 (N_1159,N_889,N_15);
and U1160 (N_1160,N_275,N_907);
and U1161 (N_1161,N_775,N_919);
and U1162 (N_1162,N_427,N_879);
and U1163 (N_1163,N_750,N_962);
nor U1164 (N_1164,N_515,N_894);
nand U1165 (N_1165,N_82,N_33);
and U1166 (N_1166,N_273,N_284);
or U1167 (N_1167,N_117,N_4);
and U1168 (N_1168,N_205,N_778);
nand U1169 (N_1169,N_699,N_143);
nand U1170 (N_1170,N_139,N_644);
xnor U1171 (N_1171,N_625,N_201);
nor U1172 (N_1172,N_748,N_460);
or U1173 (N_1173,N_351,N_385);
nor U1174 (N_1174,N_627,N_664);
and U1175 (N_1175,N_495,N_30);
and U1176 (N_1176,N_908,N_715);
nand U1177 (N_1177,N_887,N_469);
or U1178 (N_1178,N_318,N_713);
or U1179 (N_1179,N_740,N_31);
nor U1180 (N_1180,N_164,N_559);
nand U1181 (N_1181,N_925,N_594);
and U1182 (N_1182,N_414,N_859);
or U1183 (N_1183,N_595,N_816);
or U1184 (N_1184,N_102,N_784);
nand U1185 (N_1185,N_49,N_328);
nand U1186 (N_1186,N_985,N_949);
and U1187 (N_1187,N_123,N_670);
and U1188 (N_1188,N_343,N_767);
nand U1189 (N_1189,N_646,N_403);
nor U1190 (N_1190,N_272,N_96);
nor U1191 (N_1191,N_821,N_165);
nor U1192 (N_1192,N_590,N_801);
or U1193 (N_1193,N_822,N_523);
nor U1194 (N_1194,N_867,N_365);
nor U1195 (N_1195,N_974,N_727);
nor U1196 (N_1196,N_430,N_86);
or U1197 (N_1197,N_313,N_711);
nor U1198 (N_1198,N_408,N_654);
nand U1199 (N_1199,N_915,N_255);
nand U1200 (N_1200,N_560,N_840);
xor U1201 (N_1201,N_448,N_45);
nand U1202 (N_1202,N_344,N_917);
and U1203 (N_1203,N_983,N_329);
nor U1204 (N_1204,N_861,N_573);
nand U1205 (N_1205,N_244,N_669);
and U1206 (N_1206,N_839,N_327);
nand U1207 (N_1207,N_391,N_466);
nor U1208 (N_1208,N_234,N_836);
nor U1209 (N_1209,N_524,N_762);
nor U1210 (N_1210,N_54,N_489);
nor U1211 (N_1211,N_944,N_119);
nand U1212 (N_1212,N_979,N_231);
and U1213 (N_1213,N_938,N_432);
and U1214 (N_1214,N_151,N_843);
nor U1215 (N_1215,N_486,N_18);
or U1216 (N_1216,N_939,N_114);
nand U1217 (N_1217,N_384,N_239);
nand U1218 (N_1218,N_527,N_263);
xor U1219 (N_1219,N_849,N_528);
nor U1220 (N_1220,N_198,N_297);
nand U1221 (N_1221,N_918,N_604);
and U1222 (N_1222,N_690,N_216);
and U1223 (N_1223,N_912,N_65);
and U1224 (N_1224,N_677,N_200);
or U1225 (N_1225,N_738,N_586);
nand U1226 (N_1226,N_57,N_707);
nor U1227 (N_1227,N_766,N_916);
nand U1228 (N_1228,N_519,N_845);
and U1229 (N_1229,N_270,N_496);
nand U1230 (N_1230,N_145,N_682);
and U1231 (N_1231,N_336,N_757);
nand U1232 (N_1232,N_657,N_374);
nor U1233 (N_1233,N_361,N_467);
xnor U1234 (N_1234,N_135,N_761);
nor U1235 (N_1235,N_616,N_315);
and U1236 (N_1236,N_479,N_372);
or U1237 (N_1237,N_356,N_724);
xor U1238 (N_1238,N_903,N_946);
nand U1239 (N_1239,N_826,N_730);
nand U1240 (N_1240,N_659,N_777);
nand U1241 (N_1241,N_647,N_444);
or U1242 (N_1242,N_877,N_470);
nand U1243 (N_1243,N_91,N_108);
and U1244 (N_1244,N_340,N_539);
nand U1245 (N_1245,N_183,N_103);
nor U1246 (N_1246,N_98,N_923);
and U1247 (N_1247,N_529,N_462);
and U1248 (N_1248,N_825,N_932);
or U1249 (N_1249,N_28,N_989);
nor U1250 (N_1250,N_789,N_621);
nor U1251 (N_1251,N_505,N_484);
or U1252 (N_1252,N_43,N_731);
and U1253 (N_1253,N_888,N_299);
nor U1254 (N_1254,N_858,N_697);
nand U1255 (N_1255,N_620,N_712);
or U1256 (N_1256,N_490,N_132);
nand U1257 (N_1257,N_803,N_491);
nor U1258 (N_1258,N_575,N_904);
nand U1259 (N_1259,N_218,N_250);
xnor U1260 (N_1260,N_37,N_436);
and U1261 (N_1261,N_367,N_540);
nand U1262 (N_1262,N_608,N_138);
or U1263 (N_1263,N_305,N_100);
or U1264 (N_1264,N_814,N_751);
or U1265 (N_1265,N_640,N_747);
nor U1266 (N_1266,N_734,N_358);
xnor U1267 (N_1267,N_222,N_851);
xor U1268 (N_1268,N_709,N_947);
nor U1269 (N_1269,N_655,N_68);
or U1270 (N_1270,N_591,N_41);
and U1271 (N_1271,N_756,N_21);
nand U1272 (N_1272,N_815,N_307);
and U1273 (N_1273,N_426,N_671);
nor U1274 (N_1274,N_639,N_301);
and U1275 (N_1275,N_247,N_88);
or U1276 (N_1276,N_421,N_835);
nor U1277 (N_1277,N_435,N_692);
nor U1278 (N_1278,N_97,N_927);
nand U1279 (N_1279,N_934,N_675);
nor U1280 (N_1280,N_848,N_945);
nor U1281 (N_1281,N_113,N_593);
and U1282 (N_1282,N_548,N_922);
or U1283 (N_1283,N_998,N_857);
nand U1284 (N_1284,N_862,N_443);
nor U1285 (N_1285,N_377,N_864);
or U1286 (N_1286,N_416,N_589);
and U1287 (N_1287,N_667,N_454);
nor U1288 (N_1288,N_542,N_953);
nand U1289 (N_1289,N_791,N_445);
or U1290 (N_1290,N_514,N_520);
nor U1291 (N_1291,N_763,N_422);
and U1292 (N_1292,N_613,N_314);
nand U1293 (N_1293,N_149,N_459);
nand U1294 (N_1294,N_173,N_603);
or U1295 (N_1295,N_886,N_536);
nor U1296 (N_1296,N_832,N_901);
and U1297 (N_1297,N_189,N_592);
or U1298 (N_1298,N_684,N_338);
nand U1299 (N_1299,N_770,N_311);
and U1300 (N_1300,N_335,N_798);
and U1301 (N_1301,N_196,N_499);
or U1302 (N_1302,N_206,N_892);
and U1303 (N_1303,N_556,N_582);
nand U1304 (N_1304,N_502,N_402);
nor U1305 (N_1305,N_492,N_688);
nand U1306 (N_1306,N_461,N_70);
nor U1307 (N_1307,N_253,N_754);
or U1308 (N_1308,N_881,N_856);
and U1309 (N_1309,N_36,N_300);
nand U1310 (N_1310,N_510,N_75);
nor U1311 (N_1311,N_966,N_991);
and U1312 (N_1312,N_446,N_10);
and U1313 (N_1313,N_287,N_381);
nand U1314 (N_1314,N_187,N_14);
nand U1315 (N_1315,N_662,N_482);
nand U1316 (N_1316,N_978,N_370);
xnor U1317 (N_1317,N_229,N_172);
or U1318 (N_1318,N_199,N_35);
nand U1319 (N_1319,N_525,N_203);
and U1320 (N_1320,N_429,N_530);
xnor U1321 (N_1321,N_828,N_577);
nor U1322 (N_1322,N_931,N_977);
and U1323 (N_1323,N_279,N_665);
nand U1324 (N_1324,N_142,N_442);
xnor U1325 (N_1325,N_417,N_133);
or U1326 (N_1326,N_549,N_280);
and U1327 (N_1327,N_245,N_375);
and U1328 (N_1328,N_566,N_648);
nor U1329 (N_1329,N_194,N_389);
and U1330 (N_1330,N_269,N_190);
and U1331 (N_1331,N_708,N_792);
or U1332 (N_1332,N_334,N_508);
nand U1333 (N_1333,N_99,N_457);
nor U1334 (N_1334,N_179,N_516);
nand U1335 (N_1335,N_605,N_478);
and U1336 (N_1336,N_695,N_267);
nand U1337 (N_1337,N_781,N_27);
nand U1338 (N_1338,N_494,N_116);
nand U1339 (N_1339,N_511,N_453);
and U1340 (N_1340,N_332,N_676);
and U1341 (N_1341,N_352,N_153);
nor U1342 (N_1342,N_746,N_541);
or U1343 (N_1343,N_405,N_558);
nand U1344 (N_1344,N_290,N_897);
nand U1345 (N_1345,N_764,N_434);
and U1346 (N_1346,N_588,N_380);
nand U1347 (N_1347,N_769,N_76);
and U1348 (N_1348,N_574,N_261);
or U1349 (N_1349,N_191,N_980);
nand U1350 (N_1350,N_192,N_350);
nand U1351 (N_1351,N_180,N_129);
nor U1352 (N_1352,N_476,N_428);
nor U1353 (N_1353,N_9,N_79);
or U1354 (N_1354,N_140,N_241);
nor U1355 (N_1355,N_506,N_652);
or U1356 (N_1356,N_532,N_230);
and U1357 (N_1357,N_61,N_366);
or U1358 (N_1358,N_759,N_933);
nand U1359 (N_1359,N_587,N_753);
or U1360 (N_1360,N_406,N_723);
and U1361 (N_1361,N_884,N_468);
or U1362 (N_1362,N_166,N_571);
nor U1363 (N_1363,N_106,N_811);
nand U1364 (N_1364,N_321,N_565);
nand U1365 (N_1365,N_521,N_875);
xor U1366 (N_1366,N_394,N_661);
nand U1367 (N_1367,N_282,N_631);
nand U1368 (N_1368,N_53,N_52);
and U1369 (N_1369,N_50,N_11);
and U1370 (N_1370,N_900,N_400);
or U1371 (N_1371,N_493,N_383);
xor U1372 (N_1372,N_93,N_824);
nor U1373 (N_1373,N_710,N_893);
and U1374 (N_1374,N_137,N_885);
nor U1375 (N_1375,N_758,N_686);
nand U1376 (N_1376,N_441,N_292);
nand U1377 (N_1377,N_210,N_650);
or U1378 (N_1378,N_360,N_813);
nor U1379 (N_1379,N_118,N_225);
nor U1380 (N_1380,N_171,N_262);
and U1381 (N_1381,N_288,N_207);
xnor U1382 (N_1382,N_464,N_683);
xor U1383 (N_1383,N_871,N_704);
and U1384 (N_1384,N_899,N_649);
and U1385 (N_1385,N_768,N_745);
nand U1386 (N_1386,N_450,N_772);
nand U1387 (N_1387,N_969,N_509);
or U1388 (N_1388,N_551,N_398);
and U1389 (N_1389,N_698,N_175);
or U1390 (N_1390,N_178,N_679);
nand U1391 (N_1391,N_238,N_126);
and U1392 (N_1392,N_485,N_232);
or U1393 (N_1393,N_800,N_555);
and U1394 (N_1394,N_719,N_578);
nand U1395 (N_1395,N_463,N_226);
and U1396 (N_1396,N_480,N_948);
and U1397 (N_1397,N_197,N_596);
or U1398 (N_1398,N_347,N_628);
nor U1399 (N_1399,N_926,N_184);
and U1400 (N_1400,N_412,N_986);
or U1401 (N_1401,N_833,N_584);
nor U1402 (N_1402,N_981,N_24);
or U1403 (N_1403,N_249,N_357);
xnor U1404 (N_1404,N_774,N_228);
or U1405 (N_1405,N_51,N_729);
and U1406 (N_1406,N_128,N_354);
nor U1407 (N_1407,N_557,N_865);
or U1408 (N_1408,N_689,N_972);
nor U1409 (N_1409,N_823,N_531);
or U1410 (N_1410,N_609,N_911);
or U1411 (N_1411,N_55,N_209);
nor U1412 (N_1412,N_304,N_411);
or U1413 (N_1413,N_988,N_952);
and U1414 (N_1414,N_876,N_941);
xor U1415 (N_1415,N_693,N_812);
nor U1416 (N_1416,N_56,N_552);
nor U1417 (N_1417,N_185,N_891);
nand U1418 (N_1418,N_802,N_449);
nand U1419 (N_1419,N_543,N_219);
and U1420 (N_1420,N_438,N_319);
and U1421 (N_1421,N_497,N_107);
and U1422 (N_1422,N_316,N_852);
or U1423 (N_1423,N_737,N_155);
and U1424 (N_1424,N_193,N_618);
or U1425 (N_1425,N_274,N_92);
or U1426 (N_1426,N_399,N_104);
xnor U1427 (N_1427,N_346,N_266);
or U1428 (N_1428,N_418,N_376);
nor U1429 (N_1429,N_518,N_77);
nand U1430 (N_1430,N_534,N_242);
xor U1431 (N_1431,N_818,N_25);
nand U1432 (N_1432,N_214,N_830);
or U1433 (N_1433,N_42,N_285);
nand U1434 (N_1434,N_614,N_706);
or U1435 (N_1435,N_264,N_401);
nor U1436 (N_1436,N_642,N_873);
or U1437 (N_1437,N_452,N_928);
and U1438 (N_1438,N_585,N_501);
and U1439 (N_1439,N_965,N_606);
or U1440 (N_1440,N_795,N_567);
nor U1441 (N_1441,N_455,N_156);
nor U1442 (N_1442,N_373,N_488);
nand U1443 (N_1443,N_159,N_612);
nand U1444 (N_1444,N_863,N_16);
and U1445 (N_1445,N_773,N_645);
and U1446 (N_1446,N_526,N_660);
nor U1447 (N_1447,N_167,N_583);
nor U1448 (N_1448,N_935,N_914);
nor U1449 (N_1449,N_937,N_359);
nand U1450 (N_1450,N_535,N_744);
and U1451 (N_1451,N_910,N_728);
nor U1452 (N_1452,N_95,N_60);
and U1453 (N_1453,N_598,N_309);
and U1454 (N_1454,N_547,N_413);
nand U1455 (N_1455,N_725,N_880);
nor U1456 (N_1456,N_844,N_834);
nor U1457 (N_1457,N_672,N_364);
and U1458 (N_1458,N_437,N_580);
and U1459 (N_1459,N_136,N_905);
or U1460 (N_1460,N_150,N_277);
nor U1461 (N_1461,N_902,N_44);
nor U1462 (N_1462,N_1,N_419);
and U1463 (N_1463,N_600,N_999);
nor U1464 (N_1464,N_921,N_553);
nor U1465 (N_1465,N_841,N_787);
and U1466 (N_1466,N_141,N_386);
nor U1467 (N_1467,N_188,N_726);
nand U1468 (N_1468,N_160,N_162);
nor U1469 (N_1469,N_793,N_630);
or U1470 (N_1470,N_805,N_456);
nor U1471 (N_1471,N_913,N_658);
xor U1472 (N_1472,N_739,N_237);
nor U1473 (N_1473,N_440,N_258);
nor U1474 (N_1474,N_72,N_34);
or U1475 (N_1475,N_122,N_248);
and U1476 (N_1476,N_85,N_512);
xnor U1477 (N_1477,N_829,N_39);
and U1478 (N_1478,N_388,N_673);
nor U1479 (N_1479,N_212,N_330);
or U1480 (N_1480,N_101,N_257);
nor U1481 (N_1481,N_742,N_23);
nand U1482 (N_1482,N_853,N_517);
xor U1483 (N_1483,N_970,N_780);
and U1484 (N_1484,N_810,N_87);
xnor U1485 (N_1485,N_796,N_371);
or U1486 (N_1486,N_984,N_749);
nand U1487 (N_1487,N_611,N_601);
nand U1488 (N_1488,N_629,N_633);
or U1489 (N_1489,N_533,N_235);
nand U1490 (N_1490,N_131,N_392);
or U1491 (N_1491,N_544,N_168);
nor U1492 (N_1492,N_538,N_855);
and U1493 (N_1493,N_735,N_817);
and U1494 (N_1494,N_838,N_651);
nor U1495 (N_1495,N_337,N_420);
nand U1496 (N_1496,N_837,N_929);
xnor U1497 (N_1497,N_211,N_345);
and U1498 (N_1498,N_38,N_221);
nand U1499 (N_1499,N_0,N_687);
nand U1500 (N_1500,N_752,N_985);
or U1501 (N_1501,N_713,N_327);
nor U1502 (N_1502,N_398,N_808);
and U1503 (N_1503,N_194,N_163);
and U1504 (N_1504,N_64,N_89);
nand U1505 (N_1505,N_25,N_45);
nor U1506 (N_1506,N_235,N_16);
xnor U1507 (N_1507,N_53,N_702);
and U1508 (N_1508,N_507,N_493);
nand U1509 (N_1509,N_592,N_658);
xor U1510 (N_1510,N_84,N_927);
nand U1511 (N_1511,N_852,N_732);
nand U1512 (N_1512,N_406,N_226);
xnor U1513 (N_1513,N_2,N_681);
nand U1514 (N_1514,N_420,N_821);
nand U1515 (N_1515,N_157,N_625);
nand U1516 (N_1516,N_677,N_543);
nor U1517 (N_1517,N_417,N_92);
xnor U1518 (N_1518,N_698,N_692);
and U1519 (N_1519,N_503,N_540);
and U1520 (N_1520,N_716,N_394);
and U1521 (N_1521,N_43,N_266);
nand U1522 (N_1522,N_711,N_672);
or U1523 (N_1523,N_826,N_231);
nand U1524 (N_1524,N_668,N_356);
and U1525 (N_1525,N_291,N_329);
and U1526 (N_1526,N_56,N_556);
or U1527 (N_1527,N_557,N_263);
or U1528 (N_1528,N_406,N_545);
and U1529 (N_1529,N_560,N_568);
or U1530 (N_1530,N_938,N_934);
or U1531 (N_1531,N_354,N_299);
or U1532 (N_1532,N_563,N_756);
xnor U1533 (N_1533,N_344,N_652);
or U1534 (N_1534,N_885,N_154);
nand U1535 (N_1535,N_819,N_295);
or U1536 (N_1536,N_761,N_30);
and U1537 (N_1537,N_609,N_261);
nor U1538 (N_1538,N_633,N_505);
nand U1539 (N_1539,N_541,N_713);
or U1540 (N_1540,N_564,N_794);
and U1541 (N_1541,N_189,N_13);
nand U1542 (N_1542,N_503,N_157);
nor U1543 (N_1543,N_331,N_241);
and U1544 (N_1544,N_153,N_702);
or U1545 (N_1545,N_752,N_587);
nor U1546 (N_1546,N_163,N_771);
nand U1547 (N_1547,N_21,N_494);
or U1548 (N_1548,N_380,N_888);
nand U1549 (N_1549,N_596,N_346);
or U1550 (N_1550,N_349,N_763);
nand U1551 (N_1551,N_238,N_780);
nor U1552 (N_1552,N_287,N_261);
nor U1553 (N_1553,N_203,N_346);
and U1554 (N_1554,N_352,N_150);
and U1555 (N_1555,N_62,N_583);
or U1556 (N_1556,N_575,N_4);
nand U1557 (N_1557,N_544,N_976);
xor U1558 (N_1558,N_972,N_653);
or U1559 (N_1559,N_229,N_720);
nor U1560 (N_1560,N_89,N_568);
nand U1561 (N_1561,N_174,N_847);
and U1562 (N_1562,N_318,N_110);
xnor U1563 (N_1563,N_143,N_19);
and U1564 (N_1564,N_311,N_478);
nor U1565 (N_1565,N_645,N_332);
and U1566 (N_1566,N_116,N_453);
nor U1567 (N_1567,N_453,N_522);
or U1568 (N_1568,N_929,N_388);
xor U1569 (N_1569,N_142,N_360);
or U1570 (N_1570,N_879,N_146);
nand U1571 (N_1571,N_716,N_392);
xor U1572 (N_1572,N_681,N_958);
or U1573 (N_1573,N_499,N_340);
nor U1574 (N_1574,N_907,N_625);
or U1575 (N_1575,N_413,N_575);
nor U1576 (N_1576,N_365,N_849);
nand U1577 (N_1577,N_467,N_474);
and U1578 (N_1578,N_399,N_798);
xor U1579 (N_1579,N_321,N_119);
or U1580 (N_1580,N_952,N_377);
and U1581 (N_1581,N_251,N_751);
or U1582 (N_1582,N_115,N_62);
nand U1583 (N_1583,N_655,N_194);
nand U1584 (N_1584,N_830,N_50);
or U1585 (N_1585,N_617,N_278);
xnor U1586 (N_1586,N_425,N_255);
xor U1587 (N_1587,N_563,N_86);
or U1588 (N_1588,N_548,N_543);
or U1589 (N_1589,N_165,N_638);
and U1590 (N_1590,N_707,N_750);
nor U1591 (N_1591,N_662,N_216);
and U1592 (N_1592,N_357,N_536);
nand U1593 (N_1593,N_258,N_771);
nand U1594 (N_1594,N_410,N_10);
and U1595 (N_1595,N_549,N_13);
nand U1596 (N_1596,N_683,N_970);
and U1597 (N_1597,N_467,N_50);
nand U1598 (N_1598,N_375,N_212);
nor U1599 (N_1599,N_294,N_310);
and U1600 (N_1600,N_270,N_581);
nor U1601 (N_1601,N_812,N_929);
xnor U1602 (N_1602,N_145,N_681);
or U1603 (N_1603,N_78,N_541);
nor U1604 (N_1604,N_978,N_225);
nand U1605 (N_1605,N_84,N_248);
nand U1606 (N_1606,N_198,N_933);
nand U1607 (N_1607,N_215,N_533);
xnor U1608 (N_1608,N_300,N_303);
xnor U1609 (N_1609,N_563,N_948);
xor U1610 (N_1610,N_93,N_345);
nand U1611 (N_1611,N_567,N_719);
nor U1612 (N_1612,N_227,N_726);
and U1613 (N_1613,N_948,N_994);
xor U1614 (N_1614,N_245,N_268);
and U1615 (N_1615,N_193,N_995);
or U1616 (N_1616,N_880,N_824);
nand U1617 (N_1617,N_498,N_742);
or U1618 (N_1618,N_835,N_130);
or U1619 (N_1619,N_951,N_842);
and U1620 (N_1620,N_353,N_803);
and U1621 (N_1621,N_578,N_138);
or U1622 (N_1622,N_198,N_95);
nor U1623 (N_1623,N_395,N_81);
nor U1624 (N_1624,N_859,N_493);
nor U1625 (N_1625,N_728,N_95);
nand U1626 (N_1626,N_837,N_544);
or U1627 (N_1627,N_73,N_173);
xor U1628 (N_1628,N_630,N_46);
or U1629 (N_1629,N_621,N_807);
and U1630 (N_1630,N_113,N_604);
nor U1631 (N_1631,N_668,N_273);
or U1632 (N_1632,N_768,N_359);
xnor U1633 (N_1633,N_967,N_100);
xnor U1634 (N_1634,N_940,N_217);
or U1635 (N_1635,N_323,N_31);
nand U1636 (N_1636,N_593,N_326);
nand U1637 (N_1637,N_299,N_707);
or U1638 (N_1638,N_627,N_500);
and U1639 (N_1639,N_489,N_579);
xor U1640 (N_1640,N_767,N_268);
and U1641 (N_1641,N_178,N_471);
and U1642 (N_1642,N_210,N_314);
nor U1643 (N_1643,N_793,N_639);
or U1644 (N_1644,N_320,N_481);
nor U1645 (N_1645,N_766,N_710);
or U1646 (N_1646,N_352,N_887);
and U1647 (N_1647,N_779,N_449);
or U1648 (N_1648,N_443,N_191);
nand U1649 (N_1649,N_21,N_432);
xor U1650 (N_1650,N_366,N_920);
nand U1651 (N_1651,N_239,N_189);
xnor U1652 (N_1652,N_155,N_812);
and U1653 (N_1653,N_725,N_278);
and U1654 (N_1654,N_160,N_521);
or U1655 (N_1655,N_422,N_581);
or U1656 (N_1656,N_806,N_670);
nand U1657 (N_1657,N_542,N_690);
or U1658 (N_1658,N_564,N_53);
and U1659 (N_1659,N_296,N_617);
nand U1660 (N_1660,N_211,N_704);
nand U1661 (N_1661,N_345,N_429);
and U1662 (N_1662,N_902,N_145);
and U1663 (N_1663,N_706,N_47);
and U1664 (N_1664,N_844,N_866);
xor U1665 (N_1665,N_802,N_960);
or U1666 (N_1666,N_573,N_903);
nand U1667 (N_1667,N_810,N_251);
nor U1668 (N_1668,N_374,N_290);
nand U1669 (N_1669,N_480,N_43);
and U1670 (N_1670,N_109,N_713);
and U1671 (N_1671,N_163,N_997);
nor U1672 (N_1672,N_225,N_677);
nor U1673 (N_1673,N_804,N_20);
and U1674 (N_1674,N_439,N_546);
nand U1675 (N_1675,N_815,N_944);
nor U1676 (N_1676,N_262,N_272);
nor U1677 (N_1677,N_427,N_797);
xnor U1678 (N_1678,N_182,N_783);
nand U1679 (N_1679,N_524,N_409);
nor U1680 (N_1680,N_676,N_281);
nand U1681 (N_1681,N_189,N_976);
or U1682 (N_1682,N_362,N_612);
xor U1683 (N_1683,N_191,N_471);
nor U1684 (N_1684,N_670,N_778);
or U1685 (N_1685,N_30,N_813);
and U1686 (N_1686,N_315,N_416);
nand U1687 (N_1687,N_377,N_258);
nand U1688 (N_1688,N_291,N_459);
nand U1689 (N_1689,N_93,N_671);
xnor U1690 (N_1690,N_498,N_764);
or U1691 (N_1691,N_72,N_71);
and U1692 (N_1692,N_590,N_425);
or U1693 (N_1693,N_491,N_482);
nand U1694 (N_1694,N_334,N_291);
and U1695 (N_1695,N_95,N_956);
nor U1696 (N_1696,N_521,N_294);
nor U1697 (N_1697,N_207,N_946);
or U1698 (N_1698,N_433,N_629);
and U1699 (N_1699,N_763,N_359);
or U1700 (N_1700,N_916,N_682);
or U1701 (N_1701,N_527,N_605);
nand U1702 (N_1702,N_464,N_761);
nor U1703 (N_1703,N_296,N_855);
and U1704 (N_1704,N_422,N_857);
nor U1705 (N_1705,N_30,N_802);
nand U1706 (N_1706,N_914,N_895);
xnor U1707 (N_1707,N_197,N_910);
nor U1708 (N_1708,N_715,N_926);
or U1709 (N_1709,N_58,N_135);
nand U1710 (N_1710,N_44,N_758);
and U1711 (N_1711,N_361,N_595);
nand U1712 (N_1712,N_798,N_991);
nor U1713 (N_1713,N_995,N_566);
xor U1714 (N_1714,N_948,N_951);
or U1715 (N_1715,N_429,N_204);
nor U1716 (N_1716,N_204,N_855);
xnor U1717 (N_1717,N_805,N_479);
and U1718 (N_1718,N_377,N_72);
and U1719 (N_1719,N_218,N_839);
or U1720 (N_1720,N_872,N_254);
or U1721 (N_1721,N_322,N_947);
and U1722 (N_1722,N_953,N_334);
nor U1723 (N_1723,N_889,N_80);
and U1724 (N_1724,N_902,N_700);
and U1725 (N_1725,N_875,N_109);
nor U1726 (N_1726,N_854,N_137);
and U1727 (N_1727,N_264,N_456);
nor U1728 (N_1728,N_694,N_590);
or U1729 (N_1729,N_321,N_575);
nand U1730 (N_1730,N_590,N_203);
or U1731 (N_1731,N_195,N_14);
or U1732 (N_1732,N_400,N_809);
xor U1733 (N_1733,N_737,N_35);
and U1734 (N_1734,N_239,N_998);
nand U1735 (N_1735,N_756,N_901);
or U1736 (N_1736,N_72,N_264);
nor U1737 (N_1737,N_730,N_234);
nand U1738 (N_1738,N_456,N_110);
nor U1739 (N_1739,N_150,N_838);
nand U1740 (N_1740,N_969,N_153);
nand U1741 (N_1741,N_91,N_258);
or U1742 (N_1742,N_238,N_798);
nor U1743 (N_1743,N_73,N_114);
xnor U1744 (N_1744,N_168,N_449);
nor U1745 (N_1745,N_530,N_709);
or U1746 (N_1746,N_616,N_410);
and U1747 (N_1747,N_398,N_358);
nor U1748 (N_1748,N_966,N_128);
xor U1749 (N_1749,N_568,N_464);
and U1750 (N_1750,N_708,N_289);
xor U1751 (N_1751,N_539,N_266);
or U1752 (N_1752,N_323,N_298);
and U1753 (N_1753,N_814,N_598);
and U1754 (N_1754,N_41,N_425);
or U1755 (N_1755,N_270,N_797);
and U1756 (N_1756,N_434,N_771);
and U1757 (N_1757,N_293,N_546);
and U1758 (N_1758,N_707,N_793);
nor U1759 (N_1759,N_963,N_495);
and U1760 (N_1760,N_903,N_211);
and U1761 (N_1761,N_93,N_360);
nor U1762 (N_1762,N_994,N_141);
and U1763 (N_1763,N_225,N_787);
nor U1764 (N_1764,N_932,N_149);
or U1765 (N_1765,N_841,N_228);
or U1766 (N_1766,N_453,N_852);
nand U1767 (N_1767,N_275,N_679);
or U1768 (N_1768,N_398,N_220);
and U1769 (N_1769,N_303,N_486);
nand U1770 (N_1770,N_617,N_107);
and U1771 (N_1771,N_737,N_359);
nor U1772 (N_1772,N_100,N_990);
nor U1773 (N_1773,N_32,N_99);
nand U1774 (N_1774,N_825,N_739);
and U1775 (N_1775,N_254,N_946);
xor U1776 (N_1776,N_923,N_621);
nand U1777 (N_1777,N_342,N_973);
and U1778 (N_1778,N_536,N_515);
or U1779 (N_1779,N_59,N_36);
xnor U1780 (N_1780,N_739,N_711);
nand U1781 (N_1781,N_780,N_634);
nand U1782 (N_1782,N_272,N_785);
nand U1783 (N_1783,N_128,N_993);
and U1784 (N_1784,N_194,N_797);
xor U1785 (N_1785,N_595,N_608);
nand U1786 (N_1786,N_66,N_408);
xor U1787 (N_1787,N_899,N_953);
and U1788 (N_1788,N_258,N_493);
or U1789 (N_1789,N_651,N_150);
xnor U1790 (N_1790,N_164,N_28);
nand U1791 (N_1791,N_997,N_910);
or U1792 (N_1792,N_862,N_993);
or U1793 (N_1793,N_547,N_394);
and U1794 (N_1794,N_498,N_497);
xor U1795 (N_1795,N_689,N_943);
nand U1796 (N_1796,N_856,N_589);
nand U1797 (N_1797,N_935,N_822);
nor U1798 (N_1798,N_361,N_230);
nor U1799 (N_1799,N_737,N_870);
or U1800 (N_1800,N_745,N_71);
nand U1801 (N_1801,N_675,N_299);
or U1802 (N_1802,N_694,N_473);
or U1803 (N_1803,N_832,N_969);
nor U1804 (N_1804,N_444,N_154);
nand U1805 (N_1805,N_956,N_498);
and U1806 (N_1806,N_472,N_651);
xor U1807 (N_1807,N_609,N_545);
or U1808 (N_1808,N_112,N_778);
or U1809 (N_1809,N_532,N_71);
nor U1810 (N_1810,N_307,N_218);
and U1811 (N_1811,N_285,N_625);
and U1812 (N_1812,N_502,N_342);
nand U1813 (N_1813,N_543,N_395);
and U1814 (N_1814,N_889,N_579);
nand U1815 (N_1815,N_656,N_352);
nor U1816 (N_1816,N_764,N_81);
nor U1817 (N_1817,N_561,N_208);
nor U1818 (N_1818,N_150,N_757);
or U1819 (N_1819,N_490,N_348);
xor U1820 (N_1820,N_255,N_487);
nor U1821 (N_1821,N_205,N_344);
or U1822 (N_1822,N_208,N_778);
and U1823 (N_1823,N_4,N_124);
nand U1824 (N_1824,N_713,N_447);
xnor U1825 (N_1825,N_455,N_49);
and U1826 (N_1826,N_791,N_156);
or U1827 (N_1827,N_675,N_886);
nand U1828 (N_1828,N_435,N_129);
xnor U1829 (N_1829,N_31,N_938);
nand U1830 (N_1830,N_903,N_142);
nor U1831 (N_1831,N_410,N_233);
xnor U1832 (N_1832,N_523,N_675);
and U1833 (N_1833,N_694,N_739);
or U1834 (N_1834,N_727,N_840);
or U1835 (N_1835,N_748,N_733);
xnor U1836 (N_1836,N_29,N_163);
nand U1837 (N_1837,N_979,N_196);
and U1838 (N_1838,N_472,N_284);
xnor U1839 (N_1839,N_972,N_120);
xor U1840 (N_1840,N_942,N_127);
or U1841 (N_1841,N_512,N_53);
nand U1842 (N_1842,N_725,N_372);
or U1843 (N_1843,N_36,N_875);
and U1844 (N_1844,N_667,N_592);
xor U1845 (N_1845,N_97,N_852);
and U1846 (N_1846,N_848,N_14);
and U1847 (N_1847,N_85,N_726);
nand U1848 (N_1848,N_206,N_890);
nor U1849 (N_1849,N_3,N_65);
nor U1850 (N_1850,N_510,N_357);
nand U1851 (N_1851,N_617,N_383);
nor U1852 (N_1852,N_762,N_123);
and U1853 (N_1853,N_898,N_61);
and U1854 (N_1854,N_458,N_720);
nand U1855 (N_1855,N_650,N_23);
nor U1856 (N_1856,N_226,N_19);
and U1857 (N_1857,N_942,N_673);
and U1858 (N_1858,N_2,N_462);
nand U1859 (N_1859,N_483,N_595);
nand U1860 (N_1860,N_315,N_619);
nor U1861 (N_1861,N_3,N_415);
nand U1862 (N_1862,N_830,N_977);
or U1863 (N_1863,N_738,N_446);
xor U1864 (N_1864,N_892,N_278);
or U1865 (N_1865,N_401,N_420);
nand U1866 (N_1866,N_51,N_638);
or U1867 (N_1867,N_47,N_815);
xnor U1868 (N_1868,N_850,N_138);
or U1869 (N_1869,N_521,N_986);
and U1870 (N_1870,N_977,N_161);
nand U1871 (N_1871,N_544,N_51);
nor U1872 (N_1872,N_38,N_530);
nand U1873 (N_1873,N_90,N_123);
nor U1874 (N_1874,N_497,N_319);
or U1875 (N_1875,N_761,N_5);
nor U1876 (N_1876,N_31,N_679);
nand U1877 (N_1877,N_194,N_828);
nand U1878 (N_1878,N_556,N_236);
nand U1879 (N_1879,N_8,N_764);
nor U1880 (N_1880,N_706,N_144);
or U1881 (N_1881,N_867,N_685);
nand U1882 (N_1882,N_388,N_340);
nor U1883 (N_1883,N_636,N_380);
or U1884 (N_1884,N_358,N_590);
and U1885 (N_1885,N_925,N_534);
and U1886 (N_1886,N_575,N_16);
and U1887 (N_1887,N_179,N_278);
xnor U1888 (N_1888,N_603,N_854);
and U1889 (N_1889,N_310,N_545);
nand U1890 (N_1890,N_563,N_113);
or U1891 (N_1891,N_152,N_863);
or U1892 (N_1892,N_994,N_999);
nand U1893 (N_1893,N_368,N_212);
nand U1894 (N_1894,N_369,N_212);
nor U1895 (N_1895,N_827,N_15);
nand U1896 (N_1896,N_103,N_464);
nand U1897 (N_1897,N_391,N_963);
or U1898 (N_1898,N_576,N_365);
nand U1899 (N_1899,N_939,N_310);
and U1900 (N_1900,N_901,N_217);
or U1901 (N_1901,N_274,N_771);
nor U1902 (N_1902,N_835,N_669);
nand U1903 (N_1903,N_568,N_852);
and U1904 (N_1904,N_329,N_283);
or U1905 (N_1905,N_724,N_293);
or U1906 (N_1906,N_99,N_527);
and U1907 (N_1907,N_869,N_650);
or U1908 (N_1908,N_163,N_419);
nand U1909 (N_1909,N_103,N_158);
xor U1910 (N_1910,N_391,N_245);
or U1911 (N_1911,N_147,N_419);
nand U1912 (N_1912,N_218,N_442);
and U1913 (N_1913,N_935,N_162);
or U1914 (N_1914,N_727,N_454);
and U1915 (N_1915,N_352,N_120);
or U1916 (N_1916,N_150,N_577);
nor U1917 (N_1917,N_245,N_494);
or U1918 (N_1918,N_556,N_546);
and U1919 (N_1919,N_761,N_372);
nand U1920 (N_1920,N_601,N_646);
xnor U1921 (N_1921,N_250,N_430);
and U1922 (N_1922,N_509,N_290);
nor U1923 (N_1923,N_674,N_396);
and U1924 (N_1924,N_827,N_136);
nor U1925 (N_1925,N_827,N_169);
or U1926 (N_1926,N_546,N_543);
or U1927 (N_1927,N_913,N_909);
nand U1928 (N_1928,N_130,N_161);
nand U1929 (N_1929,N_146,N_610);
or U1930 (N_1930,N_795,N_373);
or U1931 (N_1931,N_30,N_730);
nand U1932 (N_1932,N_123,N_888);
nor U1933 (N_1933,N_751,N_829);
nand U1934 (N_1934,N_337,N_330);
or U1935 (N_1935,N_828,N_787);
or U1936 (N_1936,N_297,N_281);
or U1937 (N_1937,N_691,N_704);
nor U1938 (N_1938,N_721,N_345);
or U1939 (N_1939,N_606,N_855);
xor U1940 (N_1940,N_183,N_685);
xnor U1941 (N_1941,N_786,N_46);
or U1942 (N_1942,N_524,N_260);
nand U1943 (N_1943,N_393,N_36);
nor U1944 (N_1944,N_907,N_187);
or U1945 (N_1945,N_909,N_450);
xnor U1946 (N_1946,N_94,N_352);
xnor U1947 (N_1947,N_863,N_559);
nand U1948 (N_1948,N_266,N_315);
and U1949 (N_1949,N_859,N_129);
and U1950 (N_1950,N_257,N_865);
nand U1951 (N_1951,N_527,N_781);
and U1952 (N_1952,N_735,N_880);
nor U1953 (N_1953,N_392,N_671);
nand U1954 (N_1954,N_46,N_860);
and U1955 (N_1955,N_139,N_523);
nor U1956 (N_1956,N_466,N_502);
nand U1957 (N_1957,N_738,N_987);
xnor U1958 (N_1958,N_88,N_25);
nor U1959 (N_1959,N_840,N_432);
and U1960 (N_1960,N_367,N_459);
nand U1961 (N_1961,N_461,N_955);
nand U1962 (N_1962,N_163,N_259);
nor U1963 (N_1963,N_950,N_768);
nand U1964 (N_1964,N_491,N_490);
nand U1965 (N_1965,N_443,N_911);
nor U1966 (N_1966,N_900,N_662);
nand U1967 (N_1967,N_519,N_196);
or U1968 (N_1968,N_76,N_479);
or U1969 (N_1969,N_327,N_326);
nand U1970 (N_1970,N_443,N_419);
nand U1971 (N_1971,N_50,N_810);
nand U1972 (N_1972,N_509,N_200);
and U1973 (N_1973,N_536,N_841);
or U1974 (N_1974,N_559,N_994);
nand U1975 (N_1975,N_296,N_716);
xor U1976 (N_1976,N_13,N_89);
nand U1977 (N_1977,N_609,N_221);
or U1978 (N_1978,N_556,N_135);
nand U1979 (N_1979,N_726,N_383);
and U1980 (N_1980,N_560,N_967);
nor U1981 (N_1981,N_341,N_973);
xnor U1982 (N_1982,N_639,N_491);
nor U1983 (N_1983,N_603,N_411);
nor U1984 (N_1984,N_315,N_92);
and U1985 (N_1985,N_572,N_520);
and U1986 (N_1986,N_640,N_651);
xor U1987 (N_1987,N_639,N_3);
or U1988 (N_1988,N_73,N_773);
or U1989 (N_1989,N_156,N_131);
nor U1990 (N_1990,N_370,N_509);
nand U1991 (N_1991,N_620,N_663);
nor U1992 (N_1992,N_984,N_563);
nand U1993 (N_1993,N_774,N_486);
nor U1994 (N_1994,N_844,N_225);
nor U1995 (N_1995,N_919,N_261);
nor U1996 (N_1996,N_861,N_427);
xor U1997 (N_1997,N_20,N_999);
nor U1998 (N_1998,N_450,N_3);
or U1999 (N_1999,N_681,N_305);
xor U2000 (N_2000,N_1863,N_1041);
or U2001 (N_2001,N_1764,N_1837);
nor U2002 (N_2002,N_1016,N_1752);
and U2003 (N_2003,N_1651,N_1091);
nor U2004 (N_2004,N_1670,N_1613);
or U2005 (N_2005,N_1423,N_1065);
nand U2006 (N_2006,N_1482,N_1384);
xor U2007 (N_2007,N_1378,N_1108);
and U2008 (N_2008,N_1832,N_1687);
and U2009 (N_2009,N_1516,N_1821);
nand U2010 (N_2010,N_1351,N_1424);
or U2011 (N_2011,N_1481,N_1627);
nand U2012 (N_2012,N_1930,N_1553);
nand U2013 (N_2013,N_1509,N_1330);
nor U2014 (N_2014,N_1508,N_1476);
and U2015 (N_2015,N_1845,N_1013);
and U2016 (N_2016,N_1021,N_1409);
nor U2017 (N_2017,N_1878,N_1223);
or U2018 (N_2018,N_1083,N_1831);
and U2019 (N_2019,N_1357,N_1211);
and U2020 (N_2020,N_1625,N_1214);
nor U2021 (N_2021,N_1182,N_1253);
and U2022 (N_2022,N_1990,N_1734);
and U2023 (N_2023,N_1779,N_1800);
or U2024 (N_2024,N_1790,N_1912);
or U2025 (N_2025,N_1344,N_1604);
and U2026 (N_2026,N_1166,N_1979);
and U2027 (N_2027,N_1588,N_1009);
nand U2028 (N_2028,N_1871,N_1581);
and U2029 (N_2029,N_1289,N_1291);
nand U2030 (N_2030,N_1269,N_1197);
or U2031 (N_2031,N_1266,N_1228);
xnor U2032 (N_2032,N_1319,N_1071);
nand U2033 (N_2033,N_1006,N_1402);
or U2034 (N_2034,N_1763,N_1203);
nor U2035 (N_2035,N_1964,N_1154);
xnor U2036 (N_2036,N_1600,N_1052);
and U2037 (N_2037,N_1852,N_1786);
xor U2038 (N_2038,N_1237,N_1301);
nand U2039 (N_2039,N_1726,N_1561);
nand U2040 (N_2040,N_1709,N_1717);
or U2041 (N_2041,N_1498,N_1787);
nand U2042 (N_2042,N_1865,N_1032);
nor U2043 (N_2043,N_1989,N_1418);
nand U2044 (N_2044,N_1387,N_1112);
and U2045 (N_2045,N_1707,N_1278);
and U2046 (N_2046,N_1365,N_1967);
and U2047 (N_2047,N_1288,N_1132);
and U2048 (N_2048,N_1973,N_1860);
nor U2049 (N_2049,N_1873,N_1927);
nor U2050 (N_2050,N_1320,N_1754);
nand U2051 (N_2051,N_1459,N_1363);
nand U2052 (N_2052,N_1596,N_1685);
and U2053 (N_2053,N_1829,N_1222);
and U2054 (N_2054,N_1673,N_1130);
nor U2055 (N_2055,N_1444,N_1060);
nand U2056 (N_2056,N_1161,N_1123);
and U2057 (N_2057,N_1259,N_1885);
nand U2058 (N_2058,N_1172,N_1514);
nand U2059 (N_2059,N_1759,N_1274);
nor U2060 (N_2060,N_1827,N_1235);
nand U2061 (N_2061,N_1024,N_1640);
or U2062 (N_2062,N_1910,N_1567);
nor U2063 (N_2063,N_1290,N_1408);
and U2064 (N_2064,N_1252,N_1884);
or U2065 (N_2065,N_1391,N_1814);
xor U2066 (N_2066,N_1251,N_1750);
or U2067 (N_2067,N_1544,N_1436);
xor U2068 (N_2068,N_1120,N_1028);
or U2069 (N_2069,N_1245,N_1807);
nand U2070 (N_2070,N_1057,N_1719);
nand U2071 (N_2071,N_1072,N_1614);
and U2072 (N_2072,N_1026,N_1883);
xnor U2073 (N_2073,N_1683,N_1977);
or U2074 (N_2074,N_1318,N_1943);
and U2075 (N_2075,N_1043,N_1417);
and U2076 (N_2076,N_1522,N_1577);
nor U2077 (N_2077,N_1535,N_1103);
or U2078 (N_2078,N_1901,N_1102);
and U2079 (N_2079,N_1493,N_1899);
or U2080 (N_2080,N_1062,N_1796);
nand U2081 (N_2081,N_1087,N_1322);
nor U2082 (N_2082,N_1637,N_1386);
and U2083 (N_2083,N_1333,N_1358);
nor U2084 (N_2084,N_1563,N_1044);
nor U2085 (N_2085,N_1618,N_1745);
nand U2086 (N_2086,N_1480,N_1519);
nor U2087 (N_2087,N_1904,N_1657);
or U2088 (N_2088,N_1746,N_1847);
and U2089 (N_2089,N_1128,N_1226);
or U2090 (N_2090,N_1833,N_1601);
nor U2091 (N_2091,N_1089,N_1830);
or U2092 (N_2092,N_1215,N_1762);
nand U2093 (N_2093,N_1986,N_1810);
nor U2094 (N_2094,N_1435,N_1525);
nand U2095 (N_2095,N_1623,N_1820);
nor U2096 (N_2096,N_1373,N_1031);
nand U2097 (N_2097,N_1771,N_1502);
nor U2098 (N_2098,N_1097,N_1099);
or U2099 (N_2099,N_1620,N_1335);
nor U2100 (N_2100,N_1850,N_1282);
xor U2101 (N_2101,N_1433,N_1573);
xnor U2102 (N_2102,N_1708,N_1729);
or U2103 (N_2103,N_1954,N_1149);
nand U2104 (N_2104,N_1626,N_1109);
and U2105 (N_2105,N_1504,N_1490);
xor U2106 (N_2106,N_1926,N_1570);
nand U2107 (N_2107,N_1050,N_1711);
or U2108 (N_2108,N_1950,N_1115);
nand U2109 (N_2109,N_1700,N_1915);
and U2110 (N_2110,N_1732,N_1841);
nand U2111 (N_2111,N_1201,N_1395);
and U2112 (N_2112,N_1866,N_1280);
xnor U2113 (N_2113,N_1248,N_1793);
or U2114 (N_2114,N_1994,N_1054);
or U2115 (N_2115,N_1145,N_1969);
or U2116 (N_2116,N_1876,N_1879);
and U2117 (N_2117,N_1710,N_1157);
xnor U2118 (N_2118,N_1377,N_1985);
nor U2119 (N_2119,N_1350,N_1388);
nand U2120 (N_2120,N_1527,N_1208);
nand U2121 (N_2121,N_1869,N_1010);
nand U2122 (N_2122,N_1716,N_1467);
or U2123 (N_2123,N_1944,N_1162);
nand U2124 (N_2124,N_1469,N_1422);
nand U2125 (N_2125,N_1066,N_1250);
xnor U2126 (N_2126,N_1738,N_1174);
nor U2127 (N_2127,N_1919,N_1339);
nor U2128 (N_2128,N_1501,N_1606);
or U2129 (N_2129,N_1325,N_1594);
nor U2130 (N_2130,N_1720,N_1406);
nor U2131 (N_2131,N_1015,N_1554);
nand U2132 (N_2132,N_1894,N_1156);
and U2133 (N_2133,N_1767,N_1928);
and U2134 (N_2134,N_1880,N_1652);
and U2135 (N_2135,N_1835,N_1073);
nand U2136 (N_2136,N_1101,N_1534);
or U2137 (N_2137,N_1539,N_1536);
nand U2138 (N_2138,N_1564,N_1968);
nor U2139 (N_2139,N_1124,N_1499);
nor U2140 (N_2140,N_1586,N_1692);
or U2141 (N_2141,N_1633,N_1017);
and U2142 (N_2142,N_1659,N_1077);
or U2143 (N_2143,N_1664,N_1788);
nand U2144 (N_2144,N_1440,N_1857);
nor U2145 (N_2145,N_1797,N_1029);
nand U2146 (N_2146,N_1486,N_1188);
and U2147 (N_2147,N_1524,N_1941);
or U2148 (N_2148,N_1047,N_1439);
nand U2149 (N_2149,N_1119,N_1287);
nor U2150 (N_2150,N_1371,N_1195);
nand U2151 (N_2151,N_1328,N_1261);
and U2152 (N_2152,N_1457,N_1945);
or U2153 (N_2153,N_1234,N_1911);
and U2154 (N_2154,N_1048,N_1728);
nor U2155 (N_2155,N_1589,N_1960);
nand U2156 (N_2156,N_1428,N_1765);
nand U2157 (N_2157,N_1809,N_1681);
nor U2158 (N_2158,N_1714,N_1667);
nand U2159 (N_2159,N_1909,N_1741);
nor U2160 (N_2160,N_1547,N_1111);
nor U2161 (N_2161,N_1961,N_1191);
nor U2162 (N_2162,N_1691,N_1742);
nand U2163 (N_2163,N_1263,N_1920);
and U2164 (N_2164,N_1264,N_1560);
nand U2165 (N_2165,N_1432,N_1137);
and U2166 (N_2166,N_1022,N_1329);
nand U2167 (N_2167,N_1931,N_1996);
nand U2168 (N_2168,N_1987,N_1584);
nor U2169 (N_2169,N_1170,N_1727);
or U2170 (N_2170,N_1038,N_1760);
or U2171 (N_2171,N_1310,N_1503);
nand U2172 (N_2172,N_1982,N_1689);
nand U2173 (N_2173,N_1296,N_1220);
nor U2174 (N_2174,N_1792,N_1549);
nand U2175 (N_2175,N_1348,N_1705);
or U2176 (N_2176,N_1557,N_1020);
and U2177 (N_2177,N_1874,N_1193);
nor U2178 (N_2178,N_1908,N_1891);
nor U2179 (N_2179,N_1221,N_1352);
or U2180 (N_2180,N_1970,N_1392);
nor U2181 (N_2181,N_1389,N_1336);
nor U2182 (N_2182,N_1654,N_1974);
and U2183 (N_2183,N_1933,N_1247);
nor U2184 (N_2184,N_1362,N_1815);
and U2185 (N_2185,N_1064,N_1270);
and U2186 (N_2186,N_1634,N_1403);
and U2187 (N_2187,N_1401,N_1802);
and U2188 (N_2188,N_1587,N_1962);
or U2189 (N_2189,N_1311,N_1458);
and U2190 (N_2190,N_1569,N_1307);
or U2191 (N_2191,N_1992,N_1199);
nor U2192 (N_2192,N_1558,N_1998);
and U2193 (N_2193,N_1396,N_1308);
or U2194 (N_2194,N_1256,N_1817);
nor U2195 (N_2195,N_1593,N_1345);
nand U2196 (N_2196,N_1168,N_1441);
nand U2197 (N_2197,N_1924,N_1114);
nor U2198 (N_2198,N_1513,N_1599);
nor U2199 (N_2199,N_1794,N_1079);
xnor U2200 (N_2200,N_1971,N_1862);
nor U2201 (N_2201,N_1347,N_1437);
nor U2202 (N_2202,N_1725,N_1046);
nor U2203 (N_2203,N_1090,N_1138);
and U2204 (N_2204,N_1552,N_1948);
nor U2205 (N_2205,N_1636,N_1551);
and U2206 (N_2206,N_1698,N_1421);
nor U2207 (N_2207,N_1206,N_1903);
nor U2208 (N_2208,N_1317,N_1148);
nand U2209 (N_2209,N_1446,N_1327);
and U2210 (N_2210,N_1142,N_1812);
or U2211 (N_2211,N_1394,N_1184);
and U2212 (N_2212,N_1475,N_1216);
nand U2213 (N_2213,N_1740,N_1828);
or U2214 (N_2214,N_1976,N_1202);
and U2215 (N_2215,N_1495,N_1382);
or U2216 (N_2216,N_1292,N_1438);
and U2217 (N_2217,N_1568,N_1559);
or U2218 (N_2218,N_1429,N_1121);
or U2219 (N_2219,N_1379,N_1823);
nor U2220 (N_2220,N_1597,N_1611);
nand U2221 (N_2221,N_1929,N_1783);
nand U2222 (N_2222,N_1003,N_1163);
nand U2223 (N_2223,N_1694,N_1940);
nor U2224 (N_2224,N_1743,N_1074);
nor U2225 (N_2225,N_1095,N_1477);
nor U2226 (N_2226,N_1294,N_1556);
nand U2227 (N_2227,N_1646,N_1521);
and U2228 (N_2228,N_1360,N_1639);
nor U2229 (N_2229,N_1081,N_1037);
nor U2230 (N_2230,N_1663,N_1179);
or U2231 (N_2231,N_1136,N_1981);
nor U2232 (N_2232,N_1285,N_1466);
or U2233 (N_2233,N_1398,N_1368);
nand U2234 (N_2234,N_1096,N_1537);
nand U2235 (N_2235,N_1231,N_1949);
or U2236 (N_2236,N_1795,N_1260);
nor U2237 (N_2237,N_1025,N_1619);
nand U2238 (N_2238,N_1205,N_1002);
nand U2239 (N_2239,N_1085,N_1431);
nor U2240 (N_2240,N_1106,N_1590);
nor U2241 (N_2241,N_1622,N_1739);
nand U2242 (N_2242,N_1736,N_1712);
nand U2243 (N_2243,N_1785,N_1164);
nand U2244 (N_2244,N_1907,N_1230);
nand U2245 (N_2245,N_1775,N_1917);
or U2246 (N_2246,N_1846,N_1861);
nand U2247 (N_2247,N_1592,N_1133);
or U2248 (N_2248,N_1479,N_1848);
nor U2249 (N_2249,N_1000,N_1737);
nand U2250 (N_2250,N_1233,N_1877);
and U2251 (N_2251,N_1058,N_1733);
or U2252 (N_2252,N_1147,N_1171);
nor U2253 (N_2253,N_1608,N_1520);
and U2254 (N_2254,N_1454,N_1213);
xnor U2255 (N_2255,N_1343,N_1151);
nand U2256 (N_2256,N_1882,N_1238);
or U2257 (N_2257,N_1204,N_1655);
nand U2258 (N_2258,N_1178,N_1975);
nor U2259 (N_2259,N_1631,N_1104);
and U2260 (N_2260,N_1621,N_1442);
and U2261 (N_2261,N_1784,N_1789);
nand U2262 (N_2262,N_1956,N_1190);
or U2263 (N_2263,N_1781,N_1898);
and U2264 (N_2264,N_1375,N_1366);
and U2265 (N_2265,N_1067,N_1946);
nor U2266 (N_2266,N_1840,N_1316);
or U2267 (N_2267,N_1565,N_1959);
nor U2268 (N_2268,N_1407,N_1932);
nand U2269 (N_2269,N_1942,N_1571);
and U2270 (N_2270,N_1735,N_1851);
or U2271 (N_2271,N_1897,N_1751);
and U2272 (N_2272,N_1843,N_1413);
or U2273 (N_2273,N_1094,N_1488);
nand U2274 (N_2274,N_1704,N_1724);
and U2275 (N_2275,N_1925,N_1131);
and U2276 (N_2276,N_1540,N_1049);
nand U2277 (N_2277,N_1984,N_1696);
nand U2278 (N_2278,N_1334,N_1666);
or U2279 (N_2279,N_1240,N_1453);
and U2280 (N_2280,N_1872,N_1011);
nand U2281 (N_2281,N_1239,N_1465);
nor U2282 (N_2282,N_1279,N_1092);
xnor U2283 (N_2283,N_1224,N_1780);
or U2284 (N_2284,N_1965,N_1776);
xor U2285 (N_2285,N_1675,N_1957);
nor U2286 (N_2286,N_1669,N_1098);
and U2287 (N_2287,N_1913,N_1210);
and U2288 (N_2288,N_1517,N_1298);
or U2289 (N_2289,N_1053,N_1511);
nor U2290 (N_2290,N_1483,N_1273);
and U2291 (N_2291,N_1181,N_1721);
or U2292 (N_2292,N_1257,N_1773);
xnor U2293 (N_2293,N_1277,N_1472);
and U2294 (N_2294,N_1566,N_1027);
nand U2295 (N_2295,N_1005,N_1275);
nand U2296 (N_2296,N_1905,N_1088);
and U2297 (N_2297,N_1854,N_1546);
and U2298 (N_2298,N_1699,N_1629);
or U2299 (N_2299,N_1595,N_1855);
and U2300 (N_2300,N_1411,N_1447);
and U2301 (N_2301,N_1598,N_1532);
nand U2302 (N_2302,N_1198,N_1951);
xor U2303 (N_2303,N_1448,N_1135);
nand U2304 (N_2304,N_1864,N_1212);
or U2305 (N_2305,N_1701,N_1575);
and U2306 (N_2306,N_1338,N_1955);
nand U2307 (N_2307,N_1243,N_1471);
or U2308 (N_2308,N_1150,N_1755);
nand U2309 (N_2309,N_1660,N_1232);
nand U2310 (N_2310,N_1947,N_1326);
nand U2311 (N_2311,N_1196,N_1676);
or U2312 (N_2312,N_1747,N_1452);
and U2313 (N_2313,N_1550,N_1420);
and U2314 (N_2314,N_1176,N_1018);
nor U2315 (N_2315,N_1769,N_1314);
nand U2316 (N_2316,N_1070,N_1693);
and U2317 (N_2317,N_1649,N_1342);
and U2318 (N_2318,N_1890,N_1507);
nand U2319 (N_2319,N_1555,N_1404);
or U2320 (N_2320,N_1093,N_1055);
and U2321 (N_2321,N_1591,N_1510);
xnor U2322 (N_2322,N_1836,N_1680);
and U2323 (N_2323,N_1068,N_1116);
and U2324 (N_2324,N_1768,N_1798);
and U2325 (N_2325,N_1144,N_1080);
nand U2326 (N_2326,N_1679,N_1141);
or U2327 (N_2327,N_1538,N_1194);
and U2328 (N_2328,N_1023,N_1935);
or U2329 (N_2329,N_1642,N_1084);
or U2330 (N_2330,N_1372,N_1997);
and U2331 (N_2331,N_1332,N_1478);
nand U2332 (N_2332,N_1671,N_1125);
nand U2333 (N_2333,N_1803,N_1939);
xnor U2334 (N_2334,N_1474,N_1265);
nor U2335 (N_2335,N_1173,N_1610);
and U2336 (N_2336,N_1051,N_1868);
nor U2337 (N_2337,N_1906,N_1999);
nand U2338 (N_2338,N_1648,N_1934);
nor U2339 (N_2339,N_1293,N_1331);
nand U2340 (N_2340,N_1470,N_1295);
nor U2341 (N_2341,N_1460,N_1838);
or U2342 (N_2342,N_1246,N_1778);
nor U2343 (N_2343,N_1530,N_1019);
or U2344 (N_2344,N_1430,N_1451);
xnor U2345 (N_2345,N_1272,N_1122);
and U2346 (N_2346,N_1219,N_1304);
nor U2347 (N_2347,N_1826,N_1127);
or U2348 (N_2348,N_1952,N_1881);
nor U2349 (N_2349,N_1461,N_1918);
and U2350 (N_2350,N_1677,N_1405);
nor U2351 (N_2351,N_1152,N_1140);
nand U2352 (N_2352,N_1443,N_1662);
nand U2353 (N_2353,N_1818,N_1574);
and U2354 (N_2354,N_1034,N_1076);
or U2355 (N_2355,N_1390,N_1545);
nor U2356 (N_2356,N_1217,N_1464);
nor U2357 (N_2357,N_1886,N_1991);
or U2358 (N_2358,N_1346,N_1192);
and U2359 (N_2359,N_1922,N_1518);
and U2360 (N_2360,N_1858,N_1412);
xor U2361 (N_2361,N_1489,N_1853);
xor U2362 (N_2362,N_1007,N_1374);
nand U2363 (N_2363,N_1731,N_1229);
or U2364 (N_2364,N_1983,N_1808);
nor U2365 (N_2365,N_1271,N_1533);
nand U2366 (N_2366,N_1582,N_1766);
or U2367 (N_2367,N_1806,N_1207);
nor U2368 (N_2368,N_1572,N_1782);
and U2369 (N_2369,N_1936,N_1494);
or U2370 (N_2370,N_1523,N_1040);
nand U2371 (N_2371,N_1463,N_1889);
and U2372 (N_2372,N_1241,N_1528);
nand U2373 (N_2373,N_1980,N_1585);
or U2374 (N_2374,N_1155,N_1001);
nor U2375 (N_2375,N_1605,N_1867);
nor U2376 (N_2376,N_1169,N_1644);
and U2377 (N_2377,N_1356,N_1487);
xor U2378 (N_2378,N_1895,N_1035);
nand U2379 (N_2379,N_1813,N_1761);
nand U2380 (N_2380,N_1300,N_1526);
nor U2381 (N_2381,N_1856,N_1512);
nand U2382 (N_2382,N_1146,N_1086);
nor U2383 (N_2383,N_1607,N_1126);
and U2384 (N_2384,N_1110,N_1938);
and U2385 (N_2385,N_1609,N_1297);
or U2386 (N_2386,N_1628,N_1069);
nand U2387 (N_2387,N_1914,N_1748);
or U2388 (N_2388,N_1383,N_1129);
or U2389 (N_2389,N_1160,N_1749);
and U2390 (N_2390,N_1937,N_1177);
nor U2391 (N_2391,N_1658,N_1500);
and U2392 (N_2392,N_1183,N_1225);
nand U2393 (N_2393,N_1875,N_1686);
or U2394 (N_2394,N_1697,N_1118);
or U2395 (N_2395,N_1834,N_1972);
nor U2396 (N_2396,N_1449,N_1399);
nor U2397 (N_2397,N_1236,N_1218);
nand U2398 (N_2398,N_1647,N_1723);
nor U2399 (N_2399,N_1030,N_1653);
nand U2400 (N_2400,N_1603,N_1036);
nand U2401 (N_2401,N_1617,N_1753);
nand U2402 (N_2402,N_1187,N_1059);
nand U2403 (N_2403,N_1995,N_1988);
or U2404 (N_2404,N_1615,N_1324);
or U2405 (N_2405,N_1337,N_1180);
or U2406 (N_2406,N_1299,N_1576);
nor U2407 (N_2407,N_1805,N_1715);
nor U2408 (N_2408,N_1276,N_1822);
and U2409 (N_2409,N_1113,N_1900);
or U2410 (N_2410,N_1529,N_1923);
or U2411 (N_2411,N_1167,N_1774);
xnor U2412 (N_2412,N_1004,N_1284);
and U2413 (N_2413,N_1381,N_1713);
and U2414 (N_2414,N_1415,N_1730);
nand U2415 (N_2415,N_1770,N_1963);
or U2416 (N_2416,N_1485,N_1665);
nor U2417 (N_2417,N_1249,N_1758);
nor U2418 (N_2418,N_1416,N_1650);
nor U2419 (N_2419,N_1376,N_1811);
and U2420 (N_2420,N_1757,N_1313);
nand U2421 (N_2421,N_1638,N_1117);
or U2422 (N_2422,N_1953,N_1254);
nand U2423 (N_2423,N_1075,N_1369);
nor U2424 (N_2424,N_1893,N_1824);
or U2425 (N_2425,N_1258,N_1801);
nor U2426 (N_2426,N_1283,N_1888);
nand U2427 (N_2427,N_1777,N_1309);
nor U2428 (N_2428,N_1242,N_1531);
and U2429 (N_2429,N_1370,N_1839);
or U2430 (N_2430,N_1426,N_1042);
nor U2431 (N_2431,N_1039,N_1656);
nor U2432 (N_2432,N_1303,N_1816);
or U2433 (N_2433,N_1340,N_1185);
and U2434 (N_2434,N_1542,N_1578);
and U2435 (N_2435,N_1842,N_1008);
nand U2436 (N_2436,N_1722,N_1302);
or U2437 (N_2437,N_1354,N_1012);
nor U2438 (N_2438,N_1690,N_1804);
nor U2439 (N_2439,N_1966,N_1543);
and U2440 (N_2440,N_1364,N_1756);
and U2441 (N_2441,N_1419,N_1455);
and U2442 (N_2442,N_1158,N_1393);
and U2443 (N_2443,N_1014,N_1462);
or U2444 (N_2444,N_1791,N_1958);
nor U2445 (N_2445,N_1427,N_1630);
nand U2446 (N_2446,N_1844,N_1562);
and U2447 (N_2447,N_1921,N_1580);
nor U2448 (N_2448,N_1643,N_1414);
or U2449 (N_2449,N_1255,N_1143);
nor U2450 (N_2450,N_1583,N_1492);
and U2451 (N_2451,N_1175,N_1668);
and U2452 (N_2452,N_1353,N_1772);
xnor U2453 (N_2453,N_1315,N_1916);
or U2454 (N_2454,N_1702,N_1703);
or U2455 (N_2455,N_1397,N_1200);
nor U2456 (N_2456,N_1641,N_1678);
xor U2457 (N_2457,N_1312,N_1892);
nand U2458 (N_2458,N_1870,N_1456);
and U2459 (N_2459,N_1159,N_1262);
nand U2460 (N_2460,N_1045,N_1267);
or U2461 (N_2461,N_1579,N_1849);
or U2462 (N_2462,N_1186,N_1902);
and U2463 (N_2463,N_1497,N_1410);
xnor U2464 (N_2464,N_1695,N_1107);
or U2465 (N_2465,N_1491,N_1268);
or U2466 (N_2466,N_1061,N_1359);
and U2467 (N_2467,N_1468,N_1367);
nor U2468 (N_2468,N_1744,N_1323);
nand U2469 (N_2469,N_1286,N_1684);
and U2470 (N_2470,N_1033,N_1859);
xor U2471 (N_2471,N_1819,N_1672);
nand U2472 (N_2472,N_1635,N_1993);
or U2473 (N_2473,N_1799,N_1134);
or U2474 (N_2474,N_1506,N_1645);
and U2475 (N_2475,N_1473,N_1349);
and U2476 (N_2476,N_1380,N_1505);
or U2477 (N_2477,N_1434,N_1887);
nand U2478 (N_2478,N_1189,N_1281);
xor U2479 (N_2479,N_1209,N_1305);
and U2480 (N_2480,N_1624,N_1632);
nand U2481 (N_2481,N_1450,N_1105);
and U2482 (N_2482,N_1361,N_1718);
nand U2483 (N_2483,N_1165,N_1445);
xnor U2484 (N_2484,N_1661,N_1400);
and U2485 (N_2485,N_1244,N_1385);
nor U2486 (N_2486,N_1548,N_1602);
nor U2487 (N_2487,N_1056,N_1978);
nand U2488 (N_2488,N_1425,N_1612);
or U2489 (N_2489,N_1825,N_1227);
nand U2490 (N_2490,N_1496,N_1139);
nor U2491 (N_2491,N_1896,N_1682);
nand U2492 (N_2492,N_1688,N_1306);
nand U2493 (N_2493,N_1341,N_1706);
nor U2494 (N_2494,N_1100,N_1484);
nor U2495 (N_2495,N_1541,N_1078);
and U2496 (N_2496,N_1321,N_1515);
and U2497 (N_2497,N_1153,N_1674);
and U2498 (N_2498,N_1616,N_1082);
or U2499 (N_2499,N_1063,N_1355);
or U2500 (N_2500,N_1604,N_1320);
or U2501 (N_2501,N_1278,N_1241);
xnor U2502 (N_2502,N_1381,N_1812);
nor U2503 (N_2503,N_1541,N_1776);
nand U2504 (N_2504,N_1366,N_1736);
or U2505 (N_2505,N_1069,N_1991);
nand U2506 (N_2506,N_1804,N_1581);
or U2507 (N_2507,N_1196,N_1633);
and U2508 (N_2508,N_1450,N_1985);
or U2509 (N_2509,N_1548,N_1536);
or U2510 (N_2510,N_1898,N_1003);
xnor U2511 (N_2511,N_1438,N_1098);
nor U2512 (N_2512,N_1266,N_1581);
nor U2513 (N_2513,N_1874,N_1843);
xnor U2514 (N_2514,N_1960,N_1237);
nand U2515 (N_2515,N_1910,N_1230);
or U2516 (N_2516,N_1237,N_1508);
nor U2517 (N_2517,N_1839,N_1301);
nand U2518 (N_2518,N_1986,N_1930);
or U2519 (N_2519,N_1389,N_1689);
or U2520 (N_2520,N_1718,N_1196);
and U2521 (N_2521,N_1443,N_1110);
or U2522 (N_2522,N_1520,N_1369);
and U2523 (N_2523,N_1284,N_1713);
or U2524 (N_2524,N_1551,N_1859);
and U2525 (N_2525,N_1690,N_1305);
xor U2526 (N_2526,N_1818,N_1816);
nand U2527 (N_2527,N_1204,N_1353);
nand U2528 (N_2528,N_1347,N_1075);
or U2529 (N_2529,N_1973,N_1901);
nand U2530 (N_2530,N_1127,N_1843);
and U2531 (N_2531,N_1431,N_1095);
or U2532 (N_2532,N_1881,N_1423);
nand U2533 (N_2533,N_1608,N_1248);
xor U2534 (N_2534,N_1624,N_1552);
or U2535 (N_2535,N_1701,N_1715);
nand U2536 (N_2536,N_1282,N_1953);
and U2537 (N_2537,N_1685,N_1416);
nor U2538 (N_2538,N_1540,N_1692);
nor U2539 (N_2539,N_1156,N_1747);
or U2540 (N_2540,N_1413,N_1217);
or U2541 (N_2541,N_1180,N_1868);
nor U2542 (N_2542,N_1835,N_1683);
or U2543 (N_2543,N_1903,N_1135);
or U2544 (N_2544,N_1625,N_1093);
and U2545 (N_2545,N_1693,N_1803);
nor U2546 (N_2546,N_1110,N_1701);
nand U2547 (N_2547,N_1541,N_1471);
xnor U2548 (N_2548,N_1289,N_1228);
nor U2549 (N_2549,N_1300,N_1705);
nand U2550 (N_2550,N_1115,N_1657);
and U2551 (N_2551,N_1861,N_1043);
nand U2552 (N_2552,N_1174,N_1708);
or U2553 (N_2553,N_1877,N_1372);
nand U2554 (N_2554,N_1202,N_1782);
nand U2555 (N_2555,N_1636,N_1994);
nand U2556 (N_2556,N_1082,N_1656);
nand U2557 (N_2557,N_1916,N_1105);
nor U2558 (N_2558,N_1202,N_1753);
nor U2559 (N_2559,N_1242,N_1961);
xnor U2560 (N_2560,N_1130,N_1346);
nor U2561 (N_2561,N_1556,N_1060);
and U2562 (N_2562,N_1424,N_1850);
or U2563 (N_2563,N_1191,N_1852);
nor U2564 (N_2564,N_1023,N_1469);
or U2565 (N_2565,N_1302,N_1956);
and U2566 (N_2566,N_1984,N_1913);
or U2567 (N_2567,N_1479,N_1486);
or U2568 (N_2568,N_1391,N_1880);
nand U2569 (N_2569,N_1109,N_1964);
nor U2570 (N_2570,N_1089,N_1953);
nor U2571 (N_2571,N_1121,N_1873);
nand U2572 (N_2572,N_1221,N_1629);
and U2573 (N_2573,N_1532,N_1010);
nand U2574 (N_2574,N_1753,N_1047);
and U2575 (N_2575,N_1440,N_1715);
nand U2576 (N_2576,N_1688,N_1913);
nand U2577 (N_2577,N_1609,N_1864);
nor U2578 (N_2578,N_1170,N_1532);
nor U2579 (N_2579,N_1398,N_1388);
and U2580 (N_2580,N_1959,N_1012);
nor U2581 (N_2581,N_1093,N_1004);
or U2582 (N_2582,N_1465,N_1336);
nand U2583 (N_2583,N_1931,N_1544);
nor U2584 (N_2584,N_1540,N_1284);
and U2585 (N_2585,N_1377,N_1817);
nand U2586 (N_2586,N_1166,N_1882);
nor U2587 (N_2587,N_1583,N_1331);
or U2588 (N_2588,N_1619,N_1526);
xnor U2589 (N_2589,N_1157,N_1780);
and U2590 (N_2590,N_1291,N_1764);
nor U2591 (N_2591,N_1215,N_1729);
or U2592 (N_2592,N_1709,N_1576);
nand U2593 (N_2593,N_1206,N_1358);
and U2594 (N_2594,N_1403,N_1362);
and U2595 (N_2595,N_1795,N_1985);
nor U2596 (N_2596,N_1042,N_1090);
or U2597 (N_2597,N_1171,N_1767);
and U2598 (N_2598,N_1316,N_1484);
nor U2599 (N_2599,N_1593,N_1346);
nor U2600 (N_2600,N_1429,N_1858);
xor U2601 (N_2601,N_1328,N_1296);
and U2602 (N_2602,N_1320,N_1777);
or U2603 (N_2603,N_1490,N_1962);
and U2604 (N_2604,N_1639,N_1701);
xor U2605 (N_2605,N_1818,N_1893);
and U2606 (N_2606,N_1514,N_1077);
and U2607 (N_2607,N_1662,N_1813);
nor U2608 (N_2608,N_1090,N_1368);
and U2609 (N_2609,N_1838,N_1306);
or U2610 (N_2610,N_1702,N_1110);
nor U2611 (N_2611,N_1101,N_1529);
nand U2612 (N_2612,N_1578,N_1330);
or U2613 (N_2613,N_1613,N_1878);
and U2614 (N_2614,N_1691,N_1390);
and U2615 (N_2615,N_1955,N_1433);
nand U2616 (N_2616,N_1150,N_1405);
xor U2617 (N_2617,N_1709,N_1313);
xnor U2618 (N_2618,N_1536,N_1259);
and U2619 (N_2619,N_1041,N_1396);
and U2620 (N_2620,N_1367,N_1371);
and U2621 (N_2621,N_1280,N_1787);
and U2622 (N_2622,N_1892,N_1039);
or U2623 (N_2623,N_1773,N_1512);
nand U2624 (N_2624,N_1546,N_1700);
nand U2625 (N_2625,N_1540,N_1999);
or U2626 (N_2626,N_1143,N_1909);
nor U2627 (N_2627,N_1328,N_1685);
and U2628 (N_2628,N_1993,N_1896);
nor U2629 (N_2629,N_1873,N_1366);
and U2630 (N_2630,N_1111,N_1123);
or U2631 (N_2631,N_1695,N_1271);
nand U2632 (N_2632,N_1614,N_1283);
xnor U2633 (N_2633,N_1869,N_1707);
or U2634 (N_2634,N_1162,N_1150);
and U2635 (N_2635,N_1252,N_1227);
and U2636 (N_2636,N_1492,N_1972);
or U2637 (N_2637,N_1349,N_1640);
or U2638 (N_2638,N_1490,N_1170);
xnor U2639 (N_2639,N_1768,N_1958);
nand U2640 (N_2640,N_1240,N_1606);
or U2641 (N_2641,N_1265,N_1890);
and U2642 (N_2642,N_1989,N_1498);
nor U2643 (N_2643,N_1273,N_1377);
nor U2644 (N_2644,N_1544,N_1169);
or U2645 (N_2645,N_1946,N_1355);
xor U2646 (N_2646,N_1809,N_1438);
nor U2647 (N_2647,N_1163,N_1335);
or U2648 (N_2648,N_1917,N_1815);
or U2649 (N_2649,N_1531,N_1661);
and U2650 (N_2650,N_1729,N_1832);
nand U2651 (N_2651,N_1768,N_1201);
xor U2652 (N_2652,N_1857,N_1445);
xor U2653 (N_2653,N_1281,N_1945);
or U2654 (N_2654,N_1678,N_1843);
nor U2655 (N_2655,N_1511,N_1699);
xnor U2656 (N_2656,N_1947,N_1618);
and U2657 (N_2657,N_1280,N_1432);
or U2658 (N_2658,N_1026,N_1817);
xnor U2659 (N_2659,N_1034,N_1388);
nor U2660 (N_2660,N_1558,N_1564);
nand U2661 (N_2661,N_1350,N_1994);
and U2662 (N_2662,N_1554,N_1002);
or U2663 (N_2663,N_1292,N_1784);
nor U2664 (N_2664,N_1447,N_1014);
or U2665 (N_2665,N_1258,N_1166);
xnor U2666 (N_2666,N_1049,N_1175);
and U2667 (N_2667,N_1772,N_1344);
nand U2668 (N_2668,N_1760,N_1020);
nor U2669 (N_2669,N_1683,N_1801);
or U2670 (N_2670,N_1894,N_1674);
and U2671 (N_2671,N_1417,N_1456);
and U2672 (N_2672,N_1217,N_1876);
nor U2673 (N_2673,N_1224,N_1971);
or U2674 (N_2674,N_1561,N_1248);
nor U2675 (N_2675,N_1816,N_1474);
and U2676 (N_2676,N_1225,N_1537);
nor U2677 (N_2677,N_1002,N_1808);
and U2678 (N_2678,N_1279,N_1433);
nand U2679 (N_2679,N_1324,N_1793);
nand U2680 (N_2680,N_1988,N_1723);
xnor U2681 (N_2681,N_1137,N_1112);
and U2682 (N_2682,N_1520,N_1746);
nor U2683 (N_2683,N_1495,N_1177);
or U2684 (N_2684,N_1336,N_1535);
xor U2685 (N_2685,N_1546,N_1098);
nor U2686 (N_2686,N_1114,N_1696);
and U2687 (N_2687,N_1053,N_1043);
and U2688 (N_2688,N_1471,N_1201);
nor U2689 (N_2689,N_1768,N_1206);
and U2690 (N_2690,N_1786,N_1187);
nand U2691 (N_2691,N_1162,N_1634);
nor U2692 (N_2692,N_1768,N_1727);
nor U2693 (N_2693,N_1564,N_1284);
or U2694 (N_2694,N_1402,N_1257);
or U2695 (N_2695,N_1209,N_1807);
or U2696 (N_2696,N_1210,N_1729);
and U2697 (N_2697,N_1751,N_1333);
nor U2698 (N_2698,N_1658,N_1236);
nor U2699 (N_2699,N_1262,N_1437);
and U2700 (N_2700,N_1712,N_1271);
nand U2701 (N_2701,N_1546,N_1978);
or U2702 (N_2702,N_1063,N_1681);
and U2703 (N_2703,N_1990,N_1420);
xor U2704 (N_2704,N_1100,N_1104);
nor U2705 (N_2705,N_1625,N_1847);
and U2706 (N_2706,N_1823,N_1189);
nand U2707 (N_2707,N_1582,N_1665);
xnor U2708 (N_2708,N_1900,N_1311);
xor U2709 (N_2709,N_1149,N_1913);
nand U2710 (N_2710,N_1678,N_1171);
and U2711 (N_2711,N_1461,N_1749);
xnor U2712 (N_2712,N_1710,N_1025);
nand U2713 (N_2713,N_1760,N_1731);
nor U2714 (N_2714,N_1926,N_1099);
nor U2715 (N_2715,N_1121,N_1152);
nand U2716 (N_2716,N_1131,N_1834);
nand U2717 (N_2717,N_1028,N_1952);
and U2718 (N_2718,N_1138,N_1814);
nand U2719 (N_2719,N_1370,N_1092);
nor U2720 (N_2720,N_1440,N_1680);
nor U2721 (N_2721,N_1610,N_1843);
nand U2722 (N_2722,N_1320,N_1061);
xor U2723 (N_2723,N_1795,N_1144);
or U2724 (N_2724,N_1696,N_1071);
nor U2725 (N_2725,N_1604,N_1514);
nor U2726 (N_2726,N_1136,N_1813);
nand U2727 (N_2727,N_1958,N_1059);
or U2728 (N_2728,N_1563,N_1274);
nand U2729 (N_2729,N_1516,N_1605);
or U2730 (N_2730,N_1097,N_1071);
nand U2731 (N_2731,N_1623,N_1519);
nor U2732 (N_2732,N_1153,N_1267);
xor U2733 (N_2733,N_1502,N_1836);
xnor U2734 (N_2734,N_1809,N_1192);
xor U2735 (N_2735,N_1852,N_1533);
xnor U2736 (N_2736,N_1010,N_1816);
or U2737 (N_2737,N_1703,N_1717);
nand U2738 (N_2738,N_1302,N_1418);
nand U2739 (N_2739,N_1068,N_1108);
xnor U2740 (N_2740,N_1583,N_1200);
and U2741 (N_2741,N_1130,N_1394);
and U2742 (N_2742,N_1801,N_1030);
or U2743 (N_2743,N_1247,N_1528);
nor U2744 (N_2744,N_1773,N_1551);
nand U2745 (N_2745,N_1528,N_1137);
or U2746 (N_2746,N_1903,N_1405);
nand U2747 (N_2747,N_1771,N_1870);
and U2748 (N_2748,N_1981,N_1971);
nand U2749 (N_2749,N_1872,N_1104);
nand U2750 (N_2750,N_1273,N_1631);
and U2751 (N_2751,N_1602,N_1080);
nor U2752 (N_2752,N_1777,N_1887);
nand U2753 (N_2753,N_1478,N_1728);
nor U2754 (N_2754,N_1186,N_1263);
and U2755 (N_2755,N_1227,N_1594);
nand U2756 (N_2756,N_1339,N_1883);
and U2757 (N_2757,N_1276,N_1092);
xnor U2758 (N_2758,N_1830,N_1513);
nand U2759 (N_2759,N_1887,N_1206);
or U2760 (N_2760,N_1542,N_1205);
nor U2761 (N_2761,N_1006,N_1383);
xnor U2762 (N_2762,N_1319,N_1456);
nor U2763 (N_2763,N_1617,N_1341);
or U2764 (N_2764,N_1968,N_1048);
and U2765 (N_2765,N_1042,N_1087);
nor U2766 (N_2766,N_1899,N_1690);
nand U2767 (N_2767,N_1545,N_1035);
or U2768 (N_2768,N_1371,N_1465);
nand U2769 (N_2769,N_1309,N_1245);
nand U2770 (N_2770,N_1141,N_1604);
or U2771 (N_2771,N_1693,N_1894);
and U2772 (N_2772,N_1247,N_1559);
and U2773 (N_2773,N_1038,N_1308);
nor U2774 (N_2774,N_1497,N_1593);
or U2775 (N_2775,N_1955,N_1263);
xnor U2776 (N_2776,N_1761,N_1945);
nor U2777 (N_2777,N_1016,N_1167);
or U2778 (N_2778,N_1005,N_1714);
or U2779 (N_2779,N_1466,N_1476);
nor U2780 (N_2780,N_1880,N_1724);
or U2781 (N_2781,N_1612,N_1491);
and U2782 (N_2782,N_1505,N_1838);
nor U2783 (N_2783,N_1879,N_1112);
nor U2784 (N_2784,N_1897,N_1188);
and U2785 (N_2785,N_1325,N_1926);
or U2786 (N_2786,N_1219,N_1367);
nor U2787 (N_2787,N_1439,N_1926);
nand U2788 (N_2788,N_1426,N_1845);
nand U2789 (N_2789,N_1091,N_1849);
or U2790 (N_2790,N_1574,N_1650);
xnor U2791 (N_2791,N_1077,N_1975);
nor U2792 (N_2792,N_1971,N_1615);
nand U2793 (N_2793,N_1299,N_1597);
and U2794 (N_2794,N_1999,N_1294);
xor U2795 (N_2795,N_1122,N_1807);
nand U2796 (N_2796,N_1248,N_1882);
or U2797 (N_2797,N_1086,N_1026);
nor U2798 (N_2798,N_1957,N_1725);
nand U2799 (N_2799,N_1202,N_1099);
xnor U2800 (N_2800,N_1254,N_1887);
xnor U2801 (N_2801,N_1432,N_1056);
or U2802 (N_2802,N_1630,N_1908);
nand U2803 (N_2803,N_1830,N_1035);
nor U2804 (N_2804,N_1571,N_1005);
nor U2805 (N_2805,N_1966,N_1838);
or U2806 (N_2806,N_1714,N_1498);
and U2807 (N_2807,N_1497,N_1797);
nor U2808 (N_2808,N_1386,N_1766);
nor U2809 (N_2809,N_1260,N_1928);
xnor U2810 (N_2810,N_1452,N_1635);
nand U2811 (N_2811,N_1285,N_1821);
nor U2812 (N_2812,N_1746,N_1625);
and U2813 (N_2813,N_1522,N_1349);
or U2814 (N_2814,N_1942,N_1608);
and U2815 (N_2815,N_1225,N_1835);
nand U2816 (N_2816,N_1484,N_1329);
and U2817 (N_2817,N_1633,N_1106);
xnor U2818 (N_2818,N_1302,N_1244);
nand U2819 (N_2819,N_1554,N_1129);
nand U2820 (N_2820,N_1165,N_1561);
or U2821 (N_2821,N_1265,N_1154);
or U2822 (N_2822,N_1717,N_1323);
and U2823 (N_2823,N_1201,N_1802);
nor U2824 (N_2824,N_1491,N_1560);
or U2825 (N_2825,N_1665,N_1894);
or U2826 (N_2826,N_1766,N_1281);
nor U2827 (N_2827,N_1523,N_1555);
nand U2828 (N_2828,N_1377,N_1049);
or U2829 (N_2829,N_1481,N_1577);
xor U2830 (N_2830,N_1541,N_1514);
and U2831 (N_2831,N_1511,N_1933);
xnor U2832 (N_2832,N_1991,N_1263);
nor U2833 (N_2833,N_1102,N_1616);
xor U2834 (N_2834,N_1199,N_1498);
nand U2835 (N_2835,N_1867,N_1119);
nand U2836 (N_2836,N_1633,N_1902);
or U2837 (N_2837,N_1499,N_1616);
xnor U2838 (N_2838,N_1209,N_1504);
nor U2839 (N_2839,N_1246,N_1608);
or U2840 (N_2840,N_1051,N_1258);
nor U2841 (N_2841,N_1762,N_1676);
and U2842 (N_2842,N_1990,N_1887);
and U2843 (N_2843,N_1547,N_1312);
or U2844 (N_2844,N_1574,N_1000);
or U2845 (N_2845,N_1366,N_1030);
nand U2846 (N_2846,N_1666,N_1105);
nand U2847 (N_2847,N_1833,N_1294);
and U2848 (N_2848,N_1233,N_1281);
nand U2849 (N_2849,N_1323,N_1610);
nand U2850 (N_2850,N_1760,N_1006);
xor U2851 (N_2851,N_1769,N_1186);
nand U2852 (N_2852,N_1915,N_1845);
nand U2853 (N_2853,N_1923,N_1215);
and U2854 (N_2854,N_1560,N_1793);
and U2855 (N_2855,N_1248,N_1598);
nor U2856 (N_2856,N_1068,N_1595);
nand U2857 (N_2857,N_1194,N_1046);
or U2858 (N_2858,N_1603,N_1331);
and U2859 (N_2859,N_1715,N_1544);
nor U2860 (N_2860,N_1404,N_1915);
and U2861 (N_2861,N_1128,N_1338);
xor U2862 (N_2862,N_1888,N_1572);
nand U2863 (N_2863,N_1862,N_1714);
and U2864 (N_2864,N_1233,N_1041);
nor U2865 (N_2865,N_1005,N_1236);
or U2866 (N_2866,N_1150,N_1246);
and U2867 (N_2867,N_1809,N_1267);
and U2868 (N_2868,N_1533,N_1735);
nand U2869 (N_2869,N_1437,N_1913);
nor U2870 (N_2870,N_1384,N_1039);
nor U2871 (N_2871,N_1495,N_1203);
xor U2872 (N_2872,N_1797,N_1440);
nand U2873 (N_2873,N_1026,N_1279);
or U2874 (N_2874,N_1166,N_1147);
nand U2875 (N_2875,N_1160,N_1775);
nand U2876 (N_2876,N_1886,N_1658);
nand U2877 (N_2877,N_1756,N_1498);
nor U2878 (N_2878,N_1423,N_1122);
nand U2879 (N_2879,N_1394,N_1070);
nand U2880 (N_2880,N_1100,N_1538);
xnor U2881 (N_2881,N_1092,N_1513);
nor U2882 (N_2882,N_1214,N_1322);
nand U2883 (N_2883,N_1769,N_1342);
nor U2884 (N_2884,N_1178,N_1664);
and U2885 (N_2885,N_1296,N_1127);
nand U2886 (N_2886,N_1017,N_1376);
nor U2887 (N_2887,N_1525,N_1842);
and U2888 (N_2888,N_1726,N_1821);
nor U2889 (N_2889,N_1573,N_1706);
nand U2890 (N_2890,N_1643,N_1611);
nand U2891 (N_2891,N_1746,N_1180);
nand U2892 (N_2892,N_1989,N_1343);
or U2893 (N_2893,N_1314,N_1899);
nand U2894 (N_2894,N_1533,N_1877);
or U2895 (N_2895,N_1860,N_1762);
nor U2896 (N_2896,N_1006,N_1584);
nand U2897 (N_2897,N_1469,N_1636);
and U2898 (N_2898,N_1591,N_1336);
nand U2899 (N_2899,N_1754,N_1377);
and U2900 (N_2900,N_1804,N_1873);
nand U2901 (N_2901,N_1704,N_1630);
xor U2902 (N_2902,N_1506,N_1851);
xor U2903 (N_2903,N_1569,N_1938);
or U2904 (N_2904,N_1540,N_1960);
nor U2905 (N_2905,N_1118,N_1848);
or U2906 (N_2906,N_1344,N_1304);
and U2907 (N_2907,N_1620,N_1515);
or U2908 (N_2908,N_1985,N_1314);
xnor U2909 (N_2909,N_1402,N_1837);
nand U2910 (N_2910,N_1792,N_1985);
nand U2911 (N_2911,N_1333,N_1408);
and U2912 (N_2912,N_1859,N_1009);
nand U2913 (N_2913,N_1615,N_1808);
nand U2914 (N_2914,N_1652,N_1245);
and U2915 (N_2915,N_1905,N_1964);
nand U2916 (N_2916,N_1222,N_1126);
nand U2917 (N_2917,N_1982,N_1930);
or U2918 (N_2918,N_1307,N_1867);
nor U2919 (N_2919,N_1398,N_1632);
nor U2920 (N_2920,N_1499,N_1931);
nand U2921 (N_2921,N_1214,N_1744);
or U2922 (N_2922,N_1012,N_1329);
nand U2923 (N_2923,N_1202,N_1443);
or U2924 (N_2924,N_1009,N_1348);
or U2925 (N_2925,N_1196,N_1497);
and U2926 (N_2926,N_1073,N_1410);
or U2927 (N_2927,N_1711,N_1598);
nand U2928 (N_2928,N_1405,N_1790);
and U2929 (N_2929,N_1149,N_1938);
and U2930 (N_2930,N_1554,N_1796);
nor U2931 (N_2931,N_1641,N_1598);
nor U2932 (N_2932,N_1626,N_1097);
nand U2933 (N_2933,N_1691,N_1314);
and U2934 (N_2934,N_1257,N_1923);
nor U2935 (N_2935,N_1523,N_1281);
or U2936 (N_2936,N_1965,N_1994);
nand U2937 (N_2937,N_1622,N_1031);
nand U2938 (N_2938,N_1910,N_1988);
or U2939 (N_2939,N_1867,N_1856);
nor U2940 (N_2940,N_1982,N_1911);
and U2941 (N_2941,N_1777,N_1589);
and U2942 (N_2942,N_1756,N_1017);
nand U2943 (N_2943,N_1152,N_1439);
nor U2944 (N_2944,N_1514,N_1723);
nand U2945 (N_2945,N_1966,N_1687);
nand U2946 (N_2946,N_1308,N_1935);
and U2947 (N_2947,N_1196,N_1437);
xor U2948 (N_2948,N_1854,N_1778);
xor U2949 (N_2949,N_1734,N_1748);
and U2950 (N_2950,N_1509,N_1894);
or U2951 (N_2951,N_1043,N_1328);
or U2952 (N_2952,N_1823,N_1367);
and U2953 (N_2953,N_1285,N_1476);
or U2954 (N_2954,N_1513,N_1860);
or U2955 (N_2955,N_1596,N_1221);
nand U2956 (N_2956,N_1571,N_1309);
and U2957 (N_2957,N_1978,N_1357);
or U2958 (N_2958,N_1127,N_1041);
nand U2959 (N_2959,N_1707,N_1977);
or U2960 (N_2960,N_1632,N_1928);
nor U2961 (N_2961,N_1061,N_1112);
nor U2962 (N_2962,N_1763,N_1636);
nand U2963 (N_2963,N_1936,N_1998);
or U2964 (N_2964,N_1669,N_1089);
nand U2965 (N_2965,N_1118,N_1097);
or U2966 (N_2966,N_1354,N_1833);
nor U2967 (N_2967,N_1806,N_1852);
xor U2968 (N_2968,N_1078,N_1441);
nor U2969 (N_2969,N_1925,N_1505);
or U2970 (N_2970,N_1561,N_1884);
and U2971 (N_2971,N_1031,N_1608);
xor U2972 (N_2972,N_1445,N_1475);
nand U2973 (N_2973,N_1018,N_1072);
and U2974 (N_2974,N_1359,N_1557);
and U2975 (N_2975,N_1146,N_1283);
nor U2976 (N_2976,N_1391,N_1847);
and U2977 (N_2977,N_1496,N_1037);
nand U2978 (N_2978,N_1656,N_1878);
nand U2979 (N_2979,N_1056,N_1106);
nor U2980 (N_2980,N_1131,N_1154);
or U2981 (N_2981,N_1625,N_1410);
nor U2982 (N_2982,N_1811,N_1774);
xnor U2983 (N_2983,N_1222,N_1094);
or U2984 (N_2984,N_1351,N_1149);
nor U2985 (N_2985,N_1498,N_1440);
and U2986 (N_2986,N_1029,N_1073);
nor U2987 (N_2987,N_1581,N_1628);
and U2988 (N_2988,N_1988,N_1173);
or U2989 (N_2989,N_1564,N_1696);
and U2990 (N_2990,N_1920,N_1314);
and U2991 (N_2991,N_1997,N_1901);
and U2992 (N_2992,N_1314,N_1413);
or U2993 (N_2993,N_1279,N_1018);
nand U2994 (N_2994,N_1228,N_1980);
nor U2995 (N_2995,N_1363,N_1096);
and U2996 (N_2996,N_1535,N_1270);
and U2997 (N_2997,N_1635,N_1299);
or U2998 (N_2998,N_1739,N_1668);
and U2999 (N_2999,N_1577,N_1321);
nor U3000 (N_3000,N_2581,N_2912);
and U3001 (N_3001,N_2558,N_2448);
nor U3002 (N_3002,N_2780,N_2699);
and U3003 (N_3003,N_2734,N_2915);
nand U3004 (N_3004,N_2668,N_2958);
or U3005 (N_3005,N_2034,N_2367);
nor U3006 (N_3006,N_2960,N_2049);
nor U3007 (N_3007,N_2128,N_2902);
nand U3008 (N_3008,N_2313,N_2098);
or U3009 (N_3009,N_2106,N_2062);
or U3010 (N_3010,N_2634,N_2556);
nor U3011 (N_3011,N_2302,N_2197);
or U3012 (N_3012,N_2240,N_2369);
nor U3013 (N_3013,N_2767,N_2501);
nand U3014 (N_3014,N_2251,N_2717);
nand U3015 (N_3015,N_2702,N_2771);
nand U3016 (N_3016,N_2199,N_2346);
nand U3017 (N_3017,N_2803,N_2113);
and U3018 (N_3018,N_2030,N_2656);
and U3019 (N_3019,N_2461,N_2330);
and U3020 (N_3020,N_2286,N_2715);
nand U3021 (N_3021,N_2575,N_2765);
and U3022 (N_3022,N_2292,N_2898);
nand U3023 (N_3023,N_2833,N_2573);
nand U3024 (N_3024,N_2447,N_2431);
xnor U3025 (N_3025,N_2621,N_2570);
and U3026 (N_3026,N_2123,N_2936);
or U3027 (N_3027,N_2489,N_2255);
and U3028 (N_3028,N_2498,N_2937);
or U3029 (N_3029,N_2995,N_2513);
nor U3030 (N_3030,N_2867,N_2801);
xor U3031 (N_3031,N_2409,N_2836);
nand U3032 (N_3032,N_2551,N_2081);
xnor U3033 (N_3033,N_2644,N_2817);
nor U3034 (N_3034,N_2515,N_2307);
and U3035 (N_3035,N_2185,N_2942);
xor U3036 (N_3036,N_2507,N_2872);
nand U3037 (N_3037,N_2746,N_2444);
nand U3038 (N_3038,N_2097,N_2273);
nand U3039 (N_3039,N_2257,N_2336);
nor U3040 (N_3040,N_2474,N_2052);
and U3041 (N_3041,N_2871,N_2743);
or U3042 (N_3042,N_2661,N_2149);
or U3043 (N_3043,N_2481,N_2163);
nor U3044 (N_3044,N_2617,N_2101);
xnor U3045 (N_3045,N_2844,N_2798);
or U3046 (N_3046,N_2815,N_2546);
and U3047 (N_3047,N_2945,N_2250);
nand U3048 (N_3048,N_2529,N_2204);
nor U3049 (N_3049,N_2851,N_2610);
and U3050 (N_3050,N_2266,N_2228);
xor U3051 (N_3051,N_2839,N_2229);
and U3052 (N_3052,N_2643,N_2165);
or U3053 (N_3053,N_2190,N_2506);
nand U3054 (N_3054,N_2954,N_2125);
nand U3055 (N_3055,N_2858,N_2335);
nand U3056 (N_3056,N_2516,N_2522);
nand U3057 (N_3057,N_2903,N_2027);
nor U3058 (N_3058,N_2597,N_2276);
or U3059 (N_3059,N_2278,N_2768);
and U3060 (N_3060,N_2990,N_2400);
nand U3061 (N_3061,N_2753,N_2539);
nand U3062 (N_3062,N_2907,N_2929);
or U3063 (N_3063,N_2533,N_2417);
nor U3064 (N_3064,N_2395,N_2701);
and U3065 (N_3065,N_2641,N_2994);
nor U3066 (N_3066,N_2488,N_2137);
nor U3067 (N_3067,N_2534,N_2398);
xnor U3068 (N_3068,N_2982,N_2951);
or U3069 (N_3069,N_2875,N_2855);
and U3070 (N_3070,N_2665,N_2158);
and U3071 (N_3071,N_2382,N_2747);
nor U3072 (N_3072,N_2452,N_2892);
nor U3073 (N_3073,N_2523,N_2118);
nand U3074 (N_3074,N_2209,N_2852);
nand U3075 (N_3075,N_2399,N_2735);
nor U3076 (N_3076,N_2207,N_2384);
nand U3077 (N_3077,N_2719,N_2018);
nor U3078 (N_3078,N_2394,N_2365);
or U3079 (N_3079,N_2985,N_2993);
nand U3080 (N_3080,N_2880,N_2244);
and U3081 (N_3081,N_2879,N_2467);
nor U3082 (N_3082,N_2940,N_2761);
nand U3083 (N_3083,N_2638,N_2047);
nor U3084 (N_3084,N_2624,N_2808);
nor U3085 (N_3085,N_2778,N_2944);
and U3086 (N_3086,N_2700,N_2662);
or U3087 (N_3087,N_2174,N_2325);
or U3088 (N_3088,N_2107,N_2349);
nand U3089 (N_3089,N_2970,N_2675);
and U3090 (N_3090,N_2923,N_2202);
nand U3091 (N_3091,N_2237,N_2595);
nor U3092 (N_3092,N_2950,N_2166);
xor U3093 (N_3093,N_2967,N_2732);
nor U3094 (N_3094,N_2419,N_2730);
nand U3095 (N_3095,N_2249,N_2494);
and U3096 (N_3096,N_2949,N_2913);
and U3097 (N_3097,N_2345,N_2390);
nor U3098 (N_3098,N_2195,N_2025);
or U3099 (N_3099,N_2979,N_2070);
nand U3100 (N_3100,N_2305,N_2866);
nor U3101 (N_3101,N_2385,N_2846);
or U3102 (N_3102,N_2530,N_2019);
or U3103 (N_3103,N_2807,N_2147);
nand U3104 (N_3104,N_2964,N_2233);
nand U3105 (N_3105,N_2178,N_2164);
and U3106 (N_3106,N_2391,N_2776);
or U3107 (N_3107,N_2961,N_2598);
nand U3108 (N_3108,N_2777,N_2426);
nand U3109 (N_3109,N_2075,N_2989);
xor U3110 (N_3110,N_2405,N_2469);
and U3111 (N_3111,N_2526,N_2442);
or U3112 (N_3112,N_2517,N_2230);
nor U3113 (N_3113,N_2594,N_2572);
nand U3114 (N_3114,N_2463,N_2591);
and U3115 (N_3115,N_2122,N_2381);
or U3116 (N_3116,N_2117,N_2001);
nand U3117 (N_3117,N_2800,N_2583);
xnor U3118 (N_3118,N_2876,N_2681);
or U3119 (N_3119,N_2383,N_2059);
and U3120 (N_3120,N_2087,N_2766);
nor U3121 (N_3121,N_2115,N_2468);
nor U3122 (N_3122,N_2562,N_2235);
nand U3123 (N_3123,N_2068,N_2022);
nand U3124 (N_3124,N_2193,N_2248);
nand U3125 (N_3125,N_2180,N_2810);
nor U3126 (N_3126,N_2672,N_2525);
and U3127 (N_3127,N_2181,N_2794);
or U3128 (N_3128,N_2042,N_2457);
nand U3129 (N_3129,N_2553,N_2883);
xor U3130 (N_3130,N_2368,N_2015);
nor U3131 (N_3131,N_2718,N_2366);
nand U3132 (N_3132,N_2884,N_2514);
and U3133 (N_3133,N_2601,N_2757);
and U3134 (N_3134,N_2509,N_2911);
nand U3135 (N_3135,N_2031,N_2016);
nand U3136 (N_3136,N_2231,N_2756);
or U3137 (N_3137,N_2592,N_2375);
or U3138 (N_3138,N_2535,N_2840);
or U3139 (N_3139,N_2003,N_2243);
or U3140 (N_3140,N_2804,N_2978);
and U3141 (N_3141,N_2722,N_2543);
nand U3142 (N_3142,N_2714,N_2626);
nor U3143 (N_3143,N_2955,N_2011);
nor U3144 (N_3144,N_2565,N_2704);
nand U3145 (N_3145,N_2261,N_2969);
or U3146 (N_3146,N_2222,N_2479);
xnor U3147 (N_3147,N_2088,N_2758);
or U3148 (N_3148,N_2491,N_2008);
and U3149 (N_3149,N_2932,N_2301);
nor U3150 (N_3150,N_2999,N_2609);
and U3151 (N_3151,N_2168,N_2897);
or U3152 (N_3152,N_2121,N_2139);
nand U3153 (N_3153,N_2607,N_2845);
nand U3154 (N_3154,N_2264,N_2211);
or U3155 (N_3155,N_2772,N_2373);
nor U3156 (N_3156,N_2434,N_2737);
nand U3157 (N_3157,N_2439,N_2537);
nand U3158 (N_3158,N_2731,N_2420);
nor U3159 (N_3159,N_2371,N_2557);
and U3160 (N_3160,N_2239,N_2425);
or U3161 (N_3161,N_2020,N_2520);
nand U3162 (N_3162,N_2318,N_2895);
nand U3163 (N_3163,N_2299,N_2397);
or U3164 (N_3164,N_2411,N_2484);
nor U3165 (N_3165,N_2716,N_2099);
xor U3166 (N_3166,N_2900,N_2012);
or U3167 (N_3167,N_2374,N_2406);
or U3168 (N_3168,N_2423,N_2647);
or U3169 (N_3169,N_2933,N_2724);
or U3170 (N_3170,N_2182,N_2187);
and U3171 (N_3171,N_2928,N_2194);
or U3172 (N_3172,N_2709,N_2496);
or U3173 (N_3173,N_2613,N_2502);
and U3174 (N_3174,N_2486,N_2683);
and U3175 (N_3175,N_2536,N_2192);
nand U3176 (N_3176,N_2612,N_2429);
or U3177 (N_3177,N_2450,N_2674);
and U3178 (N_3178,N_2952,N_2487);
nor U3179 (N_3179,N_2069,N_2823);
nor U3180 (N_3180,N_2646,N_2627);
and U3181 (N_3181,N_2449,N_2162);
nand U3182 (N_3182,N_2339,N_2310);
nand U3183 (N_3183,N_2331,N_2749);
nand U3184 (N_3184,N_2210,N_2454);
nor U3185 (N_3185,N_2303,N_2850);
nand U3186 (N_3186,N_2669,N_2762);
nor U3187 (N_3187,N_2973,N_2322);
and U3188 (N_3188,N_2268,N_2976);
nor U3189 (N_3189,N_2280,N_2129);
or U3190 (N_3190,N_2215,N_2790);
and U3191 (N_3191,N_2329,N_2917);
nor U3192 (N_3192,N_2023,N_2205);
nor U3193 (N_3193,N_2721,N_2309);
nor U3194 (N_3194,N_2853,N_2102);
nand U3195 (N_3195,N_2010,N_2750);
or U3196 (N_3196,N_2291,N_2363);
xor U3197 (N_3197,N_2584,N_2116);
and U3198 (N_3198,N_2380,N_2065);
or U3199 (N_3199,N_2671,N_2651);
nor U3200 (N_3200,N_2652,N_2208);
nor U3201 (N_3201,N_2130,N_2588);
and U3202 (N_3202,N_2044,N_2014);
and U3203 (N_3203,N_2890,N_2868);
xnor U3204 (N_3204,N_2682,N_2054);
and U3205 (N_3205,N_2242,N_2860);
or U3206 (N_3206,N_2095,N_2337);
nor U3207 (N_3207,N_2080,N_2298);
nor U3208 (N_3208,N_2818,N_2300);
or U3209 (N_3209,N_2143,N_2376);
nor U3210 (N_3210,N_2378,N_2133);
or U3211 (N_3211,N_2691,N_2623);
nand U3212 (N_3212,N_2596,N_2629);
xor U3213 (N_3213,N_2848,N_2692);
or U3214 (N_3214,N_2874,N_2896);
or U3215 (N_3215,N_2495,N_2763);
and U3216 (N_3216,N_2492,N_2813);
and U3217 (N_3217,N_2548,N_2028);
or U3218 (N_3218,N_2500,N_2538);
nand U3219 (N_3219,N_2091,N_2304);
or U3220 (N_3220,N_2580,N_2996);
nand U3221 (N_3221,N_2408,N_2684);
and U3222 (N_3222,N_2972,N_2909);
nor U3223 (N_3223,N_2407,N_2574);
nand U3224 (N_3224,N_2549,N_2635);
nand U3225 (N_3225,N_2865,N_2480);
nor U3226 (N_3226,N_2687,N_2939);
nand U3227 (N_3227,N_2512,N_2555);
nor U3228 (N_3228,N_2105,N_2029);
xor U3229 (N_3229,N_2916,N_2055);
or U3230 (N_3230,N_2071,N_2477);
and U3231 (N_3231,N_2728,N_2333);
xor U3232 (N_3232,N_2100,N_2037);
nor U3233 (N_3233,N_2048,N_2482);
or U3234 (N_3234,N_2812,N_2402);
and U3235 (N_3235,N_2720,N_2177);
xor U3236 (N_3236,N_2152,N_2111);
nor U3237 (N_3237,N_2751,N_2931);
nor U3238 (N_3238,N_2649,N_2830);
nand U3239 (N_3239,N_2882,N_2567);
nor U3240 (N_3240,N_2770,N_2791);
nor U3241 (N_3241,N_2578,N_2259);
nor U3242 (N_3242,N_2981,N_2676);
nand U3243 (N_3243,N_2155,N_2446);
nor U3244 (N_3244,N_2938,N_2806);
or U3245 (N_3245,N_2103,N_2350);
and U3246 (N_3246,N_2991,N_2109);
and U3247 (N_3247,N_2424,N_2899);
and U3248 (N_3248,N_2358,N_2258);
xor U3249 (N_3249,N_2053,N_2473);
and U3250 (N_3250,N_2711,N_2466);
or U3251 (N_3251,N_2279,N_2490);
and U3252 (N_3252,N_2593,N_2579);
or U3253 (N_3253,N_2033,N_2849);
and U3254 (N_3254,N_2505,N_2114);
and U3255 (N_3255,N_2201,N_2364);
and U3256 (N_3256,N_2393,N_2415);
nor U3257 (N_3257,N_2078,N_2226);
and U3258 (N_3258,N_2157,N_2926);
or U3259 (N_3259,N_2148,N_2645);
nand U3260 (N_3260,N_2223,N_2614);
nor U3261 (N_3261,N_2703,N_2108);
or U3262 (N_3262,N_2540,N_2901);
and U3263 (N_3263,N_2733,N_2348);
nand U3264 (N_3264,N_2904,N_2126);
nor U3265 (N_3265,N_2156,N_2306);
nor U3266 (N_3266,N_2908,N_2485);
and U3267 (N_3267,N_2021,N_2561);
xor U3268 (N_3268,N_2503,N_2564);
and U3269 (N_3269,N_2922,N_2738);
nand U3270 (N_3270,N_2631,N_2093);
nand U3271 (N_3271,N_2524,N_2270);
nor U3272 (N_3272,N_2064,N_2657);
nor U3273 (N_3273,N_2172,N_2056);
and U3274 (N_3274,N_2045,N_2041);
nand U3275 (N_3275,N_2074,N_2294);
and U3276 (N_3276,N_2079,N_2063);
or U3277 (N_3277,N_2317,N_2616);
nand U3278 (N_3278,N_2712,N_2443);
or U3279 (N_3279,N_2925,N_2959);
and U3280 (N_3280,N_2814,N_2372);
and U3281 (N_3281,N_2472,N_2677);
and U3282 (N_3282,N_2698,N_2060);
or U3283 (N_3283,N_2618,N_2404);
and U3284 (N_3284,N_2504,N_2269);
or U3285 (N_3285,N_2795,N_2356);
or U3286 (N_3286,N_2965,N_2630);
nor U3287 (N_3287,N_2764,N_2387);
nor U3288 (N_3288,N_2986,N_2962);
or U3289 (N_3289,N_2013,N_2067);
nand U3290 (N_3290,N_2234,N_2038);
nor U3291 (N_3291,N_2664,N_2566);
and U3292 (N_3292,N_2953,N_2963);
and U3293 (N_3293,N_2835,N_2024);
or U3294 (N_3294,N_2092,N_2948);
and U3295 (N_3295,N_2686,N_2151);
nor U3296 (N_3296,N_2706,N_2328);
or U3297 (N_3297,N_2773,N_2998);
nor U3298 (N_3298,N_2769,N_2396);
nor U3299 (N_3299,N_2218,N_2587);
or U3300 (N_3300,N_2464,N_2401);
nor U3301 (N_3301,N_2083,N_2983);
nand U3302 (N_3302,N_2822,N_2666);
and U3303 (N_3303,N_2797,N_2220);
and U3304 (N_3304,N_2825,N_2873);
or U3305 (N_3305,N_2497,N_2935);
nand U3306 (N_3306,N_2085,N_2914);
nor U3307 (N_3307,N_2726,N_2341);
nor U3308 (N_3308,N_2082,N_2253);
nand U3309 (N_3309,N_2971,N_2988);
nor U3310 (N_3310,N_2673,N_2351);
nor U3311 (N_3311,N_2475,N_2975);
nand U3312 (N_3312,N_2412,N_2314);
or U3313 (N_3313,N_2427,N_2799);
and U3314 (N_3314,N_2238,N_2416);
and U3315 (N_3315,N_2046,N_2422);
and U3316 (N_3316,N_2527,N_2453);
or U3317 (N_3317,N_2589,N_2094);
xnor U3318 (N_3318,N_2744,N_2343);
or U3319 (N_3319,N_2216,N_2430);
xnor U3320 (N_3320,N_2334,N_2550);
nor U3321 (N_3321,N_2816,N_2077);
nand U3322 (N_3322,N_2569,N_2110);
nand U3323 (N_3323,N_2340,N_2256);
nor U3324 (N_3324,N_2323,N_2219);
nand U3325 (N_3325,N_2277,N_2586);
nor U3326 (N_3326,N_2531,N_2619);
xor U3327 (N_3327,N_2811,N_2282);
or U3328 (N_3328,N_2377,N_2140);
xnor U3329 (N_3329,N_2347,N_2252);
or U3330 (N_3330,N_2135,N_2161);
nand U3331 (N_3331,N_2186,N_2984);
or U3332 (N_3332,N_2386,N_2842);
nand U3333 (N_3333,N_2805,N_2320);
or U3334 (N_3334,N_2642,N_2315);
or U3335 (N_3335,N_2154,N_2774);
nand U3336 (N_3336,N_2779,N_2740);
or U3337 (N_3337,N_2311,N_2392);
and U3338 (N_3338,N_2221,N_2000);
nor U3339 (N_3339,N_2946,N_2032);
xnor U3340 (N_3340,N_2957,N_2036);
nand U3341 (N_3341,N_2820,N_2232);
and U3342 (N_3342,N_2285,N_2039);
or U3343 (N_3343,N_2889,N_2650);
and U3344 (N_3344,N_2150,N_2659);
nor U3345 (N_3345,N_2653,N_2212);
xnor U3346 (N_3346,N_2752,N_2679);
and U3347 (N_3347,N_2002,N_2321);
and U3348 (N_3348,N_2196,N_2217);
nand U3349 (N_3349,N_2793,N_2974);
nor U3350 (N_3350,N_2528,N_2729);
and U3351 (N_3351,N_2437,N_2227);
and U3352 (N_3352,N_2863,N_2354);
and U3353 (N_3353,N_2061,N_2224);
xor U3354 (N_3354,N_2727,N_2361);
xor U3355 (N_3355,N_2802,N_2782);
or U3356 (N_3356,N_2355,N_2748);
or U3357 (N_3357,N_2678,N_2456);
or U3358 (N_3358,N_2854,N_2870);
xor U3359 (N_3359,N_2357,N_2824);
nand U3360 (N_3360,N_2127,N_2784);
and U3361 (N_3361,N_2312,N_2544);
and U3362 (N_3362,N_2585,N_2606);
or U3363 (N_3363,N_2342,N_2086);
or U3364 (N_3364,N_2834,N_2200);
nor U3365 (N_3365,N_2176,N_2435);
or U3366 (N_3366,N_2987,N_2009);
xor U3367 (N_3367,N_2066,N_2171);
nor U3368 (N_3368,N_2035,N_2519);
nand U3369 (N_3369,N_2745,N_2919);
nand U3370 (N_3370,N_2465,N_2017);
nor U3371 (N_3371,N_2175,N_2636);
nand U3372 (N_3372,N_2640,N_2690);
or U3373 (N_3373,N_2451,N_2831);
nor U3374 (N_3374,N_2796,N_2203);
and U3375 (N_3375,N_2620,N_2877);
nor U3376 (N_3376,N_2254,N_2179);
nor U3377 (N_3377,N_2421,N_2295);
nor U3378 (N_3378,N_2605,N_2787);
or U3379 (N_3379,N_2247,N_2198);
nor U3380 (N_3380,N_2563,N_2124);
nor U3381 (N_3381,N_2775,N_2138);
and U3382 (N_3382,N_2142,N_2288);
xnor U3383 (N_3383,N_2847,N_2146);
and U3384 (N_3384,N_2697,N_2460);
nand U3385 (N_3385,N_2582,N_2881);
and U3386 (N_3386,N_2602,N_2338);
nor U3387 (N_3387,N_2696,N_2947);
or U3388 (N_3388,N_2878,N_2708);
nand U3389 (N_3389,N_2966,N_2600);
and U3390 (N_3390,N_2861,N_2783);
nor U3391 (N_3391,N_2693,N_2603);
nor U3392 (N_3392,N_2441,N_2508);
or U3393 (N_3393,N_2471,N_2167);
nand U3394 (N_3394,N_2459,N_2262);
or U3395 (N_3395,N_2326,N_2590);
nor U3396 (N_3396,N_2189,N_2921);
xnor U3397 (N_3397,N_2622,N_2759);
and U3398 (N_3398,N_2159,N_2319);
or U3399 (N_3399,N_2272,N_2275);
and U3400 (N_3400,N_2433,N_2785);
nor U3401 (N_3401,N_2841,N_2639);
nand U3402 (N_3402,N_2827,N_2414);
xnor U3403 (N_3403,N_2284,N_2308);
xor U3404 (N_3404,N_2265,N_2418);
nand U3405 (N_3405,N_2120,N_2051);
nand U3406 (N_3406,N_2511,N_2478);
or U3407 (N_3407,N_2930,N_2436);
xnor U3408 (N_3408,N_2483,N_2560);
or U3409 (N_3409,N_2510,N_2723);
or U3410 (N_3410,N_2821,N_2005);
and U3411 (N_3411,N_2760,N_2058);
nor U3412 (N_3412,N_2689,N_2173);
nor U3413 (N_3413,N_2568,N_2943);
and U3414 (N_3414,N_2287,N_2741);
and U3415 (N_3415,N_2910,N_2297);
or U3416 (N_3416,N_2455,N_2260);
or U3417 (N_3417,N_2043,N_2541);
nor U3418 (N_3418,N_2552,N_2476);
and U3419 (N_3419,N_2633,N_2316);
nor U3420 (N_3420,N_2905,N_2694);
or U3421 (N_3421,N_2445,N_2353);
nand U3422 (N_3422,N_2428,N_2007);
nor U3423 (N_3423,N_2352,N_2296);
and U3424 (N_3424,N_2611,N_2742);
xnor U3425 (N_3425,N_2183,N_2112);
and U3426 (N_3426,N_2332,N_2924);
or U3427 (N_3427,N_2707,N_2559);
nand U3428 (N_3428,N_2263,N_2856);
or U3429 (N_3429,N_2888,N_2660);
xnor U3430 (N_3430,N_2119,N_2688);
nand U3431 (N_3431,N_2236,N_2680);
nor U3432 (N_3432,N_2134,N_2104);
and U3433 (N_3433,N_2887,N_2245);
or U3434 (N_3434,N_2050,N_2755);
nand U3435 (N_3435,N_2281,N_2927);
nand U3436 (N_3436,N_2184,N_2084);
nor U3437 (N_3437,N_2632,N_2090);
nand U3438 (N_3438,N_2293,N_2739);
and U3439 (N_3439,N_2379,N_2843);
nand U3440 (N_3440,N_2359,N_2781);
nand U3441 (N_3441,N_2710,N_2289);
xor U3442 (N_3442,N_2153,N_2792);
xnor U3443 (N_3443,N_2956,N_2545);
xor U3444 (N_3444,N_2625,N_2499);
nand U3445 (N_3445,N_2169,N_2615);
nand U3446 (N_3446,N_2470,N_2885);
nor U3447 (N_3447,N_2413,N_2283);
and U3448 (N_3448,N_2918,N_2004);
nor U3449 (N_3449,N_2191,N_2225);
nand U3450 (N_3450,N_2089,N_2992);
nand U3451 (N_3451,N_2862,N_2997);
xnor U3452 (N_3452,N_2073,N_2206);
and U3453 (N_3453,N_2705,N_2829);
and U3454 (N_3454,N_2389,N_2655);
nor U3455 (N_3455,N_2886,N_2542);
or U3456 (N_3456,N_2026,N_2663);
and U3457 (N_3457,N_2754,N_2170);
nor U3458 (N_3458,N_2713,N_2554);
and U3459 (N_3459,N_2132,N_2214);
nor U3460 (N_3460,N_2685,N_2920);
nand U3461 (N_3461,N_2906,N_2869);
and U3462 (N_3462,N_2144,N_2628);
nand U3463 (N_3463,N_2271,N_2637);
nor U3464 (N_3464,N_2968,N_2327);
and U3465 (N_3465,N_2324,N_2891);
and U3466 (N_3466,N_2136,N_2388);
xnor U3467 (N_3467,N_2608,N_2599);
or U3468 (N_3468,N_2438,N_2577);
and U3469 (N_3469,N_2072,N_2658);
and U3470 (N_3470,N_2362,N_2076);
and U3471 (N_3471,N_2246,N_2789);
nor U3472 (N_3472,N_2518,N_2547);
and U3473 (N_3473,N_2370,N_2893);
nor U3474 (N_3474,N_2828,N_2440);
nor U3475 (N_3475,N_2141,N_2654);
xor U3476 (N_3476,N_2096,N_2667);
and U3477 (N_3477,N_2213,N_2725);
nor U3478 (N_3478,N_2838,N_2403);
nand U3479 (N_3479,N_2571,N_2040);
nor U3480 (N_3480,N_2410,N_2462);
nor U3481 (N_3481,N_2521,N_2648);
and U3482 (N_3482,N_2934,N_2532);
or U3483 (N_3483,N_2006,N_2131);
or U3484 (N_3484,N_2941,N_2057);
and U3485 (N_3485,N_2576,N_2360);
nand U3486 (N_3486,N_2695,N_2857);
or U3487 (N_3487,N_2980,N_2826);
or U3488 (N_3488,N_2432,N_2837);
or U3489 (N_3489,N_2160,N_2894);
nand U3490 (N_3490,N_2832,N_2788);
or U3491 (N_3491,N_2977,N_2864);
and U3492 (N_3492,N_2493,N_2290);
nor U3493 (N_3493,N_2145,N_2458);
and U3494 (N_3494,N_2786,N_2274);
and U3495 (N_3495,N_2670,N_2267);
nor U3496 (N_3496,N_2604,N_2809);
and U3497 (N_3497,N_2344,N_2241);
nand U3498 (N_3498,N_2819,N_2859);
nor U3499 (N_3499,N_2736,N_2188);
nor U3500 (N_3500,N_2970,N_2792);
nor U3501 (N_3501,N_2207,N_2935);
nor U3502 (N_3502,N_2568,N_2698);
nor U3503 (N_3503,N_2965,N_2981);
and U3504 (N_3504,N_2438,N_2581);
nor U3505 (N_3505,N_2650,N_2699);
and U3506 (N_3506,N_2850,N_2731);
or U3507 (N_3507,N_2237,N_2317);
nor U3508 (N_3508,N_2253,N_2283);
nor U3509 (N_3509,N_2030,N_2760);
and U3510 (N_3510,N_2277,N_2235);
xor U3511 (N_3511,N_2283,N_2337);
xor U3512 (N_3512,N_2215,N_2343);
nand U3513 (N_3513,N_2380,N_2443);
nand U3514 (N_3514,N_2958,N_2667);
or U3515 (N_3515,N_2864,N_2528);
nor U3516 (N_3516,N_2074,N_2758);
nand U3517 (N_3517,N_2955,N_2924);
or U3518 (N_3518,N_2440,N_2702);
and U3519 (N_3519,N_2196,N_2892);
nor U3520 (N_3520,N_2555,N_2467);
nor U3521 (N_3521,N_2893,N_2398);
or U3522 (N_3522,N_2494,N_2336);
or U3523 (N_3523,N_2207,N_2799);
nor U3524 (N_3524,N_2198,N_2167);
nor U3525 (N_3525,N_2733,N_2016);
nor U3526 (N_3526,N_2618,N_2446);
nor U3527 (N_3527,N_2919,N_2644);
or U3528 (N_3528,N_2909,N_2727);
nor U3529 (N_3529,N_2761,N_2695);
and U3530 (N_3530,N_2916,N_2419);
or U3531 (N_3531,N_2122,N_2697);
nand U3532 (N_3532,N_2483,N_2556);
and U3533 (N_3533,N_2176,N_2654);
nand U3534 (N_3534,N_2757,N_2699);
xor U3535 (N_3535,N_2524,N_2138);
nor U3536 (N_3536,N_2409,N_2669);
and U3537 (N_3537,N_2245,N_2877);
and U3538 (N_3538,N_2601,N_2526);
nor U3539 (N_3539,N_2210,N_2417);
nand U3540 (N_3540,N_2776,N_2028);
nand U3541 (N_3541,N_2704,N_2939);
nor U3542 (N_3542,N_2790,N_2185);
or U3543 (N_3543,N_2999,N_2135);
nor U3544 (N_3544,N_2813,N_2339);
nand U3545 (N_3545,N_2312,N_2185);
nor U3546 (N_3546,N_2442,N_2837);
and U3547 (N_3547,N_2183,N_2959);
nor U3548 (N_3548,N_2779,N_2385);
nor U3549 (N_3549,N_2526,N_2763);
nor U3550 (N_3550,N_2238,N_2146);
or U3551 (N_3551,N_2629,N_2221);
or U3552 (N_3552,N_2662,N_2122);
nand U3553 (N_3553,N_2400,N_2154);
nor U3554 (N_3554,N_2279,N_2633);
nand U3555 (N_3555,N_2223,N_2791);
nand U3556 (N_3556,N_2248,N_2232);
and U3557 (N_3557,N_2276,N_2539);
and U3558 (N_3558,N_2468,N_2328);
or U3559 (N_3559,N_2543,N_2878);
and U3560 (N_3560,N_2395,N_2511);
xnor U3561 (N_3561,N_2687,N_2478);
nor U3562 (N_3562,N_2896,N_2872);
nand U3563 (N_3563,N_2592,N_2632);
or U3564 (N_3564,N_2881,N_2549);
or U3565 (N_3565,N_2075,N_2055);
and U3566 (N_3566,N_2788,N_2130);
nand U3567 (N_3567,N_2171,N_2476);
xor U3568 (N_3568,N_2661,N_2792);
nor U3569 (N_3569,N_2460,N_2114);
and U3570 (N_3570,N_2330,N_2719);
nor U3571 (N_3571,N_2056,N_2197);
xor U3572 (N_3572,N_2704,N_2397);
nand U3573 (N_3573,N_2584,N_2071);
xor U3574 (N_3574,N_2030,N_2970);
and U3575 (N_3575,N_2202,N_2397);
nand U3576 (N_3576,N_2020,N_2264);
nand U3577 (N_3577,N_2674,N_2138);
or U3578 (N_3578,N_2747,N_2472);
and U3579 (N_3579,N_2196,N_2675);
nand U3580 (N_3580,N_2677,N_2517);
and U3581 (N_3581,N_2985,N_2908);
and U3582 (N_3582,N_2278,N_2314);
and U3583 (N_3583,N_2428,N_2144);
or U3584 (N_3584,N_2420,N_2121);
xor U3585 (N_3585,N_2911,N_2653);
or U3586 (N_3586,N_2719,N_2406);
nor U3587 (N_3587,N_2378,N_2846);
nand U3588 (N_3588,N_2615,N_2382);
nor U3589 (N_3589,N_2994,N_2687);
nand U3590 (N_3590,N_2565,N_2343);
xor U3591 (N_3591,N_2592,N_2535);
nor U3592 (N_3592,N_2333,N_2984);
and U3593 (N_3593,N_2375,N_2800);
or U3594 (N_3594,N_2692,N_2974);
nor U3595 (N_3595,N_2006,N_2166);
or U3596 (N_3596,N_2733,N_2410);
or U3597 (N_3597,N_2653,N_2108);
and U3598 (N_3598,N_2459,N_2137);
nand U3599 (N_3599,N_2098,N_2993);
nand U3600 (N_3600,N_2165,N_2176);
nor U3601 (N_3601,N_2209,N_2518);
xor U3602 (N_3602,N_2047,N_2883);
or U3603 (N_3603,N_2283,N_2939);
or U3604 (N_3604,N_2464,N_2274);
or U3605 (N_3605,N_2966,N_2439);
xor U3606 (N_3606,N_2280,N_2961);
or U3607 (N_3607,N_2723,N_2809);
or U3608 (N_3608,N_2731,N_2715);
or U3609 (N_3609,N_2175,N_2155);
or U3610 (N_3610,N_2025,N_2524);
xnor U3611 (N_3611,N_2346,N_2569);
or U3612 (N_3612,N_2058,N_2977);
nor U3613 (N_3613,N_2677,N_2645);
or U3614 (N_3614,N_2772,N_2928);
or U3615 (N_3615,N_2389,N_2091);
nor U3616 (N_3616,N_2543,N_2749);
or U3617 (N_3617,N_2075,N_2117);
and U3618 (N_3618,N_2310,N_2755);
nand U3619 (N_3619,N_2804,N_2458);
and U3620 (N_3620,N_2982,N_2679);
nand U3621 (N_3621,N_2132,N_2307);
or U3622 (N_3622,N_2446,N_2370);
and U3623 (N_3623,N_2340,N_2242);
nor U3624 (N_3624,N_2148,N_2485);
nand U3625 (N_3625,N_2771,N_2391);
or U3626 (N_3626,N_2105,N_2811);
nand U3627 (N_3627,N_2231,N_2687);
and U3628 (N_3628,N_2195,N_2866);
or U3629 (N_3629,N_2255,N_2250);
and U3630 (N_3630,N_2777,N_2928);
nand U3631 (N_3631,N_2688,N_2359);
nand U3632 (N_3632,N_2259,N_2251);
and U3633 (N_3633,N_2165,N_2531);
xnor U3634 (N_3634,N_2838,N_2641);
nand U3635 (N_3635,N_2581,N_2888);
nand U3636 (N_3636,N_2818,N_2991);
nor U3637 (N_3637,N_2731,N_2431);
nor U3638 (N_3638,N_2445,N_2462);
nor U3639 (N_3639,N_2828,N_2499);
or U3640 (N_3640,N_2667,N_2133);
nor U3641 (N_3641,N_2314,N_2629);
nor U3642 (N_3642,N_2955,N_2850);
xor U3643 (N_3643,N_2763,N_2999);
or U3644 (N_3644,N_2148,N_2625);
nor U3645 (N_3645,N_2352,N_2854);
nor U3646 (N_3646,N_2658,N_2950);
and U3647 (N_3647,N_2475,N_2085);
xnor U3648 (N_3648,N_2282,N_2464);
or U3649 (N_3649,N_2946,N_2085);
or U3650 (N_3650,N_2598,N_2324);
xnor U3651 (N_3651,N_2474,N_2745);
xor U3652 (N_3652,N_2692,N_2163);
nand U3653 (N_3653,N_2542,N_2366);
and U3654 (N_3654,N_2179,N_2800);
or U3655 (N_3655,N_2885,N_2692);
and U3656 (N_3656,N_2494,N_2984);
and U3657 (N_3657,N_2119,N_2137);
or U3658 (N_3658,N_2528,N_2661);
and U3659 (N_3659,N_2084,N_2611);
and U3660 (N_3660,N_2084,N_2575);
nand U3661 (N_3661,N_2628,N_2288);
nor U3662 (N_3662,N_2266,N_2570);
and U3663 (N_3663,N_2010,N_2853);
nor U3664 (N_3664,N_2022,N_2710);
or U3665 (N_3665,N_2556,N_2924);
or U3666 (N_3666,N_2225,N_2483);
or U3667 (N_3667,N_2800,N_2103);
nand U3668 (N_3668,N_2100,N_2278);
and U3669 (N_3669,N_2575,N_2944);
nand U3670 (N_3670,N_2262,N_2853);
or U3671 (N_3671,N_2223,N_2901);
nor U3672 (N_3672,N_2911,N_2635);
or U3673 (N_3673,N_2760,N_2782);
nand U3674 (N_3674,N_2101,N_2208);
or U3675 (N_3675,N_2674,N_2430);
xor U3676 (N_3676,N_2553,N_2230);
or U3677 (N_3677,N_2088,N_2867);
nor U3678 (N_3678,N_2088,N_2045);
or U3679 (N_3679,N_2093,N_2661);
nand U3680 (N_3680,N_2618,N_2044);
or U3681 (N_3681,N_2366,N_2374);
nand U3682 (N_3682,N_2621,N_2139);
and U3683 (N_3683,N_2632,N_2230);
or U3684 (N_3684,N_2429,N_2338);
nand U3685 (N_3685,N_2526,N_2162);
and U3686 (N_3686,N_2129,N_2138);
or U3687 (N_3687,N_2465,N_2418);
and U3688 (N_3688,N_2171,N_2228);
nand U3689 (N_3689,N_2760,N_2678);
or U3690 (N_3690,N_2420,N_2385);
nand U3691 (N_3691,N_2274,N_2056);
or U3692 (N_3692,N_2829,N_2174);
nand U3693 (N_3693,N_2013,N_2708);
xnor U3694 (N_3694,N_2684,N_2171);
and U3695 (N_3695,N_2886,N_2396);
nand U3696 (N_3696,N_2741,N_2217);
nor U3697 (N_3697,N_2444,N_2048);
nor U3698 (N_3698,N_2002,N_2149);
or U3699 (N_3699,N_2328,N_2276);
nand U3700 (N_3700,N_2800,N_2865);
nor U3701 (N_3701,N_2040,N_2529);
nand U3702 (N_3702,N_2847,N_2912);
or U3703 (N_3703,N_2418,N_2711);
or U3704 (N_3704,N_2281,N_2630);
or U3705 (N_3705,N_2432,N_2612);
nor U3706 (N_3706,N_2599,N_2414);
or U3707 (N_3707,N_2770,N_2190);
or U3708 (N_3708,N_2607,N_2203);
nand U3709 (N_3709,N_2619,N_2140);
nand U3710 (N_3710,N_2011,N_2636);
nand U3711 (N_3711,N_2623,N_2150);
or U3712 (N_3712,N_2885,N_2900);
and U3713 (N_3713,N_2977,N_2910);
and U3714 (N_3714,N_2671,N_2889);
nor U3715 (N_3715,N_2905,N_2663);
or U3716 (N_3716,N_2161,N_2327);
and U3717 (N_3717,N_2029,N_2423);
or U3718 (N_3718,N_2667,N_2468);
nand U3719 (N_3719,N_2462,N_2708);
xor U3720 (N_3720,N_2279,N_2710);
or U3721 (N_3721,N_2672,N_2024);
or U3722 (N_3722,N_2586,N_2013);
nor U3723 (N_3723,N_2175,N_2711);
nor U3724 (N_3724,N_2239,N_2206);
and U3725 (N_3725,N_2563,N_2394);
nand U3726 (N_3726,N_2786,N_2154);
or U3727 (N_3727,N_2770,N_2118);
or U3728 (N_3728,N_2941,N_2878);
and U3729 (N_3729,N_2205,N_2755);
nor U3730 (N_3730,N_2882,N_2117);
nor U3731 (N_3731,N_2865,N_2292);
nand U3732 (N_3732,N_2414,N_2065);
or U3733 (N_3733,N_2705,N_2421);
xnor U3734 (N_3734,N_2493,N_2861);
nand U3735 (N_3735,N_2799,N_2505);
and U3736 (N_3736,N_2511,N_2023);
and U3737 (N_3737,N_2322,N_2336);
and U3738 (N_3738,N_2686,N_2330);
or U3739 (N_3739,N_2383,N_2361);
and U3740 (N_3740,N_2771,N_2108);
and U3741 (N_3741,N_2262,N_2483);
nand U3742 (N_3742,N_2647,N_2378);
nand U3743 (N_3743,N_2632,N_2847);
nand U3744 (N_3744,N_2122,N_2650);
and U3745 (N_3745,N_2575,N_2702);
and U3746 (N_3746,N_2238,N_2873);
xnor U3747 (N_3747,N_2555,N_2960);
and U3748 (N_3748,N_2629,N_2142);
xor U3749 (N_3749,N_2280,N_2078);
and U3750 (N_3750,N_2057,N_2007);
nor U3751 (N_3751,N_2911,N_2599);
nor U3752 (N_3752,N_2412,N_2636);
nor U3753 (N_3753,N_2342,N_2559);
or U3754 (N_3754,N_2507,N_2698);
nor U3755 (N_3755,N_2669,N_2310);
nor U3756 (N_3756,N_2509,N_2615);
xnor U3757 (N_3757,N_2529,N_2950);
or U3758 (N_3758,N_2439,N_2360);
nand U3759 (N_3759,N_2872,N_2806);
and U3760 (N_3760,N_2951,N_2150);
or U3761 (N_3761,N_2726,N_2697);
xnor U3762 (N_3762,N_2295,N_2676);
xor U3763 (N_3763,N_2839,N_2070);
nand U3764 (N_3764,N_2026,N_2811);
and U3765 (N_3765,N_2015,N_2688);
nand U3766 (N_3766,N_2940,N_2120);
and U3767 (N_3767,N_2079,N_2262);
nor U3768 (N_3768,N_2113,N_2777);
and U3769 (N_3769,N_2621,N_2536);
nand U3770 (N_3770,N_2572,N_2411);
xor U3771 (N_3771,N_2082,N_2351);
or U3772 (N_3772,N_2185,N_2781);
xnor U3773 (N_3773,N_2754,N_2432);
and U3774 (N_3774,N_2881,N_2761);
nor U3775 (N_3775,N_2973,N_2535);
nor U3776 (N_3776,N_2616,N_2331);
nor U3777 (N_3777,N_2436,N_2363);
and U3778 (N_3778,N_2790,N_2130);
or U3779 (N_3779,N_2437,N_2888);
or U3780 (N_3780,N_2687,N_2004);
nand U3781 (N_3781,N_2808,N_2709);
and U3782 (N_3782,N_2938,N_2773);
nor U3783 (N_3783,N_2736,N_2134);
or U3784 (N_3784,N_2432,N_2522);
nor U3785 (N_3785,N_2794,N_2063);
and U3786 (N_3786,N_2463,N_2805);
nand U3787 (N_3787,N_2094,N_2316);
and U3788 (N_3788,N_2324,N_2535);
and U3789 (N_3789,N_2810,N_2181);
and U3790 (N_3790,N_2554,N_2900);
nor U3791 (N_3791,N_2155,N_2614);
or U3792 (N_3792,N_2273,N_2475);
xor U3793 (N_3793,N_2204,N_2647);
nand U3794 (N_3794,N_2422,N_2262);
or U3795 (N_3795,N_2133,N_2758);
and U3796 (N_3796,N_2283,N_2784);
and U3797 (N_3797,N_2998,N_2131);
or U3798 (N_3798,N_2009,N_2264);
and U3799 (N_3799,N_2646,N_2778);
or U3800 (N_3800,N_2185,N_2076);
and U3801 (N_3801,N_2875,N_2937);
or U3802 (N_3802,N_2170,N_2685);
nand U3803 (N_3803,N_2086,N_2617);
nor U3804 (N_3804,N_2829,N_2276);
nor U3805 (N_3805,N_2255,N_2315);
or U3806 (N_3806,N_2208,N_2221);
and U3807 (N_3807,N_2268,N_2135);
xor U3808 (N_3808,N_2625,N_2863);
or U3809 (N_3809,N_2153,N_2922);
nor U3810 (N_3810,N_2611,N_2479);
nor U3811 (N_3811,N_2913,N_2391);
and U3812 (N_3812,N_2724,N_2837);
nor U3813 (N_3813,N_2835,N_2130);
xnor U3814 (N_3814,N_2590,N_2697);
and U3815 (N_3815,N_2362,N_2211);
xor U3816 (N_3816,N_2024,N_2295);
nand U3817 (N_3817,N_2198,N_2016);
and U3818 (N_3818,N_2411,N_2294);
nand U3819 (N_3819,N_2650,N_2314);
and U3820 (N_3820,N_2890,N_2479);
nand U3821 (N_3821,N_2278,N_2464);
nor U3822 (N_3822,N_2667,N_2003);
and U3823 (N_3823,N_2749,N_2383);
and U3824 (N_3824,N_2690,N_2110);
nand U3825 (N_3825,N_2645,N_2816);
or U3826 (N_3826,N_2169,N_2572);
nor U3827 (N_3827,N_2065,N_2706);
xnor U3828 (N_3828,N_2489,N_2388);
nor U3829 (N_3829,N_2855,N_2191);
and U3830 (N_3830,N_2508,N_2469);
or U3831 (N_3831,N_2736,N_2366);
and U3832 (N_3832,N_2089,N_2777);
nor U3833 (N_3833,N_2900,N_2663);
and U3834 (N_3834,N_2165,N_2067);
or U3835 (N_3835,N_2491,N_2215);
and U3836 (N_3836,N_2993,N_2575);
and U3837 (N_3837,N_2559,N_2817);
and U3838 (N_3838,N_2375,N_2314);
nor U3839 (N_3839,N_2752,N_2389);
and U3840 (N_3840,N_2799,N_2385);
nand U3841 (N_3841,N_2909,N_2974);
nor U3842 (N_3842,N_2971,N_2613);
nand U3843 (N_3843,N_2936,N_2260);
nand U3844 (N_3844,N_2608,N_2863);
xnor U3845 (N_3845,N_2135,N_2610);
nand U3846 (N_3846,N_2563,N_2184);
nor U3847 (N_3847,N_2871,N_2022);
nand U3848 (N_3848,N_2252,N_2570);
or U3849 (N_3849,N_2359,N_2473);
or U3850 (N_3850,N_2578,N_2927);
or U3851 (N_3851,N_2638,N_2318);
nor U3852 (N_3852,N_2546,N_2346);
nand U3853 (N_3853,N_2713,N_2083);
or U3854 (N_3854,N_2662,N_2469);
nand U3855 (N_3855,N_2000,N_2284);
nor U3856 (N_3856,N_2054,N_2317);
nand U3857 (N_3857,N_2416,N_2717);
xor U3858 (N_3858,N_2759,N_2490);
nand U3859 (N_3859,N_2216,N_2517);
and U3860 (N_3860,N_2173,N_2860);
or U3861 (N_3861,N_2166,N_2039);
nand U3862 (N_3862,N_2808,N_2917);
and U3863 (N_3863,N_2755,N_2253);
nand U3864 (N_3864,N_2034,N_2014);
or U3865 (N_3865,N_2876,N_2394);
or U3866 (N_3866,N_2410,N_2708);
or U3867 (N_3867,N_2238,N_2986);
nand U3868 (N_3868,N_2685,N_2683);
or U3869 (N_3869,N_2294,N_2382);
and U3870 (N_3870,N_2731,N_2085);
nor U3871 (N_3871,N_2688,N_2710);
nor U3872 (N_3872,N_2981,N_2645);
and U3873 (N_3873,N_2740,N_2698);
or U3874 (N_3874,N_2578,N_2637);
nor U3875 (N_3875,N_2995,N_2494);
nor U3876 (N_3876,N_2173,N_2808);
and U3877 (N_3877,N_2059,N_2812);
xnor U3878 (N_3878,N_2805,N_2434);
and U3879 (N_3879,N_2317,N_2461);
nand U3880 (N_3880,N_2724,N_2220);
or U3881 (N_3881,N_2261,N_2753);
nand U3882 (N_3882,N_2976,N_2402);
xor U3883 (N_3883,N_2555,N_2561);
nand U3884 (N_3884,N_2631,N_2227);
and U3885 (N_3885,N_2821,N_2138);
nand U3886 (N_3886,N_2947,N_2984);
nor U3887 (N_3887,N_2985,N_2917);
nand U3888 (N_3888,N_2447,N_2779);
nor U3889 (N_3889,N_2731,N_2511);
xor U3890 (N_3890,N_2730,N_2381);
and U3891 (N_3891,N_2665,N_2850);
nor U3892 (N_3892,N_2509,N_2629);
and U3893 (N_3893,N_2699,N_2419);
nand U3894 (N_3894,N_2453,N_2941);
nand U3895 (N_3895,N_2023,N_2093);
nor U3896 (N_3896,N_2128,N_2097);
or U3897 (N_3897,N_2502,N_2956);
and U3898 (N_3898,N_2918,N_2223);
or U3899 (N_3899,N_2561,N_2017);
nand U3900 (N_3900,N_2206,N_2832);
and U3901 (N_3901,N_2047,N_2751);
nand U3902 (N_3902,N_2071,N_2653);
nand U3903 (N_3903,N_2857,N_2684);
or U3904 (N_3904,N_2830,N_2378);
nor U3905 (N_3905,N_2683,N_2451);
or U3906 (N_3906,N_2843,N_2336);
or U3907 (N_3907,N_2162,N_2976);
nand U3908 (N_3908,N_2591,N_2149);
or U3909 (N_3909,N_2391,N_2871);
nor U3910 (N_3910,N_2655,N_2214);
or U3911 (N_3911,N_2436,N_2107);
or U3912 (N_3912,N_2842,N_2652);
and U3913 (N_3913,N_2973,N_2163);
nand U3914 (N_3914,N_2261,N_2422);
and U3915 (N_3915,N_2429,N_2170);
and U3916 (N_3916,N_2328,N_2092);
xor U3917 (N_3917,N_2097,N_2975);
and U3918 (N_3918,N_2085,N_2766);
and U3919 (N_3919,N_2128,N_2952);
and U3920 (N_3920,N_2705,N_2792);
or U3921 (N_3921,N_2840,N_2353);
nor U3922 (N_3922,N_2659,N_2071);
xnor U3923 (N_3923,N_2142,N_2066);
nor U3924 (N_3924,N_2088,N_2582);
xor U3925 (N_3925,N_2038,N_2229);
and U3926 (N_3926,N_2294,N_2060);
nand U3927 (N_3927,N_2477,N_2605);
nand U3928 (N_3928,N_2052,N_2391);
nor U3929 (N_3929,N_2642,N_2600);
and U3930 (N_3930,N_2107,N_2118);
or U3931 (N_3931,N_2031,N_2010);
and U3932 (N_3932,N_2277,N_2372);
and U3933 (N_3933,N_2748,N_2770);
nand U3934 (N_3934,N_2651,N_2010);
and U3935 (N_3935,N_2631,N_2418);
or U3936 (N_3936,N_2211,N_2748);
nor U3937 (N_3937,N_2184,N_2339);
or U3938 (N_3938,N_2956,N_2118);
or U3939 (N_3939,N_2163,N_2394);
nor U3940 (N_3940,N_2746,N_2385);
or U3941 (N_3941,N_2010,N_2377);
and U3942 (N_3942,N_2362,N_2892);
nand U3943 (N_3943,N_2336,N_2832);
and U3944 (N_3944,N_2036,N_2180);
xor U3945 (N_3945,N_2359,N_2097);
xnor U3946 (N_3946,N_2564,N_2135);
and U3947 (N_3947,N_2070,N_2396);
or U3948 (N_3948,N_2491,N_2785);
nand U3949 (N_3949,N_2847,N_2943);
and U3950 (N_3950,N_2102,N_2452);
nand U3951 (N_3951,N_2100,N_2979);
and U3952 (N_3952,N_2246,N_2831);
nand U3953 (N_3953,N_2242,N_2446);
or U3954 (N_3954,N_2731,N_2775);
nand U3955 (N_3955,N_2252,N_2758);
nand U3956 (N_3956,N_2674,N_2466);
xor U3957 (N_3957,N_2113,N_2319);
xnor U3958 (N_3958,N_2703,N_2960);
nor U3959 (N_3959,N_2901,N_2847);
nand U3960 (N_3960,N_2131,N_2667);
nand U3961 (N_3961,N_2293,N_2401);
or U3962 (N_3962,N_2389,N_2860);
and U3963 (N_3963,N_2156,N_2265);
nand U3964 (N_3964,N_2035,N_2640);
xnor U3965 (N_3965,N_2993,N_2119);
xor U3966 (N_3966,N_2431,N_2898);
nor U3967 (N_3967,N_2562,N_2731);
nor U3968 (N_3968,N_2019,N_2708);
xor U3969 (N_3969,N_2538,N_2473);
xnor U3970 (N_3970,N_2859,N_2100);
or U3971 (N_3971,N_2129,N_2275);
and U3972 (N_3972,N_2821,N_2028);
nand U3973 (N_3973,N_2404,N_2268);
or U3974 (N_3974,N_2724,N_2735);
and U3975 (N_3975,N_2040,N_2744);
and U3976 (N_3976,N_2408,N_2462);
or U3977 (N_3977,N_2129,N_2186);
or U3978 (N_3978,N_2422,N_2548);
nand U3979 (N_3979,N_2248,N_2722);
nor U3980 (N_3980,N_2293,N_2415);
nor U3981 (N_3981,N_2487,N_2798);
xnor U3982 (N_3982,N_2852,N_2118);
nand U3983 (N_3983,N_2898,N_2662);
nand U3984 (N_3984,N_2785,N_2607);
xor U3985 (N_3985,N_2028,N_2446);
and U3986 (N_3986,N_2815,N_2900);
nand U3987 (N_3987,N_2318,N_2553);
nand U3988 (N_3988,N_2743,N_2159);
and U3989 (N_3989,N_2097,N_2348);
nand U3990 (N_3990,N_2971,N_2711);
or U3991 (N_3991,N_2155,N_2409);
or U3992 (N_3992,N_2418,N_2114);
and U3993 (N_3993,N_2454,N_2775);
xor U3994 (N_3994,N_2367,N_2352);
xor U3995 (N_3995,N_2315,N_2258);
nand U3996 (N_3996,N_2757,N_2995);
or U3997 (N_3997,N_2425,N_2646);
xor U3998 (N_3998,N_2447,N_2006);
nand U3999 (N_3999,N_2699,N_2723);
or U4000 (N_4000,N_3687,N_3260);
nor U4001 (N_4001,N_3399,N_3437);
nand U4002 (N_4002,N_3182,N_3164);
or U4003 (N_4003,N_3178,N_3404);
nand U4004 (N_4004,N_3357,N_3822);
or U4005 (N_4005,N_3225,N_3762);
and U4006 (N_4006,N_3813,N_3317);
nor U4007 (N_4007,N_3018,N_3415);
nand U4008 (N_4008,N_3603,N_3942);
nand U4009 (N_4009,N_3433,N_3533);
nand U4010 (N_4010,N_3914,N_3755);
nand U4011 (N_4011,N_3016,N_3551);
nand U4012 (N_4012,N_3382,N_3778);
nand U4013 (N_4013,N_3936,N_3593);
nand U4014 (N_4014,N_3445,N_3535);
nand U4015 (N_4015,N_3974,N_3147);
nor U4016 (N_4016,N_3229,N_3076);
or U4017 (N_4017,N_3262,N_3792);
or U4018 (N_4018,N_3060,N_3666);
nand U4019 (N_4019,N_3042,N_3215);
nand U4020 (N_4020,N_3814,N_3347);
or U4021 (N_4021,N_3746,N_3854);
nand U4022 (N_4022,N_3572,N_3150);
or U4023 (N_4023,N_3568,N_3406);
or U4024 (N_4024,N_3155,N_3723);
nor U4025 (N_4025,N_3876,N_3092);
nand U4026 (N_4026,N_3311,N_3906);
or U4027 (N_4027,N_3167,N_3017);
and U4028 (N_4028,N_3096,N_3693);
and U4029 (N_4029,N_3239,N_3964);
nand U4030 (N_4030,N_3629,N_3313);
nand U4031 (N_4031,N_3475,N_3349);
and U4032 (N_4032,N_3645,N_3634);
or U4033 (N_4033,N_3102,N_3495);
nand U4034 (N_4034,N_3704,N_3412);
and U4035 (N_4035,N_3385,N_3486);
and U4036 (N_4036,N_3230,N_3049);
or U4037 (N_4037,N_3789,N_3391);
nand U4038 (N_4038,N_3536,N_3576);
nor U4039 (N_4039,N_3829,N_3488);
xor U4040 (N_4040,N_3882,N_3885);
xor U4041 (N_4041,N_3968,N_3756);
xor U4042 (N_4042,N_3440,N_3760);
nor U4043 (N_4043,N_3994,N_3900);
or U4044 (N_4044,N_3548,N_3569);
and U4045 (N_4045,N_3821,N_3432);
and U4046 (N_4046,N_3923,N_3967);
nor U4047 (N_4047,N_3483,N_3720);
nor U4048 (N_4048,N_3421,N_3013);
nor U4049 (N_4049,N_3872,N_3101);
and U4050 (N_4050,N_3851,N_3428);
or U4051 (N_4051,N_3545,N_3157);
nand U4052 (N_4052,N_3636,N_3958);
nor U4053 (N_4053,N_3052,N_3701);
nand U4054 (N_4054,N_3862,N_3615);
and U4055 (N_4055,N_3716,N_3749);
xor U4056 (N_4056,N_3763,N_3894);
nand U4057 (N_4057,N_3090,N_3099);
nand U4058 (N_4058,N_3361,N_3857);
and U4059 (N_4059,N_3933,N_3546);
nor U4060 (N_4060,N_3087,N_3422);
nor U4061 (N_4061,N_3863,N_3330);
or U4062 (N_4062,N_3920,N_3118);
nand U4063 (N_4063,N_3142,N_3633);
and U4064 (N_4064,N_3670,N_3580);
nor U4065 (N_4065,N_3761,N_3237);
and U4066 (N_4066,N_3158,N_3075);
or U4067 (N_4067,N_3318,N_3344);
or U4068 (N_4068,N_3736,N_3590);
nor U4069 (N_4069,N_3977,N_3714);
nand U4070 (N_4070,N_3310,N_3588);
or U4071 (N_4071,N_3125,N_3040);
xnor U4072 (N_4072,N_3825,N_3655);
xnor U4073 (N_4073,N_3992,N_3915);
nand U4074 (N_4074,N_3784,N_3146);
nor U4075 (N_4075,N_3035,N_3517);
nor U4076 (N_4076,N_3667,N_3256);
nor U4077 (N_4077,N_3812,N_3613);
and U4078 (N_4078,N_3774,N_3355);
or U4079 (N_4079,N_3343,N_3441);
xor U4080 (N_4080,N_3161,N_3932);
or U4081 (N_4081,N_3029,N_3168);
or U4082 (N_4082,N_3115,N_3531);
or U4083 (N_4083,N_3238,N_3631);
and U4084 (N_4084,N_3520,N_3621);
and U4085 (N_4085,N_3703,N_3485);
nor U4086 (N_4086,N_3446,N_3254);
and U4087 (N_4087,N_3316,N_3975);
or U4088 (N_4088,N_3773,N_3322);
or U4089 (N_4089,N_3165,N_3985);
and U4090 (N_4090,N_3053,N_3148);
and U4091 (N_4091,N_3650,N_3356);
and U4092 (N_4092,N_3348,N_3541);
xnor U4093 (N_4093,N_3328,N_3635);
nor U4094 (N_4094,N_3242,N_3396);
and U4095 (N_4095,N_3031,N_3791);
and U4096 (N_4096,N_3700,N_3103);
or U4097 (N_4097,N_3695,N_3525);
xnor U4098 (N_4098,N_3561,N_3392);
nand U4099 (N_4099,N_3290,N_3886);
nand U4100 (N_4100,N_3847,N_3279);
or U4101 (N_4101,N_3608,N_3518);
and U4102 (N_4102,N_3033,N_3506);
and U4103 (N_4103,N_3649,N_3278);
or U4104 (N_4104,N_3001,N_3221);
nor U4105 (N_4105,N_3307,N_3516);
and U4106 (N_4106,N_3071,N_3481);
xor U4107 (N_4107,N_3637,N_3869);
and U4108 (N_4108,N_3331,N_3418);
nand U4109 (N_4109,N_3827,N_3524);
and U4110 (N_4110,N_3450,N_3617);
nor U4111 (N_4111,N_3837,N_3680);
nor U4112 (N_4112,N_3039,N_3939);
nand U4113 (N_4113,N_3751,N_3627);
nor U4114 (N_4114,N_3610,N_3258);
xor U4115 (N_4115,N_3362,N_3091);
and U4116 (N_4116,N_3934,N_3803);
and U4117 (N_4117,N_3032,N_3339);
xor U4118 (N_4118,N_3235,N_3000);
or U4119 (N_4119,N_3351,N_3757);
or U4120 (N_4120,N_3086,N_3259);
nor U4121 (N_4121,N_3494,N_3137);
and U4122 (N_4122,N_3389,N_3319);
or U4123 (N_4123,N_3298,N_3810);
or U4124 (N_4124,N_3771,N_3336);
nor U4125 (N_4125,N_3009,N_3194);
and U4126 (N_4126,N_3346,N_3998);
nand U4127 (N_4127,N_3873,N_3891);
and U4128 (N_4128,N_3304,N_3175);
nand U4129 (N_4129,N_3456,N_3640);
and U4130 (N_4130,N_3400,N_3880);
and U4131 (N_4131,N_3881,N_3135);
and U4132 (N_4132,N_3870,N_3947);
nor U4133 (N_4133,N_3973,N_3542);
nor U4134 (N_4134,N_3180,N_3529);
nor U4135 (N_4135,N_3962,N_3941);
nor U4136 (N_4136,N_3474,N_3677);
nor U4137 (N_4137,N_3832,N_3471);
or U4138 (N_4138,N_3735,N_3333);
and U4139 (N_4139,N_3373,N_3315);
or U4140 (N_4140,N_3149,N_3989);
nand U4141 (N_4141,N_3372,N_3390);
nand U4142 (N_4142,N_3275,N_3019);
xnor U4143 (N_4143,N_3402,N_3370);
nor U4144 (N_4144,N_3758,N_3713);
nor U4145 (N_4145,N_3338,N_3671);
nand U4146 (N_4146,N_3583,N_3850);
nand U4147 (N_4147,N_3381,N_3438);
xnor U4148 (N_4148,N_3658,N_3079);
nor U4149 (N_4149,N_3276,N_3856);
nor U4150 (N_4150,N_3470,N_3683);
nand U4151 (N_4151,N_3765,N_3136);
and U4152 (N_4152,N_3253,N_3011);
or U4153 (N_4153,N_3151,N_3416);
xnor U4154 (N_4154,N_3543,N_3782);
or U4155 (N_4155,N_3449,N_3620);
and U4156 (N_4156,N_3114,N_3405);
and U4157 (N_4157,N_3597,N_3377);
nor U4158 (N_4158,N_3638,N_3503);
nor U4159 (N_4159,N_3741,N_3309);
and U4160 (N_4160,N_3965,N_3661);
or U4161 (N_4161,N_3840,N_3606);
nor U4162 (N_4162,N_3820,N_3860);
and U4163 (N_4163,N_3795,N_3173);
nor U4164 (N_4164,N_3398,N_3823);
nor U4165 (N_4165,N_3224,N_3783);
nand U4166 (N_4166,N_3705,N_3190);
nand U4167 (N_4167,N_3248,N_3826);
nand U4168 (N_4168,N_3255,N_3679);
nor U4169 (N_4169,N_3499,N_3896);
nand U4170 (N_4170,N_3501,N_3243);
xor U4171 (N_4171,N_3326,N_3464);
nand U4172 (N_4172,N_3508,N_3984);
or U4173 (N_4173,N_3996,N_3707);
nor U4174 (N_4174,N_3497,N_3916);
and U4175 (N_4175,N_3754,N_3830);
nor U4176 (N_4176,N_3133,N_3271);
xor U4177 (N_4177,N_3805,N_3043);
and U4178 (N_4178,N_3628,N_3024);
nor U4179 (N_4179,N_3244,N_3554);
or U4180 (N_4180,N_3417,N_3345);
nand U4181 (N_4181,N_3106,N_3077);
and U4182 (N_4182,N_3653,N_3815);
nand U4183 (N_4183,N_3489,N_3144);
or U4184 (N_4184,N_3866,N_3630);
and U4185 (N_4185,N_3972,N_3786);
and U4186 (N_4186,N_3948,N_3265);
and U4187 (N_4187,N_3817,N_3552);
nand U4188 (N_4188,N_3510,N_3919);
nor U4189 (N_4189,N_3112,N_3549);
nor U4190 (N_4190,N_3393,N_3200);
and U4191 (N_4191,N_3387,N_3193);
and U4192 (N_4192,N_3469,N_3587);
and U4193 (N_4193,N_3420,N_3080);
and U4194 (N_4194,N_3512,N_3515);
nand U4195 (N_4195,N_3216,N_3245);
nand U4196 (N_4196,N_3970,N_3544);
or U4197 (N_4197,N_3988,N_3409);
nor U4198 (N_4198,N_3879,N_3883);
nand U4199 (N_4199,N_3166,N_3159);
nor U4200 (N_4200,N_3663,N_3287);
and U4201 (N_4201,N_3240,N_3884);
and U4202 (N_4202,N_3505,N_3971);
xor U4203 (N_4203,N_3204,N_3066);
or U4204 (N_4204,N_3849,N_3668);
nand U4205 (N_4205,N_3824,N_3777);
nor U4206 (N_4206,N_3674,N_3284);
and U4207 (N_4207,N_3601,N_3926);
nand U4208 (N_4208,N_3946,N_3526);
and U4209 (N_4209,N_3726,N_3776);
nand U4210 (N_4210,N_3547,N_3123);
nor U4211 (N_4211,N_3500,N_3156);
and U4212 (N_4212,N_3599,N_3027);
and U4213 (N_4213,N_3108,N_3838);
and U4214 (N_4214,N_3051,N_3478);
xnor U4215 (N_4215,N_3111,N_3472);
and U4216 (N_4216,N_3227,N_3797);
and U4217 (N_4217,N_3183,N_3068);
nand U4218 (N_4218,N_3145,N_3902);
and U4219 (N_4219,N_3767,N_3203);
nand U4220 (N_4220,N_3129,N_3314);
or U4221 (N_4221,N_3431,N_3944);
xor U4222 (N_4222,N_3711,N_3274);
nand U4223 (N_4223,N_3796,N_3565);
nand U4224 (N_4224,N_3046,N_3069);
and U4225 (N_4225,N_3047,N_3575);
or U4226 (N_4226,N_3192,N_3467);
nand U4227 (N_4227,N_3045,N_3555);
and U4228 (N_4228,N_3198,N_3234);
and U4229 (N_4229,N_3350,N_3249);
nor U4230 (N_4230,N_3898,N_3586);
nor U4231 (N_4231,N_3689,N_3522);
and U4232 (N_4232,N_3953,N_3266);
nor U4233 (N_4233,N_3940,N_3727);
nor U4234 (N_4234,N_3878,N_3935);
and U4235 (N_4235,N_3913,N_3448);
and U4236 (N_4236,N_3537,N_3960);
nor U4237 (N_4237,N_3864,N_3181);
nand U4238 (N_4238,N_3081,N_3063);
nand U4239 (N_4239,N_3745,N_3162);
or U4240 (N_4240,N_3380,N_3987);
xor U4241 (N_4241,N_3577,N_3956);
or U4242 (N_4242,N_3834,N_3798);
nand U4243 (N_4243,N_3624,N_3534);
and U4244 (N_4244,N_3458,N_3366);
and U4245 (N_4245,N_3059,N_3995);
or U4246 (N_4246,N_3859,N_3731);
or U4247 (N_4247,N_3335,N_3766);
nand U4248 (N_4248,N_3187,N_3951);
or U4249 (N_4249,N_3116,N_3360);
xor U4250 (N_4250,N_3073,N_3020);
xnor U4251 (N_4251,N_3616,N_3408);
and U4252 (N_4252,N_3447,N_3223);
and U4253 (N_4253,N_3574,N_3899);
and U4254 (N_4254,N_3799,N_3868);
xnor U4255 (N_4255,N_3890,N_3006);
or U4256 (N_4256,N_3539,N_3528);
or U4257 (N_4257,N_3744,N_3130);
and U4258 (N_4258,N_3261,N_3787);
xnor U4259 (N_4259,N_3476,N_3591);
or U4260 (N_4260,N_3678,N_3191);
and U4261 (N_4261,N_3365,N_3186);
nor U4262 (N_4262,N_3589,N_3806);
xor U4263 (N_4263,N_3003,N_3981);
nor U4264 (N_4264,N_3270,N_3690);
and U4265 (N_4265,N_3300,N_3490);
nand U4266 (N_4266,N_3341,N_3600);
nand U4267 (N_4267,N_3930,N_3665);
nand U4268 (N_4268,N_3918,N_3169);
nor U4269 (N_4269,N_3607,N_3354);
or U4270 (N_4270,N_3559,N_3581);
and U4271 (N_4271,N_3550,N_3057);
and U4272 (N_4272,N_3131,N_3231);
nand U4273 (N_4273,N_3504,N_3295);
nand U4274 (N_4274,N_3005,N_3044);
nor U4275 (N_4275,N_3945,N_3436);
nor U4276 (N_4276,N_3853,N_3014);
nor U4277 (N_4277,N_3519,N_3836);
xor U4278 (N_4278,N_3289,N_3811);
or U4279 (N_4279,N_3395,N_3263);
xnor U4280 (N_4280,N_3435,N_3807);
nor U4281 (N_4281,N_3513,N_3054);
nand U4282 (N_4282,N_3511,N_3124);
or U4283 (N_4283,N_3493,N_3160);
nand U4284 (N_4284,N_3764,N_3434);
or U4285 (N_4285,N_3062,N_3648);
and U4286 (N_4286,N_3222,N_3922);
nor U4287 (N_4287,N_3685,N_3457);
nand U4288 (N_4288,N_3277,N_3728);
nand U4289 (N_4289,N_3604,N_3562);
or U4290 (N_4290,N_3329,N_3775);
nor U4291 (N_4291,N_3943,N_3122);
xor U4292 (N_4292,N_3911,N_3904);
nand U4293 (N_4293,N_3285,N_3491);
xnor U4294 (N_4294,N_3925,N_3921);
nand U4295 (N_4295,N_3781,N_3502);
or U4296 (N_4296,N_3770,N_3573);
xor U4297 (N_4297,N_3403,N_3163);
and U4298 (N_4298,N_3938,N_3273);
xnor U4299 (N_4299,N_3595,N_3578);
nor U4300 (N_4300,N_3927,N_3246);
and U4301 (N_4301,N_3117,N_3734);
or U4302 (N_4302,N_3219,N_3492);
or U4303 (N_4303,N_3733,N_3107);
or U4304 (N_4304,N_3041,N_3632);
or U4305 (N_4305,N_3672,N_3895);
nor U4306 (N_4306,N_3785,N_3247);
nor U4307 (N_4307,N_3819,N_3954);
nand U4308 (N_4308,N_3909,N_3109);
or U4309 (N_4309,N_3657,N_3937);
nor U4310 (N_4310,N_3132,N_3455);
or U4311 (N_4311,N_3839,N_3769);
nand U4312 (N_4312,N_3852,N_3557);
and U4313 (N_4313,N_3523,N_3702);
and U4314 (N_4314,N_3401,N_3719);
nand U4315 (N_4315,N_3082,N_3567);
nor U4316 (N_4316,N_3089,N_3012);
or U4317 (N_4317,N_3085,N_3384);
nand U4318 (N_4318,N_3217,N_3056);
or U4319 (N_4319,N_3291,N_3722);
xor U4320 (N_4320,N_3748,N_3461);
nand U4321 (N_4321,N_3367,N_3507);
and U4322 (N_4322,N_3451,N_3571);
or U4323 (N_4323,N_3188,N_3997);
nand U4324 (N_4324,N_3171,N_3842);
nor U4325 (N_4325,N_3639,N_3718);
and U4326 (N_4326,N_3538,N_3496);
nand U4327 (N_4327,N_3065,N_3966);
nor U4328 (N_4328,N_3980,N_3364);
nor U4329 (N_4329,N_3058,N_3871);
and U4330 (N_4330,N_3865,N_3780);
nor U4331 (N_4331,N_3250,N_3267);
nand U4332 (N_4332,N_3023,N_3208);
and U4333 (N_4333,N_3477,N_3321);
or U4334 (N_4334,N_3213,N_3293);
nand U4335 (N_4335,N_3730,N_3473);
nand U4336 (N_4336,N_3397,N_3721);
xor U4337 (N_4337,N_3206,N_3297);
nor U4338 (N_4338,N_3582,N_3241);
nand U4339 (N_4339,N_3750,N_3197);
or U4340 (N_4340,N_3908,N_3479);
and U4341 (N_4341,N_3596,N_3498);
or U4342 (N_4342,N_3306,N_3611);
nand U4343 (N_4343,N_3463,N_3867);
or U4344 (N_4344,N_3609,N_3026);
nor U4345 (N_4345,N_3623,N_3753);
nand U4346 (N_4346,N_3742,N_3154);
nand U4347 (N_4347,N_3729,N_3585);
nor U4348 (N_4348,N_3682,N_3050);
and U4349 (N_4349,N_3236,N_3592);
or U4350 (N_4350,N_3738,N_3218);
xnor U4351 (N_4351,N_3694,N_3978);
nor U4352 (N_4352,N_3715,N_3022);
nand U4353 (N_4353,N_3340,N_3959);
xnor U4354 (N_4354,N_3453,N_3861);
nor U4355 (N_4355,N_3579,N_3374);
or U4356 (N_4356,N_3618,N_3654);
and U4357 (N_4357,N_3647,N_3028);
or U4358 (N_4358,N_3901,N_3675);
and U4359 (N_4359,N_3211,N_3696);
and U4360 (N_4360,N_3907,N_3929);
and U4361 (N_4361,N_3303,N_3025);
and U4362 (N_4362,N_3570,N_3686);
xor U4363 (N_4363,N_3425,N_3207);
and U4364 (N_4364,N_3369,N_3527);
and U4365 (N_4365,N_3015,N_3443);
or U4366 (N_4366,N_3681,N_3323);
xnor U4367 (N_4367,N_3530,N_3413);
and U4368 (N_4368,N_3036,N_3961);
nand U4369 (N_4369,N_3414,N_3843);
nor U4370 (N_4370,N_3252,N_3324);
or U4371 (N_4371,N_3835,N_3113);
and U4372 (N_4372,N_3100,N_3141);
xor U4373 (N_4373,N_3622,N_3706);
nand U4374 (N_4374,N_3305,N_3281);
nor U4375 (N_4375,N_3912,N_3893);
xnor U4376 (N_4376,N_3359,N_3386);
or U4377 (N_4377,N_3626,N_3790);
or U4378 (N_4378,N_3083,N_3688);
and U4379 (N_4379,N_3692,N_3875);
xnor U4380 (N_4380,N_3201,N_3139);
or U4381 (N_4381,N_3283,N_3427);
nand U4382 (N_4382,N_3272,N_3802);
or U4383 (N_4383,N_3002,N_3625);
or U4384 (N_4384,N_3352,N_3462);
or U4385 (N_4385,N_3072,N_3388);
nor U4386 (N_4386,N_3264,N_3656);
or U4387 (N_4387,N_3383,N_3659);
xor U4388 (N_4388,N_3067,N_3325);
nor U4389 (N_4389,N_3845,N_3743);
nor U4390 (N_4390,N_3664,N_3566);
xor U4391 (N_4391,N_3917,N_3378);
nor U4392 (N_4392,N_3286,N_3642);
nor U4393 (N_4393,N_3710,N_3999);
or U4394 (N_4394,N_3982,N_3084);
and U4395 (N_4395,N_3292,N_3140);
or U4396 (N_4396,N_3509,N_3152);
or U4397 (N_4397,N_3897,N_3119);
or U4398 (N_4398,N_3482,N_3189);
and U4399 (N_4399,N_3521,N_3093);
and U4400 (N_4400,N_3128,N_3794);
and U4401 (N_4401,N_3430,N_3220);
nand U4402 (N_4402,N_3717,N_3732);
and U4403 (N_4403,N_3233,N_3174);
xnor U4404 (N_4404,N_3444,N_3110);
or U4405 (N_4405,N_3480,N_3979);
or U4406 (N_4406,N_3127,N_3889);
and U4407 (N_4407,N_3251,N_3368);
or U4408 (N_4408,N_3134,N_3143);
nand U4409 (N_4409,N_3739,N_3419);
nand U4410 (N_4410,N_3514,N_3487);
nand U4411 (N_4411,N_3021,N_3088);
nand U4412 (N_4412,N_3800,N_3594);
and U4413 (N_4413,N_3424,N_3963);
nand U4414 (N_4414,N_3990,N_3818);
or U4415 (N_4415,N_3848,N_3226);
xnor U4416 (N_4416,N_3691,N_3740);
nand U4417 (N_4417,N_3429,N_3185);
or U4418 (N_4418,N_3153,N_3358);
nor U4419 (N_4419,N_3724,N_3905);
nor U4420 (N_4420,N_3651,N_3120);
nand U4421 (N_4421,N_3268,N_3176);
nor U4422 (N_4422,N_3643,N_3179);
nand U4423 (N_4423,N_3983,N_3804);
nor U4424 (N_4424,N_3737,N_3196);
or U4425 (N_4425,N_3676,N_3342);
or U4426 (N_4426,N_3708,N_3602);
nand U4427 (N_4427,N_3646,N_3105);
nand U4428 (N_4428,N_3375,N_3327);
nand U4429 (N_4429,N_3652,N_3928);
xor U4430 (N_4430,N_3210,N_3888);
xor U4431 (N_4431,N_3055,N_3465);
nor U4432 (N_4432,N_3949,N_3779);
nand U4433 (N_4433,N_3170,N_3078);
or U4434 (N_4434,N_3184,N_3684);
or U4435 (N_4435,N_3007,N_3121);
nand U4436 (N_4436,N_3376,N_3070);
and U4437 (N_4437,N_3008,N_3752);
or U4438 (N_4438,N_3903,N_3605);
and U4439 (N_4439,N_3048,N_3712);
nor U4440 (N_4440,N_3104,N_3556);
or U4441 (N_4441,N_3379,N_3950);
xnor U4442 (N_4442,N_3177,N_3038);
nand U4443 (N_4443,N_3788,N_3612);
and U4444 (N_4444,N_3332,N_3484);
or U4445 (N_4445,N_3308,N_3199);
nand U4446 (N_4446,N_3614,N_3288);
or U4447 (N_4447,N_3097,N_3660);
nor U4448 (N_4448,N_3363,N_3172);
or U4449 (N_4449,N_3353,N_3010);
and U4450 (N_4450,N_3337,N_3976);
or U4451 (N_4451,N_3558,N_3924);
or U4452 (N_4452,N_3801,N_3004);
or U4453 (N_4453,N_3299,N_3892);
and U4454 (N_4454,N_3296,N_3410);
or U4455 (N_4455,N_3808,N_3202);
nor U4456 (N_4456,N_3816,N_3887);
nand U4457 (N_4457,N_3910,N_3301);
and U4458 (N_4458,N_3697,N_3991);
and U4459 (N_4459,N_3619,N_3257);
xnor U4460 (N_4460,N_3931,N_3641);
nor U4461 (N_4461,N_3772,N_3699);
nand U4462 (N_4462,N_3138,N_3560);
nor U4463 (N_4463,N_3439,N_3282);
xor U4464 (N_4464,N_3371,N_3747);
nor U4465 (N_4465,N_3205,N_3669);
or U4466 (N_4466,N_3294,N_3334);
nor U4467 (N_4467,N_3759,N_3563);
or U4468 (N_4468,N_3540,N_3232);
and U4469 (N_4469,N_3662,N_3095);
nor U4470 (N_4470,N_3320,N_3874);
and U4471 (N_4471,N_3407,N_3828);
nor U4472 (N_4472,N_3986,N_3037);
nand U4473 (N_4473,N_3459,N_3809);
nand U4474 (N_4474,N_3228,N_3877);
nor U4475 (N_4475,N_3466,N_3831);
and U4476 (N_4476,N_3768,N_3030);
and U4477 (N_4477,N_3725,N_3855);
nor U4478 (N_4478,N_3454,N_3841);
nand U4479 (N_4479,N_3426,N_3969);
nor U4480 (N_4480,N_3064,N_3993);
and U4481 (N_4481,N_3844,N_3564);
nand U4482 (N_4482,N_3452,N_3644);
nand U4483 (N_4483,N_3858,N_3074);
and U4484 (N_4484,N_3955,N_3098);
xor U4485 (N_4485,N_3957,N_3411);
nor U4486 (N_4486,N_3269,N_3673);
and U4487 (N_4487,N_3312,N_3302);
xnor U4488 (N_4488,N_3553,N_3212);
or U4489 (N_4489,N_3094,N_3280);
and U4490 (N_4490,N_3460,N_3061);
nand U4491 (N_4491,N_3846,N_3423);
and U4492 (N_4492,N_3195,N_3442);
or U4493 (N_4493,N_3598,N_3532);
nor U4494 (N_4494,N_3034,N_3214);
nand U4495 (N_4495,N_3126,N_3209);
nor U4496 (N_4496,N_3833,N_3394);
xnor U4497 (N_4497,N_3698,N_3468);
nand U4498 (N_4498,N_3709,N_3952);
and U4499 (N_4499,N_3793,N_3584);
nor U4500 (N_4500,N_3279,N_3961);
nor U4501 (N_4501,N_3004,N_3207);
nand U4502 (N_4502,N_3350,N_3729);
nand U4503 (N_4503,N_3830,N_3812);
nor U4504 (N_4504,N_3004,N_3470);
nor U4505 (N_4505,N_3110,N_3891);
nor U4506 (N_4506,N_3285,N_3334);
or U4507 (N_4507,N_3694,N_3085);
nor U4508 (N_4508,N_3451,N_3785);
nand U4509 (N_4509,N_3988,N_3433);
or U4510 (N_4510,N_3375,N_3231);
and U4511 (N_4511,N_3390,N_3285);
nor U4512 (N_4512,N_3775,N_3151);
or U4513 (N_4513,N_3990,N_3885);
or U4514 (N_4514,N_3078,N_3525);
or U4515 (N_4515,N_3394,N_3659);
and U4516 (N_4516,N_3234,N_3000);
nand U4517 (N_4517,N_3327,N_3539);
nand U4518 (N_4518,N_3941,N_3410);
and U4519 (N_4519,N_3331,N_3271);
nor U4520 (N_4520,N_3721,N_3573);
nand U4521 (N_4521,N_3932,N_3073);
nor U4522 (N_4522,N_3627,N_3048);
nand U4523 (N_4523,N_3996,N_3817);
and U4524 (N_4524,N_3174,N_3903);
xor U4525 (N_4525,N_3710,N_3554);
nor U4526 (N_4526,N_3409,N_3418);
and U4527 (N_4527,N_3658,N_3331);
and U4528 (N_4528,N_3985,N_3008);
or U4529 (N_4529,N_3848,N_3079);
nand U4530 (N_4530,N_3666,N_3436);
and U4531 (N_4531,N_3645,N_3315);
and U4532 (N_4532,N_3206,N_3746);
and U4533 (N_4533,N_3917,N_3314);
xor U4534 (N_4534,N_3420,N_3880);
nor U4535 (N_4535,N_3051,N_3739);
nor U4536 (N_4536,N_3219,N_3052);
and U4537 (N_4537,N_3398,N_3715);
nor U4538 (N_4538,N_3041,N_3749);
and U4539 (N_4539,N_3847,N_3351);
and U4540 (N_4540,N_3541,N_3148);
and U4541 (N_4541,N_3411,N_3047);
nor U4542 (N_4542,N_3742,N_3572);
or U4543 (N_4543,N_3424,N_3245);
xnor U4544 (N_4544,N_3968,N_3117);
xnor U4545 (N_4545,N_3245,N_3971);
xnor U4546 (N_4546,N_3271,N_3544);
or U4547 (N_4547,N_3681,N_3156);
and U4548 (N_4548,N_3365,N_3744);
and U4549 (N_4549,N_3460,N_3251);
nand U4550 (N_4550,N_3043,N_3295);
nor U4551 (N_4551,N_3897,N_3273);
xor U4552 (N_4552,N_3701,N_3535);
nand U4553 (N_4553,N_3899,N_3872);
nand U4554 (N_4554,N_3803,N_3135);
or U4555 (N_4555,N_3523,N_3032);
nand U4556 (N_4556,N_3568,N_3912);
or U4557 (N_4557,N_3268,N_3322);
and U4558 (N_4558,N_3712,N_3286);
nor U4559 (N_4559,N_3537,N_3371);
or U4560 (N_4560,N_3726,N_3160);
and U4561 (N_4561,N_3976,N_3289);
nor U4562 (N_4562,N_3635,N_3699);
nand U4563 (N_4563,N_3318,N_3445);
nor U4564 (N_4564,N_3039,N_3210);
and U4565 (N_4565,N_3738,N_3755);
and U4566 (N_4566,N_3896,N_3206);
nor U4567 (N_4567,N_3983,N_3751);
nor U4568 (N_4568,N_3538,N_3486);
and U4569 (N_4569,N_3998,N_3219);
nand U4570 (N_4570,N_3406,N_3484);
or U4571 (N_4571,N_3894,N_3493);
xnor U4572 (N_4572,N_3636,N_3582);
xor U4573 (N_4573,N_3530,N_3471);
or U4574 (N_4574,N_3548,N_3130);
nand U4575 (N_4575,N_3244,N_3490);
xnor U4576 (N_4576,N_3254,N_3821);
nand U4577 (N_4577,N_3712,N_3042);
and U4578 (N_4578,N_3287,N_3079);
and U4579 (N_4579,N_3687,N_3116);
nor U4580 (N_4580,N_3664,N_3863);
nand U4581 (N_4581,N_3047,N_3139);
and U4582 (N_4582,N_3985,N_3494);
nand U4583 (N_4583,N_3921,N_3462);
nor U4584 (N_4584,N_3722,N_3731);
and U4585 (N_4585,N_3276,N_3918);
nor U4586 (N_4586,N_3400,N_3467);
nand U4587 (N_4587,N_3850,N_3590);
and U4588 (N_4588,N_3216,N_3197);
xor U4589 (N_4589,N_3750,N_3349);
nand U4590 (N_4590,N_3722,N_3399);
nor U4591 (N_4591,N_3468,N_3748);
or U4592 (N_4592,N_3975,N_3554);
xor U4593 (N_4593,N_3404,N_3358);
and U4594 (N_4594,N_3746,N_3278);
and U4595 (N_4595,N_3162,N_3848);
or U4596 (N_4596,N_3626,N_3296);
or U4597 (N_4597,N_3391,N_3780);
or U4598 (N_4598,N_3315,N_3614);
and U4599 (N_4599,N_3882,N_3226);
nor U4600 (N_4600,N_3359,N_3778);
and U4601 (N_4601,N_3904,N_3408);
or U4602 (N_4602,N_3596,N_3147);
nand U4603 (N_4603,N_3335,N_3603);
nand U4604 (N_4604,N_3598,N_3892);
xnor U4605 (N_4605,N_3618,N_3122);
or U4606 (N_4606,N_3296,N_3189);
nand U4607 (N_4607,N_3832,N_3819);
nand U4608 (N_4608,N_3865,N_3530);
nand U4609 (N_4609,N_3063,N_3716);
nand U4610 (N_4610,N_3875,N_3174);
nor U4611 (N_4611,N_3295,N_3213);
and U4612 (N_4612,N_3670,N_3764);
nor U4613 (N_4613,N_3071,N_3195);
nand U4614 (N_4614,N_3931,N_3907);
nand U4615 (N_4615,N_3035,N_3864);
nand U4616 (N_4616,N_3409,N_3867);
nand U4617 (N_4617,N_3594,N_3698);
xnor U4618 (N_4618,N_3674,N_3173);
nand U4619 (N_4619,N_3942,N_3312);
nand U4620 (N_4620,N_3016,N_3783);
xor U4621 (N_4621,N_3755,N_3766);
and U4622 (N_4622,N_3034,N_3412);
nor U4623 (N_4623,N_3327,N_3444);
and U4624 (N_4624,N_3183,N_3187);
nand U4625 (N_4625,N_3547,N_3566);
nand U4626 (N_4626,N_3008,N_3934);
and U4627 (N_4627,N_3584,N_3977);
and U4628 (N_4628,N_3128,N_3015);
and U4629 (N_4629,N_3917,N_3935);
xnor U4630 (N_4630,N_3537,N_3413);
and U4631 (N_4631,N_3088,N_3375);
or U4632 (N_4632,N_3996,N_3057);
nand U4633 (N_4633,N_3158,N_3168);
nor U4634 (N_4634,N_3347,N_3949);
or U4635 (N_4635,N_3941,N_3366);
or U4636 (N_4636,N_3783,N_3967);
and U4637 (N_4637,N_3492,N_3805);
nor U4638 (N_4638,N_3495,N_3325);
and U4639 (N_4639,N_3749,N_3341);
and U4640 (N_4640,N_3172,N_3747);
or U4641 (N_4641,N_3830,N_3411);
or U4642 (N_4642,N_3968,N_3093);
or U4643 (N_4643,N_3582,N_3202);
nor U4644 (N_4644,N_3099,N_3698);
nor U4645 (N_4645,N_3985,N_3208);
and U4646 (N_4646,N_3945,N_3876);
nand U4647 (N_4647,N_3220,N_3208);
xor U4648 (N_4648,N_3392,N_3971);
or U4649 (N_4649,N_3575,N_3781);
nand U4650 (N_4650,N_3446,N_3564);
xnor U4651 (N_4651,N_3254,N_3527);
and U4652 (N_4652,N_3344,N_3529);
nand U4653 (N_4653,N_3374,N_3008);
nand U4654 (N_4654,N_3491,N_3795);
nor U4655 (N_4655,N_3725,N_3226);
nand U4656 (N_4656,N_3544,N_3968);
nand U4657 (N_4657,N_3386,N_3885);
nand U4658 (N_4658,N_3361,N_3582);
xor U4659 (N_4659,N_3853,N_3984);
and U4660 (N_4660,N_3474,N_3067);
nand U4661 (N_4661,N_3705,N_3049);
nand U4662 (N_4662,N_3682,N_3178);
nand U4663 (N_4663,N_3688,N_3829);
nor U4664 (N_4664,N_3610,N_3124);
nand U4665 (N_4665,N_3927,N_3202);
nor U4666 (N_4666,N_3768,N_3472);
or U4667 (N_4667,N_3214,N_3208);
nand U4668 (N_4668,N_3242,N_3864);
or U4669 (N_4669,N_3778,N_3953);
nor U4670 (N_4670,N_3108,N_3512);
xor U4671 (N_4671,N_3997,N_3436);
or U4672 (N_4672,N_3150,N_3686);
nor U4673 (N_4673,N_3666,N_3489);
or U4674 (N_4674,N_3797,N_3160);
nor U4675 (N_4675,N_3816,N_3953);
nand U4676 (N_4676,N_3838,N_3681);
nor U4677 (N_4677,N_3746,N_3717);
nor U4678 (N_4678,N_3681,N_3555);
nand U4679 (N_4679,N_3518,N_3823);
xnor U4680 (N_4680,N_3758,N_3159);
nand U4681 (N_4681,N_3942,N_3964);
and U4682 (N_4682,N_3441,N_3405);
nand U4683 (N_4683,N_3066,N_3975);
nor U4684 (N_4684,N_3764,N_3324);
xnor U4685 (N_4685,N_3546,N_3754);
nor U4686 (N_4686,N_3653,N_3746);
nand U4687 (N_4687,N_3197,N_3288);
nor U4688 (N_4688,N_3319,N_3065);
or U4689 (N_4689,N_3596,N_3132);
nand U4690 (N_4690,N_3088,N_3383);
or U4691 (N_4691,N_3745,N_3465);
xnor U4692 (N_4692,N_3638,N_3692);
and U4693 (N_4693,N_3590,N_3508);
and U4694 (N_4694,N_3702,N_3981);
xnor U4695 (N_4695,N_3589,N_3972);
or U4696 (N_4696,N_3620,N_3985);
nand U4697 (N_4697,N_3854,N_3982);
nor U4698 (N_4698,N_3348,N_3517);
nor U4699 (N_4699,N_3937,N_3189);
nor U4700 (N_4700,N_3212,N_3763);
xor U4701 (N_4701,N_3523,N_3931);
or U4702 (N_4702,N_3225,N_3973);
and U4703 (N_4703,N_3719,N_3484);
nor U4704 (N_4704,N_3742,N_3504);
or U4705 (N_4705,N_3480,N_3198);
and U4706 (N_4706,N_3639,N_3756);
or U4707 (N_4707,N_3262,N_3102);
nor U4708 (N_4708,N_3010,N_3031);
nand U4709 (N_4709,N_3672,N_3465);
nor U4710 (N_4710,N_3365,N_3868);
or U4711 (N_4711,N_3106,N_3168);
nand U4712 (N_4712,N_3939,N_3358);
xor U4713 (N_4713,N_3574,N_3716);
or U4714 (N_4714,N_3268,N_3590);
xor U4715 (N_4715,N_3059,N_3927);
or U4716 (N_4716,N_3983,N_3163);
nor U4717 (N_4717,N_3549,N_3581);
nor U4718 (N_4718,N_3786,N_3101);
nor U4719 (N_4719,N_3793,N_3086);
nor U4720 (N_4720,N_3557,N_3436);
or U4721 (N_4721,N_3027,N_3689);
nand U4722 (N_4722,N_3356,N_3476);
or U4723 (N_4723,N_3319,N_3440);
nor U4724 (N_4724,N_3025,N_3850);
nor U4725 (N_4725,N_3378,N_3102);
xor U4726 (N_4726,N_3617,N_3972);
nand U4727 (N_4727,N_3153,N_3955);
and U4728 (N_4728,N_3519,N_3647);
nand U4729 (N_4729,N_3002,N_3835);
and U4730 (N_4730,N_3065,N_3913);
and U4731 (N_4731,N_3860,N_3159);
nand U4732 (N_4732,N_3172,N_3098);
and U4733 (N_4733,N_3958,N_3950);
or U4734 (N_4734,N_3172,N_3650);
xnor U4735 (N_4735,N_3409,N_3305);
and U4736 (N_4736,N_3249,N_3912);
or U4737 (N_4737,N_3732,N_3448);
and U4738 (N_4738,N_3483,N_3080);
nand U4739 (N_4739,N_3738,N_3318);
nor U4740 (N_4740,N_3733,N_3310);
nand U4741 (N_4741,N_3936,N_3953);
or U4742 (N_4742,N_3237,N_3597);
nand U4743 (N_4743,N_3388,N_3026);
or U4744 (N_4744,N_3816,N_3307);
and U4745 (N_4745,N_3783,N_3229);
nand U4746 (N_4746,N_3254,N_3925);
nor U4747 (N_4747,N_3614,N_3793);
nor U4748 (N_4748,N_3336,N_3099);
and U4749 (N_4749,N_3786,N_3580);
nand U4750 (N_4750,N_3957,N_3326);
nand U4751 (N_4751,N_3522,N_3519);
nor U4752 (N_4752,N_3944,N_3885);
nor U4753 (N_4753,N_3625,N_3217);
nand U4754 (N_4754,N_3229,N_3540);
xor U4755 (N_4755,N_3191,N_3394);
or U4756 (N_4756,N_3271,N_3440);
xor U4757 (N_4757,N_3565,N_3767);
nand U4758 (N_4758,N_3395,N_3022);
nor U4759 (N_4759,N_3330,N_3490);
or U4760 (N_4760,N_3039,N_3305);
or U4761 (N_4761,N_3490,N_3449);
nand U4762 (N_4762,N_3052,N_3709);
nand U4763 (N_4763,N_3931,N_3716);
and U4764 (N_4764,N_3198,N_3608);
or U4765 (N_4765,N_3198,N_3308);
nor U4766 (N_4766,N_3662,N_3792);
and U4767 (N_4767,N_3797,N_3681);
nand U4768 (N_4768,N_3111,N_3682);
and U4769 (N_4769,N_3050,N_3658);
or U4770 (N_4770,N_3640,N_3110);
nand U4771 (N_4771,N_3648,N_3841);
xnor U4772 (N_4772,N_3119,N_3714);
xnor U4773 (N_4773,N_3464,N_3792);
or U4774 (N_4774,N_3156,N_3264);
or U4775 (N_4775,N_3845,N_3658);
or U4776 (N_4776,N_3185,N_3448);
and U4777 (N_4777,N_3058,N_3832);
nand U4778 (N_4778,N_3502,N_3348);
or U4779 (N_4779,N_3404,N_3823);
nor U4780 (N_4780,N_3768,N_3663);
xor U4781 (N_4781,N_3325,N_3351);
nor U4782 (N_4782,N_3045,N_3217);
nor U4783 (N_4783,N_3131,N_3641);
or U4784 (N_4784,N_3758,N_3536);
nand U4785 (N_4785,N_3345,N_3933);
nor U4786 (N_4786,N_3522,N_3042);
and U4787 (N_4787,N_3446,N_3089);
or U4788 (N_4788,N_3832,N_3461);
nor U4789 (N_4789,N_3357,N_3346);
and U4790 (N_4790,N_3057,N_3093);
or U4791 (N_4791,N_3451,N_3946);
or U4792 (N_4792,N_3730,N_3951);
and U4793 (N_4793,N_3366,N_3792);
xor U4794 (N_4794,N_3408,N_3495);
and U4795 (N_4795,N_3232,N_3098);
or U4796 (N_4796,N_3781,N_3542);
nand U4797 (N_4797,N_3427,N_3020);
xor U4798 (N_4798,N_3914,N_3322);
or U4799 (N_4799,N_3775,N_3793);
or U4800 (N_4800,N_3638,N_3031);
xor U4801 (N_4801,N_3481,N_3812);
nor U4802 (N_4802,N_3501,N_3772);
nor U4803 (N_4803,N_3281,N_3575);
nand U4804 (N_4804,N_3972,N_3740);
nand U4805 (N_4805,N_3931,N_3643);
nand U4806 (N_4806,N_3824,N_3672);
or U4807 (N_4807,N_3893,N_3590);
nand U4808 (N_4808,N_3227,N_3925);
or U4809 (N_4809,N_3418,N_3261);
nor U4810 (N_4810,N_3976,N_3637);
or U4811 (N_4811,N_3474,N_3882);
xnor U4812 (N_4812,N_3113,N_3358);
or U4813 (N_4813,N_3704,N_3583);
and U4814 (N_4814,N_3912,N_3418);
and U4815 (N_4815,N_3124,N_3650);
xnor U4816 (N_4816,N_3862,N_3954);
and U4817 (N_4817,N_3777,N_3979);
and U4818 (N_4818,N_3907,N_3274);
and U4819 (N_4819,N_3149,N_3732);
and U4820 (N_4820,N_3102,N_3834);
nor U4821 (N_4821,N_3511,N_3293);
nand U4822 (N_4822,N_3144,N_3970);
nor U4823 (N_4823,N_3932,N_3646);
nand U4824 (N_4824,N_3772,N_3176);
nor U4825 (N_4825,N_3713,N_3248);
nand U4826 (N_4826,N_3095,N_3764);
and U4827 (N_4827,N_3712,N_3430);
nor U4828 (N_4828,N_3371,N_3249);
and U4829 (N_4829,N_3869,N_3382);
and U4830 (N_4830,N_3543,N_3511);
nor U4831 (N_4831,N_3913,N_3301);
or U4832 (N_4832,N_3969,N_3502);
nand U4833 (N_4833,N_3179,N_3704);
or U4834 (N_4834,N_3530,N_3165);
or U4835 (N_4835,N_3752,N_3538);
and U4836 (N_4836,N_3629,N_3058);
and U4837 (N_4837,N_3691,N_3877);
or U4838 (N_4838,N_3809,N_3022);
nor U4839 (N_4839,N_3711,N_3966);
nand U4840 (N_4840,N_3814,N_3963);
and U4841 (N_4841,N_3379,N_3943);
xnor U4842 (N_4842,N_3031,N_3517);
xnor U4843 (N_4843,N_3303,N_3804);
xnor U4844 (N_4844,N_3750,N_3269);
nor U4845 (N_4845,N_3004,N_3433);
and U4846 (N_4846,N_3851,N_3289);
and U4847 (N_4847,N_3993,N_3670);
nor U4848 (N_4848,N_3801,N_3493);
nor U4849 (N_4849,N_3395,N_3585);
nand U4850 (N_4850,N_3776,N_3813);
xor U4851 (N_4851,N_3882,N_3174);
nor U4852 (N_4852,N_3920,N_3430);
xor U4853 (N_4853,N_3003,N_3271);
and U4854 (N_4854,N_3228,N_3189);
nand U4855 (N_4855,N_3285,N_3183);
or U4856 (N_4856,N_3628,N_3676);
and U4857 (N_4857,N_3319,N_3124);
and U4858 (N_4858,N_3085,N_3891);
and U4859 (N_4859,N_3755,N_3999);
and U4860 (N_4860,N_3415,N_3033);
nand U4861 (N_4861,N_3311,N_3046);
or U4862 (N_4862,N_3088,N_3358);
or U4863 (N_4863,N_3388,N_3614);
nor U4864 (N_4864,N_3686,N_3103);
or U4865 (N_4865,N_3782,N_3460);
or U4866 (N_4866,N_3963,N_3039);
nand U4867 (N_4867,N_3702,N_3556);
or U4868 (N_4868,N_3548,N_3109);
xor U4869 (N_4869,N_3679,N_3464);
xnor U4870 (N_4870,N_3877,N_3694);
xor U4871 (N_4871,N_3949,N_3606);
or U4872 (N_4872,N_3608,N_3689);
xor U4873 (N_4873,N_3331,N_3688);
and U4874 (N_4874,N_3182,N_3877);
and U4875 (N_4875,N_3451,N_3603);
nand U4876 (N_4876,N_3430,N_3612);
nor U4877 (N_4877,N_3877,N_3046);
nor U4878 (N_4878,N_3992,N_3279);
nand U4879 (N_4879,N_3588,N_3733);
and U4880 (N_4880,N_3999,N_3294);
nand U4881 (N_4881,N_3523,N_3055);
nand U4882 (N_4882,N_3673,N_3644);
nor U4883 (N_4883,N_3908,N_3474);
nor U4884 (N_4884,N_3530,N_3316);
nand U4885 (N_4885,N_3074,N_3804);
nor U4886 (N_4886,N_3615,N_3885);
nand U4887 (N_4887,N_3838,N_3871);
xnor U4888 (N_4888,N_3065,N_3565);
nor U4889 (N_4889,N_3634,N_3620);
and U4890 (N_4890,N_3944,N_3287);
nand U4891 (N_4891,N_3245,N_3940);
and U4892 (N_4892,N_3997,N_3626);
or U4893 (N_4893,N_3643,N_3604);
nand U4894 (N_4894,N_3599,N_3443);
nand U4895 (N_4895,N_3398,N_3058);
or U4896 (N_4896,N_3776,N_3929);
nand U4897 (N_4897,N_3899,N_3644);
nor U4898 (N_4898,N_3508,N_3162);
or U4899 (N_4899,N_3759,N_3213);
and U4900 (N_4900,N_3492,N_3831);
nor U4901 (N_4901,N_3661,N_3176);
nor U4902 (N_4902,N_3113,N_3706);
or U4903 (N_4903,N_3048,N_3461);
nand U4904 (N_4904,N_3209,N_3687);
and U4905 (N_4905,N_3005,N_3895);
or U4906 (N_4906,N_3511,N_3281);
nor U4907 (N_4907,N_3383,N_3268);
nor U4908 (N_4908,N_3193,N_3565);
or U4909 (N_4909,N_3066,N_3490);
and U4910 (N_4910,N_3153,N_3510);
nand U4911 (N_4911,N_3126,N_3493);
nand U4912 (N_4912,N_3590,N_3742);
nor U4913 (N_4913,N_3466,N_3450);
and U4914 (N_4914,N_3867,N_3350);
and U4915 (N_4915,N_3144,N_3630);
nor U4916 (N_4916,N_3486,N_3407);
or U4917 (N_4917,N_3042,N_3985);
xnor U4918 (N_4918,N_3110,N_3604);
xnor U4919 (N_4919,N_3170,N_3455);
nand U4920 (N_4920,N_3538,N_3202);
and U4921 (N_4921,N_3798,N_3541);
or U4922 (N_4922,N_3108,N_3500);
xor U4923 (N_4923,N_3131,N_3062);
nor U4924 (N_4924,N_3731,N_3073);
nand U4925 (N_4925,N_3100,N_3287);
and U4926 (N_4926,N_3968,N_3492);
nand U4927 (N_4927,N_3873,N_3573);
or U4928 (N_4928,N_3563,N_3721);
or U4929 (N_4929,N_3375,N_3008);
and U4930 (N_4930,N_3568,N_3989);
and U4931 (N_4931,N_3524,N_3908);
and U4932 (N_4932,N_3257,N_3940);
nor U4933 (N_4933,N_3850,N_3706);
or U4934 (N_4934,N_3243,N_3225);
and U4935 (N_4935,N_3846,N_3009);
or U4936 (N_4936,N_3242,N_3344);
nand U4937 (N_4937,N_3639,N_3382);
nand U4938 (N_4938,N_3536,N_3683);
and U4939 (N_4939,N_3373,N_3516);
nor U4940 (N_4940,N_3241,N_3824);
or U4941 (N_4941,N_3870,N_3814);
and U4942 (N_4942,N_3634,N_3793);
xnor U4943 (N_4943,N_3735,N_3812);
or U4944 (N_4944,N_3776,N_3114);
and U4945 (N_4945,N_3874,N_3740);
and U4946 (N_4946,N_3273,N_3231);
xor U4947 (N_4947,N_3944,N_3852);
or U4948 (N_4948,N_3816,N_3355);
nor U4949 (N_4949,N_3837,N_3696);
nor U4950 (N_4950,N_3247,N_3676);
nand U4951 (N_4951,N_3861,N_3700);
xor U4952 (N_4952,N_3800,N_3416);
xor U4953 (N_4953,N_3300,N_3533);
and U4954 (N_4954,N_3029,N_3540);
or U4955 (N_4955,N_3500,N_3469);
or U4956 (N_4956,N_3646,N_3204);
nor U4957 (N_4957,N_3725,N_3675);
and U4958 (N_4958,N_3964,N_3928);
nor U4959 (N_4959,N_3272,N_3726);
nand U4960 (N_4960,N_3247,N_3109);
and U4961 (N_4961,N_3636,N_3477);
and U4962 (N_4962,N_3111,N_3800);
nor U4963 (N_4963,N_3965,N_3239);
nand U4964 (N_4964,N_3700,N_3073);
nor U4965 (N_4965,N_3825,N_3423);
and U4966 (N_4966,N_3323,N_3988);
or U4967 (N_4967,N_3183,N_3794);
nand U4968 (N_4968,N_3930,N_3325);
or U4969 (N_4969,N_3526,N_3970);
or U4970 (N_4970,N_3325,N_3916);
and U4971 (N_4971,N_3424,N_3637);
nand U4972 (N_4972,N_3096,N_3423);
or U4973 (N_4973,N_3535,N_3733);
nand U4974 (N_4974,N_3106,N_3467);
or U4975 (N_4975,N_3881,N_3616);
nand U4976 (N_4976,N_3640,N_3311);
nor U4977 (N_4977,N_3182,N_3255);
nand U4978 (N_4978,N_3495,N_3388);
or U4979 (N_4979,N_3430,N_3563);
nand U4980 (N_4980,N_3449,N_3678);
or U4981 (N_4981,N_3184,N_3109);
nor U4982 (N_4982,N_3963,N_3241);
nand U4983 (N_4983,N_3789,N_3604);
or U4984 (N_4984,N_3803,N_3625);
and U4985 (N_4985,N_3095,N_3847);
xor U4986 (N_4986,N_3591,N_3510);
nor U4987 (N_4987,N_3500,N_3486);
nand U4988 (N_4988,N_3131,N_3530);
nor U4989 (N_4989,N_3582,N_3281);
or U4990 (N_4990,N_3868,N_3945);
nor U4991 (N_4991,N_3184,N_3801);
and U4992 (N_4992,N_3729,N_3423);
and U4993 (N_4993,N_3868,N_3809);
nor U4994 (N_4994,N_3025,N_3423);
and U4995 (N_4995,N_3451,N_3857);
nand U4996 (N_4996,N_3708,N_3060);
nor U4997 (N_4997,N_3342,N_3356);
and U4998 (N_4998,N_3547,N_3175);
and U4999 (N_4999,N_3116,N_3438);
or U5000 (N_5000,N_4358,N_4264);
and U5001 (N_5001,N_4217,N_4610);
nor U5002 (N_5002,N_4129,N_4307);
nand U5003 (N_5003,N_4112,N_4750);
nor U5004 (N_5004,N_4919,N_4484);
nand U5005 (N_5005,N_4970,N_4493);
nor U5006 (N_5006,N_4131,N_4442);
nor U5007 (N_5007,N_4446,N_4203);
and U5008 (N_5008,N_4943,N_4086);
xnor U5009 (N_5009,N_4069,N_4398);
nor U5010 (N_5010,N_4714,N_4092);
nor U5011 (N_5011,N_4257,N_4087);
nor U5012 (N_5012,N_4882,N_4439);
nand U5013 (N_5013,N_4539,N_4713);
and U5014 (N_5014,N_4804,N_4921);
xnor U5015 (N_5015,N_4572,N_4565);
or U5016 (N_5016,N_4595,N_4085);
xor U5017 (N_5017,N_4428,N_4334);
or U5018 (N_5018,N_4298,N_4959);
and U5019 (N_5019,N_4695,N_4044);
nor U5020 (N_5020,N_4424,N_4095);
or U5021 (N_5021,N_4792,N_4930);
nor U5022 (N_5022,N_4228,N_4248);
nand U5023 (N_5023,N_4956,N_4599);
nand U5024 (N_5024,N_4200,N_4250);
nor U5025 (N_5025,N_4474,N_4642);
xor U5026 (N_5026,N_4392,N_4693);
and U5027 (N_5027,N_4444,N_4522);
or U5028 (N_5028,N_4765,N_4616);
nor U5029 (N_5029,N_4404,N_4806);
and U5030 (N_5030,N_4329,N_4586);
nor U5031 (N_5031,N_4362,N_4831);
nand U5032 (N_5032,N_4518,N_4353);
and U5033 (N_5033,N_4467,N_4053);
nand U5034 (N_5034,N_4012,N_4189);
nor U5035 (N_5035,N_4662,N_4598);
nor U5036 (N_5036,N_4281,N_4304);
nor U5037 (N_5037,N_4426,N_4858);
nand U5038 (N_5038,N_4555,N_4551);
or U5039 (N_5039,N_4976,N_4238);
or U5040 (N_5040,N_4715,N_4547);
nand U5041 (N_5041,N_4732,N_4822);
and U5042 (N_5042,N_4960,N_4164);
or U5043 (N_5043,N_4074,N_4508);
xnor U5044 (N_5044,N_4784,N_4854);
or U5045 (N_5045,N_4267,N_4370);
and U5046 (N_5046,N_4051,N_4411);
or U5047 (N_5047,N_4675,N_4656);
nor U5048 (N_5048,N_4450,N_4585);
nor U5049 (N_5049,N_4157,N_4350);
or U5050 (N_5050,N_4670,N_4782);
and U5051 (N_5051,N_4139,N_4581);
and U5052 (N_5052,N_4277,N_4316);
nor U5053 (N_5053,N_4048,N_4192);
nand U5054 (N_5054,N_4883,N_4206);
and U5055 (N_5055,N_4688,N_4376);
and U5056 (N_5056,N_4721,N_4745);
nor U5057 (N_5057,N_4159,N_4753);
nor U5058 (N_5058,N_4512,N_4730);
nor U5059 (N_5059,N_4691,N_4867);
nand U5060 (N_5060,N_4541,N_4634);
nand U5061 (N_5061,N_4643,N_4673);
nor U5062 (N_5062,N_4696,N_4503);
nand U5063 (N_5063,N_4078,N_4229);
nor U5064 (N_5064,N_4099,N_4807);
nor U5065 (N_5065,N_4319,N_4749);
xnor U5066 (N_5066,N_4593,N_4031);
nor U5067 (N_5067,N_4817,N_4607);
nand U5068 (N_5068,N_4234,N_4460);
or U5069 (N_5069,N_4184,N_4116);
or U5070 (N_5070,N_4191,N_4396);
xnor U5071 (N_5071,N_4660,N_4577);
and U5072 (N_5072,N_4063,N_4866);
nand U5073 (N_5073,N_4395,N_4770);
or U5074 (N_5074,N_4725,N_4355);
xnor U5075 (N_5075,N_4456,N_4107);
and U5076 (N_5076,N_4140,N_4669);
or U5077 (N_5077,N_4712,N_4755);
and U5078 (N_5078,N_4818,N_4222);
or U5079 (N_5079,N_4330,N_4364);
nand U5080 (N_5080,N_4174,N_4747);
nor U5081 (N_5081,N_4357,N_4757);
nand U5082 (N_5082,N_4751,N_4678);
nor U5083 (N_5083,N_4361,N_4744);
and U5084 (N_5084,N_4470,N_4220);
and U5085 (N_5085,N_4346,N_4325);
and U5086 (N_5086,N_4072,N_4386);
and U5087 (N_5087,N_4705,N_4954);
nand U5088 (N_5088,N_4387,N_4080);
nand U5089 (N_5089,N_4038,N_4615);
or U5090 (N_5090,N_4957,N_4285);
nor U5091 (N_5091,N_4556,N_4423);
and U5092 (N_5092,N_4440,N_4499);
xor U5093 (N_5093,N_4618,N_4797);
or U5094 (N_5094,N_4024,N_4368);
nand U5095 (N_5095,N_4594,N_4901);
nor U5096 (N_5096,N_4632,N_4352);
nand U5097 (N_5097,N_4686,N_4596);
or U5098 (N_5098,N_4903,N_4528);
nor U5099 (N_5099,N_4195,N_4557);
nor U5100 (N_5100,N_4791,N_4653);
nand U5101 (N_5101,N_4698,N_4559);
xor U5102 (N_5102,N_4090,N_4886);
or U5103 (N_5103,N_4451,N_4253);
and U5104 (N_5104,N_4526,N_4150);
and U5105 (N_5105,N_4046,N_4065);
and U5106 (N_5106,N_4758,N_4597);
or U5107 (N_5107,N_4432,N_4168);
nand U5108 (N_5108,N_4059,N_4991);
or U5109 (N_5109,N_4079,N_4412);
xnor U5110 (N_5110,N_4067,N_4216);
or U5111 (N_5111,N_4198,N_4629);
or U5112 (N_5112,N_4852,N_4627);
and U5113 (N_5113,N_4938,N_4701);
nand U5114 (N_5114,N_4233,N_4500);
nand U5115 (N_5115,N_4413,N_4517);
nand U5116 (N_5116,N_4839,N_4975);
nor U5117 (N_5117,N_4231,N_4472);
nor U5118 (N_5118,N_4625,N_4734);
xor U5119 (N_5119,N_4360,N_4834);
nor U5120 (N_5120,N_4796,N_4431);
nand U5121 (N_5121,N_4601,N_4374);
and U5122 (N_5122,N_4082,N_4741);
and U5123 (N_5123,N_4527,N_4225);
nor U5124 (N_5124,N_4617,N_4057);
nor U5125 (N_5125,N_4863,N_4535);
nand U5126 (N_5126,N_4433,N_4710);
and U5127 (N_5127,N_4936,N_4182);
nor U5128 (N_5128,N_4335,N_4505);
nor U5129 (N_5129,N_4926,N_4153);
nor U5130 (N_5130,N_4382,N_4322);
nand U5131 (N_5131,N_4853,N_4469);
xnor U5132 (N_5132,N_4702,N_4015);
and U5133 (N_5133,N_4731,N_4454);
xor U5134 (N_5134,N_4911,N_4354);
xnor U5135 (N_5135,N_4972,N_4378);
nor U5136 (N_5136,N_4384,N_4449);
nor U5137 (N_5137,N_4981,N_4084);
nand U5138 (N_5138,N_4158,N_4996);
nor U5139 (N_5139,N_4125,N_4888);
nor U5140 (N_5140,N_4850,N_4210);
nor U5141 (N_5141,N_4733,N_4156);
nor U5142 (N_5142,N_4317,N_4754);
nor U5143 (N_5143,N_4992,N_4590);
xor U5144 (N_5144,N_4789,N_4054);
or U5145 (N_5145,N_4121,N_4922);
and U5146 (N_5146,N_4300,N_4416);
nand U5147 (N_5147,N_4978,N_4312);
nor U5148 (N_5148,N_4485,N_4194);
nand U5149 (N_5149,N_4504,N_4788);
xor U5150 (N_5150,N_4891,N_4737);
nor U5151 (N_5151,N_4743,N_4836);
nand U5152 (N_5152,N_4717,N_4331);
and U5153 (N_5153,N_4471,N_4811);
or U5154 (N_5154,N_4968,N_4644);
nor U5155 (N_5155,N_4964,N_4582);
or U5156 (N_5156,N_4016,N_4561);
nand U5157 (N_5157,N_4434,N_4639);
nand U5158 (N_5158,N_4939,N_4826);
nor U5159 (N_5159,N_4224,N_4829);
and U5160 (N_5160,N_4980,N_4127);
nand U5161 (N_5161,N_4342,N_4984);
or U5162 (N_5162,N_4814,N_4910);
nor U5163 (N_5163,N_4906,N_4628);
xor U5164 (N_5164,N_4830,N_4306);
or U5165 (N_5165,N_4613,N_4196);
and U5166 (N_5166,N_4260,N_4923);
nor U5167 (N_5167,N_4949,N_4025);
nand U5168 (N_5168,N_4998,N_4483);
or U5169 (N_5169,N_4815,N_4240);
or U5170 (N_5170,N_4133,N_4008);
xnor U5171 (N_5171,N_4833,N_4385);
or U5172 (N_5172,N_4985,N_4648);
and U5173 (N_5173,N_4963,N_4403);
xor U5174 (N_5174,N_4269,N_4847);
nand U5175 (N_5175,N_4511,N_4542);
nand U5176 (N_5176,N_4671,N_4429);
nor U5177 (N_5177,N_4066,N_4775);
nand U5178 (N_5178,N_4869,N_4408);
and U5179 (N_5179,N_4529,N_4945);
and U5180 (N_5180,N_4383,N_4783);
nand U5181 (N_5181,N_4029,N_4138);
nand U5182 (N_5182,N_4032,N_4679);
or U5183 (N_5183,N_4047,N_4146);
nor U5184 (N_5184,N_4772,N_4562);
nand U5185 (N_5185,N_4167,N_4605);
and U5186 (N_5186,N_4611,N_4962);
and U5187 (N_5187,N_4875,N_4974);
or U5188 (N_5188,N_4563,N_4844);
and U5189 (N_5189,N_4893,N_4247);
xnor U5190 (N_5190,N_4645,N_4707);
nand U5191 (N_5191,N_4659,N_4263);
or U5192 (N_5192,N_4668,N_4553);
and U5193 (N_5193,N_4213,N_4909);
xnor U5194 (N_5194,N_4672,N_4418);
or U5195 (N_5195,N_4952,N_4487);
and U5196 (N_5196,N_4083,N_4543);
nand U5197 (N_5197,N_4738,N_4437);
or U5198 (N_5198,N_4160,N_4583);
or U5199 (N_5199,N_4872,N_4941);
nor U5200 (N_5200,N_4301,N_4144);
nand U5201 (N_5201,N_4638,N_4173);
xnor U5202 (N_5202,N_4389,N_4574);
xnor U5203 (N_5203,N_4005,N_4478);
nand U5204 (N_5204,N_4391,N_4916);
and U5205 (N_5205,N_4103,N_4899);
and U5206 (N_5206,N_4820,N_4546);
nand U5207 (N_5207,N_4489,N_4873);
nor U5208 (N_5208,N_4457,N_4291);
and U5209 (N_5209,N_4179,N_4030);
nor U5210 (N_5210,N_4027,N_4925);
nand U5211 (N_5211,N_4718,N_4380);
and U5212 (N_5212,N_4245,N_4060);
xnor U5213 (N_5213,N_4096,N_4988);
nor U5214 (N_5214,N_4236,N_4934);
nand U5215 (N_5215,N_4631,N_4884);
or U5216 (N_5216,N_4533,N_4294);
or U5217 (N_5217,N_4415,N_4636);
nand U5218 (N_5218,N_4207,N_4163);
xor U5219 (N_5219,N_4777,N_4664);
or U5220 (N_5220,N_4455,N_4262);
xnor U5221 (N_5221,N_4037,N_4573);
nor U5222 (N_5222,N_4172,N_4023);
nor U5223 (N_5223,N_4193,N_4892);
nand U5224 (N_5224,N_4482,N_4958);
nand U5225 (N_5225,N_4538,N_4468);
nor U5226 (N_5226,N_4406,N_4843);
or U5227 (N_5227,N_4340,N_4697);
nand U5228 (N_5228,N_4190,N_4343);
nand U5229 (N_5229,N_4977,N_4676);
nor U5230 (N_5230,N_4677,N_4278);
nand U5231 (N_5231,N_4303,N_4861);
and U5232 (N_5232,N_4902,N_4812);
or U5233 (N_5233,N_4381,N_4983);
nand U5234 (N_5234,N_4049,N_4286);
or U5235 (N_5235,N_4622,N_4232);
xor U5236 (N_5236,N_4685,N_4104);
nand U5237 (N_5237,N_4390,N_4274);
or U5238 (N_5238,N_4525,N_4452);
nor U5239 (N_5239,N_4524,N_4108);
or U5240 (N_5240,N_4859,N_4935);
xnor U5241 (N_5241,N_4756,N_4600);
nor U5242 (N_5242,N_4033,N_4953);
xnor U5243 (N_5243,N_4620,N_4397);
xnor U5244 (N_5244,N_4036,N_4742);
and U5245 (N_5245,N_4205,N_4020);
or U5246 (N_5246,N_4762,N_4532);
nor U5247 (N_5247,N_4993,N_4706);
nand U5248 (N_5248,N_4689,N_4273);
nand U5249 (N_5249,N_4359,N_4897);
nor U5250 (N_5250,N_4202,N_4145);
nand U5251 (N_5251,N_4841,N_4105);
xor U5252 (N_5252,N_4865,N_4453);
xor U5253 (N_5253,N_4568,N_4979);
nand U5254 (N_5254,N_4043,N_4739);
nor U5255 (N_5255,N_4045,N_4375);
and U5256 (N_5256,N_4223,N_4513);
nor U5257 (N_5257,N_4100,N_4802);
nor U5258 (N_5258,N_4351,N_4914);
xnor U5259 (N_5259,N_4709,N_4333);
and U5260 (N_5260,N_4327,N_4227);
nor U5261 (N_5261,N_4272,N_4409);
and U5262 (N_5262,N_4619,N_4124);
or U5263 (N_5263,N_4746,N_4279);
and U5264 (N_5264,N_4769,N_4781);
and U5265 (N_5265,N_4969,N_4204);
nand U5266 (N_5266,N_4723,N_4479);
and U5267 (N_5267,N_4441,N_4035);
nand U5268 (N_5268,N_4249,N_4509);
nand U5269 (N_5269,N_4091,N_4399);
nand U5270 (N_5270,N_4780,N_4515);
and U5271 (N_5271,N_4134,N_4908);
nand U5272 (N_5272,N_4896,N_4177);
and U5273 (N_5273,N_4799,N_4497);
xnor U5274 (N_5274,N_4401,N_4915);
or U5275 (N_5275,N_4890,N_4845);
xor U5276 (N_5276,N_4349,N_4661);
nand U5277 (N_5277,N_4176,N_4900);
nor U5278 (N_5278,N_4315,N_4481);
and U5279 (N_5279,N_4680,N_4186);
nor U5280 (N_5280,N_4209,N_4514);
and U5281 (N_5281,N_4477,N_4641);
nand U5282 (N_5282,N_4215,N_4603);
xor U5283 (N_5283,N_4328,N_4933);
nor U5284 (N_5284,N_4237,N_4268);
nand U5285 (N_5285,N_4001,N_4724);
or U5286 (N_5286,N_4123,N_4075);
or U5287 (N_5287,N_4010,N_4283);
nor U5288 (N_5288,N_4161,N_4466);
nor U5289 (N_5289,N_4438,N_4379);
and U5290 (N_5290,N_4647,N_4877);
and U5291 (N_5291,N_4218,N_4735);
nand U5292 (N_5292,N_4425,N_4323);
nand U5293 (N_5293,N_4009,N_4621);
and U5294 (N_5294,N_4071,N_4690);
and U5295 (N_5295,N_4039,N_4637);
nor U5296 (N_5296,N_4870,N_4510);
and U5297 (N_5297,N_4427,N_4885);
or U5298 (N_5298,N_4109,N_4447);
nand U5299 (N_5299,N_4868,N_4825);
nor U5300 (N_5300,N_4904,N_4280);
nand U5301 (N_5301,N_4295,N_4986);
or U5302 (N_5302,N_4394,N_4989);
nand U5303 (N_5303,N_4462,N_4779);
nand U5304 (N_5304,N_4289,N_4492);
and U5305 (N_5305,N_4609,N_4912);
or U5306 (N_5306,N_4494,N_4475);
or U5307 (N_5307,N_4549,N_4019);
nor U5308 (N_5308,N_4275,N_4097);
xor U5309 (N_5309,N_4951,N_4464);
or U5310 (N_5310,N_4309,N_4230);
or U5311 (N_5311,N_4995,N_4363);
and U5312 (N_5312,N_4488,N_4917);
xnor U5313 (N_5313,N_4171,N_4531);
nand U5314 (N_5314,N_4373,N_4014);
and U5315 (N_5315,N_4860,N_4928);
nand U5316 (N_5316,N_4252,N_4716);
or U5317 (N_5317,N_4658,N_4534);
or U5318 (N_5318,N_4258,N_4626);
or U5319 (N_5319,N_4417,N_4683);
nand U5320 (N_5320,N_4259,N_4496);
or U5321 (N_5321,N_4170,N_4271);
nand U5322 (N_5322,N_4835,N_4459);
and U5323 (N_5323,N_4569,N_4320);
and U5324 (N_5324,N_4838,N_4388);
nor U5325 (N_5325,N_4567,N_4366);
nor U5326 (N_5326,N_4365,N_4965);
nand U5327 (N_5327,N_4824,N_4864);
nor U5328 (N_5328,N_4026,N_4341);
nor U5329 (N_5329,N_4786,N_4821);
nor U5330 (N_5330,N_4666,N_4550);
or U5331 (N_5331,N_4495,N_4407);
nor U5332 (N_5332,N_4851,N_4808);
and U5333 (N_5333,N_4879,N_4136);
nor U5334 (N_5334,N_4110,N_4076);
nor U5335 (N_5335,N_4007,N_4266);
nor U5336 (N_5336,N_4219,N_4655);
nand U5337 (N_5337,N_4183,N_4652);
and U5338 (N_5338,N_4663,N_4188);
and U5339 (N_5339,N_4332,N_4458);
or U5340 (N_5340,N_4130,N_4937);
nor U5341 (N_5341,N_4768,N_4564);
and U5342 (N_5342,N_4840,N_4443);
nand U5343 (N_5343,N_4501,N_4421);
and U5344 (N_5344,N_4313,N_4299);
nand U5345 (N_5345,N_4135,N_4848);
and U5346 (N_5346,N_4665,N_4187);
nand U5347 (N_5347,N_4516,N_4519);
and U5348 (N_5348,N_4119,N_4088);
or U5349 (N_5349,N_4729,N_4305);
xor U5350 (N_5350,N_4552,N_4151);
or U5351 (N_5351,N_4239,N_4752);
nor U5352 (N_5352,N_4113,N_4790);
nand U5353 (N_5353,N_4197,N_4767);
xnor U5354 (N_5354,N_4034,N_4640);
and U5355 (N_5355,N_4290,N_4764);
nand U5356 (N_5356,N_4785,N_4711);
nor U5357 (N_5357,N_4115,N_4261);
nor U5358 (N_5358,N_4654,N_4803);
nand U5359 (N_5359,N_4165,N_4293);
nand U5360 (N_5360,N_4558,N_4208);
xnor U5361 (N_5361,N_4147,N_4420);
nor U5362 (N_5362,N_4308,N_4310);
xor U5363 (N_5363,N_4297,N_4226);
xor U5364 (N_5364,N_4128,N_4874);
nand U5365 (N_5365,N_4805,N_4827);
and U5366 (N_5366,N_4093,N_4011);
nor U5367 (N_5367,N_4338,N_4571);
and U5368 (N_5368,N_4946,N_4324);
nand U5369 (N_5369,N_4918,N_4548);
nor U5370 (N_5370,N_4898,N_4056);
xnor U5371 (N_5371,N_4727,N_4606);
or U5372 (N_5372,N_4740,N_4728);
or U5373 (N_5373,N_4070,N_4212);
or U5374 (N_5374,N_4521,N_4842);
nor U5375 (N_5375,N_4646,N_4265);
and U5376 (N_5376,N_4061,N_4448);
and U5377 (N_5377,N_4703,N_4422);
or U5378 (N_5378,N_4624,N_4498);
nor U5379 (N_5379,N_4651,N_4246);
nand U5380 (N_5380,N_4955,N_4181);
or U5381 (N_5381,N_4720,N_4878);
nand U5382 (N_5382,N_4924,N_4486);
and U5383 (N_5383,N_4773,N_4787);
nor U5384 (N_5384,N_4132,N_4169);
and U5385 (N_5385,N_4126,N_4318);
nand U5386 (N_5386,N_4339,N_4201);
nor U5387 (N_5387,N_4942,N_4270);
nor U5388 (N_5388,N_4377,N_4588);
nand U5389 (N_5389,N_4759,N_4166);
and U5390 (N_5390,N_4578,N_4345);
or U5391 (N_5391,N_4846,N_4288);
xnor U5392 (N_5392,N_4856,N_4887);
nor U5393 (N_5393,N_4292,N_4947);
or U5394 (N_5394,N_4681,N_4667);
and U5395 (N_5395,N_4570,N_4592);
nor U5396 (N_5396,N_4871,N_4410);
or U5397 (N_5397,N_4967,N_4591);
and U5398 (N_5398,N_4684,N_4491);
and U5399 (N_5399,N_4221,N_4154);
nand U5400 (N_5400,N_4623,N_4372);
nor U5401 (N_5401,N_4137,N_4336);
nor U5402 (N_5402,N_4004,N_4021);
and U5403 (N_5403,N_4502,N_4296);
nand U5404 (N_5404,N_4114,N_4920);
nor U5405 (N_5405,N_4931,N_4576);
or U5406 (N_5406,N_4089,N_4687);
nor U5407 (N_5407,N_4180,N_4929);
nand U5408 (N_5408,N_4302,N_4774);
or U5409 (N_5409,N_4763,N_4604);
or U5410 (N_5410,N_4994,N_4143);
xor U5411 (N_5411,N_4445,N_4402);
or U5412 (N_5412,N_4722,N_4905);
nand U5413 (N_5413,N_4073,N_4400);
and U5414 (N_5414,N_4895,N_4950);
nor U5415 (N_5415,N_4614,N_4987);
nand U5416 (N_5416,N_4055,N_4540);
xnor U5417 (N_5417,N_4162,N_4098);
nor U5418 (N_5418,N_4507,N_4017);
nor U5419 (N_5419,N_4344,N_4175);
nand U5420 (N_5420,N_4211,N_4013);
nor U5421 (N_5421,N_4436,N_4694);
nor U5422 (N_5422,N_4256,N_4042);
or U5423 (N_5423,N_4849,N_4241);
and U5424 (N_5424,N_4894,N_4966);
nand U5425 (N_5425,N_4708,N_4214);
nor U5426 (N_5426,N_4000,N_4028);
and U5427 (N_5427,N_4798,N_4760);
nor U5428 (N_5428,N_4430,N_4052);
xnor U5429 (N_5429,N_4794,N_4480);
xnor U5430 (N_5430,N_4094,N_4371);
and U5431 (N_5431,N_4700,N_4699);
or U5432 (N_5432,N_4321,N_4649);
and U5433 (N_5433,N_4832,N_4287);
or U5434 (N_5434,N_4657,N_4337);
nor U5435 (N_5435,N_4748,N_4490);
nor U5436 (N_5436,N_4006,N_4635);
nor U5437 (N_5437,N_4149,N_4022);
and U5438 (N_5438,N_4465,N_4587);
or U5439 (N_5439,N_4579,N_4520);
nand U5440 (N_5440,N_4932,N_4122);
or U5441 (N_5441,N_4117,N_4771);
nor U5442 (N_5442,N_4463,N_4155);
or U5443 (N_5443,N_4536,N_4999);
nand U5444 (N_5444,N_4692,N_4178);
and U5445 (N_5445,N_4889,N_4199);
or U5446 (N_5446,N_4704,N_4414);
or U5447 (N_5447,N_4102,N_4816);
or U5448 (N_5448,N_4793,N_4506);
or U5449 (N_5449,N_4682,N_4837);
xnor U5450 (N_5450,N_4393,N_4726);
nand U5451 (N_5451,N_4356,N_4284);
and U5452 (N_5452,N_4800,N_4855);
nor U5453 (N_5453,N_4566,N_4064);
or U5454 (N_5454,N_4326,N_4120);
nor U5455 (N_5455,N_4584,N_4761);
nand U5456 (N_5456,N_4058,N_4880);
nand U5457 (N_5457,N_4602,N_4367);
xnor U5458 (N_5458,N_4118,N_4018);
nand U5459 (N_5459,N_4111,N_4244);
nor U5460 (N_5460,N_4255,N_4537);
nor U5461 (N_5461,N_4369,N_4142);
xnor U5462 (N_5462,N_4062,N_4476);
or U5463 (N_5463,N_4948,N_4242);
nor U5464 (N_5464,N_4990,N_4907);
nand U5465 (N_5465,N_4940,N_4348);
and U5466 (N_5466,N_4612,N_4560);
nor U5467 (N_5467,N_4152,N_4971);
nand U5468 (N_5468,N_4650,N_4674);
nor U5469 (N_5469,N_4311,N_4461);
and U5470 (N_5470,N_4068,N_4589);
or U5471 (N_5471,N_4003,N_4435);
or U5472 (N_5472,N_4795,N_4002);
nand U5473 (N_5473,N_4040,N_4554);
xor U5474 (N_5474,N_4801,N_4575);
xnor U5475 (N_5475,N_4185,N_4077);
nand U5476 (N_5476,N_4819,N_4251);
xnor U5477 (N_5477,N_4544,N_4141);
and U5478 (N_5478,N_4314,N_4881);
nand U5479 (N_5479,N_4828,N_4050);
or U5480 (N_5480,N_4608,N_4997);
or U5481 (N_5481,N_4927,N_4106);
nand U5482 (N_5482,N_4719,N_4347);
nand U5483 (N_5483,N_4913,N_4405);
nor U5484 (N_5484,N_4254,N_4736);
and U5485 (N_5485,N_4276,N_4810);
nor U5486 (N_5486,N_4813,N_4876);
nand U5487 (N_5487,N_4961,N_4419);
nor U5488 (N_5488,N_4766,N_4523);
xnor U5489 (N_5489,N_4823,N_4973);
xnor U5490 (N_5490,N_4630,N_4944);
xnor U5491 (N_5491,N_4776,N_4857);
and U5492 (N_5492,N_4778,N_4235);
and U5493 (N_5493,N_4148,N_4041);
nand U5494 (N_5494,N_4282,N_4809);
nand U5495 (N_5495,N_4862,N_4545);
xnor U5496 (N_5496,N_4081,N_4473);
or U5497 (N_5497,N_4101,N_4633);
nor U5498 (N_5498,N_4580,N_4243);
xnor U5499 (N_5499,N_4982,N_4530);
and U5500 (N_5500,N_4852,N_4790);
and U5501 (N_5501,N_4784,N_4873);
nand U5502 (N_5502,N_4066,N_4016);
nand U5503 (N_5503,N_4185,N_4412);
or U5504 (N_5504,N_4356,N_4906);
and U5505 (N_5505,N_4593,N_4475);
xor U5506 (N_5506,N_4295,N_4623);
nand U5507 (N_5507,N_4024,N_4659);
or U5508 (N_5508,N_4571,N_4787);
xor U5509 (N_5509,N_4469,N_4660);
nand U5510 (N_5510,N_4965,N_4275);
or U5511 (N_5511,N_4707,N_4070);
nor U5512 (N_5512,N_4221,N_4606);
or U5513 (N_5513,N_4467,N_4305);
or U5514 (N_5514,N_4771,N_4613);
nor U5515 (N_5515,N_4057,N_4442);
nand U5516 (N_5516,N_4265,N_4545);
nand U5517 (N_5517,N_4319,N_4690);
xnor U5518 (N_5518,N_4286,N_4894);
nor U5519 (N_5519,N_4659,N_4287);
and U5520 (N_5520,N_4384,N_4007);
nand U5521 (N_5521,N_4236,N_4032);
nand U5522 (N_5522,N_4976,N_4220);
or U5523 (N_5523,N_4822,N_4538);
and U5524 (N_5524,N_4462,N_4954);
xor U5525 (N_5525,N_4064,N_4173);
or U5526 (N_5526,N_4517,N_4167);
nand U5527 (N_5527,N_4136,N_4260);
or U5528 (N_5528,N_4159,N_4588);
and U5529 (N_5529,N_4196,N_4726);
nor U5530 (N_5530,N_4800,N_4213);
nand U5531 (N_5531,N_4949,N_4632);
xnor U5532 (N_5532,N_4143,N_4542);
or U5533 (N_5533,N_4669,N_4053);
nor U5534 (N_5534,N_4900,N_4583);
nor U5535 (N_5535,N_4794,N_4312);
and U5536 (N_5536,N_4234,N_4395);
and U5537 (N_5537,N_4018,N_4914);
xnor U5538 (N_5538,N_4332,N_4021);
nand U5539 (N_5539,N_4414,N_4169);
xor U5540 (N_5540,N_4155,N_4457);
or U5541 (N_5541,N_4723,N_4622);
or U5542 (N_5542,N_4521,N_4064);
xnor U5543 (N_5543,N_4828,N_4444);
nand U5544 (N_5544,N_4633,N_4755);
nand U5545 (N_5545,N_4841,N_4207);
nand U5546 (N_5546,N_4329,N_4821);
xnor U5547 (N_5547,N_4142,N_4062);
nand U5548 (N_5548,N_4693,N_4584);
and U5549 (N_5549,N_4836,N_4879);
nand U5550 (N_5550,N_4539,N_4654);
or U5551 (N_5551,N_4215,N_4138);
or U5552 (N_5552,N_4160,N_4030);
or U5553 (N_5553,N_4549,N_4061);
and U5554 (N_5554,N_4022,N_4232);
and U5555 (N_5555,N_4763,N_4370);
and U5556 (N_5556,N_4838,N_4853);
or U5557 (N_5557,N_4487,N_4686);
or U5558 (N_5558,N_4298,N_4019);
nand U5559 (N_5559,N_4052,N_4246);
nor U5560 (N_5560,N_4311,N_4621);
nand U5561 (N_5561,N_4713,N_4955);
and U5562 (N_5562,N_4023,N_4678);
or U5563 (N_5563,N_4450,N_4484);
nor U5564 (N_5564,N_4262,N_4239);
nor U5565 (N_5565,N_4544,N_4011);
or U5566 (N_5566,N_4457,N_4785);
and U5567 (N_5567,N_4659,N_4365);
nor U5568 (N_5568,N_4111,N_4382);
or U5569 (N_5569,N_4093,N_4242);
nor U5570 (N_5570,N_4580,N_4011);
nor U5571 (N_5571,N_4385,N_4005);
or U5572 (N_5572,N_4456,N_4211);
nand U5573 (N_5573,N_4296,N_4072);
nor U5574 (N_5574,N_4382,N_4352);
or U5575 (N_5575,N_4962,N_4181);
and U5576 (N_5576,N_4211,N_4657);
and U5577 (N_5577,N_4000,N_4198);
nand U5578 (N_5578,N_4466,N_4493);
nor U5579 (N_5579,N_4946,N_4081);
or U5580 (N_5580,N_4181,N_4840);
nand U5581 (N_5581,N_4166,N_4640);
nand U5582 (N_5582,N_4822,N_4764);
xor U5583 (N_5583,N_4718,N_4149);
nand U5584 (N_5584,N_4713,N_4186);
nor U5585 (N_5585,N_4594,N_4837);
nand U5586 (N_5586,N_4996,N_4550);
nand U5587 (N_5587,N_4208,N_4665);
nand U5588 (N_5588,N_4444,N_4042);
nand U5589 (N_5589,N_4618,N_4733);
xor U5590 (N_5590,N_4119,N_4154);
or U5591 (N_5591,N_4000,N_4784);
or U5592 (N_5592,N_4158,N_4942);
nor U5593 (N_5593,N_4091,N_4824);
nand U5594 (N_5594,N_4435,N_4737);
nand U5595 (N_5595,N_4429,N_4831);
nand U5596 (N_5596,N_4382,N_4279);
and U5597 (N_5597,N_4369,N_4513);
and U5598 (N_5598,N_4419,N_4991);
and U5599 (N_5599,N_4082,N_4715);
nor U5600 (N_5600,N_4086,N_4571);
and U5601 (N_5601,N_4565,N_4368);
and U5602 (N_5602,N_4709,N_4325);
and U5603 (N_5603,N_4822,N_4466);
xor U5604 (N_5604,N_4022,N_4874);
nand U5605 (N_5605,N_4951,N_4334);
nand U5606 (N_5606,N_4162,N_4602);
nand U5607 (N_5607,N_4344,N_4934);
and U5608 (N_5608,N_4430,N_4315);
nor U5609 (N_5609,N_4405,N_4963);
and U5610 (N_5610,N_4506,N_4940);
nor U5611 (N_5611,N_4223,N_4322);
and U5612 (N_5612,N_4457,N_4689);
and U5613 (N_5613,N_4058,N_4631);
nand U5614 (N_5614,N_4256,N_4828);
or U5615 (N_5615,N_4399,N_4610);
or U5616 (N_5616,N_4834,N_4087);
and U5617 (N_5617,N_4370,N_4772);
nor U5618 (N_5618,N_4104,N_4073);
or U5619 (N_5619,N_4458,N_4540);
nor U5620 (N_5620,N_4642,N_4366);
xor U5621 (N_5621,N_4937,N_4308);
nand U5622 (N_5622,N_4464,N_4317);
or U5623 (N_5623,N_4659,N_4997);
or U5624 (N_5624,N_4285,N_4283);
and U5625 (N_5625,N_4911,N_4478);
or U5626 (N_5626,N_4927,N_4034);
xnor U5627 (N_5627,N_4214,N_4438);
nand U5628 (N_5628,N_4069,N_4735);
nor U5629 (N_5629,N_4478,N_4031);
or U5630 (N_5630,N_4159,N_4120);
nand U5631 (N_5631,N_4966,N_4404);
or U5632 (N_5632,N_4421,N_4787);
nand U5633 (N_5633,N_4528,N_4682);
xor U5634 (N_5634,N_4484,N_4220);
and U5635 (N_5635,N_4260,N_4456);
nor U5636 (N_5636,N_4097,N_4875);
and U5637 (N_5637,N_4057,N_4546);
nand U5638 (N_5638,N_4203,N_4763);
or U5639 (N_5639,N_4182,N_4235);
nand U5640 (N_5640,N_4515,N_4574);
and U5641 (N_5641,N_4846,N_4956);
xnor U5642 (N_5642,N_4965,N_4825);
nand U5643 (N_5643,N_4089,N_4524);
or U5644 (N_5644,N_4264,N_4680);
nand U5645 (N_5645,N_4231,N_4331);
and U5646 (N_5646,N_4367,N_4057);
or U5647 (N_5647,N_4709,N_4312);
and U5648 (N_5648,N_4513,N_4145);
nand U5649 (N_5649,N_4919,N_4775);
and U5650 (N_5650,N_4285,N_4207);
nand U5651 (N_5651,N_4433,N_4735);
nor U5652 (N_5652,N_4882,N_4221);
nand U5653 (N_5653,N_4326,N_4141);
nand U5654 (N_5654,N_4506,N_4206);
nor U5655 (N_5655,N_4519,N_4065);
nand U5656 (N_5656,N_4124,N_4170);
and U5657 (N_5657,N_4016,N_4705);
or U5658 (N_5658,N_4072,N_4694);
nor U5659 (N_5659,N_4843,N_4148);
and U5660 (N_5660,N_4300,N_4304);
nor U5661 (N_5661,N_4884,N_4511);
nand U5662 (N_5662,N_4546,N_4618);
and U5663 (N_5663,N_4189,N_4030);
and U5664 (N_5664,N_4055,N_4563);
or U5665 (N_5665,N_4398,N_4980);
xor U5666 (N_5666,N_4959,N_4329);
nand U5667 (N_5667,N_4281,N_4399);
or U5668 (N_5668,N_4505,N_4769);
and U5669 (N_5669,N_4560,N_4861);
nor U5670 (N_5670,N_4713,N_4398);
or U5671 (N_5671,N_4113,N_4570);
or U5672 (N_5672,N_4592,N_4378);
nand U5673 (N_5673,N_4671,N_4157);
nor U5674 (N_5674,N_4786,N_4753);
nor U5675 (N_5675,N_4779,N_4658);
nor U5676 (N_5676,N_4497,N_4304);
nor U5677 (N_5677,N_4097,N_4198);
nor U5678 (N_5678,N_4462,N_4301);
nor U5679 (N_5679,N_4767,N_4910);
or U5680 (N_5680,N_4839,N_4722);
or U5681 (N_5681,N_4239,N_4337);
or U5682 (N_5682,N_4031,N_4365);
nor U5683 (N_5683,N_4135,N_4003);
nor U5684 (N_5684,N_4951,N_4911);
nand U5685 (N_5685,N_4150,N_4654);
or U5686 (N_5686,N_4617,N_4409);
nor U5687 (N_5687,N_4880,N_4016);
and U5688 (N_5688,N_4456,N_4182);
and U5689 (N_5689,N_4005,N_4938);
and U5690 (N_5690,N_4151,N_4557);
or U5691 (N_5691,N_4531,N_4705);
or U5692 (N_5692,N_4224,N_4792);
nand U5693 (N_5693,N_4232,N_4905);
or U5694 (N_5694,N_4438,N_4329);
xnor U5695 (N_5695,N_4010,N_4681);
and U5696 (N_5696,N_4218,N_4722);
and U5697 (N_5697,N_4789,N_4362);
nand U5698 (N_5698,N_4135,N_4590);
nand U5699 (N_5699,N_4693,N_4931);
or U5700 (N_5700,N_4546,N_4143);
nand U5701 (N_5701,N_4919,N_4754);
nand U5702 (N_5702,N_4871,N_4478);
and U5703 (N_5703,N_4938,N_4505);
xnor U5704 (N_5704,N_4234,N_4295);
xnor U5705 (N_5705,N_4351,N_4210);
and U5706 (N_5706,N_4841,N_4165);
nand U5707 (N_5707,N_4058,N_4783);
and U5708 (N_5708,N_4270,N_4305);
nand U5709 (N_5709,N_4374,N_4304);
nor U5710 (N_5710,N_4695,N_4016);
nor U5711 (N_5711,N_4276,N_4383);
and U5712 (N_5712,N_4387,N_4995);
nand U5713 (N_5713,N_4351,N_4137);
xnor U5714 (N_5714,N_4532,N_4621);
nor U5715 (N_5715,N_4252,N_4416);
xor U5716 (N_5716,N_4460,N_4778);
and U5717 (N_5717,N_4519,N_4085);
nor U5718 (N_5718,N_4778,N_4137);
nand U5719 (N_5719,N_4344,N_4076);
nand U5720 (N_5720,N_4198,N_4508);
or U5721 (N_5721,N_4103,N_4772);
or U5722 (N_5722,N_4886,N_4494);
nand U5723 (N_5723,N_4428,N_4120);
xnor U5724 (N_5724,N_4659,N_4982);
and U5725 (N_5725,N_4151,N_4636);
nor U5726 (N_5726,N_4167,N_4488);
nand U5727 (N_5727,N_4444,N_4846);
or U5728 (N_5728,N_4664,N_4546);
and U5729 (N_5729,N_4873,N_4943);
xnor U5730 (N_5730,N_4369,N_4702);
nand U5731 (N_5731,N_4588,N_4254);
and U5732 (N_5732,N_4050,N_4518);
nand U5733 (N_5733,N_4644,N_4893);
nand U5734 (N_5734,N_4581,N_4815);
nor U5735 (N_5735,N_4376,N_4617);
nor U5736 (N_5736,N_4505,N_4288);
nor U5737 (N_5737,N_4412,N_4439);
and U5738 (N_5738,N_4451,N_4401);
and U5739 (N_5739,N_4390,N_4588);
nand U5740 (N_5740,N_4195,N_4597);
nor U5741 (N_5741,N_4486,N_4414);
and U5742 (N_5742,N_4475,N_4089);
nand U5743 (N_5743,N_4382,N_4549);
xnor U5744 (N_5744,N_4325,N_4535);
and U5745 (N_5745,N_4364,N_4382);
xnor U5746 (N_5746,N_4847,N_4876);
nor U5747 (N_5747,N_4996,N_4272);
and U5748 (N_5748,N_4709,N_4370);
or U5749 (N_5749,N_4956,N_4176);
nor U5750 (N_5750,N_4062,N_4253);
and U5751 (N_5751,N_4098,N_4980);
and U5752 (N_5752,N_4960,N_4644);
and U5753 (N_5753,N_4758,N_4829);
nor U5754 (N_5754,N_4239,N_4585);
nand U5755 (N_5755,N_4347,N_4363);
nor U5756 (N_5756,N_4052,N_4065);
nor U5757 (N_5757,N_4025,N_4372);
nor U5758 (N_5758,N_4094,N_4038);
nand U5759 (N_5759,N_4624,N_4126);
nand U5760 (N_5760,N_4354,N_4431);
and U5761 (N_5761,N_4714,N_4479);
nor U5762 (N_5762,N_4978,N_4548);
and U5763 (N_5763,N_4744,N_4756);
xor U5764 (N_5764,N_4725,N_4490);
nand U5765 (N_5765,N_4610,N_4042);
or U5766 (N_5766,N_4230,N_4921);
and U5767 (N_5767,N_4654,N_4597);
and U5768 (N_5768,N_4067,N_4988);
nand U5769 (N_5769,N_4954,N_4987);
and U5770 (N_5770,N_4072,N_4470);
xnor U5771 (N_5771,N_4772,N_4110);
xor U5772 (N_5772,N_4339,N_4783);
xor U5773 (N_5773,N_4846,N_4826);
nor U5774 (N_5774,N_4931,N_4098);
nor U5775 (N_5775,N_4158,N_4152);
or U5776 (N_5776,N_4359,N_4125);
and U5777 (N_5777,N_4058,N_4285);
nor U5778 (N_5778,N_4563,N_4207);
and U5779 (N_5779,N_4205,N_4815);
or U5780 (N_5780,N_4870,N_4426);
or U5781 (N_5781,N_4668,N_4069);
xnor U5782 (N_5782,N_4455,N_4771);
and U5783 (N_5783,N_4029,N_4677);
nor U5784 (N_5784,N_4178,N_4440);
or U5785 (N_5785,N_4328,N_4785);
or U5786 (N_5786,N_4791,N_4926);
nor U5787 (N_5787,N_4556,N_4155);
nand U5788 (N_5788,N_4829,N_4916);
nand U5789 (N_5789,N_4880,N_4668);
nor U5790 (N_5790,N_4841,N_4335);
nor U5791 (N_5791,N_4289,N_4695);
and U5792 (N_5792,N_4286,N_4079);
or U5793 (N_5793,N_4150,N_4414);
or U5794 (N_5794,N_4380,N_4415);
nor U5795 (N_5795,N_4704,N_4808);
and U5796 (N_5796,N_4396,N_4898);
nor U5797 (N_5797,N_4737,N_4056);
and U5798 (N_5798,N_4288,N_4947);
nor U5799 (N_5799,N_4157,N_4563);
and U5800 (N_5800,N_4773,N_4102);
nand U5801 (N_5801,N_4777,N_4807);
xnor U5802 (N_5802,N_4319,N_4580);
or U5803 (N_5803,N_4985,N_4365);
xor U5804 (N_5804,N_4437,N_4715);
and U5805 (N_5805,N_4512,N_4999);
xor U5806 (N_5806,N_4840,N_4635);
or U5807 (N_5807,N_4882,N_4311);
and U5808 (N_5808,N_4776,N_4010);
and U5809 (N_5809,N_4930,N_4125);
and U5810 (N_5810,N_4417,N_4968);
and U5811 (N_5811,N_4272,N_4835);
xnor U5812 (N_5812,N_4689,N_4336);
and U5813 (N_5813,N_4117,N_4512);
nand U5814 (N_5814,N_4920,N_4359);
nand U5815 (N_5815,N_4023,N_4239);
nand U5816 (N_5816,N_4659,N_4908);
nor U5817 (N_5817,N_4791,N_4779);
nand U5818 (N_5818,N_4701,N_4384);
nand U5819 (N_5819,N_4296,N_4902);
and U5820 (N_5820,N_4565,N_4328);
nor U5821 (N_5821,N_4625,N_4148);
and U5822 (N_5822,N_4665,N_4150);
nand U5823 (N_5823,N_4073,N_4062);
nand U5824 (N_5824,N_4465,N_4820);
or U5825 (N_5825,N_4884,N_4693);
and U5826 (N_5826,N_4475,N_4839);
and U5827 (N_5827,N_4723,N_4291);
and U5828 (N_5828,N_4301,N_4000);
nor U5829 (N_5829,N_4102,N_4409);
and U5830 (N_5830,N_4294,N_4005);
xor U5831 (N_5831,N_4336,N_4221);
xnor U5832 (N_5832,N_4971,N_4806);
xor U5833 (N_5833,N_4218,N_4944);
or U5834 (N_5834,N_4631,N_4730);
nor U5835 (N_5835,N_4826,N_4444);
nor U5836 (N_5836,N_4414,N_4330);
and U5837 (N_5837,N_4537,N_4567);
nand U5838 (N_5838,N_4064,N_4981);
and U5839 (N_5839,N_4549,N_4053);
nor U5840 (N_5840,N_4830,N_4490);
nor U5841 (N_5841,N_4916,N_4768);
or U5842 (N_5842,N_4894,N_4382);
nor U5843 (N_5843,N_4120,N_4897);
xor U5844 (N_5844,N_4480,N_4051);
or U5845 (N_5845,N_4942,N_4576);
or U5846 (N_5846,N_4600,N_4382);
and U5847 (N_5847,N_4274,N_4560);
nor U5848 (N_5848,N_4724,N_4382);
nor U5849 (N_5849,N_4497,N_4258);
and U5850 (N_5850,N_4170,N_4636);
nor U5851 (N_5851,N_4785,N_4423);
xnor U5852 (N_5852,N_4916,N_4502);
nor U5853 (N_5853,N_4483,N_4269);
nand U5854 (N_5854,N_4786,N_4553);
and U5855 (N_5855,N_4269,N_4260);
and U5856 (N_5856,N_4568,N_4836);
nand U5857 (N_5857,N_4187,N_4584);
nor U5858 (N_5858,N_4857,N_4613);
nor U5859 (N_5859,N_4883,N_4001);
or U5860 (N_5860,N_4610,N_4977);
nor U5861 (N_5861,N_4766,N_4879);
nor U5862 (N_5862,N_4238,N_4871);
and U5863 (N_5863,N_4155,N_4351);
nand U5864 (N_5864,N_4616,N_4585);
nand U5865 (N_5865,N_4266,N_4320);
nor U5866 (N_5866,N_4674,N_4671);
nand U5867 (N_5867,N_4157,N_4072);
nand U5868 (N_5868,N_4503,N_4090);
and U5869 (N_5869,N_4658,N_4867);
or U5870 (N_5870,N_4378,N_4660);
or U5871 (N_5871,N_4195,N_4721);
and U5872 (N_5872,N_4590,N_4516);
nor U5873 (N_5873,N_4457,N_4262);
or U5874 (N_5874,N_4549,N_4579);
nor U5875 (N_5875,N_4424,N_4764);
xor U5876 (N_5876,N_4048,N_4885);
and U5877 (N_5877,N_4896,N_4856);
nor U5878 (N_5878,N_4350,N_4139);
xor U5879 (N_5879,N_4570,N_4100);
or U5880 (N_5880,N_4566,N_4445);
nor U5881 (N_5881,N_4254,N_4605);
or U5882 (N_5882,N_4262,N_4305);
nand U5883 (N_5883,N_4481,N_4748);
and U5884 (N_5884,N_4339,N_4999);
nor U5885 (N_5885,N_4734,N_4216);
or U5886 (N_5886,N_4010,N_4842);
or U5887 (N_5887,N_4246,N_4910);
or U5888 (N_5888,N_4253,N_4531);
nand U5889 (N_5889,N_4674,N_4619);
xor U5890 (N_5890,N_4824,N_4528);
nor U5891 (N_5891,N_4834,N_4254);
nor U5892 (N_5892,N_4041,N_4101);
nor U5893 (N_5893,N_4561,N_4683);
and U5894 (N_5894,N_4695,N_4129);
or U5895 (N_5895,N_4298,N_4767);
or U5896 (N_5896,N_4608,N_4896);
or U5897 (N_5897,N_4139,N_4160);
and U5898 (N_5898,N_4877,N_4759);
nand U5899 (N_5899,N_4662,N_4783);
nor U5900 (N_5900,N_4888,N_4599);
nor U5901 (N_5901,N_4045,N_4464);
nor U5902 (N_5902,N_4567,N_4130);
and U5903 (N_5903,N_4942,N_4274);
or U5904 (N_5904,N_4112,N_4733);
and U5905 (N_5905,N_4400,N_4933);
or U5906 (N_5906,N_4323,N_4868);
nor U5907 (N_5907,N_4329,N_4748);
or U5908 (N_5908,N_4365,N_4488);
xnor U5909 (N_5909,N_4356,N_4824);
and U5910 (N_5910,N_4787,N_4925);
or U5911 (N_5911,N_4270,N_4661);
and U5912 (N_5912,N_4383,N_4775);
nand U5913 (N_5913,N_4735,N_4206);
nor U5914 (N_5914,N_4147,N_4350);
nor U5915 (N_5915,N_4691,N_4626);
nor U5916 (N_5916,N_4127,N_4885);
or U5917 (N_5917,N_4264,N_4871);
nor U5918 (N_5918,N_4067,N_4704);
nor U5919 (N_5919,N_4767,N_4374);
and U5920 (N_5920,N_4622,N_4107);
or U5921 (N_5921,N_4897,N_4971);
nor U5922 (N_5922,N_4954,N_4049);
and U5923 (N_5923,N_4729,N_4713);
and U5924 (N_5924,N_4886,N_4470);
xnor U5925 (N_5925,N_4182,N_4564);
and U5926 (N_5926,N_4000,N_4304);
xor U5927 (N_5927,N_4937,N_4565);
and U5928 (N_5928,N_4047,N_4094);
nor U5929 (N_5929,N_4870,N_4247);
and U5930 (N_5930,N_4303,N_4565);
or U5931 (N_5931,N_4148,N_4225);
nor U5932 (N_5932,N_4383,N_4917);
xor U5933 (N_5933,N_4625,N_4438);
or U5934 (N_5934,N_4424,N_4079);
nand U5935 (N_5935,N_4636,N_4702);
nand U5936 (N_5936,N_4368,N_4749);
nor U5937 (N_5937,N_4801,N_4032);
or U5938 (N_5938,N_4584,N_4744);
nand U5939 (N_5939,N_4017,N_4966);
or U5940 (N_5940,N_4459,N_4749);
nor U5941 (N_5941,N_4593,N_4286);
nand U5942 (N_5942,N_4428,N_4088);
nand U5943 (N_5943,N_4367,N_4506);
or U5944 (N_5944,N_4370,N_4183);
xnor U5945 (N_5945,N_4354,N_4606);
nand U5946 (N_5946,N_4316,N_4052);
xor U5947 (N_5947,N_4174,N_4866);
or U5948 (N_5948,N_4306,N_4282);
or U5949 (N_5949,N_4288,N_4578);
or U5950 (N_5950,N_4832,N_4449);
nand U5951 (N_5951,N_4715,N_4817);
or U5952 (N_5952,N_4331,N_4422);
or U5953 (N_5953,N_4245,N_4608);
and U5954 (N_5954,N_4016,N_4105);
or U5955 (N_5955,N_4031,N_4169);
and U5956 (N_5956,N_4628,N_4495);
or U5957 (N_5957,N_4051,N_4436);
or U5958 (N_5958,N_4540,N_4617);
xor U5959 (N_5959,N_4461,N_4363);
and U5960 (N_5960,N_4438,N_4409);
nand U5961 (N_5961,N_4248,N_4826);
nor U5962 (N_5962,N_4912,N_4092);
and U5963 (N_5963,N_4378,N_4089);
nand U5964 (N_5964,N_4612,N_4723);
or U5965 (N_5965,N_4855,N_4411);
or U5966 (N_5966,N_4270,N_4166);
and U5967 (N_5967,N_4972,N_4412);
nor U5968 (N_5968,N_4774,N_4231);
and U5969 (N_5969,N_4040,N_4694);
xor U5970 (N_5970,N_4014,N_4562);
nor U5971 (N_5971,N_4045,N_4116);
nor U5972 (N_5972,N_4523,N_4144);
nand U5973 (N_5973,N_4672,N_4951);
nand U5974 (N_5974,N_4374,N_4355);
or U5975 (N_5975,N_4211,N_4486);
nand U5976 (N_5976,N_4450,N_4682);
nand U5977 (N_5977,N_4500,N_4182);
or U5978 (N_5978,N_4585,N_4974);
nand U5979 (N_5979,N_4540,N_4113);
and U5980 (N_5980,N_4445,N_4929);
nand U5981 (N_5981,N_4351,N_4853);
and U5982 (N_5982,N_4599,N_4889);
or U5983 (N_5983,N_4204,N_4598);
and U5984 (N_5984,N_4473,N_4168);
nor U5985 (N_5985,N_4421,N_4989);
and U5986 (N_5986,N_4429,N_4715);
xor U5987 (N_5987,N_4961,N_4554);
xnor U5988 (N_5988,N_4760,N_4483);
and U5989 (N_5989,N_4233,N_4067);
and U5990 (N_5990,N_4775,N_4821);
or U5991 (N_5991,N_4176,N_4879);
and U5992 (N_5992,N_4695,N_4851);
nand U5993 (N_5993,N_4487,N_4348);
xor U5994 (N_5994,N_4201,N_4922);
nand U5995 (N_5995,N_4785,N_4832);
and U5996 (N_5996,N_4671,N_4455);
and U5997 (N_5997,N_4444,N_4071);
or U5998 (N_5998,N_4274,N_4270);
or U5999 (N_5999,N_4921,N_4291);
and U6000 (N_6000,N_5152,N_5367);
nor U6001 (N_6001,N_5538,N_5450);
or U6002 (N_6002,N_5886,N_5357);
xor U6003 (N_6003,N_5487,N_5230);
nand U6004 (N_6004,N_5856,N_5278);
nand U6005 (N_6005,N_5848,N_5446);
nor U6006 (N_6006,N_5244,N_5297);
nor U6007 (N_6007,N_5322,N_5902);
nor U6008 (N_6008,N_5997,N_5277);
nand U6009 (N_6009,N_5341,N_5161);
or U6010 (N_6010,N_5876,N_5967);
and U6011 (N_6011,N_5928,N_5257);
and U6012 (N_6012,N_5234,N_5620);
or U6013 (N_6013,N_5016,N_5781);
nand U6014 (N_6014,N_5145,N_5226);
and U6015 (N_6015,N_5518,N_5738);
nand U6016 (N_6016,N_5466,N_5169);
or U6017 (N_6017,N_5205,N_5001);
nor U6018 (N_6018,N_5599,N_5535);
nor U6019 (N_6019,N_5042,N_5994);
nand U6020 (N_6020,N_5422,N_5885);
or U6021 (N_6021,N_5568,N_5028);
nor U6022 (N_6022,N_5936,N_5319);
nand U6023 (N_6023,N_5067,N_5378);
xor U6024 (N_6024,N_5424,N_5999);
nand U6025 (N_6025,N_5709,N_5521);
nand U6026 (N_6026,N_5937,N_5491);
or U6027 (N_6027,N_5340,N_5094);
and U6028 (N_6028,N_5249,N_5229);
xnor U6029 (N_6029,N_5517,N_5123);
or U6030 (N_6030,N_5023,N_5681);
nor U6031 (N_6031,N_5726,N_5460);
xnor U6032 (N_6032,N_5805,N_5283);
nor U6033 (N_6033,N_5577,N_5444);
or U6034 (N_6034,N_5966,N_5592);
and U6035 (N_6035,N_5807,N_5414);
nand U6036 (N_6036,N_5492,N_5267);
nand U6037 (N_6037,N_5076,N_5000);
nor U6038 (N_6038,N_5833,N_5552);
or U6039 (N_6039,N_5497,N_5514);
nor U6040 (N_6040,N_5273,N_5220);
xnor U6041 (N_6041,N_5306,N_5132);
and U6042 (N_6042,N_5509,N_5455);
or U6043 (N_6043,N_5558,N_5124);
or U6044 (N_6044,N_5636,N_5878);
or U6045 (N_6045,N_5930,N_5537);
nand U6046 (N_6046,N_5053,N_5772);
nor U6047 (N_6047,N_5139,N_5512);
or U6048 (N_6048,N_5810,N_5170);
nand U6049 (N_6049,N_5079,N_5173);
and U6050 (N_6050,N_5549,N_5188);
or U6051 (N_6051,N_5349,N_5111);
nor U6052 (N_6052,N_5536,N_5405);
or U6053 (N_6053,N_5945,N_5125);
xor U6054 (N_6054,N_5347,N_5740);
xnor U6055 (N_6055,N_5073,N_5468);
and U6056 (N_6056,N_5210,N_5701);
nor U6057 (N_6057,N_5473,N_5652);
nor U6058 (N_6058,N_5311,N_5873);
and U6059 (N_6059,N_5964,N_5853);
xnor U6060 (N_6060,N_5780,N_5732);
nor U6061 (N_6061,N_5179,N_5369);
or U6062 (N_6062,N_5985,N_5419);
nor U6063 (N_6063,N_5838,N_5974);
nor U6064 (N_6064,N_5486,N_5003);
xor U6065 (N_6065,N_5806,N_5065);
or U6066 (N_6066,N_5741,N_5191);
nor U6067 (N_6067,N_5934,N_5852);
nor U6068 (N_6068,N_5721,N_5617);
or U6069 (N_6069,N_5370,N_5903);
nor U6070 (N_6070,N_5742,N_5890);
and U6071 (N_6071,N_5063,N_5891);
nand U6072 (N_6072,N_5630,N_5961);
nand U6073 (N_6073,N_5379,N_5661);
and U6074 (N_6074,N_5298,N_5488);
xnor U6075 (N_6075,N_5138,N_5386);
and U6076 (N_6076,N_5397,N_5587);
nor U6077 (N_6077,N_5544,N_5476);
nand U6078 (N_6078,N_5904,N_5127);
and U6079 (N_6079,N_5368,N_5581);
nor U6080 (N_6080,N_5477,N_5449);
nand U6081 (N_6081,N_5583,N_5019);
nor U6082 (N_6082,N_5602,N_5133);
xnor U6083 (N_6083,N_5018,N_5789);
and U6084 (N_6084,N_5716,N_5889);
nand U6085 (N_6085,N_5749,N_5197);
or U6086 (N_6086,N_5295,N_5321);
nor U6087 (N_6087,N_5515,N_5922);
nand U6088 (N_6088,N_5432,N_5777);
and U6089 (N_6089,N_5899,N_5782);
or U6090 (N_6090,N_5401,N_5808);
and U6091 (N_6091,N_5005,N_5631);
nor U6092 (N_6092,N_5008,N_5024);
nand U6093 (N_6093,N_5645,N_5182);
and U6094 (N_6094,N_5639,N_5383);
nand U6095 (N_6095,N_5457,N_5122);
nor U6096 (N_6096,N_5567,N_5119);
or U6097 (N_6097,N_5157,N_5540);
or U6098 (N_6098,N_5253,N_5823);
nand U6099 (N_6099,N_5569,N_5305);
nor U6100 (N_6100,N_5025,N_5183);
and U6101 (N_6101,N_5007,N_5348);
or U6102 (N_6102,N_5235,N_5693);
nand U6103 (N_6103,N_5241,N_5164);
or U6104 (N_6104,N_5785,N_5700);
nand U6105 (N_6105,N_5570,N_5375);
and U6106 (N_6106,N_5657,N_5135);
nand U6107 (N_6107,N_5692,N_5917);
xor U6108 (N_6108,N_5925,N_5299);
nand U6109 (N_6109,N_5009,N_5771);
or U6110 (N_6110,N_5364,N_5648);
nand U6111 (N_6111,N_5409,N_5747);
and U6112 (N_6112,N_5088,N_5216);
xor U6113 (N_6113,N_5864,N_5187);
or U6114 (N_6114,N_5835,N_5167);
nand U6115 (N_6115,N_5333,N_5503);
xnor U6116 (N_6116,N_5097,N_5117);
nor U6117 (N_6117,N_5787,N_5983);
nor U6118 (N_6118,N_5354,N_5068);
and U6119 (N_6119,N_5745,N_5715);
xor U6120 (N_6120,N_5705,N_5394);
or U6121 (N_6121,N_5238,N_5213);
and U6122 (N_6122,N_5279,N_5080);
or U6123 (N_6123,N_5980,N_5776);
xor U6124 (N_6124,N_5478,N_5523);
nor U6125 (N_6125,N_5439,N_5201);
nor U6126 (N_6126,N_5353,N_5573);
xnor U6127 (N_6127,N_5935,N_5723);
xnor U6128 (N_6128,N_5165,N_5799);
nor U6129 (N_6129,N_5339,N_5734);
and U6130 (N_6130,N_5373,N_5699);
and U6131 (N_6131,N_5642,N_5438);
and U6132 (N_6132,N_5398,N_5166);
nand U6133 (N_6133,N_5108,N_5107);
and U6134 (N_6134,N_5718,N_5236);
or U6135 (N_6135,N_5707,N_5365);
and U6136 (N_6136,N_5546,N_5098);
and U6137 (N_6137,N_5109,N_5362);
or U6138 (N_6138,N_5996,N_5291);
nor U6139 (N_6139,N_5725,N_5096);
nand U6140 (N_6140,N_5040,N_5729);
nor U6141 (N_6141,N_5637,N_5194);
or U6142 (N_6142,N_5763,N_5046);
and U6143 (N_6143,N_5739,N_5323);
xnor U6144 (N_6144,N_5957,N_5453);
and U6145 (N_6145,N_5564,N_5774);
nand U6146 (N_6146,N_5162,N_5938);
xor U6147 (N_6147,N_5309,N_5672);
nand U6148 (N_6148,N_5020,N_5027);
or U6149 (N_6149,N_5982,N_5104);
nand U6150 (N_6150,N_5877,N_5614);
nand U6151 (N_6151,N_5494,N_5621);
nor U6152 (N_6152,N_5619,N_5812);
and U6153 (N_6153,N_5786,N_5268);
nor U6154 (N_6154,N_5318,N_5095);
and U6155 (N_6155,N_5842,N_5859);
nand U6156 (N_6156,N_5010,N_5381);
nor U6157 (N_6157,N_5649,N_5371);
nor U6158 (N_6158,N_5817,N_5184);
nand U6159 (N_6159,N_5428,N_5824);
or U6160 (N_6160,N_5857,N_5467);
nor U6161 (N_6161,N_5972,N_5443);
or U6162 (N_6162,N_5655,N_5626);
nor U6163 (N_6163,N_5221,N_5193);
or U6164 (N_6164,N_5499,N_5272);
nor U6165 (N_6165,N_5541,N_5261);
or U6166 (N_6166,N_5704,N_5624);
xnor U6167 (N_6167,N_5758,N_5667);
or U6168 (N_6168,N_5962,N_5662);
nand U6169 (N_6169,N_5352,N_5035);
or U6170 (N_6170,N_5588,N_5905);
and U6171 (N_6171,N_5960,N_5265);
nor U6172 (N_6172,N_5209,N_5887);
or U6173 (N_6173,N_5832,N_5604);
or U6174 (N_6174,N_5976,N_5571);
nand U6175 (N_6175,N_5836,N_5659);
nor U6176 (N_6176,N_5388,N_5811);
nor U6177 (N_6177,N_5500,N_5479);
nor U6178 (N_6178,N_5330,N_5463);
nor U6179 (N_6179,N_5384,N_5361);
or U6180 (N_6180,N_5850,N_5137);
or U6181 (N_6181,N_5783,N_5411);
nand U6182 (N_6182,N_5071,N_5189);
and U6183 (N_6183,N_5923,N_5214);
nand U6184 (N_6184,N_5075,N_5670);
nor U6185 (N_6185,N_5324,N_5565);
xor U6186 (N_6186,N_5456,N_5489);
or U6187 (N_6187,N_5128,N_5134);
or U6188 (N_6188,N_5402,N_5327);
nor U6189 (N_6189,N_5860,N_5641);
or U6190 (N_6190,N_5346,N_5882);
nor U6191 (N_6191,N_5360,N_5579);
nor U6192 (N_6192,N_5501,N_5181);
nand U6193 (N_6193,N_5580,N_5447);
xor U6194 (N_6194,N_5207,N_5440);
nor U6195 (N_6195,N_5310,N_5055);
xor U6196 (N_6196,N_5459,N_5174);
nand U6197 (N_6197,N_5144,N_5312);
xor U6198 (N_6198,N_5927,N_5643);
nor U6199 (N_6199,N_5773,N_5441);
or U6200 (N_6200,N_5968,N_5678);
nor U6201 (N_6201,N_5276,N_5633);
nor U6202 (N_6202,N_5151,N_5425);
nor U6203 (N_6203,N_5884,N_5550);
nand U6204 (N_6204,N_5513,N_5120);
or U6205 (N_6205,N_5675,N_5663);
nor U6206 (N_6206,N_5858,N_5556);
or U6207 (N_6207,N_5798,N_5710);
nand U6208 (N_6208,N_5998,N_5610);
and U6209 (N_6209,N_5290,N_5574);
or U6210 (N_6210,N_5078,N_5192);
or U6211 (N_6211,N_5613,N_5022);
or U6212 (N_6212,N_5706,N_5239);
nor U6213 (N_6213,N_5072,N_5416);
or U6214 (N_6214,N_5585,N_5228);
or U6215 (N_6215,N_5907,N_5351);
nor U6216 (N_6216,N_5851,N_5646);
xnor U6217 (N_6217,N_5262,N_5089);
or U6218 (N_6218,N_5595,N_5149);
nor U6219 (N_6219,N_5981,N_5155);
and U6220 (N_6220,N_5493,N_5286);
and U6221 (N_6221,N_5036,N_5870);
nand U6222 (N_6222,N_5644,N_5429);
nand U6223 (N_6223,N_5240,N_5387);
nor U6224 (N_6224,N_5761,N_5301);
nand U6225 (N_6225,N_5625,N_5083);
nand U6226 (N_6226,N_5287,N_5282);
nand U6227 (N_6227,N_5534,N_5284);
or U6228 (N_6228,N_5952,N_5731);
nand U6229 (N_6229,N_5926,N_5250);
nor U6230 (N_6230,N_5176,N_5408);
and U6231 (N_6231,N_5908,N_5437);
nor U6232 (N_6232,N_5325,N_5237);
xor U6233 (N_6233,N_5190,N_5914);
and U6234 (N_6234,N_5606,N_5694);
nor U6235 (N_6235,N_5628,N_5754);
or U6236 (N_6236,N_5472,N_5849);
nor U6237 (N_6237,N_5211,N_5975);
nand U6238 (N_6238,N_5147,N_5775);
nor U6239 (N_6239,N_5413,N_5006);
or U6240 (N_6240,N_5400,N_5246);
nor U6241 (N_6241,N_5334,N_5746);
nand U6242 (N_6242,N_5021,N_5991);
nand U6243 (N_6243,N_5545,N_5868);
or U6244 (N_6244,N_5059,N_5532);
nor U6245 (N_6245,N_5888,N_5591);
nand U6246 (N_6246,N_5356,N_5436);
nand U6247 (N_6247,N_5664,N_5863);
or U6248 (N_6248,N_5215,N_5920);
or U6249 (N_6249,N_5304,N_5315);
or U6250 (N_6250,N_5389,N_5854);
xor U6251 (N_6251,N_5590,N_5177);
nor U6252 (N_6252,N_5126,N_5947);
nor U6253 (N_6253,N_5730,N_5114);
nor U6254 (N_6254,N_5049,N_5392);
nand U6255 (N_6255,N_5092,N_5047);
nor U6256 (N_6256,N_5158,N_5474);
nand U6257 (N_6257,N_5665,N_5751);
or U6258 (N_6258,N_5737,N_5430);
nand U6259 (N_6259,N_5622,N_5461);
or U6260 (N_6260,N_5185,N_5690);
nor U6261 (N_6261,N_5978,N_5159);
or U6262 (N_6262,N_5482,N_5061);
nor U6263 (N_6263,N_5762,N_5115);
or U6264 (N_6264,N_5522,N_5669);
nand U6265 (N_6265,N_5252,N_5553);
nand U6266 (N_6266,N_5435,N_5847);
nand U6267 (N_6267,N_5524,N_5099);
and U6268 (N_6268,N_5320,N_5017);
and U6269 (N_6269,N_5802,N_5575);
and U6270 (N_6270,N_5171,N_5576);
or U6271 (N_6271,N_5893,N_5566);
nand U6272 (N_6272,N_5898,N_5756);
and U6273 (N_6273,N_5531,N_5691);
nand U6274 (N_6274,N_5650,N_5508);
nand U6275 (N_6275,N_5862,N_5469);
or U6276 (N_6276,N_5303,N_5004);
xnor U6277 (N_6277,N_5407,N_5562);
xnor U6278 (N_6278,N_5281,N_5377);
xnor U6279 (N_6279,N_5223,N_5970);
nand U6280 (N_6280,N_5338,N_5530);
or U6281 (N_6281,N_5933,N_5682);
or U6282 (N_6282,N_5300,N_5990);
or U6283 (N_6283,N_5412,N_5560);
and U6284 (N_6284,N_5154,N_5874);
or U6285 (N_6285,N_5778,N_5733);
or U6286 (N_6286,N_5837,N_5766);
and U6287 (N_6287,N_5979,N_5684);
or U6288 (N_6288,N_5855,N_5415);
nor U6289 (N_6289,N_5224,N_5589);
nor U6290 (N_6290,N_5484,N_5110);
or U6291 (N_6291,N_5342,N_5526);
and U6292 (N_6292,N_5288,N_5924);
xnor U6293 (N_6293,N_5584,N_5462);
or U6294 (N_6294,N_5826,N_5168);
and U6295 (N_6295,N_5698,N_5434);
or U6296 (N_6296,N_5148,N_5302);
or U6297 (N_6297,N_5984,N_5527);
nand U6298 (N_6298,N_5198,N_5054);
or U6299 (N_6299,N_5271,N_5623);
or U6300 (N_6300,N_5100,N_5728);
nor U6301 (N_6301,N_5607,N_5769);
and U6302 (N_6302,N_5951,N_5359);
or U6303 (N_6303,N_5328,N_5759);
and U6304 (N_6304,N_5085,N_5516);
xor U6305 (N_6305,N_5551,N_5506);
or U6306 (N_6306,N_5222,N_5547);
nor U6307 (N_6307,N_5175,N_5396);
nand U6308 (N_6308,N_5172,N_5112);
nor U6309 (N_6309,N_5129,N_5308);
nand U6310 (N_6310,N_5615,N_5875);
nor U6311 (N_6311,N_5895,N_5744);
xor U6312 (N_6312,N_5685,N_5445);
nand U6313 (N_6313,N_5495,N_5867);
nor U6314 (N_6314,N_5793,N_5647);
nor U6315 (N_6315,N_5792,N_5317);
or U6316 (N_6316,N_5683,N_5116);
and U6317 (N_6317,N_5247,N_5121);
or U6318 (N_6318,N_5376,N_5233);
or U6319 (N_6319,N_5616,N_5827);
and U6320 (N_6320,N_5048,N_5727);
nand U6321 (N_6321,N_5293,N_5029);
nand U6322 (N_6322,N_5421,N_5480);
and U6323 (N_6323,N_5395,N_5160);
xor U6324 (N_6324,N_5218,N_5634);
nor U6325 (N_6325,N_5753,N_5307);
nor U6326 (N_6326,N_5195,N_5217);
xnor U6327 (N_6327,N_5840,N_5956);
or U6328 (N_6328,N_5454,N_5638);
or U6329 (N_6329,N_5906,N_5433);
nor U6330 (N_6330,N_5764,N_5600);
or U6331 (N_6331,N_5912,N_5041);
xor U6332 (N_6332,N_5543,N_5343);
or U6333 (N_6333,N_5130,N_5034);
xnor U6334 (N_6334,N_5066,N_5274);
nor U6335 (N_6335,N_5426,N_5712);
and U6336 (N_6336,N_5345,N_5866);
nor U6337 (N_6337,N_5481,N_5533);
nand U6338 (N_6338,N_5724,N_5289);
nand U6339 (N_6339,N_5519,N_5861);
xnor U6340 (N_6340,N_5828,N_5654);
or U6341 (N_6341,N_5929,N_5784);
and U6342 (N_6342,N_5143,N_5788);
and U6343 (N_6343,N_5916,N_5225);
xor U6344 (N_6344,N_5910,N_5988);
or U6345 (N_6345,N_5963,N_5498);
or U6346 (N_6346,N_5880,N_5032);
xnor U6347 (N_6347,N_5163,N_5948);
or U6348 (N_6348,N_5911,N_5410);
nand U6349 (N_6349,N_5470,N_5037);
and U6350 (N_6350,N_5881,N_5314);
xnor U6351 (N_6351,N_5070,N_5743);
nand U6352 (N_6352,N_5668,N_5091);
nand U6353 (N_6353,N_5797,N_5921);
nand U6354 (N_6354,N_5131,N_5374);
nand U6355 (N_6355,N_5760,N_5485);
xnor U6356 (N_6356,N_5813,N_5033);
xor U6357 (N_6357,N_5140,N_5941);
nand U6358 (N_6358,N_5977,N_5831);
nor U6359 (N_6359,N_5475,N_5958);
and U6360 (N_6360,N_5232,N_5865);
nor U6361 (N_6361,N_5081,N_5618);
or U6362 (N_6362,N_5679,N_5755);
nand U6363 (N_6363,N_5872,N_5015);
or U6364 (N_6364,N_5993,N_5366);
nand U6365 (N_6365,N_5069,N_5082);
nor U6366 (N_6366,N_5292,N_5748);
xor U6367 (N_6367,N_5794,N_5915);
xnor U6368 (N_6368,N_5056,N_5399);
nor U6369 (N_6369,N_5103,N_5186);
or U6370 (N_6370,N_5719,N_5084);
nor U6371 (N_6371,N_5118,N_5834);
and U6372 (N_6372,N_5955,N_5629);
nand U6373 (N_6373,N_5464,N_5593);
and U6374 (N_6374,N_5057,N_5062);
or U6375 (N_6375,N_5026,N_5490);
nand U6376 (N_6376,N_5586,N_5919);
or U6377 (N_6377,N_5971,N_5953);
and U6378 (N_6378,N_5879,N_5427);
nand U6379 (N_6379,N_5231,N_5254);
nor U6380 (N_6380,N_5030,N_5313);
nand U6381 (N_6381,N_5316,N_5989);
xnor U6382 (N_6382,N_5597,N_5779);
nand U6383 (N_6383,N_5791,N_5336);
or U6384 (N_6384,N_5796,N_5263);
nor U6385 (N_6385,N_5548,N_5942);
and U6386 (N_6386,N_5954,N_5932);
xnor U6387 (N_6387,N_5757,N_5913);
and U6388 (N_6388,N_5418,N_5869);
or U6389 (N_6389,N_5382,N_5656);
xor U6390 (N_6390,N_5051,N_5448);
nand U6391 (N_6391,N_5736,N_5156);
nor U6392 (N_6392,N_5843,N_5039);
nand U6393 (N_6393,N_5363,N_5946);
nand U6394 (N_6394,N_5845,N_5901);
nand U6395 (N_6395,N_5578,N_5245);
and U6396 (N_6396,N_5871,N_5821);
or U6397 (N_6397,N_5417,N_5973);
nor U6398 (N_6398,N_5391,N_5511);
nor U6399 (N_6399,N_5202,N_5203);
nand U6400 (N_6400,N_5206,N_5270);
and U6401 (N_6401,N_5332,N_5087);
nor U6402 (N_6402,N_5093,N_5212);
and U6403 (N_6403,N_5529,N_5819);
or U6404 (N_6404,N_5703,N_5605);
nor U6405 (N_6405,N_5180,N_5940);
and U6406 (N_6406,N_5052,N_5702);
or U6407 (N_6407,N_5248,N_5809);
nor U6408 (N_6408,N_5259,N_5451);
nor U6409 (N_6409,N_5582,N_5897);
and U6410 (N_6410,N_5086,N_5839);
and U6411 (N_6411,N_5038,N_5825);
and U6412 (N_6412,N_5077,N_5064);
or U6413 (N_6413,N_5750,N_5594);
nor U6414 (N_6414,N_5204,N_5720);
or U6415 (N_6415,N_5818,N_5014);
nor U6416 (N_6416,N_5815,N_5200);
nand U6417 (N_6417,N_5931,N_5502);
xor U6418 (N_6418,N_5687,N_5385);
and U6419 (N_6419,N_5520,N_5596);
xnor U6420 (N_6420,N_5102,N_5950);
or U6421 (N_6421,N_5909,N_5695);
nand U6422 (N_6422,N_5141,N_5572);
nor U6423 (N_6423,N_5329,N_5651);
and U6424 (N_6424,N_5803,N_5767);
nor U6425 (N_6425,N_5708,N_5561);
nand U6426 (N_6426,N_5074,N_5752);
nand U6427 (N_6427,N_5528,N_5559);
nand U6428 (N_6428,N_5714,N_5403);
and U6429 (N_6429,N_5260,N_5563);
and U6430 (N_6430,N_5894,N_5722);
nor U6431 (N_6431,N_5680,N_5106);
nor U6432 (N_6432,N_5986,N_5830);
nand U6433 (N_6433,N_5697,N_5790);
nand U6434 (N_6434,N_5471,N_5465);
nand U6435 (N_6435,N_5804,N_5243);
and U6436 (N_6436,N_5280,N_5442);
nand U6437 (N_6437,N_5542,N_5992);
and U6438 (N_6438,N_5673,N_5969);
and U6439 (N_6439,N_5711,N_5632);
nor U6440 (N_6440,N_5380,N_5653);
and U6441 (N_6441,N_5452,N_5770);
and U6442 (N_6442,N_5671,N_5331);
nand U6443 (N_6443,N_5153,N_5601);
and U6444 (N_6444,N_5717,N_5255);
xnor U6445 (N_6445,N_5900,N_5688);
nor U6446 (N_6446,N_5136,N_5355);
and U6447 (N_6447,N_5326,N_5058);
nor U6448 (N_6448,N_5258,N_5603);
nand U6449 (N_6449,N_5372,N_5674);
or U6450 (N_6450,N_5251,N_5660);
and U6451 (N_6451,N_5294,N_5199);
xor U6452 (N_6452,N_5113,N_5892);
and U6453 (N_6453,N_5987,N_5696);
nor U6454 (N_6454,N_5390,N_5045);
nand U6455 (N_6455,N_5800,N_5949);
nor U6456 (N_6456,N_5196,N_5814);
or U6457 (N_6457,N_5505,N_5609);
nor U6458 (N_6458,N_5918,N_5256);
nor U6459 (N_6459,N_5677,N_5829);
xor U6460 (N_6460,N_5735,N_5423);
or U6461 (N_6461,N_5612,N_5939);
or U6462 (N_6462,N_5011,N_5142);
and U6463 (N_6463,N_5611,N_5795);
or U6464 (N_6464,N_5350,N_5598);
nor U6465 (N_6465,N_5208,N_5816);
nand U6466 (N_6466,N_5608,N_5496);
and U6467 (N_6467,N_5554,N_5344);
nand U6468 (N_6468,N_5995,N_5101);
or U6469 (N_6469,N_5676,N_5844);
nand U6470 (N_6470,N_5146,N_5959);
and U6471 (N_6471,N_5090,N_5285);
xor U6472 (N_6472,N_5105,N_5266);
nand U6473 (N_6473,N_5635,N_5557);
and U6474 (N_6474,N_5896,N_5943);
and U6475 (N_6475,N_5765,N_5504);
nand U6476 (N_6476,N_5846,N_5012);
nor U6477 (N_6477,N_5510,N_5713);
nand U6478 (N_6478,N_5883,N_5337);
xnor U6479 (N_6479,N_5640,N_5275);
or U6480 (N_6480,N_5404,N_5539);
and U6481 (N_6481,N_5335,N_5841);
nor U6482 (N_6482,N_5483,N_5525);
or U6483 (N_6483,N_5031,N_5666);
xnor U6484 (N_6484,N_5264,N_5555);
or U6485 (N_6485,N_5178,N_5420);
or U6486 (N_6486,N_5043,N_5269);
and U6487 (N_6487,N_5219,N_5013);
and U6488 (N_6488,N_5431,N_5458);
or U6489 (N_6489,N_5507,N_5801);
nor U6490 (N_6490,N_5358,N_5820);
nor U6491 (N_6491,N_5627,N_5050);
or U6492 (N_6492,N_5768,N_5060);
and U6493 (N_6493,N_5689,N_5150);
or U6494 (N_6494,N_5242,N_5965);
nand U6495 (N_6495,N_5686,N_5406);
nor U6496 (N_6496,N_5296,N_5944);
or U6497 (N_6497,N_5002,N_5227);
and U6498 (N_6498,N_5822,N_5393);
xnor U6499 (N_6499,N_5044,N_5658);
or U6500 (N_6500,N_5854,N_5134);
nand U6501 (N_6501,N_5153,N_5841);
and U6502 (N_6502,N_5309,N_5633);
or U6503 (N_6503,N_5510,N_5001);
nor U6504 (N_6504,N_5957,N_5355);
or U6505 (N_6505,N_5932,N_5824);
nor U6506 (N_6506,N_5524,N_5876);
or U6507 (N_6507,N_5045,N_5205);
nor U6508 (N_6508,N_5158,N_5964);
and U6509 (N_6509,N_5775,N_5381);
nor U6510 (N_6510,N_5302,N_5268);
xor U6511 (N_6511,N_5040,N_5196);
nor U6512 (N_6512,N_5267,N_5731);
or U6513 (N_6513,N_5607,N_5214);
nand U6514 (N_6514,N_5733,N_5569);
nand U6515 (N_6515,N_5502,N_5978);
or U6516 (N_6516,N_5085,N_5732);
nor U6517 (N_6517,N_5390,N_5159);
nor U6518 (N_6518,N_5070,N_5301);
or U6519 (N_6519,N_5983,N_5869);
or U6520 (N_6520,N_5028,N_5180);
and U6521 (N_6521,N_5423,N_5726);
and U6522 (N_6522,N_5918,N_5120);
nand U6523 (N_6523,N_5310,N_5715);
and U6524 (N_6524,N_5911,N_5507);
nor U6525 (N_6525,N_5376,N_5168);
or U6526 (N_6526,N_5441,N_5640);
or U6527 (N_6527,N_5340,N_5444);
nand U6528 (N_6528,N_5739,N_5362);
or U6529 (N_6529,N_5233,N_5384);
and U6530 (N_6530,N_5411,N_5614);
or U6531 (N_6531,N_5818,N_5402);
and U6532 (N_6532,N_5498,N_5306);
nand U6533 (N_6533,N_5624,N_5397);
nor U6534 (N_6534,N_5194,N_5574);
nand U6535 (N_6535,N_5801,N_5949);
and U6536 (N_6536,N_5300,N_5847);
nand U6537 (N_6537,N_5256,N_5972);
and U6538 (N_6538,N_5762,N_5641);
nor U6539 (N_6539,N_5906,N_5488);
nor U6540 (N_6540,N_5491,N_5275);
and U6541 (N_6541,N_5372,N_5499);
nor U6542 (N_6542,N_5064,N_5246);
nand U6543 (N_6543,N_5962,N_5086);
or U6544 (N_6544,N_5726,N_5207);
xnor U6545 (N_6545,N_5032,N_5675);
xor U6546 (N_6546,N_5255,N_5283);
or U6547 (N_6547,N_5218,N_5646);
and U6548 (N_6548,N_5516,N_5668);
nand U6549 (N_6549,N_5248,N_5099);
nor U6550 (N_6550,N_5272,N_5725);
nor U6551 (N_6551,N_5138,N_5902);
and U6552 (N_6552,N_5269,N_5179);
nor U6553 (N_6553,N_5808,N_5095);
and U6554 (N_6554,N_5273,N_5107);
xnor U6555 (N_6555,N_5910,N_5334);
nor U6556 (N_6556,N_5674,N_5943);
nor U6557 (N_6557,N_5868,N_5294);
or U6558 (N_6558,N_5838,N_5402);
or U6559 (N_6559,N_5895,N_5572);
nand U6560 (N_6560,N_5935,N_5842);
nand U6561 (N_6561,N_5295,N_5328);
or U6562 (N_6562,N_5888,N_5441);
nand U6563 (N_6563,N_5746,N_5804);
and U6564 (N_6564,N_5924,N_5858);
or U6565 (N_6565,N_5242,N_5220);
nor U6566 (N_6566,N_5289,N_5300);
nand U6567 (N_6567,N_5529,N_5401);
xnor U6568 (N_6568,N_5948,N_5083);
and U6569 (N_6569,N_5710,N_5262);
or U6570 (N_6570,N_5662,N_5828);
or U6571 (N_6571,N_5656,N_5396);
and U6572 (N_6572,N_5460,N_5224);
and U6573 (N_6573,N_5555,N_5307);
xor U6574 (N_6574,N_5855,N_5858);
or U6575 (N_6575,N_5211,N_5388);
xnor U6576 (N_6576,N_5785,N_5957);
nand U6577 (N_6577,N_5315,N_5519);
or U6578 (N_6578,N_5501,N_5359);
or U6579 (N_6579,N_5308,N_5495);
nor U6580 (N_6580,N_5611,N_5083);
or U6581 (N_6581,N_5104,N_5258);
nor U6582 (N_6582,N_5724,N_5741);
nor U6583 (N_6583,N_5520,N_5020);
nand U6584 (N_6584,N_5195,N_5958);
or U6585 (N_6585,N_5837,N_5262);
nand U6586 (N_6586,N_5813,N_5461);
or U6587 (N_6587,N_5658,N_5449);
and U6588 (N_6588,N_5799,N_5821);
nand U6589 (N_6589,N_5151,N_5689);
or U6590 (N_6590,N_5682,N_5989);
or U6591 (N_6591,N_5845,N_5149);
and U6592 (N_6592,N_5280,N_5268);
nand U6593 (N_6593,N_5878,N_5000);
xnor U6594 (N_6594,N_5711,N_5873);
and U6595 (N_6595,N_5529,N_5864);
nand U6596 (N_6596,N_5209,N_5920);
or U6597 (N_6597,N_5561,N_5572);
and U6598 (N_6598,N_5869,N_5935);
nor U6599 (N_6599,N_5050,N_5608);
nand U6600 (N_6600,N_5674,N_5445);
nor U6601 (N_6601,N_5446,N_5064);
nand U6602 (N_6602,N_5392,N_5727);
nor U6603 (N_6603,N_5679,N_5507);
nor U6604 (N_6604,N_5203,N_5732);
nor U6605 (N_6605,N_5157,N_5738);
and U6606 (N_6606,N_5129,N_5057);
nand U6607 (N_6607,N_5054,N_5340);
or U6608 (N_6608,N_5497,N_5766);
nor U6609 (N_6609,N_5618,N_5979);
and U6610 (N_6610,N_5814,N_5022);
or U6611 (N_6611,N_5586,N_5207);
nor U6612 (N_6612,N_5527,N_5090);
and U6613 (N_6613,N_5906,N_5361);
nor U6614 (N_6614,N_5699,N_5040);
nor U6615 (N_6615,N_5707,N_5318);
nor U6616 (N_6616,N_5769,N_5906);
xor U6617 (N_6617,N_5556,N_5639);
or U6618 (N_6618,N_5330,N_5788);
nor U6619 (N_6619,N_5394,N_5411);
and U6620 (N_6620,N_5446,N_5578);
xor U6621 (N_6621,N_5281,N_5657);
nor U6622 (N_6622,N_5450,N_5719);
nor U6623 (N_6623,N_5734,N_5295);
or U6624 (N_6624,N_5415,N_5932);
nand U6625 (N_6625,N_5796,N_5916);
nand U6626 (N_6626,N_5977,N_5975);
nor U6627 (N_6627,N_5410,N_5540);
nand U6628 (N_6628,N_5937,N_5713);
or U6629 (N_6629,N_5505,N_5830);
or U6630 (N_6630,N_5833,N_5612);
nor U6631 (N_6631,N_5430,N_5216);
xnor U6632 (N_6632,N_5390,N_5730);
or U6633 (N_6633,N_5005,N_5269);
nand U6634 (N_6634,N_5733,N_5079);
nand U6635 (N_6635,N_5408,N_5605);
nand U6636 (N_6636,N_5925,N_5002);
or U6637 (N_6637,N_5459,N_5693);
nor U6638 (N_6638,N_5444,N_5439);
and U6639 (N_6639,N_5716,N_5030);
or U6640 (N_6640,N_5976,N_5152);
or U6641 (N_6641,N_5662,N_5785);
nor U6642 (N_6642,N_5819,N_5451);
nand U6643 (N_6643,N_5662,N_5727);
nor U6644 (N_6644,N_5215,N_5392);
nand U6645 (N_6645,N_5110,N_5702);
or U6646 (N_6646,N_5972,N_5323);
xor U6647 (N_6647,N_5468,N_5391);
nor U6648 (N_6648,N_5312,N_5705);
or U6649 (N_6649,N_5841,N_5485);
nand U6650 (N_6650,N_5764,N_5036);
xnor U6651 (N_6651,N_5097,N_5641);
nor U6652 (N_6652,N_5987,N_5895);
and U6653 (N_6653,N_5905,N_5387);
nand U6654 (N_6654,N_5388,N_5543);
and U6655 (N_6655,N_5216,N_5534);
nor U6656 (N_6656,N_5592,N_5718);
and U6657 (N_6657,N_5403,N_5128);
or U6658 (N_6658,N_5012,N_5680);
nor U6659 (N_6659,N_5304,N_5425);
xor U6660 (N_6660,N_5355,N_5360);
or U6661 (N_6661,N_5508,N_5774);
or U6662 (N_6662,N_5799,N_5996);
and U6663 (N_6663,N_5344,N_5200);
or U6664 (N_6664,N_5406,N_5616);
or U6665 (N_6665,N_5387,N_5174);
or U6666 (N_6666,N_5468,N_5040);
and U6667 (N_6667,N_5109,N_5413);
and U6668 (N_6668,N_5050,N_5047);
xnor U6669 (N_6669,N_5271,N_5664);
nor U6670 (N_6670,N_5276,N_5656);
nor U6671 (N_6671,N_5136,N_5810);
nand U6672 (N_6672,N_5689,N_5154);
xnor U6673 (N_6673,N_5317,N_5901);
or U6674 (N_6674,N_5537,N_5459);
or U6675 (N_6675,N_5254,N_5223);
nor U6676 (N_6676,N_5020,N_5098);
and U6677 (N_6677,N_5998,N_5100);
or U6678 (N_6678,N_5438,N_5207);
and U6679 (N_6679,N_5529,N_5845);
nor U6680 (N_6680,N_5816,N_5015);
nor U6681 (N_6681,N_5406,N_5436);
and U6682 (N_6682,N_5046,N_5074);
nor U6683 (N_6683,N_5250,N_5960);
and U6684 (N_6684,N_5508,N_5990);
and U6685 (N_6685,N_5407,N_5172);
nor U6686 (N_6686,N_5941,N_5308);
or U6687 (N_6687,N_5466,N_5892);
nor U6688 (N_6688,N_5925,N_5571);
xnor U6689 (N_6689,N_5238,N_5942);
nand U6690 (N_6690,N_5363,N_5079);
nor U6691 (N_6691,N_5204,N_5278);
xnor U6692 (N_6692,N_5337,N_5066);
nand U6693 (N_6693,N_5304,N_5710);
nand U6694 (N_6694,N_5530,N_5816);
and U6695 (N_6695,N_5502,N_5539);
or U6696 (N_6696,N_5903,N_5849);
nand U6697 (N_6697,N_5709,N_5051);
nand U6698 (N_6698,N_5827,N_5874);
and U6699 (N_6699,N_5673,N_5210);
and U6700 (N_6700,N_5708,N_5494);
and U6701 (N_6701,N_5560,N_5552);
nand U6702 (N_6702,N_5387,N_5597);
and U6703 (N_6703,N_5047,N_5920);
nor U6704 (N_6704,N_5068,N_5869);
or U6705 (N_6705,N_5254,N_5202);
nand U6706 (N_6706,N_5617,N_5917);
and U6707 (N_6707,N_5753,N_5395);
and U6708 (N_6708,N_5981,N_5517);
nor U6709 (N_6709,N_5180,N_5188);
and U6710 (N_6710,N_5690,N_5242);
and U6711 (N_6711,N_5233,N_5070);
or U6712 (N_6712,N_5747,N_5400);
nand U6713 (N_6713,N_5325,N_5809);
and U6714 (N_6714,N_5430,N_5537);
and U6715 (N_6715,N_5769,N_5982);
nand U6716 (N_6716,N_5141,N_5069);
or U6717 (N_6717,N_5677,N_5913);
nand U6718 (N_6718,N_5299,N_5342);
xor U6719 (N_6719,N_5855,N_5007);
nand U6720 (N_6720,N_5239,N_5233);
and U6721 (N_6721,N_5570,N_5889);
and U6722 (N_6722,N_5560,N_5292);
and U6723 (N_6723,N_5526,N_5503);
and U6724 (N_6724,N_5285,N_5642);
or U6725 (N_6725,N_5616,N_5115);
or U6726 (N_6726,N_5159,N_5592);
and U6727 (N_6727,N_5930,N_5624);
nand U6728 (N_6728,N_5678,N_5344);
and U6729 (N_6729,N_5009,N_5764);
nor U6730 (N_6730,N_5367,N_5443);
nand U6731 (N_6731,N_5342,N_5730);
and U6732 (N_6732,N_5674,N_5982);
and U6733 (N_6733,N_5033,N_5464);
or U6734 (N_6734,N_5042,N_5468);
and U6735 (N_6735,N_5477,N_5157);
and U6736 (N_6736,N_5964,N_5652);
nor U6737 (N_6737,N_5387,N_5604);
nand U6738 (N_6738,N_5876,N_5746);
and U6739 (N_6739,N_5049,N_5345);
nor U6740 (N_6740,N_5474,N_5463);
nand U6741 (N_6741,N_5713,N_5582);
xor U6742 (N_6742,N_5218,N_5847);
nor U6743 (N_6743,N_5005,N_5729);
nand U6744 (N_6744,N_5425,N_5983);
nand U6745 (N_6745,N_5176,N_5009);
nor U6746 (N_6746,N_5766,N_5928);
nand U6747 (N_6747,N_5723,N_5251);
xor U6748 (N_6748,N_5020,N_5969);
nand U6749 (N_6749,N_5855,N_5206);
nand U6750 (N_6750,N_5568,N_5899);
and U6751 (N_6751,N_5226,N_5242);
nor U6752 (N_6752,N_5262,N_5369);
nand U6753 (N_6753,N_5266,N_5090);
nand U6754 (N_6754,N_5818,N_5023);
xnor U6755 (N_6755,N_5578,N_5645);
or U6756 (N_6756,N_5868,N_5331);
and U6757 (N_6757,N_5955,N_5082);
or U6758 (N_6758,N_5314,N_5327);
xor U6759 (N_6759,N_5342,N_5721);
nor U6760 (N_6760,N_5389,N_5348);
nor U6761 (N_6761,N_5138,N_5702);
nand U6762 (N_6762,N_5300,N_5476);
nand U6763 (N_6763,N_5174,N_5798);
xor U6764 (N_6764,N_5057,N_5454);
or U6765 (N_6765,N_5887,N_5654);
and U6766 (N_6766,N_5080,N_5775);
nor U6767 (N_6767,N_5313,N_5446);
xor U6768 (N_6768,N_5036,N_5981);
and U6769 (N_6769,N_5526,N_5970);
nand U6770 (N_6770,N_5769,N_5736);
and U6771 (N_6771,N_5954,N_5938);
nor U6772 (N_6772,N_5583,N_5942);
and U6773 (N_6773,N_5514,N_5753);
and U6774 (N_6774,N_5360,N_5264);
nand U6775 (N_6775,N_5241,N_5078);
or U6776 (N_6776,N_5062,N_5460);
and U6777 (N_6777,N_5029,N_5590);
xor U6778 (N_6778,N_5005,N_5939);
nor U6779 (N_6779,N_5817,N_5172);
nor U6780 (N_6780,N_5970,N_5626);
nor U6781 (N_6781,N_5469,N_5992);
nor U6782 (N_6782,N_5764,N_5169);
nand U6783 (N_6783,N_5125,N_5863);
nand U6784 (N_6784,N_5819,N_5687);
nand U6785 (N_6785,N_5378,N_5142);
nand U6786 (N_6786,N_5103,N_5020);
and U6787 (N_6787,N_5766,N_5429);
or U6788 (N_6788,N_5352,N_5283);
nor U6789 (N_6789,N_5180,N_5557);
and U6790 (N_6790,N_5347,N_5411);
nand U6791 (N_6791,N_5026,N_5806);
nand U6792 (N_6792,N_5969,N_5613);
and U6793 (N_6793,N_5043,N_5169);
nor U6794 (N_6794,N_5480,N_5007);
and U6795 (N_6795,N_5823,N_5268);
or U6796 (N_6796,N_5464,N_5217);
nor U6797 (N_6797,N_5146,N_5714);
nor U6798 (N_6798,N_5115,N_5530);
nand U6799 (N_6799,N_5915,N_5938);
nor U6800 (N_6800,N_5529,N_5897);
nor U6801 (N_6801,N_5725,N_5182);
or U6802 (N_6802,N_5933,N_5261);
nand U6803 (N_6803,N_5392,N_5585);
and U6804 (N_6804,N_5238,N_5617);
or U6805 (N_6805,N_5452,N_5272);
nor U6806 (N_6806,N_5175,N_5162);
nand U6807 (N_6807,N_5977,N_5707);
nor U6808 (N_6808,N_5218,N_5561);
or U6809 (N_6809,N_5205,N_5294);
xor U6810 (N_6810,N_5545,N_5898);
nand U6811 (N_6811,N_5325,N_5860);
nor U6812 (N_6812,N_5621,N_5711);
nor U6813 (N_6813,N_5686,N_5843);
and U6814 (N_6814,N_5128,N_5095);
nor U6815 (N_6815,N_5912,N_5883);
xnor U6816 (N_6816,N_5717,N_5137);
and U6817 (N_6817,N_5186,N_5755);
nor U6818 (N_6818,N_5596,N_5228);
xnor U6819 (N_6819,N_5420,N_5269);
nor U6820 (N_6820,N_5489,N_5505);
and U6821 (N_6821,N_5929,N_5197);
and U6822 (N_6822,N_5155,N_5567);
nor U6823 (N_6823,N_5517,N_5070);
nor U6824 (N_6824,N_5589,N_5892);
and U6825 (N_6825,N_5330,N_5161);
xor U6826 (N_6826,N_5582,N_5964);
nand U6827 (N_6827,N_5192,N_5044);
nor U6828 (N_6828,N_5076,N_5167);
nand U6829 (N_6829,N_5072,N_5387);
xor U6830 (N_6830,N_5483,N_5570);
and U6831 (N_6831,N_5383,N_5763);
or U6832 (N_6832,N_5459,N_5926);
or U6833 (N_6833,N_5652,N_5504);
or U6834 (N_6834,N_5127,N_5655);
nand U6835 (N_6835,N_5939,N_5548);
nor U6836 (N_6836,N_5293,N_5631);
xor U6837 (N_6837,N_5930,N_5771);
xnor U6838 (N_6838,N_5980,N_5546);
and U6839 (N_6839,N_5666,N_5925);
nand U6840 (N_6840,N_5414,N_5684);
nor U6841 (N_6841,N_5615,N_5706);
xnor U6842 (N_6842,N_5022,N_5415);
nand U6843 (N_6843,N_5762,N_5864);
and U6844 (N_6844,N_5980,N_5884);
or U6845 (N_6845,N_5667,N_5887);
and U6846 (N_6846,N_5383,N_5922);
and U6847 (N_6847,N_5225,N_5781);
xnor U6848 (N_6848,N_5580,N_5736);
or U6849 (N_6849,N_5665,N_5817);
and U6850 (N_6850,N_5530,N_5153);
or U6851 (N_6851,N_5101,N_5609);
and U6852 (N_6852,N_5877,N_5885);
or U6853 (N_6853,N_5757,N_5584);
nand U6854 (N_6854,N_5904,N_5167);
nand U6855 (N_6855,N_5595,N_5516);
or U6856 (N_6856,N_5250,N_5102);
or U6857 (N_6857,N_5567,N_5912);
nor U6858 (N_6858,N_5620,N_5484);
and U6859 (N_6859,N_5013,N_5413);
or U6860 (N_6860,N_5145,N_5555);
xor U6861 (N_6861,N_5242,N_5267);
nor U6862 (N_6862,N_5635,N_5249);
nand U6863 (N_6863,N_5009,N_5271);
and U6864 (N_6864,N_5518,N_5350);
or U6865 (N_6865,N_5112,N_5755);
or U6866 (N_6866,N_5877,N_5183);
nor U6867 (N_6867,N_5223,N_5367);
nor U6868 (N_6868,N_5987,N_5524);
nor U6869 (N_6869,N_5910,N_5381);
nand U6870 (N_6870,N_5135,N_5383);
or U6871 (N_6871,N_5347,N_5961);
nand U6872 (N_6872,N_5963,N_5455);
and U6873 (N_6873,N_5059,N_5268);
or U6874 (N_6874,N_5763,N_5107);
nand U6875 (N_6875,N_5384,N_5111);
and U6876 (N_6876,N_5229,N_5951);
nand U6877 (N_6877,N_5797,N_5756);
nor U6878 (N_6878,N_5525,N_5773);
and U6879 (N_6879,N_5192,N_5357);
or U6880 (N_6880,N_5125,N_5407);
nand U6881 (N_6881,N_5456,N_5636);
and U6882 (N_6882,N_5183,N_5559);
nor U6883 (N_6883,N_5296,N_5441);
nand U6884 (N_6884,N_5475,N_5405);
and U6885 (N_6885,N_5545,N_5251);
nor U6886 (N_6886,N_5818,N_5156);
or U6887 (N_6887,N_5011,N_5546);
nor U6888 (N_6888,N_5452,N_5743);
nor U6889 (N_6889,N_5040,N_5924);
and U6890 (N_6890,N_5814,N_5289);
or U6891 (N_6891,N_5997,N_5915);
nor U6892 (N_6892,N_5953,N_5081);
and U6893 (N_6893,N_5362,N_5703);
or U6894 (N_6894,N_5539,N_5263);
nor U6895 (N_6895,N_5494,N_5213);
nor U6896 (N_6896,N_5067,N_5775);
xnor U6897 (N_6897,N_5734,N_5465);
nor U6898 (N_6898,N_5267,N_5420);
and U6899 (N_6899,N_5936,N_5533);
and U6900 (N_6900,N_5276,N_5450);
nor U6901 (N_6901,N_5102,N_5078);
or U6902 (N_6902,N_5213,N_5503);
and U6903 (N_6903,N_5398,N_5648);
and U6904 (N_6904,N_5451,N_5396);
xor U6905 (N_6905,N_5712,N_5694);
or U6906 (N_6906,N_5161,N_5417);
nor U6907 (N_6907,N_5425,N_5807);
nor U6908 (N_6908,N_5533,N_5995);
xnor U6909 (N_6909,N_5239,N_5763);
nor U6910 (N_6910,N_5373,N_5963);
and U6911 (N_6911,N_5044,N_5599);
or U6912 (N_6912,N_5871,N_5149);
or U6913 (N_6913,N_5524,N_5674);
and U6914 (N_6914,N_5730,N_5666);
or U6915 (N_6915,N_5897,N_5420);
and U6916 (N_6916,N_5151,N_5817);
nor U6917 (N_6917,N_5035,N_5426);
nor U6918 (N_6918,N_5911,N_5712);
nor U6919 (N_6919,N_5881,N_5264);
nand U6920 (N_6920,N_5125,N_5296);
nor U6921 (N_6921,N_5812,N_5243);
xor U6922 (N_6922,N_5090,N_5499);
nand U6923 (N_6923,N_5267,N_5340);
nor U6924 (N_6924,N_5963,N_5950);
and U6925 (N_6925,N_5937,N_5755);
nand U6926 (N_6926,N_5384,N_5746);
and U6927 (N_6927,N_5340,N_5268);
or U6928 (N_6928,N_5142,N_5725);
xnor U6929 (N_6929,N_5089,N_5847);
nor U6930 (N_6930,N_5265,N_5916);
and U6931 (N_6931,N_5699,N_5327);
nor U6932 (N_6932,N_5410,N_5841);
or U6933 (N_6933,N_5246,N_5577);
nor U6934 (N_6934,N_5390,N_5897);
and U6935 (N_6935,N_5057,N_5353);
nor U6936 (N_6936,N_5921,N_5012);
nand U6937 (N_6937,N_5049,N_5467);
nor U6938 (N_6938,N_5598,N_5832);
or U6939 (N_6939,N_5046,N_5535);
or U6940 (N_6940,N_5105,N_5849);
and U6941 (N_6941,N_5017,N_5878);
nor U6942 (N_6942,N_5706,N_5803);
or U6943 (N_6943,N_5178,N_5288);
nor U6944 (N_6944,N_5044,N_5288);
nor U6945 (N_6945,N_5250,N_5016);
nand U6946 (N_6946,N_5204,N_5692);
nor U6947 (N_6947,N_5641,N_5619);
nand U6948 (N_6948,N_5669,N_5699);
and U6949 (N_6949,N_5813,N_5258);
and U6950 (N_6950,N_5113,N_5390);
nand U6951 (N_6951,N_5486,N_5255);
nor U6952 (N_6952,N_5542,N_5363);
nor U6953 (N_6953,N_5547,N_5103);
nand U6954 (N_6954,N_5435,N_5282);
nor U6955 (N_6955,N_5762,N_5723);
nor U6956 (N_6956,N_5275,N_5218);
nand U6957 (N_6957,N_5612,N_5641);
nand U6958 (N_6958,N_5869,N_5311);
nand U6959 (N_6959,N_5216,N_5558);
and U6960 (N_6960,N_5583,N_5593);
nor U6961 (N_6961,N_5406,N_5061);
or U6962 (N_6962,N_5862,N_5513);
xor U6963 (N_6963,N_5990,N_5175);
nand U6964 (N_6964,N_5673,N_5203);
or U6965 (N_6965,N_5786,N_5285);
and U6966 (N_6966,N_5591,N_5681);
and U6967 (N_6967,N_5930,N_5611);
xnor U6968 (N_6968,N_5972,N_5740);
nand U6969 (N_6969,N_5066,N_5435);
or U6970 (N_6970,N_5630,N_5805);
nand U6971 (N_6971,N_5551,N_5479);
nand U6972 (N_6972,N_5371,N_5920);
or U6973 (N_6973,N_5259,N_5093);
or U6974 (N_6974,N_5902,N_5574);
nand U6975 (N_6975,N_5468,N_5352);
nor U6976 (N_6976,N_5710,N_5951);
and U6977 (N_6977,N_5966,N_5315);
nor U6978 (N_6978,N_5967,N_5046);
and U6979 (N_6979,N_5814,N_5887);
and U6980 (N_6980,N_5327,N_5095);
nand U6981 (N_6981,N_5566,N_5927);
xor U6982 (N_6982,N_5889,N_5852);
nand U6983 (N_6983,N_5688,N_5133);
nor U6984 (N_6984,N_5992,N_5493);
and U6985 (N_6985,N_5298,N_5095);
nand U6986 (N_6986,N_5536,N_5022);
or U6987 (N_6987,N_5923,N_5192);
nand U6988 (N_6988,N_5338,N_5973);
or U6989 (N_6989,N_5053,N_5594);
and U6990 (N_6990,N_5477,N_5750);
or U6991 (N_6991,N_5517,N_5850);
nor U6992 (N_6992,N_5047,N_5963);
nor U6993 (N_6993,N_5981,N_5525);
nor U6994 (N_6994,N_5305,N_5817);
nand U6995 (N_6995,N_5547,N_5388);
xnor U6996 (N_6996,N_5607,N_5945);
nand U6997 (N_6997,N_5443,N_5685);
xnor U6998 (N_6998,N_5421,N_5163);
or U6999 (N_6999,N_5593,N_5838);
and U7000 (N_7000,N_6265,N_6826);
or U7001 (N_7001,N_6627,N_6909);
or U7002 (N_7002,N_6078,N_6861);
xnor U7003 (N_7003,N_6105,N_6577);
xor U7004 (N_7004,N_6772,N_6456);
and U7005 (N_7005,N_6677,N_6704);
nor U7006 (N_7006,N_6457,N_6428);
xor U7007 (N_7007,N_6696,N_6431);
or U7008 (N_7008,N_6363,N_6328);
nor U7009 (N_7009,N_6816,N_6572);
xor U7010 (N_7010,N_6857,N_6998);
nor U7011 (N_7011,N_6322,N_6372);
nor U7012 (N_7012,N_6036,N_6808);
nor U7013 (N_7013,N_6586,N_6634);
nand U7014 (N_7014,N_6256,N_6158);
nand U7015 (N_7015,N_6992,N_6921);
or U7016 (N_7016,N_6181,N_6805);
and U7017 (N_7017,N_6811,N_6734);
nor U7018 (N_7018,N_6050,N_6932);
and U7019 (N_7019,N_6842,N_6668);
xnor U7020 (N_7020,N_6370,N_6700);
xnor U7021 (N_7021,N_6818,N_6764);
or U7022 (N_7022,N_6641,N_6989);
nand U7023 (N_7023,N_6447,N_6832);
nor U7024 (N_7024,N_6865,N_6217);
nand U7025 (N_7025,N_6664,N_6613);
nand U7026 (N_7026,N_6883,N_6578);
and U7027 (N_7027,N_6895,N_6305);
nor U7028 (N_7028,N_6748,N_6547);
or U7029 (N_7029,N_6040,N_6488);
or U7030 (N_7030,N_6144,N_6569);
or U7031 (N_7031,N_6039,N_6684);
nor U7032 (N_7032,N_6557,N_6168);
nand U7033 (N_7033,N_6096,N_6203);
nand U7034 (N_7034,N_6853,N_6373);
or U7035 (N_7035,N_6012,N_6837);
or U7036 (N_7036,N_6450,N_6443);
nand U7037 (N_7037,N_6133,N_6983);
or U7038 (N_7038,N_6283,N_6874);
nand U7039 (N_7039,N_6219,N_6064);
or U7040 (N_7040,N_6500,N_6136);
xnor U7041 (N_7041,N_6121,N_6714);
nor U7042 (N_7042,N_6946,N_6942);
and U7043 (N_7043,N_6884,N_6379);
or U7044 (N_7044,N_6900,N_6108);
and U7045 (N_7045,N_6002,N_6615);
or U7046 (N_7046,N_6384,N_6342);
or U7047 (N_7047,N_6828,N_6100);
and U7048 (N_7048,N_6898,N_6427);
xnor U7049 (N_7049,N_6730,N_6074);
nand U7050 (N_7050,N_6391,N_6639);
or U7051 (N_7051,N_6389,N_6424);
nor U7052 (N_7052,N_6863,N_6513);
nand U7053 (N_7053,N_6997,N_6119);
or U7054 (N_7054,N_6381,N_6423);
nor U7055 (N_7055,N_6887,N_6545);
and U7056 (N_7056,N_6127,N_6749);
and U7057 (N_7057,N_6830,N_6101);
and U7058 (N_7058,N_6049,N_6231);
and U7059 (N_7059,N_6948,N_6798);
and U7060 (N_7060,N_6258,N_6114);
or U7061 (N_7061,N_6848,N_6924);
nand U7062 (N_7062,N_6622,N_6580);
xnor U7063 (N_7063,N_6439,N_6938);
and U7064 (N_7064,N_6233,N_6838);
or U7065 (N_7065,N_6282,N_6972);
nand U7066 (N_7066,N_6367,N_6732);
and U7067 (N_7067,N_6169,N_6802);
and U7068 (N_7068,N_6555,N_6927);
nand U7069 (N_7069,N_6279,N_6962);
or U7070 (N_7070,N_6628,N_6341);
xor U7071 (N_7071,N_6046,N_6966);
xor U7072 (N_7072,N_6027,N_6584);
or U7073 (N_7073,N_6623,N_6479);
and U7074 (N_7074,N_6534,N_6891);
xnor U7075 (N_7075,N_6089,N_6564);
and U7076 (N_7076,N_6284,N_6204);
or U7077 (N_7077,N_6184,N_6030);
and U7078 (N_7078,N_6971,N_6020);
nor U7079 (N_7079,N_6230,N_6394);
or U7080 (N_7080,N_6174,N_6182);
and U7081 (N_7081,N_6892,N_6978);
nor U7082 (N_7082,N_6669,N_6385);
and U7083 (N_7083,N_6822,N_6129);
or U7084 (N_7084,N_6657,N_6916);
nand U7085 (N_7085,N_6464,N_6750);
and U7086 (N_7086,N_6435,N_6031);
xnor U7087 (N_7087,N_6227,N_6480);
nand U7088 (N_7088,N_6316,N_6467);
nor U7089 (N_7089,N_6761,N_6654);
xnor U7090 (N_7090,N_6566,N_6088);
nand U7091 (N_7091,N_6984,N_6446);
or U7092 (N_7092,N_6197,N_6701);
or U7093 (N_7093,N_6980,N_6324);
nor U7094 (N_7094,N_6721,N_6516);
nor U7095 (N_7095,N_6484,N_6693);
nor U7096 (N_7096,N_6487,N_6619);
xnor U7097 (N_7097,N_6453,N_6071);
nor U7098 (N_7098,N_6413,N_6263);
nand U7099 (N_7099,N_6570,N_6678);
nand U7100 (N_7100,N_6225,N_6683);
and U7101 (N_7101,N_6821,N_6719);
nor U7102 (N_7102,N_6731,N_6825);
nand U7103 (N_7103,N_6106,N_6662);
nor U7104 (N_7104,N_6589,N_6189);
nor U7105 (N_7105,N_6244,N_6800);
and U7106 (N_7106,N_6999,N_6608);
nand U7107 (N_7107,N_6058,N_6094);
nand U7108 (N_7108,N_6616,N_6000);
or U7109 (N_7109,N_6164,N_6458);
or U7110 (N_7110,N_6786,N_6486);
nor U7111 (N_7111,N_6820,N_6343);
nor U7112 (N_7112,N_6315,N_6499);
nor U7113 (N_7113,N_6539,N_6354);
or U7114 (N_7114,N_6939,N_6271);
nand U7115 (N_7115,N_6943,N_6845);
and U7116 (N_7116,N_6494,N_6777);
and U7117 (N_7117,N_6157,N_6102);
nor U7118 (N_7118,N_6801,N_6796);
or U7119 (N_7119,N_6173,N_6124);
and U7120 (N_7120,N_6056,N_6298);
nand U7121 (N_7121,N_6743,N_6773);
or U7122 (N_7122,N_6523,N_6833);
or U7123 (N_7123,N_6493,N_6620);
nand U7124 (N_7124,N_6625,N_6449);
or U7125 (N_7125,N_6161,N_6744);
and U7126 (N_7126,N_6188,N_6596);
or U7127 (N_7127,N_6255,N_6793);
nor U7128 (N_7128,N_6065,N_6374);
nand U7129 (N_7129,N_6880,N_6126);
xor U7130 (N_7130,N_6288,N_6763);
or U7131 (N_7131,N_6725,N_6913);
nor U7132 (N_7132,N_6809,N_6167);
and U7133 (N_7133,N_6485,N_6261);
and U7134 (N_7134,N_6658,N_6336);
or U7135 (N_7135,N_6959,N_6930);
nand U7136 (N_7136,N_6420,N_6736);
or U7137 (N_7137,N_6746,N_6470);
or U7138 (N_7138,N_6741,N_6010);
nand U7139 (N_7139,N_6593,N_6390);
nand U7140 (N_7140,N_6112,N_6517);
or U7141 (N_7141,N_6185,N_6951);
or U7142 (N_7142,N_6314,N_6070);
and U7143 (N_7143,N_6468,N_6080);
and U7144 (N_7144,N_6195,N_6996);
and U7145 (N_7145,N_6242,N_6005);
or U7146 (N_7146,N_6007,N_6856);
and U7147 (N_7147,N_6785,N_6695);
and U7148 (N_7148,N_6257,N_6154);
and U7149 (N_7149,N_6462,N_6273);
or U7150 (N_7150,N_6116,N_6923);
xnor U7151 (N_7151,N_6813,N_6024);
nand U7152 (N_7152,N_6482,N_6788);
nand U7153 (N_7153,N_6630,N_6934);
and U7154 (N_7154,N_6015,N_6521);
nor U7155 (N_7155,N_6053,N_6200);
nand U7156 (N_7156,N_6091,N_6310);
or U7157 (N_7157,N_6819,N_6047);
and U7158 (N_7158,N_6063,N_6952);
nor U7159 (N_7159,N_6723,N_6395);
and U7160 (N_7160,N_6098,N_6670);
nand U7161 (N_7161,N_6844,N_6403);
or U7162 (N_7162,N_6776,N_6835);
and U7163 (N_7163,N_6665,N_6624);
nor U7164 (N_7164,N_6375,N_6382);
nor U7165 (N_7165,N_6532,N_6568);
nand U7166 (N_7166,N_6211,N_6626);
and U7167 (N_7167,N_6588,N_6912);
or U7168 (N_7168,N_6292,N_6210);
or U7169 (N_7169,N_6594,N_6095);
nand U7170 (N_7170,N_6442,N_6950);
or U7171 (N_7171,N_6293,N_6426);
and U7172 (N_7172,N_6947,N_6510);
nor U7173 (N_7173,N_6803,N_6176);
nor U7174 (N_7174,N_6705,N_6334);
or U7175 (N_7175,N_6371,N_6082);
and U7176 (N_7176,N_6910,N_6143);
or U7177 (N_7177,N_6032,N_6974);
or U7178 (N_7178,N_6636,N_6659);
or U7179 (N_7179,N_6365,N_6524);
nand U7180 (N_7180,N_6113,N_6149);
nand U7181 (N_7181,N_6536,N_6708);
nor U7182 (N_7182,N_6084,N_6740);
or U7183 (N_7183,N_6514,N_6025);
nand U7184 (N_7184,N_6881,N_6006);
or U7185 (N_7185,N_6383,N_6151);
nor U7186 (N_7186,N_6476,N_6787);
nand U7187 (N_7187,N_6198,N_6792);
nand U7188 (N_7188,N_6882,N_6232);
or U7189 (N_7189,N_6944,N_6407);
and U7190 (N_7190,N_6790,N_6663);
xor U7191 (N_7191,N_6223,N_6868);
nand U7192 (N_7192,N_6421,N_6915);
nor U7193 (N_7193,N_6737,N_6783);
and U7194 (N_7194,N_6937,N_6515);
nor U7195 (N_7195,N_6504,N_6520);
nor U7196 (N_7196,N_6533,N_6827);
xnor U7197 (N_7197,N_6765,N_6226);
nand U7198 (N_7198,N_6357,N_6858);
nand U7199 (N_7199,N_6672,N_6638);
nor U7200 (N_7200,N_6306,N_6175);
or U7201 (N_7201,N_6068,N_6526);
xor U7202 (N_7202,N_6631,N_6496);
or U7203 (N_7203,N_6976,N_6460);
and U7204 (N_7204,N_6400,N_6501);
or U7205 (N_7205,N_6933,N_6576);
nand U7206 (N_7206,N_6142,N_6222);
nand U7207 (N_7207,N_6190,N_6445);
and U7208 (N_7208,N_6935,N_6239);
and U7209 (N_7209,N_6878,N_6477);
or U7210 (N_7210,N_6307,N_6795);
nor U7211 (N_7211,N_6926,N_6141);
or U7212 (N_7212,N_6183,N_6396);
xor U7213 (N_7213,N_6208,N_6262);
nand U7214 (N_7214,N_6187,N_6440);
nor U7215 (N_7215,N_6558,N_6556);
or U7216 (N_7216,N_6302,N_6869);
or U7217 (N_7217,N_6617,N_6377);
xnor U7218 (N_7218,N_6337,N_6807);
nand U7219 (N_7219,N_6340,N_6351);
xor U7220 (N_7220,N_6437,N_6872);
nand U7221 (N_7221,N_6804,N_6922);
and U7222 (N_7222,N_6691,N_6252);
xor U7223 (N_7223,N_6834,N_6717);
and U7224 (N_7224,N_6729,N_6320);
nand U7225 (N_7225,N_6072,N_6455);
nand U7226 (N_7226,N_6682,N_6945);
or U7227 (N_7227,N_6964,N_6987);
or U7228 (N_7228,N_6685,N_6756);
nand U7229 (N_7229,N_6864,N_6212);
nor U7230 (N_7230,N_6410,N_6170);
nor U7231 (N_7231,N_6846,N_6893);
nand U7232 (N_7232,N_6018,N_6137);
nor U7233 (N_7233,N_6270,N_6364);
or U7234 (N_7234,N_6724,N_6461);
and U7235 (N_7235,N_6205,N_6522);
nor U7236 (N_7236,N_6917,N_6794);
nand U7237 (N_7237,N_6327,N_6452);
and U7238 (N_7238,N_6247,N_6414);
xor U7239 (N_7239,N_6412,N_6599);
xor U7240 (N_7240,N_6041,N_6117);
and U7241 (N_7241,N_6901,N_6530);
and U7242 (N_7242,N_6931,N_6561);
or U7243 (N_7243,N_6733,N_6552);
or U7244 (N_7244,N_6574,N_6254);
nor U7245 (N_7245,N_6076,N_6299);
nand U7246 (N_7246,N_6936,N_6335);
xor U7247 (N_7247,N_6311,N_6378);
xor U7248 (N_7248,N_6349,N_6851);
nor U7249 (N_7249,N_6042,N_6598);
nand U7250 (N_7250,N_6229,N_6652);
or U7251 (N_7251,N_6512,N_6988);
nand U7252 (N_7252,N_6213,N_6637);
and U7253 (N_7253,N_6304,N_6266);
nor U7254 (N_7254,N_6862,N_6043);
nor U7255 (N_7255,N_6591,N_6519);
nor U7256 (N_7256,N_6465,N_6399);
nor U7257 (N_7257,N_6285,N_6345);
and U7258 (N_7258,N_6518,N_6034);
or U7259 (N_7259,N_6528,N_6860);
and U7260 (N_7260,N_6728,N_6768);
nor U7261 (N_7261,N_6406,N_6352);
or U7262 (N_7262,N_6152,N_6199);
and U7263 (N_7263,N_6960,N_6755);
nand U7264 (N_7264,N_6873,N_6722);
nand U7265 (N_7265,N_6680,N_6323);
and U7266 (N_7266,N_6703,N_6907);
or U7267 (N_7267,N_6267,N_6961);
or U7268 (N_7268,N_6333,N_6438);
nor U7269 (N_7269,N_6416,N_6321);
and U7270 (N_7270,N_6604,N_6287);
and U7271 (N_7271,N_6739,N_6754);
nor U7272 (N_7272,N_6497,N_6602);
and U7273 (N_7273,N_6876,N_6954);
nand U7274 (N_7274,N_6920,N_6535);
or U7275 (N_7275,N_6769,N_6673);
and U7276 (N_7276,N_6138,N_6104);
and U7277 (N_7277,N_6035,N_6286);
or U7278 (N_7278,N_6193,N_6432);
or U7279 (N_7279,N_6474,N_6055);
nand U7280 (N_7280,N_6128,N_6767);
and U7281 (N_7281,N_6051,N_6331);
nor U7282 (N_7282,N_6894,N_6671);
and U7283 (N_7283,N_6778,N_6150);
nand U7284 (N_7284,N_6289,N_6186);
xnor U7285 (N_7285,N_6348,N_6234);
nor U7286 (N_7286,N_6013,N_6565);
nor U7287 (N_7287,N_6906,N_6645);
and U7288 (N_7288,N_6159,N_6411);
nor U7289 (N_7289,N_6774,N_6726);
and U7290 (N_7290,N_6201,N_6361);
nand U7291 (N_7291,N_6344,N_6489);
nand U7292 (N_7292,N_6009,N_6103);
and U7293 (N_7293,N_6118,N_6902);
nand U7294 (N_7294,N_6029,N_6646);
or U7295 (N_7295,N_6326,N_6979);
nor U7296 (N_7296,N_6269,N_6481);
nor U7297 (N_7297,N_6206,N_6023);
and U7298 (N_7298,N_6597,N_6587);
and U7299 (N_7299,N_6238,N_6008);
and U7300 (N_7300,N_6220,N_6471);
and U7301 (N_7301,N_6814,N_6393);
or U7302 (N_7302,N_6674,N_6240);
or U7303 (N_7303,N_6661,N_6218);
xor U7304 (N_7304,N_6405,N_6318);
or U7305 (N_7305,N_6779,N_6148);
nand U7306 (N_7306,N_6537,N_6264);
or U7307 (N_7307,N_6248,N_6981);
xor U7308 (N_7308,N_6949,N_6649);
or U7309 (N_7309,N_6014,N_6918);
nand U7310 (N_7310,N_6702,N_6970);
and U7311 (N_7311,N_6849,N_6380);
nand U7312 (N_7312,N_6162,N_6109);
nor U7313 (N_7313,N_6752,N_6694);
or U7314 (N_7314,N_6870,N_6260);
or U7315 (N_7315,N_6581,N_6123);
or U7316 (N_7316,N_6635,N_6855);
and U7317 (N_7317,N_6506,N_6977);
or U7318 (N_7318,N_6559,N_6045);
nand U7319 (N_7319,N_6824,N_6823);
nor U7320 (N_7320,N_6276,N_6011);
xnor U7321 (N_7321,N_6120,N_6235);
nor U7322 (N_7322,N_6425,N_6245);
and U7323 (N_7323,N_6134,N_6742);
xnor U7324 (N_7324,N_6956,N_6308);
or U7325 (N_7325,N_6560,N_6990);
nand U7326 (N_7326,N_6953,N_6679);
nor U7327 (N_7327,N_6829,N_6171);
nor U7328 (N_7328,N_6582,N_6610);
nand U7329 (N_7329,N_6300,N_6643);
and U7330 (N_7330,N_6451,N_6840);
nand U7331 (N_7331,N_6590,N_6651);
and U7332 (N_7332,N_6711,N_6727);
nand U7333 (N_7333,N_6301,N_6178);
nand U7334 (N_7334,N_6650,N_6492);
and U7335 (N_7335,N_6221,N_6710);
or U7336 (N_7336,N_6441,N_6139);
nor U7337 (N_7337,N_6066,N_6177);
nor U7338 (N_7338,N_6402,N_6090);
and U7339 (N_7339,N_6629,N_6319);
xor U7340 (N_7340,N_6549,N_6360);
and U7341 (N_7341,N_6667,N_6111);
xnor U7342 (N_7342,N_6309,N_6914);
nor U7343 (N_7343,N_6339,N_6692);
or U7344 (N_7344,N_6359,N_6982);
nor U7345 (N_7345,N_6274,N_6601);
nand U7346 (N_7346,N_6275,N_6356);
xnor U7347 (N_7347,N_6888,N_6033);
nand U7348 (N_7348,N_6817,N_6022);
or U7349 (N_7349,N_6083,N_6122);
nor U7350 (N_7350,N_6202,N_6969);
or U7351 (N_7351,N_6745,N_6563);
or U7352 (N_7352,N_6115,N_6236);
nand U7353 (N_7353,N_6527,N_6965);
nor U7354 (N_7354,N_6553,N_6338);
or U7355 (N_7355,N_6277,N_6747);
nor U7356 (N_7356,N_6885,N_6697);
and U7357 (N_7357,N_6583,N_6166);
xor U7358 (N_7358,N_6054,N_6831);
nand U7359 (N_7359,N_6329,N_6686);
nand U7360 (N_7360,N_6463,N_6886);
or U7361 (N_7361,N_6272,N_6075);
or U7362 (N_7362,N_6125,N_6758);
nand U7363 (N_7363,N_6508,N_6551);
nor U7364 (N_7364,N_6797,N_6368);
and U7365 (N_7365,N_6436,N_6478);
or U7366 (N_7366,N_6567,N_6017);
or U7367 (N_7367,N_6294,N_6618);
nand U7368 (N_7368,N_6995,N_6069);
or U7369 (N_7369,N_6409,N_6259);
or U7370 (N_7370,N_6044,N_6085);
nand U7371 (N_7371,N_6607,N_6542);
or U7372 (N_7372,N_6350,N_6156);
nor U7373 (N_7373,N_6214,N_6019);
or U7374 (N_7374,N_6155,N_6993);
nand U7375 (N_7375,N_6709,N_6086);
nor U7376 (N_7376,N_6789,N_6268);
nor U7377 (N_7377,N_6147,N_6196);
and U7378 (N_7378,N_6606,N_6799);
nand U7379 (N_7379,N_6430,N_6466);
and U7380 (N_7380,N_6433,N_6699);
or U7381 (N_7381,N_6062,N_6498);
nand U7382 (N_7382,N_6757,N_6941);
nor U7383 (N_7383,N_6905,N_6771);
nand U7384 (N_7384,N_6016,N_6550);
or U7385 (N_7385,N_6592,N_6548);
or U7386 (N_7386,N_6780,N_6940);
xor U7387 (N_7387,N_6454,N_6073);
nand U7388 (N_7388,N_6850,N_6052);
xor U7389 (N_7389,N_6642,N_6791);
and U7390 (N_7390,N_6388,N_6146);
nor U7391 (N_7391,N_6163,N_6280);
nor U7392 (N_7392,N_6782,N_6716);
and U7393 (N_7393,N_6718,N_6753);
nor U7394 (N_7394,N_6540,N_6495);
and U7395 (N_7395,N_6093,N_6422);
xor U7396 (N_7396,N_6975,N_6621);
nor U7397 (N_7397,N_6854,N_6491);
nand U7398 (N_7398,N_6107,N_6770);
and U7399 (N_7399,N_6097,N_6417);
and U7400 (N_7400,N_6419,N_6573);
nand U7401 (N_7401,N_6291,N_6775);
and U7402 (N_7402,N_6473,N_6110);
xor U7403 (N_7403,N_6140,N_6666);
and U7404 (N_7404,N_6037,N_6919);
nor U7405 (N_7405,N_6644,N_6810);
nor U7406 (N_7406,N_6689,N_6525);
or U7407 (N_7407,N_6048,N_6655);
nand U7408 (N_7408,N_6908,N_6544);
or U7409 (N_7409,N_6541,N_6812);
xor U7410 (N_7410,N_6571,N_6612);
nand U7411 (N_7411,N_6503,N_6192);
nand U7412 (N_7412,N_6179,N_6330);
or U7413 (N_7413,N_6759,N_6611);
or U7414 (N_7414,N_6057,N_6676);
nand U7415 (N_7415,N_6967,N_6687);
or U7416 (N_7416,N_6224,N_6397);
nor U7417 (N_7417,N_6562,N_6165);
or U7418 (N_7418,N_6366,N_6502);
or U7419 (N_7419,N_6720,N_6735);
nand U7420 (N_7420,N_6688,N_6632);
and U7421 (N_7421,N_6296,N_6890);
nor U7422 (N_7422,N_6418,N_6713);
or U7423 (N_7423,N_6038,N_6781);
nand U7424 (N_7424,N_6595,N_6459);
nand U7425 (N_7425,N_6099,N_6448);
nor U7426 (N_7426,N_6404,N_6973);
nor U7427 (N_7427,N_6281,N_6246);
and U7428 (N_7428,N_6911,N_6579);
or U7429 (N_7429,N_6215,N_6191);
nand U7430 (N_7430,N_6963,N_6609);
nor U7431 (N_7431,N_6871,N_6836);
nor U7432 (N_7432,N_6207,N_6067);
or U7433 (N_7433,N_6538,N_6325);
or U7434 (N_7434,N_6889,N_6386);
or U7435 (N_7435,N_6605,N_6092);
nand U7436 (N_7436,N_6332,N_6194);
nor U7437 (N_7437,N_6751,N_6859);
nand U7438 (N_7438,N_6968,N_6766);
nor U7439 (N_7439,N_6575,N_6434);
or U7440 (N_7440,N_6698,N_6681);
nand U7441 (N_7441,N_6505,N_6243);
and U7442 (N_7442,N_6660,N_6656);
and U7443 (N_7443,N_6132,N_6852);
nand U7444 (N_7444,N_6640,N_6295);
nand U7445 (N_7445,N_6877,N_6003);
nor U7446 (N_7446,N_6429,N_6715);
xnor U7447 (N_7447,N_6806,N_6986);
xor U7448 (N_7448,N_6472,N_6760);
and U7449 (N_7449,N_6841,N_6529);
or U7450 (N_7450,N_6237,N_6955);
and U7451 (N_7451,N_6369,N_6077);
nor U7452 (N_7452,N_6647,N_6028);
or U7453 (N_7453,N_6957,N_6153);
and U7454 (N_7454,N_6839,N_6249);
nand U7455 (N_7455,N_6633,N_6059);
and U7456 (N_7456,N_6899,N_6362);
nor U7457 (N_7457,N_6896,N_6847);
and U7458 (N_7458,N_6843,N_6347);
or U7459 (N_7459,N_6398,N_6585);
nor U7460 (N_7460,N_6543,N_6690);
or U7461 (N_7461,N_6507,N_6303);
or U7462 (N_7462,N_6290,N_6250);
xnor U7463 (N_7463,N_6228,N_6707);
or U7464 (N_7464,N_6021,N_6358);
nand U7465 (N_7465,N_6738,N_6081);
and U7466 (N_7466,N_6490,N_6145);
nor U7467 (N_7467,N_6180,N_6511);
or U7468 (N_7468,N_6241,N_6614);
and U7469 (N_7469,N_6985,N_6904);
nor U7470 (N_7470,N_6653,N_6130);
xnor U7471 (N_7471,N_6531,N_6346);
nor U7472 (N_7472,N_6312,N_6415);
xor U7473 (N_7473,N_6712,N_6762);
or U7474 (N_7474,N_6313,N_6160);
or U7475 (N_7475,N_6866,N_6004);
or U7476 (N_7476,N_6297,N_6928);
nor U7477 (N_7477,N_6879,N_6875);
nor U7478 (N_7478,N_6675,N_6172);
nand U7479 (N_7479,N_6026,N_6469);
and U7480 (N_7480,N_6387,N_6991);
or U7481 (N_7481,N_6546,N_6603);
xor U7482 (N_7482,N_6925,N_6131);
or U7483 (N_7483,N_6408,N_6897);
nand U7484 (N_7484,N_6353,N_6392);
and U7485 (N_7485,N_6251,N_6135);
nand U7486 (N_7486,N_6376,N_6079);
xnor U7487 (N_7487,N_6001,N_6060);
nor U7488 (N_7488,N_6815,N_6278);
nor U7489 (N_7489,N_6509,N_6648);
or U7490 (N_7490,N_6958,N_6209);
or U7491 (N_7491,N_6061,N_6554);
or U7492 (N_7492,N_6401,N_6253);
and U7493 (N_7493,N_6903,N_6994);
xor U7494 (N_7494,N_6216,N_6706);
xnor U7495 (N_7495,N_6355,N_6483);
or U7496 (N_7496,N_6475,N_6867);
and U7497 (N_7497,N_6087,N_6600);
nor U7498 (N_7498,N_6444,N_6929);
nor U7499 (N_7499,N_6317,N_6784);
nand U7500 (N_7500,N_6416,N_6463);
nor U7501 (N_7501,N_6663,N_6050);
xor U7502 (N_7502,N_6602,N_6422);
nor U7503 (N_7503,N_6670,N_6277);
xor U7504 (N_7504,N_6662,N_6356);
nor U7505 (N_7505,N_6599,N_6418);
or U7506 (N_7506,N_6288,N_6429);
xor U7507 (N_7507,N_6419,N_6695);
and U7508 (N_7508,N_6626,N_6708);
or U7509 (N_7509,N_6860,N_6246);
and U7510 (N_7510,N_6735,N_6240);
nor U7511 (N_7511,N_6092,N_6735);
nor U7512 (N_7512,N_6564,N_6202);
xnor U7513 (N_7513,N_6988,N_6671);
nor U7514 (N_7514,N_6606,N_6270);
and U7515 (N_7515,N_6300,N_6620);
nand U7516 (N_7516,N_6205,N_6843);
nor U7517 (N_7517,N_6988,N_6778);
nor U7518 (N_7518,N_6518,N_6724);
xnor U7519 (N_7519,N_6064,N_6939);
or U7520 (N_7520,N_6445,N_6129);
xnor U7521 (N_7521,N_6390,N_6582);
or U7522 (N_7522,N_6019,N_6836);
or U7523 (N_7523,N_6271,N_6772);
and U7524 (N_7524,N_6969,N_6663);
nor U7525 (N_7525,N_6894,N_6938);
or U7526 (N_7526,N_6266,N_6797);
nand U7527 (N_7527,N_6086,N_6507);
or U7528 (N_7528,N_6515,N_6116);
xnor U7529 (N_7529,N_6041,N_6148);
and U7530 (N_7530,N_6260,N_6847);
and U7531 (N_7531,N_6522,N_6690);
nand U7532 (N_7532,N_6853,N_6887);
xor U7533 (N_7533,N_6622,N_6142);
nand U7534 (N_7534,N_6538,N_6529);
xor U7535 (N_7535,N_6518,N_6621);
nand U7536 (N_7536,N_6926,N_6165);
nor U7537 (N_7537,N_6995,N_6112);
nand U7538 (N_7538,N_6651,N_6125);
and U7539 (N_7539,N_6267,N_6168);
and U7540 (N_7540,N_6222,N_6414);
nor U7541 (N_7541,N_6809,N_6094);
nor U7542 (N_7542,N_6539,N_6467);
or U7543 (N_7543,N_6897,N_6881);
and U7544 (N_7544,N_6699,N_6244);
or U7545 (N_7545,N_6293,N_6918);
nor U7546 (N_7546,N_6738,N_6863);
nor U7547 (N_7547,N_6637,N_6765);
or U7548 (N_7548,N_6162,N_6383);
nor U7549 (N_7549,N_6864,N_6843);
and U7550 (N_7550,N_6002,N_6387);
and U7551 (N_7551,N_6599,N_6382);
xnor U7552 (N_7552,N_6507,N_6349);
or U7553 (N_7553,N_6932,N_6268);
or U7554 (N_7554,N_6861,N_6033);
and U7555 (N_7555,N_6293,N_6356);
and U7556 (N_7556,N_6613,N_6459);
nand U7557 (N_7557,N_6749,N_6199);
xnor U7558 (N_7558,N_6464,N_6508);
nand U7559 (N_7559,N_6502,N_6032);
nor U7560 (N_7560,N_6449,N_6143);
or U7561 (N_7561,N_6688,N_6208);
or U7562 (N_7562,N_6444,N_6900);
nor U7563 (N_7563,N_6810,N_6876);
nor U7564 (N_7564,N_6596,N_6637);
and U7565 (N_7565,N_6079,N_6873);
and U7566 (N_7566,N_6821,N_6012);
and U7567 (N_7567,N_6964,N_6962);
nand U7568 (N_7568,N_6597,N_6058);
xnor U7569 (N_7569,N_6824,N_6932);
or U7570 (N_7570,N_6088,N_6214);
nand U7571 (N_7571,N_6848,N_6109);
or U7572 (N_7572,N_6480,N_6070);
and U7573 (N_7573,N_6982,N_6203);
or U7574 (N_7574,N_6502,N_6293);
and U7575 (N_7575,N_6451,N_6025);
and U7576 (N_7576,N_6779,N_6585);
and U7577 (N_7577,N_6254,N_6899);
and U7578 (N_7578,N_6816,N_6474);
nand U7579 (N_7579,N_6700,N_6154);
nand U7580 (N_7580,N_6400,N_6086);
nand U7581 (N_7581,N_6990,N_6330);
and U7582 (N_7582,N_6019,N_6180);
or U7583 (N_7583,N_6845,N_6955);
and U7584 (N_7584,N_6851,N_6622);
nor U7585 (N_7585,N_6749,N_6830);
and U7586 (N_7586,N_6900,N_6142);
nor U7587 (N_7587,N_6461,N_6163);
and U7588 (N_7588,N_6142,N_6228);
or U7589 (N_7589,N_6350,N_6499);
nor U7590 (N_7590,N_6532,N_6569);
nor U7591 (N_7591,N_6809,N_6108);
nand U7592 (N_7592,N_6156,N_6690);
nand U7593 (N_7593,N_6919,N_6971);
nand U7594 (N_7594,N_6792,N_6651);
nand U7595 (N_7595,N_6448,N_6102);
and U7596 (N_7596,N_6948,N_6182);
nand U7597 (N_7597,N_6601,N_6697);
and U7598 (N_7598,N_6626,N_6786);
nand U7599 (N_7599,N_6357,N_6440);
nor U7600 (N_7600,N_6176,N_6380);
or U7601 (N_7601,N_6835,N_6389);
nand U7602 (N_7602,N_6409,N_6370);
and U7603 (N_7603,N_6811,N_6528);
nor U7604 (N_7604,N_6739,N_6424);
nand U7605 (N_7605,N_6146,N_6957);
and U7606 (N_7606,N_6598,N_6187);
xnor U7607 (N_7607,N_6613,N_6289);
nand U7608 (N_7608,N_6862,N_6202);
and U7609 (N_7609,N_6240,N_6419);
or U7610 (N_7610,N_6378,N_6356);
nand U7611 (N_7611,N_6570,N_6608);
xnor U7612 (N_7612,N_6734,N_6712);
xnor U7613 (N_7613,N_6807,N_6795);
xor U7614 (N_7614,N_6496,N_6603);
nand U7615 (N_7615,N_6080,N_6379);
nand U7616 (N_7616,N_6452,N_6696);
and U7617 (N_7617,N_6819,N_6084);
nor U7618 (N_7618,N_6888,N_6017);
and U7619 (N_7619,N_6572,N_6085);
nand U7620 (N_7620,N_6789,N_6798);
nor U7621 (N_7621,N_6323,N_6393);
nor U7622 (N_7622,N_6651,N_6360);
nand U7623 (N_7623,N_6806,N_6667);
or U7624 (N_7624,N_6280,N_6830);
nand U7625 (N_7625,N_6843,N_6665);
nand U7626 (N_7626,N_6534,N_6014);
nor U7627 (N_7627,N_6843,N_6417);
nor U7628 (N_7628,N_6498,N_6544);
nor U7629 (N_7629,N_6709,N_6881);
xnor U7630 (N_7630,N_6634,N_6027);
or U7631 (N_7631,N_6971,N_6406);
and U7632 (N_7632,N_6460,N_6479);
nand U7633 (N_7633,N_6043,N_6680);
or U7634 (N_7634,N_6020,N_6751);
nor U7635 (N_7635,N_6209,N_6014);
nor U7636 (N_7636,N_6479,N_6018);
nor U7637 (N_7637,N_6437,N_6736);
and U7638 (N_7638,N_6578,N_6412);
and U7639 (N_7639,N_6631,N_6088);
or U7640 (N_7640,N_6041,N_6675);
nor U7641 (N_7641,N_6406,N_6404);
nand U7642 (N_7642,N_6017,N_6659);
nor U7643 (N_7643,N_6856,N_6107);
or U7644 (N_7644,N_6089,N_6005);
and U7645 (N_7645,N_6300,N_6770);
nor U7646 (N_7646,N_6863,N_6974);
nor U7647 (N_7647,N_6560,N_6904);
or U7648 (N_7648,N_6627,N_6519);
or U7649 (N_7649,N_6373,N_6714);
nor U7650 (N_7650,N_6605,N_6685);
and U7651 (N_7651,N_6393,N_6885);
and U7652 (N_7652,N_6073,N_6263);
nand U7653 (N_7653,N_6159,N_6757);
nand U7654 (N_7654,N_6960,N_6243);
nor U7655 (N_7655,N_6902,N_6036);
nand U7656 (N_7656,N_6388,N_6826);
nand U7657 (N_7657,N_6879,N_6970);
and U7658 (N_7658,N_6224,N_6038);
nor U7659 (N_7659,N_6443,N_6073);
xnor U7660 (N_7660,N_6564,N_6741);
nand U7661 (N_7661,N_6326,N_6901);
nand U7662 (N_7662,N_6683,N_6602);
and U7663 (N_7663,N_6796,N_6541);
xor U7664 (N_7664,N_6389,N_6368);
nor U7665 (N_7665,N_6533,N_6627);
or U7666 (N_7666,N_6943,N_6644);
and U7667 (N_7667,N_6758,N_6450);
and U7668 (N_7668,N_6025,N_6216);
xor U7669 (N_7669,N_6085,N_6959);
and U7670 (N_7670,N_6263,N_6381);
nand U7671 (N_7671,N_6238,N_6807);
nand U7672 (N_7672,N_6042,N_6173);
and U7673 (N_7673,N_6125,N_6845);
nor U7674 (N_7674,N_6791,N_6306);
xnor U7675 (N_7675,N_6215,N_6711);
and U7676 (N_7676,N_6656,N_6779);
and U7677 (N_7677,N_6551,N_6504);
or U7678 (N_7678,N_6835,N_6430);
or U7679 (N_7679,N_6682,N_6666);
nor U7680 (N_7680,N_6411,N_6723);
nand U7681 (N_7681,N_6785,N_6027);
or U7682 (N_7682,N_6735,N_6398);
or U7683 (N_7683,N_6887,N_6695);
and U7684 (N_7684,N_6576,N_6480);
and U7685 (N_7685,N_6469,N_6011);
or U7686 (N_7686,N_6460,N_6306);
or U7687 (N_7687,N_6155,N_6056);
nand U7688 (N_7688,N_6767,N_6692);
nor U7689 (N_7689,N_6860,N_6723);
nor U7690 (N_7690,N_6983,N_6172);
nand U7691 (N_7691,N_6186,N_6894);
or U7692 (N_7692,N_6287,N_6179);
or U7693 (N_7693,N_6184,N_6721);
or U7694 (N_7694,N_6320,N_6978);
nor U7695 (N_7695,N_6898,N_6541);
and U7696 (N_7696,N_6093,N_6726);
and U7697 (N_7697,N_6871,N_6283);
and U7698 (N_7698,N_6214,N_6722);
nand U7699 (N_7699,N_6701,N_6531);
nand U7700 (N_7700,N_6111,N_6228);
xnor U7701 (N_7701,N_6757,N_6138);
nor U7702 (N_7702,N_6653,N_6358);
or U7703 (N_7703,N_6394,N_6739);
or U7704 (N_7704,N_6632,N_6156);
nand U7705 (N_7705,N_6837,N_6431);
xor U7706 (N_7706,N_6703,N_6111);
xnor U7707 (N_7707,N_6922,N_6164);
nor U7708 (N_7708,N_6201,N_6979);
and U7709 (N_7709,N_6453,N_6340);
xor U7710 (N_7710,N_6252,N_6036);
or U7711 (N_7711,N_6278,N_6748);
and U7712 (N_7712,N_6538,N_6223);
nand U7713 (N_7713,N_6950,N_6469);
nor U7714 (N_7714,N_6535,N_6309);
nor U7715 (N_7715,N_6255,N_6516);
or U7716 (N_7716,N_6196,N_6205);
nor U7717 (N_7717,N_6672,N_6629);
xnor U7718 (N_7718,N_6290,N_6147);
and U7719 (N_7719,N_6858,N_6720);
nand U7720 (N_7720,N_6342,N_6751);
and U7721 (N_7721,N_6815,N_6094);
or U7722 (N_7722,N_6774,N_6399);
xor U7723 (N_7723,N_6457,N_6635);
nor U7724 (N_7724,N_6426,N_6149);
nand U7725 (N_7725,N_6006,N_6721);
xor U7726 (N_7726,N_6793,N_6655);
nand U7727 (N_7727,N_6825,N_6172);
and U7728 (N_7728,N_6045,N_6330);
xor U7729 (N_7729,N_6988,N_6912);
nor U7730 (N_7730,N_6535,N_6151);
nand U7731 (N_7731,N_6192,N_6404);
or U7732 (N_7732,N_6845,N_6712);
nand U7733 (N_7733,N_6880,N_6198);
nor U7734 (N_7734,N_6373,N_6415);
nand U7735 (N_7735,N_6391,N_6077);
or U7736 (N_7736,N_6238,N_6614);
nand U7737 (N_7737,N_6949,N_6701);
and U7738 (N_7738,N_6908,N_6311);
nand U7739 (N_7739,N_6161,N_6484);
and U7740 (N_7740,N_6885,N_6637);
or U7741 (N_7741,N_6746,N_6507);
xnor U7742 (N_7742,N_6199,N_6278);
nand U7743 (N_7743,N_6552,N_6366);
and U7744 (N_7744,N_6212,N_6312);
or U7745 (N_7745,N_6568,N_6601);
and U7746 (N_7746,N_6859,N_6092);
nor U7747 (N_7747,N_6531,N_6761);
nor U7748 (N_7748,N_6949,N_6648);
or U7749 (N_7749,N_6328,N_6230);
and U7750 (N_7750,N_6846,N_6185);
or U7751 (N_7751,N_6875,N_6830);
and U7752 (N_7752,N_6158,N_6135);
nor U7753 (N_7753,N_6431,N_6800);
nor U7754 (N_7754,N_6577,N_6618);
or U7755 (N_7755,N_6127,N_6467);
nor U7756 (N_7756,N_6883,N_6623);
and U7757 (N_7757,N_6815,N_6595);
and U7758 (N_7758,N_6200,N_6667);
nand U7759 (N_7759,N_6590,N_6421);
or U7760 (N_7760,N_6739,N_6324);
or U7761 (N_7761,N_6400,N_6350);
or U7762 (N_7762,N_6952,N_6241);
nand U7763 (N_7763,N_6069,N_6697);
or U7764 (N_7764,N_6333,N_6310);
nand U7765 (N_7765,N_6878,N_6572);
or U7766 (N_7766,N_6833,N_6042);
or U7767 (N_7767,N_6005,N_6131);
or U7768 (N_7768,N_6325,N_6251);
and U7769 (N_7769,N_6551,N_6288);
xor U7770 (N_7770,N_6403,N_6762);
and U7771 (N_7771,N_6659,N_6858);
nor U7772 (N_7772,N_6560,N_6539);
and U7773 (N_7773,N_6535,N_6416);
nand U7774 (N_7774,N_6358,N_6105);
and U7775 (N_7775,N_6025,N_6317);
and U7776 (N_7776,N_6786,N_6394);
nor U7777 (N_7777,N_6538,N_6720);
nand U7778 (N_7778,N_6553,N_6256);
or U7779 (N_7779,N_6875,N_6092);
nand U7780 (N_7780,N_6171,N_6183);
and U7781 (N_7781,N_6884,N_6955);
nand U7782 (N_7782,N_6212,N_6284);
or U7783 (N_7783,N_6661,N_6700);
nand U7784 (N_7784,N_6052,N_6237);
or U7785 (N_7785,N_6226,N_6580);
and U7786 (N_7786,N_6991,N_6972);
nor U7787 (N_7787,N_6748,N_6103);
nor U7788 (N_7788,N_6156,N_6131);
and U7789 (N_7789,N_6491,N_6359);
xnor U7790 (N_7790,N_6550,N_6096);
or U7791 (N_7791,N_6503,N_6968);
and U7792 (N_7792,N_6989,N_6372);
nand U7793 (N_7793,N_6369,N_6496);
nor U7794 (N_7794,N_6715,N_6173);
or U7795 (N_7795,N_6533,N_6492);
or U7796 (N_7796,N_6517,N_6408);
nand U7797 (N_7797,N_6477,N_6651);
and U7798 (N_7798,N_6251,N_6267);
nand U7799 (N_7799,N_6949,N_6391);
and U7800 (N_7800,N_6342,N_6974);
nor U7801 (N_7801,N_6767,N_6733);
nand U7802 (N_7802,N_6226,N_6206);
nor U7803 (N_7803,N_6588,N_6834);
nor U7804 (N_7804,N_6389,N_6987);
and U7805 (N_7805,N_6929,N_6088);
nand U7806 (N_7806,N_6144,N_6864);
nand U7807 (N_7807,N_6423,N_6072);
or U7808 (N_7808,N_6133,N_6065);
or U7809 (N_7809,N_6143,N_6018);
and U7810 (N_7810,N_6741,N_6342);
nor U7811 (N_7811,N_6604,N_6779);
nand U7812 (N_7812,N_6620,N_6901);
or U7813 (N_7813,N_6600,N_6717);
xnor U7814 (N_7814,N_6390,N_6818);
nand U7815 (N_7815,N_6548,N_6878);
nor U7816 (N_7816,N_6044,N_6843);
nor U7817 (N_7817,N_6090,N_6305);
and U7818 (N_7818,N_6492,N_6578);
xnor U7819 (N_7819,N_6669,N_6328);
and U7820 (N_7820,N_6841,N_6506);
and U7821 (N_7821,N_6607,N_6141);
and U7822 (N_7822,N_6794,N_6658);
and U7823 (N_7823,N_6961,N_6426);
or U7824 (N_7824,N_6732,N_6202);
and U7825 (N_7825,N_6373,N_6734);
nor U7826 (N_7826,N_6730,N_6004);
nand U7827 (N_7827,N_6520,N_6181);
or U7828 (N_7828,N_6565,N_6842);
xnor U7829 (N_7829,N_6191,N_6888);
or U7830 (N_7830,N_6910,N_6385);
nor U7831 (N_7831,N_6147,N_6548);
nor U7832 (N_7832,N_6776,N_6815);
nor U7833 (N_7833,N_6740,N_6173);
nand U7834 (N_7834,N_6054,N_6771);
nor U7835 (N_7835,N_6653,N_6614);
and U7836 (N_7836,N_6506,N_6807);
nor U7837 (N_7837,N_6027,N_6560);
nor U7838 (N_7838,N_6734,N_6624);
and U7839 (N_7839,N_6665,N_6090);
nand U7840 (N_7840,N_6571,N_6379);
nor U7841 (N_7841,N_6280,N_6604);
or U7842 (N_7842,N_6225,N_6597);
nand U7843 (N_7843,N_6207,N_6910);
nand U7844 (N_7844,N_6305,N_6995);
and U7845 (N_7845,N_6009,N_6327);
and U7846 (N_7846,N_6442,N_6914);
or U7847 (N_7847,N_6344,N_6594);
and U7848 (N_7848,N_6026,N_6087);
and U7849 (N_7849,N_6355,N_6277);
nand U7850 (N_7850,N_6637,N_6389);
and U7851 (N_7851,N_6568,N_6998);
and U7852 (N_7852,N_6901,N_6892);
nor U7853 (N_7853,N_6520,N_6370);
nand U7854 (N_7854,N_6669,N_6707);
and U7855 (N_7855,N_6340,N_6820);
and U7856 (N_7856,N_6362,N_6934);
nor U7857 (N_7857,N_6054,N_6059);
and U7858 (N_7858,N_6008,N_6665);
xor U7859 (N_7859,N_6779,N_6780);
nand U7860 (N_7860,N_6568,N_6905);
or U7861 (N_7861,N_6796,N_6821);
nor U7862 (N_7862,N_6528,N_6144);
nand U7863 (N_7863,N_6354,N_6457);
and U7864 (N_7864,N_6336,N_6558);
nand U7865 (N_7865,N_6267,N_6643);
and U7866 (N_7866,N_6120,N_6276);
xnor U7867 (N_7867,N_6249,N_6309);
nand U7868 (N_7868,N_6364,N_6238);
xnor U7869 (N_7869,N_6289,N_6659);
or U7870 (N_7870,N_6119,N_6879);
and U7871 (N_7871,N_6047,N_6719);
nor U7872 (N_7872,N_6214,N_6883);
or U7873 (N_7873,N_6939,N_6040);
nor U7874 (N_7874,N_6563,N_6681);
nor U7875 (N_7875,N_6278,N_6783);
nand U7876 (N_7876,N_6169,N_6617);
nor U7877 (N_7877,N_6011,N_6804);
nand U7878 (N_7878,N_6877,N_6791);
or U7879 (N_7879,N_6795,N_6338);
or U7880 (N_7880,N_6771,N_6483);
nand U7881 (N_7881,N_6885,N_6600);
xnor U7882 (N_7882,N_6002,N_6684);
nor U7883 (N_7883,N_6089,N_6732);
or U7884 (N_7884,N_6300,N_6407);
and U7885 (N_7885,N_6522,N_6959);
and U7886 (N_7886,N_6280,N_6615);
nor U7887 (N_7887,N_6265,N_6832);
nand U7888 (N_7888,N_6960,N_6970);
nand U7889 (N_7889,N_6416,N_6053);
or U7890 (N_7890,N_6075,N_6666);
xor U7891 (N_7891,N_6316,N_6201);
xor U7892 (N_7892,N_6438,N_6145);
nor U7893 (N_7893,N_6707,N_6153);
nor U7894 (N_7894,N_6474,N_6289);
or U7895 (N_7895,N_6913,N_6746);
nor U7896 (N_7896,N_6979,N_6289);
and U7897 (N_7897,N_6365,N_6384);
and U7898 (N_7898,N_6043,N_6827);
and U7899 (N_7899,N_6093,N_6834);
and U7900 (N_7900,N_6567,N_6247);
nor U7901 (N_7901,N_6936,N_6749);
xnor U7902 (N_7902,N_6579,N_6763);
nand U7903 (N_7903,N_6832,N_6939);
or U7904 (N_7904,N_6579,N_6756);
and U7905 (N_7905,N_6817,N_6125);
and U7906 (N_7906,N_6797,N_6299);
and U7907 (N_7907,N_6359,N_6444);
or U7908 (N_7908,N_6274,N_6560);
nor U7909 (N_7909,N_6793,N_6555);
nor U7910 (N_7910,N_6722,N_6993);
or U7911 (N_7911,N_6105,N_6696);
nor U7912 (N_7912,N_6097,N_6473);
nand U7913 (N_7913,N_6568,N_6135);
nand U7914 (N_7914,N_6108,N_6691);
nand U7915 (N_7915,N_6352,N_6594);
nor U7916 (N_7916,N_6724,N_6007);
nand U7917 (N_7917,N_6365,N_6269);
nand U7918 (N_7918,N_6199,N_6463);
and U7919 (N_7919,N_6118,N_6855);
nor U7920 (N_7920,N_6327,N_6012);
nor U7921 (N_7921,N_6992,N_6929);
or U7922 (N_7922,N_6528,N_6593);
xnor U7923 (N_7923,N_6634,N_6434);
nor U7924 (N_7924,N_6714,N_6864);
and U7925 (N_7925,N_6020,N_6221);
nor U7926 (N_7926,N_6777,N_6890);
and U7927 (N_7927,N_6261,N_6598);
and U7928 (N_7928,N_6635,N_6243);
or U7929 (N_7929,N_6227,N_6181);
nand U7930 (N_7930,N_6586,N_6314);
xor U7931 (N_7931,N_6132,N_6423);
or U7932 (N_7932,N_6408,N_6822);
nand U7933 (N_7933,N_6786,N_6971);
xor U7934 (N_7934,N_6138,N_6430);
nand U7935 (N_7935,N_6642,N_6657);
and U7936 (N_7936,N_6145,N_6282);
nand U7937 (N_7937,N_6608,N_6631);
and U7938 (N_7938,N_6791,N_6454);
xor U7939 (N_7939,N_6960,N_6016);
nor U7940 (N_7940,N_6695,N_6319);
nand U7941 (N_7941,N_6936,N_6915);
or U7942 (N_7942,N_6933,N_6582);
nor U7943 (N_7943,N_6490,N_6203);
nand U7944 (N_7944,N_6347,N_6395);
or U7945 (N_7945,N_6110,N_6517);
xnor U7946 (N_7946,N_6931,N_6336);
nand U7947 (N_7947,N_6293,N_6814);
and U7948 (N_7948,N_6334,N_6246);
or U7949 (N_7949,N_6964,N_6275);
and U7950 (N_7950,N_6627,N_6355);
or U7951 (N_7951,N_6214,N_6734);
and U7952 (N_7952,N_6753,N_6907);
nand U7953 (N_7953,N_6762,N_6362);
or U7954 (N_7954,N_6132,N_6337);
and U7955 (N_7955,N_6461,N_6471);
nand U7956 (N_7956,N_6207,N_6811);
nand U7957 (N_7957,N_6226,N_6048);
xor U7958 (N_7958,N_6521,N_6108);
nor U7959 (N_7959,N_6903,N_6603);
or U7960 (N_7960,N_6758,N_6969);
or U7961 (N_7961,N_6643,N_6845);
nor U7962 (N_7962,N_6437,N_6270);
nor U7963 (N_7963,N_6574,N_6858);
nor U7964 (N_7964,N_6390,N_6774);
nor U7965 (N_7965,N_6000,N_6074);
xor U7966 (N_7966,N_6237,N_6952);
or U7967 (N_7967,N_6073,N_6709);
or U7968 (N_7968,N_6620,N_6766);
or U7969 (N_7969,N_6667,N_6465);
or U7970 (N_7970,N_6173,N_6893);
and U7971 (N_7971,N_6918,N_6921);
nand U7972 (N_7972,N_6471,N_6858);
nor U7973 (N_7973,N_6515,N_6015);
nor U7974 (N_7974,N_6117,N_6957);
nand U7975 (N_7975,N_6711,N_6786);
nand U7976 (N_7976,N_6714,N_6994);
and U7977 (N_7977,N_6523,N_6126);
nand U7978 (N_7978,N_6544,N_6576);
nor U7979 (N_7979,N_6825,N_6209);
and U7980 (N_7980,N_6237,N_6441);
xnor U7981 (N_7981,N_6803,N_6482);
or U7982 (N_7982,N_6673,N_6236);
nand U7983 (N_7983,N_6799,N_6675);
xor U7984 (N_7984,N_6915,N_6393);
nand U7985 (N_7985,N_6748,N_6159);
nand U7986 (N_7986,N_6070,N_6045);
or U7987 (N_7987,N_6585,N_6595);
and U7988 (N_7988,N_6102,N_6894);
or U7989 (N_7989,N_6501,N_6917);
nor U7990 (N_7990,N_6788,N_6269);
nor U7991 (N_7991,N_6783,N_6594);
nor U7992 (N_7992,N_6751,N_6645);
xnor U7993 (N_7993,N_6489,N_6582);
xor U7994 (N_7994,N_6047,N_6200);
and U7995 (N_7995,N_6905,N_6526);
or U7996 (N_7996,N_6868,N_6543);
or U7997 (N_7997,N_6886,N_6087);
nand U7998 (N_7998,N_6794,N_6137);
nand U7999 (N_7999,N_6254,N_6867);
and U8000 (N_8000,N_7744,N_7332);
or U8001 (N_8001,N_7128,N_7064);
and U8002 (N_8002,N_7366,N_7132);
and U8003 (N_8003,N_7328,N_7330);
or U8004 (N_8004,N_7071,N_7404);
nor U8005 (N_8005,N_7793,N_7612);
and U8006 (N_8006,N_7705,N_7577);
nor U8007 (N_8007,N_7698,N_7928);
or U8008 (N_8008,N_7658,N_7760);
and U8009 (N_8009,N_7509,N_7798);
or U8010 (N_8010,N_7822,N_7037);
or U8011 (N_8011,N_7893,N_7180);
nor U8012 (N_8012,N_7364,N_7283);
nor U8013 (N_8013,N_7756,N_7339);
nand U8014 (N_8014,N_7007,N_7270);
xnor U8015 (N_8015,N_7380,N_7986);
nand U8016 (N_8016,N_7149,N_7592);
nor U8017 (N_8017,N_7348,N_7373);
nand U8018 (N_8018,N_7941,N_7595);
nand U8019 (N_8019,N_7832,N_7726);
nand U8020 (N_8020,N_7011,N_7492);
nand U8021 (N_8021,N_7346,N_7356);
nand U8022 (N_8022,N_7152,N_7068);
nand U8023 (N_8023,N_7160,N_7441);
and U8024 (N_8024,N_7255,N_7102);
nand U8025 (N_8025,N_7890,N_7514);
or U8026 (N_8026,N_7681,N_7925);
and U8027 (N_8027,N_7268,N_7845);
xnor U8028 (N_8028,N_7746,N_7718);
and U8029 (N_8029,N_7762,N_7956);
nor U8030 (N_8030,N_7367,N_7975);
nand U8031 (N_8031,N_7554,N_7653);
xnor U8032 (N_8032,N_7545,N_7032);
or U8033 (N_8033,N_7403,N_7119);
and U8034 (N_8034,N_7720,N_7561);
nand U8035 (N_8035,N_7660,N_7922);
nor U8036 (N_8036,N_7578,N_7954);
or U8037 (N_8037,N_7159,N_7549);
nand U8038 (N_8038,N_7258,N_7379);
and U8039 (N_8039,N_7461,N_7186);
nor U8040 (N_8040,N_7087,N_7801);
nand U8041 (N_8041,N_7778,N_7725);
nand U8042 (N_8042,N_7389,N_7636);
or U8043 (N_8043,N_7854,N_7569);
and U8044 (N_8044,N_7027,N_7645);
nor U8045 (N_8045,N_7033,N_7579);
or U8046 (N_8046,N_7467,N_7126);
and U8047 (N_8047,N_7520,N_7304);
nand U8048 (N_8048,N_7010,N_7525);
or U8049 (N_8049,N_7099,N_7177);
nor U8050 (N_8050,N_7316,N_7075);
nand U8051 (N_8051,N_7296,N_7158);
nand U8052 (N_8052,N_7903,N_7459);
nand U8053 (N_8053,N_7532,N_7387);
xnor U8054 (N_8054,N_7082,N_7533);
or U8055 (N_8055,N_7232,N_7086);
nand U8056 (N_8056,N_7342,N_7182);
nor U8057 (N_8057,N_7302,N_7222);
or U8058 (N_8058,N_7606,N_7081);
or U8059 (N_8059,N_7513,N_7743);
nor U8060 (N_8060,N_7805,N_7910);
or U8061 (N_8061,N_7717,N_7786);
nand U8062 (N_8062,N_7148,N_7345);
xnor U8063 (N_8063,N_7629,N_7924);
nor U8064 (N_8064,N_7305,N_7966);
and U8065 (N_8065,N_7708,N_7942);
or U8066 (N_8066,N_7065,N_7278);
nand U8067 (N_8067,N_7162,N_7411);
and U8068 (N_8068,N_7819,N_7529);
or U8069 (N_8069,N_7432,N_7239);
nor U8070 (N_8070,N_7115,N_7567);
and U8071 (N_8071,N_7051,N_7013);
and U8072 (N_8072,N_7498,N_7862);
and U8073 (N_8073,N_7308,N_7484);
nand U8074 (N_8074,N_7818,N_7881);
nor U8075 (N_8075,N_7934,N_7497);
and U8076 (N_8076,N_7883,N_7557);
or U8077 (N_8077,N_7321,N_7455);
xor U8078 (N_8078,N_7378,N_7097);
nor U8079 (N_8079,N_7123,N_7619);
or U8080 (N_8080,N_7029,N_7673);
nor U8081 (N_8081,N_7950,N_7889);
and U8082 (N_8082,N_7517,N_7669);
nor U8083 (N_8083,N_7362,N_7865);
or U8084 (N_8084,N_7482,N_7622);
nand U8085 (N_8085,N_7614,N_7624);
nand U8086 (N_8086,N_7164,N_7953);
nor U8087 (N_8087,N_7044,N_7390);
xor U8088 (N_8088,N_7092,N_7074);
nand U8089 (N_8089,N_7277,N_7063);
xor U8090 (N_8090,N_7654,N_7769);
or U8091 (N_8091,N_7078,N_7548);
or U8092 (N_8092,N_7217,N_7814);
or U8093 (N_8093,N_7927,N_7641);
nor U8094 (N_8094,N_7847,N_7117);
xor U8095 (N_8095,N_7703,N_7856);
or U8096 (N_8096,N_7035,N_7273);
or U8097 (N_8097,N_7145,N_7430);
nor U8098 (N_8098,N_7187,N_7830);
or U8099 (N_8099,N_7486,N_7325);
and U8100 (N_8100,N_7943,N_7633);
and U8101 (N_8101,N_7812,N_7562);
and U8102 (N_8102,N_7080,N_7958);
xor U8103 (N_8103,N_7853,N_7473);
xor U8104 (N_8104,N_7426,N_7596);
and U8105 (N_8105,N_7407,N_7113);
xnor U8106 (N_8106,N_7110,N_7704);
and U8107 (N_8107,N_7253,N_7571);
xor U8108 (N_8108,N_7827,N_7458);
or U8109 (N_8109,N_7091,N_7189);
or U8110 (N_8110,N_7695,N_7872);
and U8111 (N_8111,N_7154,N_7488);
and U8112 (N_8112,N_7952,N_7860);
nand U8113 (N_8113,N_7552,N_7949);
or U8114 (N_8114,N_7671,N_7803);
nor U8115 (N_8115,N_7314,N_7911);
nor U8116 (N_8116,N_7478,N_7285);
xnor U8117 (N_8117,N_7556,N_7324);
and U8118 (N_8118,N_7083,N_7133);
nor U8119 (N_8119,N_7898,N_7931);
nor U8120 (N_8120,N_7228,N_7310);
or U8121 (N_8121,N_7539,N_7331);
nand U8122 (N_8122,N_7166,N_7381);
and U8123 (N_8123,N_7023,N_7917);
nor U8124 (N_8124,N_7777,N_7406);
nand U8125 (N_8125,N_7623,N_7299);
nand U8126 (N_8126,N_7333,N_7440);
nand U8127 (N_8127,N_7017,N_7940);
nor U8128 (N_8128,N_7833,N_7598);
xor U8129 (N_8129,N_7794,N_7352);
and U8130 (N_8130,N_7738,N_7930);
nand U8131 (N_8131,N_7608,N_7503);
nor U8132 (N_8132,N_7098,N_7499);
xor U8133 (N_8133,N_7506,N_7522);
and U8134 (N_8134,N_7871,N_7020);
nor U8135 (N_8135,N_7468,N_7518);
nand U8136 (N_8136,N_7059,N_7524);
nand U8137 (N_8137,N_7997,N_7944);
or U8138 (N_8138,N_7611,N_7863);
nor U8139 (N_8139,N_7683,N_7427);
or U8140 (N_8140,N_7840,N_7060);
xor U8141 (N_8141,N_7684,N_7260);
or U8142 (N_8142,N_7919,N_7019);
nor U8143 (N_8143,N_7295,N_7784);
and U8144 (N_8144,N_7237,N_7878);
or U8145 (N_8145,N_7457,N_7572);
nor U8146 (N_8146,N_7587,N_7101);
nor U8147 (N_8147,N_7600,N_7991);
xor U8148 (N_8148,N_7904,N_7693);
and U8149 (N_8149,N_7179,N_7625);
and U8150 (N_8150,N_7825,N_7907);
or U8151 (N_8151,N_7796,N_7679);
nor U8152 (N_8152,N_7836,N_7343);
and U8153 (N_8153,N_7615,N_7724);
xnor U8154 (N_8154,N_7365,N_7982);
or U8155 (N_8155,N_7984,N_7672);
nand U8156 (N_8156,N_7588,N_7811);
nor U8157 (N_8157,N_7680,N_7519);
and U8158 (N_8158,N_7014,N_7885);
nand U8159 (N_8159,N_7398,N_7772);
xnor U8160 (N_8160,N_7837,N_7359);
nor U8161 (N_8161,N_7489,N_7477);
nor U8162 (N_8162,N_7480,N_7084);
nand U8163 (N_8163,N_7315,N_7790);
nand U8164 (N_8164,N_7580,N_7834);
nor U8165 (N_8165,N_7912,N_7460);
and U8166 (N_8166,N_7212,N_7251);
nand U8167 (N_8167,N_7347,N_7028);
nand U8168 (N_8168,N_7573,N_7586);
nand U8169 (N_8169,N_7575,N_7800);
xnor U8170 (N_8170,N_7985,N_7436);
nor U8171 (N_8171,N_7111,N_7742);
nand U8172 (N_8172,N_7008,N_7281);
nand U8173 (N_8173,N_7218,N_7445);
nor U8174 (N_8174,N_7353,N_7388);
and U8175 (N_8175,N_7916,N_7897);
or U8176 (N_8176,N_7291,N_7104);
nand U8177 (N_8177,N_7055,N_7320);
xnor U8178 (N_8178,N_7057,N_7495);
or U8179 (N_8179,N_7230,N_7740);
and U8180 (N_8180,N_7842,N_7076);
nand U8181 (N_8181,N_7161,N_7361);
and U8182 (N_8182,N_7939,N_7979);
nor U8183 (N_8183,N_7402,N_7349);
and U8184 (N_8184,N_7234,N_7209);
and U8185 (N_8185,N_7399,N_7583);
xnor U8186 (N_8186,N_7647,N_7405);
nand U8187 (N_8187,N_7874,N_7470);
nand U8188 (N_8188,N_7905,N_7297);
xor U8189 (N_8189,N_7948,N_7265);
or U8190 (N_8190,N_7947,N_7504);
and U8191 (N_8191,N_7298,N_7142);
or U8192 (N_8192,N_7327,N_7197);
or U8193 (N_8193,N_7538,N_7808);
or U8194 (N_8194,N_7039,N_7634);
nor U8195 (N_8195,N_7392,N_7085);
nand U8196 (N_8196,N_7329,N_7921);
and U8197 (N_8197,N_7763,N_7699);
or U8198 (N_8198,N_7946,N_7914);
and U8199 (N_8199,N_7536,N_7650);
or U8200 (N_8200,N_7377,N_7073);
or U8201 (N_8201,N_7038,N_7867);
nor U8202 (N_8202,N_7809,N_7134);
and U8203 (N_8203,N_7424,N_7058);
nor U8204 (N_8204,N_7555,N_7072);
and U8205 (N_8205,N_7971,N_7279);
nor U8206 (N_8206,N_7621,N_7355);
nor U8207 (N_8207,N_7668,N_7200);
and U8208 (N_8208,N_7560,N_7521);
nand U8209 (N_8209,N_7275,N_7512);
and U8210 (N_8210,N_7959,N_7244);
or U8211 (N_8211,N_7932,N_7835);
nor U8212 (N_8212,N_7205,N_7307);
or U8213 (N_8213,N_7481,N_7886);
or U8214 (N_8214,N_7690,N_7609);
and U8215 (N_8215,N_7848,N_7438);
nand U8216 (N_8216,N_7670,N_7995);
nor U8217 (N_8217,N_7382,N_7312);
nor U8218 (N_8218,N_7747,N_7516);
or U8219 (N_8219,N_7021,N_7216);
and U8220 (N_8220,N_7088,N_7689);
nand U8221 (N_8221,N_7607,N_7601);
nand U8222 (N_8222,N_7861,N_7748);
nand U8223 (N_8223,N_7899,N_7428);
xor U8224 (N_8224,N_7929,N_7233);
or U8225 (N_8225,N_7593,N_7354);
nand U8226 (N_8226,N_7371,N_7184);
and U8227 (N_8227,N_7715,N_7891);
or U8228 (N_8228,N_7707,N_7391);
xor U8229 (N_8229,N_7311,N_7433);
xor U8230 (N_8230,N_7866,N_7688);
nand U8231 (N_8231,N_7876,N_7155);
nor U8232 (N_8232,N_7095,N_7602);
nor U8233 (N_8233,N_7821,N_7697);
xnor U8234 (N_8234,N_7728,N_7293);
and U8235 (N_8235,N_7289,N_7219);
nand U8236 (N_8236,N_7737,N_7213);
nand U8237 (N_8237,N_7207,N_7173);
or U8238 (N_8238,N_7651,N_7879);
nor U8239 (N_8239,N_7198,N_7262);
or U8240 (N_8240,N_7630,N_7807);
and U8241 (N_8241,N_7214,N_7242);
or U8242 (N_8242,N_7386,N_7449);
nor U8243 (N_8243,N_7618,N_7201);
nand U8244 (N_8244,N_7224,N_7714);
xnor U8245 (N_8245,N_7241,N_7204);
or U8246 (N_8246,N_7828,N_7574);
or U8247 (N_8247,N_7920,N_7375);
nand U8248 (N_8248,N_7661,N_7906);
nand U8249 (N_8249,N_7616,N_7558);
nand U8250 (N_8250,N_7576,N_7016);
or U8251 (N_8251,N_7195,N_7464);
and U8252 (N_8252,N_7419,N_7317);
and U8253 (N_8253,N_7795,N_7852);
or U8254 (N_8254,N_7351,N_7804);
nor U8255 (N_8255,N_7272,N_7843);
and U8256 (N_8256,N_7712,N_7626);
nor U8257 (N_8257,N_7472,N_7700);
or U8258 (N_8258,N_7753,N_7036);
and U8259 (N_8259,N_7018,N_7147);
nor U8260 (N_8260,N_7442,N_7632);
nand U8261 (N_8261,N_7534,N_7857);
and U8262 (N_8262,N_7880,N_7168);
and U8263 (N_8263,N_7306,N_7376);
xnor U8264 (N_8264,N_7118,N_7393);
and U8265 (N_8265,N_7701,N_7108);
nor U8266 (N_8266,N_7485,N_7523);
and U8267 (N_8267,N_7450,N_7250);
xor U8268 (N_8268,N_7463,N_7140);
nor U8269 (N_8269,N_7873,N_7999);
nor U8270 (N_8270,N_7069,N_7962);
nand U8271 (N_8271,N_7103,N_7590);
nor U8272 (N_8272,N_7969,N_7188);
xnor U8273 (N_8273,N_7882,N_7096);
nand U8274 (N_8274,N_7719,N_7716);
nand U8275 (N_8275,N_7826,N_7431);
nor U8276 (N_8276,N_7146,N_7261);
nand U8277 (N_8277,N_7869,N_7423);
and U8278 (N_8278,N_7901,N_7181);
and U8279 (N_8279,N_7475,N_7884);
nand U8280 (N_8280,N_7729,N_7937);
or U8281 (N_8281,N_7501,N_7026);
and U8282 (N_8282,N_7271,N_7502);
or U8283 (N_8283,N_7444,N_7066);
or U8284 (N_8284,N_7395,N_7409);
nor U8285 (N_8285,N_7977,N_7792);
and U8286 (N_8286,N_7163,N_7300);
nand U8287 (N_8287,N_7220,N_7049);
nor U8288 (N_8288,N_7245,N_7003);
and U8289 (N_8289,N_7192,N_7806);
nand U8290 (N_8290,N_7603,N_7964);
xnor U8291 (N_8291,N_7227,N_7368);
and U8292 (N_8292,N_7175,N_7370);
and U8293 (N_8293,N_7323,N_7313);
nand U8294 (N_8294,N_7540,N_7276);
and U8295 (N_8295,N_7053,N_7183);
nor U8296 (N_8296,N_7256,N_7739);
and U8297 (N_8297,N_7435,N_7437);
xor U8298 (N_8298,N_7938,N_7752);
or U8299 (N_8299,N_7675,N_7462);
and U8300 (N_8300,N_7226,N_7282);
or U8301 (N_8301,N_7052,N_7960);
nor U8302 (N_8302,N_7259,N_7781);
nand U8303 (N_8303,N_7787,N_7638);
and U8304 (N_8304,N_7171,N_7820);
nor U8305 (N_8305,N_7094,N_7408);
xor U8306 (N_8306,N_7544,N_7363);
nor U8307 (N_8307,N_7543,N_7105);
nand U8308 (N_8308,N_7550,N_7635);
nand U8309 (N_8309,N_7429,N_7425);
and U8310 (N_8310,N_7056,N_7963);
or U8311 (N_8311,N_7535,N_7568);
and U8312 (N_8312,N_7372,N_7150);
or U8313 (N_8313,N_7537,N_7210);
and U8314 (N_8314,N_7945,N_7676);
xor U8315 (N_8315,N_7422,N_7079);
xnor U8316 (N_8316,N_7061,N_7730);
and U8317 (N_8317,N_7120,N_7090);
nand U8318 (N_8318,N_7526,N_7961);
and U8319 (N_8319,N_7465,N_7170);
nand U8320 (N_8320,N_7846,N_7508);
nand U8321 (N_8321,N_7788,N_7691);
xnor U8322 (N_8322,N_7267,N_7735);
nor U8323 (N_8323,N_7264,N_7996);
or U8324 (N_8324,N_7246,N_7721);
or U8325 (N_8325,N_7062,N_7269);
xnor U8326 (N_8326,N_7597,N_7476);
nand U8327 (N_8327,N_7319,N_7817);
nor U8328 (N_8328,N_7687,N_7733);
and U8329 (N_8329,N_7604,N_7723);
or U8330 (N_8330,N_7015,N_7143);
and U8331 (N_8331,N_7107,N_7448);
nand U8332 (N_8332,N_7420,N_7564);
nand U8333 (N_8333,N_7418,N_7570);
nand U8334 (N_8334,N_7868,N_7559);
and U8335 (N_8335,N_7093,N_7736);
and U8336 (N_8336,N_7479,N_7456);
or U8337 (N_8337,N_7350,N_7617);
nand U8338 (N_8338,N_7401,N_7374);
and U8339 (N_8339,N_7089,N_7169);
nor U8340 (N_8340,N_7751,N_7046);
and U8341 (N_8341,N_7713,N_7453);
nor U8342 (N_8342,N_7610,N_7613);
xor U8343 (N_8343,N_7301,N_7292);
nand U8344 (N_8344,N_7770,N_7421);
nand U8345 (N_8345,N_7667,N_7682);
and U8346 (N_8346,N_7994,N_7240);
or U8347 (N_8347,N_7988,N_7439);
nor U8348 (N_8348,N_7655,N_7211);
nand U8349 (N_8349,N_7384,N_7034);
and U8350 (N_8350,N_7254,N_7722);
or U8351 (N_8351,N_7396,N_7892);
nand U8352 (N_8352,N_7659,N_7754);
nand U8353 (N_8353,N_7417,N_7040);
or U8354 (N_8354,N_7434,N_7208);
xor U8355 (N_8355,N_7631,N_7993);
nor U8356 (N_8356,N_7839,N_7664);
and U8357 (N_8357,N_7983,N_7045);
nor U8358 (N_8358,N_7344,N_7895);
and U8359 (N_8359,N_7247,N_7176);
nor U8360 (N_8360,N_7178,N_7193);
nor U8361 (N_8361,N_7563,N_7791);
or U8362 (N_8362,N_7774,N_7757);
xnor U8363 (N_8363,N_7000,N_7799);
and U8364 (N_8364,N_7005,N_7710);
and U8365 (N_8365,N_7335,N_7900);
nand U8366 (N_8366,N_7410,N_7678);
nand U8367 (N_8367,N_7646,N_7491);
or U8368 (N_8368,N_7507,N_7235);
and U8369 (N_8369,N_7584,N_7841);
or U8370 (N_8370,N_7591,N_7965);
or U8371 (N_8371,N_7511,N_7412);
nor U8372 (N_8372,N_7542,N_7303);
nand U8373 (N_8373,N_7990,N_7454);
xor U8374 (N_8374,N_7202,N_7662);
nand U8375 (N_8375,N_7340,N_7686);
nand U8376 (N_8376,N_7706,N_7196);
nand U8377 (N_8377,N_7136,N_7338);
nand U8378 (N_8378,N_7987,N_7127);
nand U8379 (N_8379,N_7980,N_7553);
and U8380 (N_8380,N_7414,N_7585);
xnor U8381 (N_8381,N_7048,N_7446);
nand U8382 (N_8382,N_7582,N_7165);
xnor U8383 (N_8383,N_7864,N_7709);
and U8384 (N_8384,N_7124,N_7813);
and U8385 (N_8385,N_7185,N_7894);
nand U8386 (N_8386,N_7452,N_7322);
nand U8387 (N_8387,N_7731,N_7581);
or U8388 (N_8388,N_7989,N_7199);
or U8389 (N_8389,N_7823,N_7077);
nand U8390 (N_8390,N_7047,N_7829);
nor U8391 (N_8391,N_7050,N_7547);
nand U8392 (N_8392,N_7231,N_7755);
and U8393 (N_8393,N_7957,N_7215);
and U8394 (N_8394,N_7968,N_7926);
nor U8395 (N_8395,N_7628,N_7810);
and U8396 (N_8396,N_7493,N_7153);
nand U8397 (N_8397,N_7992,N_7334);
xnor U8398 (N_8398,N_7483,N_7494);
nand U8399 (N_8399,N_7223,N_7648);
or U8400 (N_8400,N_7109,N_7229);
and U8401 (N_8401,N_7649,N_7114);
nor U8402 (N_8402,N_7138,N_7067);
nand U8403 (N_8403,N_7877,N_7326);
nand U8404 (N_8404,N_7816,N_7252);
or U8405 (N_8405,N_7775,N_7850);
or U8406 (N_8406,N_7773,N_7531);
nand U8407 (N_8407,N_7274,N_7221);
nand U8408 (N_8408,N_7413,N_7385);
and U8409 (N_8409,N_7527,N_7913);
or U8410 (N_8410,N_7666,N_7469);
and U8411 (N_8411,N_7702,N_7783);
or U8412 (N_8412,N_7054,N_7510);
nand U8413 (N_8413,N_7789,N_7656);
and U8414 (N_8414,N_7369,N_7973);
nor U8415 (N_8415,N_7318,N_7070);
xnor U8416 (N_8416,N_7443,N_7759);
or U8417 (N_8417,N_7637,N_7257);
and U8418 (N_8418,N_7902,N_7998);
and U8419 (N_8419,N_7824,N_7766);
nor U8420 (N_8420,N_7970,N_7474);
xnor U8421 (N_8421,N_7838,N_7167);
and U8422 (N_8422,N_7263,N_7266);
nand U8423 (N_8423,N_7248,N_7357);
nand U8424 (N_8424,N_7505,N_7280);
or U8425 (N_8425,N_7785,N_7031);
and U8426 (N_8426,N_7627,N_7002);
nand U8427 (N_8427,N_7546,N_7206);
nand U8428 (N_8428,N_7674,N_7768);
nand U8429 (N_8429,N_7172,N_7741);
or U8430 (N_8430,N_7711,N_7337);
nand U8431 (N_8431,N_7551,N_7870);
or U8432 (N_8432,N_7121,N_7851);
and U8433 (N_8433,N_7758,N_7122);
and U8434 (N_8434,N_7336,N_7288);
nor U8435 (N_8435,N_7383,N_7129);
or U8436 (N_8436,N_7236,N_7530);
or U8437 (N_8437,N_7284,N_7692);
nor U8438 (N_8438,N_7203,N_7776);
and U8439 (N_8439,N_7400,N_7394);
xor U8440 (N_8440,N_7025,N_7001);
nor U8441 (N_8441,N_7887,N_7685);
and U8442 (N_8442,N_7243,N_7130);
nor U8443 (N_8443,N_7447,N_7566);
nand U8444 (N_8444,N_7663,N_7896);
or U8445 (N_8445,N_7487,N_7605);
nor U8446 (N_8446,N_7238,N_7599);
nand U8447 (N_8447,N_7009,N_7831);
and U8448 (N_8448,N_7750,N_7022);
or U8449 (N_8449,N_7125,N_7131);
and U8450 (N_8450,N_7652,N_7734);
or U8451 (N_8451,N_7802,N_7643);
nand U8452 (N_8452,N_7194,N_7908);
xor U8453 (N_8453,N_7849,N_7761);
or U8454 (N_8454,N_7644,N_7665);
nand U8455 (N_8455,N_7749,N_7225);
nand U8456 (N_8456,N_7844,N_7451);
or U8457 (N_8457,N_7620,N_7972);
or U8458 (N_8458,N_7918,N_7042);
or U8459 (N_8459,N_7797,N_7141);
xor U8460 (N_8460,N_7135,N_7727);
or U8461 (N_8461,N_7541,N_7030);
and U8462 (N_8462,N_7936,N_7677);
nand U8463 (N_8463,N_7144,N_7286);
nor U8464 (N_8464,N_7594,N_7190);
nor U8465 (N_8465,N_7978,N_7360);
or U8466 (N_8466,N_7100,N_7490);
nand U8467 (N_8467,N_7151,N_7358);
and U8468 (N_8468,N_7294,N_7782);
or U8469 (N_8469,N_7191,N_7967);
nor U8470 (N_8470,N_7780,N_7767);
or U8471 (N_8471,N_7642,N_7341);
nor U8472 (N_8472,N_7528,N_7858);
and U8473 (N_8473,N_7981,N_7976);
xor U8474 (N_8474,N_7951,N_7309);
and U8475 (N_8475,N_7745,N_7875);
nor U8476 (N_8476,N_7696,N_7915);
or U8477 (N_8477,N_7174,N_7639);
and U8478 (N_8478,N_7933,N_7466);
or U8479 (N_8479,N_7137,N_7156);
xor U8480 (N_8480,N_7157,N_7496);
and U8481 (N_8481,N_7024,N_7290);
and U8482 (N_8482,N_7565,N_7004);
nand U8483 (N_8483,N_7471,N_7888);
nand U8484 (N_8484,N_7694,N_7923);
nand U8485 (N_8485,N_7640,N_7955);
and U8486 (N_8486,N_7287,N_7006);
nor U8487 (N_8487,N_7765,N_7657);
and U8488 (N_8488,N_7859,N_7106);
and U8489 (N_8489,N_7500,N_7515);
and U8490 (N_8490,N_7012,N_7771);
nand U8491 (N_8491,N_7779,N_7974);
xor U8492 (N_8492,N_7732,N_7855);
or U8493 (N_8493,N_7416,N_7397);
and U8494 (N_8494,N_7041,N_7815);
nor U8495 (N_8495,N_7112,N_7764);
nand U8496 (N_8496,N_7043,N_7139);
or U8497 (N_8497,N_7589,N_7909);
nor U8498 (N_8498,N_7935,N_7415);
nand U8499 (N_8499,N_7116,N_7249);
xor U8500 (N_8500,N_7984,N_7219);
nor U8501 (N_8501,N_7359,N_7024);
nor U8502 (N_8502,N_7433,N_7118);
nand U8503 (N_8503,N_7946,N_7987);
nor U8504 (N_8504,N_7721,N_7751);
nor U8505 (N_8505,N_7601,N_7337);
nor U8506 (N_8506,N_7936,N_7907);
nor U8507 (N_8507,N_7301,N_7888);
or U8508 (N_8508,N_7100,N_7690);
nand U8509 (N_8509,N_7793,N_7152);
nand U8510 (N_8510,N_7031,N_7103);
and U8511 (N_8511,N_7020,N_7437);
nand U8512 (N_8512,N_7917,N_7805);
and U8513 (N_8513,N_7822,N_7167);
nor U8514 (N_8514,N_7857,N_7768);
or U8515 (N_8515,N_7299,N_7502);
nor U8516 (N_8516,N_7809,N_7667);
nor U8517 (N_8517,N_7149,N_7976);
nor U8518 (N_8518,N_7696,N_7690);
nand U8519 (N_8519,N_7274,N_7495);
nor U8520 (N_8520,N_7352,N_7286);
xnor U8521 (N_8521,N_7695,N_7624);
nor U8522 (N_8522,N_7861,N_7608);
nand U8523 (N_8523,N_7302,N_7234);
and U8524 (N_8524,N_7297,N_7097);
and U8525 (N_8525,N_7259,N_7112);
nand U8526 (N_8526,N_7521,N_7335);
and U8527 (N_8527,N_7751,N_7072);
nand U8528 (N_8528,N_7009,N_7463);
nand U8529 (N_8529,N_7299,N_7732);
and U8530 (N_8530,N_7009,N_7771);
and U8531 (N_8531,N_7729,N_7171);
xnor U8532 (N_8532,N_7741,N_7139);
nand U8533 (N_8533,N_7622,N_7993);
and U8534 (N_8534,N_7201,N_7151);
nand U8535 (N_8535,N_7389,N_7144);
nand U8536 (N_8536,N_7299,N_7167);
and U8537 (N_8537,N_7067,N_7180);
or U8538 (N_8538,N_7755,N_7838);
nand U8539 (N_8539,N_7105,N_7000);
nand U8540 (N_8540,N_7162,N_7406);
nor U8541 (N_8541,N_7904,N_7760);
nand U8542 (N_8542,N_7803,N_7146);
nor U8543 (N_8543,N_7522,N_7217);
nand U8544 (N_8544,N_7754,N_7979);
or U8545 (N_8545,N_7956,N_7298);
and U8546 (N_8546,N_7937,N_7702);
or U8547 (N_8547,N_7915,N_7119);
nand U8548 (N_8548,N_7894,N_7579);
and U8549 (N_8549,N_7819,N_7382);
or U8550 (N_8550,N_7352,N_7841);
nor U8551 (N_8551,N_7867,N_7086);
and U8552 (N_8552,N_7650,N_7133);
nand U8553 (N_8553,N_7352,N_7127);
or U8554 (N_8554,N_7648,N_7173);
and U8555 (N_8555,N_7008,N_7589);
nor U8556 (N_8556,N_7091,N_7312);
and U8557 (N_8557,N_7179,N_7468);
xnor U8558 (N_8558,N_7313,N_7432);
nor U8559 (N_8559,N_7345,N_7582);
and U8560 (N_8560,N_7775,N_7439);
nand U8561 (N_8561,N_7090,N_7220);
nor U8562 (N_8562,N_7868,N_7184);
or U8563 (N_8563,N_7459,N_7414);
and U8564 (N_8564,N_7932,N_7998);
nor U8565 (N_8565,N_7892,N_7163);
nor U8566 (N_8566,N_7187,N_7527);
nand U8567 (N_8567,N_7629,N_7454);
or U8568 (N_8568,N_7399,N_7784);
nand U8569 (N_8569,N_7086,N_7670);
or U8570 (N_8570,N_7319,N_7499);
or U8571 (N_8571,N_7926,N_7626);
or U8572 (N_8572,N_7100,N_7335);
and U8573 (N_8573,N_7932,N_7241);
nor U8574 (N_8574,N_7151,N_7773);
and U8575 (N_8575,N_7115,N_7020);
nand U8576 (N_8576,N_7410,N_7155);
xor U8577 (N_8577,N_7921,N_7673);
and U8578 (N_8578,N_7319,N_7339);
nor U8579 (N_8579,N_7113,N_7621);
and U8580 (N_8580,N_7942,N_7060);
and U8581 (N_8581,N_7336,N_7139);
nor U8582 (N_8582,N_7009,N_7999);
and U8583 (N_8583,N_7703,N_7711);
or U8584 (N_8584,N_7281,N_7080);
nor U8585 (N_8585,N_7698,N_7675);
xnor U8586 (N_8586,N_7787,N_7331);
and U8587 (N_8587,N_7799,N_7995);
nand U8588 (N_8588,N_7129,N_7546);
xor U8589 (N_8589,N_7343,N_7984);
and U8590 (N_8590,N_7935,N_7220);
and U8591 (N_8591,N_7177,N_7310);
and U8592 (N_8592,N_7792,N_7254);
and U8593 (N_8593,N_7347,N_7026);
or U8594 (N_8594,N_7480,N_7441);
nand U8595 (N_8595,N_7975,N_7404);
and U8596 (N_8596,N_7821,N_7234);
nand U8597 (N_8597,N_7914,N_7217);
nor U8598 (N_8598,N_7406,N_7395);
or U8599 (N_8599,N_7613,N_7865);
or U8600 (N_8600,N_7248,N_7626);
nand U8601 (N_8601,N_7227,N_7028);
nor U8602 (N_8602,N_7727,N_7697);
nand U8603 (N_8603,N_7721,N_7316);
and U8604 (N_8604,N_7535,N_7670);
or U8605 (N_8605,N_7958,N_7061);
and U8606 (N_8606,N_7281,N_7385);
nor U8607 (N_8607,N_7207,N_7526);
nand U8608 (N_8608,N_7769,N_7714);
nand U8609 (N_8609,N_7407,N_7971);
and U8610 (N_8610,N_7685,N_7229);
or U8611 (N_8611,N_7790,N_7535);
nor U8612 (N_8612,N_7293,N_7843);
nand U8613 (N_8613,N_7637,N_7948);
or U8614 (N_8614,N_7740,N_7275);
or U8615 (N_8615,N_7044,N_7456);
or U8616 (N_8616,N_7354,N_7984);
or U8617 (N_8617,N_7519,N_7655);
nand U8618 (N_8618,N_7908,N_7004);
nand U8619 (N_8619,N_7819,N_7917);
xnor U8620 (N_8620,N_7016,N_7152);
xor U8621 (N_8621,N_7614,N_7478);
xor U8622 (N_8622,N_7692,N_7603);
and U8623 (N_8623,N_7460,N_7049);
or U8624 (N_8624,N_7138,N_7908);
nor U8625 (N_8625,N_7122,N_7919);
nor U8626 (N_8626,N_7609,N_7154);
and U8627 (N_8627,N_7848,N_7658);
and U8628 (N_8628,N_7324,N_7065);
xor U8629 (N_8629,N_7600,N_7028);
nor U8630 (N_8630,N_7325,N_7885);
nor U8631 (N_8631,N_7584,N_7457);
or U8632 (N_8632,N_7723,N_7734);
nor U8633 (N_8633,N_7173,N_7324);
nor U8634 (N_8634,N_7096,N_7932);
and U8635 (N_8635,N_7005,N_7516);
and U8636 (N_8636,N_7426,N_7494);
and U8637 (N_8637,N_7198,N_7189);
and U8638 (N_8638,N_7394,N_7330);
or U8639 (N_8639,N_7036,N_7586);
nand U8640 (N_8640,N_7964,N_7494);
nor U8641 (N_8641,N_7798,N_7439);
and U8642 (N_8642,N_7372,N_7137);
nand U8643 (N_8643,N_7774,N_7669);
nand U8644 (N_8644,N_7918,N_7611);
or U8645 (N_8645,N_7158,N_7655);
nor U8646 (N_8646,N_7677,N_7545);
nand U8647 (N_8647,N_7479,N_7032);
or U8648 (N_8648,N_7598,N_7417);
xnor U8649 (N_8649,N_7711,N_7737);
and U8650 (N_8650,N_7413,N_7669);
xor U8651 (N_8651,N_7823,N_7902);
nand U8652 (N_8652,N_7759,N_7940);
nand U8653 (N_8653,N_7511,N_7060);
nor U8654 (N_8654,N_7084,N_7344);
xor U8655 (N_8655,N_7003,N_7192);
nand U8656 (N_8656,N_7162,N_7169);
or U8657 (N_8657,N_7715,N_7943);
nand U8658 (N_8658,N_7740,N_7555);
and U8659 (N_8659,N_7157,N_7996);
nor U8660 (N_8660,N_7812,N_7337);
nand U8661 (N_8661,N_7863,N_7944);
nor U8662 (N_8662,N_7560,N_7467);
xor U8663 (N_8663,N_7524,N_7119);
or U8664 (N_8664,N_7057,N_7454);
or U8665 (N_8665,N_7619,N_7239);
or U8666 (N_8666,N_7445,N_7211);
or U8667 (N_8667,N_7279,N_7594);
xnor U8668 (N_8668,N_7471,N_7224);
and U8669 (N_8669,N_7571,N_7730);
nand U8670 (N_8670,N_7649,N_7566);
and U8671 (N_8671,N_7489,N_7724);
or U8672 (N_8672,N_7281,N_7682);
nor U8673 (N_8673,N_7952,N_7337);
and U8674 (N_8674,N_7641,N_7647);
or U8675 (N_8675,N_7245,N_7699);
and U8676 (N_8676,N_7708,N_7187);
nor U8677 (N_8677,N_7817,N_7281);
nand U8678 (N_8678,N_7006,N_7267);
xor U8679 (N_8679,N_7959,N_7281);
nand U8680 (N_8680,N_7999,N_7945);
or U8681 (N_8681,N_7203,N_7052);
xnor U8682 (N_8682,N_7453,N_7268);
or U8683 (N_8683,N_7771,N_7458);
or U8684 (N_8684,N_7782,N_7973);
nand U8685 (N_8685,N_7722,N_7679);
xor U8686 (N_8686,N_7690,N_7987);
or U8687 (N_8687,N_7784,N_7833);
nand U8688 (N_8688,N_7418,N_7095);
nand U8689 (N_8689,N_7915,N_7866);
or U8690 (N_8690,N_7968,N_7100);
xor U8691 (N_8691,N_7703,N_7071);
nor U8692 (N_8692,N_7679,N_7914);
xnor U8693 (N_8693,N_7549,N_7074);
xor U8694 (N_8694,N_7528,N_7471);
nand U8695 (N_8695,N_7681,N_7840);
or U8696 (N_8696,N_7354,N_7889);
or U8697 (N_8697,N_7550,N_7253);
nand U8698 (N_8698,N_7492,N_7294);
nor U8699 (N_8699,N_7670,N_7810);
and U8700 (N_8700,N_7439,N_7454);
nand U8701 (N_8701,N_7275,N_7349);
and U8702 (N_8702,N_7074,N_7345);
or U8703 (N_8703,N_7603,N_7390);
nand U8704 (N_8704,N_7256,N_7104);
and U8705 (N_8705,N_7938,N_7779);
or U8706 (N_8706,N_7478,N_7198);
and U8707 (N_8707,N_7696,N_7487);
nand U8708 (N_8708,N_7236,N_7164);
nand U8709 (N_8709,N_7999,N_7262);
or U8710 (N_8710,N_7804,N_7588);
and U8711 (N_8711,N_7019,N_7596);
nand U8712 (N_8712,N_7845,N_7909);
nor U8713 (N_8713,N_7906,N_7869);
xnor U8714 (N_8714,N_7406,N_7719);
xnor U8715 (N_8715,N_7286,N_7626);
or U8716 (N_8716,N_7901,N_7028);
nand U8717 (N_8717,N_7038,N_7749);
or U8718 (N_8718,N_7582,N_7627);
nor U8719 (N_8719,N_7489,N_7975);
nor U8720 (N_8720,N_7215,N_7288);
nand U8721 (N_8721,N_7119,N_7628);
or U8722 (N_8722,N_7997,N_7491);
or U8723 (N_8723,N_7416,N_7006);
nor U8724 (N_8724,N_7955,N_7290);
nand U8725 (N_8725,N_7185,N_7920);
nand U8726 (N_8726,N_7613,N_7241);
nand U8727 (N_8727,N_7269,N_7288);
or U8728 (N_8728,N_7338,N_7107);
nor U8729 (N_8729,N_7845,N_7061);
nor U8730 (N_8730,N_7499,N_7652);
or U8731 (N_8731,N_7825,N_7776);
and U8732 (N_8732,N_7766,N_7893);
nor U8733 (N_8733,N_7050,N_7412);
or U8734 (N_8734,N_7861,N_7080);
nand U8735 (N_8735,N_7488,N_7737);
nor U8736 (N_8736,N_7710,N_7365);
and U8737 (N_8737,N_7328,N_7471);
or U8738 (N_8738,N_7959,N_7895);
nand U8739 (N_8739,N_7848,N_7949);
nor U8740 (N_8740,N_7774,N_7390);
nand U8741 (N_8741,N_7382,N_7601);
or U8742 (N_8742,N_7886,N_7645);
nand U8743 (N_8743,N_7842,N_7014);
or U8744 (N_8744,N_7309,N_7078);
nor U8745 (N_8745,N_7705,N_7500);
and U8746 (N_8746,N_7577,N_7173);
nor U8747 (N_8747,N_7973,N_7886);
nand U8748 (N_8748,N_7735,N_7908);
nor U8749 (N_8749,N_7000,N_7973);
nor U8750 (N_8750,N_7814,N_7762);
xor U8751 (N_8751,N_7457,N_7981);
nand U8752 (N_8752,N_7100,N_7414);
xor U8753 (N_8753,N_7057,N_7128);
or U8754 (N_8754,N_7245,N_7140);
nand U8755 (N_8755,N_7791,N_7682);
and U8756 (N_8756,N_7823,N_7775);
and U8757 (N_8757,N_7377,N_7844);
and U8758 (N_8758,N_7886,N_7670);
or U8759 (N_8759,N_7088,N_7034);
xnor U8760 (N_8760,N_7565,N_7439);
or U8761 (N_8761,N_7496,N_7128);
xnor U8762 (N_8762,N_7344,N_7685);
nor U8763 (N_8763,N_7812,N_7504);
and U8764 (N_8764,N_7454,N_7429);
or U8765 (N_8765,N_7740,N_7049);
nand U8766 (N_8766,N_7759,N_7247);
and U8767 (N_8767,N_7244,N_7375);
nand U8768 (N_8768,N_7867,N_7332);
and U8769 (N_8769,N_7467,N_7305);
nor U8770 (N_8770,N_7578,N_7886);
and U8771 (N_8771,N_7030,N_7658);
nand U8772 (N_8772,N_7268,N_7520);
nor U8773 (N_8773,N_7201,N_7358);
nor U8774 (N_8774,N_7237,N_7459);
and U8775 (N_8775,N_7756,N_7220);
nand U8776 (N_8776,N_7708,N_7589);
nor U8777 (N_8777,N_7086,N_7318);
nor U8778 (N_8778,N_7091,N_7322);
nor U8779 (N_8779,N_7113,N_7155);
xnor U8780 (N_8780,N_7638,N_7001);
nand U8781 (N_8781,N_7541,N_7232);
xnor U8782 (N_8782,N_7617,N_7564);
or U8783 (N_8783,N_7727,N_7600);
xnor U8784 (N_8784,N_7811,N_7015);
nor U8785 (N_8785,N_7583,N_7024);
nor U8786 (N_8786,N_7664,N_7208);
nand U8787 (N_8787,N_7197,N_7307);
nand U8788 (N_8788,N_7117,N_7402);
and U8789 (N_8789,N_7857,N_7417);
or U8790 (N_8790,N_7901,N_7958);
nor U8791 (N_8791,N_7994,N_7533);
nor U8792 (N_8792,N_7823,N_7263);
nor U8793 (N_8793,N_7827,N_7719);
nor U8794 (N_8794,N_7330,N_7922);
nand U8795 (N_8795,N_7275,N_7973);
nor U8796 (N_8796,N_7447,N_7192);
and U8797 (N_8797,N_7769,N_7579);
or U8798 (N_8798,N_7667,N_7835);
xor U8799 (N_8799,N_7164,N_7349);
or U8800 (N_8800,N_7323,N_7967);
and U8801 (N_8801,N_7080,N_7994);
and U8802 (N_8802,N_7222,N_7735);
and U8803 (N_8803,N_7991,N_7407);
nor U8804 (N_8804,N_7419,N_7263);
xor U8805 (N_8805,N_7002,N_7131);
nand U8806 (N_8806,N_7511,N_7602);
or U8807 (N_8807,N_7445,N_7831);
nand U8808 (N_8808,N_7210,N_7751);
nor U8809 (N_8809,N_7963,N_7444);
and U8810 (N_8810,N_7550,N_7978);
and U8811 (N_8811,N_7248,N_7748);
xnor U8812 (N_8812,N_7357,N_7608);
or U8813 (N_8813,N_7066,N_7122);
nor U8814 (N_8814,N_7288,N_7846);
nor U8815 (N_8815,N_7042,N_7236);
and U8816 (N_8816,N_7140,N_7038);
or U8817 (N_8817,N_7931,N_7389);
nor U8818 (N_8818,N_7752,N_7918);
and U8819 (N_8819,N_7036,N_7736);
nand U8820 (N_8820,N_7730,N_7340);
xor U8821 (N_8821,N_7207,N_7064);
or U8822 (N_8822,N_7053,N_7674);
nand U8823 (N_8823,N_7648,N_7711);
nand U8824 (N_8824,N_7017,N_7605);
nor U8825 (N_8825,N_7201,N_7330);
nor U8826 (N_8826,N_7262,N_7055);
or U8827 (N_8827,N_7477,N_7600);
and U8828 (N_8828,N_7864,N_7413);
nand U8829 (N_8829,N_7472,N_7423);
or U8830 (N_8830,N_7679,N_7345);
nand U8831 (N_8831,N_7003,N_7071);
nand U8832 (N_8832,N_7518,N_7008);
or U8833 (N_8833,N_7173,N_7611);
nor U8834 (N_8834,N_7235,N_7614);
xor U8835 (N_8835,N_7990,N_7181);
nand U8836 (N_8836,N_7815,N_7755);
nand U8837 (N_8837,N_7835,N_7153);
nor U8838 (N_8838,N_7819,N_7759);
nand U8839 (N_8839,N_7633,N_7177);
or U8840 (N_8840,N_7872,N_7456);
and U8841 (N_8841,N_7748,N_7783);
nand U8842 (N_8842,N_7179,N_7514);
and U8843 (N_8843,N_7354,N_7576);
xor U8844 (N_8844,N_7370,N_7403);
and U8845 (N_8845,N_7264,N_7752);
or U8846 (N_8846,N_7333,N_7660);
nor U8847 (N_8847,N_7132,N_7578);
xor U8848 (N_8848,N_7045,N_7189);
nand U8849 (N_8849,N_7356,N_7389);
nand U8850 (N_8850,N_7288,N_7499);
and U8851 (N_8851,N_7634,N_7151);
nor U8852 (N_8852,N_7545,N_7026);
or U8853 (N_8853,N_7282,N_7186);
or U8854 (N_8854,N_7777,N_7715);
nand U8855 (N_8855,N_7633,N_7204);
nand U8856 (N_8856,N_7251,N_7148);
or U8857 (N_8857,N_7357,N_7891);
and U8858 (N_8858,N_7157,N_7519);
or U8859 (N_8859,N_7709,N_7687);
nor U8860 (N_8860,N_7331,N_7955);
nand U8861 (N_8861,N_7429,N_7552);
nor U8862 (N_8862,N_7902,N_7225);
nand U8863 (N_8863,N_7284,N_7317);
and U8864 (N_8864,N_7080,N_7717);
xor U8865 (N_8865,N_7868,N_7467);
xor U8866 (N_8866,N_7105,N_7154);
nor U8867 (N_8867,N_7549,N_7757);
xnor U8868 (N_8868,N_7509,N_7361);
nand U8869 (N_8869,N_7455,N_7995);
nor U8870 (N_8870,N_7648,N_7602);
nand U8871 (N_8871,N_7419,N_7762);
nor U8872 (N_8872,N_7830,N_7387);
nor U8873 (N_8873,N_7792,N_7681);
nor U8874 (N_8874,N_7327,N_7610);
and U8875 (N_8875,N_7461,N_7575);
nor U8876 (N_8876,N_7350,N_7298);
nor U8877 (N_8877,N_7490,N_7053);
and U8878 (N_8878,N_7449,N_7124);
or U8879 (N_8879,N_7179,N_7116);
and U8880 (N_8880,N_7515,N_7163);
xor U8881 (N_8881,N_7766,N_7145);
and U8882 (N_8882,N_7408,N_7124);
nand U8883 (N_8883,N_7754,N_7210);
xor U8884 (N_8884,N_7067,N_7643);
or U8885 (N_8885,N_7153,N_7237);
nand U8886 (N_8886,N_7949,N_7775);
nor U8887 (N_8887,N_7348,N_7901);
or U8888 (N_8888,N_7954,N_7362);
and U8889 (N_8889,N_7336,N_7129);
nand U8890 (N_8890,N_7452,N_7733);
nor U8891 (N_8891,N_7091,N_7859);
nand U8892 (N_8892,N_7555,N_7940);
or U8893 (N_8893,N_7683,N_7284);
nand U8894 (N_8894,N_7233,N_7290);
xor U8895 (N_8895,N_7851,N_7201);
or U8896 (N_8896,N_7374,N_7920);
nor U8897 (N_8897,N_7151,N_7455);
nor U8898 (N_8898,N_7002,N_7483);
nor U8899 (N_8899,N_7361,N_7631);
and U8900 (N_8900,N_7049,N_7267);
nand U8901 (N_8901,N_7880,N_7221);
xor U8902 (N_8902,N_7076,N_7370);
nand U8903 (N_8903,N_7621,N_7811);
nor U8904 (N_8904,N_7268,N_7694);
nor U8905 (N_8905,N_7061,N_7023);
nand U8906 (N_8906,N_7713,N_7076);
nand U8907 (N_8907,N_7909,N_7959);
or U8908 (N_8908,N_7997,N_7638);
and U8909 (N_8909,N_7815,N_7343);
and U8910 (N_8910,N_7160,N_7756);
nand U8911 (N_8911,N_7161,N_7557);
nor U8912 (N_8912,N_7316,N_7934);
nand U8913 (N_8913,N_7720,N_7649);
nand U8914 (N_8914,N_7149,N_7999);
or U8915 (N_8915,N_7332,N_7572);
nor U8916 (N_8916,N_7347,N_7059);
nand U8917 (N_8917,N_7265,N_7871);
and U8918 (N_8918,N_7449,N_7832);
xnor U8919 (N_8919,N_7104,N_7184);
nand U8920 (N_8920,N_7258,N_7670);
or U8921 (N_8921,N_7889,N_7488);
or U8922 (N_8922,N_7853,N_7343);
nor U8923 (N_8923,N_7605,N_7306);
nand U8924 (N_8924,N_7909,N_7344);
or U8925 (N_8925,N_7389,N_7042);
nand U8926 (N_8926,N_7648,N_7835);
and U8927 (N_8927,N_7491,N_7792);
xnor U8928 (N_8928,N_7713,N_7800);
xor U8929 (N_8929,N_7200,N_7290);
xnor U8930 (N_8930,N_7594,N_7497);
and U8931 (N_8931,N_7294,N_7350);
and U8932 (N_8932,N_7424,N_7479);
and U8933 (N_8933,N_7480,N_7354);
nor U8934 (N_8934,N_7527,N_7101);
nand U8935 (N_8935,N_7271,N_7244);
or U8936 (N_8936,N_7240,N_7204);
xor U8937 (N_8937,N_7959,N_7913);
and U8938 (N_8938,N_7487,N_7301);
nand U8939 (N_8939,N_7959,N_7366);
and U8940 (N_8940,N_7415,N_7679);
xor U8941 (N_8941,N_7451,N_7846);
nor U8942 (N_8942,N_7814,N_7014);
nor U8943 (N_8943,N_7813,N_7037);
and U8944 (N_8944,N_7492,N_7583);
and U8945 (N_8945,N_7382,N_7033);
or U8946 (N_8946,N_7399,N_7512);
or U8947 (N_8947,N_7742,N_7140);
or U8948 (N_8948,N_7364,N_7703);
or U8949 (N_8949,N_7413,N_7794);
nand U8950 (N_8950,N_7803,N_7017);
nand U8951 (N_8951,N_7012,N_7277);
nor U8952 (N_8952,N_7922,N_7251);
and U8953 (N_8953,N_7478,N_7579);
or U8954 (N_8954,N_7459,N_7990);
nand U8955 (N_8955,N_7338,N_7202);
and U8956 (N_8956,N_7328,N_7141);
nand U8957 (N_8957,N_7646,N_7726);
xor U8958 (N_8958,N_7431,N_7489);
nand U8959 (N_8959,N_7850,N_7331);
xor U8960 (N_8960,N_7214,N_7668);
nand U8961 (N_8961,N_7072,N_7363);
nand U8962 (N_8962,N_7482,N_7929);
nand U8963 (N_8963,N_7319,N_7568);
nand U8964 (N_8964,N_7640,N_7685);
nand U8965 (N_8965,N_7030,N_7480);
or U8966 (N_8966,N_7862,N_7346);
and U8967 (N_8967,N_7061,N_7059);
nand U8968 (N_8968,N_7471,N_7687);
xnor U8969 (N_8969,N_7487,N_7039);
nor U8970 (N_8970,N_7969,N_7686);
or U8971 (N_8971,N_7668,N_7877);
or U8972 (N_8972,N_7485,N_7681);
nor U8973 (N_8973,N_7419,N_7216);
and U8974 (N_8974,N_7986,N_7013);
or U8975 (N_8975,N_7893,N_7822);
or U8976 (N_8976,N_7482,N_7855);
nor U8977 (N_8977,N_7124,N_7894);
and U8978 (N_8978,N_7153,N_7947);
or U8979 (N_8979,N_7166,N_7480);
nand U8980 (N_8980,N_7752,N_7288);
and U8981 (N_8981,N_7027,N_7547);
nor U8982 (N_8982,N_7400,N_7968);
nand U8983 (N_8983,N_7546,N_7585);
nor U8984 (N_8984,N_7216,N_7378);
or U8985 (N_8985,N_7407,N_7058);
nor U8986 (N_8986,N_7136,N_7493);
nor U8987 (N_8987,N_7809,N_7735);
xnor U8988 (N_8988,N_7679,N_7147);
or U8989 (N_8989,N_7404,N_7703);
nand U8990 (N_8990,N_7560,N_7317);
and U8991 (N_8991,N_7927,N_7021);
and U8992 (N_8992,N_7766,N_7606);
nor U8993 (N_8993,N_7357,N_7918);
nor U8994 (N_8994,N_7390,N_7559);
xor U8995 (N_8995,N_7210,N_7005);
nor U8996 (N_8996,N_7050,N_7682);
nor U8997 (N_8997,N_7598,N_7647);
and U8998 (N_8998,N_7049,N_7602);
nand U8999 (N_8999,N_7549,N_7534);
nor U9000 (N_9000,N_8452,N_8680);
nand U9001 (N_9001,N_8160,N_8659);
xor U9002 (N_9002,N_8396,N_8145);
nand U9003 (N_9003,N_8942,N_8669);
or U9004 (N_9004,N_8360,N_8662);
nand U9005 (N_9005,N_8989,N_8523);
and U9006 (N_9006,N_8799,N_8291);
nand U9007 (N_9007,N_8032,N_8563);
nand U9008 (N_9008,N_8244,N_8566);
nand U9009 (N_9009,N_8941,N_8255);
xnor U9010 (N_9010,N_8748,N_8629);
nand U9011 (N_9011,N_8029,N_8358);
nor U9012 (N_9012,N_8636,N_8077);
nor U9013 (N_9013,N_8637,N_8097);
nor U9014 (N_9014,N_8499,N_8818);
and U9015 (N_9015,N_8509,N_8290);
and U9016 (N_9016,N_8492,N_8897);
and U9017 (N_9017,N_8567,N_8908);
and U9018 (N_9018,N_8790,N_8046);
xor U9019 (N_9019,N_8640,N_8119);
nand U9020 (N_9020,N_8473,N_8342);
and U9021 (N_9021,N_8053,N_8139);
and U9022 (N_9022,N_8524,N_8346);
or U9023 (N_9023,N_8470,N_8453);
nand U9024 (N_9024,N_8088,N_8898);
and U9025 (N_9025,N_8374,N_8208);
nor U9026 (N_9026,N_8683,N_8067);
nand U9027 (N_9027,N_8540,N_8394);
nand U9028 (N_9028,N_8630,N_8154);
nand U9029 (N_9029,N_8658,N_8875);
or U9030 (N_9030,N_8366,N_8924);
or U9031 (N_9031,N_8901,N_8089);
nor U9032 (N_9032,N_8831,N_8857);
nand U9033 (N_9033,N_8546,N_8580);
or U9034 (N_9034,N_8064,N_8214);
nand U9035 (N_9035,N_8638,N_8239);
nor U9036 (N_9036,N_8568,N_8825);
and U9037 (N_9037,N_8118,N_8036);
or U9038 (N_9038,N_8450,N_8604);
or U9039 (N_9039,N_8850,N_8059);
and U9040 (N_9040,N_8371,N_8350);
or U9041 (N_9041,N_8186,N_8593);
xnor U9042 (N_9042,N_8550,N_8795);
or U9043 (N_9043,N_8802,N_8721);
nor U9044 (N_9044,N_8851,N_8312);
or U9045 (N_9045,N_8287,N_8080);
or U9046 (N_9046,N_8623,N_8933);
or U9047 (N_9047,N_8307,N_8297);
and U9048 (N_9048,N_8755,N_8914);
nand U9049 (N_9049,N_8133,N_8275);
nor U9050 (N_9050,N_8798,N_8811);
and U9051 (N_9051,N_8416,N_8175);
nor U9052 (N_9052,N_8494,N_8939);
nor U9053 (N_9053,N_8425,N_8664);
or U9054 (N_9054,N_8896,N_8206);
and U9055 (N_9055,N_8201,N_8986);
xnor U9056 (N_9056,N_8073,N_8316);
and U9057 (N_9057,N_8174,N_8966);
nand U9058 (N_9058,N_8180,N_8899);
nor U9059 (N_9059,N_8672,N_8243);
nor U9060 (N_9060,N_8171,N_8824);
and U9061 (N_9061,N_8838,N_8752);
nor U9062 (N_9062,N_8226,N_8987);
or U9063 (N_9063,N_8065,N_8935);
nand U9064 (N_9064,N_8022,N_8797);
nor U9065 (N_9065,N_8969,N_8707);
nand U9066 (N_9066,N_8903,N_8819);
or U9067 (N_9067,N_8197,N_8793);
and U9068 (N_9068,N_8729,N_8852);
and U9069 (N_9069,N_8227,N_8515);
nand U9070 (N_9070,N_8199,N_8500);
nand U9071 (N_9071,N_8009,N_8872);
and U9072 (N_9072,N_8808,N_8855);
xor U9073 (N_9073,N_8161,N_8098);
nand U9074 (N_9074,N_8198,N_8796);
nand U9075 (N_9075,N_8289,N_8355);
or U9076 (N_9076,N_8422,N_8002);
and U9077 (N_9077,N_8684,N_8541);
and U9078 (N_9078,N_8462,N_8578);
or U9079 (N_9079,N_8222,N_8397);
nor U9080 (N_9080,N_8308,N_8443);
and U9081 (N_9081,N_8948,N_8836);
and U9082 (N_9082,N_8419,N_8106);
xnor U9083 (N_9083,N_8958,N_8574);
and U9084 (N_9084,N_8950,N_8779);
nor U9085 (N_9085,N_8368,N_8887);
xor U9086 (N_9086,N_8114,N_8362);
xor U9087 (N_9087,N_8026,N_8900);
or U9088 (N_9088,N_8225,N_8019);
nand U9089 (N_9089,N_8033,N_8497);
and U9090 (N_9090,N_8367,N_8305);
or U9091 (N_9091,N_8188,N_8311);
nand U9092 (N_9092,N_8582,N_8863);
or U9093 (N_9093,N_8946,N_8881);
or U9094 (N_9094,N_8953,N_8163);
or U9095 (N_9095,N_8873,N_8276);
nand U9096 (N_9096,N_8714,N_8364);
nand U9097 (N_9097,N_8639,N_8781);
and U9098 (N_9098,N_8572,N_8870);
and U9099 (N_9099,N_8438,N_8038);
and U9100 (N_9100,N_8344,N_8705);
and U9101 (N_9101,N_8040,N_8733);
nor U9102 (N_9102,N_8528,N_8934);
or U9103 (N_9103,N_8666,N_8359);
xnor U9104 (N_9104,N_8159,N_8951);
and U9105 (N_9105,N_8379,N_8339);
and U9106 (N_9106,N_8151,N_8054);
or U9107 (N_9107,N_8738,N_8542);
xnor U9108 (N_9108,N_8888,N_8940);
and U9109 (N_9109,N_8232,N_8103);
nand U9110 (N_9110,N_8332,N_8189);
nand U9111 (N_9111,N_8746,N_8783);
or U9112 (N_9112,N_8150,N_8284);
nor U9113 (N_9113,N_8162,N_8608);
or U9114 (N_9114,N_8235,N_8107);
and U9115 (N_9115,N_8137,N_8156);
nand U9116 (N_9116,N_8879,N_8111);
or U9117 (N_9117,N_8943,N_8561);
and U9118 (N_9118,N_8476,N_8912);
nor U9119 (N_9119,N_8600,N_8677);
nor U9120 (N_9120,N_8092,N_8166);
and U9121 (N_9121,N_8084,N_8045);
and U9122 (N_9122,N_8442,N_8909);
nand U9123 (N_9123,N_8341,N_8230);
xnor U9124 (N_9124,N_8979,N_8164);
or U9125 (N_9125,N_8110,N_8502);
xnor U9126 (N_9126,N_8081,N_8329);
nand U9127 (N_9127,N_8196,N_8937);
and U9128 (N_9128,N_8085,N_8252);
xor U9129 (N_9129,N_8423,N_8005);
nor U9130 (N_9130,N_8330,N_8384);
nor U9131 (N_9131,N_8758,N_8884);
or U9132 (N_9132,N_8400,N_8792);
nand U9133 (N_9133,N_8468,N_8789);
or U9134 (N_9134,N_8913,N_8478);
xnor U9135 (N_9135,N_8635,N_8285);
and U9136 (N_9136,N_8778,N_8925);
nor U9137 (N_9137,N_8410,N_8292);
or U9138 (N_9138,N_8181,N_8559);
xor U9139 (N_9139,N_8667,N_8813);
or U9140 (N_9140,N_8585,N_8069);
or U9141 (N_9141,N_8015,N_8712);
and U9142 (N_9142,N_8218,N_8221);
or U9143 (N_9143,N_8929,N_8345);
nand U9144 (N_9144,N_8253,N_8869);
nand U9145 (N_9145,N_8126,N_8217);
nand U9146 (N_9146,N_8723,N_8931);
or U9147 (N_9147,N_8169,N_8433);
nor U9148 (N_9148,N_8759,N_8724);
nand U9149 (N_9149,N_8762,N_8775);
nand U9150 (N_9150,N_8245,N_8039);
and U9151 (N_9151,N_8628,N_8482);
and U9152 (N_9152,N_8518,N_8261);
nand U9153 (N_9153,N_8391,N_8978);
or U9154 (N_9154,N_8657,N_8093);
nor U9155 (N_9155,N_8765,N_8105);
nand U9156 (N_9156,N_8668,N_8320);
and U9157 (N_9157,N_8554,N_8434);
or U9158 (N_9158,N_8573,N_8907);
nand U9159 (N_9159,N_8076,N_8317);
and U9160 (N_9160,N_8385,N_8956);
nand U9161 (N_9161,N_8975,N_8099);
or U9162 (N_9162,N_8418,N_8340);
and U9163 (N_9163,N_8735,N_8140);
or U9164 (N_9164,N_8516,N_8203);
and U9165 (N_9165,N_8314,N_8272);
or U9166 (N_9166,N_8801,N_8277);
nand U9167 (N_9167,N_8063,N_8674);
nor U9168 (N_9168,N_8378,N_8094);
or U9169 (N_9169,N_8967,N_8124);
nor U9170 (N_9170,N_8372,N_8902);
nand U9171 (N_9171,N_8743,N_8459);
or U9172 (N_9172,N_8766,N_8671);
xor U9173 (N_9173,N_8552,N_8395);
xor U9174 (N_9174,N_8176,N_8837);
nand U9175 (N_9175,N_8689,N_8483);
and U9176 (N_9176,N_8382,N_8963);
nand U9177 (N_9177,N_8619,N_8172);
nor U9178 (N_9178,N_8158,N_8056);
or U9179 (N_9179,N_8555,N_8965);
and U9180 (N_9180,N_8938,N_8503);
nand U9181 (N_9181,N_8142,N_8457);
or U9182 (N_9182,N_8467,N_8806);
or U9183 (N_9183,N_8233,N_8420);
nor U9184 (N_9184,N_8890,N_8918);
nand U9185 (N_9185,N_8977,N_8694);
nand U9186 (N_9186,N_8034,N_8061);
and U9187 (N_9187,N_8547,N_8242);
and U9188 (N_9188,N_8370,N_8356);
nand U9189 (N_9189,N_8115,N_8445);
nor U9190 (N_9190,N_8835,N_8012);
xor U9191 (N_9191,N_8584,N_8999);
nor U9192 (N_9192,N_8266,N_8731);
nand U9193 (N_9193,N_8876,N_8464);
and U9194 (N_9194,N_8024,N_8335);
and U9195 (N_9195,N_8794,N_8363);
or U9196 (N_9196,N_8834,N_8407);
and U9197 (N_9197,N_8011,N_8651);
or U9198 (N_9198,N_8429,N_8220);
xor U9199 (N_9199,N_8772,N_8010);
nor U9200 (N_9200,N_8641,N_8016);
and U9201 (N_9201,N_8071,N_8083);
nand U9202 (N_9202,N_8532,N_8644);
xor U9203 (N_9203,N_8670,N_8613);
or U9204 (N_9204,N_8463,N_8602);
nor U9205 (N_9205,N_8178,N_8601);
or U9206 (N_9206,N_8507,N_8191);
nand U9207 (N_9207,N_8592,N_8751);
and U9208 (N_9208,N_8823,N_8534);
or U9209 (N_9209,N_8720,N_8116);
and U9210 (N_9210,N_8262,N_8001);
and U9211 (N_9211,N_8096,N_8553);
or U9212 (N_9212,N_8771,N_8513);
or U9213 (N_9213,N_8496,N_8611);
nand U9214 (N_9214,N_8321,N_8776);
or U9215 (N_9215,N_8860,N_8066);
or U9216 (N_9216,N_8971,N_8047);
and U9217 (N_9217,N_8803,N_8343);
or U9218 (N_9218,N_8859,N_8996);
or U9219 (N_9219,N_8068,N_8589);
or U9220 (N_9220,N_8179,N_8926);
nor U9221 (N_9221,N_8195,N_8136);
nor U9222 (N_9222,N_8968,N_8642);
nor U9223 (N_9223,N_8815,N_8928);
or U9224 (N_9224,N_8231,N_8849);
or U9225 (N_9225,N_8440,N_8558);
xnor U9226 (N_9226,N_8624,N_8104);
xnor U9227 (N_9227,N_8216,N_8121);
nor U9228 (N_9228,N_8294,N_8535);
nor U9229 (N_9229,N_8165,N_8021);
nand U9230 (N_9230,N_8460,N_8742);
or U9231 (N_9231,N_8280,N_8544);
and U9232 (N_9232,N_8338,N_8247);
nor U9233 (N_9233,N_8577,N_8660);
and U9234 (N_9234,N_8536,N_8152);
and U9235 (N_9235,N_8980,N_8764);
and U9236 (N_9236,N_8679,N_8525);
nand U9237 (N_9237,N_8351,N_8389);
nand U9238 (N_9238,N_8204,N_8006);
nor U9239 (N_9239,N_8143,N_8148);
nor U9240 (N_9240,N_8543,N_8424);
nand U9241 (N_9241,N_8974,N_8052);
nand U9242 (N_9242,N_8474,N_8529);
or U9243 (N_9243,N_8932,N_8549);
nand U9244 (N_9244,N_8883,N_8281);
nor U9245 (N_9245,N_8557,N_8769);
nand U9246 (N_9246,N_8484,N_8210);
and U9247 (N_9247,N_8004,N_8736);
nor U9248 (N_9248,N_8380,N_8194);
and U9249 (N_9249,N_8739,N_8828);
or U9250 (N_9250,N_8533,N_8606);
and U9251 (N_9251,N_8990,N_8517);
nand U9252 (N_9252,N_8882,N_8185);
and U9253 (N_9253,N_8787,N_8030);
or U9254 (N_9254,N_8605,N_8548);
or U9255 (N_9255,N_8538,N_8248);
nand U9256 (N_9256,N_8961,N_8822);
nor U9257 (N_9257,N_8927,N_8877);
and U9258 (N_9258,N_8257,N_8477);
and U9259 (N_9259,N_8295,N_8962);
nand U9260 (N_9260,N_8153,N_8991);
and U9261 (N_9261,N_8774,N_8387);
and U9262 (N_9262,N_8028,N_8530);
nor U9263 (N_9263,N_8401,N_8035);
nand U9264 (N_9264,N_8784,N_8955);
nor U9265 (N_9265,N_8101,N_8236);
and U9266 (N_9266,N_8665,N_8414);
and U9267 (N_9267,N_8936,N_8072);
nand U9268 (N_9268,N_8632,N_8493);
nor U9269 (N_9269,N_8841,N_8686);
xor U9270 (N_9270,N_8631,N_8487);
nor U9271 (N_9271,N_8113,N_8485);
nand U9272 (N_9272,N_8108,N_8000);
and U9273 (N_9273,N_8596,N_8479);
nand U9274 (N_9274,N_8594,N_8565);
or U9275 (N_9275,N_8983,N_8708);
nand U9276 (N_9276,N_8435,N_8273);
or U9277 (N_9277,N_8480,N_8048);
and U9278 (N_9278,N_8082,N_8481);
and U9279 (N_9279,N_8267,N_8504);
and U9280 (N_9280,N_8120,N_8322);
nor U9281 (N_9281,N_8695,N_8747);
or U9282 (N_9282,N_8182,N_8168);
or U9283 (N_9283,N_8144,N_8209);
or U9284 (N_9284,N_8810,N_8475);
nand U9285 (N_9285,N_8564,N_8981);
nand U9286 (N_9286,N_8885,N_8620);
or U9287 (N_9287,N_8597,N_8390);
or U9288 (N_9288,N_8122,N_8131);
and U9289 (N_9289,N_8049,N_8649);
nor U9290 (N_9290,N_8313,N_8087);
nor U9291 (N_9291,N_8134,N_8854);
nand U9292 (N_9292,N_8972,N_8023);
and U9293 (N_9293,N_8719,N_8675);
and U9294 (N_9294,N_8676,N_8112);
and U9295 (N_9295,N_8466,N_8471);
nand U9296 (N_9296,N_8519,N_8760);
and U9297 (N_9297,N_8691,N_8610);
or U9298 (N_9298,N_8603,N_8698);
or U9299 (N_9299,N_8415,N_8693);
xor U9300 (N_9300,N_8782,N_8439);
nand U9301 (N_9301,N_8997,N_8058);
nand U9302 (N_9302,N_8861,N_8051);
nand U9303 (N_9303,N_8283,N_8522);
nand U9304 (N_9304,N_8428,N_8491);
nor U9305 (N_9305,N_8498,N_8654);
nand U9306 (N_9306,N_8044,N_8512);
nor U9307 (N_9307,N_8095,N_8309);
and U9308 (N_9308,N_8944,N_8167);
and U9309 (N_9309,N_8386,N_8376);
and U9310 (N_9310,N_8985,N_8399);
or U9311 (N_9311,N_8617,N_8791);
nand U9312 (N_9312,N_8263,N_8856);
nor U9313 (N_9313,N_8832,N_8070);
and U9314 (N_9314,N_8612,N_8408);
nor U9315 (N_9315,N_8703,N_8973);
nor U9316 (N_9316,N_8412,N_8469);
and U9317 (N_9317,N_8258,N_8993);
xor U9318 (N_9318,N_8609,N_8265);
nand U9319 (N_9319,N_8352,N_8296);
or U9320 (N_9320,N_8060,N_8207);
and U9321 (N_9321,N_8816,N_8090);
or U9322 (N_9322,N_8741,N_8920);
nor U9323 (N_9323,N_8527,N_8922);
and U9324 (N_9324,N_8687,N_8886);
nor U9325 (N_9325,N_8685,N_8431);
nor U9326 (N_9326,N_8506,N_8757);
nor U9327 (N_9327,N_8375,N_8696);
nor U9328 (N_9328,N_8269,N_8055);
and U9329 (N_9329,N_8017,N_8681);
and U9330 (N_9330,N_8353,N_8446);
and U9331 (N_9331,N_8960,N_8994);
xor U9332 (N_9332,N_8461,N_8615);
nand U9333 (N_9333,N_8043,N_8328);
nor U9334 (N_9334,N_8270,N_8146);
and U9335 (N_9335,N_8279,N_8906);
nand U9336 (N_9336,N_8393,N_8411);
and U9337 (N_9337,N_8732,N_8020);
or U9338 (N_9338,N_8616,N_8773);
nand U9339 (N_9339,N_8531,N_8777);
nand U9340 (N_9340,N_8868,N_8436);
nand U9341 (N_9341,N_8880,N_8373);
nand U9342 (N_9342,N_8298,N_8805);
nand U9343 (N_9343,N_8228,N_8817);
nor U9344 (N_9344,N_8652,N_8599);
or U9345 (N_9345,N_8354,N_8646);
nand U9346 (N_9346,N_8916,N_8141);
or U9347 (N_9347,N_8614,N_8347);
nand U9348 (N_9348,N_8734,N_8587);
nand U9349 (N_9349,N_8234,N_8753);
or U9350 (N_9350,N_8398,N_8318);
and U9351 (N_9351,N_8132,N_8042);
or U9352 (N_9352,N_8581,N_8964);
nand U9353 (N_9353,N_8193,N_8304);
or U9354 (N_9354,N_8062,N_8643);
nand U9355 (N_9355,N_8455,N_8840);
nor U9356 (N_9356,N_8212,N_8634);
or U9357 (N_9357,N_8930,N_8821);
nor U9358 (N_9358,N_8853,N_8571);
xor U9359 (N_9359,N_8403,N_8315);
nand U9360 (N_9360,N_8844,N_8337);
and U9361 (N_9361,N_8319,N_8895);
nand U9362 (N_9362,N_8891,N_8079);
or U9363 (N_9363,N_8770,N_8598);
nand U9364 (N_9364,N_8947,N_8240);
or U9365 (N_9365,N_8357,N_8656);
or U9366 (N_9366,N_8745,N_8688);
nand U9367 (N_9367,N_8911,N_8713);
and U9368 (N_9368,N_8183,N_8763);
nand U9369 (N_9369,N_8545,N_8505);
and U9370 (N_9370,N_8075,N_8100);
nand U9371 (N_9371,N_8383,N_8488);
nor U9372 (N_9372,N_8444,N_8264);
nor U9373 (N_9373,N_8648,N_8187);
or U9374 (N_9374,N_8490,N_8867);
xnor U9375 (N_9375,N_8678,N_8976);
and U9376 (N_9376,N_8388,N_8846);
and U9377 (N_9377,N_8756,N_8814);
nand U9378 (N_9378,N_8893,N_8915);
xor U9379 (N_9379,N_8673,N_8905);
or U9380 (N_9380,N_8702,N_8710);
and U9381 (N_9381,N_8537,N_8726);
and U9382 (N_9382,N_8954,N_8421);
nor U9383 (N_9383,N_8878,N_8406);
or U9384 (N_9384,N_8224,N_8447);
nand U9385 (N_9385,N_8449,N_8441);
xnor U9386 (N_9386,N_8833,N_8249);
nor U9387 (N_9387,N_8008,N_8586);
and U9388 (N_9388,N_8278,N_8570);
or U9389 (N_9389,N_8510,N_8219);
nor U9390 (N_9390,N_8091,N_8331);
xor U9391 (N_9391,N_8626,N_8377);
or U9392 (N_9392,N_8725,N_8740);
and U9393 (N_9393,N_8800,N_8995);
and U9394 (N_9394,N_8129,N_8303);
and U9395 (N_9395,N_8716,N_8402);
nand U9396 (N_9396,N_8192,N_8715);
and U9397 (N_9397,N_8501,N_8865);
or U9398 (N_9398,N_8551,N_8690);
nand U9399 (N_9399,N_8826,N_8959);
and U9400 (N_9400,N_8301,N_8699);
nand U9401 (N_9401,N_8286,N_8361);
xnor U9402 (N_9402,N_8454,N_8750);
or U9403 (N_9403,N_8157,N_8575);
or U9404 (N_9404,N_8405,N_8205);
nand U9405 (N_9405,N_8919,N_8871);
or U9406 (N_9406,N_8299,N_8730);
nor U9407 (N_9407,N_8845,N_8706);
and U9408 (N_9408,N_8917,N_8013);
and U9409 (N_9409,N_8709,N_8842);
and U9410 (N_9410,N_8588,N_8495);
nor U9411 (N_9411,N_8237,N_8737);
and U9412 (N_9412,N_8591,N_8300);
and U9413 (N_9413,N_8014,N_8663);
nor U9414 (N_9414,N_8562,N_8190);
or U9415 (N_9415,N_8768,N_8788);
nor U9416 (N_9416,N_8583,N_8923);
and U9417 (N_9417,N_8829,N_8025);
nand U9418 (N_9418,N_8704,N_8874);
or U9419 (N_9419,N_8744,N_8256);
and U9420 (N_9420,N_8569,N_8489);
xor U9421 (N_9421,N_8866,N_8627);
nand U9422 (N_9422,N_8381,N_8050);
or U9423 (N_9423,N_8982,N_8722);
nand U9424 (N_9424,N_8456,N_8430);
and U9425 (N_9425,N_8125,N_8348);
or U9426 (N_9426,N_8647,N_8655);
and U9427 (N_9427,N_8369,N_8451);
and U9428 (N_9428,N_8123,N_8645);
or U9429 (N_9429,N_8149,N_8754);
nand U9430 (N_9430,N_8211,N_8173);
and U9431 (N_9431,N_8780,N_8892);
nor U9432 (N_9432,N_8254,N_8988);
and U9433 (N_9433,N_8250,N_8238);
nor U9434 (N_9434,N_8692,N_8334);
and U9435 (N_9435,N_8520,N_8984);
nand U9436 (N_9436,N_8945,N_8392);
xor U9437 (N_9437,N_8310,N_8306);
or U9438 (N_9438,N_8785,N_8894);
xnor U9439 (N_9439,N_8809,N_8260);
or U9440 (N_9440,N_8807,N_8268);
or U9441 (N_9441,N_8184,N_8147);
or U9442 (N_9442,N_8018,N_8078);
and U9443 (N_9443,N_8701,N_8661);
and U9444 (N_9444,N_8223,N_8843);
or U9445 (N_9445,N_8427,N_8700);
or U9446 (N_9446,N_8633,N_8508);
or U9447 (N_9447,N_8847,N_8618);
or U9448 (N_9448,N_8526,N_8711);
or U9449 (N_9449,N_8576,N_8830);
or U9450 (N_9450,N_8992,N_8007);
nor U9451 (N_9451,N_8417,N_8697);
or U9452 (N_9452,N_8625,N_8130);
nand U9453 (N_9453,N_8458,N_8595);
or U9454 (N_9454,N_8349,N_8579);
nor U9455 (N_9455,N_8448,N_8426);
or U9456 (N_9456,N_8622,N_8336);
xnor U9457 (N_9457,N_8117,N_8325);
and U9458 (N_9458,N_8003,N_8213);
nor U9459 (N_9459,N_8998,N_8202);
nand U9460 (N_9460,N_8259,N_8511);
nand U9461 (N_9461,N_8102,N_8952);
or U9462 (N_9462,N_8889,N_8607);
or U9463 (N_9463,N_8404,N_8864);
nor U9464 (N_9464,N_8718,N_8653);
or U9465 (N_9465,N_8282,N_8432);
or U9466 (N_9466,N_8293,N_8109);
and U9467 (N_9467,N_8302,N_8215);
nor U9468 (N_9468,N_8086,N_8177);
xnor U9469 (N_9469,N_8949,N_8074);
and U9470 (N_9470,N_8170,N_8155);
and U9471 (N_9471,N_8057,N_8804);
nor U9472 (N_9472,N_8413,N_8970);
nor U9473 (N_9473,N_8128,N_8727);
and U9474 (N_9474,N_8326,N_8858);
nand U9475 (N_9475,N_8037,N_8041);
nand U9476 (N_9476,N_8241,N_8274);
nand U9477 (N_9477,N_8465,N_8323);
or U9478 (N_9478,N_8728,N_8786);
nor U9479 (N_9479,N_8812,N_8324);
and U9480 (N_9480,N_8472,N_8717);
nand U9481 (N_9481,N_8138,N_8031);
and U9482 (N_9482,N_8848,N_8027);
nor U9483 (N_9483,N_8365,N_8910);
xnor U9484 (N_9484,N_8621,N_8904);
nand U9485 (N_9485,N_8820,N_8437);
nor U9486 (N_9486,N_8288,N_8539);
or U9487 (N_9487,N_8590,N_8827);
xor U9488 (N_9488,N_8409,N_8514);
or U9489 (N_9489,N_8246,N_8560);
nor U9490 (N_9490,N_8327,N_8486);
nor U9491 (N_9491,N_8271,N_8749);
or U9492 (N_9492,N_8251,N_8200);
or U9493 (N_9493,N_8650,N_8862);
or U9494 (N_9494,N_8521,N_8127);
and U9495 (N_9495,N_8767,N_8921);
nor U9496 (N_9496,N_8333,N_8839);
nor U9497 (N_9497,N_8556,N_8135);
nand U9498 (N_9498,N_8761,N_8229);
nor U9499 (N_9499,N_8682,N_8957);
nand U9500 (N_9500,N_8573,N_8138);
and U9501 (N_9501,N_8841,N_8265);
nor U9502 (N_9502,N_8520,N_8281);
and U9503 (N_9503,N_8321,N_8884);
nand U9504 (N_9504,N_8124,N_8931);
or U9505 (N_9505,N_8151,N_8436);
and U9506 (N_9506,N_8184,N_8481);
and U9507 (N_9507,N_8424,N_8404);
nor U9508 (N_9508,N_8154,N_8273);
xnor U9509 (N_9509,N_8672,N_8351);
nand U9510 (N_9510,N_8291,N_8744);
nand U9511 (N_9511,N_8198,N_8883);
xnor U9512 (N_9512,N_8503,N_8891);
or U9513 (N_9513,N_8778,N_8149);
nor U9514 (N_9514,N_8200,N_8018);
nand U9515 (N_9515,N_8520,N_8546);
nor U9516 (N_9516,N_8572,N_8250);
or U9517 (N_9517,N_8471,N_8111);
xnor U9518 (N_9518,N_8296,N_8189);
xor U9519 (N_9519,N_8348,N_8258);
nand U9520 (N_9520,N_8492,N_8481);
nor U9521 (N_9521,N_8675,N_8651);
nor U9522 (N_9522,N_8792,N_8421);
nand U9523 (N_9523,N_8648,N_8092);
nor U9524 (N_9524,N_8118,N_8891);
nor U9525 (N_9525,N_8868,N_8844);
or U9526 (N_9526,N_8947,N_8313);
xor U9527 (N_9527,N_8251,N_8649);
nand U9528 (N_9528,N_8949,N_8941);
and U9529 (N_9529,N_8630,N_8723);
or U9530 (N_9530,N_8516,N_8806);
and U9531 (N_9531,N_8386,N_8204);
and U9532 (N_9532,N_8304,N_8487);
xnor U9533 (N_9533,N_8385,N_8052);
and U9534 (N_9534,N_8496,N_8633);
nand U9535 (N_9535,N_8810,N_8500);
or U9536 (N_9536,N_8107,N_8083);
nand U9537 (N_9537,N_8031,N_8912);
and U9538 (N_9538,N_8161,N_8459);
nand U9539 (N_9539,N_8215,N_8083);
xor U9540 (N_9540,N_8620,N_8306);
and U9541 (N_9541,N_8631,N_8068);
nand U9542 (N_9542,N_8848,N_8091);
or U9543 (N_9543,N_8843,N_8157);
or U9544 (N_9544,N_8379,N_8316);
and U9545 (N_9545,N_8822,N_8702);
and U9546 (N_9546,N_8562,N_8668);
nor U9547 (N_9547,N_8823,N_8564);
nand U9548 (N_9548,N_8990,N_8280);
or U9549 (N_9549,N_8705,N_8975);
or U9550 (N_9550,N_8390,N_8989);
xor U9551 (N_9551,N_8048,N_8358);
nand U9552 (N_9552,N_8323,N_8642);
nand U9553 (N_9553,N_8875,N_8215);
nand U9554 (N_9554,N_8380,N_8128);
and U9555 (N_9555,N_8922,N_8779);
nor U9556 (N_9556,N_8133,N_8735);
nor U9557 (N_9557,N_8406,N_8208);
nand U9558 (N_9558,N_8202,N_8949);
or U9559 (N_9559,N_8466,N_8489);
nor U9560 (N_9560,N_8479,N_8545);
and U9561 (N_9561,N_8147,N_8822);
nor U9562 (N_9562,N_8894,N_8386);
xnor U9563 (N_9563,N_8397,N_8179);
or U9564 (N_9564,N_8810,N_8364);
nor U9565 (N_9565,N_8243,N_8835);
or U9566 (N_9566,N_8131,N_8799);
xnor U9567 (N_9567,N_8409,N_8698);
or U9568 (N_9568,N_8781,N_8769);
and U9569 (N_9569,N_8216,N_8889);
nand U9570 (N_9570,N_8643,N_8850);
or U9571 (N_9571,N_8238,N_8972);
and U9572 (N_9572,N_8487,N_8694);
and U9573 (N_9573,N_8106,N_8454);
and U9574 (N_9574,N_8577,N_8330);
or U9575 (N_9575,N_8399,N_8720);
or U9576 (N_9576,N_8876,N_8916);
nand U9577 (N_9577,N_8466,N_8724);
xor U9578 (N_9578,N_8114,N_8782);
and U9579 (N_9579,N_8807,N_8407);
or U9580 (N_9580,N_8638,N_8097);
xnor U9581 (N_9581,N_8050,N_8755);
or U9582 (N_9582,N_8447,N_8197);
nand U9583 (N_9583,N_8321,N_8630);
or U9584 (N_9584,N_8344,N_8507);
nor U9585 (N_9585,N_8617,N_8216);
xor U9586 (N_9586,N_8621,N_8588);
nand U9587 (N_9587,N_8620,N_8167);
and U9588 (N_9588,N_8510,N_8768);
xnor U9589 (N_9589,N_8078,N_8000);
and U9590 (N_9590,N_8753,N_8809);
nor U9591 (N_9591,N_8193,N_8010);
or U9592 (N_9592,N_8661,N_8009);
or U9593 (N_9593,N_8318,N_8581);
and U9594 (N_9594,N_8594,N_8550);
nor U9595 (N_9595,N_8977,N_8196);
or U9596 (N_9596,N_8201,N_8125);
or U9597 (N_9597,N_8111,N_8627);
and U9598 (N_9598,N_8048,N_8765);
nand U9599 (N_9599,N_8866,N_8652);
nand U9600 (N_9600,N_8443,N_8118);
nand U9601 (N_9601,N_8711,N_8548);
nor U9602 (N_9602,N_8394,N_8553);
or U9603 (N_9603,N_8179,N_8719);
nor U9604 (N_9604,N_8658,N_8080);
nand U9605 (N_9605,N_8820,N_8541);
or U9606 (N_9606,N_8547,N_8878);
nor U9607 (N_9607,N_8690,N_8571);
or U9608 (N_9608,N_8075,N_8161);
nand U9609 (N_9609,N_8497,N_8748);
nand U9610 (N_9610,N_8510,N_8123);
nor U9611 (N_9611,N_8238,N_8123);
nor U9612 (N_9612,N_8803,N_8146);
and U9613 (N_9613,N_8691,N_8292);
nor U9614 (N_9614,N_8849,N_8005);
xor U9615 (N_9615,N_8731,N_8893);
nand U9616 (N_9616,N_8770,N_8652);
xnor U9617 (N_9617,N_8602,N_8242);
or U9618 (N_9618,N_8670,N_8589);
xnor U9619 (N_9619,N_8582,N_8558);
and U9620 (N_9620,N_8897,N_8562);
xnor U9621 (N_9621,N_8101,N_8476);
nand U9622 (N_9622,N_8998,N_8513);
and U9623 (N_9623,N_8784,N_8602);
nand U9624 (N_9624,N_8993,N_8855);
nor U9625 (N_9625,N_8051,N_8034);
xnor U9626 (N_9626,N_8024,N_8342);
nor U9627 (N_9627,N_8798,N_8701);
and U9628 (N_9628,N_8380,N_8381);
and U9629 (N_9629,N_8619,N_8493);
xnor U9630 (N_9630,N_8714,N_8234);
nor U9631 (N_9631,N_8816,N_8310);
xnor U9632 (N_9632,N_8742,N_8659);
xor U9633 (N_9633,N_8522,N_8280);
nor U9634 (N_9634,N_8545,N_8213);
nor U9635 (N_9635,N_8184,N_8392);
or U9636 (N_9636,N_8710,N_8797);
nand U9637 (N_9637,N_8188,N_8625);
xnor U9638 (N_9638,N_8989,N_8434);
nand U9639 (N_9639,N_8730,N_8555);
nand U9640 (N_9640,N_8688,N_8727);
nand U9641 (N_9641,N_8238,N_8049);
nand U9642 (N_9642,N_8240,N_8319);
nor U9643 (N_9643,N_8059,N_8209);
nand U9644 (N_9644,N_8444,N_8985);
and U9645 (N_9645,N_8791,N_8334);
xor U9646 (N_9646,N_8606,N_8269);
nor U9647 (N_9647,N_8761,N_8167);
nor U9648 (N_9648,N_8489,N_8089);
or U9649 (N_9649,N_8795,N_8650);
nand U9650 (N_9650,N_8082,N_8490);
nand U9651 (N_9651,N_8230,N_8375);
nor U9652 (N_9652,N_8447,N_8635);
or U9653 (N_9653,N_8174,N_8048);
xor U9654 (N_9654,N_8511,N_8627);
xor U9655 (N_9655,N_8678,N_8452);
nand U9656 (N_9656,N_8999,N_8807);
nand U9657 (N_9657,N_8913,N_8533);
and U9658 (N_9658,N_8769,N_8879);
nand U9659 (N_9659,N_8087,N_8562);
and U9660 (N_9660,N_8999,N_8835);
or U9661 (N_9661,N_8029,N_8387);
nor U9662 (N_9662,N_8603,N_8883);
xnor U9663 (N_9663,N_8199,N_8735);
nor U9664 (N_9664,N_8110,N_8669);
or U9665 (N_9665,N_8875,N_8607);
and U9666 (N_9666,N_8498,N_8239);
and U9667 (N_9667,N_8403,N_8180);
or U9668 (N_9668,N_8963,N_8259);
xor U9669 (N_9669,N_8818,N_8152);
or U9670 (N_9670,N_8845,N_8295);
nand U9671 (N_9671,N_8506,N_8259);
and U9672 (N_9672,N_8059,N_8828);
or U9673 (N_9673,N_8003,N_8824);
or U9674 (N_9674,N_8815,N_8510);
nor U9675 (N_9675,N_8367,N_8576);
xor U9676 (N_9676,N_8375,N_8150);
and U9677 (N_9677,N_8064,N_8304);
and U9678 (N_9678,N_8442,N_8750);
nand U9679 (N_9679,N_8102,N_8358);
nor U9680 (N_9680,N_8577,N_8529);
or U9681 (N_9681,N_8200,N_8104);
nor U9682 (N_9682,N_8763,N_8385);
and U9683 (N_9683,N_8754,N_8392);
nand U9684 (N_9684,N_8882,N_8888);
or U9685 (N_9685,N_8183,N_8719);
nor U9686 (N_9686,N_8402,N_8446);
nand U9687 (N_9687,N_8524,N_8317);
and U9688 (N_9688,N_8630,N_8807);
nor U9689 (N_9689,N_8975,N_8291);
nand U9690 (N_9690,N_8607,N_8528);
nor U9691 (N_9691,N_8364,N_8203);
or U9692 (N_9692,N_8818,N_8881);
or U9693 (N_9693,N_8582,N_8484);
nor U9694 (N_9694,N_8091,N_8570);
and U9695 (N_9695,N_8646,N_8316);
and U9696 (N_9696,N_8800,N_8389);
and U9697 (N_9697,N_8505,N_8294);
or U9698 (N_9698,N_8951,N_8681);
nor U9699 (N_9699,N_8437,N_8420);
or U9700 (N_9700,N_8376,N_8334);
or U9701 (N_9701,N_8603,N_8713);
or U9702 (N_9702,N_8956,N_8864);
nand U9703 (N_9703,N_8410,N_8261);
and U9704 (N_9704,N_8160,N_8588);
or U9705 (N_9705,N_8528,N_8592);
or U9706 (N_9706,N_8979,N_8800);
and U9707 (N_9707,N_8711,N_8596);
or U9708 (N_9708,N_8040,N_8422);
nand U9709 (N_9709,N_8720,N_8033);
or U9710 (N_9710,N_8552,N_8365);
xor U9711 (N_9711,N_8073,N_8502);
nor U9712 (N_9712,N_8701,N_8238);
and U9713 (N_9713,N_8385,N_8841);
nor U9714 (N_9714,N_8979,N_8884);
or U9715 (N_9715,N_8943,N_8946);
and U9716 (N_9716,N_8973,N_8827);
or U9717 (N_9717,N_8370,N_8234);
or U9718 (N_9718,N_8877,N_8588);
nand U9719 (N_9719,N_8409,N_8243);
nand U9720 (N_9720,N_8693,N_8219);
and U9721 (N_9721,N_8916,N_8595);
or U9722 (N_9722,N_8756,N_8507);
nand U9723 (N_9723,N_8761,N_8553);
or U9724 (N_9724,N_8681,N_8234);
nand U9725 (N_9725,N_8618,N_8263);
nand U9726 (N_9726,N_8139,N_8860);
and U9727 (N_9727,N_8467,N_8670);
and U9728 (N_9728,N_8212,N_8449);
and U9729 (N_9729,N_8214,N_8900);
nand U9730 (N_9730,N_8148,N_8353);
and U9731 (N_9731,N_8813,N_8676);
nor U9732 (N_9732,N_8215,N_8087);
and U9733 (N_9733,N_8463,N_8328);
or U9734 (N_9734,N_8266,N_8661);
or U9735 (N_9735,N_8581,N_8284);
nand U9736 (N_9736,N_8863,N_8686);
nand U9737 (N_9737,N_8181,N_8741);
or U9738 (N_9738,N_8346,N_8827);
xnor U9739 (N_9739,N_8468,N_8067);
or U9740 (N_9740,N_8762,N_8069);
xnor U9741 (N_9741,N_8463,N_8206);
and U9742 (N_9742,N_8237,N_8215);
or U9743 (N_9743,N_8581,N_8514);
and U9744 (N_9744,N_8678,N_8067);
and U9745 (N_9745,N_8245,N_8083);
and U9746 (N_9746,N_8318,N_8719);
nor U9747 (N_9747,N_8419,N_8031);
nand U9748 (N_9748,N_8701,N_8341);
or U9749 (N_9749,N_8862,N_8267);
and U9750 (N_9750,N_8960,N_8329);
and U9751 (N_9751,N_8788,N_8296);
or U9752 (N_9752,N_8634,N_8979);
nor U9753 (N_9753,N_8432,N_8143);
and U9754 (N_9754,N_8037,N_8379);
nand U9755 (N_9755,N_8595,N_8507);
or U9756 (N_9756,N_8839,N_8509);
and U9757 (N_9757,N_8867,N_8922);
nand U9758 (N_9758,N_8350,N_8349);
or U9759 (N_9759,N_8833,N_8136);
nand U9760 (N_9760,N_8115,N_8110);
or U9761 (N_9761,N_8218,N_8641);
and U9762 (N_9762,N_8348,N_8829);
xor U9763 (N_9763,N_8253,N_8556);
nand U9764 (N_9764,N_8752,N_8490);
nand U9765 (N_9765,N_8425,N_8139);
or U9766 (N_9766,N_8014,N_8606);
nand U9767 (N_9767,N_8393,N_8761);
and U9768 (N_9768,N_8546,N_8771);
nand U9769 (N_9769,N_8380,N_8156);
nor U9770 (N_9770,N_8703,N_8665);
nand U9771 (N_9771,N_8539,N_8088);
or U9772 (N_9772,N_8937,N_8339);
xnor U9773 (N_9773,N_8411,N_8801);
or U9774 (N_9774,N_8892,N_8645);
or U9775 (N_9775,N_8406,N_8611);
or U9776 (N_9776,N_8673,N_8991);
and U9777 (N_9777,N_8781,N_8599);
nand U9778 (N_9778,N_8691,N_8618);
or U9779 (N_9779,N_8921,N_8116);
or U9780 (N_9780,N_8420,N_8081);
xnor U9781 (N_9781,N_8158,N_8425);
or U9782 (N_9782,N_8769,N_8380);
nor U9783 (N_9783,N_8725,N_8857);
nand U9784 (N_9784,N_8341,N_8248);
and U9785 (N_9785,N_8007,N_8086);
or U9786 (N_9786,N_8528,N_8501);
nand U9787 (N_9787,N_8691,N_8402);
nor U9788 (N_9788,N_8654,N_8750);
nor U9789 (N_9789,N_8129,N_8407);
and U9790 (N_9790,N_8244,N_8452);
nand U9791 (N_9791,N_8488,N_8017);
nand U9792 (N_9792,N_8787,N_8267);
or U9793 (N_9793,N_8373,N_8388);
nor U9794 (N_9794,N_8052,N_8863);
nor U9795 (N_9795,N_8136,N_8811);
and U9796 (N_9796,N_8693,N_8159);
or U9797 (N_9797,N_8939,N_8518);
and U9798 (N_9798,N_8600,N_8267);
and U9799 (N_9799,N_8871,N_8219);
and U9800 (N_9800,N_8250,N_8995);
nor U9801 (N_9801,N_8377,N_8155);
or U9802 (N_9802,N_8204,N_8646);
nand U9803 (N_9803,N_8591,N_8792);
nand U9804 (N_9804,N_8444,N_8193);
or U9805 (N_9805,N_8517,N_8602);
or U9806 (N_9806,N_8600,N_8051);
nor U9807 (N_9807,N_8966,N_8944);
nor U9808 (N_9808,N_8249,N_8197);
or U9809 (N_9809,N_8351,N_8937);
or U9810 (N_9810,N_8003,N_8339);
and U9811 (N_9811,N_8124,N_8216);
nor U9812 (N_9812,N_8382,N_8511);
nand U9813 (N_9813,N_8112,N_8337);
or U9814 (N_9814,N_8901,N_8204);
nor U9815 (N_9815,N_8022,N_8609);
nand U9816 (N_9816,N_8110,N_8971);
xnor U9817 (N_9817,N_8663,N_8547);
and U9818 (N_9818,N_8483,N_8270);
xor U9819 (N_9819,N_8565,N_8296);
xor U9820 (N_9820,N_8827,N_8146);
nor U9821 (N_9821,N_8567,N_8407);
or U9822 (N_9822,N_8053,N_8759);
and U9823 (N_9823,N_8334,N_8558);
or U9824 (N_9824,N_8842,N_8327);
and U9825 (N_9825,N_8961,N_8823);
nor U9826 (N_9826,N_8481,N_8400);
and U9827 (N_9827,N_8932,N_8261);
xor U9828 (N_9828,N_8250,N_8313);
and U9829 (N_9829,N_8592,N_8473);
xnor U9830 (N_9830,N_8661,N_8093);
nand U9831 (N_9831,N_8744,N_8245);
nand U9832 (N_9832,N_8360,N_8703);
nor U9833 (N_9833,N_8734,N_8099);
and U9834 (N_9834,N_8783,N_8136);
xor U9835 (N_9835,N_8971,N_8408);
nand U9836 (N_9836,N_8297,N_8612);
xnor U9837 (N_9837,N_8264,N_8762);
nor U9838 (N_9838,N_8711,N_8308);
nor U9839 (N_9839,N_8527,N_8253);
and U9840 (N_9840,N_8999,N_8275);
nand U9841 (N_9841,N_8938,N_8964);
nand U9842 (N_9842,N_8419,N_8878);
or U9843 (N_9843,N_8438,N_8385);
nand U9844 (N_9844,N_8176,N_8168);
nor U9845 (N_9845,N_8491,N_8332);
nor U9846 (N_9846,N_8272,N_8912);
nor U9847 (N_9847,N_8896,N_8291);
and U9848 (N_9848,N_8658,N_8220);
or U9849 (N_9849,N_8895,N_8443);
xor U9850 (N_9850,N_8759,N_8619);
xnor U9851 (N_9851,N_8822,N_8380);
nor U9852 (N_9852,N_8574,N_8363);
nand U9853 (N_9853,N_8831,N_8877);
nor U9854 (N_9854,N_8438,N_8550);
and U9855 (N_9855,N_8702,N_8992);
nand U9856 (N_9856,N_8277,N_8959);
xnor U9857 (N_9857,N_8857,N_8674);
and U9858 (N_9858,N_8162,N_8925);
or U9859 (N_9859,N_8589,N_8575);
or U9860 (N_9860,N_8859,N_8579);
or U9861 (N_9861,N_8811,N_8067);
nand U9862 (N_9862,N_8878,N_8405);
nor U9863 (N_9863,N_8011,N_8080);
xor U9864 (N_9864,N_8237,N_8390);
or U9865 (N_9865,N_8559,N_8956);
nand U9866 (N_9866,N_8284,N_8412);
or U9867 (N_9867,N_8102,N_8934);
and U9868 (N_9868,N_8821,N_8127);
nor U9869 (N_9869,N_8494,N_8792);
and U9870 (N_9870,N_8456,N_8865);
nor U9871 (N_9871,N_8016,N_8309);
or U9872 (N_9872,N_8852,N_8457);
nand U9873 (N_9873,N_8270,N_8482);
xor U9874 (N_9874,N_8133,N_8301);
nand U9875 (N_9875,N_8590,N_8060);
xnor U9876 (N_9876,N_8979,N_8568);
or U9877 (N_9877,N_8769,N_8021);
or U9878 (N_9878,N_8392,N_8435);
and U9879 (N_9879,N_8626,N_8183);
nor U9880 (N_9880,N_8043,N_8344);
nor U9881 (N_9881,N_8013,N_8055);
or U9882 (N_9882,N_8982,N_8692);
or U9883 (N_9883,N_8792,N_8746);
xor U9884 (N_9884,N_8235,N_8700);
or U9885 (N_9885,N_8062,N_8597);
or U9886 (N_9886,N_8332,N_8481);
nand U9887 (N_9887,N_8308,N_8287);
nand U9888 (N_9888,N_8309,N_8230);
nor U9889 (N_9889,N_8657,N_8130);
or U9890 (N_9890,N_8911,N_8826);
nand U9891 (N_9891,N_8737,N_8854);
and U9892 (N_9892,N_8588,N_8226);
nor U9893 (N_9893,N_8292,N_8524);
and U9894 (N_9894,N_8216,N_8784);
nand U9895 (N_9895,N_8442,N_8787);
and U9896 (N_9896,N_8520,N_8159);
or U9897 (N_9897,N_8300,N_8814);
or U9898 (N_9898,N_8529,N_8217);
and U9899 (N_9899,N_8539,N_8307);
nand U9900 (N_9900,N_8475,N_8974);
nor U9901 (N_9901,N_8211,N_8946);
xnor U9902 (N_9902,N_8294,N_8189);
xnor U9903 (N_9903,N_8268,N_8372);
or U9904 (N_9904,N_8338,N_8549);
or U9905 (N_9905,N_8529,N_8193);
and U9906 (N_9906,N_8415,N_8322);
or U9907 (N_9907,N_8870,N_8555);
and U9908 (N_9908,N_8941,N_8227);
xor U9909 (N_9909,N_8008,N_8776);
xnor U9910 (N_9910,N_8546,N_8409);
nand U9911 (N_9911,N_8800,N_8649);
nand U9912 (N_9912,N_8137,N_8949);
nor U9913 (N_9913,N_8771,N_8726);
nand U9914 (N_9914,N_8672,N_8895);
or U9915 (N_9915,N_8397,N_8994);
nor U9916 (N_9916,N_8223,N_8741);
and U9917 (N_9917,N_8764,N_8542);
or U9918 (N_9918,N_8924,N_8796);
xor U9919 (N_9919,N_8167,N_8034);
xnor U9920 (N_9920,N_8626,N_8061);
and U9921 (N_9921,N_8244,N_8117);
and U9922 (N_9922,N_8023,N_8277);
or U9923 (N_9923,N_8998,N_8699);
nand U9924 (N_9924,N_8389,N_8788);
nor U9925 (N_9925,N_8945,N_8190);
xor U9926 (N_9926,N_8635,N_8784);
and U9927 (N_9927,N_8503,N_8677);
nand U9928 (N_9928,N_8357,N_8384);
xor U9929 (N_9929,N_8502,N_8151);
nand U9930 (N_9930,N_8297,N_8625);
nand U9931 (N_9931,N_8161,N_8470);
nand U9932 (N_9932,N_8373,N_8340);
nor U9933 (N_9933,N_8603,N_8534);
or U9934 (N_9934,N_8507,N_8406);
or U9935 (N_9935,N_8648,N_8048);
nand U9936 (N_9936,N_8804,N_8012);
and U9937 (N_9937,N_8519,N_8027);
nand U9938 (N_9938,N_8663,N_8210);
nor U9939 (N_9939,N_8666,N_8939);
or U9940 (N_9940,N_8860,N_8626);
nor U9941 (N_9941,N_8139,N_8118);
or U9942 (N_9942,N_8775,N_8722);
nor U9943 (N_9943,N_8444,N_8129);
xnor U9944 (N_9944,N_8160,N_8229);
nand U9945 (N_9945,N_8066,N_8391);
and U9946 (N_9946,N_8258,N_8136);
or U9947 (N_9947,N_8093,N_8768);
nor U9948 (N_9948,N_8041,N_8146);
nand U9949 (N_9949,N_8852,N_8983);
nand U9950 (N_9950,N_8560,N_8968);
and U9951 (N_9951,N_8954,N_8276);
and U9952 (N_9952,N_8329,N_8612);
nor U9953 (N_9953,N_8722,N_8106);
nand U9954 (N_9954,N_8105,N_8391);
and U9955 (N_9955,N_8372,N_8003);
and U9956 (N_9956,N_8128,N_8798);
or U9957 (N_9957,N_8378,N_8409);
and U9958 (N_9958,N_8737,N_8606);
and U9959 (N_9959,N_8987,N_8016);
or U9960 (N_9960,N_8122,N_8019);
or U9961 (N_9961,N_8054,N_8598);
and U9962 (N_9962,N_8993,N_8428);
and U9963 (N_9963,N_8269,N_8378);
nor U9964 (N_9964,N_8629,N_8688);
xnor U9965 (N_9965,N_8160,N_8948);
and U9966 (N_9966,N_8305,N_8986);
nand U9967 (N_9967,N_8188,N_8391);
or U9968 (N_9968,N_8607,N_8148);
nor U9969 (N_9969,N_8974,N_8292);
nand U9970 (N_9970,N_8828,N_8390);
or U9971 (N_9971,N_8190,N_8910);
nand U9972 (N_9972,N_8224,N_8162);
xor U9973 (N_9973,N_8104,N_8757);
nand U9974 (N_9974,N_8066,N_8181);
or U9975 (N_9975,N_8474,N_8328);
and U9976 (N_9976,N_8327,N_8555);
nand U9977 (N_9977,N_8109,N_8938);
and U9978 (N_9978,N_8381,N_8080);
nand U9979 (N_9979,N_8249,N_8575);
and U9980 (N_9980,N_8261,N_8258);
or U9981 (N_9981,N_8263,N_8956);
nor U9982 (N_9982,N_8391,N_8340);
nor U9983 (N_9983,N_8634,N_8314);
and U9984 (N_9984,N_8930,N_8631);
or U9985 (N_9985,N_8013,N_8530);
nand U9986 (N_9986,N_8073,N_8260);
and U9987 (N_9987,N_8919,N_8339);
nand U9988 (N_9988,N_8027,N_8236);
and U9989 (N_9989,N_8862,N_8438);
nand U9990 (N_9990,N_8459,N_8876);
xnor U9991 (N_9991,N_8668,N_8751);
nor U9992 (N_9992,N_8674,N_8755);
nor U9993 (N_9993,N_8538,N_8945);
and U9994 (N_9994,N_8338,N_8363);
nor U9995 (N_9995,N_8523,N_8344);
xnor U9996 (N_9996,N_8551,N_8786);
nor U9997 (N_9997,N_8268,N_8096);
nor U9998 (N_9998,N_8650,N_8189);
nor U9999 (N_9999,N_8815,N_8054);
or UO_0 (O_0,N_9907,N_9876);
nand UO_1 (O_1,N_9118,N_9098);
or UO_2 (O_2,N_9846,N_9038);
nor UO_3 (O_3,N_9799,N_9933);
nand UO_4 (O_4,N_9247,N_9204);
and UO_5 (O_5,N_9935,N_9823);
xnor UO_6 (O_6,N_9684,N_9558);
and UO_7 (O_7,N_9710,N_9365);
nor UO_8 (O_8,N_9533,N_9553);
and UO_9 (O_9,N_9664,N_9912);
xor UO_10 (O_10,N_9295,N_9244);
and UO_11 (O_11,N_9028,N_9720);
nand UO_12 (O_12,N_9181,N_9769);
xor UO_13 (O_13,N_9721,N_9438);
nor UO_14 (O_14,N_9406,N_9063);
and UO_15 (O_15,N_9851,N_9812);
nor UO_16 (O_16,N_9497,N_9747);
and UO_17 (O_17,N_9178,N_9580);
nor UO_18 (O_18,N_9530,N_9635);
nor UO_19 (O_19,N_9871,N_9566);
nand UO_20 (O_20,N_9427,N_9976);
or UO_21 (O_21,N_9877,N_9766);
and UO_22 (O_22,N_9674,N_9361);
or UO_23 (O_23,N_9188,N_9571);
xnor UO_24 (O_24,N_9627,N_9453);
or UO_25 (O_25,N_9158,N_9528);
and UO_26 (O_26,N_9486,N_9650);
or UO_27 (O_27,N_9875,N_9210);
or UO_28 (O_28,N_9140,N_9013);
nor UO_29 (O_29,N_9516,N_9101);
nand UO_30 (O_30,N_9565,N_9661);
nand UO_31 (O_31,N_9080,N_9602);
nand UO_32 (O_32,N_9646,N_9541);
and UO_33 (O_33,N_9053,N_9043);
or UO_34 (O_34,N_9155,N_9977);
xnor UO_35 (O_35,N_9417,N_9032);
nand UO_36 (O_36,N_9454,N_9613);
xor UO_37 (O_37,N_9508,N_9416);
nor UO_38 (O_38,N_9714,N_9440);
nor UO_39 (O_39,N_9238,N_9501);
and UO_40 (O_40,N_9536,N_9148);
nand UO_41 (O_41,N_9578,N_9256);
nor UO_42 (O_42,N_9874,N_9751);
nor UO_43 (O_43,N_9514,N_9425);
nand UO_44 (O_44,N_9112,N_9084);
or UO_45 (O_45,N_9544,N_9227);
xnor UO_46 (O_46,N_9384,N_9311);
nand UO_47 (O_47,N_9243,N_9066);
nor UO_48 (O_48,N_9444,N_9722);
nor UO_49 (O_49,N_9670,N_9415);
or UO_50 (O_50,N_9120,N_9756);
nand UO_51 (O_51,N_9249,N_9269);
nor UO_52 (O_52,N_9363,N_9209);
nor UO_53 (O_53,N_9930,N_9401);
or UO_54 (O_54,N_9164,N_9442);
nor UO_55 (O_55,N_9147,N_9764);
or UO_56 (O_56,N_9435,N_9740);
nor UO_57 (O_57,N_9498,N_9446);
nor UO_58 (O_58,N_9064,N_9470);
nand UO_59 (O_59,N_9506,N_9608);
or UO_60 (O_60,N_9889,N_9377);
and UO_61 (O_61,N_9046,N_9932);
or UO_62 (O_62,N_9070,N_9582);
xor UO_63 (O_63,N_9898,N_9847);
or UO_64 (O_64,N_9995,N_9037);
nand UO_65 (O_65,N_9494,N_9001);
xnor UO_66 (O_66,N_9944,N_9869);
and UO_67 (O_67,N_9459,N_9213);
or UO_68 (O_68,N_9585,N_9610);
and UO_69 (O_69,N_9719,N_9184);
xnor UO_70 (O_70,N_9093,N_9936);
or UO_71 (O_71,N_9653,N_9414);
nor UO_72 (O_72,N_9789,N_9838);
and UO_73 (O_73,N_9814,N_9021);
and UO_74 (O_74,N_9094,N_9810);
nor UO_75 (O_75,N_9018,N_9180);
or UO_76 (O_76,N_9839,N_9681);
nor UO_77 (O_77,N_9683,N_9150);
nand UO_78 (O_78,N_9781,N_9531);
xor UO_79 (O_79,N_9090,N_9012);
and UO_80 (O_80,N_9752,N_9696);
or UO_81 (O_81,N_9010,N_9011);
or UO_82 (O_82,N_9423,N_9629);
nor UO_83 (O_83,N_9062,N_9518);
nand UO_84 (O_84,N_9822,N_9845);
or UO_85 (O_85,N_9100,N_9928);
xnor UO_86 (O_86,N_9014,N_9281);
nand UO_87 (O_87,N_9475,N_9405);
nand UO_88 (O_88,N_9149,N_9689);
nand UO_89 (O_89,N_9702,N_9123);
and UO_90 (O_90,N_9165,N_9892);
nor UO_91 (O_91,N_9618,N_9463);
and UO_92 (O_92,N_9016,N_9589);
or UO_93 (O_93,N_9154,N_9717);
nor UO_94 (O_94,N_9412,N_9085);
nor UO_95 (O_95,N_9404,N_9774);
nand UO_96 (O_96,N_9598,N_9611);
and UO_97 (O_97,N_9260,N_9476);
nor UO_98 (O_98,N_9586,N_9744);
xor UO_99 (O_99,N_9366,N_9904);
or UO_100 (O_100,N_9286,N_9590);
nor UO_101 (O_101,N_9132,N_9153);
or UO_102 (O_102,N_9335,N_9946);
or UO_103 (O_103,N_9216,N_9189);
and UO_104 (O_104,N_9757,N_9220);
and UO_105 (O_105,N_9305,N_9102);
nor UO_106 (O_106,N_9929,N_9663);
or UO_107 (O_107,N_9786,N_9246);
nand UO_108 (O_108,N_9262,N_9041);
or UO_109 (O_109,N_9142,N_9829);
nand UO_110 (O_110,N_9357,N_9020);
nand UO_111 (O_111,N_9002,N_9739);
nor UO_112 (O_112,N_9901,N_9821);
nor UO_113 (O_113,N_9293,N_9096);
or UO_114 (O_114,N_9346,N_9251);
and UO_115 (O_115,N_9315,N_9772);
xnor UO_116 (O_116,N_9700,N_9073);
nor UO_117 (O_117,N_9467,N_9560);
nand UO_118 (O_118,N_9226,N_9283);
or UO_119 (O_119,N_9171,N_9382);
nor UO_120 (O_120,N_9489,N_9524);
xor UO_121 (O_121,N_9354,N_9051);
nand UO_122 (O_122,N_9999,N_9274);
or UO_123 (O_123,N_9979,N_9833);
and UO_124 (O_124,N_9206,N_9665);
or UO_125 (O_125,N_9538,N_9801);
or UO_126 (O_126,N_9701,N_9919);
or UO_127 (O_127,N_9818,N_9909);
or UO_128 (O_128,N_9997,N_9430);
and UO_129 (O_129,N_9658,N_9135);
nor UO_130 (O_130,N_9044,N_9968);
nand UO_131 (O_131,N_9368,N_9673);
nor UO_132 (O_132,N_9609,N_9765);
or UO_133 (O_133,N_9107,N_9439);
and UO_134 (O_134,N_9499,N_9873);
or UO_135 (O_135,N_9923,N_9277);
or UO_136 (O_136,N_9452,N_9854);
or UO_137 (O_137,N_9397,N_9219);
and UO_138 (O_138,N_9694,N_9978);
xor UO_139 (O_139,N_9513,N_9174);
nand UO_140 (O_140,N_9308,N_9706);
nand UO_141 (O_141,N_9965,N_9761);
nor UO_142 (O_142,N_9421,N_9119);
and UO_143 (O_143,N_9742,N_9324);
or UO_144 (O_144,N_9160,N_9278);
or UO_145 (O_145,N_9607,N_9144);
nor UO_146 (O_146,N_9299,N_9647);
nand UO_147 (O_147,N_9688,N_9481);
nor UO_148 (O_148,N_9623,N_9592);
or UO_149 (O_149,N_9852,N_9556);
nor UO_150 (O_150,N_9849,N_9985);
or UO_151 (O_151,N_9321,N_9035);
nor UO_152 (O_152,N_9614,N_9922);
nand UO_153 (O_153,N_9325,N_9850);
nor UO_154 (O_154,N_9285,N_9802);
nand UO_155 (O_155,N_9167,N_9895);
xor UO_156 (O_156,N_9581,N_9782);
or UO_157 (O_157,N_9369,N_9819);
and UO_158 (O_158,N_9125,N_9455);
nand UO_159 (O_159,N_9179,N_9078);
nand UO_160 (O_160,N_9803,N_9908);
nor UO_161 (O_161,N_9191,N_9334);
nor UO_162 (O_162,N_9076,N_9272);
nor UO_163 (O_163,N_9199,N_9236);
nor UO_164 (O_164,N_9034,N_9783);
xnor UO_165 (O_165,N_9356,N_9104);
and UO_166 (O_166,N_9773,N_9047);
nor UO_167 (O_167,N_9955,N_9151);
and UO_168 (O_168,N_9679,N_9329);
or UO_169 (O_169,N_9519,N_9413);
xor UO_170 (O_170,N_9040,N_9079);
nor UO_171 (O_171,N_9996,N_9925);
nor UO_172 (O_172,N_9579,N_9370);
nand UO_173 (O_173,N_9450,N_9660);
nor UO_174 (O_174,N_9250,N_9115);
or UO_175 (O_175,N_9254,N_9309);
nor UO_176 (O_176,N_9264,N_9126);
nand UO_177 (O_177,N_9622,N_9350);
and UO_178 (O_178,N_9987,N_9728);
or UO_179 (O_179,N_9716,N_9193);
nand UO_180 (O_180,N_9162,N_9795);
or UO_181 (O_181,N_9616,N_9509);
and UO_182 (O_182,N_9641,N_9828);
or UO_183 (O_183,N_9958,N_9320);
nor UO_184 (O_184,N_9619,N_9460);
nor UO_185 (O_185,N_9059,N_9279);
nand UO_186 (O_186,N_9668,N_9548);
nand UO_187 (O_187,N_9240,N_9403);
nand UO_188 (O_188,N_9464,N_9072);
nor UO_189 (O_189,N_9883,N_9723);
and UO_190 (O_190,N_9832,N_9143);
nor UO_191 (O_191,N_9737,N_9750);
or UO_192 (O_192,N_9022,N_9626);
nor UO_193 (O_193,N_9339,N_9811);
xnor UO_194 (O_194,N_9634,N_9826);
nor UO_195 (O_195,N_9344,N_9291);
nor UO_196 (O_196,N_9768,N_9310);
or UO_197 (O_197,N_9082,N_9915);
nor UO_198 (O_198,N_9594,N_9593);
or UO_199 (O_199,N_9878,N_9157);
nand UO_200 (O_200,N_9961,N_9492);
nand UO_201 (O_201,N_9201,N_9190);
nand UO_202 (O_202,N_9232,N_9834);
and UO_203 (O_203,N_9225,N_9746);
or UO_204 (O_204,N_9025,N_9307);
nand UO_205 (O_205,N_9083,N_9615);
and UO_206 (O_206,N_9606,N_9715);
and UO_207 (O_207,N_9758,N_9228);
nand UO_208 (O_208,N_9888,N_9116);
or UO_209 (O_209,N_9437,N_9815);
nand UO_210 (O_210,N_9303,N_9292);
and UO_211 (O_211,N_9974,N_9632);
and UO_212 (O_212,N_9378,N_9557);
nand UO_213 (O_213,N_9848,N_9205);
nor UO_214 (O_214,N_9420,N_9948);
or UO_215 (O_215,N_9526,N_9515);
nand UO_216 (O_216,N_9584,N_9337);
nand UO_217 (O_217,N_9872,N_9994);
nand UO_218 (O_218,N_9825,N_9316);
and UO_219 (O_219,N_9091,N_9328);
or UO_220 (O_220,N_9234,N_9966);
nor UO_221 (O_221,N_9255,N_9379);
or UO_222 (O_222,N_9559,N_9237);
nand UO_223 (O_223,N_9488,N_9890);
nand UO_224 (O_224,N_9657,N_9648);
and UO_225 (O_225,N_9669,N_9671);
and UO_226 (O_226,N_9755,N_9788);
xnor UO_227 (O_227,N_9859,N_9807);
or UO_228 (O_228,N_9468,N_9937);
or UO_229 (O_229,N_9759,N_9990);
and UO_230 (O_230,N_9068,N_9345);
nand UO_231 (O_231,N_9418,N_9857);
nand UO_232 (O_232,N_9860,N_9398);
nand UO_233 (O_233,N_9218,N_9945);
and UO_234 (O_234,N_9336,N_9196);
and UO_235 (O_235,N_9884,N_9709);
nor UO_236 (O_236,N_9798,N_9124);
nor UO_237 (O_237,N_9270,N_9229);
and UO_238 (O_238,N_9141,N_9731);
xor UO_239 (O_239,N_9482,N_9804);
nand UO_240 (O_240,N_9621,N_9779);
or UO_241 (O_241,N_9882,N_9267);
nor UO_242 (O_242,N_9282,N_9207);
and UO_243 (O_243,N_9362,N_9263);
or UO_244 (O_244,N_9732,N_9175);
nand UO_245 (O_245,N_9241,N_9790);
and UO_246 (O_246,N_9776,N_9067);
and UO_247 (O_247,N_9003,N_9187);
or UO_248 (O_248,N_9982,N_9527);
nor UO_249 (O_249,N_9649,N_9957);
nand UO_250 (O_250,N_9451,N_9865);
nand UO_251 (O_251,N_9676,N_9131);
and UO_252 (O_252,N_9323,N_9654);
or UO_253 (O_253,N_9298,N_9917);
xnor UO_254 (O_254,N_9631,N_9485);
nand UO_255 (O_255,N_9549,N_9914);
nand UO_256 (O_256,N_9726,N_9659);
nand UO_257 (O_257,N_9698,N_9521);
nor UO_258 (O_258,N_9760,N_9941);
nor UO_259 (O_259,N_9351,N_9113);
and UO_260 (O_260,N_9920,N_9972);
or UO_261 (O_261,N_9695,N_9092);
xnor UO_262 (O_262,N_9396,N_9312);
nor UO_263 (O_263,N_9372,N_9169);
nand UO_264 (O_264,N_9666,N_9729);
and UO_265 (O_265,N_9458,N_9371);
and UO_266 (O_266,N_9152,N_9926);
nor UO_267 (O_267,N_9806,N_9745);
nor UO_268 (O_268,N_9712,N_9387);
xnor UO_269 (O_269,N_9170,N_9655);
nand UO_270 (O_270,N_9880,N_9261);
nor UO_271 (O_271,N_9692,N_9741);
and UO_272 (O_272,N_9708,N_9831);
and UO_273 (O_273,N_9749,N_9449);
nor UO_274 (O_274,N_9938,N_9099);
and UO_275 (O_275,N_9503,N_9562);
or UO_276 (O_276,N_9287,N_9603);
xor UO_277 (O_277,N_9678,N_9574);
nand UO_278 (O_278,N_9984,N_9886);
or UO_279 (O_279,N_9525,N_9894);
and UO_280 (O_280,N_9844,N_9636);
nand UO_281 (O_281,N_9231,N_9887);
nor UO_282 (O_282,N_9951,N_9953);
or UO_283 (O_283,N_9029,N_9624);
or UO_284 (O_284,N_9642,N_9036);
and UO_285 (O_285,N_9258,N_9704);
and UO_286 (O_286,N_9870,N_9400);
and UO_287 (O_287,N_9973,N_9088);
nand UO_288 (O_288,N_9257,N_9058);
and UO_289 (O_289,N_9991,N_9122);
nor UO_290 (O_290,N_9591,N_9855);
or UO_291 (O_291,N_9302,N_9338);
or UO_292 (O_292,N_9322,N_9568);
or UO_293 (O_293,N_9472,N_9434);
nand UO_294 (O_294,N_9546,N_9381);
and UO_295 (O_295,N_9358,N_9841);
or UO_296 (O_296,N_9478,N_9097);
and UO_297 (O_297,N_9049,N_9600);
nand UO_298 (O_298,N_9791,N_9461);
nand UO_299 (O_299,N_9332,N_9637);
nand UO_300 (O_300,N_9327,N_9800);
xor UO_301 (O_301,N_9300,N_9331);
and UO_302 (O_302,N_9563,N_9754);
nand UO_303 (O_303,N_9504,N_9724);
nor UO_304 (O_304,N_9333,N_9612);
or UO_305 (O_305,N_9419,N_9426);
nor UO_306 (O_306,N_9364,N_9597);
nand UO_307 (O_307,N_9071,N_9993);
or UO_308 (O_308,N_9436,N_9939);
nor UO_309 (O_309,N_9490,N_9496);
nor UO_310 (O_310,N_9348,N_9510);
nand UO_311 (O_311,N_9052,N_9547);
or UO_312 (O_312,N_9317,N_9522);
nand UO_313 (O_313,N_9711,N_9964);
and UO_314 (O_314,N_9137,N_9656);
nor UO_315 (O_315,N_9778,N_9129);
xor UO_316 (O_316,N_9667,N_9075);
xnor UO_317 (O_317,N_9820,N_9542);
nor UO_318 (O_318,N_9583,N_9484);
or UO_319 (O_319,N_9794,N_9858);
nor UO_320 (O_320,N_9156,N_9587);
nand UO_321 (O_321,N_9087,N_9687);
and UO_322 (O_322,N_9395,N_9388);
or UO_323 (O_323,N_9359,N_9026);
xor UO_324 (O_324,N_9893,N_9159);
xnor UO_325 (O_325,N_9447,N_9114);
and UO_326 (O_326,N_9899,N_9195);
or UO_327 (O_327,N_9952,N_9730);
or UO_328 (O_328,N_9896,N_9736);
xnor UO_329 (O_329,N_9856,N_9176);
nand UO_330 (O_330,N_9391,N_9000);
and UO_331 (O_331,N_9375,N_9863);
and UO_332 (O_332,N_9644,N_9106);
xnor UO_333 (O_333,N_9265,N_9743);
nor UO_334 (O_334,N_9373,N_9523);
nor UO_335 (O_335,N_9707,N_9500);
nor UO_336 (O_336,N_9424,N_9009);
nor UO_337 (O_337,N_9787,N_9208);
nand UO_338 (O_338,N_9314,N_9551);
nor UO_339 (O_339,N_9770,N_9564);
or UO_340 (O_340,N_9005,N_9897);
or UO_341 (O_341,N_9431,N_9198);
nor UO_342 (O_342,N_9383,N_9428);
xnor UO_343 (O_343,N_9474,N_9048);
and UO_344 (O_344,N_9879,N_9203);
nand UO_345 (O_345,N_9089,N_9962);
nand UO_346 (O_346,N_9060,N_9975);
or UO_347 (O_347,N_9540,N_9318);
nand UO_348 (O_348,N_9573,N_9816);
nor UO_349 (O_349,N_9921,N_9853);
nand UO_350 (O_350,N_9477,N_9588);
and UO_351 (O_351,N_9469,N_9493);
or UO_352 (O_352,N_9306,N_9617);
or UO_353 (O_353,N_9605,N_9224);
nand UO_354 (O_354,N_9399,N_9843);
nand UO_355 (O_355,N_9462,N_9045);
nand UO_356 (O_356,N_9215,N_9223);
nor UO_357 (O_357,N_9824,N_9296);
or UO_358 (O_358,N_9360,N_9271);
nor UO_359 (O_359,N_9146,N_9480);
nor UO_360 (O_360,N_9192,N_9577);
nand UO_361 (O_361,N_9214,N_9081);
xor UO_362 (O_362,N_9409,N_9685);
or UO_363 (O_363,N_9652,N_9567);
and UO_364 (O_364,N_9030,N_9927);
nand UO_365 (O_365,N_9466,N_9949);
nand UO_366 (O_366,N_9110,N_9024);
xnor UO_367 (O_367,N_9545,N_9221);
nor UO_368 (O_368,N_9386,N_9520);
nand UO_369 (O_369,N_9956,N_9868);
or UO_370 (O_370,N_9569,N_9491);
or UO_371 (O_371,N_9507,N_9342);
and UO_372 (O_372,N_9866,N_9969);
and UO_373 (O_373,N_9862,N_9916);
or UO_374 (O_374,N_9771,N_9677);
or UO_375 (O_375,N_9039,N_9502);
nand UO_376 (O_376,N_9197,N_9903);
and UO_377 (O_377,N_9077,N_9103);
or UO_378 (O_378,N_9202,N_9572);
nor UO_379 (O_379,N_9235,N_9233);
nand UO_380 (O_380,N_9942,N_9947);
nor UO_381 (O_381,N_9343,N_9552);
nand UO_382 (O_382,N_9861,N_9628);
nor UO_383 (O_383,N_9762,N_9109);
nand UO_384 (O_384,N_9906,N_9266);
or UO_385 (O_385,N_9033,N_9133);
xnor UO_386 (O_386,N_9121,N_9433);
and UO_387 (O_387,N_9885,N_9517);
or UO_388 (O_388,N_9830,N_9686);
nor UO_389 (O_389,N_9988,N_9422);
nand UO_390 (O_390,N_9289,N_9127);
and UO_391 (O_391,N_9630,N_9840);
and UO_392 (O_392,N_9604,N_9313);
or UO_393 (O_393,N_9330,N_9705);
nand UO_394 (O_394,N_9487,N_9367);
nand UO_395 (O_395,N_9050,N_9057);
nor UO_396 (O_396,N_9891,N_9633);
nand UO_397 (O_397,N_9963,N_9352);
and UO_398 (O_398,N_9355,N_9554);
nor UO_399 (O_399,N_9211,N_9836);
and UO_400 (O_400,N_9134,N_9471);
nor UO_401 (O_401,N_9341,N_9456);
nor UO_402 (O_402,N_9753,N_9505);
nand UO_403 (O_403,N_9411,N_9069);
or UO_404 (O_404,N_9183,N_9473);
and UO_405 (O_405,N_9620,N_9017);
nor UO_406 (O_406,N_9640,N_9835);
or UO_407 (O_407,N_9108,N_9534);
xnor UO_408 (O_408,N_9443,N_9407);
and UO_409 (O_409,N_9913,N_9775);
or UO_410 (O_410,N_9748,N_9376);
and UO_411 (O_411,N_9900,N_9651);
nor UO_412 (O_412,N_9304,N_9576);
nand UO_413 (O_413,N_9074,N_9242);
or UO_414 (O_414,N_9738,N_9319);
nor UO_415 (O_415,N_9643,N_9284);
and UO_416 (O_416,N_9182,N_9027);
and UO_417 (O_417,N_9349,N_9217);
nand UO_418 (O_418,N_9275,N_9511);
and UO_419 (O_419,N_9495,N_9983);
or UO_420 (O_420,N_9867,N_9163);
and UO_421 (O_421,N_9970,N_9599);
or UO_422 (O_422,N_9902,N_9280);
nand UO_423 (O_423,N_9539,N_9239);
and UO_424 (O_424,N_9252,N_9380);
and UO_425 (O_425,N_9796,N_9532);
nand UO_426 (O_426,N_9672,N_9967);
nand UO_427 (O_427,N_9943,N_9596);
nand UO_428 (O_428,N_9168,N_9161);
nor UO_429 (O_429,N_9777,N_9797);
nor UO_430 (O_430,N_9145,N_9347);
or UO_431 (O_431,N_9940,N_9725);
nand UO_432 (O_432,N_9086,N_9483);
or UO_433 (O_433,N_9301,N_9245);
and UO_434 (O_434,N_9986,N_9645);
or UO_435 (O_435,N_9055,N_9699);
nor UO_436 (O_436,N_9276,N_9054);
nand UO_437 (O_437,N_9784,N_9924);
nor UO_438 (O_438,N_9733,N_9138);
or UO_439 (O_439,N_9555,N_9735);
and UO_440 (O_440,N_9056,N_9512);
and UO_441 (O_441,N_9105,N_9992);
or UO_442 (O_442,N_9065,N_9326);
and UO_443 (O_443,N_9817,N_9805);
nor UO_444 (O_444,N_9031,N_9340);
and UO_445 (O_445,N_9785,N_9465);
nor UO_446 (O_446,N_9529,N_9410);
and UO_447 (O_447,N_9186,N_9959);
and UO_448 (O_448,N_9393,N_9543);
xor UO_449 (O_449,N_9809,N_9389);
nor UO_450 (O_450,N_9268,N_9934);
nand UO_451 (O_451,N_9989,N_9248);
or UO_452 (O_452,N_9172,N_9960);
nor UO_453 (O_453,N_9703,N_9980);
nor UO_454 (O_454,N_9061,N_9128);
and UO_455 (O_455,N_9595,N_9998);
nor UO_456 (O_456,N_9639,N_9718);
and UO_457 (O_457,N_9200,N_9918);
and UO_458 (O_458,N_9166,N_9950);
nand UO_459 (O_459,N_9550,N_9290);
or UO_460 (O_460,N_9259,N_9808);
nand UO_461 (O_461,N_9911,N_9910);
and UO_462 (O_462,N_9139,N_9691);
nor UO_463 (O_463,N_9625,N_9780);
nor UO_464 (O_464,N_9601,N_9402);
nor UO_465 (O_465,N_9008,N_9288);
nand UO_466 (O_466,N_9006,N_9385);
nor UO_467 (O_467,N_9682,N_9353);
nor UO_468 (O_468,N_9697,N_9837);
or UO_469 (O_469,N_9793,N_9638);
nand UO_470 (O_470,N_9297,N_9570);
nand UO_471 (O_471,N_9675,N_9561);
xnor UO_472 (O_472,N_9095,N_9662);
or UO_473 (O_473,N_9394,N_9457);
nand UO_474 (O_474,N_9194,N_9727);
and UO_475 (O_475,N_9827,N_9680);
xnor UO_476 (O_476,N_9173,N_9693);
nand UO_477 (O_477,N_9273,N_9117);
or UO_478 (O_478,N_9023,N_9981);
nor UO_479 (O_479,N_9813,N_9713);
or UO_480 (O_480,N_9015,N_9432);
and UO_481 (O_481,N_9429,N_9185);
xor UO_482 (O_482,N_9864,N_9537);
or UO_483 (O_483,N_9479,N_9448);
nand UO_484 (O_484,N_9222,N_9177);
and UO_485 (O_485,N_9212,N_9575);
and UO_486 (O_486,N_9763,N_9792);
or UO_487 (O_487,N_9971,N_9019);
or UO_488 (O_488,N_9690,N_9734);
and UO_489 (O_489,N_9007,N_9111);
nor UO_490 (O_490,N_9042,N_9408);
or UO_491 (O_491,N_9253,N_9004);
nor UO_492 (O_492,N_9130,N_9374);
or UO_493 (O_493,N_9931,N_9445);
or UO_494 (O_494,N_9905,N_9392);
xor UO_495 (O_495,N_9767,N_9881);
xor UO_496 (O_496,N_9535,N_9294);
and UO_497 (O_497,N_9954,N_9230);
or UO_498 (O_498,N_9390,N_9136);
xor UO_499 (O_499,N_9441,N_9842);
nor UO_500 (O_500,N_9814,N_9424);
nor UO_501 (O_501,N_9005,N_9113);
or UO_502 (O_502,N_9413,N_9556);
and UO_503 (O_503,N_9010,N_9125);
nand UO_504 (O_504,N_9203,N_9389);
and UO_505 (O_505,N_9615,N_9624);
nor UO_506 (O_506,N_9747,N_9717);
nor UO_507 (O_507,N_9641,N_9904);
xor UO_508 (O_508,N_9234,N_9717);
or UO_509 (O_509,N_9707,N_9723);
nor UO_510 (O_510,N_9682,N_9720);
xor UO_511 (O_511,N_9004,N_9570);
xnor UO_512 (O_512,N_9828,N_9405);
and UO_513 (O_513,N_9824,N_9036);
nand UO_514 (O_514,N_9219,N_9075);
and UO_515 (O_515,N_9164,N_9683);
nor UO_516 (O_516,N_9310,N_9958);
xor UO_517 (O_517,N_9215,N_9010);
and UO_518 (O_518,N_9557,N_9925);
nand UO_519 (O_519,N_9371,N_9805);
nor UO_520 (O_520,N_9338,N_9190);
nor UO_521 (O_521,N_9653,N_9875);
or UO_522 (O_522,N_9919,N_9252);
and UO_523 (O_523,N_9166,N_9085);
xnor UO_524 (O_524,N_9021,N_9956);
or UO_525 (O_525,N_9921,N_9888);
nand UO_526 (O_526,N_9671,N_9265);
nor UO_527 (O_527,N_9836,N_9574);
nor UO_528 (O_528,N_9030,N_9586);
or UO_529 (O_529,N_9347,N_9558);
nand UO_530 (O_530,N_9372,N_9791);
nand UO_531 (O_531,N_9782,N_9977);
and UO_532 (O_532,N_9903,N_9777);
nand UO_533 (O_533,N_9860,N_9417);
and UO_534 (O_534,N_9321,N_9016);
xor UO_535 (O_535,N_9274,N_9123);
xnor UO_536 (O_536,N_9038,N_9639);
nand UO_537 (O_537,N_9827,N_9117);
xnor UO_538 (O_538,N_9918,N_9704);
and UO_539 (O_539,N_9720,N_9149);
and UO_540 (O_540,N_9477,N_9554);
or UO_541 (O_541,N_9883,N_9125);
nand UO_542 (O_542,N_9736,N_9310);
nand UO_543 (O_543,N_9259,N_9072);
nor UO_544 (O_544,N_9688,N_9279);
and UO_545 (O_545,N_9298,N_9713);
and UO_546 (O_546,N_9915,N_9614);
or UO_547 (O_547,N_9170,N_9488);
or UO_548 (O_548,N_9291,N_9948);
nor UO_549 (O_549,N_9020,N_9412);
and UO_550 (O_550,N_9456,N_9805);
or UO_551 (O_551,N_9464,N_9199);
or UO_552 (O_552,N_9212,N_9485);
or UO_553 (O_553,N_9146,N_9922);
and UO_554 (O_554,N_9356,N_9483);
nor UO_555 (O_555,N_9420,N_9702);
and UO_556 (O_556,N_9801,N_9132);
and UO_557 (O_557,N_9385,N_9470);
nor UO_558 (O_558,N_9618,N_9038);
and UO_559 (O_559,N_9275,N_9639);
xnor UO_560 (O_560,N_9148,N_9421);
nor UO_561 (O_561,N_9665,N_9520);
nor UO_562 (O_562,N_9818,N_9123);
or UO_563 (O_563,N_9565,N_9692);
xor UO_564 (O_564,N_9206,N_9362);
and UO_565 (O_565,N_9617,N_9639);
or UO_566 (O_566,N_9744,N_9542);
and UO_567 (O_567,N_9723,N_9286);
nand UO_568 (O_568,N_9551,N_9240);
or UO_569 (O_569,N_9092,N_9320);
nand UO_570 (O_570,N_9763,N_9464);
nand UO_571 (O_571,N_9120,N_9084);
and UO_572 (O_572,N_9581,N_9630);
xor UO_573 (O_573,N_9642,N_9241);
nor UO_574 (O_574,N_9942,N_9841);
xnor UO_575 (O_575,N_9074,N_9960);
xnor UO_576 (O_576,N_9683,N_9608);
nor UO_577 (O_577,N_9687,N_9516);
and UO_578 (O_578,N_9064,N_9066);
and UO_579 (O_579,N_9952,N_9448);
nor UO_580 (O_580,N_9629,N_9771);
nand UO_581 (O_581,N_9400,N_9334);
nor UO_582 (O_582,N_9479,N_9713);
or UO_583 (O_583,N_9616,N_9762);
nor UO_584 (O_584,N_9844,N_9617);
nor UO_585 (O_585,N_9822,N_9584);
or UO_586 (O_586,N_9970,N_9893);
nor UO_587 (O_587,N_9749,N_9739);
nor UO_588 (O_588,N_9593,N_9908);
and UO_589 (O_589,N_9867,N_9004);
or UO_590 (O_590,N_9215,N_9858);
and UO_591 (O_591,N_9516,N_9405);
and UO_592 (O_592,N_9139,N_9939);
xor UO_593 (O_593,N_9772,N_9065);
and UO_594 (O_594,N_9608,N_9661);
or UO_595 (O_595,N_9320,N_9091);
and UO_596 (O_596,N_9387,N_9431);
or UO_597 (O_597,N_9894,N_9847);
nor UO_598 (O_598,N_9099,N_9574);
and UO_599 (O_599,N_9900,N_9391);
nand UO_600 (O_600,N_9175,N_9164);
or UO_601 (O_601,N_9514,N_9270);
and UO_602 (O_602,N_9383,N_9349);
nor UO_603 (O_603,N_9631,N_9929);
nor UO_604 (O_604,N_9726,N_9850);
and UO_605 (O_605,N_9662,N_9911);
nand UO_606 (O_606,N_9973,N_9101);
and UO_607 (O_607,N_9084,N_9744);
nand UO_608 (O_608,N_9451,N_9064);
nand UO_609 (O_609,N_9165,N_9993);
or UO_610 (O_610,N_9412,N_9951);
nor UO_611 (O_611,N_9256,N_9753);
xnor UO_612 (O_612,N_9345,N_9650);
or UO_613 (O_613,N_9851,N_9024);
and UO_614 (O_614,N_9521,N_9301);
or UO_615 (O_615,N_9837,N_9790);
nor UO_616 (O_616,N_9197,N_9473);
xnor UO_617 (O_617,N_9621,N_9370);
or UO_618 (O_618,N_9455,N_9274);
xnor UO_619 (O_619,N_9927,N_9015);
or UO_620 (O_620,N_9715,N_9328);
xnor UO_621 (O_621,N_9419,N_9159);
and UO_622 (O_622,N_9948,N_9317);
xnor UO_623 (O_623,N_9179,N_9137);
and UO_624 (O_624,N_9304,N_9442);
nand UO_625 (O_625,N_9288,N_9311);
nand UO_626 (O_626,N_9059,N_9371);
nor UO_627 (O_627,N_9386,N_9043);
nand UO_628 (O_628,N_9591,N_9202);
nor UO_629 (O_629,N_9749,N_9669);
and UO_630 (O_630,N_9383,N_9997);
xnor UO_631 (O_631,N_9611,N_9833);
or UO_632 (O_632,N_9730,N_9988);
or UO_633 (O_633,N_9049,N_9353);
nand UO_634 (O_634,N_9183,N_9998);
and UO_635 (O_635,N_9530,N_9954);
or UO_636 (O_636,N_9739,N_9114);
xor UO_637 (O_637,N_9504,N_9621);
or UO_638 (O_638,N_9591,N_9543);
nor UO_639 (O_639,N_9362,N_9140);
nand UO_640 (O_640,N_9203,N_9235);
nand UO_641 (O_641,N_9392,N_9112);
or UO_642 (O_642,N_9810,N_9404);
nor UO_643 (O_643,N_9729,N_9829);
xnor UO_644 (O_644,N_9136,N_9857);
xnor UO_645 (O_645,N_9053,N_9809);
or UO_646 (O_646,N_9496,N_9961);
and UO_647 (O_647,N_9757,N_9176);
xor UO_648 (O_648,N_9778,N_9016);
nor UO_649 (O_649,N_9976,N_9831);
nor UO_650 (O_650,N_9167,N_9215);
nor UO_651 (O_651,N_9261,N_9572);
and UO_652 (O_652,N_9388,N_9687);
nor UO_653 (O_653,N_9971,N_9618);
xnor UO_654 (O_654,N_9660,N_9031);
nor UO_655 (O_655,N_9564,N_9403);
nor UO_656 (O_656,N_9815,N_9624);
and UO_657 (O_657,N_9747,N_9921);
and UO_658 (O_658,N_9367,N_9186);
xnor UO_659 (O_659,N_9231,N_9430);
and UO_660 (O_660,N_9747,N_9644);
nand UO_661 (O_661,N_9408,N_9856);
and UO_662 (O_662,N_9018,N_9222);
xnor UO_663 (O_663,N_9162,N_9646);
nor UO_664 (O_664,N_9660,N_9629);
xnor UO_665 (O_665,N_9736,N_9175);
or UO_666 (O_666,N_9282,N_9041);
nor UO_667 (O_667,N_9120,N_9722);
nand UO_668 (O_668,N_9036,N_9431);
and UO_669 (O_669,N_9187,N_9063);
nand UO_670 (O_670,N_9556,N_9392);
or UO_671 (O_671,N_9757,N_9311);
xnor UO_672 (O_672,N_9024,N_9523);
nand UO_673 (O_673,N_9071,N_9920);
or UO_674 (O_674,N_9237,N_9653);
nor UO_675 (O_675,N_9112,N_9460);
or UO_676 (O_676,N_9383,N_9615);
or UO_677 (O_677,N_9175,N_9140);
xor UO_678 (O_678,N_9241,N_9260);
and UO_679 (O_679,N_9064,N_9450);
nand UO_680 (O_680,N_9056,N_9803);
nand UO_681 (O_681,N_9454,N_9540);
nor UO_682 (O_682,N_9102,N_9257);
nor UO_683 (O_683,N_9561,N_9968);
and UO_684 (O_684,N_9289,N_9128);
xor UO_685 (O_685,N_9654,N_9231);
and UO_686 (O_686,N_9524,N_9898);
nor UO_687 (O_687,N_9089,N_9984);
nor UO_688 (O_688,N_9425,N_9731);
and UO_689 (O_689,N_9040,N_9781);
or UO_690 (O_690,N_9803,N_9005);
nor UO_691 (O_691,N_9471,N_9076);
and UO_692 (O_692,N_9132,N_9998);
or UO_693 (O_693,N_9829,N_9082);
xor UO_694 (O_694,N_9684,N_9341);
nand UO_695 (O_695,N_9124,N_9464);
nand UO_696 (O_696,N_9718,N_9732);
xnor UO_697 (O_697,N_9778,N_9433);
or UO_698 (O_698,N_9504,N_9119);
nor UO_699 (O_699,N_9171,N_9647);
nand UO_700 (O_700,N_9521,N_9768);
and UO_701 (O_701,N_9851,N_9240);
nand UO_702 (O_702,N_9279,N_9577);
and UO_703 (O_703,N_9050,N_9926);
nor UO_704 (O_704,N_9687,N_9076);
nor UO_705 (O_705,N_9039,N_9810);
or UO_706 (O_706,N_9937,N_9140);
nor UO_707 (O_707,N_9420,N_9529);
nor UO_708 (O_708,N_9169,N_9240);
nor UO_709 (O_709,N_9826,N_9641);
nand UO_710 (O_710,N_9339,N_9395);
and UO_711 (O_711,N_9374,N_9395);
or UO_712 (O_712,N_9796,N_9411);
or UO_713 (O_713,N_9701,N_9518);
or UO_714 (O_714,N_9799,N_9659);
xnor UO_715 (O_715,N_9888,N_9356);
nor UO_716 (O_716,N_9464,N_9614);
nor UO_717 (O_717,N_9091,N_9522);
or UO_718 (O_718,N_9244,N_9882);
nand UO_719 (O_719,N_9083,N_9495);
xor UO_720 (O_720,N_9391,N_9434);
or UO_721 (O_721,N_9820,N_9884);
xor UO_722 (O_722,N_9294,N_9963);
nor UO_723 (O_723,N_9359,N_9818);
or UO_724 (O_724,N_9792,N_9092);
nor UO_725 (O_725,N_9233,N_9524);
and UO_726 (O_726,N_9959,N_9835);
nor UO_727 (O_727,N_9253,N_9958);
nor UO_728 (O_728,N_9440,N_9315);
nand UO_729 (O_729,N_9298,N_9288);
or UO_730 (O_730,N_9544,N_9884);
or UO_731 (O_731,N_9908,N_9853);
or UO_732 (O_732,N_9929,N_9821);
nor UO_733 (O_733,N_9054,N_9137);
and UO_734 (O_734,N_9468,N_9826);
or UO_735 (O_735,N_9774,N_9287);
and UO_736 (O_736,N_9833,N_9433);
and UO_737 (O_737,N_9153,N_9366);
and UO_738 (O_738,N_9814,N_9615);
and UO_739 (O_739,N_9887,N_9493);
and UO_740 (O_740,N_9623,N_9555);
or UO_741 (O_741,N_9042,N_9493);
or UO_742 (O_742,N_9602,N_9748);
xor UO_743 (O_743,N_9756,N_9087);
and UO_744 (O_744,N_9702,N_9960);
nand UO_745 (O_745,N_9349,N_9040);
or UO_746 (O_746,N_9234,N_9677);
nand UO_747 (O_747,N_9666,N_9584);
nor UO_748 (O_748,N_9760,N_9858);
nor UO_749 (O_749,N_9991,N_9117);
or UO_750 (O_750,N_9294,N_9805);
nand UO_751 (O_751,N_9064,N_9554);
nand UO_752 (O_752,N_9977,N_9621);
or UO_753 (O_753,N_9533,N_9318);
xnor UO_754 (O_754,N_9804,N_9984);
or UO_755 (O_755,N_9646,N_9714);
nor UO_756 (O_756,N_9794,N_9180);
nand UO_757 (O_757,N_9277,N_9040);
and UO_758 (O_758,N_9470,N_9086);
or UO_759 (O_759,N_9242,N_9389);
xor UO_760 (O_760,N_9273,N_9906);
nor UO_761 (O_761,N_9290,N_9803);
nor UO_762 (O_762,N_9535,N_9059);
nand UO_763 (O_763,N_9233,N_9266);
nand UO_764 (O_764,N_9055,N_9868);
and UO_765 (O_765,N_9389,N_9845);
or UO_766 (O_766,N_9482,N_9031);
or UO_767 (O_767,N_9714,N_9382);
nand UO_768 (O_768,N_9098,N_9418);
and UO_769 (O_769,N_9951,N_9940);
or UO_770 (O_770,N_9727,N_9933);
nor UO_771 (O_771,N_9644,N_9466);
nand UO_772 (O_772,N_9664,N_9070);
and UO_773 (O_773,N_9064,N_9080);
nand UO_774 (O_774,N_9166,N_9513);
or UO_775 (O_775,N_9049,N_9950);
or UO_776 (O_776,N_9806,N_9994);
and UO_777 (O_777,N_9976,N_9041);
xnor UO_778 (O_778,N_9953,N_9126);
or UO_779 (O_779,N_9446,N_9507);
nor UO_780 (O_780,N_9185,N_9713);
nand UO_781 (O_781,N_9884,N_9965);
or UO_782 (O_782,N_9306,N_9371);
or UO_783 (O_783,N_9972,N_9125);
nor UO_784 (O_784,N_9846,N_9991);
and UO_785 (O_785,N_9546,N_9289);
or UO_786 (O_786,N_9362,N_9880);
nand UO_787 (O_787,N_9183,N_9655);
xnor UO_788 (O_788,N_9980,N_9100);
or UO_789 (O_789,N_9491,N_9005);
and UO_790 (O_790,N_9645,N_9574);
or UO_791 (O_791,N_9458,N_9712);
nand UO_792 (O_792,N_9101,N_9027);
and UO_793 (O_793,N_9001,N_9900);
nand UO_794 (O_794,N_9284,N_9956);
and UO_795 (O_795,N_9875,N_9209);
and UO_796 (O_796,N_9710,N_9971);
nor UO_797 (O_797,N_9218,N_9037);
nor UO_798 (O_798,N_9597,N_9271);
and UO_799 (O_799,N_9993,N_9747);
nor UO_800 (O_800,N_9067,N_9603);
or UO_801 (O_801,N_9496,N_9489);
xnor UO_802 (O_802,N_9184,N_9127);
or UO_803 (O_803,N_9334,N_9842);
nor UO_804 (O_804,N_9451,N_9911);
or UO_805 (O_805,N_9471,N_9446);
nor UO_806 (O_806,N_9504,N_9056);
and UO_807 (O_807,N_9418,N_9298);
and UO_808 (O_808,N_9010,N_9066);
nor UO_809 (O_809,N_9349,N_9471);
nand UO_810 (O_810,N_9537,N_9961);
and UO_811 (O_811,N_9594,N_9135);
and UO_812 (O_812,N_9377,N_9830);
nand UO_813 (O_813,N_9775,N_9965);
xnor UO_814 (O_814,N_9076,N_9680);
nand UO_815 (O_815,N_9347,N_9805);
and UO_816 (O_816,N_9975,N_9637);
or UO_817 (O_817,N_9544,N_9909);
xor UO_818 (O_818,N_9348,N_9779);
or UO_819 (O_819,N_9229,N_9146);
or UO_820 (O_820,N_9991,N_9242);
and UO_821 (O_821,N_9065,N_9089);
nand UO_822 (O_822,N_9572,N_9789);
nand UO_823 (O_823,N_9165,N_9023);
nand UO_824 (O_824,N_9883,N_9819);
nand UO_825 (O_825,N_9979,N_9303);
or UO_826 (O_826,N_9744,N_9925);
or UO_827 (O_827,N_9083,N_9753);
and UO_828 (O_828,N_9476,N_9935);
or UO_829 (O_829,N_9445,N_9081);
and UO_830 (O_830,N_9890,N_9107);
nor UO_831 (O_831,N_9422,N_9426);
nand UO_832 (O_832,N_9863,N_9469);
or UO_833 (O_833,N_9574,N_9705);
or UO_834 (O_834,N_9010,N_9343);
nand UO_835 (O_835,N_9321,N_9978);
nor UO_836 (O_836,N_9687,N_9910);
nor UO_837 (O_837,N_9845,N_9873);
or UO_838 (O_838,N_9208,N_9791);
nor UO_839 (O_839,N_9102,N_9921);
or UO_840 (O_840,N_9779,N_9802);
or UO_841 (O_841,N_9569,N_9379);
and UO_842 (O_842,N_9159,N_9115);
or UO_843 (O_843,N_9630,N_9648);
nand UO_844 (O_844,N_9330,N_9493);
and UO_845 (O_845,N_9175,N_9249);
xor UO_846 (O_846,N_9725,N_9363);
or UO_847 (O_847,N_9042,N_9393);
or UO_848 (O_848,N_9751,N_9893);
nor UO_849 (O_849,N_9160,N_9435);
nor UO_850 (O_850,N_9536,N_9796);
nand UO_851 (O_851,N_9759,N_9076);
and UO_852 (O_852,N_9084,N_9278);
and UO_853 (O_853,N_9143,N_9359);
or UO_854 (O_854,N_9889,N_9658);
and UO_855 (O_855,N_9576,N_9107);
nand UO_856 (O_856,N_9859,N_9735);
nor UO_857 (O_857,N_9579,N_9187);
nand UO_858 (O_858,N_9347,N_9133);
or UO_859 (O_859,N_9905,N_9486);
and UO_860 (O_860,N_9010,N_9243);
and UO_861 (O_861,N_9683,N_9651);
and UO_862 (O_862,N_9971,N_9438);
and UO_863 (O_863,N_9128,N_9303);
or UO_864 (O_864,N_9611,N_9067);
or UO_865 (O_865,N_9850,N_9591);
or UO_866 (O_866,N_9405,N_9930);
or UO_867 (O_867,N_9049,N_9136);
or UO_868 (O_868,N_9234,N_9109);
nand UO_869 (O_869,N_9921,N_9820);
xnor UO_870 (O_870,N_9899,N_9383);
and UO_871 (O_871,N_9645,N_9532);
or UO_872 (O_872,N_9485,N_9315);
or UO_873 (O_873,N_9668,N_9728);
xnor UO_874 (O_874,N_9776,N_9405);
nand UO_875 (O_875,N_9523,N_9759);
nor UO_876 (O_876,N_9316,N_9189);
nor UO_877 (O_877,N_9608,N_9216);
and UO_878 (O_878,N_9619,N_9122);
nand UO_879 (O_879,N_9880,N_9658);
nor UO_880 (O_880,N_9631,N_9570);
or UO_881 (O_881,N_9517,N_9055);
nand UO_882 (O_882,N_9376,N_9435);
nor UO_883 (O_883,N_9938,N_9482);
and UO_884 (O_884,N_9680,N_9995);
or UO_885 (O_885,N_9358,N_9807);
nand UO_886 (O_886,N_9651,N_9014);
or UO_887 (O_887,N_9228,N_9027);
or UO_888 (O_888,N_9690,N_9622);
or UO_889 (O_889,N_9585,N_9823);
nand UO_890 (O_890,N_9348,N_9782);
nand UO_891 (O_891,N_9908,N_9130);
xor UO_892 (O_892,N_9439,N_9092);
nand UO_893 (O_893,N_9124,N_9150);
or UO_894 (O_894,N_9344,N_9646);
or UO_895 (O_895,N_9285,N_9925);
or UO_896 (O_896,N_9055,N_9103);
nor UO_897 (O_897,N_9175,N_9062);
nor UO_898 (O_898,N_9306,N_9046);
nand UO_899 (O_899,N_9766,N_9421);
nand UO_900 (O_900,N_9569,N_9179);
nor UO_901 (O_901,N_9456,N_9001);
or UO_902 (O_902,N_9775,N_9141);
nand UO_903 (O_903,N_9278,N_9998);
and UO_904 (O_904,N_9673,N_9648);
nand UO_905 (O_905,N_9266,N_9748);
or UO_906 (O_906,N_9569,N_9272);
xnor UO_907 (O_907,N_9710,N_9946);
xor UO_908 (O_908,N_9178,N_9549);
xnor UO_909 (O_909,N_9361,N_9635);
nand UO_910 (O_910,N_9557,N_9301);
or UO_911 (O_911,N_9226,N_9870);
or UO_912 (O_912,N_9790,N_9899);
or UO_913 (O_913,N_9820,N_9773);
and UO_914 (O_914,N_9752,N_9888);
or UO_915 (O_915,N_9568,N_9381);
or UO_916 (O_916,N_9736,N_9344);
nor UO_917 (O_917,N_9237,N_9387);
and UO_918 (O_918,N_9269,N_9032);
and UO_919 (O_919,N_9119,N_9198);
and UO_920 (O_920,N_9704,N_9479);
xor UO_921 (O_921,N_9137,N_9739);
nand UO_922 (O_922,N_9989,N_9374);
or UO_923 (O_923,N_9581,N_9244);
and UO_924 (O_924,N_9872,N_9951);
or UO_925 (O_925,N_9983,N_9290);
or UO_926 (O_926,N_9999,N_9408);
or UO_927 (O_927,N_9757,N_9241);
xor UO_928 (O_928,N_9794,N_9060);
or UO_929 (O_929,N_9093,N_9774);
and UO_930 (O_930,N_9989,N_9138);
nand UO_931 (O_931,N_9207,N_9518);
or UO_932 (O_932,N_9003,N_9364);
nand UO_933 (O_933,N_9572,N_9296);
nor UO_934 (O_934,N_9171,N_9823);
nor UO_935 (O_935,N_9758,N_9524);
or UO_936 (O_936,N_9501,N_9195);
nand UO_937 (O_937,N_9265,N_9296);
nand UO_938 (O_938,N_9593,N_9790);
and UO_939 (O_939,N_9240,N_9822);
and UO_940 (O_940,N_9064,N_9219);
nand UO_941 (O_941,N_9185,N_9843);
xnor UO_942 (O_942,N_9168,N_9066);
and UO_943 (O_943,N_9422,N_9805);
nand UO_944 (O_944,N_9274,N_9153);
and UO_945 (O_945,N_9909,N_9300);
and UO_946 (O_946,N_9485,N_9100);
nand UO_947 (O_947,N_9240,N_9861);
and UO_948 (O_948,N_9492,N_9118);
nor UO_949 (O_949,N_9012,N_9401);
and UO_950 (O_950,N_9410,N_9645);
nor UO_951 (O_951,N_9761,N_9856);
xor UO_952 (O_952,N_9770,N_9091);
nor UO_953 (O_953,N_9232,N_9036);
and UO_954 (O_954,N_9696,N_9666);
nand UO_955 (O_955,N_9345,N_9126);
and UO_956 (O_956,N_9473,N_9434);
or UO_957 (O_957,N_9299,N_9184);
nand UO_958 (O_958,N_9075,N_9236);
and UO_959 (O_959,N_9542,N_9587);
nor UO_960 (O_960,N_9941,N_9747);
xor UO_961 (O_961,N_9653,N_9340);
or UO_962 (O_962,N_9000,N_9966);
or UO_963 (O_963,N_9193,N_9171);
or UO_964 (O_964,N_9321,N_9270);
nand UO_965 (O_965,N_9477,N_9040);
nand UO_966 (O_966,N_9568,N_9368);
xnor UO_967 (O_967,N_9156,N_9188);
xnor UO_968 (O_968,N_9613,N_9961);
nor UO_969 (O_969,N_9181,N_9310);
nor UO_970 (O_970,N_9471,N_9956);
xnor UO_971 (O_971,N_9649,N_9168);
nor UO_972 (O_972,N_9038,N_9499);
nor UO_973 (O_973,N_9634,N_9441);
and UO_974 (O_974,N_9211,N_9939);
nand UO_975 (O_975,N_9968,N_9972);
or UO_976 (O_976,N_9508,N_9244);
nand UO_977 (O_977,N_9691,N_9589);
and UO_978 (O_978,N_9595,N_9479);
nand UO_979 (O_979,N_9700,N_9680);
nor UO_980 (O_980,N_9145,N_9071);
nor UO_981 (O_981,N_9317,N_9367);
or UO_982 (O_982,N_9614,N_9491);
nor UO_983 (O_983,N_9140,N_9467);
nand UO_984 (O_984,N_9089,N_9666);
nand UO_985 (O_985,N_9235,N_9154);
or UO_986 (O_986,N_9364,N_9715);
nor UO_987 (O_987,N_9124,N_9156);
and UO_988 (O_988,N_9022,N_9958);
or UO_989 (O_989,N_9229,N_9309);
nor UO_990 (O_990,N_9992,N_9531);
nor UO_991 (O_991,N_9547,N_9058);
nand UO_992 (O_992,N_9072,N_9211);
and UO_993 (O_993,N_9221,N_9212);
nand UO_994 (O_994,N_9370,N_9985);
or UO_995 (O_995,N_9921,N_9451);
or UO_996 (O_996,N_9342,N_9891);
and UO_997 (O_997,N_9058,N_9652);
nand UO_998 (O_998,N_9151,N_9086);
nand UO_999 (O_999,N_9987,N_9002);
and UO_1000 (O_1000,N_9235,N_9726);
or UO_1001 (O_1001,N_9764,N_9868);
and UO_1002 (O_1002,N_9570,N_9229);
xnor UO_1003 (O_1003,N_9469,N_9291);
or UO_1004 (O_1004,N_9372,N_9366);
and UO_1005 (O_1005,N_9760,N_9539);
or UO_1006 (O_1006,N_9458,N_9675);
nand UO_1007 (O_1007,N_9179,N_9520);
or UO_1008 (O_1008,N_9821,N_9510);
or UO_1009 (O_1009,N_9299,N_9988);
xnor UO_1010 (O_1010,N_9738,N_9003);
or UO_1011 (O_1011,N_9506,N_9682);
and UO_1012 (O_1012,N_9937,N_9659);
and UO_1013 (O_1013,N_9637,N_9714);
nand UO_1014 (O_1014,N_9991,N_9315);
or UO_1015 (O_1015,N_9553,N_9548);
nand UO_1016 (O_1016,N_9784,N_9629);
nand UO_1017 (O_1017,N_9577,N_9491);
or UO_1018 (O_1018,N_9203,N_9304);
xor UO_1019 (O_1019,N_9680,N_9912);
nor UO_1020 (O_1020,N_9821,N_9663);
or UO_1021 (O_1021,N_9098,N_9512);
and UO_1022 (O_1022,N_9984,N_9460);
xnor UO_1023 (O_1023,N_9820,N_9819);
or UO_1024 (O_1024,N_9736,N_9493);
or UO_1025 (O_1025,N_9813,N_9473);
or UO_1026 (O_1026,N_9665,N_9656);
nand UO_1027 (O_1027,N_9635,N_9237);
and UO_1028 (O_1028,N_9807,N_9514);
nor UO_1029 (O_1029,N_9318,N_9759);
and UO_1030 (O_1030,N_9964,N_9290);
nand UO_1031 (O_1031,N_9222,N_9378);
nor UO_1032 (O_1032,N_9608,N_9319);
or UO_1033 (O_1033,N_9787,N_9446);
nand UO_1034 (O_1034,N_9574,N_9985);
xor UO_1035 (O_1035,N_9470,N_9643);
and UO_1036 (O_1036,N_9380,N_9147);
and UO_1037 (O_1037,N_9094,N_9101);
xor UO_1038 (O_1038,N_9201,N_9836);
nand UO_1039 (O_1039,N_9867,N_9575);
nand UO_1040 (O_1040,N_9562,N_9519);
nor UO_1041 (O_1041,N_9538,N_9184);
and UO_1042 (O_1042,N_9640,N_9539);
xnor UO_1043 (O_1043,N_9979,N_9785);
or UO_1044 (O_1044,N_9892,N_9375);
or UO_1045 (O_1045,N_9763,N_9831);
nor UO_1046 (O_1046,N_9764,N_9632);
nand UO_1047 (O_1047,N_9759,N_9970);
or UO_1048 (O_1048,N_9718,N_9983);
and UO_1049 (O_1049,N_9070,N_9217);
xor UO_1050 (O_1050,N_9514,N_9408);
and UO_1051 (O_1051,N_9579,N_9456);
xor UO_1052 (O_1052,N_9360,N_9160);
nor UO_1053 (O_1053,N_9103,N_9847);
nand UO_1054 (O_1054,N_9281,N_9763);
xor UO_1055 (O_1055,N_9313,N_9501);
nor UO_1056 (O_1056,N_9486,N_9538);
and UO_1057 (O_1057,N_9714,N_9166);
or UO_1058 (O_1058,N_9962,N_9824);
or UO_1059 (O_1059,N_9158,N_9287);
or UO_1060 (O_1060,N_9999,N_9110);
and UO_1061 (O_1061,N_9009,N_9249);
and UO_1062 (O_1062,N_9611,N_9062);
nor UO_1063 (O_1063,N_9455,N_9852);
or UO_1064 (O_1064,N_9432,N_9048);
nor UO_1065 (O_1065,N_9843,N_9152);
or UO_1066 (O_1066,N_9930,N_9498);
nor UO_1067 (O_1067,N_9944,N_9673);
and UO_1068 (O_1068,N_9754,N_9418);
nand UO_1069 (O_1069,N_9902,N_9627);
xor UO_1070 (O_1070,N_9103,N_9172);
nor UO_1071 (O_1071,N_9313,N_9433);
nand UO_1072 (O_1072,N_9351,N_9460);
nand UO_1073 (O_1073,N_9266,N_9320);
or UO_1074 (O_1074,N_9807,N_9133);
and UO_1075 (O_1075,N_9639,N_9902);
nand UO_1076 (O_1076,N_9900,N_9871);
nor UO_1077 (O_1077,N_9947,N_9299);
and UO_1078 (O_1078,N_9949,N_9787);
and UO_1079 (O_1079,N_9573,N_9730);
nand UO_1080 (O_1080,N_9423,N_9830);
or UO_1081 (O_1081,N_9765,N_9059);
or UO_1082 (O_1082,N_9901,N_9904);
nand UO_1083 (O_1083,N_9192,N_9023);
nand UO_1084 (O_1084,N_9007,N_9100);
xor UO_1085 (O_1085,N_9864,N_9241);
nor UO_1086 (O_1086,N_9064,N_9689);
nand UO_1087 (O_1087,N_9117,N_9579);
or UO_1088 (O_1088,N_9522,N_9258);
nand UO_1089 (O_1089,N_9450,N_9178);
and UO_1090 (O_1090,N_9828,N_9114);
and UO_1091 (O_1091,N_9026,N_9854);
xnor UO_1092 (O_1092,N_9357,N_9683);
nand UO_1093 (O_1093,N_9277,N_9754);
and UO_1094 (O_1094,N_9399,N_9481);
or UO_1095 (O_1095,N_9143,N_9270);
and UO_1096 (O_1096,N_9375,N_9115);
xnor UO_1097 (O_1097,N_9677,N_9587);
nand UO_1098 (O_1098,N_9944,N_9470);
nand UO_1099 (O_1099,N_9368,N_9526);
nor UO_1100 (O_1100,N_9851,N_9819);
or UO_1101 (O_1101,N_9345,N_9006);
nor UO_1102 (O_1102,N_9102,N_9956);
nor UO_1103 (O_1103,N_9562,N_9967);
nor UO_1104 (O_1104,N_9905,N_9475);
nand UO_1105 (O_1105,N_9670,N_9100);
xor UO_1106 (O_1106,N_9082,N_9804);
xor UO_1107 (O_1107,N_9537,N_9550);
and UO_1108 (O_1108,N_9106,N_9339);
or UO_1109 (O_1109,N_9301,N_9446);
nand UO_1110 (O_1110,N_9163,N_9369);
or UO_1111 (O_1111,N_9642,N_9734);
nor UO_1112 (O_1112,N_9829,N_9121);
and UO_1113 (O_1113,N_9884,N_9609);
and UO_1114 (O_1114,N_9157,N_9222);
and UO_1115 (O_1115,N_9041,N_9648);
nor UO_1116 (O_1116,N_9798,N_9171);
nor UO_1117 (O_1117,N_9248,N_9759);
and UO_1118 (O_1118,N_9539,N_9341);
and UO_1119 (O_1119,N_9813,N_9386);
nand UO_1120 (O_1120,N_9868,N_9103);
and UO_1121 (O_1121,N_9062,N_9386);
nor UO_1122 (O_1122,N_9901,N_9589);
nand UO_1123 (O_1123,N_9068,N_9256);
nor UO_1124 (O_1124,N_9795,N_9761);
or UO_1125 (O_1125,N_9618,N_9449);
nand UO_1126 (O_1126,N_9128,N_9417);
nor UO_1127 (O_1127,N_9547,N_9302);
and UO_1128 (O_1128,N_9449,N_9027);
and UO_1129 (O_1129,N_9528,N_9329);
nand UO_1130 (O_1130,N_9964,N_9248);
and UO_1131 (O_1131,N_9281,N_9831);
and UO_1132 (O_1132,N_9612,N_9827);
nor UO_1133 (O_1133,N_9625,N_9010);
or UO_1134 (O_1134,N_9721,N_9085);
nand UO_1135 (O_1135,N_9182,N_9390);
nand UO_1136 (O_1136,N_9147,N_9590);
nand UO_1137 (O_1137,N_9460,N_9057);
or UO_1138 (O_1138,N_9077,N_9453);
and UO_1139 (O_1139,N_9211,N_9823);
or UO_1140 (O_1140,N_9071,N_9357);
and UO_1141 (O_1141,N_9485,N_9786);
nor UO_1142 (O_1142,N_9808,N_9936);
xnor UO_1143 (O_1143,N_9221,N_9786);
or UO_1144 (O_1144,N_9025,N_9831);
xor UO_1145 (O_1145,N_9918,N_9593);
or UO_1146 (O_1146,N_9695,N_9195);
xor UO_1147 (O_1147,N_9034,N_9049);
or UO_1148 (O_1148,N_9248,N_9921);
nand UO_1149 (O_1149,N_9852,N_9146);
nand UO_1150 (O_1150,N_9766,N_9672);
or UO_1151 (O_1151,N_9746,N_9081);
nand UO_1152 (O_1152,N_9745,N_9171);
and UO_1153 (O_1153,N_9379,N_9364);
xnor UO_1154 (O_1154,N_9633,N_9970);
nor UO_1155 (O_1155,N_9385,N_9695);
or UO_1156 (O_1156,N_9060,N_9866);
nand UO_1157 (O_1157,N_9171,N_9094);
and UO_1158 (O_1158,N_9271,N_9830);
nor UO_1159 (O_1159,N_9771,N_9324);
or UO_1160 (O_1160,N_9668,N_9993);
nand UO_1161 (O_1161,N_9984,N_9710);
nand UO_1162 (O_1162,N_9523,N_9461);
or UO_1163 (O_1163,N_9079,N_9358);
or UO_1164 (O_1164,N_9525,N_9330);
and UO_1165 (O_1165,N_9008,N_9196);
and UO_1166 (O_1166,N_9925,N_9898);
xor UO_1167 (O_1167,N_9880,N_9539);
or UO_1168 (O_1168,N_9800,N_9729);
or UO_1169 (O_1169,N_9864,N_9529);
nand UO_1170 (O_1170,N_9689,N_9332);
and UO_1171 (O_1171,N_9346,N_9724);
nor UO_1172 (O_1172,N_9908,N_9897);
or UO_1173 (O_1173,N_9405,N_9197);
and UO_1174 (O_1174,N_9542,N_9326);
or UO_1175 (O_1175,N_9780,N_9291);
nand UO_1176 (O_1176,N_9363,N_9548);
nor UO_1177 (O_1177,N_9290,N_9528);
and UO_1178 (O_1178,N_9113,N_9909);
nor UO_1179 (O_1179,N_9217,N_9513);
nand UO_1180 (O_1180,N_9049,N_9603);
nor UO_1181 (O_1181,N_9433,N_9906);
and UO_1182 (O_1182,N_9183,N_9449);
and UO_1183 (O_1183,N_9707,N_9298);
nand UO_1184 (O_1184,N_9459,N_9050);
nor UO_1185 (O_1185,N_9916,N_9708);
nand UO_1186 (O_1186,N_9120,N_9027);
and UO_1187 (O_1187,N_9354,N_9174);
and UO_1188 (O_1188,N_9137,N_9374);
and UO_1189 (O_1189,N_9597,N_9661);
or UO_1190 (O_1190,N_9585,N_9272);
or UO_1191 (O_1191,N_9510,N_9892);
nor UO_1192 (O_1192,N_9132,N_9727);
or UO_1193 (O_1193,N_9798,N_9334);
nand UO_1194 (O_1194,N_9910,N_9015);
and UO_1195 (O_1195,N_9070,N_9525);
xor UO_1196 (O_1196,N_9674,N_9243);
and UO_1197 (O_1197,N_9131,N_9293);
nor UO_1198 (O_1198,N_9230,N_9200);
nor UO_1199 (O_1199,N_9429,N_9357);
or UO_1200 (O_1200,N_9792,N_9914);
xor UO_1201 (O_1201,N_9628,N_9998);
or UO_1202 (O_1202,N_9277,N_9953);
nor UO_1203 (O_1203,N_9248,N_9407);
nor UO_1204 (O_1204,N_9888,N_9883);
xor UO_1205 (O_1205,N_9262,N_9417);
nor UO_1206 (O_1206,N_9234,N_9997);
nand UO_1207 (O_1207,N_9313,N_9924);
or UO_1208 (O_1208,N_9796,N_9643);
and UO_1209 (O_1209,N_9856,N_9267);
or UO_1210 (O_1210,N_9710,N_9066);
and UO_1211 (O_1211,N_9264,N_9544);
nor UO_1212 (O_1212,N_9467,N_9928);
and UO_1213 (O_1213,N_9447,N_9182);
and UO_1214 (O_1214,N_9270,N_9754);
nor UO_1215 (O_1215,N_9583,N_9616);
nor UO_1216 (O_1216,N_9092,N_9335);
xor UO_1217 (O_1217,N_9316,N_9280);
nor UO_1218 (O_1218,N_9540,N_9291);
xnor UO_1219 (O_1219,N_9240,N_9929);
and UO_1220 (O_1220,N_9432,N_9137);
and UO_1221 (O_1221,N_9401,N_9853);
xnor UO_1222 (O_1222,N_9648,N_9105);
and UO_1223 (O_1223,N_9324,N_9097);
or UO_1224 (O_1224,N_9608,N_9396);
and UO_1225 (O_1225,N_9680,N_9892);
and UO_1226 (O_1226,N_9801,N_9433);
and UO_1227 (O_1227,N_9360,N_9632);
and UO_1228 (O_1228,N_9960,N_9425);
and UO_1229 (O_1229,N_9323,N_9249);
or UO_1230 (O_1230,N_9663,N_9999);
and UO_1231 (O_1231,N_9657,N_9399);
nor UO_1232 (O_1232,N_9417,N_9990);
nor UO_1233 (O_1233,N_9463,N_9122);
nor UO_1234 (O_1234,N_9236,N_9669);
nor UO_1235 (O_1235,N_9710,N_9515);
xor UO_1236 (O_1236,N_9665,N_9243);
or UO_1237 (O_1237,N_9565,N_9750);
nand UO_1238 (O_1238,N_9366,N_9553);
nor UO_1239 (O_1239,N_9992,N_9112);
nand UO_1240 (O_1240,N_9859,N_9719);
xor UO_1241 (O_1241,N_9868,N_9145);
nor UO_1242 (O_1242,N_9976,N_9491);
nor UO_1243 (O_1243,N_9242,N_9111);
and UO_1244 (O_1244,N_9120,N_9801);
or UO_1245 (O_1245,N_9959,N_9207);
and UO_1246 (O_1246,N_9358,N_9334);
xor UO_1247 (O_1247,N_9431,N_9201);
nand UO_1248 (O_1248,N_9694,N_9611);
nor UO_1249 (O_1249,N_9541,N_9606);
nand UO_1250 (O_1250,N_9611,N_9648);
xor UO_1251 (O_1251,N_9403,N_9492);
xor UO_1252 (O_1252,N_9651,N_9426);
nor UO_1253 (O_1253,N_9326,N_9437);
xnor UO_1254 (O_1254,N_9480,N_9105);
or UO_1255 (O_1255,N_9997,N_9857);
nand UO_1256 (O_1256,N_9165,N_9956);
or UO_1257 (O_1257,N_9737,N_9448);
and UO_1258 (O_1258,N_9420,N_9277);
or UO_1259 (O_1259,N_9048,N_9158);
nor UO_1260 (O_1260,N_9721,N_9152);
and UO_1261 (O_1261,N_9900,N_9242);
and UO_1262 (O_1262,N_9941,N_9996);
nor UO_1263 (O_1263,N_9373,N_9989);
nand UO_1264 (O_1264,N_9502,N_9240);
xnor UO_1265 (O_1265,N_9638,N_9372);
nor UO_1266 (O_1266,N_9386,N_9239);
nand UO_1267 (O_1267,N_9499,N_9715);
or UO_1268 (O_1268,N_9201,N_9434);
and UO_1269 (O_1269,N_9464,N_9579);
nor UO_1270 (O_1270,N_9887,N_9094);
nor UO_1271 (O_1271,N_9747,N_9344);
or UO_1272 (O_1272,N_9325,N_9994);
xor UO_1273 (O_1273,N_9132,N_9738);
or UO_1274 (O_1274,N_9422,N_9090);
nand UO_1275 (O_1275,N_9757,N_9824);
or UO_1276 (O_1276,N_9793,N_9850);
nand UO_1277 (O_1277,N_9564,N_9491);
and UO_1278 (O_1278,N_9116,N_9743);
nand UO_1279 (O_1279,N_9988,N_9246);
xnor UO_1280 (O_1280,N_9069,N_9979);
xor UO_1281 (O_1281,N_9603,N_9475);
xor UO_1282 (O_1282,N_9896,N_9782);
nor UO_1283 (O_1283,N_9687,N_9896);
and UO_1284 (O_1284,N_9788,N_9883);
xor UO_1285 (O_1285,N_9650,N_9255);
or UO_1286 (O_1286,N_9736,N_9885);
and UO_1287 (O_1287,N_9212,N_9739);
nand UO_1288 (O_1288,N_9288,N_9342);
and UO_1289 (O_1289,N_9855,N_9961);
or UO_1290 (O_1290,N_9568,N_9608);
nand UO_1291 (O_1291,N_9434,N_9704);
or UO_1292 (O_1292,N_9028,N_9918);
nor UO_1293 (O_1293,N_9284,N_9762);
and UO_1294 (O_1294,N_9595,N_9749);
nand UO_1295 (O_1295,N_9218,N_9001);
nor UO_1296 (O_1296,N_9310,N_9727);
nor UO_1297 (O_1297,N_9392,N_9466);
or UO_1298 (O_1298,N_9360,N_9408);
nand UO_1299 (O_1299,N_9987,N_9628);
or UO_1300 (O_1300,N_9478,N_9228);
nor UO_1301 (O_1301,N_9723,N_9656);
nand UO_1302 (O_1302,N_9146,N_9415);
or UO_1303 (O_1303,N_9177,N_9438);
nand UO_1304 (O_1304,N_9770,N_9210);
and UO_1305 (O_1305,N_9874,N_9029);
xor UO_1306 (O_1306,N_9859,N_9434);
or UO_1307 (O_1307,N_9003,N_9068);
and UO_1308 (O_1308,N_9400,N_9421);
and UO_1309 (O_1309,N_9310,N_9863);
xor UO_1310 (O_1310,N_9748,N_9206);
and UO_1311 (O_1311,N_9809,N_9332);
nor UO_1312 (O_1312,N_9902,N_9069);
nor UO_1313 (O_1313,N_9366,N_9632);
and UO_1314 (O_1314,N_9776,N_9662);
nor UO_1315 (O_1315,N_9267,N_9726);
or UO_1316 (O_1316,N_9391,N_9351);
nor UO_1317 (O_1317,N_9347,N_9612);
and UO_1318 (O_1318,N_9131,N_9634);
nand UO_1319 (O_1319,N_9208,N_9715);
and UO_1320 (O_1320,N_9172,N_9830);
or UO_1321 (O_1321,N_9899,N_9067);
or UO_1322 (O_1322,N_9122,N_9368);
xor UO_1323 (O_1323,N_9058,N_9169);
nor UO_1324 (O_1324,N_9639,N_9989);
xor UO_1325 (O_1325,N_9659,N_9277);
nand UO_1326 (O_1326,N_9831,N_9920);
nand UO_1327 (O_1327,N_9533,N_9246);
and UO_1328 (O_1328,N_9365,N_9314);
or UO_1329 (O_1329,N_9980,N_9776);
and UO_1330 (O_1330,N_9946,N_9585);
or UO_1331 (O_1331,N_9438,N_9031);
nor UO_1332 (O_1332,N_9338,N_9592);
nand UO_1333 (O_1333,N_9954,N_9340);
or UO_1334 (O_1334,N_9138,N_9066);
and UO_1335 (O_1335,N_9226,N_9378);
or UO_1336 (O_1336,N_9621,N_9909);
nor UO_1337 (O_1337,N_9348,N_9448);
nor UO_1338 (O_1338,N_9519,N_9608);
and UO_1339 (O_1339,N_9375,N_9555);
and UO_1340 (O_1340,N_9871,N_9551);
or UO_1341 (O_1341,N_9695,N_9721);
nor UO_1342 (O_1342,N_9164,N_9410);
nor UO_1343 (O_1343,N_9668,N_9708);
nor UO_1344 (O_1344,N_9176,N_9921);
and UO_1345 (O_1345,N_9460,N_9780);
or UO_1346 (O_1346,N_9634,N_9213);
and UO_1347 (O_1347,N_9478,N_9344);
and UO_1348 (O_1348,N_9801,N_9386);
and UO_1349 (O_1349,N_9924,N_9170);
nand UO_1350 (O_1350,N_9952,N_9487);
nor UO_1351 (O_1351,N_9595,N_9865);
or UO_1352 (O_1352,N_9122,N_9039);
nor UO_1353 (O_1353,N_9167,N_9202);
and UO_1354 (O_1354,N_9852,N_9372);
nand UO_1355 (O_1355,N_9394,N_9327);
nor UO_1356 (O_1356,N_9166,N_9532);
or UO_1357 (O_1357,N_9487,N_9289);
and UO_1358 (O_1358,N_9987,N_9159);
nand UO_1359 (O_1359,N_9545,N_9409);
or UO_1360 (O_1360,N_9450,N_9458);
nand UO_1361 (O_1361,N_9991,N_9898);
xnor UO_1362 (O_1362,N_9407,N_9906);
nand UO_1363 (O_1363,N_9596,N_9403);
and UO_1364 (O_1364,N_9834,N_9765);
or UO_1365 (O_1365,N_9686,N_9092);
nor UO_1366 (O_1366,N_9753,N_9210);
nand UO_1367 (O_1367,N_9773,N_9444);
xor UO_1368 (O_1368,N_9654,N_9635);
or UO_1369 (O_1369,N_9582,N_9475);
nand UO_1370 (O_1370,N_9697,N_9513);
or UO_1371 (O_1371,N_9230,N_9286);
nor UO_1372 (O_1372,N_9183,N_9696);
nand UO_1373 (O_1373,N_9873,N_9780);
nor UO_1374 (O_1374,N_9528,N_9647);
or UO_1375 (O_1375,N_9123,N_9902);
nor UO_1376 (O_1376,N_9886,N_9851);
nand UO_1377 (O_1377,N_9520,N_9060);
nand UO_1378 (O_1378,N_9194,N_9803);
nor UO_1379 (O_1379,N_9704,N_9368);
xor UO_1380 (O_1380,N_9932,N_9535);
or UO_1381 (O_1381,N_9642,N_9082);
nor UO_1382 (O_1382,N_9031,N_9350);
and UO_1383 (O_1383,N_9926,N_9524);
and UO_1384 (O_1384,N_9096,N_9389);
and UO_1385 (O_1385,N_9962,N_9603);
and UO_1386 (O_1386,N_9488,N_9091);
nor UO_1387 (O_1387,N_9802,N_9989);
nor UO_1388 (O_1388,N_9909,N_9938);
and UO_1389 (O_1389,N_9121,N_9079);
nor UO_1390 (O_1390,N_9120,N_9274);
nand UO_1391 (O_1391,N_9849,N_9502);
nand UO_1392 (O_1392,N_9767,N_9394);
xor UO_1393 (O_1393,N_9817,N_9217);
or UO_1394 (O_1394,N_9240,N_9465);
xor UO_1395 (O_1395,N_9836,N_9623);
xnor UO_1396 (O_1396,N_9893,N_9449);
and UO_1397 (O_1397,N_9250,N_9932);
and UO_1398 (O_1398,N_9032,N_9196);
or UO_1399 (O_1399,N_9405,N_9528);
or UO_1400 (O_1400,N_9067,N_9257);
nor UO_1401 (O_1401,N_9937,N_9997);
and UO_1402 (O_1402,N_9369,N_9151);
or UO_1403 (O_1403,N_9546,N_9711);
or UO_1404 (O_1404,N_9625,N_9753);
nor UO_1405 (O_1405,N_9346,N_9565);
nor UO_1406 (O_1406,N_9568,N_9013);
and UO_1407 (O_1407,N_9604,N_9678);
and UO_1408 (O_1408,N_9179,N_9882);
nand UO_1409 (O_1409,N_9126,N_9270);
or UO_1410 (O_1410,N_9868,N_9384);
or UO_1411 (O_1411,N_9964,N_9766);
or UO_1412 (O_1412,N_9108,N_9022);
and UO_1413 (O_1413,N_9708,N_9372);
or UO_1414 (O_1414,N_9221,N_9737);
or UO_1415 (O_1415,N_9528,N_9474);
or UO_1416 (O_1416,N_9662,N_9774);
and UO_1417 (O_1417,N_9170,N_9852);
or UO_1418 (O_1418,N_9566,N_9121);
xor UO_1419 (O_1419,N_9077,N_9728);
xor UO_1420 (O_1420,N_9258,N_9701);
nor UO_1421 (O_1421,N_9353,N_9979);
and UO_1422 (O_1422,N_9994,N_9400);
nand UO_1423 (O_1423,N_9319,N_9717);
and UO_1424 (O_1424,N_9826,N_9527);
or UO_1425 (O_1425,N_9030,N_9065);
nor UO_1426 (O_1426,N_9345,N_9410);
xor UO_1427 (O_1427,N_9798,N_9831);
or UO_1428 (O_1428,N_9747,N_9253);
nand UO_1429 (O_1429,N_9597,N_9522);
or UO_1430 (O_1430,N_9590,N_9976);
or UO_1431 (O_1431,N_9785,N_9795);
or UO_1432 (O_1432,N_9954,N_9850);
and UO_1433 (O_1433,N_9783,N_9898);
or UO_1434 (O_1434,N_9750,N_9263);
or UO_1435 (O_1435,N_9261,N_9944);
and UO_1436 (O_1436,N_9437,N_9611);
and UO_1437 (O_1437,N_9356,N_9157);
nand UO_1438 (O_1438,N_9354,N_9130);
or UO_1439 (O_1439,N_9021,N_9606);
xor UO_1440 (O_1440,N_9632,N_9181);
nand UO_1441 (O_1441,N_9261,N_9949);
nand UO_1442 (O_1442,N_9728,N_9473);
nand UO_1443 (O_1443,N_9672,N_9574);
or UO_1444 (O_1444,N_9043,N_9597);
and UO_1445 (O_1445,N_9144,N_9715);
or UO_1446 (O_1446,N_9881,N_9279);
nand UO_1447 (O_1447,N_9712,N_9357);
nand UO_1448 (O_1448,N_9167,N_9950);
nand UO_1449 (O_1449,N_9457,N_9504);
and UO_1450 (O_1450,N_9854,N_9398);
and UO_1451 (O_1451,N_9641,N_9308);
and UO_1452 (O_1452,N_9924,N_9473);
nor UO_1453 (O_1453,N_9400,N_9579);
xnor UO_1454 (O_1454,N_9349,N_9693);
or UO_1455 (O_1455,N_9101,N_9243);
nor UO_1456 (O_1456,N_9523,N_9462);
nand UO_1457 (O_1457,N_9975,N_9881);
and UO_1458 (O_1458,N_9690,N_9248);
and UO_1459 (O_1459,N_9150,N_9481);
and UO_1460 (O_1460,N_9526,N_9071);
or UO_1461 (O_1461,N_9999,N_9685);
nor UO_1462 (O_1462,N_9266,N_9345);
nand UO_1463 (O_1463,N_9442,N_9981);
or UO_1464 (O_1464,N_9556,N_9139);
nor UO_1465 (O_1465,N_9744,N_9482);
or UO_1466 (O_1466,N_9473,N_9056);
and UO_1467 (O_1467,N_9013,N_9809);
or UO_1468 (O_1468,N_9725,N_9793);
and UO_1469 (O_1469,N_9561,N_9687);
nand UO_1470 (O_1470,N_9542,N_9053);
xor UO_1471 (O_1471,N_9839,N_9594);
nor UO_1472 (O_1472,N_9538,N_9493);
or UO_1473 (O_1473,N_9057,N_9023);
or UO_1474 (O_1474,N_9723,N_9316);
nor UO_1475 (O_1475,N_9511,N_9382);
and UO_1476 (O_1476,N_9294,N_9854);
xnor UO_1477 (O_1477,N_9517,N_9400);
or UO_1478 (O_1478,N_9753,N_9183);
or UO_1479 (O_1479,N_9801,N_9024);
xnor UO_1480 (O_1480,N_9969,N_9209);
nor UO_1481 (O_1481,N_9498,N_9979);
nand UO_1482 (O_1482,N_9974,N_9328);
nor UO_1483 (O_1483,N_9934,N_9127);
or UO_1484 (O_1484,N_9869,N_9893);
or UO_1485 (O_1485,N_9343,N_9521);
nand UO_1486 (O_1486,N_9573,N_9381);
and UO_1487 (O_1487,N_9189,N_9608);
and UO_1488 (O_1488,N_9796,N_9038);
xnor UO_1489 (O_1489,N_9256,N_9257);
nor UO_1490 (O_1490,N_9401,N_9087);
or UO_1491 (O_1491,N_9592,N_9235);
nor UO_1492 (O_1492,N_9439,N_9719);
and UO_1493 (O_1493,N_9989,N_9402);
and UO_1494 (O_1494,N_9457,N_9544);
nor UO_1495 (O_1495,N_9630,N_9737);
nor UO_1496 (O_1496,N_9765,N_9870);
or UO_1497 (O_1497,N_9686,N_9346);
xor UO_1498 (O_1498,N_9577,N_9188);
or UO_1499 (O_1499,N_9352,N_9296);
endmodule