module basic_3000_30000_3500_50_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
and U0 (N_0,In_2810,In_1537);
nand U1 (N_1,In_879,In_0);
or U2 (N_2,In_1420,In_105);
and U3 (N_3,In_2340,In_1193);
or U4 (N_4,In_2416,In_442);
nor U5 (N_5,In_1817,In_962);
xnor U6 (N_6,In_410,In_334);
xnor U7 (N_7,In_2087,In_2440);
nand U8 (N_8,In_2335,In_544);
or U9 (N_9,In_138,In_2849);
and U10 (N_10,In_2140,In_158);
nand U11 (N_11,In_1578,In_2013);
nand U12 (N_12,In_2762,In_2631);
and U13 (N_13,In_1490,In_1112);
nor U14 (N_14,In_2693,In_1172);
nand U15 (N_15,In_235,In_2374);
xnor U16 (N_16,In_2461,In_1706);
nor U17 (N_17,In_1318,In_1688);
nor U18 (N_18,In_1027,In_1801);
and U19 (N_19,In_220,In_2081);
or U20 (N_20,In_1534,In_806);
nand U21 (N_21,In_655,In_286);
or U22 (N_22,In_1292,In_255);
or U23 (N_23,In_1152,In_1224);
or U24 (N_24,In_1447,In_2732);
or U25 (N_25,In_1245,In_350);
nor U26 (N_26,In_2407,In_581);
xnor U27 (N_27,In_271,In_2551);
nor U28 (N_28,In_307,In_2537);
xnor U29 (N_29,In_876,In_1048);
or U30 (N_30,In_2609,In_990);
nor U31 (N_31,In_2687,In_2896);
nor U32 (N_32,In_1491,In_1994);
nor U33 (N_33,In_819,In_1339);
or U34 (N_34,In_308,In_1654);
nand U35 (N_35,In_2510,In_2878);
or U36 (N_36,In_277,In_306);
nor U37 (N_37,In_2520,In_101);
or U38 (N_38,In_2691,In_2563);
or U39 (N_39,In_1361,In_1100);
nand U40 (N_40,In_1041,In_1820);
or U41 (N_41,In_2095,In_2198);
or U42 (N_42,In_2851,In_2581);
and U43 (N_43,In_1657,In_1297);
nor U44 (N_44,In_2493,In_2304);
xnor U45 (N_45,In_2937,In_1922);
nor U46 (N_46,In_2589,In_752);
nand U47 (N_47,In_1990,In_69);
nand U48 (N_48,In_2587,In_1570);
nand U49 (N_49,In_413,In_1767);
nor U50 (N_50,In_2828,In_1958);
and U51 (N_51,In_1781,In_2492);
xor U52 (N_52,In_2248,In_2153);
nor U53 (N_53,In_1487,In_328);
nand U54 (N_54,In_2477,In_1583);
or U55 (N_55,In_2506,In_1686);
nor U56 (N_56,In_18,In_1009);
nand U57 (N_57,In_731,In_2848);
nand U58 (N_58,In_567,In_718);
nand U59 (N_59,In_199,In_911);
nand U60 (N_60,In_1705,In_1492);
xor U61 (N_61,In_1113,In_2194);
xnor U62 (N_62,In_1819,In_2858);
or U63 (N_63,In_2627,In_945);
nand U64 (N_64,In_1612,In_603);
nand U65 (N_65,In_119,In_681);
nand U66 (N_66,In_2402,In_904);
or U67 (N_67,In_2452,In_965);
xor U68 (N_68,In_1093,In_1911);
or U69 (N_69,In_154,In_1625);
nand U70 (N_70,In_1671,In_530);
xnor U71 (N_71,In_658,In_829);
or U72 (N_72,In_778,In_800);
nor U73 (N_73,In_999,In_2611);
nand U74 (N_74,In_2604,In_2953);
xor U75 (N_75,In_2593,In_2912);
nand U76 (N_76,In_985,In_1236);
or U77 (N_77,In_802,In_510);
or U78 (N_78,In_550,In_2145);
xnor U79 (N_79,In_327,In_211);
and U80 (N_80,In_2429,In_2926);
or U81 (N_81,In_318,In_2496);
or U82 (N_82,In_99,In_1164);
and U83 (N_83,In_2790,In_1878);
xor U84 (N_84,In_2472,In_1195);
nand U85 (N_85,In_2641,In_2777);
xor U86 (N_86,In_363,In_1645);
and U87 (N_87,In_2205,In_556);
nand U88 (N_88,In_2773,In_1453);
xor U89 (N_89,In_709,In_2916);
nor U90 (N_90,In_48,In_989);
xnor U91 (N_91,In_2874,In_2605);
nand U92 (N_92,In_414,In_2332);
nor U93 (N_93,In_299,In_1040);
or U94 (N_94,In_2987,In_2224);
nor U95 (N_95,In_2617,In_699);
nor U96 (N_96,In_1983,In_729);
nor U97 (N_97,In_2705,In_1146);
and U98 (N_98,In_950,In_424);
or U99 (N_99,In_881,In_1187);
nor U100 (N_100,In_604,In_148);
nor U101 (N_101,In_2623,In_1914);
nor U102 (N_102,In_1374,In_2888);
xnor U103 (N_103,In_1350,In_1023);
xor U104 (N_104,In_1376,In_2458);
xnor U105 (N_105,In_2033,In_517);
nor U106 (N_106,In_1504,In_1475);
nor U107 (N_107,In_944,In_1921);
or U108 (N_108,In_102,In_228);
nor U109 (N_109,In_1988,In_9);
nand U110 (N_110,In_1127,In_2917);
and U111 (N_111,In_1346,In_2695);
xor U112 (N_112,In_1594,In_229);
nor U113 (N_113,In_863,In_1078);
or U114 (N_114,In_1904,In_724);
and U115 (N_115,In_1201,In_1280);
nand U116 (N_116,In_2495,In_2067);
and U117 (N_117,In_2821,In_449);
and U118 (N_118,In_847,In_2804);
or U119 (N_119,In_2323,In_2977);
nand U120 (N_120,In_2583,In_1565);
xnor U121 (N_121,In_978,In_1549);
xnor U122 (N_122,In_2522,In_1162);
xor U123 (N_123,In_2988,In_1936);
nor U124 (N_124,In_78,In_464);
and U125 (N_125,In_2731,In_1235);
xnor U126 (N_126,In_2980,In_723);
or U127 (N_127,In_1906,In_656);
nand U128 (N_128,In_725,In_1118);
xor U129 (N_129,In_2512,In_1160);
and U130 (N_130,In_2908,In_592);
or U131 (N_131,In_2843,In_2803);
xnor U132 (N_132,In_2590,In_1282);
and U133 (N_133,In_2668,In_213);
nor U134 (N_134,In_364,In_1227);
or U135 (N_135,In_2613,In_354);
nor U136 (N_136,In_1584,In_2638);
nor U137 (N_137,In_2594,In_2230);
and U138 (N_138,In_2771,In_2329);
or U139 (N_139,In_2626,In_1883);
nand U140 (N_140,In_1055,In_2383);
and U141 (N_141,In_909,In_1577);
and U142 (N_142,In_1046,In_2904);
xor U143 (N_143,In_391,In_524);
xnor U144 (N_144,In_2303,In_1111);
xor U145 (N_145,In_2475,In_1156);
or U146 (N_146,In_2503,In_2368);
and U147 (N_147,In_2381,In_2357);
and U148 (N_148,In_1711,In_874);
nand U149 (N_149,In_1013,In_941);
or U150 (N_150,In_720,In_637);
xor U151 (N_151,In_2713,In_2183);
and U152 (N_152,In_2229,In_1818);
xnor U153 (N_153,In_2714,In_118);
or U154 (N_154,In_2666,In_260);
nor U155 (N_155,In_1553,In_852);
or U156 (N_156,In_804,In_2826);
or U157 (N_157,In_2756,In_2339);
or U158 (N_158,In_1895,In_773);
or U159 (N_159,In_2065,In_1868);
or U160 (N_160,In_2349,In_129);
or U161 (N_161,In_1793,In_823);
or U162 (N_162,In_1949,In_2723);
nor U163 (N_163,In_1629,In_2123);
xnor U164 (N_164,In_2263,In_2288);
xnor U165 (N_165,In_2514,In_1879);
nor U166 (N_166,In_1776,In_461);
xnor U167 (N_167,In_2394,In_1989);
xnor U168 (N_168,In_1255,In_64);
nor U169 (N_169,In_1807,In_1377);
and U170 (N_170,In_951,In_1016);
xnor U171 (N_171,In_1267,In_1951);
nand U172 (N_172,In_1708,In_1909);
and U173 (N_173,In_1473,In_1098);
xor U174 (N_174,In_34,In_2507);
nand U175 (N_175,In_1017,In_2539);
nand U176 (N_176,In_1669,In_1344);
nor U177 (N_177,In_2943,In_2062);
nor U178 (N_178,In_2859,In_813);
and U179 (N_179,In_13,In_234);
and U180 (N_180,In_858,In_2659);
and U181 (N_181,In_607,In_2361);
nand U182 (N_182,In_1269,In_2989);
or U183 (N_183,In_1387,In_1137);
and U184 (N_184,In_855,In_356);
and U185 (N_185,In_2029,In_304);
xor U186 (N_186,In_281,In_993);
nor U187 (N_187,In_2865,In_1823);
xor U188 (N_188,In_1701,In_505);
nor U189 (N_189,In_253,In_559);
nor U190 (N_190,In_736,In_2560);
nor U191 (N_191,In_849,In_1770);
or U192 (N_192,In_2390,In_1802);
xnor U193 (N_193,In_240,In_1950);
nand U194 (N_194,In_1219,In_2573);
and U195 (N_195,In_342,In_135);
nor U196 (N_196,In_2354,In_2270);
or U197 (N_197,In_2203,In_1147);
or U198 (N_198,In_1059,In_61);
nor U199 (N_199,In_1486,In_221);
nand U200 (N_200,In_846,In_1329);
xnor U201 (N_201,In_593,In_21);
and U202 (N_202,In_2376,In_1470);
and U203 (N_203,In_1020,In_1799);
and U204 (N_204,In_507,In_2176);
and U205 (N_205,In_1782,In_1448);
nor U206 (N_206,In_2995,In_623);
nor U207 (N_207,In_2491,In_1398);
and U208 (N_208,In_1321,In_1579);
and U209 (N_209,In_1190,In_2256);
nand U210 (N_210,In_42,In_1550);
xor U211 (N_211,In_2582,In_77);
xor U212 (N_212,In_2688,In_368);
xor U213 (N_213,In_2549,In_2350);
xor U214 (N_214,In_2328,In_1954);
nor U215 (N_215,In_711,In_1692);
nor U216 (N_216,In_411,In_2562);
xor U217 (N_217,In_1418,In_2929);
nand U218 (N_218,In_2375,In_2124);
and U219 (N_219,In_2296,In_2082);
and U220 (N_220,In_896,In_309);
nor U221 (N_221,In_1682,In_1797);
nand U222 (N_222,In_2423,In_2012);
nor U223 (N_223,In_1992,In_2138);
xnor U224 (N_224,In_1900,In_777);
nand U225 (N_225,In_236,In_2070);
xnor U226 (N_226,In_1691,In_1752);
xor U227 (N_227,In_2093,In_1441);
nor U228 (N_228,In_183,In_1898);
and U229 (N_229,In_261,In_1084);
xor U230 (N_230,In_1920,In_1636);
or U231 (N_231,In_1028,In_2258);
or U232 (N_232,In_2373,In_2252);
or U233 (N_233,In_1228,In_2089);
and U234 (N_234,In_1142,In_2923);
nor U235 (N_235,In_913,In_1264);
nor U236 (N_236,In_2818,In_1430);
or U237 (N_237,In_822,In_1938);
nor U238 (N_238,In_1365,In_279);
xnor U239 (N_239,In_1925,In_1757);
xnor U240 (N_240,In_476,In_2041);
or U241 (N_241,In_1996,In_1520);
and U242 (N_242,In_1004,In_2168);
xnor U243 (N_243,In_1070,In_305);
nand U244 (N_244,In_1945,In_1613);
xnor U245 (N_245,In_1639,In_1247);
nand U246 (N_246,In_1286,In_979);
nor U247 (N_247,In_2824,In_1272);
or U248 (N_248,In_1178,In_673);
nor U249 (N_249,In_2209,In_2961);
nand U250 (N_250,In_624,In_1039);
xor U251 (N_251,In_93,In_1206);
and U252 (N_252,In_2090,In_1773);
or U253 (N_253,In_212,In_685);
and U254 (N_254,In_1204,In_2106);
and U255 (N_255,In_2043,In_2184);
and U256 (N_256,In_1576,In_2715);
nand U257 (N_257,In_2892,In_738);
nand U258 (N_258,In_2311,In_2782);
nor U259 (N_259,In_2853,In_1434);
xnor U260 (N_260,In_226,In_2501);
nand U261 (N_261,In_2517,In_2728);
and U262 (N_262,In_126,In_1378);
and U263 (N_263,In_2947,In_964);
nor U264 (N_264,In_1423,In_2336);
or U265 (N_265,In_2660,In_1148);
xnor U266 (N_266,In_1080,In_1600);
and U267 (N_267,In_457,In_55);
xnor U268 (N_268,In_1853,In_1536);
or U269 (N_269,In_868,In_2628);
and U270 (N_270,In_696,In_1258);
nand U271 (N_271,In_1285,In_2286);
nor U272 (N_272,In_2457,In_2232);
nand U273 (N_273,In_1044,In_2971);
and U274 (N_274,In_2162,In_159);
or U275 (N_275,In_2314,In_2518);
or U276 (N_276,In_2164,In_2318);
nand U277 (N_277,In_582,In_1959);
nand U278 (N_278,In_1675,In_668);
xor U279 (N_279,In_1122,In_899);
or U280 (N_280,In_2442,In_2753);
nand U281 (N_281,In_735,In_1533);
nor U282 (N_282,In_2603,In_982);
xnor U283 (N_283,In_303,In_416);
or U284 (N_284,In_661,In_689);
or U285 (N_285,In_1062,In_1665);
xnor U286 (N_286,In_1305,In_2956);
nand U287 (N_287,In_1850,In_977);
xnor U288 (N_288,In_1031,In_1591);
or U289 (N_289,In_1754,In_2262);
nor U290 (N_290,In_1566,In_625);
nand U291 (N_291,In_1465,In_1144);
and U292 (N_292,In_2778,In_590);
and U293 (N_293,In_43,In_2978);
xnor U294 (N_294,In_2212,In_1170);
and U295 (N_295,In_1860,In_586);
nand U296 (N_296,In_938,In_917);
xnor U297 (N_297,In_1208,In_998);
nand U298 (N_298,In_186,In_2271);
xor U299 (N_299,In_572,In_293);
nand U300 (N_300,In_355,In_705);
nand U301 (N_301,In_2983,In_552);
and U302 (N_302,In_1859,In_1722);
or U303 (N_303,In_276,In_906);
xnor U304 (N_304,In_929,In_2453);
and U305 (N_305,In_830,In_2684);
xor U306 (N_306,In_2355,In_2307);
and U307 (N_307,In_1231,In_1116);
nand U308 (N_308,In_1923,In_875);
xor U309 (N_309,In_934,In_2298);
and U310 (N_310,In_1335,In_2763);
nand U311 (N_311,In_2201,In_2774);
nand U312 (N_312,In_1741,In_301);
nand U313 (N_313,In_1791,In_149);
xnor U314 (N_314,In_2612,In_2088);
nor U315 (N_315,In_2692,In_1667);
xnor U316 (N_316,In_203,In_2064);
and U317 (N_317,In_2542,In_1015);
and U318 (N_318,In_1238,In_2255);
and U319 (N_319,In_2797,In_1733);
or U320 (N_320,In_794,In_2422);
nor U321 (N_321,In_797,In_2727);
xor U322 (N_322,In_2806,In_139);
nand U323 (N_323,In_323,In_971);
or U324 (N_324,In_1391,In_2873);
nor U325 (N_325,In_1239,In_2338);
nand U326 (N_326,In_1413,In_1857);
or U327 (N_327,In_722,In_1425);
xor U328 (N_328,In_1596,In_85);
and U329 (N_329,In_2913,In_754);
nor U330 (N_330,In_1840,In_2552);
xnor U331 (N_331,In_1766,In_2607);
xnor U332 (N_332,In_2524,In_691);
and U333 (N_333,In_1944,In_2955);
xnor U334 (N_334,In_1088,In_2285);
nor U335 (N_335,In_2530,In_2750);
and U336 (N_336,In_6,In_1697);
nor U337 (N_337,In_1428,In_2595);
and U338 (N_338,In_2827,In_1186);
and U339 (N_339,In_2866,In_1276);
nor U340 (N_340,In_2941,In_1869);
nor U341 (N_341,In_2984,In_2042);
and U342 (N_342,In_2333,In_1975);
nand U343 (N_343,In_2238,In_1888);
or U344 (N_344,In_2584,In_836);
xor U345 (N_345,In_2559,In_390);
nor U346 (N_346,In_1341,In_1702);
and U347 (N_347,In_1035,In_2173);
nand U348 (N_348,In_833,In_895);
nor U349 (N_349,In_1198,In_378);
xnor U350 (N_350,In_2276,In_1829);
and U351 (N_351,In_181,In_20);
and U352 (N_352,In_1135,In_2720);
xnor U353 (N_353,In_1568,In_1472);
and U354 (N_354,In_447,In_97);
xnor U355 (N_355,In_2272,In_1010);
nor U356 (N_356,In_988,In_883);
or U357 (N_357,In_1556,In_2689);
xor U358 (N_358,In_436,In_1582);
and U359 (N_359,In_994,In_520);
xor U360 (N_360,In_2768,In_175);
xnor U361 (N_361,In_2190,In_2384);
nor U362 (N_362,In_1354,In_1191);
xnor U363 (N_363,In_1502,In_1256);
and U364 (N_364,In_1542,In_2253);
nor U365 (N_365,In_2898,In_145);
or U366 (N_366,In_1415,In_1953);
nand U367 (N_367,In_134,In_456);
xor U368 (N_368,In_1694,In_782);
or U369 (N_369,In_1471,In_2282);
or U370 (N_370,In_2654,In_956);
or U371 (N_371,In_278,In_1734);
and U372 (N_372,In_815,In_2066);
and U373 (N_373,In_1735,In_2385);
nand U374 (N_374,In_1887,In_1557);
and U375 (N_375,In_687,In_621);
and U376 (N_376,In_2137,In_1246);
and U377 (N_377,In_1086,In_2856);
and U378 (N_378,In_2791,In_1446);
xor U379 (N_379,In_2981,In_2949);
xor U380 (N_380,In_2893,In_1476);
nor U381 (N_381,In_345,In_1466);
nand U382 (N_382,In_2950,In_237);
xor U383 (N_383,In_1503,In_2134);
xor U384 (N_384,In_2108,In_2885);
xnor U385 (N_385,In_173,In_2277);
and U386 (N_386,In_367,In_179);
nor U387 (N_387,In_2553,In_515);
nor U388 (N_388,In_2125,In_1403);
xnor U389 (N_389,In_2967,In_2497);
nor U390 (N_390,In_666,In_2001);
nor U391 (N_391,In_1772,In_2504);
nor U392 (N_392,In_2743,In_1952);
xor U393 (N_393,In_2789,In_1574);
xor U394 (N_394,In_143,In_787);
and U395 (N_395,In_1459,In_799);
or U396 (N_396,In_2269,In_443);
or U397 (N_397,In_1333,In_2571);
and U398 (N_398,In_1729,In_1787);
and U399 (N_399,In_1194,In_1966);
xor U400 (N_400,In_2397,In_1998);
nand U401 (N_401,In_2048,In_2588);
nor U402 (N_402,In_2171,In_2657);
or U403 (N_403,In_289,In_486);
xnor U404 (N_404,In_1569,In_1454);
xnor U405 (N_405,In_2112,In_1631);
or U406 (N_406,In_1362,In_58);
nand U407 (N_407,In_1464,In_1514);
xor U408 (N_408,In_1867,In_71);
nand U409 (N_409,In_2356,In_2283);
or U410 (N_410,In_268,In_1544);
and U411 (N_411,In_1519,In_568);
and U412 (N_412,In_826,In_2734);
xnor U413 (N_413,In_1189,In_967);
xnor U414 (N_414,In_91,In_144);
or U415 (N_415,In_262,In_472);
xnor U416 (N_416,In_1092,In_2928);
or U417 (N_417,In_843,In_2895);
nor U418 (N_418,In_1581,In_2408);
and U419 (N_419,In_949,In_2104);
nor U420 (N_420,In_525,In_2403);
nor U421 (N_421,In_2215,In_1795);
nor U422 (N_422,In_419,In_1713);
or U423 (N_423,In_1375,In_939);
xor U424 (N_424,In_1221,In_728);
xnor U425 (N_425,In_2200,In_2651);
xor U426 (N_426,In_2841,In_543);
and U427 (N_427,In_371,In_639);
or U428 (N_428,In_249,In_250);
xnor U429 (N_429,In_2822,In_1014);
or U430 (N_430,In_2076,In_814);
or U431 (N_431,In_2960,In_2051);
or U432 (N_432,In_2807,In_2189);
and U433 (N_433,In_952,In_1687);
and U434 (N_434,In_1666,In_1664);
nor U435 (N_435,In_1678,In_1072);
and U436 (N_436,In_775,In_1724);
and U437 (N_437,In_1229,In_132);
and U438 (N_438,In_2724,In_454);
nor U439 (N_439,In_1412,In_810);
xor U440 (N_440,In_202,In_2244);
nand U441 (N_441,In_1442,In_152);
xor U442 (N_442,In_733,In_1618);
or U443 (N_443,In_12,In_49);
nand U444 (N_444,In_2109,In_2342);
nor U445 (N_445,In_2297,In_1607);
or U446 (N_446,In_2035,In_2935);
and U447 (N_447,In_1640,In_1635);
nor U448 (N_448,In_509,In_415);
nand U449 (N_449,In_2259,In_2174);
and U450 (N_450,In_1288,In_393);
and U451 (N_451,In_2877,In_1240);
or U452 (N_452,In_2922,In_23);
nand U453 (N_453,In_2557,In_2748);
nor U454 (N_454,In_201,In_1461);
and U455 (N_455,In_1901,In_2301);
nor U456 (N_456,In_1262,In_759);
or U457 (N_457,In_1609,In_538);
or U458 (N_458,In_2347,In_862);
nor U459 (N_459,In_233,In_381);
and U460 (N_460,In_2302,In_2103);
xnor U461 (N_461,In_1814,In_2868);
nand U462 (N_462,In_986,In_2681);
xor U463 (N_463,In_409,In_380);
nand U464 (N_464,In_160,In_351);
xnor U465 (N_465,In_30,In_2265);
or U466 (N_466,In_483,In_761);
and U467 (N_467,In_2694,In_1891);
nand U468 (N_468,In_995,In_2721);
xnor U469 (N_469,In_536,In_1337);
nor U470 (N_470,In_921,In_1019);
and U471 (N_471,In_1310,In_1138);
xnor U472 (N_472,In_499,In_848);
xnor U473 (N_473,In_1851,In_1680);
xor U474 (N_474,In_1668,In_2811);
xnor U475 (N_475,In_167,In_514);
nand U476 (N_476,In_2837,In_296);
nand U477 (N_477,In_1150,In_853);
xor U478 (N_478,In_743,In_5);
nor U479 (N_479,In_1424,In_2862);
xnor U480 (N_480,In_2236,In_1493);
nor U481 (N_481,In_357,In_803);
nor U482 (N_482,In_2523,In_943);
nand U483 (N_483,In_1546,In_2488);
nand U484 (N_484,In_710,In_1083);
or U485 (N_485,In_2141,In_460);
xnor U486 (N_486,In_774,In_916);
nor U487 (N_487,In_996,In_631);
and U488 (N_488,In_1474,In_627);
nor U489 (N_489,In_453,In_713);
or U490 (N_490,In_605,In_1439);
and U491 (N_491,In_1875,In_1907);
nor U492 (N_492,In_2680,In_2747);
and U493 (N_493,In_2556,In_1223);
xor U494 (N_494,In_2188,In_2759);
nand U495 (N_495,In_1979,In_2310);
or U496 (N_496,In_2234,In_2463);
or U497 (N_497,In_878,In_831);
and U498 (N_498,In_361,In_2447);
xor U499 (N_499,In_1030,In_1450);
and U500 (N_500,In_588,In_1233);
nand U501 (N_501,In_2021,In_511);
or U502 (N_502,In_2509,In_2656);
and U503 (N_503,In_2637,In_1167);
and U504 (N_504,In_2409,In_2293);
xnor U505 (N_505,In_545,In_825);
nand U506 (N_506,In_11,In_1317);
or U507 (N_507,In_1125,In_341);
nand U508 (N_508,In_2625,In_845);
xnor U509 (N_509,In_1764,In_95);
nor U510 (N_510,In_2850,In_1562);
nor U511 (N_511,In_861,In_2400);
nand U512 (N_512,In_1731,In_2091);
xnor U513 (N_513,In_267,In_548);
nor U514 (N_514,In_2471,In_1710);
nor U515 (N_515,In_2074,In_1384);
xnor U516 (N_516,In_2800,In_2316);
nand U517 (N_517,In_765,In_2380);
nand U518 (N_518,In_2606,In_2003);
nand U519 (N_519,In_1332,In_1740);
xor U520 (N_520,In_2740,In_1336);
xnor U521 (N_521,In_2578,In_2869);
nor U522 (N_522,In_539,In_1401);
nor U523 (N_523,In_1291,In_1599);
xor U524 (N_524,In_434,In_749);
nand U525 (N_525,In_513,In_2377);
or U526 (N_526,In_1289,In_2401);
nand U527 (N_527,In_2907,In_854);
xor U528 (N_528,In_2985,In_117);
xor U529 (N_529,In_1717,In_1744);
nor U530 (N_530,In_2819,In_2586);
or U531 (N_531,In_2446,In_1892);
and U532 (N_532,In_887,In_771);
and U533 (N_533,In_1849,In_2669);
nor U534 (N_534,In_1438,In_2424);
nand U535 (N_535,In_2260,In_1109);
or U536 (N_536,In_2986,In_128);
nand U537 (N_537,In_1143,In_892);
or U538 (N_538,In_1064,In_426);
nand U539 (N_539,In_209,In_1718);
nor U540 (N_540,In_1940,In_1175);
xnor U541 (N_541,In_2930,In_161);
nor U542 (N_542,In_2096,In_1155);
xnor U543 (N_543,In_1250,In_2886);
and U544 (N_544,In_417,In_1870);
and U545 (N_545,In_283,In_315);
nor U546 (N_546,In_1739,In_1094);
xor U547 (N_547,In_2736,In_177);
nand U548 (N_548,In_2951,In_2187);
nand U549 (N_549,In_2938,In_2092);
nor U550 (N_550,In_2959,In_75);
nand U551 (N_551,In_2698,In_1257);
nor U552 (N_552,In_1786,In_997);
and U553 (N_553,In_215,In_285);
nand U554 (N_554,In_1407,In_462);
nand U555 (N_555,In_302,In_682);
nor U556 (N_556,In_257,In_2208);
xor U557 (N_557,In_397,In_2119);
nand U558 (N_558,In_1852,In_2711);
nand U559 (N_559,In_1543,In_1964);
nor U560 (N_560,In_583,In_2147);
nor U561 (N_561,In_1881,In_246);
nor U562 (N_562,In_2396,In_2061);
nor U563 (N_563,In_1037,In_16);
nor U564 (N_564,In_2765,In_2334);
and U565 (N_565,In_2799,In_1349);
nor U566 (N_566,In_1856,In_1745);
xnor U567 (N_567,In_808,In_1456);
nor U568 (N_568,In_2221,In_284);
nand U569 (N_569,In_553,In_2579);
nand U570 (N_570,In_2182,In_369);
nor U571 (N_571,In_214,In_2697);
nand U572 (N_572,In_618,In_2155);
xnor U573 (N_573,In_942,In_1813);
and U574 (N_574,In_1381,In_1060);
and U575 (N_575,In_2548,In_89);
or U576 (N_576,In_400,In_1650);
or U577 (N_577,In_8,In_1129);
xor U578 (N_578,In_1273,In_2226);
nor U579 (N_579,In_835,In_2754);
xnor U580 (N_580,In_1082,In_2682);
xnor U581 (N_581,In_1032,In_2781);
and U582 (N_582,In_1271,In_739);
nor U583 (N_583,In_632,In_26);
nand U584 (N_584,In_438,In_888);
or U585 (N_585,In_1481,In_1364);
nor U586 (N_586,In_2240,In_59);
or U587 (N_587,In_535,In_657);
xor U588 (N_588,In_1939,In_312);
and U589 (N_589,In_2287,In_2887);
and U590 (N_590,In_1738,In_111);
xnor U591 (N_591,In_191,In_2925);
xnor U592 (N_592,In_1249,In_1517);
or U593 (N_593,In_360,In_1234);
nor U594 (N_594,In_1775,In_923);
and U595 (N_595,In_2418,In_918);
xnor U596 (N_596,In_1811,In_81);
nor U597 (N_597,In_2325,In_259);
nand U598 (N_598,In_1763,In_1427);
or U599 (N_599,In_1322,In_2436);
nor U600 (N_600,In_500,N_261);
and U601 (N_601,In_2973,In_924);
xnor U602 (N_602,N_537,N_173);
nand U603 (N_603,In_1184,In_2130);
nand U604 (N_604,N_567,In_1435);
and U605 (N_605,In_76,In_2970);
nand U606 (N_606,In_1843,In_348);
or U607 (N_607,In_2152,In_1278);
or U608 (N_608,In_96,In_425);
and U609 (N_609,In_2204,In_2882);
or U610 (N_610,In_2899,In_418);
nand U611 (N_611,In_1077,In_2505);
nor U612 (N_612,In_2752,In_704);
nor U613 (N_613,N_577,N_456);
and U614 (N_614,In_2889,N_357);
nor U615 (N_615,N_215,In_703);
nor U616 (N_616,In_1284,In_2798);
nand U617 (N_617,In_2114,In_2172);
nor U618 (N_618,In_1242,In_243);
or U619 (N_619,In_2404,N_88);
xnor U620 (N_620,In_107,In_2643);
nor U621 (N_621,In_497,In_2927);
or U622 (N_622,In_2900,N_143);
nand U623 (N_623,In_28,In_1999);
and U624 (N_624,N_6,In_244);
nand U625 (N_625,N_449,In_24);
nand U626 (N_626,N_298,In_2444);
nor U627 (N_627,N_218,In_2993);
and U628 (N_628,In_2558,N_312);
and U629 (N_629,N_156,In_1792);
nand U630 (N_630,In_2100,In_796);
xnor U631 (N_631,N_92,In_2099);
nor U632 (N_632,In_47,N_229);
and U633 (N_633,In_1163,In_2838);
xnor U634 (N_634,In_688,N_125);
or U635 (N_635,In_92,N_431);
or U636 (N_636,In_1107,In_1457);
nand U637 (N_637,In_468,In_2319);
nand U638 (N_638,N_410,In_204);
and U639 (N_639,N_323,In_1124);
or U640 (N_640,In_2968,In_828);
nor U641 (N_641,In_1620,N_479);
nor U642 (N_642,In_2879,In_2321);
xor U643 (N_643,In_2077,In_2614);
nor U644 (N_644,N_444,In_2801);
or U645 (N_645,N_251,In_1957);
nand U646 (N_646,In_2000,In_2535);
nor U647 (N_647,In_1552,N_344);
nand U648 (N_648,In_331,In_2365);
or U649 (N_649,In_394,In_1483);
nor U650 (N_650,In_1478,In_1930);
nand U651 (N_651,N_31,In_1316);
and U652 (N_652,In_1312,In_1825);
and U653 (N_653,In_2094,In_2704);
and U654 (N_654,In_2809,In_32);
nor U655 (N_655,In_1056,N_554);
or U656 (N_656,In_700,In_1431);
and U657 (N_657,In_232,In_157);
or U658 (N_658,In_329,In_2739);
nand U659 (N_659,In_2554,N_213);
nor U660 (N_660,N_366,In_1619);
or U661 (N_661,N_560,In_46);
and U662 (N_662,In_651,In_1732);
nor U663 (N_663,N_548,In_2330);
or U664 (N_664,In_1369,N_271);
or U665 (N_665,In_1824,In_882);
xnor U666 (N_666,In_1049,N_30);
nor U667 (N_667,In_1216,In_2143);
nand U668 (N_668,In_2464,In_987);
nor U669 (N_669,N_175,In_1501);
xor U670 (N_670,In_1326,N_230);
xor U671 (N_671,N_249,In_747);
nor U672 (N_672,In_1978,N_399);
and U673 (N_673,In_1862,N_221);
and U674 (N_674,In_901,In_912);
nand U675 (N_675,In_2309,In_2741);
or U676 (N_676,In_406,N_508);
nor U677 (N_677,In_564,In_2425);
nor U678 (N_678,N_140,N_58);
or U679 (N_679,In_540,In_195);
xor U680 (N_680,In_420,N_455);
xor U681 (N_681,In_2218,In_2620);
and U682 (N_682,In_2392,N_561);
or U683 (N_683,In_2596,In_435);
or U684 (N_684,In_1995,In_645);
and U685 (N_685,N_377,In_1161);
nand U686 (N_686,In_1079,In_1658);
and U687 (N_687,N_424,In_779);
xnor U688 (N_688,N_231,N_489);
nor U689 (N_689,In_841,In_821);
xor U690 (N_690,N_549,N_188);
or U691 (N_691,In_931,N_518);
nand U692 (N_692,In_2084,In_615);
xor U693 (N_693,In_1896,In_1075);
nand U694 (N_694,In_1134,In_1637);
or U695 (N_695,In_940,In_2405);
nand U696 (N_696,In_1165,In_2073);
or U697 (N_697,In_1230,N_361);
nor U698 (N_698,In_2737,In_1846);
nor U699 (N_699,N_396,In_1720);
nor U700 (N_700,N_17,In_2479);
xnor U701 (N_701,In_359,N_28);
nand U702 (N_702,N_106,In_2009);
and U703 (N_703,In_100,In_320);
or U704 (N_704,In_2294,In_2706);
or U705 (N_705,In_795,In_365);
nand U706 (N_706,In_313,In_294);
nand U707 (N_707,In_2213,In_322);
or U708 (N_708,In_1841,In_346);
xor U709 (N_709,N_169,In_972);
or U710 (N_710,N_159,In_1396);
or U711 (N_711,In_816,In_1522);
nand U712 (N_712,In_2284,In_408);
nor U713 (N_713,In_2144,In_14);
nor U714 (N_714,In_708,In_2717);
xor U715 (N_715,In_2915,In_217);
nand U716 (N_716,In_1460,In_619);
nand U717 (N_717,In_1753,In_2703);
nand U718 (N_718,N_432,In_558);
xor U719 (N_719,In_719,In_2028);
and U720 (N_720,In_430,N_436);
nand U721 (N_721,N_534,In_452);
nor U722 (N_722,In_2529,In_902);
nor U723 (N_723,N_382,In_1602);
or U724 (N_724,N_400,In_197);
and U725 (N_725,In_678,In_1800);
nand U726 (N_726,N_503,In_851);
and U727 (N_727,In_1025,N_598);
xnor U728 (N_728,N_395,In_22);
and U729 (N_729,In_636,In_1212);
xor U730 (N_730,In_566,N_355);
nand U731 (N_731,In_1987,N_56);
xnor U732 (N_732,N_520,N_36);
nor U733 (N_733,In_1145,In_104);
nor U734 (N_734,In_86,In_715);
nand U735 (N_735,N_433,In_1319);
xor U736 (N_736,N_329,In_1022);
and U737 (N_737,In_1894,In_2413);
xnor U738 (N_738,In_2910,In_1961);
and U739 (N_739,In_2054,In_1771);
nor U740 (N_740,In_38,N_69);
nor U741 (N_741,In_2460,In_272);
and U742 (N_742,In_1499,In_68);
and U743 (N_743,In_2306,In_1615);
nand U744 (N_744,N_314,In_1018);
and U745 (N_745,In_1213,In_446);
and U746 (N_746,In_7,In_2881);
or U747 (N_747,N_494,In_1872);
nor U748 (N_748,In_2482,In_1573);
and U749 (N_749,In_1564,In_1480);
nor U750 (N_750,N_225,In_290);
xor U751 (N_751,N_597,In_1180);
nor U752 (N_752,In_2267,In_206);
xnor U753 (N_753,In_1633,In_1762);
and U754 (N_754,In_2746,In_1437);
or U755 (N_755,In_1848,In_475);
and U756 (N_756,In_353,In_1303);
xor U757 (N_757,In_114,In_2322);
nand U758 (N_758,In_192,N_304);
xnor U759 (N_759,N_168,In_1698);
or U760 (N_760,In_1063,N_542);
and U761 (N_761,N_599,In_2489);
nor U762 (N_762,N_320,In_1496);
nand U763 (N_763,In_2770,In_1784);
nand U764 (N_764,N_319,In_440);
nor U765 (N_765,In_551,In_1844);
and U766 (N_766,N_420,In_343);
and U767 (N_767,In_2192,N_48);
nand U768 (N_768,In_2441,In_768);
nor U769 (N_769,In_2052,In_2462);
nand U770 (N_770,N_325,N_59);
nor U771 (N_771,N_16,In_1597);
nand U772 (N_772,In_2120,N_318);
nor U773 (N_773,In_1623,In_834);
xnor U774 (N_774,N_219,In_2257);
nor U775 (N_775,In_263,In_1497);
and U776 (N_776,In_1452,In_701);
and U777 (N_777,In_1672,In_321);
nand U778 (N_778,In_1128,N_281);
nand U779 (N_779,N_486,In_1357);
or U780 (N_780,In_1047,N_543);
and U781 (N_781,N_544,In_1831);
and U782 (N_782,N_85,In_2580);
xnor U783 (N_783,In_2443,In_2629);
nand U784 (N_784,In_2228,In_1399);
nand U785 (N_785,N_513,In_165);
nor U786 (N_786,In_1861,In_1899);
nor U787 (N_787,N_521,N_397);
nand U788 (N_788,In_1173,N_354);
or U789 (N_789,N_475,In_784);
nor U790 (N_790,N_47,In_2366);
and U791 (N_791,In_811,N_52);
nand U792 (N_792,In_2179,In_2618);
and U793 (N_793,In_198,N_303);
xnor U794 (N_794,N_63,In_455);
nor U795 (N_795,In_492,In_2591);
or U796 (N_796,In_2364,In_121);
nor U797 (N_797,In_519,N_256);
and U798 (N_798,In_1237,N_19);
nor U799 (N_799,N_501,In_1426);
and U800 (N_800,In_1834,In_53);
nor U801 (N_801,In_1115,In_1967);
or U802 (N_802,In_2363,In_801);
and U803 (N_803,In_1601,In_2211);
and U804 (N_804,In_2210,N_406);
and U805 (N_805,In_2430,N_147);
nand U806 (N_806,In_1789,N_102);
nand U807 (N_807,In_485,In_2036);
xnor U808 (N_808,In_1002,In_282);
or U809 (N_809,N_3,In_954);
nand U810 (N_810,In_1703,N_488);
and U811 (N_811,N_290,In_484);
xor U812 (N_812,N_13,In_450);
xor U813 (N_813,In_1808,In_1360);
or U814 (N_814,In_73,In_850);
nand U815 (N_815,In_866,In_2855);
or U816 (N_816,N_421,In_2965);
or U817 (N_817,N_524,In_2572);
nand U818 (N_818,N_50,In_501);
xnor U819 (N_819,In_790,In_2632);
nor U820 (N_820,N_286,In_2345);
xnor U821 (N_821,N_117,N_481);
xor U822 (N_822,In_1730,In_2387);
and U823 (N_823,In_1304,In_488);
nand U824 (N_824,N_44,In_2010);
nor U825 (N_825,In_785,N_33);
and U826 (N_826,N_95,N_1);
or U827 (N_827,In_2696,N_226);
and U828 (N_828,In_1149,In_469);
nand U829 (N_829,In_783,In_2421);
nor U830 (N_830,In_755,In_1743);
nand U831 (N_831,In_50,In_399);
nor U832 (N_832,N_104,In_384);
nor U833 (N_833,In_1812,In_1301);
nor U834 (N_834,In_2834,N_330);
xnor U835 (N_835,In_612,N_482);
and U836 (N_836,In_1551,In_176);
nor U837 (N_837,N_301,In_948);
or U838 (N_838,N_233,In_1997);
and U839 (N_839,In_712,In_2300);
or U840 (N_840,N_239,In_897);
or U841 (N_841,N_97,In_2540);
or U842 (N_842,N_538,In_222);
xor U843 (N_843,In_980,In_1067);
or U844 (N_844,In_90,In_1338);
nor U845 (N_845,In_1897,In_1409);
and U846 (N_846,In_1963,In_1411);
xor U847 (N_847,In_471,In_1928);
xor U848 (N_848,In_809,In_2532);
xor U849 (N_849,In_2469,In_67);
nand U850 (N_850,N_582,In_2901);
xnor U851 (N_851,In_1355,In_839);
xor U852 (N_852,In_2519,In_2050);
and U853 (N_853,In_1903,In_1343);
and U854 (N_854,In_1455,In_1674);
and U855 (N_855,In_521,In_273);
nor U856 (N_856,In_1778,In_2005);
and U857 (N_857,N_587,N_161);
xnor U858 (N_858,In_1090,In_2127);
and U859 (N_859,In_60,In_634);
xnor U860 (N_860,In_1616,In_2026);
nand U861 (N_861,In_732,N_437);
xor U862 (N_862,In_638,In_275);
nand U863 (N_863,In_707,In_79);
or U864 (N_864,N_465,In_1096);
and U865 (N_865,In_266,In_2432);
nor U866 (N_866,In_870,In_758);
or U867 (N_867,In_1595,In_2434);
nand U868 (N_868,In_907,In_2348);
nor U869 (N_869,N_187,N_162);
and U870 (N_870,In_1281,In_617);
or U871 (N_871,In_422,N_321);
or U872 (N_872,In_2467,N_42);
or U873 (N_873,In_87,In_182);
or U874 (N_874,In_1057,In_578);
xor U875 (N_875,N_84,N_530);
and U876 (N_876,In_358,In_2958);
xnor U877 (N_877,In_1810,In_2264);
nor U878 (N_878,In_2448,In_1171);
nor U879 (N_879,N_458,N_464);
xnor U880 (N_880,In_1933,In_1509);
nand U881 (N_881,N_242,N_576);
nand U882 (N_882,N_123,In_508);
nand U883 (N_883,In_151,N_250);
xor U884 (N_884,In_1641,In_2379);
and U885 (N_885,N_365,In_1404);
or U886 (N_886,N_510,In_2842);
and U887 (N_887,N_566,In_919);
xnor U888 (N_888,In_873,In_1913);
or U889 (N_889,N_201,In_1561);
or U890 (N_890,In_2158,In_180);
nand U891 (N_891,In_2249,In_714);
xor U892 (N_892,N_454,In_120);
or U893 (N_893,In_130,In_1196);
nand U894 (N_894,In_2415,In_1765);
and U895 (N_895,In_2019,In_1506);
and U896 (N_896,N_183,N_490);
or U897 (N_897,In_1660,In_531);
xnor U898 (N_898,In_494,In_2615);
nand U899 (N_899,In_57,In_598);
or U900 (N_900,In_1984,In_2921);
xor U901 (N_901,In_333,In_2994);
nand U902 (N_902,In_1074,In_1085);
or U903 (N_903,In_694,In_1498);
and U904 (N_904,In_2341,N_374);
nand U905 (N_905,In_635,In_332);
nor U906 (N_906,In_2078,In_1714);
or U907 (N_907,In_2644,In_1610);
and U908 (N_908,In_1133,In_63);
or U909 (N_909,In_2599,In_561);
nand U910 (N_910,In_1131,In_2331);
nand U911 (N_911,In_2382,N_402);
nand U912 (N_912,In_2566,In_1140);
nor U913 (N_913,In_936,In_1302);
nor U914 (N_914,In_1038,In_576);
nand U915 (N_915,N_211,N_536);
or U916 (N_916,N_166,In_991);
and U917 (N_917,N_345,In_1324);
and U918 (N_918,In_1253,In_587);
xor U919 (N_919,In_2847,N_99);
and U920 (N_920,In_1890,N_322);
nand U921 (N_921,N_267,N_174);
or U922 (N_922,In_2180,In_817);
xor U923 (N_923,In_2483,In_2243);
or U924 (N_924,N_531,N_372);
or U925 (N_925,In_2251,In_2118);
and U926 (N_926,In_1955,In_1053);
nor U927 (N_927,N_506,N_282);
nand U928 (N_928,In_1141,In_2836);
and U929 (N_929,In_2166,In_337);
xnor U930 (N_930,N_185,N_388);
xor U931 (N_931,In_1608,In_310);
xnor U932 (N_932,N_210,In_2242);
xor U933 (N_933,N_40,In_451);
xor U934 (N_934,In_2250,In_756);
nor U935 (N_935,In_1941,In_2946);
nor U936 (N_936,In_200,In_857);
and U937 (N_937,In_1532,N_568);
nor U938 (N_938,In_1306,N_160);
or U939 (N_939,N_578,In_2055);
or U940 (N_940,N_62,In_2275);
nor U941 (N_941,In_70,In_746);
nor U942 (N_942,In_169,In_751);
nand U943 (N_943,N_283,N_83);
nor U944 (N_944,In_1685,N_404);
xnor U945 (N_945,In_1419,N_197);
or U946 (N_946,In_640,In_894);
and U947 (N_947,In_110,In_1719);
nor U948 (N_948,In_1008,In_1076);
xnor U949 (N_949,In_1525,In_1181);
or U950 (N_950,In_256,In_230);
xor U951 (N_951,In_2521,In_1785);
and U952 (N_952,In_402,In_1300);
xor U953 (N_953,In_467,In_2870);
and U954 (N_954,N_463,In_1567);
and U955 (N_955,In_196,In_1756);
xor U956 (N_956,In_742,In_798);
nor U957 (N_957,N_53,In_2640);
nand U958 (N_958,In_2776,N_77);
nor U959 (N_959,In_208,In_679);
xor U960 (N_960,In_66,In_2107);
or U961 (N_961,N_558,In_2344);
nand U962 (N_962,N_109,In_1707);
nor U963 (N_963,N_335,In_1910);
and U964 (N_964,In_1222,In_730);
nor U965 (N_965,In_2150,In_2635);
xnor U966 (N_966,In_2326,In_2222);
or U967 (N_967,In_292,In_2686);
nor U968 (N_968,N_559,In_2063);
or U969 (N_969,In_2235,N_180);
nor U970 (N_970,In_2327,N_352);
nor U971 (N_971,N_435,N_403);
xnor U972 (N_972,In_1097,In_2767);
or U973 (N_973,In_662,N_150);
xor U974 (N_974,In_274,In_432);
nand U975 (N_975,In_1371,In_1924);
nand U976 (N_976,In_1956,In_2585);
or U977 (N_977,N_541,In_1511);
xnor U978 (N_978,In_219,In_2622);
or U979 (N_979,In_2025,In_142);
nand U980 (N_980,In_1931,In_1380);
nand U981 (N_981,In_2963,In_2846);
xor U982 (N_982,N_54,In_491);
and U983 (N_983,N_253,N_555);
xor U984 (N_984,N_324,In_2974);
and U985 (N_985,In_2785,In_1968);
xnor U986 (N_986,In_122,In_807);
nor U987 (N_987,N_184,In_1445);
nand U988 (N_988,N_466,In_1798);
xnor U989 (N_989,In_2624,In_155);
nand U990 (N_990,In_2207,N_473);
nor U991 (N_991,In_903,In_1854);
and U992 (N_992,In_1548,N_347);
xor U993 (N_993,In_630,In_1217);
nand U994 (N_994,N_423,N_21);
xnor U995 (N_995,In_2676,In_1295);
xnor U996 (N_996,N_516,In_1087);
and U997 (N_997,In_2619,N_198);
and U998 (N_998,In_502,In_1359);
xnor U999 (N_999,In_1309,N_522);
xnor U1000 (N_1000,In_760,In_2169);
xnor U1001 (N_1001,In_1393,In_1871);
nand U1002 (N_1002,In_1642,In_2610);
xor U1003 (N_1003,In_549,In_2449);
and U1004 (N_1004,In_2281,In_1153);
nor U1005 (N_1005,N_540,In_2481);
xnor U1006 (N_1006,In_187,In_1558);
nor U1007 (N_1007,In_2690,N_280);
or U1008 (N_1008,N_585,In_584);
nor U1009 (N_1009,In_238,In_1440);
and U1010 (N_1010,In_1606,In_571);
xnor U1011 (N_1011,N_378,In_1026);
and U1012 (N_1012,In_1603,N_177);
xnor U1013 (N_1013,N_467,In_932);
or U1014 (N_1014,In_674,In_1379);
or U1015 (N_1015,N_206,N_93);
nand U1016 (N_1016,In_526,N_70);
nand U1017 (N_1017,In_2034,N_235);
nor U1018 (N_1018,N_105,In_2914);
nor U1019 (N_1019,In_506,N_39);
nand U1020 (N_1020,In_258,In_2439);
and U1021 (N_1021,In_2749,In_1575);
or U1022 (N_1022,In_1110,N_269);
and U1023 (N_1023,In_2598,In_2008);
nor U1024 (N_1024,In_349,In_2156);
nor U1025 (N_1025,In_1746,N_333);
xnor U1026 (N_1026,In_2245,N_20);
xnor U1027 (N_1027,In_1463,In_2305);
nand U1028 (N_1028,N_119,N_358);
or U1029 (N_1029,In_2719,In_2672);
and U1030 (N_1030,In_1340,In_1033);
xnor U1031 (N_1031,N_340,N_373);
and U1032 (N_1032,In_1232,N_375);
or U1033 (N_1033,In_2450,In_94);
nand U1034 (N_1034,In_1243,In_37);
and U1035 (N_1035,In_54,In_2016);
nand U1036 (N_1036,In_140,N_474);
or U1037 (N_1037,In_479,In_1199);
nand U1038 (N_1038,In_2813,In_2545);
or U1039 (N_1039,In_1104,In_740);
nand U1040 (N_1040,In_838,In_620);
or U1041 (N_1041,In_2733,In_1174);
xnor U1042 (N_1042,N_457,In_316);
xnor U1043 (N_1043,N_11,In_767);
nor U1044 (N_1044,In_2570,In_1314);
nand U1045 (N_1045,In_171,In_753);
nor U1046 (N_1046,N_580,In_570);
and U1047 (N_1047,In_2072,N_480);
or U1048 (N_1048,N_381,In_1029);
nor U1049 (N_1049,In_1737,In_2601);
nand U1050 (N_1050,N_418,N_535);
or U1051 (N_1051,In_1761,In_2032);
and U1052 (N_1052,N_279,In_616);
or U1053 (N_1053,N_469,In_2411);
or U1054 (N_1054,In_2639,In_2786);
nand U1055 (N_1055,In_1207,In_2667);
xor U1056 (N_1056,N_278,N_337);
and U1057 (N_1057,In_602,In_1750);
and U1058 (N_1058,In_2528,In_2674);
nand U1059 (N_1059,In_1330,In_1927);
or U1060 (N_1060,In_2121,In_2738);
xor U1061 (N_1061,In_975,In_1842);
nand U1062 (N_1062,N_129,In_1410);
and U1063 (N_1063,In_398,In_2630);
and U1064 (N_1064,In_2337,In_362);
xor U1065 (N_1065,In_224,In_2362);
and U1066 (N_1066,In_388,N_359);
and U1067 (N_1067,In_2852,N_200);
nor U1068 (N_1068,In_1132,In_2037);
or U1069 (N_1069,N_67,In_1721);
nand U1070 (N_1070,N_342,In_1358);
or U1071 (N_1071,In_2435,N_583);
nand U1072 (N_1072,In_2772,N_348);
or U1073 (N_1073,In_239,N_430);
xor U1074 (N_1074,In_1943,In_1003);
nand U1075 (N_1075,In_2942,In_1311);
nand U1076 (N_1076,In_1902,In_522);
xor U1077 (N_1077,In_908,In_2431);
or U1078 (N_1078,In_2420,In_2547);
xnor U1079 (N_1079,In_2924,In_652);
xnor U1080 (N_1080,In_2634,N_80);
and U1081 (N_1081,In_247,In_2161);
xor U1082 (N_1082,In_174,In_1327);
and U1083 (N_1083,In_2470,In_1555);
nand U1084 (N_1084,N_252,In_960);
and U1085 (N_1085,In_2678,In_757);
xor U1086 (N_1086,In_766,In_1580);
or U1087 (N_1087,In_445,N_452);
or U1088 (N_1088,N_25,N_426);
nand U1089 (N_1089,In_1121,N_514);
or U1090 (N_1090,In_2237,In_2079);
nor U1091 (N_1091,In_2186,In_1433);
xnor U1092 (N_1092,In_2040,In_2057);
nand U1093 (N_1093,In_382,In_1287);
nand U1094 (N_1094,In_2006,In_347);
nand U1095 (N_1095,In_2665,In_1394);
nand U1096 (N_1096,In_2911,In_2053);
or U1097 (N_1097,N_383,In_1268);
and U1098 (N_1098,In_961,N_208);
or U1099 (N_1099,In_2102,In_298);
and U1100 (N_1100,In_1832,In_2751);
and U1101 (N_1101,In_1830,In_2663);
and U1102 (N_1102,In_585,N_8);
nand U1103 (N_1103,In_1605,In_2083);
and U1104 (N_1104,In_1709,In_1389);
nor U1105 (N_1105,N_72,In_2992);
or U1106 (N_1106,In_2395,In_1559);
xor U1107 (N_1107,In_2030,In_920);
nor U1108 (N_1108,N_511,N_157);
xor U1109 (N_1109,In_376,N_527);
xor U1110 (N_1110,In_1847,In_1621);
nand U1111 (N_1111,In_927,In_2324);
xnor U1112 (N_1112,In_614,In_2508);
nand U1113 (N_1113,In_2936,In_577);
or U1114 (N_1114,In_2997,N_75);
nor U1115 (N_1115,In_1991,In_2561);
or U1116 (N_1116,In_1816,In_395);
xnor U1117 (N_1117,In_2419,In_528);
nand U1118 (N_1118,In_670,In_2700);
or U1119 (N_1119,In_1932,In_1469);
xnor U1120 (N_1120,In_824,In_392);
xor U1121 (N_1121,In_844,In_2718);
or U1122 (N_1122,In_1611,In_1876);
nand U1123 (N_1123,N_369,N_419);
xnor U1124 (N_1124,N_307,In_820);
and U1125 (N_1125,In_1985,In_2712);
nand U1126 (N_1126,N_153,In_946);
nor U1127 (N_1127,In_1908,In_973);
nand U1128 (N_1128,N_248,N_356);
and U1129 (N_1129,In_56,In_2279);
nor U1130 (N_1130,In_1422,In_72);
nor U1131 (N_1131,In_1244,N_491);
or U1132 (N_1132,In_565,In_2151);
nand U1133 (N_1133,In_969,N_152);
nand U1134 (N_1134,In_1676,In_910);
nor U1135 (N_1135,In_2320,In_1769);
or U1136 (N_1136,In_529,In_2814);
xnor U1137 (N_1137,N_429,In_2133);
or U1138 (N_1138,N_82,In_532);
and U1139 (N_1139,In_958,In_495);
nor U1140 (N_1140,N_478,In_1488);
nor U1141 (N_1141,In_1052,In_1251);
nor U1142 (N_1142,In_1593,In_2880);
nor U1143 (N_1143,In_2291,N_29);
xnor U1144 (N_1144,N_194,In_251);
or U1145 (N_1145,In_963,In_2511);
nand U1146 (N_1146,N_592,In_2788);
xor U1147 (N_1147,In_926,In_1494);
or U1148 (N_1148,In_2056,In_745);
nand U1149 (N_1149,In_2476,In_1628);
nand U1150 (N_1150,In_172,N_110);
xor U1151 (N_1151,In_2920,In_1254);
and U1152 (N_1152,In_1261,In_1021);
nand U1153 (N_1153,In_503,In_1822);
and U1154 (N_1154,In_386,N_351);
or U1155 (N_1155,In_786,In_2280);
nand U1156 (N_1156,In_2177,In_1105);
and U1157 (N_1157,N_398,In_2175);
nand U1158 (N_1158,N_234,N_66);
and U1159 (N_1159,In_25,In_474);
and U1160 (N_1160,In_2861,In_184);
nor U1161 (N_1161,In_2494,In_1915);
or U1162 (N_1162,In_1748,In_1736);
nor U1163 (N_1163,In_1929,In_1592);
xor U1164 (N_1164,In_2944,N_199);
and U1165 (N_1165,In_2039,In_527);
xnor U1166 (N_1166,In_188,In_1101);
xor U1167 (N_1167,In_2940,In_2191);
xnor U1168 (N_1168,N_434,N_460);
nor U1169 (N_1169,In_2796,N_257);
or U1170 (N_1170,N_384,In_1477);
or U1171 (N_1171,In_959,In_706);
nor U1172 (N_1172,In_812,In_2787);
and U1173 (N_1173,In_992,In_1617);
nor U1174 (N_1174,In_930,N_512);
and U1175 (N_1175,N_146,In_1827);
and U1176 (N_1176,In_2966,In_1139);
xnor U1177 (N_1177,N_499,In_557);
nand U1178 (N_1178,N_350,In_646);
nand U1179 (N_1179,In_2129,In_1315);
or U1180 (N_1180,In_2671,In_2952);
nor U1181 (N_1181,N_367,In_1436);
xor U1182 (N_1182,N_422,In_2500);
nor U1183 (N_1183,N_51,N_32);
xnor U1184 (N_1184,In_2136,In_164);
xor U1185 (N_1185,In_2278,In_2909);
or U1186 (N_1186,In_2784,In_2312);
nor U1187 (N_1187,In_928,In_2531);
nor U1188 (N_1188,N_428,In_1120);
xnor U1189 (N_1189,In_1513,In_2661);
and U1190 (N_1190,In_2565,N_24);
nor U1191 (N_1191,N_588,In_372);
nand U1192 (N_1192,In_2254,N_222);
or U1193 (N_1193,In_2931,In_1946);
xor U1194 (N_1194,N_263,In_1646);
nor U1195 (N_1195,In_2975,In_2023);
nand U1196 (N_1196,In_2550,In_1484);
nand U1197 (N_1197,In_569,In_421);
nand U1198 (N_1198,In_1716,In_2683);
xnor U1199 (N_1199,In_2196,N_164);
or U1200 (N_1200,In_2829,N_961);
or U1201 (N_1201,N_880,In_106);
or U1202 (N_1202,In_1069,N_1043);
or U1203 (N_1203,In_2722,In_2742);
or U1204 (N_1204,N_634,N_882);
or U1205 (N_1205,In_2022,In_716);
or U1206 (N_1206,N_791,N_780);
or U1207 (N_1207,In_473,N_932);
nor U1208 (N_1208,N_858,N_1110);
and U1209 (N_1209,N_68,N_1050);
xor U1210 (N_1210,N_529,N_892);
nand U1211 (N_1211,N_617,N_684);
and U1212 (N_1212,N_1020,In_516);
nand U1213 (N_1213,N_731,In_1855);
or U1214 (N_1214,In_1518,In_2115);
nor U1215 (N_1215,N_616,N_1082);
or U1216 (N_1216,In_496,In_2378);
or U1217 (N_1217,N_795,In_2831);
nor U1218 (N_1218,N_755,N_631);
and U1219 (N_1219,N_891,In_1937);
or U1220 (N_1220,In_178,In_1521);
nor U1221 (N_1221,N_1174,N_942);
xnor U1222 (N_1222,In_2389,N_1091);
and U1223 (N_1223,N_713,In_2769);
xnor U1224 (N_1224,N_295,In_2159);
nor U1225 (N_1225,In_1366,In_340);
xor U1226 (N_1226,N_1055,N_142);
nor U1227 (N_1227,In_1489,In_2406);
or U1228 (N_1228,N_132,In_1588);
or U1229 (N_1229,In_1065,In_953);
or U1230 (N_1230,N_816,In_832);
and U1231 (N_1231,N_22,N_872);
nand U1232 (N_1232,In_2007,In_1449);
xnor U1233 (N_1233,In_2352,N_796);
nor U1234 (N_1234,In_2433,N_1051);
or U1235 (N_1235,N_601,N_37);
nor U1236 (N_1236,N_1029,In_252);
or U1237 (N_1237,N_993,N_845);
and U1238 (N_1238,In_248,N_1073);
and U1239 (N_1239,N_732,N_472);
or U1240 (N_1240,In_2353,In_1159);
or U1241 (N_1241,N_861,In_2933);
and U1242 (N_1242,N_43,In_886);
xor U1243 (N_1243,In_1524,N_1158);
or U1244 (N_1244,N_504,N_1068);
nor U1245 (N_1245,N_76,In_2116);
and U1246 (N_1246,N_1098,In_770);
or U1247 (N_1247,In_957,In_2113);
nor U1248 (N_1248,N_386,In_2502);
and U1249 (N_1249,N_931,In_2185);
nand U1250 (N_1250,In_2525,In_141);
and U1251 (N_1251,N_744,In_478);
nand U1252 (N_1252,N_862,In_2445);
xnor U1253 (N_1253,In_1505,In_2652);
xor U1254 (N_1254,In_2101,N_1173);
nand U1255 (N_1255,N_824,In_3);
and U1256 (N_1256,N_991,N_784);
or U1257 (N_1257,N_608,In_933);
xnor U1258 (N_1258,N_822,In_88);
and U1259 (N_1259,N_708,In_533);
or U1260 (N_1260,In_131,In_885);
or U1261 (N_1261,N_1089,N_607);
xor U1262 (N_1262,N_651,N_1131);
and U1263 (N_1263,In_1547,N_644);
nor U1264 (N_1264,N_4,N_407);
nand U1265 (N_1265,In_2343,N_694);
nand U1266 (N_1266,In_1299,In_1508);
xor U1267 (N_1267,In_512,N_777);
nand U1268 (N_1268,In_27,N_647);
nand U1269 (N_1269,N_370,N_986);
xor U1270 (N_1270,N_1074,In_1323);
and U1271 (N_1271,N_526,N_451);
and U1272 (N_1272,N_829,N_507);
xnor U1273 (N_1273,N_998,N_662);
nor U1274 (N_1274,In_2982,N_1159);
nand U1275 (N_1275,In_2872,N_950);
nor U1276 (N_1276,In_2426,N_1057);
nand U1277 (N_1277,N_1097,In_2792);
nand U1278 (N_1278,N_679,N_984);
and U1279 (N_1279,In_216,N_293);
nand U1280 (N_1280,In_1368,N_214);
nand U1281 (N_1281,N_96,In_1749);
nor U1282 (N_1282,In_2386,In_2217);
or U1283 (N_1283,In_2649,N_889);
or U1284 (N_1284,N_1054,In_717);
or U1285 (N_1285,In_2014,In_1308);
nor U1286 (N_1286,In_2487,N_115);
xnor U1287 (N_1287,In_789,In_223);
nand U1288 (N_1288,In_377,N_774);
nand U1289 (N_1289,In_2757,N_41);
xnor U1290 (N_1290,N_888,N_1126);
nor U1291 (N_1291,In_2241,N_1161);
nand U1292 (N_1292,In_697,N_120);
nor U1293 (N_1293,N_854,In_2650);
nand U1294 (N_1294,In_1783,N_807);
xnor U1295 (N_1295,N_1064,N_877);
nand U1296 (N_1296,In_2484,N_638);
nand U1297 (N_1297,N_154,In_1880);
nor U1298 (N_1298,In_1182,In_968);
and U1299 (N_1299,N_772,In_1972);
nand U1300 (N_1300,In_669,In_2812);
or U1301 (N_1301,In_383,N_627);
xnor U1302 (N_1302,N_1199,N_1092);
or U1303 (N_1303,In_339,N_1164);
xor U1304 (N_1304,In_1965,In_1352);
nor U1305 (N_1305,N_1053,N_91);
nor U1306 (N_1306,In_1320,N_1077);
or U1307 (N_1307,N_287,N_757);
xnor U1308 (N_1308,In_1007,In_1969);
nand U1309 (N_1309,In_379,N_232);
and U1310 (N_1310,In_466,N_116);
xor U1311 (N_1311,N_268,N_866);
nor U1312 (N_1312,N_1099,In_1183);
nor U1313 (N_1313,In_2367,In_1747);
nand U1314 (N_1314,In_2490,In_2097);
or U1315 (N_1315,In_1882,N_971);
nand U1316 (N_1316,N_205,N_939);
nor U1317 (N_1317,In_1790,In_641);
or U1318 (N_1318,In_2391,N_1115);
xor U1319 (N_1319,In_2844,In_314);
nand U1320 (N_1320,N_666,In_1947);
or U1321 (N_1321,In_2289,N_111);
and U1322 (N_1322,N_118,N_1156);
nand U1323 (N_1323,In_1679,N_596);
and U1324 (N_1324,N_1113,In_1689);
or U1325 (N_1325,N_885,In_2018);
nor U1326 (N_1326,N_1128,N_296);
nor U1327 (N_1327,In_608,In_1624);
xor U1328 (N_1328,N_415,In_2664);
nand U1329 (N_1329,In_523,In_2371);
nand U1330 (N_1330,N_1137,N_705);
and U1331 (N_1331,In_2636,N_525);
nor U1332 (N_1332,In_1804,N_837);
or U1333 (N_1333,N_1080,In_2662);
or U1334 (N_1334,In_650,In_1632);
nand U1335 (N_1335,In_1043,N_620);
xnor U1336 (N_1336,In_842,N_690);
nand U1337 (N_1337,N_202,N_167);
xnor U1338 (N_1338,In_2894,N_1177);
nand U1339 (N_1339,In_2299,In_1670);
nand U1340 (N_1340,N_751,N_835);
or U1341 (N_1341,In_2292,In_1663);
nand U1342 (N_1342,In_487,N_646);
xnor U1343 (N_1343,In_698,In_2957);
or U1344 (N_1344,N_960,In_2948);
and U1345 (N_1345,N_1135,In_1728);
xnor U1346 (N_1346,N_1008,In_1500);
or U1347 (N_1347,In_1626,In_370);
or U1348 (N_1348,In_498,N_346);
nor U1349 (N_1349,N_803,N_952);
and U1350 (N_1350,N_45,In_1889);
nor U1351 (N_1351,N_302,In_2167);
or U1352 (N_1352,In_780,N_747);
xor U1353 (N_1353,N_775,In_600);
and U1354 (N_1354,N_1124,In_1589);
nand U1355 (N_1355,In_319,N_575);
and U1356 (N_1356,In_389,In_2577);
or U1357 (N_1357,In_2225,In_1960);
nand U1358 (N_1358,N_155,N_637);
and U1359 (N_1359,N_1035,In_1259);
nor U1360 (N_1360,N_1109,In_791);
nor U1361 (N_1361,N_341,N_810);
nand U1362 (N_1362,N_812,N_254);
xnor U1363 (N_1363,In_2202,In_2555);
xor U1364 (N_1364,N_1023,In_441);
nand U1365 (N_1365,N_918,N_310);
xor U1366 (N_1366,In_884,In_1050);
nor U1367 (N_1367,N_1007,N_767);
nor U1368 (N_1368,N_672,In_1370);
nand U1369 (N_1369,In_2456,N_18);
nand U1370 (N_1370,In_1103,In_2223);
nor U1371 (N_1371,In_2538,In_51);
or U1372 (N_1372,In_647,N_745);
xnor U1373 (N_1373,N_1180,In_663);
nor U1374 (N_1374,In_1385,N_1154);
xor U1375 (N_1375,N_158,N_923);
nand U1376 (N_1376,In_1806,N_414);
xor U1377 (N_1377,N_228,In_448);
nor U1378 (N_1378,In_404,N_590);
or U1379 (N_1379,In_481,N_1056);
or U1380 (N_1380,N_258,In_966);
or U1381 (N_1381,In_2011,N_121);
nand U1382 (N_1382,N_921,In_2122);
and U1383 (N_1383,N_338,N_392);
xnor U1384 (N_1384,In_1328,In_401);
nand U1385 (N_1385,In_490,In_2808);
nor U1386 (N_1386,N_217,In_344);
nor U1387 (N_1387,N_847,N_483);
nor U1388 (N_1388,In_925,In_1935);
nand U1389 (N_1389,N_740,In_2954);
xnor U1390 (N_1390,N_959,N_60);
and U1391 (N_1391,N_523,N_179);
nor U1392 (N_1392,In_644,N_145);
nor U1393 (N_1393,In_922,N_216);
and U1394 (N_1394,In_2729,N_593);
and U1395 (N_1395,N_443,In_1815);
nor U1396 (N_1396,N_1072,In_2131);
nor U1397 (N_1397,N_640,In_1700);
nor U1398 (N_1398,N_461,N_779);
and U1399 (N_1399,In_1290,In_1839);
and U1400 (N_1400,In_115,N_987);
or U1401 (N_1401,N_255,In_1540);
nand U1402 (N_1402,In_147,N_227);
or U1403 (N_1403,N_73,In_2526);
or U1404 (N_1404,In_915,In_80);
nor U1405 (N_1405,N_911,N_1017);
and U1406 (N_1406,N_934,In_137);
or U1407 (N_1407,N_725,In_2233);
nand U1408 (N_1408,In_1005,N_313);
nand U1409 (N_1409,In_41,In_613);
and U1410 (N_1410,In_1068,In_2647);
nand U1411 (N_1411,N_291,In_2745);
nand U1412 (N_1412,N_393,In_269);
nor U1413 (N_1413,N_799,In_1760);
or U1414 (N_1414,N_193,N_976);
nor U1415 (N_1415,N_364,In_596);
and U1416 (N_1416,In_860,N_759);
nor U1417 (N_1417,N_438,In_150);
nand U1418 (N_1418,In_1673,N_935);
or U1419 (N_1419,N_741,N_834);
nor U1420 (N_1420,N_754,In_1528);
xor U1421 (N_1421,In_2783,N_746);
nand U1422 (N_1422,In_574,In_1054);
nand U1423 (N_1423,In_2833,In_622);
nor U1424 (N_1424,N_1081,N_753);
nor U1425 (N_1425,In_1704,N_852);
and U1426 (N_1426,N_979,N_1048);
or U1427 (N_1427,N_814,In_375);
xor U1428 (N_1428,In_1,In_2600);
and U1429 (N_1429,In_1919,In_867);
or U1430 (N_1430,N_865,N_1075);
and U1431 (N_1431,N_220,N_652);
and U1432 (N_1432,In_1045,N_1165);
and U1433 (N_1433,N_988,In_1214);
xor U1434 (N_1434,N_655,In_580);
xor U1435 (N_1435,In_1836,In_1942);
nor U1436 (N_1436,N_697,N_71);
or U1437 (N_1437,N_1170,N_446);
xnor U1438 (N_1438,In_185,N_417);
or U1439 (N_1439,In_2473,In_2735);
nor U1440 (N_1440,In_374,N_843);
nor U1441 (N_1441,N_528,N_1150);
xnor U1442 (N_1442,N_682,In_2359);
and U1443 (N_1443,In_2658,N_928);
xnor U1444 (N_1444,In_1185,N_792);
and U1445 (N_1445,In_1386,N_665);
xnor U1446 (N_1446,N_609,In_36);
and U1447 (N_1447,In_2451,N_898);
and U1448 (N_1448,In_1313,In_1390);
or U1449 (N_1449,N_624,N_1069);
or U1450 (N_1450,N_462,N_305);
nand U1451 (N_1451,N_496,N_1139);
or U1452 (N_1452,N_860,N_1021);
and U1453 (N_1453,In_1265,In_336);
or U1454 (N_1454,In_1690,In_2486);
nor U1455 (N_1455,In_1572,N_308);
nor U1456 (N_1456,N_1146,N_112);
or U1457 (N_1457,N_277,In_2268);
and U1458 (N_1458,N_962,N_656);
or U1459 (N_1459,N_981,N_736);
or U1460 (N_1460,In_676,N_1189);
xor U1461 (N_1461,In_1838,In_1545);
and U1462 (N_1462,N_387,N_353);
nand U1463 (N_1463,In_659,N_447);
or U1464 (N_1464,In_2648,N_1120);
and U1465 (N_1465,N_711,In_2979);
xnor U1466 (N_1466,N_833,N_244);
nor U1467 (N_1467,In_2835,N_236);
xor U1468 (N_1468,In_2273,N_768);
nor U1469 (N_1469,In_1622,In_2568);
or U1470 (N_1470,In_2498,In_871);
or U1471 (N_1471,N_701,N_9);
nand U1472 (N_1472,N_964,N_1012);
xor U1473 (N_1473,N_1031,In_2085);
or U1474 (N_1474,N_1030,In_727);
nand U1475 (N_1475,In_547,In_788);
or U1476 (N_1476,N_569,In_2414);
or U1477 (N_1477,N_937,In_970);
xor U1478 (N_1478,N_944,N_1144);
or U1479 (N_1479,N_141,N_65);
nand U1480 (N_1480,N_825,In_1837);
xor U1481 (N_1481,In_2543,In_189);
and U1482 (N_1482,In_1516,N_101);
nor U1483 (N_1483,N_306,N_726);
and U1484 (N_1484,In_518,N_893);
or U1485 (N_1485,In_889,N_224);
or U1486 (N_1486,In_1523,In_869);
or U1487 (N_1487,N_349,In_1993);
or U1488 (N_1488,N_1133,In_1169);
nor U1489 (N_1489,N_734,N_509);
nor U1490 (N_1490,In_2398,In_218);
nand U1491 (N_1491,In_872,N_1129);
or U1492 (N_1492,In_2675,N_1100);
and U1493 (N_1493,N_371,N_949);
nor U1494 (N_1494,In_1119,In_2219);
nand U1495 (N_1495,N_591,In_974);
and U1496 (N_1496,In_2024,In_396);
and U1497 (N_1497,N_628,N_668);
nand U1498 (N_1498,N_853,N_1034);
nor U1499 (N_1499,In_1177,N_1036);
nor U1500 (N_1500,N_681,N_786);
xor U1501 (N_1501,In_891,N_693);
xor U1502 (N_1502,N_100,In_1158);
nand U1503 (N_1503,In_1179,In_1293);
nand U1504 (N_1504,N_826,N_445);
nand U1505 (N_1505,In_2820,N_284);
xor U1506 (N_1506,N_702,N_683);
nand U1507 (N_1507,In_2645,In_2998);
nor U1508 (N_1508,N_1002,N_98);
or U1509 (N_1509,N_881,N_749);
xnor U1510 (N_1510,N_896,N_844);
xor U1511 (N_1511,N_1095,N_941);
nor U1512 (N_1512,In_1095,N_1127);
or U1513 (N_1513,N_678,In_2725);
and U1514 (N_1514,In_335,In_649);
xnor U1515 (N_1515,N_1106,In_1649);
and U1516 (N_1516,N_557,In_31);
xnor U1517 (N_1517,N_1176,In_2370);
nor U1518 (N_1518,N_74,In_1652);
xnor U1519 (N_1519,In_2823,In_792);
or U1520 (N_1520,In_2086,N_49);
and U1521 (N_1521,In_1383,In_2117);
and U1522 (N_1522,N_502,In_1451);
and U1523 (N_1523,N_729,N_1060);
xnor U1524 (N_1524,N_695,In_680);
nand U1525 (N_1525,N_940,N_55);
xor U1526 (N_1526,N_126,In_1225);
and U1527 (N_1527,In_1788,N_151);
nor U1528 (N_1528,N_686,In_2031);
nor U1529 (N_1529,N_887,N_851);
or U1530 (N_1530,N_603,N_890);
and U1531 (N_1531,In_1677,In_2574);
nor U1532 (N_1532,In_1200,N_773);
xnor U1533 (N_1533,In_1260,N_497);
nor U1534 (N_1534,In_534,In_2060);
xor U1535 (N_1535,N_769,N_405);
nor U1536 (N_1536,In_877,N_821);
nand U1537 (N_1537,N_487,N_241);
and U1538 (N_1538,In_2515,In_15);
nor U1539 (N_1539,N_411,N_920);
and U1540 (N_1540,N_327,N_883);
and U1541 (N_1541,In_1400,In_1796);
or U1542 (N_1542,In_2399,N_641);
and U1543 (N_1543,In_2170,N_901);
nor U1544 (N_1544,In_1468,N_605);
or U1545 (N_1545,N_1196,In_2049);
nor U1546 (N_1546,N_1118,N_600);
or U1547 (N_1547,N_875,In_1661);
nand U1548 (N_1548,In_2890,In_1585);
and U1549 (N_1549,In_626,N_207);
and U1550 (N_1550,In_1755,In_2699);
or U1551 (N_1551,N_1039,N_610);
nor U1552 (N_1552,In_865,N_972);
xor U1553 (N_1553,In_2730,N_594);
and U1554 (N_1554,N_139,In_643);
nand U1555 (N_1555,N_38,N_710);
and U1556 (N_1556,In_2597,In_1803);
nor U1557 (N_1557,In_1973,N_727);
xor U1558 (N_1558,N_968,N_869);
nor U1559 (N_1559,N_584,In_2679);
or U1560 (N_1560,N_0,In_1630);
nor U1561 (N_1561,In_1307,N_1052);
or U1562 (N_1562,N_820,N_954);
nor U1563 (N_1563,N_114,N_442);
and U1564 (N_1564,N_246,In_433);
or U1565 (N_1565,N_35,N_259);
or U1566 (N_1566,N_1041,N_871);
nand U1567 (N_1567,In_1325,In_2351);
xor U1568 (N_1568,In_2388,In_1885);
nand U1569 (N_1569,In_2437,N_572);
and U1570 (N_1570,N_771,In_242);
nor U1571 (N_1571,In_1893,N_748);
xor U1572 (N_1572,N_913,N_1090);
xor U1573 (N_1573,In_325,In_1873);
nor U1574 (N_1574,In_562,N_1079);
or U1575 (N_1575,N_274,N_1148);
nand U1576 (N_1576,N_630,In_146);
or U1577 (N_1577,N_137,In_628);
xor U1578 (N_1578,N_788,In_2932);
or U1579 (N_1579,In_245,N_1136);
or U1580 (N_1580,In_935,In_2616);
or U1581 (N_1581,N_1157,N_1111);
nor U1582 (N_1582,In_692,In_542);
nor U1583 (N_1583,In_1696,N_328);
and U1584 (N_1584,In_297,In_338);
xnor U1585 (N_1585,N_884,In_2146);
and U1586 (N_1586,N_212,N_956);
nand U1587 (N_1587,In_1874,In_2393);
and U1588 (N_1588,N_789,N_716);
or U1589 (N_1589,N_476,N_181);
xnor U1590 (N_1590,In_2015,In_827);
or U1591 (N_1591,In_1263,N_894);
and U1592 (N_1592,N_723,N_879);
nor U1593 (N_1593,N_1145,N_1037);
or U1594 (N_1594,In_1168,N_78);
xnor U1595 (N_1595,In_893,In_1863);
and U1596 (N_1596,In_1000,In_1971);
or U1597 (N_1597,N_720,N_182);
and U1598 (N_1598,In_1123,In_2867);
nand U1599 (N_1599,In_1099,N_1046);
nor U1600 (N_1600,N_667,N_955);
and U1601 (N_1601,N_1194,In_1363);
xor U1602 (N_1602,In_1560,In_98);
or U1603 (N_1603,N_966,In_1331);
xnor U1604 (N_1604,N_363,N_765);
and U1605 (N_1605,In_1071,In_1089);
xnor U1606 (N_1606,In_2863,In_684);
xnor U1607 (N_1607,N_992,N_675);
xnor U1608 (N_1608,N_390,N_735);
nor U1609 (N_1609,N_1101,In_1758);
nor U1610 (N_1610,In_1638,In_1275);
or U1611 (N_1611,In_163,In_1563);
nor U1612 (N_1612,N_969,N_1006);
nand U1613 (N_1613,In_629,In_601);
or U1614 (N_1614,In_1683,N_408);
xor U1615 (N_1615,In_2793,N_1171);
nor U1616 (N_1616,In_207,N_1114);
and U1617 (N_1617,In_1130,N_362);
and U1618 (N_1618,In_541,In_702);
and U1619 (N_1619,In_2128,N_906);
and U1620 (N_1620,In_156,In_254);
and U1621 (N_1621,In_1345,In_504);
and U1622 (N_1622,In_983,N_1187);
nor U1623 (N_1623,N_696,N_1185);
or U1624 (N_1624,N_687,In_2780);
or U1625 (N_1625,N_376,N_128);
nor U1626 (N_1626,In_1334,N_633);
xnor U1627 (N_1627,N_1122,In_190);
nor U1628 (N_1628,N_1009,In_2708);
nor U1629 (N_1629,N_468,N_532);
nor U1630 (N_1630,In_2575,In_2906);
or U1631 (N_1631,N_1047,N_1116);
or U1632 (N_1632,In_611,In_1012);
and U1633 (N_1633,N_247,N_266);
or U1634 (N_1634,N_334,N_209);
xor U1635 (N_1635,In_2455,In_1166);
nand U1636 (N_1636,In_427,In_555);
or U1637 (N_1637,N_1143,In_805);
xor U1638 (N_1638,N_240,In_280);
nand U1639 (N_1639,N_1045,N_1033);
nor U1640 (N_1640,In_762,In_2045);
xor U1641 (N_1641,N_938,In_2670);
xor U1642 (N_1642,In_905,In_1151);
nor U1643 (N_1643,In_1779,In_660);
nor U1644 (N_1644,In_2702,N_317);
nor U1645 (N_1645,N_680,In_856);
and U1646 (N_1646,N_1093,In_324);
xor U1647 (N_1647,In_1794,N_1121);
nor U1648 (N_1648,N_805,In_2642);
or U1649 (N_1649,N_7,N_448);
nand U1650 (N_1650,N_1019,In_1081);
nor U1651 (N_1651,N_622,N_983);
nand U1652 (N_1652,In_763,In_2214);
and U1653 (N_1653,N_389,In_10);
or U1654 (N_1654,N_832,In_2962);
xnor U1655 (N_1655,In_734,N_450);
or U1656 (N_1656,In_1916,N_849);
nand U1657 (N_1657,N_264,N_673);
nand U1658 (N_1658,N_782,N_766);
nor U1659 (N_1659,N_718,N_868);
nor U1660 (N_1660,N_1049,N_914);
and U1661 (N_1661,In_1644,In_2825);
xnor U1662 (N_1662,In_366,In_444);
and U1663 (N_1663,N_133,In_2905);
and U1664 (N_1664,In_1397,N_285);
and U1665 (N_1665,N_635,In_859);
or U1666 (N_1666,In_412,In_1347);
xnor U1667 (N_1667,In_1342,In_437);
xnor U1668 (N_1668,N_895,In_2315);
xor U1669 (N_1669,In_2317,N_1067);
or U1670 (N_1670,In_109,N_677);
nand U1671 (N_1671,N_838,In_1526);
xor U1672 (N_1672,In_458,In_772);
and U1673 (N_1673,In_1042,N_924);
nor U1674 (N_1674,N_108,In_2058);
nand U1675 (N_1675,In_633,N_1038);
or U1676 (N_1676,In_428,N_830);
nor U1677 (N_1677,N_203,N_709);
nand U1678 (N_1678,N_223,In_2157);
or U1679 (N_1679,In_1512,In_317);
nor U1680 (N_1680,N_192,In_1598);
or U1681 (N_1681,N_1138,In_642);
and U1682 (N_1682,In_2499,N_756);
or U1683 (N_1683,N_170,N_237);
or U1684 (N_1684,In_1554,N_300);
nand U1685 (N_1685,In_2412,In_1034);
and U1686 (N_1686,In_1541,N_839);
nor U1687 (N_1687,N_907,N_850);
nor U1688 (N_1688,N_917,N_794);
and U1689 (N_1689,N_815,In_2919);
or U1690 (N_1690,N_707,In_1157);
and U1691 (N_1691,In_2567,N_801);
nor U1692 (N_1692,In_1210,N_551);
nand U1693 (N_1693,N_23,In_1220);
nand U1694 (N_1694,N_902,In_595);
nor U1695 (N_1695,In_311,N_811);
nor U1696 (N_1696,N_642,In_1066);
nand U1697 (N_1697,N_936,In_2646);
nand U1698 (N_1698,N_899,N_87);
nor U1699 (N_1699,N_195,In_2372);
or U1700 (N_1700,In_2195,In_573);
xor U1701 (N_1701,In_599,In_2764);
and U1702 (N_1702,In_554,In_2295);
or U1703 (N_1703,N_929,N_1001);
nor U1704 (N_1704,In_1373,In_330);
or U1705 (N_1705,N_238,In_2231);
nand U1706 (N_1706,In_2744,In_19);
or U1707 (N_1707,N_1198,In_265);
and U1708 (N_1708,In_45,N_500);
or U1709 (N_1709,N_658,In_423);
and U1710 (N_1710,N_855,In_112);
nand U1711 (N_1711,In_1980,N_276);
nor U1712 (N_1712,In_864,N_867);
and U1713 (N_1713,N_1162,In_116);
or U1714 (N_1714,N_89,In_1507);
nand U1715 (N_1715,N_841,N_785);
and U1716 (N_1716,N_416,In_1864);
nor U1717 (N_1717,N_1155,N_189);
or U1718 (N_1718,In_463,N_1141);
and U1719 (N_1719,N_79,N_440);
xor U1720 (N_1720,N_1193,N_919);
nor U1721 (N_1721,In_1695,In_1530);
xor U1722 (N_1722,N_804,N_1103);
or U1723 (N_1723,In_2466,In_493);
or U1724 (N_1724,In_270,In_589);
and U1725 (N_1725,In_2569,N_492);
nand U1726 (N_1726,In_2417,N_1169);
nor U1727 (N_1727,In_210,N_1066);
nor U1728 (N_1728,N_703,In_981);
nand U1729 (N_1729,N_134,N_1027);
xnor U1730 (N_1730,N_1065,N_245);
nor U1731 (N_1731,N_571,N_122);
or U1732 (N_1732,In_2832,N_994);
nor U1733 (N_1733,In_74,N_1061);
nand U1734 (N_1734,In_84,In_1351);
nor U1735 (N_1735,In_2360,N_453);
xnor U1736 (N_1736,In_1699,N_760);
and U1737 (N_1737,In_241,N_94);
or U1738 (N_1738,In_2608,N_1025);
nand U1739 (N_1739,N_1132,N_1044);
nor U1740 (N_1740,N_953,In_1835);
nor U1741 (N_1741,In_1211,In_127);
nand U1742 (N_1742,In_2163,In_1001);
xnor U1743 (N_1743,N_2,In_288);
xnor U1744 (N_1744,In_2875,In_1495);
and U1745 (N_1745,N_1178,N_823);
and U1746 (N_1746,N_14,In_1768);
or U1747 (N_1747,N_848,N_427);
xnor U1748 (N_1748,N_908,In_890);
nand U1749 (N_1749,N_553,In_984);
and U1750 (N_1750,N_618,N_439);
or U1751 (N_1751,N_1142,N_870);
xnor U1752 (N_1752,N_1005,N_836);
nand U1753 (N_1753,N_706,N_10);
or U1754 (N_1754,N_343,In_2576);
and U1755 (N_1755,N_758,In_1444);
nand U1756 (N_1756,N_691,N_948);
nor U1757 (N_1757,N_273,N_191);
nor U1758 (N_1758,In_1684,N_970);
nand U1759 (N_1759,N_498,N_761);
nand U1760 (N_1760,In_1805,N_1188);
xnor U1761 (N_1761,In_537,In_405);
nor U1762 (N_1762,N_965,In_459);
xnor U1763 (N_1763,N_1086,In_665);
and U1764 (N_1764,In_2709,In_2080);
and U1765 (N_1765,In_2546,In_1102);
and U1766 (N_1766,In_750,N_910);
nor U1767 (N_1767,N_1107,N_614);
xor U1768 (N_1768,N_626,N_864);
or U1769 (N_1769,N_579,In_2990);
or U1770 (N_1770,In_1188,In_2266);
xnor U1771 (N_1771,N_809,N_958);
nor U1772 (N_1772,N_262,In_225);
or U1773 (N_1773,N_1104,N_574);
and U1774 (N_1774,N_27,N_289);
and U1775 (N_1775,N_564,In_1604);
xor U1776 (N_1776,N_604,In_1627);
and U1777 (N_1777,In_1024,In_470);
nor U1778 (N_1778,N_138,In_2358);
xor U1779 (N_1779,In_1414,In_648);
nand U1780 (N_1780,In_2438,N_783);
nor U1781 (N_1781,In_2766,In_52);
and U1782 (N_1782,N_1004,N_750);
nor U1783 (N_1783,In_124,In_1826);
nor U1784 (N_1784,In_2897,N_819);
and U1785 (N_1785,N_61,In_2710);
nand U1786 (N_1786,In_1443,N_86);
or U1787 (N_1787,In_1970,In_489);
xnor U1788 (N_1788,N_1160,In_205);
and U1789 (N_1789,In_2227,N_171);
xor U1790 (N_1790,N_808,N_519);
nand U1791 (N_1791,In_2802,N_1026);
and U1792 (N_1792,In_2534,N_743);
and U1793 (N_1793,In_1759,N_1078);
xnor U1794 (N_1794,In_776,In_2002);
and U1795 (N_1795,In_1858,N_1024);
or U1796 (N_1796,In_1590,In_1202);
and U1797 (N_1797,N_1166,N_700);
nor U1798 (N_1798,In_2816,N_136);
nor U1799 (N_1799,N_632,N_770);
and U1800 (N_1800,N_1422,N_1353);
nand U1801 (N_1801,In_40,N_1229);
or U1802 (N_1802,N_1147,In_1479);
or U1803 (N_1803,N_545,N_1500);
nand U1804 (N_1804,N_15,N_1772);
and U1805 (N_1805,In_291,In_33);
and U1806 (N_1806,N_1569,N_1209);
or U1807 (N_1807,N_1440,N_874);
xnor U1808 (N_1808,In_2135,N_717);
xor U1809 (N_1809,N_1766,In_2027);
xnor U1810 (N_1810,N_1243,N_1715);
and U1811 (N_1811,In_373,In_672);
or U1812 (N_1812,N_1432,N_1408);
and U1813 (N_1813,N_671,N_721);
nand U1814 (N_1814,N_1266,N_739);
or U1815 (N_1815,N_1250,N_1063);
nor U1816 (N_1816,N_46,N_1610);
and U1817 (N_1817,In_1296,N_1281);
nor U1818 (N_1818,N_425,In_2815);
xnor U1819 (N_1819,In_1662,N_1596);
nand U1820 (N_1820,N_1283,N_909);
xnor U1821 (N_1821,N_1625,In_2541);
or U1822 (N_1822,In_168,N_1262);
xor U1823 (N_1823,N_643,In_1406);
xor U1824 (N_1824,N_1427,N_1277);
nor U1825 (N_1825,In_2996,N_1511);
or U1826 (N_1826,N_1270,N_1655);
and U1827 (N_1827,N_1105,N_1497);
or U1828 (N_1828,N_1235,N_581);
nor U1829 (N_1829,N_1520,N_1558);
nor U1830 (N_1830,N_1764,N_1676);
nand U1831 (N_1831,N_1496,In_1367);
xnor U1832 (N_1832,N_1623,N_1628);
or U1833 (N_1833,In_2860,N_1588);
nand U1834 (N_1834,N_1762,In_2871);
nand U1835 (N_1835,N_1627,N_797);
xor U1836 (N_1836,N_1791,N_1321);
nand U1837 (N_1837,N_586,N_856);
nor U1838 (N_1838,N_659,N_1550);
and U1839 (N_1839,N_1507,N_1255);
and U1840 (N_1840,N_1418,N_1438);
nor U1841 (N_1841,In_653,N_1392);
xnor U1842 (N_1842,In_2346,N_1757);
xnor U1843 (N_1843,N_1014,N_1230);
and U1844 (N_1844,N_1481,N_1314);
xor U1845 (N_1845,N_570,N_1259);
or U1846 (N_1846,N_946,In_1515);
nand U1847 (N_1847,N_1672,In_741);
nor U1848 (N_1848,N_1716,N_1374);
nor U1849 (N_1849,N_859,In_1203);
nand U1850 (N_1850,N_1579,N_1202);
and U1851 (N_1851,N_1469,N_978);
nand U1852 (N_1852,N_1362,N_326);
xnor U1853 (N_1853,N_1682,In_2621);
nand U1854 (N_1854,N_1320,N_1748);
xnor U1855 (N_1855,N_1510,N_1493);
and U1856 (N_1856,N_1242,N_916);
or U1857 (N_1857,N_1223,N_1666);
nor U1858 (N_1858,N_1548,N_1697);
or U1859 (N_1859,N_1232,N_1573);
xnor U1860 (N_1860,N_621,N_1566);
nand U1861 (N_1861,N_1248,N_1317);
and U1862 (N_1862,N_927,N_1450);
nand U1863 (N_1863,In_387,N_552);
xnor U1864 (N_1864,In_690,N_1441);
xnor U1865 (N_1865,In_2206,N_1717);
xnor U1866 (N_1866,N_1375,In_1106);
nor U1867 (N_1867,N_1613,In_1780);
xor U1868 (N_1868,N_1562,N_1670);
xor U1869 (N_1869,N_742,N_1268);
xor U1870 (N_1870,In_2685,N_933);
or U1871 (N_1871,N_1779,N_1200);
nand U1872 (N_1872,N_957,N_728);
nand U1873 (N_1873,N_135,N_1788);
xnor U1874 (N_1874,N_1656,N_900);
nor U1875 (N_1875,N_905,In_1372);
or U1876 (N_1876,N_550,N_1190);
or U1877 (N_1877,N_1352,In_2854);
and U1878 (N_1878,In_385,N_1201);
and U1879 (N_1879,N_1368,In_2246);
nand U1880 (N_1880,N_1172,In_2154);
nand U1881 (N_1881,N_1334,N_1630);
xor U1882 (N_1882,N_1117,In_1348);
nor U1883 (N_1883,N_1294,N_401);
or U1884 (N_1884,N_1506,N_1743);
nand U1885 (N_1885,N_1291,In_2794);
and U1886 (N_1886,N_1179,N_1279);
xor U1887 (N_1887,In_1429,N_495);
nand U1888 (N_1888,N_1085,N_947);
nand U1889 (N_1889,N_1518,N_190);
nor U1890 (N_1890,N_699,N_1598);
or U1891 (N_1891,N_1293,N_1411);
nand U1892 (N_1892,N_1754,N_1642);
nand U1893 (N_1893,N_1222,N_1649);
or U1894 (N_1894,N_1712,N_1457);
and U1895 (N_1895,N_1312,N_1322);
and U1896 (N_1896,N_982,N_127);
xor U1897 (N_1897,N_1434,N_1533);
nor U1898 (N_1898,N_1280,In_2653);
nand U1899 (N_1899,N_1015,N_1614);
or U1900 (N_1900,N_1554,N_1648);
and U1901 (N_1901,N_1373,N_1478);
nand U1902 (N_1902,N_1704,N_733);
nand U1903 (N_1903,In_1061,In_2274);
and U1904 (N_1904,In_667,N_1378);
and U1905 (N_1905,N_612,N_1351);
xnor U1906 (N_1906,N_163,N_1247);
xnor U1907 (N_1907,N_1040,In_1986);
nor U1908 (N_1908,N_1297,N_1761);
nand U1909 (N_1909,N_1152,In_1209);
and U1910 (N_1910,N_1401,N_1601);
or U1911 (N_1911,In_597,N_316);
nand U1912 (N_1912,N_1335,N_1689);
xnor U1913 (N_1913,In_737,N_1398);
nand U1914 (N_1914,N_477,In_2165);
xor U1915 (N_1915,N_1674,N_1724);
or U1916 (N_1916,N_265,N_1546);
and U1917 (N_1917,N_1403,In_575);
nand U1918 (N_1918,N_1028,N_1424);
nand U1919 (N_1919,N_648,In_1091);
or U1920 (N_1920,In_2110,N_1382);
nand U1921 (N_1921,N_1264,In_1252);
nand U1922 (N_1922,N_639,In_1197);
or U1923 (N_1923,N_315,N_1357);
xor U1924 (N_1924,N_1622,N_1703);
or U1925 (N_1925,In_677,In_153);
nor U1926 (N_1926,N_1696,N_368);
and U1927 (N_1927,In_2069,N_1739);
or U1928 (N_1928,N_674,In_1809);
or U1929 (N_1929,N_1453,N_985);
xor U1930 (N_1930,In_2817,N_1661);
xor U1931 (N_1931,N_1760,N_1563);
nor U1932 (N_1932,In_2261,N_1216);
nor U1933 (N_1933,In_1527,N_1796);
nor U1934 (N_1934,N_1698,N_1340);
and U1935 (N_1935,N_1786,N_299);
nand U1936 (N_1936,N_1356,N_1719);
xnor U1937 (N_1937,N_1449,N_1713);
nor U1938 (N_1938,N_1700,N_1685);
xor U1939 (N_1939,N_1140,N_1084);
xor U1940 (N_1940,N_1011,In_2795);
nor U1941 (N_1941,N_64,In_465);
and U1942 (N_1942,In_2468,In_2655);
or U1943 (N_1943,N_800,N_1773);
nand U1944 (N_1944,In_2945,In_2857);
nand U1945 (N_1945,In_2139,N_1285);
and U1946 (N_1946,N_1480,N_1591);
or U1947 (N_1947,N_565,N_840);
or U1948 (N_1948,In_170,In_1833);
xor U1949 (N_1949,In_2602,N_1501);
or U1950 (N_1950,N_1276,N_1163);
nor U1951 (N_1951,N_1448,N_1551);
or U1952 (N_1952,N_897,N_243);
nand U1953 (N_1953,In_1405,N_1663);
and U1954 (N_1954,N_1436,In_103);
nor U1955 (N_1955,In_744,N_1691);
and U1956 (N_1956,In_1114,In_482);
or U1957 (N_1957,In_840,N_1758);
nor U1958 (N_1958,N_1344,N_1459);
and U1959 (N_1959,N_533,N_660);
xnor U1960 (N_1960,N_692,N_876);
and U1961 (N_1961,In_726,N_1617);
or U1962 (N_1962,N_1417,N_1515);
or U1963 (N_1963,N_1746,N_1616);
or U1964 (N_1964,N_1765,N_1301);
nor U1965 (N_1965,N_842,N_1770);
or U1966 (N_1966,N_1729,N_1337);
or U1967 (N_1967,N_1722,In_2369);
nand U1968 (N_1968,N_943,In_35);
or U1969 (N_1969,In_1279,N_1184);
or U1970 (N_1970,N_1585,In_664);
or U1971 (N_1971,In_1727,N_1463);
nand U1972 (N_1972,N_1701,N_1323);
and U1973 (N_1973,N_1304,In_2533);
nand U1974 (N_1974,N_730,N_1633);
nand U1975 (N_1975,In_2701,N_1239);
or U1976 (N_1976,N_1112,N_1205);
xnor U1977 (N_1977,N_1365,In_300);
and U1978 (N_1978,N_980,N_1652);
xnor U1979 (N_1979,N_704,N_828);
nor U1980 (N_1980,In_2197,N_1219);
nor U1981 (N_1981,N_1538,N_781);
xnor U1982 (N_1982,N_670,N_1272);
nand U1983 (N_1983,N_1664,N_989);
xnor U1984 (N_1984,N_1678,N_1191);
nand U1985 (N_1985,N_615,N_974);
nor U1986 (N_1986,N_1389,N_1502);
nand U1987 (N_1987,In_1402,N_1379);
and U1988 (N_1988,N_1699,In_1828);
or U1989 (N_1989,In_900,N_1745);
xnor U1990 (N_1990,N_1733,N_573);
xor U1991 (N_1991,N_1557,In_2047);
nor U1992 (N_1992,N_1723,N_412);
xnor U1993 (N_1993,N_1134,N_1213);
or U1994 (N_1994,In_2126,N_1567);
xnor U1995 (N_1995,N_1595,N_1319);
xnor U1996 (N_1996,In_748,N_1256);
and U1997 (N_1997,In_1586,N_1433);
or U1998 (N_1998,In_431,N_1215);
or U1999 (N_1999,N_1425,In_1634);
nand U2000 (N_2000,N_1534,In_2478);
nor U2001 (N_2001,N_1634,N_1308);
xor U2002 (N_2002,In_2142,In_769);
xor U2003 (N_2003,N_1032,N_391);
or U2004 (N_2004,N_1780,N_1261);
nor U2005 (N_2005,N_1612,N_1288);
and U2006 (N_2006,In_1777,In_1176);
nand U2007 (N_2007,N_945,N_1059);
or U2008 (N_2008,In_947,N_715);
xor U2009 (N_2009,N_1620,N_1525);
nand U2010 (N_2010,N_1549,N_1088);
and U2011 (N_2011,N_1186,In_2876);
and U2012 (N_2012,N_1751,In_2592);
xor U2013 (N_2013,In_2845,N_1727);
nor U2014 (N_2014,In_1482,N_556);
nand U2015 (N_2015,N_1350,N_1647);
xnor U2016 (N_2016,N_1168,N_1445);
and U2017 (N_2017,In_2544,N_1435);
nor U2018 (N_2018,In_2020,In_2830);
nor U2019 (N_2019,In_1538,In_162);
and U2020 (N_2020,N_493,N_1396);
or U2021 (N_2021,N_1564,N_1442);
xnor U2022 (N_2022,In_2017,N_1736);
and U2023 (N_2023,N_1367,N_1680);
and U2024 (N_2024,N_1460,N_1204);
nor U2025 (N_2025,N_763,N_1306);
and U2026 (N_2026,N_1517,N_1000);
nor U2027 (N_2027,N_1487,N_1290);
nand U2028 (N_2028,In_194,N_1690);
nor U2029 (N_2029,N_1677,N_294);
or U2030 (N_2030,N_176,N_787);
or U2031 (N_2031,N_650,In_17);
and U2032 (N_2032,N_1076,N_629);
and U2033 (N_2033,N_1547,N_1212);
nor U2034 (N_2034,N_1657,N_1671);
nor U2035 (N_2035,N_1473,N_975);
and U2036 (N_2036,N_1313,N_275);
nand U2037 (N_2037,N_1606,In_1392);
nand U2038 (N_2038,N_1466,N_1694);
xnor U2039 (N_2039,In_1712,N_752);
nand U2040 (N_2040,N_1300,N_204);
and U2041 (N_2041,N_1519,In_837);
nor U2042 (N_2042,N_1474,N_5);
nand U2043 (N_2043,N_653,In_955);
and U2044 (N_2044,N_611,N_685);
nor U2045 (N_2045,In_1277,In_62);
and U2046 (N_2046,N_1669,N_1561);
nor U2047 (N_2047,N_172,N_1597);
or U2048 (N_2048,N_1477,N_1094);
xor U2049 (N_2049,N_1265,N_1447);
and U2050 (N_2050,In_1531,N_1149);
xor U2051 (N_2051,In_2044,N_1646);
nand U2052 (N_2052,In_1408,In_1467);
or U2053 (N_2053,In_2964,N_999);
and U2054 (N_2054,N_1708,N_1681);
and U2055 (N_2055,N_1465,N_1753);
nand U2056 (N_2056,N_1071,N_1240);
and U2057 (N_2057,N_379,N_1385);
and U2058 (N_2058,In_477,N_1570);
xnor U2059 (N_2059,N_1675,N_1249);
xnor U2060 (N_2060,In_403,N_1624);
nor U2061 (N_2061,N_26,N_724);
or U2062 (N_2062,N_915,In_1918);
or U2063 (N_2063,N_1638,N_1728);
nor U2064 (N_2064,In_2758,In_2239);
or U2065 (N_2065,N_1298,N_1369);
and U2066 (N_2066,N_1741,N_1537);
xor U2067 (N_2067,N_764,In_2199);
and U2068 (N_2068,N_1404,N_1439);
xnor U2069 (N_2069,N_1325,In_1417);
nand U2070 (N_2070,In_2485,In_108);
or U2071 (N_2071,N_1516,In_2999);
or U2072 (N_2072,N_1575,In_1866);
or U2073 (N_2073,In_1126,N_1130);
and U2074 (N_2074,N_12,N_1225);
nand U2075 (N_2075,N_1512,N_1257);
xor U2076 (N_2076,In_1535,N_1730);
xor U2077 (N_2077,N_963,N_1175);
and U2078 (N_2078,N_1437,In_818);
xor U2079 (N_2079,N_1446,N_1490);
nor U2080 (N_2080,N_1241,N_1640);
nor U2081 (N_2081,In_2038,In_39);
nor U2082 (N_2082,N_1364,In_671);
xor U2083 (N_2083,In_1241,In_1298);
xnor U2084 (N_2084,N_1555,N_1621);
xor U2085 (N_2085,N_1383,In_2004);
xnor U2086 (N_2086,N_912,N_1329);
nand U2087 (N_2087,In_1036,In_1742);
xor U2088 (N_2088,N_1768,In_1715);
nor U2089 (N_2089,N_57,N_1315);
xor U2090 (N_2090,N_1233,In_439);
or U2091 (N_2091,N_1609,N_1577);
xor U2092 (N_2092,N_1635,N_1399);
xnor U2093 (N_2093,N_817,In_1218);
or U2094 (N_2094,N_1452,N_1732);
xor U2095 (N_2095,In_1886,N_409);
and U2096 (N_2096,In_2059,N_1208);
and U2097 (N_2097,N_1769,N_1426);
or U2098 (N_2098,N_1735,N_1413);
nor U2099 (N_2099,N_1284,N_1390);
nand U2100 (N_2100,N_1571,N_1543);
xnor U2101 (N_2101,In_2779,N_1289);
and U2102 (N_2102,N_1102,N_1282);
xnor U2103 (N_2103,N_1665,N_1443);
nor U2104 (N_2104,N_1429,N_1393);
and U2105 (N_2105,N_1668,N_1513);
nor U2106 (N_2106,N_1785,In_295);
nor U2107 (N_2107,In_133,N_793);
or U2108 (N_2108,In_2564,In_2480);
or U2109 (N_2109,N_922,N_802);
nand U2110 (N_2110,N_1494,N_1013);
xnor U2111 (N_2111,N_1324,N_1330);
and U2112 (N_2112,N_806,N_1333);
xor U2113 (N_2113,N_1343,N_1528);
xnor U2114 (N_2114,N_1618,In_683);
nor U2115 (N_2115,N_1400,N_1684);
nor U2116 (N_2116,N_1530,N_113);
xnor U2117 (N_2117,N_1484,N_1428);
nand U2118 (N_2118,In_1726,In_937);
nor U2119 (N_2119,In_1462,N_1087);
and U2120 (N_2120,N_1096,In_1723);
and U2121 (N_2121,In_1388,N_1252);
and U2122 (N_2122,N_689,N_1331);
and U2123 (N_2123,N_1167,N_1394);
or U2124 (N_2124,N_1207,N_1720);
nand U2125 (N_2125,N_1295,N_1583);
xnor U2126 (N_2126,N_1755,In_1656);
nand U2127 (N_2127,N_1718,N_1415);
nor U2128 (N_2128,In_1205,N_1328);
and U2129 (N_2129,In_82,N_1767);
xnor U2130 (N_2130,N_1376,In_2410);
xor U2131 (N_2131,In_231,N_613);
or U2132 (N_2132,N_1539,N_1514);
and U2133 (N_2133,N_1472,In_2760);
and U2134 (N_2134,N_1018,N_1058);
nand U2135 (N_2135,N_1794,N_778);
and U2136 (N_2136,N_394,N_1482);
xor U2137 (N_2137,N_1594,In_2474);
and U2138 (N_2138,N_762,N_1318);
or U2139 (N_2139,N_903,N_1645);
or U2140 (N_2140,N_857,In_1653);
xor U2141 (N_2141,N_1522,N_547);
nand U2142 (N_2142,N_973,In_193);
and U2143 (N_2143,N_1274,N_1341);
nand U2144 (N_2144,N_1725,In_2969);
nor U2145 (N_2145,In_579,In_2098);
nand U2146 (N_2146,N_332,N_1253);
and U2147 (N_2147,N_1744,N_1414);
xnor U2148 (N_2148,N_90,In_721);
nand U2149 (N_2149,N_1629,N_1458);
nor U2150 (N_2150,N_1775,In_125);
and U2151 (N_2151,N_1384,N_1781);
and U2152 (N_2152,N_1673,In_1485);
xor U2153 (N_2153,N_539,In_2068);
nand U2154 (N_2154,N_1412,N_1784);
xor U2155 (N_2155,N_1574,In_2891);
nand U2156 (N_2156,N_178,N_1740);
nor U2157 (N_2157,In_1912,N_1799);
xnor U2158 (N_2158,In_2459,N_1456);
and U2159 (N_2159,N_625,N_1486);
nor U2160 (N_2160,N_1119,N_1542);
nand U2161 (N_2161,N_1016,N_1683);
and U2162 (N_2162,In_2181,In_2178);
nand U2163 (N_2163,In_976,In_2840);
or U2164 (N_2164,N_292,N_331);
nor U2165 (N_2165,N_1731,N_131);
nor U2166 (N_2166,In_2290,N_562);
xor U2167 (N_2167,In_2716,N_1654);
nor U2168 (N_2168,N_1346,In_693);
xor U2169 (N_2169,In_2313,N_1192);
or U2170 (N_2170,N_1783,N_1763);
nor U2171 (N_2171,In_2536,N_1224);
or U2172 (N_2172,In_1905,N_1578);
xnor U2173 (N_2173,N_1545,N_1246);
nor U2174 (N_2174,N_1777,In_793);
xnor U2175 (N_2175,N_1658,N_1342);
and U2176 (N_2176,In_1725,In_2707);
nor U2177 (N_2177,N_1544,N_1468);
or U2178 (N_2178,In_123,N_485);
and U2179 (N_2179,N_311,In_1693);
nor U2180 (N_2180,In_2193,N_1388);
xnor U2181 (N_2181,N_1707,N_1123);
and U2182 (N_2182,N_669,N_1750);
and U2183 (N_2183,In_1648,N_1386);
nand U2184 (N_2184,N_1581,N_1527);
or U2185 (N_2185,N_738,In_560);
or U2186 (N_2186,In_2633,In_594);
nor U2187 (N_2187,N_1406,N_1366);
nand U2188 (N_2188,In_1421,In_2775);
nand U2189 (N_2189,N_1234,N_636);
nor U2190 (N_2190,N_714,N_1387);
or U2191 (N_2191,N_776,N_1377);
nor U2192 (N_2192,N_130,N_798);
and U2193 (N_2193,N_1228,N_1790);
nor U2194 (N_2194,N_1327,N_1286);
and U2195 (N_2195,N_595,N_1206);
and U2196 (N_2196,In_675,N_996);
nand U2197 (N_2197,N_1795,In_2527);
nand U2198 (N_2198,N_1636,In_2677);
or U2199 (N_2199,N_1361,N_1559);
xnor U2200 (N_2200,N_688,N_654);
or U2201 (N_2201,N_1568,In_4);
xnor U2202 (N_2202,N_1455,N_977);
xor U2203 (N_2203,N_951,In_2991);
or U2204 (N_2204,In_563,N_1605);
xor U2205 (N_2205,In_1962,N_1409);
xnor U2206 (N_2206,N_1582,N_1643);
xor U2207 (N_2207,In_2160,N_1339);
or U2208 (N_2208,N_1632,N_1607);
nand U2209 (N_2209,In_1981,In_429);
or U2210 (N_2210,In_2934,N_1789);
nand U2211 (N_2211,N_1221,N_1380);
and U2212 (N_2212,N_1326,N_1391);
or U2213 (N_2213,N_1503,N_1359);
and U2214 (N_2214,N_1505,N_505);
or U2215 (N_2215,In_1651,N_1589);
and U2216 (N_2216,In_1154,N_103);
and U2217 (N_2217,N_1263,N_1430);
nand U2218 (N_2218,N_1650,N_1419);
and U2219 (N_2219,N_649,N_1584);
nor U2220 (N_2220,N_1332,N_1358);
or U2221 (N_2221,N_1476,N_1310);
nor U2222 (N_2222,N_1316,N_1003);
nand U2223 (N_2223,N_1572,In_1416);
nand U2224 (N_2224,In_591,N_1749);
nor U2225 (N_2225,In_1587,N_1742);
or U2226 (N_2226,N_1738,In_1571);
and U2227 (N_2227,N_1451,In_654);
nand U2228 (N_2228,In_1382,N_1641);
xor U2229 (N_2229,N_1488,In_29);
nor U2230 (N_2230,N_1726,N_186);
nand U2231 (N_2231,N_1659,N_1737);
and U2232 (N_2232,N_873,N_813);
or U2233 (N_2233,N_1787,In_1458);
nor U2234 (N_2234,N_1611,N_1363);
nor U2235 (N_2235,N_1771,In_1073);
and U2236 (N_2236,N_1471,N_1354);
nor U2237 (N_2237,In_113,N_1260);
or U2238 (N_2238,N_1693,N_124);
nor U2239 (N_2239,In_609,In_1356);
and U2240 (N_2240,N_1602,N_712);
nand U2241 (N_2241,N_1461,In_1226);
nand U2242 (N_2242,In_2726,N_1532);
and U2243 (N_2243,N_1348,N_1798);
and U2244 (N_2244,N_1153,In_83);
nand U2245 (N_2245,N_1508,In_1917);
nand U2246 (N_2246,In_898,N_1560);
and U2247 (N_2247,In_2902,N_1637);
xor U2248 (N_2248,N_1553,N_1402);
and U2249 (N_2249,N_722,N_1540);
or U2250 (N_2250,In_2454,N_471);
nand U2251 (N_2251,N_1305,N_926);
or U2252 (N_2252,N_1372,In_2148);
nand U2253 (N_2253,In_1108,N_1495);
nor U2254 (N_2254,In_2075,N_1062);
nand U2255 (N_2255,N_1347,In_2972);
nor U2256 (N_2256,N_1687,In_914);
nand U2257 (N_2257,N_470,N_1211);
nand U2258 (N_2258,N_148,N_1667);
and U2259 (N_2259,N_1576,N_657);
or U2260 (N_2260,N_1483,N_1395);
nor U2261 (N_2261,N_546,In_2513);
nor U2262 (N_2262,In_695,In_1845);
nand U2263 (N_2263,N_661,N_360);
and U2264 (N_2264,In_1248,N_1504);
xnor U2265 (N_2265,N_385,In_2105);
nand U2266 (N_2266,N_676,N_1267);
or U2267 (N_2267,N_1709,N_1360);
xor U2268 (N_2268,In_2755,N_309);
or U2269 (N_2269,In_1974,In_2132);
nand U2270 (N_2270,N_1776,N_1338);
or U2271 (N_2271,In_1977,N_1336);
nand U2272 (N_2272,N_1370,N_1711);
or U2273 (N_2273,N_1734,N_1586);
and U2274 (N_2274,N_1580,N_1254);
xnor U2275 (N_2275,N_1273,N_1010);
nor U2276 (N_2276,In_606,In_2046);
or U2277 (N_2277,N_413,N_260);
nor U2278 (N_2278,N_602,N_1644);
xor U2279 (N_2279,N_165,N_1258);
nor U2280 (N_2280,N_1302,N_1631);
and U2281 (N_2281,In_2884,In_2939);
and U2282 (N_2282,In_227,In_2308);
and U2283 (N_2283,In_1395,N_1778);
or U2284 (N_2284,N_619,N_1214);
xnor U2285 (N_2285,In_1614,N_34);
nand U2286 (N_2286,N_1421,In_407);
and U2287 (N_2287,In_2516,N_1692);
nand U2288 (N_2288,In_1982,N_1509);
nor U2289 (N_2289,In_2111,N_1307);
xor U2290 (N_2290,N_1782,In_136);
nand U2291 (N_2291,In_1948,N_1407);
xnor U2292 (N_2292,N_196,In_1643);
and U2293 (N_2293,N_1756,N_1381);
nor U2294 (N_2294,N_1705,N_1593);
nand U2295 (N_2295,In_686,In_1539);
or U2296 (N_2296,N_1639,N_1679);
nand U2297 (N_2297,N_1714,N_517);
nor U2298 (N_2298,In_1877,In_1529);
xnor U2299 (N_2299,N_1195,In_2149);
nor U2300 (N_2300,N_1599,N_1238);
nor U2301 (N_2301,N_1070,N_1454);
and U2302 (N_2302,N_1489,N_1420);
nand U2303 (N_2303,N_1125,N_563);
or U2304 (N_2304,In_2427,N_1565);
nand U2305 (N_2305,In_166,N_1397);
or U2306 (N_2306,In_2,N_1182);
nor U2307 (N_2307,N_1479,N_663);
nor U2308 (N_2308,N_1526,N_1462);
nand U2309 (N_2309,In_2071,N_1292);
nor U2310 (N_2310,N_1226,N_272);
nand U2311 (N_2311,In_2903,In_1215);
nand U2312 (N_2312,N_1470,N_925);
or U2313 (N_2313,In_1117,N_1197);
and U2314 (N_2314,N_1524,N_1371);
nand U2315 (N_2315,N_1410,N_1416);
xnor U2316 (N_2316,N_846,N_719);
and U2317 (N_2317,In_2976,N_1181);
nor U2318 (N_2318,N_1793,N_1797);
nand U2319 (N_2319,N_1108,N_1220);
or U2320 (N_2320,In_2805,N_1556);
xnor U2321 (N_2321,N_1083,N_904);
or U2322 (N_2322,In_1270,N_1296);
nor U2323 (N_2323,N_1491,In_1006);
and U2324 (N_2324,N_623,In_480);
nand U2325 (N_2325,N_1752,N_1227);
nor U2326 (N_2326,N_441,In_1774);
and U2327 (N_2327,N_606,In_1294);
nand U2328 (N_2328,N_827,N_1615);
and U2329 (N_2329,N_990,N_1604);
or U2330 (N_2330,N_1151,In_1976);
xor U2331 (N_2331,N_1702,In_1926);
xnor U2332 (N_2332,N_288,N_149);
or U2333 (N_2333,N_484,N_1552);
nor U2334 (N_2334,N_967,N_1587);
and U2335 (N_2335,N_664,N_1217);
xor U2336 (N_2336,N_1349,N_380);
or U2337 (N_2337,In_610,In_352);
or U2338 (N_2338,N_1405,N_1695);
xor U2339 (N_2339,N_1237,N_1278);
nor U2340 (N_2340,N_270,In_1681);
xor U2341 (N_2341,In_546,N_1688);
nand U2342 (N_2342,N_1231,N_1203);
and U2343 (N_2343,N_1747,N_818);
and U2344 (N_2344,In_2673,In_2918);
nor U2345 (N_2345,N_831,In_2220);
or U2346 (N_2346,N_1464,In_65);
nand U2347 (N_2347,N_1721,N_1536);
nand U2348 (N_2348,N_297,N_737);
and U2349 (N_2349,N_1619,In_2761);
and U2350 (N_2350,N_459,In_1283);
xnor U2351 (N_2351,N_1355,N_1774);
or U2352 (N_2352,In_287,N_1467);
and U2353 (N_2353,N_1600,In_1865);
xnor U2354 (N_2354,In_1934,N_698);
or U2355 (N_2355,N_878,N_107);
nand U2356 (N_2356,N_1303,N_1251);
nand U2357 (N_2357,In_2428,N_339);
and U2358 (N_2358,N_1686,In_1051);
nand U2359 (N_2359,N_1521,N_1608);
or U2360 (N_2360,N_1535,N_1042);
or U2361 (N_2361,N_1236,In_2216);
xor U2362 (N_2362,N_997,N_1299);
xnor U2363 (N_2363,N_1759,In_1659);
xnor U2364 (N_2364,N_1431,N_863);
xor U2365 (N_2365,In_1821,N_1269);
xnor U2366 (N_2366,In_264,N_336);
nand U2367 (N_2367,N_1592,N_1523);
nor U2368 (N_2368,N_645,N_1022);
or U2369 (N_2369,N_1710,In_2839);
and U2370 (N_2370,N_1275,N_1531);
nor U2371 (N_2371,In_1353,N_1271);
or U2372 (N_2372,N_1541,N_1485);
nor U2373 (N_2373,N_144,In_1510);
xnor U2374 (N_2374,N_995,In_1751);
or U2375 (N_2375,N_1660,In_880);
or U2376 (N_2376,In_1266,N_1492);
nor U2377 (N_2377,N_1590,N_1287);
or U2378 (N_2378,N_930,N_1498);
and U2379 (N_2379,N_589,N_1183);
nor U2380 (N_2380,N_886,N_1423);
nor U2381 (N_2381,N_1499,N_1706);
nand U2382 (N_2382,In_2247,N_515);
and U2383 (N_2383,N_1311,In_1884);
nor U2384 (N_2384,N_1651,In_1647);
xnor U2385 (N_2385,In_2883,In_781);
xor U2386 (N_2386,In_1274,In_1655);
or U2387 (N_2387,In_2465,N_1345);
nor U2388 (N_2388,In_1011,In_1136);
nor U2389 (N_2389,N_81,N_1244);
nor U2390 (N_2390,In_44,N_1603);
xnor U2391 (N_2391,N_790,N_1309);
xor U2392 (N_2392,In_2864,N_1792);
and U2393 (N_2393,N_1218,N_1210);
xnor U2394 (N_2394,In_764,In_326);
xor U2395 (N_2395,N_1662,N_1444);
and U2396 (N_2396,In_1192,N_1626);
nor U2397 (N_2397,N_1245,In_1432);
nand U2398 (N_2398,N_1475,In_1058);
xnor U2399 (N_2399,N_1529,N_1653);
or U2400 (N_2400,N_1886,N_2347);
nor U2401 (N_2401,N_1806,N_2219);
nor U2402 (N_2402,N_2089,N_1949);
nor U2403 (N_2403,N_1891,N_2227);
xnor U2404 (N_2404,N_1866,N_2314);
xor U2405 (N_2405,N_2349,N_1901);
or U2406 (N_2406,N_2031,N_2167);
and U2407 (N_2407,N_2305,N_2085);
nand U2408 (N_2408,N_2171,N_2238);
and U2409 (N_2409,N_2166,N_1957);
and U2410 (N_2410,N_2078,N_1955);
nor U2411 (N_2411,N_2175,N_1870);
nor U2412 (N_2412,N_1965,N_2060);
xor U2413 (N_2413,N_2099,N_2006);
nand U2414 (N_2414,N_1859,N_2327);
nand U2415 (N_2415,N_1970,N_2054);
xor U2416 (N_2416,N_2244,N_1926);
nor U2417 (N_2417,N_2266,N_1823);
xnor U2418 (N_2418,N_2370,N_2053);
nand U2419 (N_2419,N_2066,N_1919);
and U2420 (N_2420,N_2178,N_1927);
nand U2421 (N_2421,N_1971,N_1967);
or U2422 (N_2422,N_1836,N_2399);
nor U2423 (N_2423,N_2058,N_1974);
xor U2424 (N_2424,N_2240,N_2016);
nor U2425 (N_2425,N_2333,N_1807);
xnor U2426 (N_2426,N_2222,N_2135);
nor U2427 (N_2427,N_1944,N_1879);
nand U2428 (N_2428,N_2228,N_1811);
xnor U2429 (N_2429,N_2036,N_2143);
nor U2430 (N_2430,N_2208,N_2179);
xnor U2431 (N_2431,N_2043,N_2077);
and U2432 (N_2432,N_2380,N_2141);
nand U2433 (N_2433,N_1890,N_1841);
xnor U2434 (N_2434,N_2273,N_2181);
nand U2435 (N_2435,N_2311,N_1882);
and U2436 (N_2436,N_2204,N_2180);
and U2437 (N_2437,N_2133,N_1952);
nand U2438 (N_2438,N_2284,N_2246);
and U2439 (N_2439,N_2280,N_1931);
and U2440 (N_2440,N_2234,N_2027);
and U2441 (N_2441,N_2325,N_2291);
xor U2442 (N_2442,N_1903,N_1816);
or U2443 (N_2443,N_2151,N_2172);
nor U2444 (N_2444,N_2187,N_1883);
nand U2445 (N_2445,N_2110,N_2081);
nor U2446 (N_2446,N_2383,N_2257);
xnor U2447 (N_2447,N_2264,N_2070);
nor U2448 (N_2448,N_2087,N_2005);
or U2449 (N_2449,N_2012,N_2357);
and U2450 (N_2450,N_2283,N_2150);
or U2451 (N_2451,N_1856,N_2119);
xor U2452 (N_2452,N_1972,N_2355);
and U2453 (N_2453,N_1851,N_2049);
xnor U2454 (N_2454,N_2338,N_2158);
or U2455 (N_2455,N_1973,N_2365);
or U2456 (N_2456,N_2366,N_2023);
nand U2457 (N_2457,N_1802,N_2071);
nor U2458 (N_2458,N_2067,N_2321);
or U2459 (N_2459,N_1954,N_2374);
or U2460 (N_2460,N_2393,N_1956);
and U2461 (N_2461,N_2214,N_1887);
nand U2462 (N_2462,N_2117,N_1850);
and U2463 (N_2463,N_1847,N_2348);
nor U2464 (N_2464,N_2358,N_2195);
nand U2465 (N_2465,N_1942,N_1939);
nor U2466 (N_2466,N_1910,N_2249);
or U2467 (N_2467,N_2254,N_2293);
or U2468 (N_2468,N_2168,N_1962);
xor U2469 (N_2469,N_2197,N_2267);
xnor U2470 (N_2470,N_1943,N_1818);
nor U2471 (N_2471,N_1913,N_2209);
xnor U2472 (N_2472,N_2044,N_2350);
nor U2473 (N_2473,N_2001,N_2161);
nand U2474 (N_2474,N_2372,N_2094);
or U2475 (N_2475,N_2302,N_2050);
and U2476 (N_2476,N_1855,N_1832);
xor U2477 (N_2477,N_2326,N_2176);
xnor U2478 (N_2478,N_1878,N_2310);
and U2479 (N_2479,N_1905,N_2295);
xnor U2480 (N_2480,N_2020,N_2155);
nand U2481 (N_2481,N_2108,N_1953);
xnor U2482 (N_2482,N_2220,N_1978);
or U2483 (N_2483,N_1898,N_2074);
xor U2484 (N_2484,N_2217,N_1868);
or U2485 (N_2485,N_2265,N_2035);
or U2486 (N_2486,N_2042,N_1852);
nor U2487 (N_2487,N_1840,N_2385);
nand U2488 (N_2488,N_1940,N_2223);
nor U2489 (N_2489,N_1895,N_2026);
nand U2490 (N_2490,N_2292,N_2361);
xnor U2491 (N_2491,N_2306,N_2336);
nor U2492 (N_2492,N_2037,N_2025);
nor U2493 (N_2493,N_1936,N_2390);
xor U2494 (N_2494,N_1843,N_2126);
or U2495 (N_2495,N_2289,N_2274);
nor U2496 (N_2496,N_2237,N_1950);
or U2497 (N_2497,N_2317,N_2194);
xnor U2498 (N_2498,N_1961,N_2236);
or U2499 (N_2499,N_1897,N_2101);
xnor U2500 (N_2500,N_2344,N_1842);
xor U2501 (N_2501,N_1872,N_1871);
and U2502 (N_2502,N_2202,N_1863);
xor U2503 (N_2503,N_2341,N_1924);
and U2504 (N_2504,N_1922,N_2029);
and U2505 (N_2505,N_2095,N_2352);
or U2506 (N_2506,N_1803,N_2201);
or U2507 (N_2507,N_2062,N_2343);
or U2508 (N_2508,N_2318,N_1857);
nand U2509 (N_2509,N_2083,N_1932);
nand U2510 (N_2510,N_2258,N_1917);
xnor U2511 (N_2511,N_2192,N_1839);
nand U2512 (N_2512,N_2225,N_1935);
and U2513 (N_2513,N_1948,N_2169);
and U2514 (N_2514,N_1844,N_2122);
nor U2515 (N_2515,N_1838,N_2387);
or U2516 (N_2516,N_2146,N_2107);
xor U2517 (N_2517,N_1986,N_1964);
nand U2518 (N_2518,N_1980,N_1861);
and U2519 (N_2519,N_2144,N_1997);
and U2520 (N_2520,N_2251,N_2268);
xnor U2521 (N_2521,N_1914,N_1815);
and U2522 (N_2522,N_2055,N_1831);
nor U2523 (N_2523,N_2324,N_2301);
nor U2524 (N_2524,N_2021,N_2015);
and U2525 (N_2525,N_2369,N_1881);
nor U2526 (N_2526,N_1826,N_2032);
nand U2527 (N_2527,N_2396,N_2235);
or U2528 (N_2528,N_1984,N_1849);
and U2529 (N_2529,N_2038,N_2079);
or U2530 (N_2530,N_2379,N_1918);
nand U2531 (N_2531,N_2183,N_1893);
nor U2532 (N_2532,N_2243,N_2353);
nand U2533 (N_2533,N_2395,N_2286);
xor U2534 (N_2534,N_1928,N_2377);
or U2535 (N_2535,N_2039,N_2392);
and U2536 (N_2536,N_2239,N_1814);
nor U2537 (N_2537,N_1805,N_1907);
nor U2538 (N_2538,N_1963,N_2138);
nor U2539 (N_2539,N_2188,N_2052);
nand U2540 (N_2540,N_2051,N_2277);
or U2541 (N_2541,N_2255,N_2090);
xor U2542 (N_2542,N_2272,N_2316);
or U2543 (N_2543,N_2278,N_2011);
nor U2544 (N_2544,N_2170,N_2088);
nor U2545 (N_2545,N_2103,N_1874);
xor U2546 (N_2546,N_2145,N_2004);
and U2547 (N_2547,N_2356,N_2231);
or U2548 (N_2548,N_2115,N_2308);
or U2549 (N_2549,N_1969,N_2382);
nand U2550 (N_2550,N_2057,N_1904);
and U2551 (N_2551,N_2339,N_2368);
nand U2552 (N_2552,N_2009,N_2022);
nand U2553 (N_2553,N_2157,N_2256);
or U2554 (N_2554,N_2084,N_2149);
nor U2555 (N_2555,N_1876,N_2073);
xnor U2556 (N_2556,N_2123,N_1912);
nand U2557 (N_2557,N_2007,N_2137);
and U2558 (N_2558,N_2048,N_2276);
nand U2559 (N_2559,N_2104,N_2299);
or U2560 (N_2560,N_2086,N_1846);
nor U2561 (N_2561,N_2270,N_2109);
nand U2562 (N_2562,N_2041,N_1801);
nor U2563 (N_2563,N_1976,N_1813);
and U2564 (N_2564,N_2364,N_1873);
nor U2565 (N_2565,N_2342,N_2247);
or U2566 (N_2566,N_2092,N_2205);
nor U2567 (N_2567,N_2386,N_2125);
and U2568 (N_2568,N_2315,N_2362);
nand U2569 (N_2569,N_2080,N_2312);
nand U2570 (N_2570,N_2165,N_2059);
or U2571 (N_2571,N_2013,N_1930);
nor U2572 (N_2572,N_1915,N_2063);
and U2573 (N_2573,N_2215,N_1830);
xor U2574 (N_2574,N_1906,N_2206);
nand U2575 (N_2575,N_1908,N_2106);
or U2576 (N_2576,N_1865,N_2152);
or U2577 (N_2577,N_1981,N_2100);
and U2578 (N_2578,N_2323,N_2064);
or U2579 (N_2579,N_1909,N_1819);
and U2580 (N_2580,N_1911,N_2120);
nand U2581 (N_2581,N_1958,N_2245);
or U2582 (N_2582,N_1921,N_1989);
or U2583 (N_2583,N_2281,N_1996);
or U2584 (N_2584,N_2093,N_2298);
and U2585 (N_2585,N_2381,N_2252);
xor U2586 (N_2586,N_1809,N_2337);
or U2587 (N_2587,N_1877,N_2345);
xnor U2588 (N_2588,N_2076,N_2394);
xor U2589 (N_2589,N_2354,N_2014);
or U2590 (N_2590,N_1941,N_2351);
nand U2591 (N_2591,N_2373,N_2329);
nor U2592 (N_2592,N_2242,N_1889);
xor U2593 (N_2593,N_2163,N_2075);
and U2594 (N_2594,N_1858,N_2233);
xnor U2595 (N_2595,N_1825,N_1812);
nand U2596 (N_2596,N_2193,N_1923);
or U2597 (N_2597,N_1833,N_2218);
nand U2598 (N_2598,N_2271,N_2360);
or U2599 (N_2599,N_2375,N_1933);
nand U2600 (N_2600,N_1867,N_2290);
nand U2601 (N_2601,N_1920,N_2072);
or U2602 (N_2602,N_1925,N_1902);
nor U2603 (N_2603,N_2269,N_1929);
or U2604 (N_2604,N_1900,N_2330);
xnor U2605 (N_2605,N_1822,N_2229);
nor U2606 (N_2606,N_1896,N_1999);
nand U2607 (N_2607,N_2154,N_1880);
nor U2608 (N_2608,N_2129,N_2174);
nor U2609 (N_2609,N_1824,N_2047);
nand U2610 (N_2610,N_2111,N_2019);
nand U2611 (N_2611,N_2297,N_2253);
and U2612 (N_2612,N_2065,N_1820);
nand U2613 (N_2613,N_1988,N_1884);
or U2614 (N_2614,N_1994,N_2232);
and U2615 (N_2615,N_1934,N_2196);
xor U2616 (N_2616,N_1854,N_2156);
or U2617 (N_2617,N_1845,N_2045);
nor U2618 (N_2618,N_2189,N_2275);
and U2619 (N_2619,N_2376,N_1945);
and U2620 (N_2620,N_1837,N_1827);
nand U2621 (N_2621,N_2177,N_2328);
and U2622 (N_2622,N_2212,N_1808);
and U2623 (N_2623,N_1938,N_2332);
xnor U2624 (N_2624,N_2282,N_2024);
xnor U2625 (N_2625,N_2335,N_2304);
or U2626 (N_2626,N_2112,N_2359);
or U2627 (N_2627,N_2142,N_2018);
and U2628 (N_2628,N_1993,N_1864);
or U2629 (N_2629,N_1987,N_2162);
xor U2630 (N_2630,N_2008,N_2263);
nand U2631 (N_2631,N_1991,N_2203);
or U2632 (N_2632,N_2248,N_2173);
and U2633 (N_2633,N_2140,N_1979);
xor U2634 (N_2634,N_2221,N_1860);
or U2635 (N_2635,N_1810,N_2182);
xnor U2636 (N_2636,N_2096,N_1998);
and U2637 (N_2637,N_2211,N_2288);
or U2638 (N_2638,N_2191,N_1899);
xor U2639 (N_2639,N_2389,N_2003);
nand U2640 (N_2640,N_2262,N_2124);
nor U2641 (N_2641,N_2033,N_2198);
nand U2642 (N_2642,N_2002,N_1990);
nor U2643 (N_2643,N_2309,N_2384);
and U2644 (N_2644,N_2069,N_2136);
nor U2645 (N_2645,N_1937,N_2307);
nor U2646 (N_2646,N_2397,N_2200);
nand U2647 (N_2647,N_2334,N_1966);
nor U2648 (N_2648,N_2331,N_2185);
nor U2649 (N_2649,N_2139,N_2132);
nand U2650 (N_2650,N_2294,N_2287);
nand U2651 (N_2651,N_2367,N_2279);
and U2652 (N_2652,N_2091,N_2128);
nand U2653 (N_2653,N_2371,N_2097);
or U2654 (N_2654,N_2224,N_1834);
nand U2655 (N_2655,N_1821,N_2046);
nand U2656 (N_2656,N_2320,N_1828);
and U2657 (N_2657,N_2388,N_2034);
xnor U2658 (N_2658,N_1946,N_1817);
or U2659 (N_2659,N_2186,N_1885);
nor U2660 (N_2660,N_1959,N_2230);
nand U2661 (N_2661,N_1888,N_2210);
or U2662 (N_2662,N_1982,N_1800);
or U2663 (N_2663,N_2398,N_1875);
nand U2664 (N_2664,N_1995,N_1804);
and U2665 (N_2665,N_1983,N_1977);
xnor U2666 (N_2666,N_2130,N_2213);
xor U2667 (N_2667,N_2116,N_2147);
or U2668 (N_2668,N_2199,N_2028);
xor U2669 (N_2669,N_1894,N_1975);
and U2670 (N_2670,N_2319,N_2113);
nand U2671 (N_2671,N_2216,N_2363);
xor U2672 (N_2672,N_2250,N_2159);
xnor U2673 (N_2673,N_1960,N_2127);
xor U2674 (N_2674,N_2164,N_1862);
and U2675 (N_2675,N_1848,N_2148);
nor U2676 (N_2676,N_2391,N_2017);
and U2677 (N_2677,N_2260,N_2030);
nand U2678 (N_2678,N_2040,N_2190);
or U2679 (N_2679,N_2313,N_2102);
nand U2680 (N_2680,N_2056,N_2184);
nand U2681 (N_2681,N_2134,N_2226);
or U2682 (N_2682,N_2153,N_2160);
nor U2683 (N_2683,N_1947,N_2207);
nor U2684 (N_2684,N_2296,N_1968);
xnor U2685 (N_2685,N_2300,N_1869);
nor U2686 (N_2686,N_2340,N_2259);
nor U2687 (N_2687,N_2241,N_2303);
xor U2688 (N_2688,N_2118,N_1916);
nor U2689 (N_2689,N_1829,N_1835);
xnor U2690 (N_2690,N_1985,N_1853);
or U2691 (N_2691,N_2000,N_2010);
nor U2692 (N_2692,N_2261,N_1892);
xnor U2693 (N_2693,N_1951,N_2082);
nand U2694 (N_2694,N_2322,N_2068);
or U2695 (N_2695,N_1992,N_2346);
or U2696 (N_2696,N_2061,N_2131);
and U2697 (N_2697,N_2105,N_2121);
xnor U2698 (N_2698,N_2114,N_2378);
xor U2699 (N_2699,N_2098,N_2285);
or U2700 (N_2700,N_2367,N_1824);
nor U2701 (N_2701,N_1881,N_2013);
or U2702 (N_2702,N_2341,N_2196);
or U2703 (N_2703,N_1939,N_1883);
xnor U2704 (N_2704,N_2024,N_2257);
nor U2705 (N_2705,N_2064,N_1834);
or U2706 (N_2706,N_2163,N_1966);
and U2707 (N_2707,N_2376,N_2179);
or U2708 (N_2708,N_2096,N_1842);
xor U2709 (N_2709,N_1805,N_2224);
and U2710 (N_2710,N_2073,N_2043);
xnor U2711 (N_2711,N_2228,N_1848);
nand U2712 (N_2712,N_2265,N_1999);
or U2713 (N_2713,N_2266,N_1920);
and U2714 (N_2714,N_1848,N_2121);
and U2715 (N_2715,N_2227,N_2251);
or U2716 (N_2716,N_1915,N_2239);
xnor U2717 (N_2717,N_2179,N_2373);
nor U2718 (N_2718,N_2057,N_2056);
nand U2719 (N_2719,N_2212,N_2127);
or U2720 (N_2720,N_2110,N_2310);
and U2721 (N_2721,N_2366,N_1823);
and U2722 (N_2722,N_2314,N_1878);
nand U2723 (N_2723,N_2330,N_2395);
nor U2724 (N_2724,N_2276,N_2299);
nand U2725 (N_2725,N_2184,N_1863);
nor U2726 (N_2726,N_1980,N_1846);
nand U2727 (N_2727,N_2361,N_1842);
nand U2728 (N_2728,N_1906,N_2166);
xor U2729 (N_2729,N_2127,N_2292);
nor U2730 (N_2730,N_2080,N_1964);
and U2731 (N_2731,N_2120,N_2102);
nor U2732 (N_2732,N_2308,N_2157);
and U2733 (N_2733,N_2331,N_1968);
nand U2734 (N_2734,N_2281,N_2282);
nor U2735 (N_2735,N_2034,N_2341);
xor U2736 (N_2736,N_1920,N_1843);
nand U2737 (N_2737,N_2167,N_2376);
nand U2738 (N_2738,N_2229,N_2221);
and U2739 (N_2739,N_2169,N_2089);
nand U2740 (N_2740,N_2093,N_1880);
xor U2741 (N_2741,N_2275,N_2337);
nor U2742 (N_2742,N_1957,N_2121);
nor U2743 (N_2743,N_1883,N_2215);
and U2744 (N_2744,N_1939,N_2337);
xnor U2745 (N_2745,N_1927,N_2135);
nand U2746 (N_2746,N_2165,N_1994);
nand U2747 (N_2747,N_2363,N_2336);
nor U2748 (N_2748,N_2062,N_2271);
nor U2749 (N_2749,N_1829,N_1844);
and U2750 (N_2750,N_1988,N_2050);
xnor U2751 (N_2751,N_1864,N_2180);
or U2752 (N_2752,N_1962,N_2330);
nor U2753 (N_2753,N_2086,N_2348);
nor U2754 (N_2754,N_2047,N_2372);
or U2755 (N_2755,N_2206,N_2088);
nand U2756 (N_2756,N_2200,N_2332);
xnor U2757 (N_2757,N_1966,N_2301);
nand U2758 (N_2758,N_2008,N_2205);
and U2759 (N_2759,N_2039,N_1807);
or U2760 (N_2760,N_2356,N_1829);
nor U2761 (N_2761,N_1965,N_2113);
nand U2762 (N_2762,N_2104,N_2349);
xor U2763 (N_2763,N_2016,N_2117);
xnor U2764 (N_2764,N_2195,N_2242);
nand U2765 (N_2765,N_2205,N_2141);
and U2766 (N_2766,N_2296,N_2083);
nor U2767 (N_2767,N_2142,N_2355);
or U2768 (N_2768,N_2058,N_2244);
xnor U2769 (N_2769,N_1824,N_2175);
nor U2770 (N_2770,N_2271,N_1986);
and U2771 (N_2771,N_2008,N_2336);
or U2772 (N_2772,N_2093,N_2338);
or U2773 (N_2773,N_1844,N_1951);
nand U2774 (N_2774,N_2012,N_1907);
and U2775 (N_2775,N_1956,N_1879);
nor U2776 (N_2776,N_2114,N_2185);
nor U2777 (N_2777,N_2190,N_1879);
or U2778 (N_2778,N_1968,N_1871);
nor U2779 (N_2779,N_2371,N_2144);
nor U2780 (N_2780,N_2191,N_2207);
xnor U2781 (N_2781,N_1993,N_1813);
and U2782 (N_2782,N_2289,N_1964);
and U2783 (N_2783,N_1961,N_1856);
nand U2784 (N_2784,N_2273,N_1934);
nand U2785 (N_2785,N_2224,N_2240);
or U2786 (N_2786,N_1817,N_2006);
nor U2787 (N_2787,N_2069,N_2234);
nor U2788 (N_2788,N_1947,N_2062);
or U2789 (N_2789,N_2301,N_2113);
and U2790 (N_2790,N_2109,N_2369);
and U2791 (N_2791,N_1895,N_2283);
xnor U2792 (N_2792,N_2346,N_1961);
nor U2793 (N_2793,N_2110,N_2135);
nor U2794 (N_2794,N_2264,N_2027);
or U2795 (N_2795,N_2137,N_2014);
and U2796 (N_2796,N_1904,N_1884);
nand U2797 (N_2797,N_2055,N_1956);
nand U2798 (N_2798,N_2349,N_1837);
and U2799 (N_2799,N_2356,N_2060);
and U2800 (N_2800,N_1904,N_1987);
or U2801 (N_2801,N_2124,N_1897);
and U2802 (N_2802,N_1873,N_1843);
and U2803 (N_2803,N_2072,N_1811);
or U2804 (N_2804,N_2093,N_2394);
nand U2805 (N_2805,N_2022,N_1894);
nand U2806 (N_2806,N_2232,N_2393);
nor U2807 (N_2807,N_2022,N_1813);
xnor U2808 (N_2808,N_1803,N_1971);
nand U2809 (N_2809,N_2028,N_1990);
xnor U2810 (N_2810,N_1978,N_2210);
xor U2811 (N_2811,N_2375,N_1808);
and U2812 (N_2812,N_2369,N_2205);
nor U2813 (N_2813,N_1834,N_2151);
nand U2814 (N_2814,N_1903,N_2133);
and U2815 (N_2815,N_2267,N_1946);
or U2816 (N_2816,N_2094,N_1926);
xnor U2817 (N_2817,N_1816,N_2391);
nor U2818 (N_2818,N_2317,N_2221);
xnor U2819 (N_2819,N_2234,N_1889);
xor U2820 (N_2820,N_2334,N_2295);
nand U2821 (N_2821,N_2276,N_1997);
xor U2822 (N_2822,N_2274,N_2053);
or U2823 (N_2823,N_2246,N_2360);
or U2824 (N_2824,N_2199,N_2184);
nor U2825 (N_2825,N_1810,N_1994);
nor U2826 (N_2826,N_2207,N_2278);
nor U2827 (N_2827,N_2252,N_2148);
nor U2828 (N_2828,N_2172,N_2045);
or U2829 (N_2829,N_2334,N_2027);
xnor U2830 (N_2830,N_1888,N_2165);
xor U2831 (N_2831,N_2087,N_2208);
xor U2832 (N_2832,N_1838,N_1809);
xnor U2833 (N_2833,N_2003,N_1973);
nor U2834 (N_2834,N_1844,N_2347);
nand U2835 (N_2835,N_1852,N_2352);
nor U2836 (N_2836,N_2018,N_1813);
xnor U2837 (N_2837,N_2114,N_2332);
xor U2838 (N_2838,N_2208,N_2032);
xor U2839 (N_2839,N_2244,N_2188);
nor U2840 (N_2840,N_2130,N_2180);
or U2841 (N_2841,N_2315,N_2368);
or U2842 (N_2842,N_2173,N_2107);
or U2843 (N_2843,N_2393,N_2041);
nor U2844 (N_2844,N_2144,N_2091);
and U2845 (N_2845,N_2193,N_2106);
nand U2846 (N_2846,N_1855,N_1809);
nand U2847 (N_2847,N_1934,N_2365);
xnor U2848 (N_2848,N_2129,N_2372);
or U2849 (N_2849,N_2130,N_2263);
xor U2850 (N_2850,N_1999,N_2353);
and U2851 (N_2851,N_1881,N_2333);
xor U2852 (N_2852,N_1910,N_1806);
and U2853 (N_2853,N_1983,N_2361);
xnor U2854 (N_2854,N_1927,N_1847);
or U2855 (N_2855,N_2040,N_2091);
and U2856 (N_2856,N_2285,N_1950);
xor U2857 (N_2857,N_2142,N_1944);
and U2858 (N_2858,N_1957,N_2072);
or U2859 (N_2859,N_1876,N_1965);
and U2860 (N_2860,N_2225,N_1882);
nand U2861 (N_2861,N_1838,N_2299);
xor U2862 (N_2862,N_2327,N_2061);
nor U2863 (N_2863,N_2336,N_2052);
or U2864 (N_2864,N_2307,N_2354);
and U2865 (N_2865,N_2211,N_1955);
nand U2866 (N_2866,N_2268,N_2376);
and U2867 (N_2867,N_2370,N_1886);
nand U2868 (N_2868,N_2099,N_1989);
xor U2869 (N_2869,N_2255,N_2195);
or U2870 (N_2870,N_2289,N_2275);
nand U2871 (N_2871,N_2159,N_1962);
or U2872 (N_2872,N_2206,N_2233);
nand U2873 (N_2873,N_2235,N_1970);
or U2874 (N_2874,N_2143,N_1894);
nand U2875 (N_2875,N_1942,N_2365);
nand U2876 (N_2876,N_2093,N_2160);
nor U2877 (N_2877,N_2108,N_2211);
and U2878 (N_2878,N_1996,N_2173);
or U2879 (N_2879,N_2374,N_2076);
and U2880 (N_2880,N_2092,N_2221);
and U2881 (N_2881,N_2244,N_2213);
nor U2882 (N_2882,N_1860,N_2272);
or U2883 (N_2883,N_2265,N_2105);
or U2884 (N_2884,N_2126,N_2075);
nor U2885 (N_2885,N_1942,N_2104);
or U2886 (N_2886,N_2068,N_1938);
or U2887 (N_2887,N_2192,N_2054);
or U2888 (N_2888,N_2397,N_2001);
nor U2889 (N_2889,N_1958,N_2267);
nor U2890 (N_2890,N_2256,N_2111);
and U2891 (N_2891,N_2065,N_1894);
or U2892 (N_2892,N_1982,N_1937);
or U2893 (N_2893,N_2274,N_2249);
and U2894 (N_2894,N_2343,N_1931);
nor U2895 (N_2895,N_2311,N_1867);
or U2896 (N_2896,N_2288,N_1960);
or U2897 (N_2897,N_2072,N_2399);
nor U2898 (N_2898,N_1835,N_2159);
nand U2899 (N_2899,N_1916,N_1858);
nand U2900 (N_2900,N_1984,N_2059);
nand U2901 (N_2901,N_2395,N_2088);
nor U2902 (N_2902,N_2204,N_2152);
nand U2903 (N_2903,N_1898,N_1982);
and U2904 (N_2904,N_1889,N_1926);
nand U2905 (N_2905,N_2176,N_2100);
or U2906 (N_2906,N_2185,N_1840);
or U2907 (N_2907,N_2071,N_2316);
nor U2908 (N_2908,N_2240,N_2359);
and U2909 (N_2909,N_2381,N_2276);
nor U2910 (N_2910,N_1868,N_2162);
nand U2911 (N_2911,N_2174,N_1903);
nor U2912 (N_2912,N_2253,N_1957);
nor U2913 (N_2913,N_2310,N_2356);
or U2914 (N_2914,N_1990,N_1967);
and U2915 (N_2915,N_1999,N_2163);
nor U2916 (N_2916,N_1804,N_2252);
nor U2917 (N_2917,N_1890,N_2159);
nand U2918 (N_2918,N_1808,N_1980);
xnor U2919 (N_2919,N_1883,N_1969);
nor U2920 (N_2920,N_2359,N_2311);
xor U2921 (N_2921,N_1843,N_1997);
xor U2922 (N_2922,N_1960,N_2017);
or U2923 (N_2923,N_2352,N_2182);
xor U2924 (N_2924,N_2060,N_1972);
and U2925 (N_2925,N_2121,N_2189);
and U2926 (N_2926,N_2165,N_1800);
nand U2927 (N_2927,N_1849,N_2143);
and U2928 (N_2928,N_1836,N_2079);
or U2929 (N_2929,N_1996,N_1891);
nor U2930 (N_2930,N_1828,N_2366);
or U2931 (N_2931,N_2184,N_2201);
and U2932 (N_2932,N_2053,N_1823);
xor U2933 (N_2933,N_1935,N_1887);
nor U2934 (N_2934,N_2203,N_1969);
and U2935 (N_2935,N_2390,N_2046);
nand U2936 (N_2936,N_1900,N_1920);
nor U2937 (N_2937,N_1972,N_2220);
xor U2938 (N_2938,N_2151,N_2128);
nor U2939 (N_2939,N_2289,N_2040);
nand U2940 (N_2940,N_2370,N_2396);
nor U2941 (N_2941,N_1917,N_2021);
nand U2942 (N_2942,N_2309,N_2079);
and U2943 (N_2943,N_1965,N_1973);
or U2944 (N_2944,N_2081,N_2049);
or U2945 (N_2945,N_1840,N_1821);
and U2946 (N_2946,N_2298,N_1819);
and U2947 (N_2947,N_2222,N_2363);
and U2948 (N_2948,N_2302,N_2247);
nor U2949 (N_2949,N_2180,N_1945);
or U2950 (N_2950,N_2120,N_1950);
xnor U2951 (N_2951,N_2369,N_1918);
xnor U2952 (N_2952,N_2028,N_1887);
or U2953 (N_2953,N_2290,N_2270);
nor U2954 (N_2954,N_1808,N_2381);
and U2955 (N_2955,N_2307,N_1805);
or U2956 (N_2956,N_2359,N_1846);
nor U2957 (N_2957,N_1956,N_2040);
and U2958 (N_2958,N_2228,N_2338);
nand U2959 (N_2959,N_2141,N_2075);
xor U2960 (N_2960,N_2281,N_2066);
xor U2961 (N_2961,N_1952,N_2318);
nand U2962 (N_2962,N_2380,N_2308);
nand U2963 (N_2963,N_2204,N_1820);
or U2964 (N_2964,N_2193,N_2074);
and U2965 (N_2965,N_2032,N_2268);
nand U2966 (N_2966,N_2349,N_2159);
nand U2967 (N_2967,N_2074,N_1890);
nor U2968 (N_2968,N_2018,N_2358);
and U2969 (N_2969,N_2202,N_1986);
and U2970 (N_2970,N_2112,N_2322);
xor U2971 (N_2971,N_1998,N_1946);
nor U2972 (N_2972,N_2143,N_1860);
or U2973 (N_2973,N_2158,N_2229);
nand U2974 (N_2974,N_2073,N_2127);
and U2975 (N_2975,N_2368,N_1908);
or U2976 (N_2976,N_2300,N_2083);
nor U2977 (N_2977,N_2234,N_2096);
and U2978 (N_2978,N_2165,N_2305);
nand U2979 (N_2979,N_2301,N_1981);
nand U2980 (N_2980,N_2374,N_2237);
and U2981 (N_2981,N_1883,N_2210);
nand U2982 (N_2982,N_2279,N_2085);
xnor U2983 (N_2983,N_2148,N_1923);
and U2984 (N_2984,N_2322,N_2392);
and U2985 (N_2985,N_2341,N_2098);
xnor U2986 (N_2986,N_1853,N_2097);
nand U2987 (N_2987,N_1963,N_1977);
xor U2988 (N_2988,N_1828,N_2365);
and U2989 (N_2989,N_2299,N_2026);
or U2990 (N_2990,N_2383,N_2202);
or U2991 (N_2991,N_2227,N_1816);
nor U2992 (N_2992,N_1837,N_1927);
or U2993 (N_2993,N_2395,N_2304);
or U2994 (N_2994,N_1922,N_1973);
and U2995 (N_2995,N_1925,N_2395);
nand U2996 (N_2996,N_2020,N_2284);
nand U2997 (N_2997,N_1849,N_1926);
nor U2998 (N_2998,N_1943,N_2047);
nor U2999 (N_2999,N_2348,N_2271);
or U3000 (N_3000,N_2572,N_2412);
nand U3001 (N_3001,N_2592,N_2687);
nor U3002 (N_3002,N_2463,N_2977);
or U3003 (N_3003,N_2996,N_2768);
or U3004 (N_3004,N_2929,N_2670);
xor U3005 (N_3005,N_2487,N_2739);
nor U3006 (N_3006,N_2881,N_2800);
and U3007 (N_3007,N_2656,N_2404);
xnor U3008 (N_3008,N_2856,N_2425);
nor U3009 (N_3009,N_2526,N_2819);
nand U3010 (N_3010,N_2461,N_2585);
nor U3011 (N_3011,N_2787,N_2569);
and U3012 (N_3012,N_2518,N_2657);
or U3013 (N_3013,N_2440,N_2565);
xor U3014 (N_3014,N_2707,N_2788);
or U3015 (N_3015,N_2980,N_2459);
xnor U3016 (N_3016,N_2488,N_2866);
or U3017 (N_3017,N_2413,N_2556);
nor U3018 (N_3018,N_2807,N_2545);
or U3019 (N_3019,N_2893,N_2988);
or U3020 (N_3020,N_2533,N_2611);
nand U3021 (N_3021,N_2916,N_2719);
xnor U3022 (N_3022,N_2780,N_2734);
and U3023 (N_3023,N_2862,N_2990);
nor U3024 (N_3024,N_2897,N_2457);
nand U3025 (N_3025,N_2955,N_2474);
nand U3026 (N_3026,N_2825,N_2653);
xor U3027 (N_3027,N_2715,N_2508);
nand U3028 (N_3028,N_2789,N_2857);
nor U3029 (N_3029,N_2541,N_2723);
xnor U3030 (N_3030,N_2965,N_2493);
xnor U3031 (N_3031,N_2671,N_2655);
nor U3032 (N_3032,N_2668,N_2675);
and U3033 (N_3033,N_2809,N_2926);
xnor U3034 (N_3034,N_2415,N_2625);
xor U3035 (N_3035,N_2626,N_2953);
nand U3036 (N_3036,N_2753,N_2843);
nor U3037 (N_3037,N_2957,N_2860);
nor U3038 (N_3038,N_2513,N_2478);
or U3039 (N_3039,N_2669,N_2535);
or U3040 (N_3040,N_2970,N_2551);
and U3041 (N_3041,N_2662,N_2797);
xnor U3042 (N_3042,N_2660,N_2839);
nand U3043 (N_3043,N_2490,N_2818);
or U3044 (N_3044,N_2554,N_2775);
xnor U3045 (N_3045,N_2760,N_2641);
xor U3046 (N_3046,N_2555,N_2450);
nand U3047 (N_3047,N_2885,N_2917);
or U3048 (N_3048,N_2959,N_2773);
or U3049 (N_3049,N_2510,N_2878);
nand U3050 (N_3050,N_2927,N_2647);
xor U3051 (N_3051,N_2920,N_2691);
or U3052 (N_3052,N_2446,N_2613);
nand U3053 (N_3053,N_2880,N_2405);
and U3054 (N_3054,N_2741,N_2979);
xor U3055 (N_3055,N_2882,N_2910);
nand U3056 (N_3056,N_2930,N_2601);
nor U3057 (N_3057,N_2582,N_2477);
nor U3058 (N_3058,N_2663,N_2874);
nand U3059 (N_3059,N_2530,N_2941);
xnor U3060 (N_3060,N_2559,N_2599);
and U3061 (N_3061,N_2690,N_2804);
nand U3062 (N_3062,N_2600,N_2672);
nor U3063 (N_3063,N_2429,N_2482);
and U3064 (N_3064,N_2875,N_2982);
xor U3065 (N_3065,N_2409,N_2822);
or U3066 (N_3066,N_2686,N_2658);
and U3067 (N_3067,N_2987,N_2496);
xor U3068 (N_3068,N_2725,N_2886);
and U3069 (N_3069,N_2749,N_2593);
or U3070 (N_3070,N_2869,N_2876);
nor U3071 (N_3071,N_2542,N_2639);
or U3072 (N_3072,N_2747,N_2603);
xor U3073 (N_3073,N_2423,N_2441);
nand U3074 (N_3074,N_2840,N_2435);
or U3075 (N_3075,N_2701,N_2735);
nand U3076 (N_3076,N_2752,N_2891);
xnor U3077 (N_3077,N_2512,N_2589);
or U3078 (N_3078,N_2769,N_2673);
or U3079 (N_3079,N_2418,N_2434);
nand U3080 (N_3080,N_2790,N_2424);
or U3081 (N_3081,N_2705,N_2850);
nand U3082 (N_3082,N_2708,N_2794);
and U3083 (N_3083,N_2894,N_2630);
xnor U3084 (N_3084,N_2448,N_2830);
nor U3085 (N_3085,N_2628,N_2938);
nand U3086 (N_3086,N_2431,N_2721);
and U3087 (N_3087,N_2740,N_2823);
and U3088 (N_3088,N_2754,N_2438);
nand U3089 (N_3089,N_2475,N_2652);
xor U3090 (N_3090,N_2607,N_2612);
nor U3091 (N_3091,N_2852,N_2619);
nor U3092 (N_3092,N_2855,N_2720);
nor U3093 (N_3093,N_2709,N_2661);
nand U3094 (N_3094,N_2810,N_2714);
or U3095 (N_3095,N_2873,N_2473);
or U3096 (N_3096,N_2956,N_2692);
or U3097 (N_3097,N_2858,N_2470);
nand U3098 (N_3098,N_2756,N_2943);
nor U3099 (N_3099,N_2727,N_2598);
nor U3100 (N_3100,N_2901,N_2617);
xnor U3101 (N_3101,N_2845,N_2932);
nor U3102 (N_3102,N_2527,N_2703);
and U3103 (N_3103,N_2900,N_2785);
and U3104 (N_3104,N_2560,N_2733);
nand U3105 (N_3105,N_2765,N_2828);
or U3106 (N_3106,N_2865,N_2937);
nand U3107 (N_3107,N_2689,N_2737);
xnor U3108 (N_3108,N_2602,N_2417);
nand U3109 (N_3109,N_2544,N_2574);
nor U3110 (N_3110,N_2934,N_2499);
nand U3111 (N_3111,N_2922,N_2525);
xnor U3112 (N_3112,N_2577,N_2514);
nor U3113 (N_3113,N_2966,N_2743);
nand U3114 (N_3114,N_2498,N_2576);
and U3115 (N_3115,N_2460,N_2581);
xor U3116 (N_3116,N_2694,N_2745);
or U3117 (N_3117,N_2835,N_2864);
nor U3118 (N_3118,N_2436,N_2651);
nor U3119 (N_3119,N_2700,N_2584);
and U3120 (N_3120,N_2587,N_2444);
nand U3121 (N_3121,N_2958,N_2933);
and U3122 (N_3122,N_2401,N_2432);
or U3123 (N_3123,N_2764,N_2468);
or U3124 (N_3124,N_2420,N_2467);
xnor U3125 (N_3125,N_2458,N_2706);
and U3126 (N_3126,N_2770,N_2763);
xnor U3127 (N_3127,N_2520,N_2515);
and U3128 (N_3128,N_2433,N_2443);
and U3129 (N_3129,N_2679,N_2967);
xnor U3130 (N_3130,N_2867,N_2791);
nand U3131 (N_3131,N_2975,N_2744);
or U3132 (N_3132,N_2954,N_2456);
and U3133 (N_3133,N_2403,N_2567);
xor U3134 (N_3134,N_2573,N_2903);
or U3135 (N_3135,N_2636,N_2447);
nor U3136 (N_3136,N_2833,N_2400);
xor U3137 (N_3137,N_2595,N_2534);
or U3138 (N_3138,N_2615,N_2995);
xnor U3139 (N_3139,N_2622,N_2761);
nand U3140 (N_3140,N_2802,N_2471);
or U3141 (N_3141,N_2472,N_2449);
nand U3142 (N_3142,N_2736,N_2469);
nand U3143 (N_3143,N_2772,N_2521);
nor U3144 (N_3144,N_2631,N_2908);
nand U3145 (N_3145,N_2476,N_2942);
xnor U3146 (N_3146,N_2563,N_2984);
nand U3147 (N_3147,N_2693,N_2517);
and U3148 (N_3148,N_2722,N_2629);
and U3149 (N_3149,N_2516,N_2604);
nand U3150 (N_3150,N_2579,N_2702);
or U3151 (N_3151,N_2522,N_2410);
or U3152 (N_3152,N_2716,N_2879);
nor U3153 (N_3153,N_2549,N_2935);
nor U3154 (N_3154,N_2774,N_2546);
and U3155 (N_3155,N_2895,N_2993);
xor U3156 (N_3156,N_2479,N_2983);
and U3157 (N_3157,N_2899,N_2624);
nor U3158 (N_3158,N_2863,N_2558);
or U3159 (N_3159,N_2590,N_2481);
and U3160 (N_3160,N_2827,N_2548);
or U3161 (N_3161,N_2884,N_2726);
nand U3162 (N_3162,N_2814,N_2644);
xor U3163 (N_3163,N_2543,N_2454);
nor U3164 (N_3164,N_2877,N_2497);
nor U3165 (N_3165,N_2906,N_2989);
nor U3166 (N_3166,N_2553,N_2519);
and U3167 (N_3167,N_2605,N_2986);
nand U3168 (N_3168,N_2883,N_2798);
or U3169 (N_3169,N_2524,N_2832);
nor U3170 (N_3170,N_2698,N_2766);
and U3171 (N_3171,N_2685,N_2750);
and U3172 (N_3172,N_2871,N_2887);
and U3173 (N_3173,N_2892,N_2480);
and U3174 (N_3174,N_2453,N_2696);
or U3175 (N_3175,N_2681,N_2568);
and U3176 (N_3176,N_2643,N_2923);
or U3177 (N_3177,N_2684,N_2466);
xnor U3178 (N_3178,N_2889,N_2495);
nor U3179 (N_3179,N_2776,N_2724);
xnor U3180 (N_3180,N_2821,N_2426);
or U3181 (N_3181,N_2596,N_2697);
or U3182 (N_3182,N_2969,N_2968);
nand U3183 (N_3183,N_2820,N_2683);
nand U3184 (N_3184,N_2783,N_2571);
nor U3185 (N_3185,N_2909,N_2610);
xnor U3186 (N_3186,N_2635,N_2637);
xnor U3187 (N_3187,N_2854,N_2914);
and U3188 (N_3188,N_2570,N_2925);
and U3189 (N_3189,N_2654,N_2915);
nand U3190 (N_3190,N_2539,N_2971);
xor U3191 (N_3191,N_2678,N_2427);
and U3192 (N_3192,N_2416,N_2936);
nor U3193 (N_3193,N_2506,N_2812);
or U3194 (N_3194,N_2841,N_2564);
or U3195 (N_3195,N_2580,N_2759);
and U3196 (N_3196,N_2547,N_2494);
or U3197 (N_3197,N_2659,N_2826);
or U3198 (N_3198,N_2552,N_2591);
or U3199 (N_3199,N_2680,N_2837);
or U3200 (N_3200,N_2575,N_2407);
or U3201 (N_3201,N_2834,N_2618);
nor U3202 (N_3202,N_2974,N_2844);
or U3203 (N_3203,N_2777,N_2674);
and U3204 (N_3204,N_2712,N_2868);
nor U3205 (N_3205,N_2921,N_2746);
nand U3206 (N_3206,N_2748,N_2949);
and U3207 (N_3207,N_2896,N_2695);
nor U3208 (N_3208,N_2406,N_2803);
nand U3209 (N_3209,N_2699,N_2588);
and U3210 (N_3210,N_2540,N_2484);
and U3211 (N_3211,N_2872,N_2911);
or U3212 (N_3212,N_2945,N_2751);
or U3213 (N_3213,N_2437,N_2642);
nor U3214 (N_3214,N_2728,N_2831);
nor U3215 (N_3215,N_2606,N_2952);
nor U3216 (N_3216,N_2985,N_2732);
and U3217 (N_3217,N_2950,N_2904);
or U3218 (N_3218,N_2946,N_2861);
nand U3219 (N_3219,N_2742,N_2963);
and U3220 (N_3220,N_2805,N_2502);
xor U3221 (N_3221,N_2561,N_2586);
xnor U3222 (N_3222,N_2489,N_2758);
and U3223 (N_3223,N_2503,N_2778);
and U3224 (N_3224,N_2870,N_2677);
or U3225 (N_3225,N_2795,N_2428);
and U3226 (N_3226,N_2729,N_2757);
nand U3227 (N_3227,N_2650,N_2710);
or U3228 (N_3228,N_2718,N_2648);
or U3229 (N_3229,N_2947,N_2851);
and U3230 (N_3230,N_2859,N_2817);
nor U3231 (N_3231,N_2492,N_2940);
nor U3232 (N_3232,N_2755,N_2597);
or U3233 (N_3233,N_2531,N_2439);
xor U3234 (N_3234,N_2638,N_2928);
nor U3235 (N_3235,N_2815,N_2731);
nor U3236 (N_3236,N_2623,N_2528);
nor U3237 (N_3237,N_2538,N_2888);
or U3238 (N_3238,N_2455,N_2537);
or U3239 (N_3239,N_2421,N_2646);
nand U3240 (N_3240,N_2848,N_2614);
and U3241 (N_3241,N_2616,N_2451);
nor U3242 (N_3242,N_2430,N_2442);
xnor U3243 (N_3243,N_2462,N_2594);
xor U3244 (N_3244,N_2813,N_2445);
nand U3245 (N_3245,N_2792,N_2847);
nor U3246 (N_3246,N_2676,N_2666);
xnor U3247 (N_3247,N_2486,N_2767);
xnor U3248 (N_3248,N_2505,N_2711);
or U3249 (N_3249,N_2717,N_2464);
and U3250 (N_3250,N_2411,N_2452);
or U3251 (N_3251,N_2529,N_2999);
and U3252 (N_3252,N_2536,N_2665);
nor U3253 (N_3253,N_2784,N_2501);
or U3254 (N_3254,N_2829,N_2890);
or U3255 (N_3255,N_2846,N_2939);
nor U3256 (N_3256,N_2924,N_2500);
and U3257 (N_3257,N_2816,N_2664);
xnor U3258 (N_3258,N_2913,N_2782);
nand U3259 (N_3259,N_2981,N_2634);
nor U3260 (N_3260,N_2557,N_2507);
xor U3261 (N_3261,N_2801,N_2978);
nor U3262 (N_3262,N_2998,N_2972);
nand U3263 (N_3263,N_2997,N_2808);
or U3264 (N_3264,N_2902,N_2912);
or U3265 (N_3265,N_2645,N_2608);
and U3266 (N_3266,N_2994,N_2562);
nand U3267 (N_3267,N_2483,N_2991);
and U3268 (N_3268,N_2771,N_2627);
nor U3269 (N_3269,N_2799,N_2640);
or U3270 (N_3270,N_2786,N_2973);
nor U3271 (N_3271,N_2849,N_2853);
and U3272 (N_3272,N_2609,N_2632);
or U3273 (N_3273,N_2649,N_2621);
nor U3274 (N_3274,N_2944,N_2465);
and U3275 (N_3275,N_2811,N_2485);
xnor U3276 (N_3276,N_2419,N_2781);
xnor U3277 (N_3277,N_2730,N_2713);
or U3278 (N_3278,N_2402,N_2620);
nand U3279 (N_3279,N_2836,N_2414);
nand U3280 (N_3280,N_2566,N_2796);
xor U3281 (N_3281,N_2704,N_2682);
or U3282 (N_3282,N_2907,N_2842);
nor U3283 (N_3283,N_2633,N_2583);
or U3284 (N_3284,N_2550,N_2779);
nand U3285 (N_3285,N_2511,N_2688);
nand U3286 (N_3286,N_2931,N_2422);
nand U3287 (N_3287,N_2948,N_2578);
nand U3288 (N_3288,N_2793,N_2960);
or U3289 (N_3289,N_2961,N_2919);
or U3290 (N_3290,N_2806,N_2509);
and U3291 (N_3291,N_2838,N_2504);
nand U3292 (N_3292,N_2824,N_2738);
or U3293 (N_3293,N_2523,N_2898);
nand U3294 (N_3294,N_2976,N_2964);
nor U3295 (N_3295,N_2762,N_2408);
xnor U3296 (N_3296,N_2667,N_2905);
nor U3297 (N_3297,N_2491,N_2992);
nor U3298 (N_3298,N_2532,N_2918);
nor U3299 (N_3299,N_2951,N_2962);
nor U3300 (N_3300,N_2558,N_2595);
or U3301 (N_3301,N_2796,N_2473);
nand U3302 (N_3302,N_2463,N_2915);
nor U3303 (N_3303,N_2914,N_2880);
and U3304 (N_3304,N_2944,N_2412);
or U3305 (N_3305,N_2606,N_2521);
or U3306 (N_3306,N_2815,N_2663);
and U3307 (N_3307,N_2414,N_2669);
or U3308 (N_3308,N_2564,N_2629);
nor U3309 (N_3309,N_2585,N_2802);
nor U3310 (N_3310,N_2900,N_2918);
nand U3311 (N_3311,N_2988,N_2663);
nand U3312 (N_3312,N_2421,N_2463);
nand U3313 (N_3313,N_2566,N_2692);
or U3314 (N_3314,N_2402,N_2828);
or U3315 (N_3315,N_2977,N_2950);
nand U3316 (N_3316,N_2655,N_2963);
and U3317 (N_3317,N_2631,N_2763);
xnor U3318 (N_3318,N_2668,N_2925);
or U3319 (N_3319,N_2998,N_2491);
nand U3320 (N_3320,N_2792,N_2855);
and U3321 (N_3321,N_2857,N_2451);
and U3322 (N_3322,N_2797,N_2811);
nand U3323 (N_3323,N_2749,N_2510);
nand U3324 (N_3324,N_2807,N_2505);
nor U3325 (N_3325,N_2954,N_2466);
xor U3326 (N_3326,N_2545,N_2971);
xor U3327 (N_3327,N_2956,N_2780);
or U3328 (N_3328,N_2421,N_2539);
or U3329 (N_3329,N_2591,N_2432);
nand U3330 (N_3330,N_2932,N_2760);
and U3331 (N_3331,N_2585,N_2514);
xnor U3332 (N_3332,N_2644,N_2612);
nor U3333 (N_3333,N_2807,N_2489);
nand U3334 (N_3334,N_2431,N_2422);
or U3335 (N_3335,N_2700,N_2872);
xor U3336 (N_3336,N_2602,N_2444);
and U3337 (N_3337,N_2960,N_2445);
and U3338 (N_3338,N_2960,N_2606);
nor U3339 (N_3339,N_2907,N_2941);
and U3340 (N_3340,N_2730,N_2573);
xnor U3341 (N_3341,N_2913,N_2793);
or U3342 (N_3342,N_2850,N_2667);
nor U3343 (N_3343,N_2618,N_2519);
or U3344 (N_3344,N_2448,N_2424);
and U3345 (N_3345,N_2816,N_2966);
xnor U3346 (N_3346,N_2445,N_2995);
nand U3347 (N_3347,N_2405,N_2571);
xnor U3348 (N_3348,N_2930,N_2780);
and U3349 (N_3349,N_2423,N_2634);
nor U3350 (N_3350,N_2511,N_2664);
xor U3351 (N_3351,N_2814,N_2908);
nand U3352 (N_3352,N_2504,N_2450);
or U3353 (N_3353,N_2801,N_2831);
and U3354 (N_3354,N_2849,N_2594);
nand U3355 (N_3355,N_2555,N_2677);
nor U3356 (N_3356,N_2708,N_2959);
nand U3357 (N_3357,N_2983,N_2508);
nand U3358 (N_3358,N_2948,N_2598);
xor U3359 (N_3359,N_2675,N_2863);
nand U3360 (N_3360,N_2456,N_2486);
or U3361 (N_3361,N_2597,N_2482);
nor U3362 (N_3362,N_2973,N_2706);
or U3363 (N_3363,N_2605,N_2733);
nor U3364 (N_3364,N_2634,N_2726);
or U3365 (N_3365,N_2887,N_2931);
xnor U3366 (N_3366,N_2433,N_2615);
and U3367 (N_3367,N_2676,N_2810);
xor U3368 (N_3368,N_2764,N_2544);
and U3369 (N_3369,N_2944,N_2978);
or U3370 (N_3370,N_2840,N_2429);
or U3371 (N_3371,N_2609,N_2513);
nand U3372 (N_3372,N_2637,N_2748);
or U3373 (N_3373,N_2794,N_2958);
and U3374 (N_3374,N_2550,N_2639);
nor U3375 (N_3375,N_2926,N_2850);
xnor U3376 (N_3376,N_2521,N_2666);
nand U3377 (N_3377,N_2553,N_2762);
nor U3378 (N_3378,N_2540,N_2562);
nor U3379 (N_3379,N_2781,N_2755);
nor U3380 (N_3380,N_2808,N_2919);
or U3381 (N_3381,N_2470,N_2899);
nand U3382 (N_3382,N_2786,N_2884);
nor U3383 (N_3383,N_2726,N_2684);
nand U3384 (N_3384,N_2501,N_2906);
nand U3385 (N_3385,N_2461,N_2811);
and U3386 (N_3386,N_2793,N_2599);
xor U3387 (N_3387,N_2962,N_2507);
or U3388 (N_3388,N_2412,N_2684);
xnor U3389 (N_3389,N_2877,N_2963);
or U3390 (N_3390,N_2499,N_2514);
or U3391 (N_3391,N_2818,N_2935);
and U3392 (N_3392,N_2667,N_2875);
and U3393 (N_3393,N_2926,N_2492);
nor U3394 (N_3394,N_2751,N_2822);
or U3395 (N_3395,N_2941,N_2875);
xor U3396 (N_3396,N_2504,N_2804);
and U3397 (N_3397,N_2771,N_2964);
nor U3398 (N_3398,N_2841,N_2829);
and U3399 (N_3399,N_2769,N_2666);
nand U3400 (N_3400,N_2792,N_2875);
and U3401 (N_3401,N_2754,N_2889);
or U3402 (N_3402,N_2535,N_2492);
nand U3403 (N_3403,N_2801,N_2945);
xor U3404 (N_3404,N_2716,N_2804);
nor U3405 (N_3405,N_2432,N_2536);
nand U3406 (N_3406,N_2413,N_2705);
and U3407 (N_3407,N_2845,N_2690);
xnor U3408 (N_3408,N_2912,N_2874);
and U3409 (N_3409,N_2861,N_2408);
and U3410 (N_3410,N_2784,N_2881);
and U3411 (N_3411,N_2996,N_2739);
or U3412 (N_3412,N_2684,N_2902);
and U3413 (N_3413,N_2628,N_2770);
or U3414 (N_3414,N_2967,N_2630);
nand U3415 (N_3415,N_2573,N_2813);
nand U3416 (N_3416,N_2564,N_2509);
and U3417 (N_3417,N_2875,N_2437);
or U3418 (N_3418,N_2431,N_2504);
nor U3419 (N_3419,N_2622,N_2985);
or U3420 (N_3420,N_2716,N_2524);
xor U3421 (N_3421,N_2736,N_2660);
or U3422 (N_3422,N_2704,N_2486);
nand U3423 (N_3423,N_2582,N_2603);
xnor U3424 (N_3424,N_2772,N_2743);
or U3425 (N_3425,N_2627,N_2886);
nor U3426 (N_3426,N_2826,N_2930);
or U3427 (N_3427,N_2455,N_2416);
nor U3428 (N_3428,N_2772,N_2607);
nor U3429 (N_3429,N_2816,N_2761);
and U3430 (N_3430,N_2689,N_2416);
and U3431 (N_3431,N_2620,N_2912);
nor U3432 (N_3432,N_2716,N_2796);
nor U3433 (N_3433,N_2458,N_2468);
or U3434 (N_3434,N_2512,N_2475);
and U3435 (N_3435,N_2727,N_2895);
nor U3436 (N_3436,N_2747,N_2977);
and U3437 (N_3437,N_2952,N_2566);
and U3438 (N_3438,N_2985,N_2572);
xor U3439 (N_3439,N_2849,N_2595);
nor U3440 (N_3440,N_2692,N_2667);
or U3441 (N_3441,N_2943,N_2426);
nor U3442 (N_3442,N_2506,N_2655);
nand U3443 (N_3443,N_2600,N_2496);
nand U3444 (N_3444,N_2706,N_2833);
or U3445 (N_3445,N_2858,N_2692);
xor U3446 (N_3446,N_2612,N_2412);
and U3447 (N_3447,N_2858,N_2733);
xor U3448 (N_3448,N_2835,N_2990);
and U3449 (N_3449,N_2763,N_2559);
nor U3450 (N_3450,N_2409,N_2499);
or U3451 (N_3451,N_2816,N_2740);
xnor U3452 (N_3452,N_2767,N_2504);
nand U3453 (N_3453,N_2735,N_2556);
nand U3454 (N_3454,N_2640,N_2993);
nand U3455 (N_3455,N_2656,N_2684);
nand U3456 (N_3456,N_2736,N_2922);
nor U3457 (N_3457,N_2456,N_2965);
nor U3458 (N_3458,N_2415,N_2480);
and U3459 (N_3459,N_2625,N_2749);
or U3460 (N_3460,N_2892,N_2872);
nand U3461 (N_3461,N_2823,N_2426);
nor U3462 (N_3462,N_2868,N_2894);
nor U3463 (N_3463,N_2455,N_2480);
nand U3464 (N_3464,N_2990,N_2942);
nor U3465 (N_3465,N_2944,N_2892);
or U3466 (N_3466,N_2793,N_2716);
nand U3467 (N_3467,N_2874,N_2453);
nand U3468 (N_3468,N_2743,N_2436);
and U3469 (N_3469,N_2742,N_2514);
and U3470 (N_3470,N_2972,N_2573);
xnor U3471 (N_3471,N_2694,N_2781);
nor U3472 (N_3472,N_2733,N_2424);
and U3473 (N_3473,N_2995,N_2460);
xnor U3474 (N_3474,N_2683,N_2460);
nor U3475 (N_3475,N_2806,N_2881);
xnor U3476 (N_3476,N_2785,N_2685);
or U3477 (N_3477,N_2834,N_2898);
nand U3478 (N_3478,N_2932,N_2540);
nand U3479 (N_3479,N_2980,N_2573);
xnor U3480 (N_3480,N_2842,N_2728);
xor U3481 (N_3481,N_2658,N_2968);
nand U3482 (N_3482,N_2837,N_2998);
xnor U3483 (N_3483,N_2765,N_2641);
and U3484 (N_3484,N_2970,N_2764);
or U3485 (N_3485,N_2836,N_2434);
and U3486 (N_3486,N_2592,N_2723);
nor U3487 (N_3487,N_2567,N_2956);
xnor U3488 (N_3488,N_2475,N_2850);
xor U3489 (N_3489,N_2882,N_2487);
and U3490 (N_3490,N_2645,N_2824);
and U3491 (N_3491,N_2791,N_2604);
nand U3492 (N_3492,N_2641,N_2909);
nor U3493 (N_3493,N_2833,N_2859);
and U3494 (N_3494,N_2749,N_2458);
nand U3495 (N_3495,N_2696,N_2675);
nor U3496 (N_3496,N_2946,N_2858);
or U3497 (N_3497,N_2718,N_2940);
nor U3498 (N_3498,N_2670,N_2644);
nand U3499 (N_3499,N_2453,N_2725);
or U3500 (N_3500,N_2412,N_2773);
nand U3501 (N_3501,N_2659,N_2424);
xor U3502 (N_3502,N_2873,N_2475);
xnor U3503 (N_3503,N_2537,N_2826);
nor U3504 (N_3504,N_2551,N_2468);
and U3505 (N_3505,N_2599,N_2786);
nor U3506 (N_3506,N_2514,N_2621);
nor U3507 (N_3507,N_2574,N_2859);
nand U3508 (N_3508,N_2754,N_2442);
and U3509 (N_3509,N_2548,N_2714);
xnor U3510 (N_3510,N_2796,N_2678);
and U3511 (N_3511,N_2858,N_2490);
or U3512 (N_3512,N_2886,N_2945);
and U3513 (N_3513,N_2576,N_2731);
or U3514 (N_3514,N_2920,N_2620);
xor U3515 (N_3515,N_2518,N_2943);
or U3516 (N_3516,N_2785,N_2626);
or U3517 (N_3517,N_2923,N_2717);
nand U3518 (N_3518,N_2757,N_2543);
xor U3519 (N_3519,N_2758,N_2854);
nand U3520 (N_3520,N_2847,N_2538);
nand U3521 (N_3521,N_2576,N_2950);
nand U3522 (N_3522,N_2422,N_2733);
and U3523 (N_3523,N_2590,N_2906);
xnor U3524 (N_3524,N_2738,N_2773);
nand U3525 (N_3525,N_2446,N_2517);
and U3526 (N_3526,N_2562,N_2895);
xor U3527 (N_3527,N_2936,N_2473);
xor U3528 (N_3528,N_2799,N_2846);
nand U3529 (N_3529,N_2848,N_2746);
nor U3530 (N_3530,N_2626,N_2805);
xor U3531 (N_3531,N_2872,N_2777);
nand U3532 (N_3532,N_2914,N_2686);
xnor U3533 (N_3533,N_2476,N_2599);
xor U3534 (N_3534,N_2782,N_2679);
or U3535 (N_3535,N_2493,N_2972);
and U3536 (N_3536,N_2626,N_2645);
nand U3537 (N_3537,N_2509,N_2977);
and U3538 (N_3538,N_2473,N_2939);
and U3539 (N_3539,N_2995,N_2687);
nand U3540 (N_3540,N_2851,N_2853);
nor U3541 (N_3541,N_2579,N_2682);
xor U3542 (N_3542,N_2452,N_2915);
or U3543 (N_3543,N_2420,N_2556);
nor U3544 (N_3544,N_2649,N_2765);
and U3545 (N_3545,N_2433,N_2590);
or U3546 (N_3546,N_2446,N_2960);
nand U3547 (N_3547,N_2715,N_2517);
nor U3548 (N_3548,N_2861,N_2497);
nand U3549 (N_3549,N_2656,N_2409);
and U3550 (N_3550,N_2695,N_2470);
nor U3551 (N_3551,N_2566,N_2975);
xnor U3552 (N_3552,N_2771,N_2416);
nor U3553 (N_3553,N_2530,N_2735);
nand U3554 (N_3554,N_2500,N_2895);
or U3555 (N_3555,N_2486,N_2682);
or U3556 (N_3556,N_2861,N_2985);
nor U3557 (N_3557,N_2846,N_2471);
or U3558 (N_3558,N_2915,N_2866);
or U3559 (N_3559,N_2635,N_2763);
xor U3560 (N_3560,N_2436,N_2792);
or U3561 (N_3561,N_2784,N_2448);
nand U3562 (N_3562,N_2716,N_2518);
and U3563 (N_3563,N_2527,N_2916);
nand U3564 (N_3564,N_2411,N_2499);
or U3565 (N_3565,N_2448,N_2414);
or U3566 (N_3566,N_2934,N_2483);
xnor U3567 (N_3567,N_2491,N_2671);
or U3568 (N_3568,N_2897,N_2817);
or U3569 (N_3569,N_2420,N_2993);
and U3570 (N_3570,N_2453,N_2522);
nor U3571 (N_3571,N_2495,N_2630);
nor U3572 (N_3572,N_2647,N_2642);
or U3573 (N_3573,N_2951,N_2579);
and U3574 (N_3574,N_2532,N_2504);
or U3575 (N_3575,N_2885,N_2604);
xnor U3576 (N_3576,N_2827,N_2620);
and U3577 (N_3577,N_2490,N_2484);
nand U3578 (N_3578,N_2562,N_2796);
nand U3579 (N_3579,N_2520,N_2862);
xor U3580 (N_3580,N_2887,N_2425);
nand U3581 (N_3581,N_2465,N_2472);
and U3582 (N_3582,N_2531,N_2832);
or U3583 (N_3583,N_2718,N_2948);
nand U3584 (N_3584,N_2892,N_2945);
nand U3585 (N_3585,N_2596,N_2583);
or U3586 (N_3586,N_2920,N_2744);
xor U3587 (N_3587,N_2624,N_2977);
xnor U3588 (N_3588,N_2540,N_2637);
or U3589 (N_3589,N_2824,N_2866);
nor U3590 (N_3590,N_2722,N_2515);
nand U3591 (N_3591,N_2920,N_2803);
nor U3592 (N_3592,N_2683,N_2428);
or U3593 (N_3593,N_2484,N_2486);
xnor U3594 (N_3594,N_2751,N_2986);
xnor U3595 (N_3595,N_2708,N_2553);
nor U3596 (N_3596,N_2421,N_2861);
or U3597 (N_3597,N_2911,N_2826);
xor U3598 (N_3598,N_2867,N_2832);
nor U3599 (N_3599,N_2998,N_2838);
xnor U3600 (N_3600,N_3249,N_3472);
xnor U3601 (N_3601,N_3113,N_3084);
nor U3602 (N_3602,N_3376,N_3117);
nand U3603 (N_3603,N_3594,N_3280);
nand U3604 (N_3604,N_3239,N_3374);
nand U3605 (N_3605,N_3212,N_3359);
and U3606 (N_3606,N_3286,N_3320);
nand U3607 (N_3607,N_3118,N_3322);
nor U3608 (N_3608,N_3290,N_3201);
nand U3609 (N_3609,N_3347,N_3399);
nor U3610 (N_3610,N_3242,N_3105);
xnor U3611 (N_3611,N_3099,N_3206);
xnor U3612 (N_3612,N_3591,N_3450);
and U3613 (N_3613,N_3024,N_3078);
nand U3614 (N_3614,N_3200,N_3298);
nand U3615 (N_3615,N_3190,N_3341);
xnor U3616 (N_3616,N_3203,N_3217);
nor U3617 (N_3617,N_3004,N_3339);
or U3618 (N_3618,N_3303,N_3060);
nor U3619 (N_3619,N_3122,N_3002);
nand U3620 (N_3620,N_3406,N_3052);
nor U3621 (N_3621,N_3037,N_3097);
and U3622 (N_3622,N_3246,N_3046);
and U3623 (N_3623,N_3373,N_3362);
and U3624 (N_3624,N_3034,N_3234);
nor U3625 (N_3625,N_3527,N_3482);
nand U3626 (N_3626,N_3486,N_3545);
nand U3627 (N_3627,N_3447,N_3181);
and U3628 (N_3628,N_3302,N_3152);
or U3629 (N_3629,N_3045,N_3567);
nand U3630 (N_3630,N_3082,N_3225);
nor U3631 (N_3631,N_3599,N_3148);
and U3632 (N_3632,N_3431,N_3142);
nand U3633 (N_3633,N_3469,N_3519);
and U3634 (N_3634,N_3087,N_3276);
nand U3635 (N_3635,N_3238,N_3353);
or U3636 (N_3636,N_3335,N_3029);
xnor U3637 (N_3637,N_3306,N_3252);
xor U3638 (N_3638,N_3005,N_3389);
xnor U3639 (N_3639,N_3429,N_3391);
xor U3640 (N_3640,N_3410,N_3357);
and U3641 (N_3641,N_3497,N_3192);
nand U3642 (N_3642,N_3436,N_3000);
nor U3643 (N_3643,N_3067,N_3479);
and U3644 (N_3644,N_3256,N_3536);
xnor U3645 (N_3645,N_3277,N_3418);
nand U3646 (N_3646,N_3430,N_3316);
nand U3647 (N_3647,N_3090,N_3275);
nor U3648 (N_3648,N_3156,N_3384);
nor U3649 (N_3649,N_3058,N_3125);
xor U3650 (N_3650,N_3270,N_3352);
and U3651 (N_3651,N_3415,N_3035);
xnor U3652 (N_3652,N_3189,N_3305);
and U3653 (N_3653,N_3514,N_3513);
and U3654 (N_3654,N_3226,N_3383);
nor U3655 (N_3655,N_3259,N_3495);
xor U3656 (N_3656,N_3008,N_3501);
or U3657 (N_3657,N_3170,N_3214);
nand U3658 (N_3658,N_3124,N_3313);
nor U3659 (N_3659,N_3108,N_3454);
nand U3660 (N_3660,N_3438,N_3414);
and U3661 (N_3661,N_3131,N_3411);
nand U3662 (N_3662,N_3565,N_3560);
nand U3663 (N_3663,N_3515,N_3315);
nand U3664 (N_3664,N_3292,N_3434);
nand U3665 (N_3665,N_3250,N_3041);
xor U3666 (N_3666,N_3523,N_3452);
nand U3667 (N_3667,N_3107,N_3100);
and U3668 (N_3668,N_3139,N_3461);
xnor U3669 (N_3669,N_3449,N_3375);
nand U3670 (N_3670,N_3123,N_3194);
or U3671 (N_3671,N_3552,N_3476);
or U3672 (N_3672,N_3173,N_3050);
or U3673 (N_3673,N_3548,N_3360);
or U3674 (N_3674,N_3288,N_3312);
xor U3675 (N_3675,N_3219,N_3584);
xor U3676 (N_3676,N_3177,N_3505);
or U3677 (N_3677,N_3392,N_3169);
nor U3678 (N_3678,N_3458,N_3554);
or U3679 (N_3679,N_3178,N_3487);
nand U3680 (N_3680,N_3355,N_3187);
nor U3681 (N_3681,N_3329,N_3585);
and U3682 (N_3682,N_3394,N_3509);
xnor U3683 (N_3683,N_3480,N_3068);
nor U3684 (N_3684,N_3174,N_3106);
nand U3685 (N_3685,N_3039,N_3126);
xor U3686 (N_3686,N_3296,N_3417);
xor U3687 (N_3687,N_3570,N_3420);
nand U3688 (N_3688,N_3525,N_3445);
xnor U3689 (N_3689,N_3295,N_3581);
and U3690 (N_3690,N_3204,N_3247);
and U3691 (N_3691,N_3556,N_3498);
xor U3692 (N_3692,N_3251,N_3018);
and U3693 (N_3693,N_3396,N_3062);
xor U3694 (N_3694,N_3561,N_3568);
nand U3695 (N_3695,N_3346,N_3587);
xnor U3696 (N_3696,N_3307,N_3356);
xor U3697 (N_3697,N_3413,N_3057);
and U3698 (N_3698,N_3530,N_3463);
xnor U3699 (N_3699,N_3390,N_3365);
nor U3700 (N_3700,N_3273,N_3340);
nand U3701 (N_3701,N_3533,N_3440);
xor U3702 (N_3702,N_3492,N_3284);
xor U3703 (N_3703,N_3236,N_3241);
nor U3704 (N_3704,N_3001,N_3317);
and U3705 (N_3705,N_3141,N_3473);
xor U3706 (N_3706,N_3208,N_3150);
or U3707 (N_3707,N_3102,N_3379);
nor U3708 (N_3708,N_3191,N_3063);
or U3709 (N_3709,N_3285,N_3083);
or U3710 (N_3710,N_3167,N_3367);
nor U3711 (N_3711,N_3453,N_3361);
and U3712 (N_3712,N_3274,N_3164);
and U3713 (N_3713,N_3381,N_3222);
and U3714 (N_3714,N_3398,N_3022);
nor U3715 (N_3715,N_3459,N_3425);
nor U3716 (N_3716,N_3428,N_3013);
xor U3717 (N_3717,N_3321,N_3582);
nand U3718 (N_3718,N_3089,N_3311);
nand U3719 (N_3719,N_3475,N_3319);
xor U3720 (N_3720,N_3331,N_3490);
nand U3721 (N_3721,N_3248,N_3223);
nand U3722 (N_3722,N_3211,N_3467);
xnor U3723 (N_3723,N_3103,N_3508);
or U3724 (N_3724,N_3385,N_3104);
nand U3725 (N_3725,N_3526,N_3129);
xnor U3726 (N_3726,N_3507,N_3073);
or U3727 (N_3727,N_3338,N_3551);
xor U3728 (N_3728,N_3363,N_3349);
nand U3729 (N_3729,N_3408,N_3337);
nor U3730 (N_3730,N_3055,N_3220);
or U3731 (N_3731,N_3334,N_3301);
nand U3732 (N_3732,N_3016,N_3184);
and U3733 (N_3733,N_3377,N_3443);
and U3734 (N_3734,N_3229,N_3564);
or U3735 (N_3735,N_3294,N_3095);
nor U3736 (N_3736,N_3109,N_3197);
xor U3737 (N_3737,N_3237,N_3233);
nor U3738 (N_3738,N_3442,N_3477);
and U3739 (N_3739,N_3308,N_3293);
nand U3740 (N_3740,N_3128,N_3589);
nand U3741 (N_3741,N_3370,N_3168);
or U3742 (N_3742,N_3172,N_3465);
or U3743 (N_3743,N_3350,N_3020);
and U3744 (N_3744,N_3166,N_3010);
xnor U3745 (N_3745,N_3146,N_3195);
nor U3746 (N_3746,N_3056,N_3216);
or U3747 (N_3747,N_3502,N_3395);
and U3748 (N_3748,N_3543,N_3091);
nor U3749 (N_3749,N_3528,N_3263);
and U3750 (N_3750,N_3221,N_3224);
nor U3751 (N_3751,N_3028,N_3038);
xnor U3752 (N_3752,N_3419,N_3470);
nor U3753 (N_3753,N_3542,N_3006);
xnor U3754 (N_3754,N_3043,N_3269);
or U3755 (N_3755,N_3145,N_3291);
nor U3756 (N_3756,N_3520,N_3009);
xnor U3757 (N_3757,N_3265,N_3205);
nand U3758 (N_3758,N_3081,N_3439);
nand U3759 (N_3759,N_3119,N_3457);
nor U3760 (N_3760,N_3262,N_3388);
nand U3761 (N_3761,N_3583,N_3299);
nor U3762 (N_3762,N_3474,N_3114);
nand U3763 (N_3763,N_3328,N_3400);
nand U3764 (N_3764,N_3456,N_3553);
nor U3765 (N_3765,N_3512,N_3380);
nor U3766 (N_3766,N_3539,N_3264);
xor U3767 (N_3767,N_3318,N_3555);
or U3768 (N_3768,N_3416,N_3143);
and U3769 (N_3769,N_3017,N_3149);
nor U3770 (N_3770,N_3557,N_3592);
and U3771 (N_3771,N_3510,N_3151);
nor U3772 (N_3772,N_3215,N_3185);
nand U3773 (N_3773,N_3048,N_3232);
nand U3774 (N_3774,N_3244,N_3521);
and U3775 (N_3775,N_3506,N_3213);
or U3776 (N_3776,N_3121,N_3230);
xnor U3777 (N_3777,N_3112,N_3163);
nor U3778 (N_3778,N_3579,N_3279);
xnor U3779 (N_3779,N_3471,N_3516);
nand U3780 (N_3780,N_3324,N_3326);
and U3781 (N_3781,N_3571,N_3441);
xor U3782 (N_3782,N_3176,N_3393);
and U3783 (N_3783,N_3433,N_3444);
and U3784 (N_3784,N_3138,N_3460);
xnor U3785 (N_3785,N_3304,N_3049);
or U3786 (N_3786,N_3210,N_3432);
nor U3787 (N_3787,N_3198,N_3023);
nand U3788 (N_3788,N_3069,N_3488);
and U3789 (N_3789,N_3183,N_3547);
nor U3790 (N_3790,N_3165,N_3562);
and U3791 (N_3791,N_3534,N_3127);
or U3792 (N_3792,N_3254,N_3569);
nor U3793 (N_3793,N_3271,N_3578);
xor U3794 (N_3794,N_3135,N_3071);
xor U3795 (N_3795,N_3021,N_3157);
and U3796 (N_3796,N_3075,N_3300);
nor U3797 (N_3797,N_3409,N_3070);
or U3798 (N_3798,N_3314,N_3209);
nor U3799 (N_3799,N_3161,N_3012);
or U3800 (N_3800,N_3202,N_3094);
xnor U3801 (N_3801,N_3297,N_3231);
and U3802 (N_3802,N_3531,N_3342);
nand U3803 (N_3803,N_3550,N_3407);
xor U3804 (N_3804,N_3524,N_3483);
nand U3805 (N_3805,N_3493,N_3544);
or U3806 (N_3806,N_3330,N_3573);
nor U3807 (N_3807,N_3086,N_3137);
nor U3808 (N_3808,N_3228,N_3132);
and U3809 (N_3809,N_3402,N_3085);
and U3810 (N_3810,N_3448,N_3537);
nand U3811 (N_3811,N_3344,N_3336);
nor U3812 (N_3812,N_3397,N_3014);
and U3813 (N_3813,N_3011,N_3496);
xnor U3814 (N_3814,N_3484,N_3588);
nor U3815 (N_3815,N_3435,N_3278);
nand U3816 (N_3816,N_3255,N_3026);
xnor U3817 (N_3817,N_3115,N_3351);
and U3818 (N_3818,N_3541,N_3160);
or U3819 (N_3819,N_3327,N_3387);
xnor U3820 (N_3820,N_3030,N_3077);
or U3821 (N_3821,N_3261,N_3033);
xnor U3822 (N_3822,N_3503,N_3378);
xor U3823 (N_3823,N_3590,N_3310);
nor U3824 (N_3824,N_3518,N_3386);
nor U3825 (N_3825,N_3093,N_3154);
nand U3826 (N_3826,N_3485,N_3019);
and U3827 (N_3827,N_3283,N_3559);
and U3828 (N_3828,N_3426,N_3500);
or U3829 (N_3829,N_3577,N_3040);
nand U3830 (N_3830,N_3369,N_3575);
or U3831 (N_3831,N_3027,N_3451);
nor U3832 (N_3832,N_3140,N_3481);
nor U3833 (N_3833,N_3382,N_3207);
or U3834 (N_3834,N_3258,N_3598);
xnor U3835 (N_3835,N_3064,N_3281);
and U3836 (N_3836,N_3532,N_3401);
nor U3837 (N_3837,N_3186,N_3044);
nand U3838 (N_3838,N_3287,N_3101);
nand U3839 (N_3839,N_3574,N_3563);
and U3840 (N_3840,N_3180,N_3066);
xnor U3841 (N_3841,N_3535,N_3193);
and U3842 (N_3842,N_3042,N_3343);
or U3843 (N_3843,N_3003,N_3289);
and U3844 (N_3844,N_3348,N_3511);
nand U3845 (N_3845,N_3421,N_3182);
or U3846 (N_3846,N_3455,N_3405);
xor U3847 (N_3847,N_3427,N_3517);
and U3848 (N_3848,N_3134,N_3257);
nand U3849 (N_3849,N_3540,N_3031);
or U3850 (N_3850,N_3345,N_3282);
xor U3851 (N_3851,N_3065,N_3053);
and U3852 (N_3852,N_3412,N_3366);
nand U3853 (N_3853,N_3098,N_3155);
xnor U3854 (N_3854,N_3199,N_3158);
xor U3855 (N_3855,N_3529,N_3175);
nor U3856 (N_3856,N_3147,N_3096);
or U3857 (N_3857,N_3489,N_3404);
and U3858 (N_3858,N_3007,N_3196);
nor U3859 (N_3859,N_3036,N_3032);
nand U3860 (N_3860,N_3245,N_3333);
or U3861 (N_3861,N_3179,N_3253);
and U3862 (N_3862,N_3332,N_3546);
nand U3863 (N_3863,N_3272,N_3136);
xor U3864 (N_3864,N_3054,N_3133);
or U3865 (N_3865,N_3538,N_3424);
nand U3866 (N_3866,N_3153,N_3437);
and U3867 (N_3867,N_3364,N_3522);
nor U3868 (N_3868,N_3323,N_3074);
nor U3869 (N_3869,N_3116,N_3576);
and U3870 (N_3870,N_3171,N_3072);
or U3871 (N_3871,N_3059,N_3499);
nand U3872 (N_3872,N_3235,N_3595);
and U3873 (N_3873,N_3325,N_3130);
or U3874 (N_3874,N_3593,N_3061);
and U3875 (N_3875,N_3243,N_3422);
nand U3876 (N_3876,N_3597,N_3309);
xor U3877 (N_3877,N_3227,N_3025);
nand U3878 (N_3878,N_3466,N_3079);
and U3879 (N_3879,N_3464,N_3110);
or U3880 (N_3880,N_3354,N_3358);
nand U3881 (N_3881,N_3268,N_3368);
and U3882 (N_3882,N_3015,N_3260);
and U3883 (N_3883,N_3423,N_3462);
xnor U3884 (N_3884,N_3468,N_3188);
xnor U3885 (N_3885,N_3159,N_3478);
nand U3886 (N_3886,N_3372,N_3266);
and U3887 (N_3887,N_3076,N_3240);
and U3888 (N_3888,N_3162,N_3111);
nor U3889 (N_3889,N_3051,N_3566);
nor U3890 (N_3890,N_3446,N_3218);
nor U3891 (N_3891,N_3080,N_3267);
and U3892 (N_3892,N_3120,N_3549);
nor U3893 (N_3893,N_3580,N_3494);
xor U3894 (N_3894,N_3572,N_3047);
xnor U3895 (N_3895,N_3558,N_3144);
nand U3896 (N_3896,N_3491,N_3403);
nor U3897 (N_3897,N_3596,N_3504);
and U3898 (N_3898,N_3092,N_3586);
xnor U3899 (N_3899,N_3371,N_3088);
and U3900 (N_3900,N_3192,N_3510);
nand U3901 (N_3901,N_3596,N_3196);
nor U3902 (N_3902,N_3248,N_3546);
or U3903 (N_3903,N_3418,N_3024);
xor U3904 (N_3904,N_3453,N_3494);
nor U3905 (N_3905,N_3439,N_3473);
and U3906 (N_3906,N_3415,N_3370);
nand U3907 (N_3907,N_3121,N_3082);
nand U3908 (N_3908,N_3379,N_3131);
and U3909 (N_3909,N_3219,N_3483);
xor U3910 (N_3910,N_3522,N_3135);
nor U3911 (N_3911,N_3308,N_3288);
xor U3912 (N_3912,N_3064,N_3224);
xor U3913 (N_3913,N_3283,N_3313);
or U3914 (N_3914,N_3040,N_3289);
nor U3915 (N_3915,N_3546,N_3073);
and U3916 (N_3916,N_3071,N_3471);
nand U3917 (N_3917,N_3253,N_3546);
xor U3918 (N_3918,N_3587,N_3195);
nand U3919 (N_3919,N_3503,N_3445);
nand U3920 (N_3920,N_3370,N_3149);
nor U3921 (N_3921,N_3000,N_3525);
nand U3922 (N_3922,N_3203,N_3021);
nor U3923 (N_3923,N_3399,N_3123);
nand U3924 (N_3924,N_3083,N_3398);
nor U3925 (N_3925,N_3420,N_3545);
and U3926 (N_3926,N_3575,N_3440);
or U3927 (N_3927,N_3540,N_3185);
or U3928 (N_3928,N_3063,N_3368);
xor U3929 (N_3929,N_3363,N_3065);
nor U3930 (N_3930,N_3387,N_3172);
or U3931 (N_3931,N_3276,N_3110);
xnor U3932 (N_3932,N_3559,N_3095);
xor U3933 (N_3933,N_3446,N_3398);
xor U3934 (N_3934,N_3538,N_3394);
and U3935 (N_3935,N_3250,N_3428);
and U3936 (N_3936,N_3593,N_3321);
nand U3937 (N_3937,N_3218,N_3430);
nor U3938 (N_3938,N_3232,N_3067);
and U3939 (N_3939,N_3543,N_3226);
and U3940 (N_3940,N_3201,N_3299);
xor U3941 (N_3941,N_3428,N_3073);
nand U3942 (N_3942,N_3101,N_3383);
xor U3943 (N_3943,N_3314,N_3588);
nor U3944 (N_3944,N_3289,N_3564);
or U3945 (N_3945,N_3280,N_3344);
or U3946 (N_3946,N_3512,N_3279);
xnor U3947 (N_3947,N_3345,N_3037);
and U3948 (N_3948,N_3378,N_3045);
or U3949 (N_3949,N_3457,N_3473);
xnor U3950 (N_3950,N_3156,N_3215);
nand U3951 (N_3951,N_3481,N_3006);
xnor U3952 (N_3952,N_3014,N_3044);
xor U3953 (N_3953,N_3407,N_3431);
and U3954 (N_3954,N_3055,N_3045);
xor U3955 (N_3955,N_3349,N_3508);
xor U3956 (N_3956,N_3107,N_3251);
and U3957 (N_3957,N_3101,N_3398);
nand U3958 (N_3958,N_3553,N_3262);
or U3959 (N_3959,N_3183,N_3226);
or U3960 (N_3960,N_3036,N_3250);
or U3961 (N_3961,N_3393,N_3435);
nand U3962 (N_3962,N_3457,N_3326);
nand U3963 (N_3963,N_3024,N_3497);
nand U3964 (N_3964,N_3109,N_3379);
xnor U3965 (N_3965,N_3027,N_3414);
xnor U3966 (N_3966,N_3581,N_3031);
xnor U3967 (N_3967,N_3448,N_3302);
and U3968 (N_3968,N_3450,N_3407);
nand U3969 (N_3969,N_3341,N_3028);
or U3970 (N_3970,N_3304,N_3208);
nand U3971 (N_3971,N_3166,N_3196);
or U3972 (N_3972,N_3244,N_3063);
nor U3973 (N_3973,N_3310,N_3417);
nor U3974 (N_3974,N_3340,N_3380);
or U3975 (N_3975,N_3202,N_3552);
nor U3976 (N_3976,N_3133,N_3161);
and U3977 (N_3977,N_3416,N_3170);
xor U3978 (N_3978,N_3470,N_3499);
nand U3979 (N_3979,N_3469,N_3387);
nor U3980 (N_3980,N_3147,N_3191);
nand U3981 (N_3981,N_3006,N_3291);
nand U3982 (N_3982,N_3536,N_3513);
or U3983 (N_3983,N_3560,N_3506);
or U3984 (N_3984,N_3537,N_3188);
or U3985 (N_3985,N_3520,N_3182);
nand U3986 (N_3986,N_3460,N_3541);
xor U3987 (N_3987,N_3027,N_3171);
nand U3988 (N_3988,N_3014,N_3496);
and U3989 (N_3989,N_3586,N_3099);
nor U3990 (N_3990,N_3458,N_3122);
nor U3991 (N_3991,N_3407,N_3203);
and U3992 (N_3992,N_3408,N_3332);
nor U3993 (N_3993,N_3578,N_3092);
nand U3994 (N_3994,N_3476,N_3211);
xnor U3995 (N_3995,N_3326,N_3262);
xor U3996 (N_3996,N_3489,N_3334);
or U3997 (N_3997,N_3454,N_3152);
nand U3998 (N_3998,N_3027,N_3373);
nor U3999 (N_3999,N_3438,N_3187);
nor U4000 (N_4000,N_3087,N_3008);
nor U4001 (N_4001,N_3470,N_3331);
and U4002 (N_4002,N_3435,N_3262);
xor U4003 (N_4003,N_3046,N_3378);
xnor U4004 (N_4004,N_3155,N_3370);
nor U4005 (N_4005,N_3164,N_3428);
and U4006 (N_4006,N_3161,N_3193);
nor U4007 (N_4007,N_3082,N_3336);
xnor U4008 (N_4008,N_3502,N_3102);
and U4009 (N_4009,N_3338,N_3243);
and U4010 (N_4010,N_3409,N_3574);
or U4011 (N_4011,N_3597,N_3012);
and U4012 (N_4012,N_3294,N_3262);
and U4013 (N_4013,N_3356,N_3206);
xnor U4014 (N_4014,N_3511,N_3476);
nand U4015 (N_4015,N_3554,N_3081);
and U4016 (N_4016,N_3043,N_3338);
nand U4017 (N_4017,N_3231,N_3476);
and U4018 (N_4018,N_3318,N_3526);
nand U4019 (N_4019,N_3237,N_3511);
or U4020 (N_4020,N_3127,N_3291);
and U4021 (N_4021,N_3244,N_3357);
xor U4022 (N_4022,N_3524,N_3225);
nand U4023 (N_4023,N_3120,N_3227);
and U4024 (N_4024,N_3081,N_3489);
and U4025 (N_4025,N_3225,N_3265);
nor U4026 (N_4026,N_3155,N_3293);
nor U4027 (N_4027,N_3309,N_3298);
or U4028 (N_4028,N_3262,N_3083);
or U4029 (N_4029,N_3587,N_3173);
or U4030 (N_4030,N_3509,N_3143);
and U4031 (N_4031,N_3252,N_3338);
or U4032 (N_4032,N_3092,N_3352);
and U4033 (N_4033,N_3224,N_3371);
nand U4034 (N_4034,N_3075,N_3313);
nand U4035 (N_4035,N_3101,N_3480);
nand U4036 (N_4036,N_3237,N_3020);
and U4037 (N_4037,N_3446,N_3552);
xnor U4038 (N_4038,N_3387,N_3023);
nor U4039 (N_4039,N_3541,N_3106);
xnor U4040 (N_4040,N_3145,N_3230);
xor U4041 (N_4041,N_3222,N_3530);
nand U4042 (N_4042,N_3495,N_3401);
or U4043 (N_4043,N_3076,N_3087);
and U4044 (N_4044,N_3377,N_3319);
xnor U4045 (N_4045,N_3445,N_3500);
nand U4046 (N_4046,N_3344,N_3050);
nand U4047 (N_4047,N_3529,N_3440);
nand U4048 (N_4048,N_3020,N_3595);
nand U4049 (N_4049,N_3551,N_3170);
nand U4050 (N_4050,N_3544,N_3215);
or U4051 (N_4051,N_3449,N_3525);
nand U4052 (N_4052,N_3209,N_3436);
nor U4053 (N_4053,N_3320,N_3042);
nor U4054 (N_4054,N_3000,N_3274);
nor U4055 (N_4055,N_3539,N_3536);
xnor U4056 (N_4056,N_3523,N_3580);
and U4057 (N_4057,N_3023,N_3341);
nor U4058 (N_4058,N_3461,N_3269);
and U4059 (N_4059,N_3147,N_3228);
xor U4060 (N_4060,N_3329,N_3265);
nand U4061 (N_4061,N_3188,N_3002);
nand U4062 (N_4062,N_3414,N_3371);
nand U4063 (N_4063,N_3243,N_3362);
nand U4064 (N_4064,N_3438,N_3522);
and U4065 (N_4065,N_3341,N_3323);
xnor U4066 (N_4066,N_3287,N_3081);
or U4067 (N_4067,N_3532,N_3218);
nand U4068 (N_4068,N_3486,N_3583);
nor U4069 (N_4069,N_3111,N_3190);
xnor U4070 (N_4070,N_3326,N_3489);
and U4071 (N_4071,N_3547,N_3094);
and U4072 (N_4072,N_3098,N_3265);
or U4073 (N_4073,N_3455,N_3051);
nand U4074 (N_4074,N_3534,N_3232);
or U4075 (N_4075,N_3231,N_3164);
nor U4076 (N_4076,N_3287,N_3050);
and U4077 (N_4077,N_3138,N_3280);
and U4078 (N_4078,N_3101,N_3410);
and U4079 (N_4079,N_3025,N_3569);
nand U4080 (N_4080,N_3505,N_3070);
or U4081 (N_4081,N_3172,N_3540);
xor U4082 (N_4082,N_3032,N_3509);
and U4083 (N_4083,N_3103,N_3099);
xor U4084 (N_4084,N_3575,N_3309);
nand U4085 (N_4085,N_3305,N_3008);
nand U4086 (N_4086,N_3420,N_3463);
nand U4087 (N_4087,N_3132,N_3113);
nor U4088 (N_4088,N_3490,N_3152);
xnor U4089 (N_4089,N_3506,N_3232);
or U4090 (N_4090,N_3039,N_3505);
and U4091 (N_4091,N_3217,N_3031);
and U4092 (N_4092,N_3581,N_3294);
and U4093 (N_4093,N_3096,N_3422);
or U4094 (N_4094,N_3321,N_3307);
or U4095 (N_4095,N_3485,N_3522);
and U4096 (N_4096,N_3530,N_3415);
nand U4097 (N_4097,N_3095,N_3395);
nor U4098 (N_4098,N_3001,N_3022);
nand U4099 (N_4099,N_3500,N_3324);
or U4100 (N_4100,N_3561,N_3594);
nor U4101 (N_4101,N_3439,N_3551);
nor U4102 (N_4102,N_3007,N_3360);
and U4103 (N_4103,N_3377,N_3102);
or U4104 (N_4104,N_3242,N_3060);
nor U4105 (N_4105,N_3018,N_3215);
nor U4106 (N_4106,N_3271,N_3325);
nand U4107 (N_4107,N_3551,N_3334);
nor U4108 (N_4108,N_3163,N_3529);
xor U4109 (N_4109,N_3127,N_3490);
and U4110 (N_4110,N_3554,N_3465);
xor U4111 (N_4111,N_3049,N_3321);
nor U4112 (N_4112,N_3213,N_3048);
nor U4113 (N_4113,N_3511,N_3543);
or U4114 (N_4114,N_3164,N_3397);
or U4115 (N_4115,N_3308,N_3515);
and U4116 (N_4116,N_3373,N_3590);
xor U4117 (N_4117,N_3140,N_3043);
nor U4118 (N_4118,N_3035,N_3407);
and U4119 (N_4119,N_3592,N_3346);
or U4120 (N_4120,N_3553,N_3321);
xnor U4121 (N_4121,N_3256,N_3315);
nand U4122 (N_4122,N_3211,N_3122);
nor U4123 (N_4123,N_3060,N_3074);
and U4124 (N_4124,N_3478,N_3129);
xnor U4125 (N_4125,N_3547,N_3435);
xor U4126 (N_4126,N_3227,N_3547);
and U4127 (N_4127,N_3028,N_3565);
xor U4128 (N_4128,N_3251,N_3577);
and U4129 (N_4129,N_3346,N_3446);
xor U4130 (N_4130,N_3509,N_3421);
xnor U4131 (N_4131,N_3585,N_3261);
nand U4132 (N_4132,N_3020,N_3579);
xnor U4133 (N_4133,N_3068,N_3430);
and U4134 (N_4134,N_3310,N_3211);
xnor U4135 (N_4135,N_3528,N_3025);
or U4136 (N_4136,N_3260,N_3386);
xor U4137 (N_4137,N_3279,N_3594);
nand U4138 (N_4138,N_3509,N_3109);
and U4139 (N_4139,N_3517,N_3148);
xnor U4140 (N_4140,N_3104,N_3522);
xnor U4141 (N_4141,N_3462,N_3185);
xnor U4142 (N_4142,N_3082,N_3554);
nand U4143 (N_4143,N_3520,N_3262);
nand U4144 (N_4144,N_3549,N_3242);
or U4145 (N_4145,N_3359,N_3032);
nand U4146 (N_4146,N_3180,N_3337);
and U4147 (N_4147,N_3449,N_3258);
and U4148 (N_4148,N_3571,N_3312);
nand U4149 (N_4149,N_3585,N_3450);
xor U4150 (N_4150,N_3542,N_3036);
or U4151 (N_4151,N_3232,N_3524);
nor U4152 (N_4152,N_3405,N_3411);
or U4153 (N_4153,N_3008,N_3240);
or U4154 (N_4154,N_3579,N_3276);
xor U4155 (N_4155,N_3433,N_3243);
and U4156 (N_4156,N_3101,N_3006);
nor U4157 (N_4157,N_3091,N_3454);
nand U4158 (N_4158,N_3497,N_3082);
xnor U4159 (N_4159,N_3153,N_3588);
nor U4160 (N_4160,N_3516,N_3519);
nor U4161 (N_4161,N_3174,N_3042);
and U4162 (N_4162,N_3445,N_3593);
nor U4163 (N_4163,N_3399,N_3390);
or U4164 (N_4164,N_3042,N_3077);
and U4165 (N_4165,N_3006,N_3160);
and U4166 (N_4166,N_3395,N_3194);
nand U4167 (N_4167,N_3108,N_3415);
and U4168 (N_4168,N_3128,N_3046);
and U4169 (N_4169,N_3558,N_3373);
nor U4170 (N_4170,N_3444,N_3100);
and U4171 (N_4171,N_3306,N_3069);
xor U4172 (N_4172,N_3220,N_3027);
and U4173 (N_4173,N_3410,N_3188);
nor U4174 (N_4174,N_3576,N_3018);
nor U4175 (N_4175,N_3057,N_3459);
nor U4176 (N_4176,N_3524,N_3093);
nor U4177 (N_4177,N_3135,N_3164);
nor U4178 (N_4178,N_3198,N_3511);
nor U4179 (N_4179,N_3480,N_3279);
nand U4180 (N_4180,N_3372,N_3366);
xnor U4181 (N_4181,N_3386,N_3394);
xor U4182 (N_4182,N_3508,N_3398);
and U4183 (N_4183,N_3313,N_3387);
nor U4184 (N_4184,N_3185,N_3249);
nor U4185 (N_4185,N_3106,N_3323);
xnor U4186 (N_4186,N_3086,N_3080);
and U4187 (N_4187,N_3173,N_3254);
or U4188 (N_4188,N_3450,N_3348);
xor U4189 (N_4189,N_3078,N_3417);
xnor U4190 (N_4190,N_3115,N_3375);
xnor U4191 (N_4191,N_3285,N_3101);
or U4192 (N_4192,N_3492,N_3092);
nor U4193 (N_4193,N_3013,N_3548);
nor U4194 (N_4194,N_3426,N_3565);
and U4195 (N_4195,N_3112,N_3080);
or U4196 (N_4196,N_3325,N_3040);
nor U4197 (N_4197,N_3095,N_3014);
nand U4198 (N_4198,N_3569,N_3382);
nor U4199 (N_4199,N_3133,N_3542);
nor U4200 (N_4200,N_3992,N_4160);
nor U4201 (N_4201,N_3722,N_3767);
xnor U4202 (N_4202,N_4155,N_3946);
nand U4203 (N_4203,N_3935,N_4126);
or U4204 (N_4204,N_4118,N_3993);
nand U4205 (N_4205,N_3602,N_3976);
or U4206 (N_4206,N_3944,N_3680);
xor U4207 (N_4207,N_3673,N_3912);
or U4208 (N_4208,N_3989,N_3832);
and U4209 (N_4209,N_3970,N_4069);
xnor U4210 (N_4210,N_3711,N_3684);
nand U4211 (N_4211,N_3887,N_4116);
nor U4212 (N_4212,N_3810,N_4052);
nor U4213 (N_4213,N_4059,N_3782);
nor U4214 (N_4214,N_3699,N_3932);
and U4215 (N_4215,N_4089,N_3803);
and U4216 (N_4216,N_3794,N_4033);
xnor U4217 (N_4217,N_3778,N_3623);
xor U4218 (N_4218,N_3888,N_3877);
nor U4219 (N_4219,N_3924,N_3876);
nor U4220 (N_4220,N_4120,N_4065);
xnor U4221 (N_4221,N_4038,N_3900);
and U4222 (N_4222,N_3762,N_3721);
nor U4223 (N_4223,N_4072,N_4097);
nor U4224 (N_4224,N_3713,N_3835);
nand U4225 (N_4225,N_3647,N_3644);
and U4226 (N_4226,N_3859,N_3652);
xnor U4227 (N_4227,N_3954,N_4164);
nand U4228 (N_4228,N_3838,N_4008);
and U4229 (N_4229,N_3689,N_4180);
nor U4230 (N_4230,N_3630,N_3829);
nand U4231 (N_4231,N_3925,N_3981);
nor U4232 (N_4232,N_4087,N_3914);
xnor U4233 (N_4233,N_4077,N_3804);
or U4234 (N_4234,N_3765,N_4098);
nand U4235 (N_4235,N_3671,N_3901);
or U4236 (N_4236,N_3800,N_3708);
nor U4237 (N_4237,N_3885,N_4189);
or U4238 (N_4238,N_3939,N_3682);
or U4239 (N_4239,N_4003,N_4016);
and U4240 (N_4240,N_3625,N_3883);
nand U4241 (N_4241,N_4158,N_4082);
nor U4242 (N_4242,N_3963,N_4144);
nor U4243 (N_4243,N_4057,N_3755);
xnor U4244 (N_4244,N_3716,N_3942);
xnor U4245 (N_4245,N_3606,N_3921);
xnor U4246 (N_4246,N_3817,N_3617);
nor U4247 (N_4247,N_3822,N_3831);
nor U4248 (N_4248,N_3881,N_4056);
nand U4249 (N_4249,N_4110,N_3789);
nand U4250 (N_4250,N_3749,N_4032);
xor U4251 (N_4251,N_3718,N_3637);
or U4252 (N_4252,N_4010,N_3839);
xor U4253 (N_4253,N_4054,N_4058);
nand U4254 (N_4254,N_3643,N_3761);
nand U4255 (N_4255,N_3678,N_3893);
xor U4256 (N_4256,N_3968,N_3626);
nand U4257 (N_4257,N_4109,N_3812);
or U4258 (N_4258,N_3702,N_3784);
xor U4259 (N_4259,N_3601,N_3751);
nor U4260 (N_4260,N_3756,N_3971);
xor U4261 (N_4261,N_3933,N_4140);
xnor U4262 (N_4262,N_3937,N_4063);
nand U4263 (N_4263,N_3801,N_4153);
and U4264 (N_4264,N_3915,N_4129);
and U4265 (N_4265,N_3999,N_4039);
xor U4266 (N_4266,N_3686,N_3654);
nor U4267 (N_4267,N_4002,N_3798);
and U4268 (N_4268,N_4167,N_3697);
and U4269 (N_4269,N_3948,N_4013);
nand U4270 (N_4270,N_4099,N_4161);
and U4271 (N_4271,N_4026,N_4159);
or U4272 (N_4272,N_3880,N_3851);
nor U4273 (N_4273,N_3650,N_4190);
and U4274 (N_4274,N_3622,N_3947);
nand U4275 (N_4275,N_3631,N_3896);
or U4276 (N_4276,N_3850,N_3977);
or U4277 (N_4277,N_3988,N_4157);
or U4278 (N_4278,N_4034,N_3941);
or U4279 (N_4279,N_3905,N_3902);
or U4280 (N_4280,N_4005,N_3764);
and U4281 (N_4281,N_3852,N_3814);
and U4282 (N_4282,N_3653,N_3873);
or U4283 (N_4283,N_4046,N_3683);
and U4284 (N_4284,N_3701,N_3791);
xor U4285 (N_4285,N_3729,N_3827);
xnor U4286 (N_4286,N_4037,N_3982);
nand U4287 (N_4287,N_3891,N_4185);
xnor U4288 (N_4288,N_3869,N_3620);
xnor U4289 (N_4289,N_3909,N_3906);
and U4290 (N_4290,N_3853,N_3928);
nand U4291 (N_4291,N_3821,N_3991);
or U4292 (N_4292,N_3813,N_4136);
or U4293 (N_4293,N_4151,N_4051);
xor U4294 (N_4294,N_3926,N_4044);
xor U4295 (N_4295,N_3709,N_3920);
xor U4296 (N_4296,N_3613,N_4122);
nor U4297 (N_4297,N_3953,N_3943);
nor U4298 (N_4298,N_3776,N_3842);
and U4299 (N_4299,N_3805,N_3670);
or U4300 (N_4300,N_3728,N_4131);
and U4301 (N_4301,N_3823,N_4123);
and U4302 (N_4302,N_3995,N_3820);
nand U4303 (N_4303,N_3641,N_3923);
or U4304 (N_4304,N_4197,N_3994);
xnor U4305 (N_4305,N_4168,N_4095);
xnor U4306 (N_4306,N_4187,N_3679);
or U4307 (N_4307,N_3903,N_3746);
nor U4308 (N_4308,N_3674,N_3719);
xor U4309 (N_4309,N_3770,N_4103);
and U4310 (N_4310,N_3786,N_3632);
xor U4311 (N_4311,N_4143,N_3826);
xor U4312 (N_4312,N_4179,N_3696);
nand U4313 (N_4313,N_4133,N_3676);
xor U4314 (N_4314,N_3837,N_4193);
nor U4315 (N_4315,N_3646,N_4107);
nor U4316 (N_4316,N_3636,N_3700);
or U4317 (N_4317,N_3754,N_3735);
nor U4318 (N_4318,N_4009,N_3750);
nor U4319 (N_4319,N_4012,N_4091);
nor U4320 (N_4320,N_4081,N_4028);
xnor U4321 (N_4321,N_4176,N_3760);
and U4322 (N_4322,N_3655,N_4023);
and U4323 (N_4323,N_3856,N_3930);
xor U4324 (N_4324,N_4076,N_3695);
and U4325 (N_4325,N_3608,N_3816);
and U4326 (N_4326,N_3918,N_3973);
or U4327 (N_4327,N_3845,N_3833);
and U4328 (N_4328,N_3707,N_4006);
nand U4329 (N_4329,N_3607,N_3922);
xor U4330 (N_4330,N_3757,N_3618);
xnor U4331 (N_4331,N_3874,N_3997);
nor U4332 (N_4332,N_3611,N_3766);
nor U4333 (N_4333,N_4111,N_4154);
xnor U4334 (N_4334,N_3895,N_3962);
or U4335 (N_4335,N_3872,N_4178);
xnor U4336 (N_4336,N_3712,N_3899);
nor U4337 (N_4337,N_4093,N_4007);
xor U4338 (N_4338,N_4067,N_4062);
or U4339 (N_4339,N_4086,N_3907);
nand U4340 (N_4340,N_3731,N_3843);
xor U4341 (N_4341,N_4186,N_3938);
xor U4342 (N_4342,N_3854,N_4146);
nor U4343 (N_4343,N_4073,N_4170);
nand U4344 (N_4344,N_4127,N_3894);
or U4345 (N_4345,N_3651,N_3956);
or U4346 (N_4346,N_3819,N_3664);
nand U4347 (N_4347,N_3704,N_3985);
nor U4348 (N_4348,N_3940,N_3871);
nand U4349 (N_4349,N_3665,N_3931);
nor U4350 (N_4350,N_4182,N_3966);
xnor U4351 (N_4351,N_3605,N_3635);
xnor U4352 (N_4352,N_4149,N_4115);
and U4353 (N_4353,N_4106,N_3744);
nor U4354 (N_4354,N_3663,N_4022);
nor U4355 (N_4355,N_4020,N_3736);
and U4356 (N_4356,N_4068,N_3958);
nand U4357 (N_4357,N_4061,N_3908);
xor U4358 (N_4358,N_4050,N_3836);
xor U4359 (N_4359,N_3733,N_3669);
and U4360 (N_4360,N_3807,N_4101);
nor U4361 (N_4361,N_3740,N_3737);
or U4362 (N_4362,N_4198,N_4114);
or U4363 (N_4363,N_3692,N_4045);
and U4364 (N_4364,N_4000,N_3884);
nor U4365 (N_4365,N_3706,N_4192);
nor U4366 (N_4366,N_3793,N_4113);
nor U4367 (N_4367,N_4102,N_3950);
or U4368 (N_4368,N_3965,N_3975);
xor U4369 (N_4369,N_3752,N_3864);
xor U4370 (N_4370,N_4142,N_4196);
nor U4371 (N_4371,N_3828,N_3825);
or U4372 (N_4372,N_3726,N_3867);
xnor U4373 (N_4373,N_4104,N_3727);
nand U4374 (N_4374,N_3629,N_3848);
nand U4375 (N_4375,N_3927,N_3609);
nor U4376 (N_4376,N_3645,N_4150);
and U4377 (N_4377,N_3863,N_3775);
nand U4378 (N_4378,N_4108,N_3818);
nand U4379 (N_4379,N_4017,N_3967);
xor U4380 (N_4380,N_3960,N_3659);
and U4381 (N_4381,N_3681,N_3668);
xnor U4382 (N_4382,N_4079,N_3790);
or U4383 (N_4383,N_3759,N_3772);
nor U4384 (N_4384,N_4169,N_4047);
nand U4385 (N_4385,N_3799,N_3773);
and U4386 (N_4386,N_3639,N_3898);
nand U4387 (N_4387,N_3612,N_4084);
nor U4388 (N_4388,N_4083,N_3844);
nor U4389 (N_4389,N_3690,N_3779);
or U4390 (N_4390,N_3792,N_4191);
and U4391 (N_4391,N_4090,N_4139);
or U4392 (N_4392,N_4064,N_3815);
nor U4393 (N_4393,N_4195,N_3732);
xnor U4394 (N_4394,N_3870,N_3886);
nand U4395 (N_4395,N_3717,N_4134);
or U4396 (N_4396,N_3806,N_3978);
and U4397 (N_4397,N_3763,N_3882);
xor U4398 (N_4398,N_4019,N_3714);
and U4399 (N_4399,N_3972,N_4141);
nand U4400 (N_4400,N_4162,N_3743);
nand U4401 (N_4401,N_3949,N_3802);
nor U4402 (N_4402,N_3667,N_3919);
xor U4403 (N_4403,N_3660,N_3703);
xnor U4404 (N_4404,N_3730,N_4125);
nand U4405 (N_4405,N_3841,N_3642);
xnor U4406 (N_4406,N_4035,N_3725);
xor U4407 (N_4407,N_3878,N_3603);
nand U4408 (N_4408,N_4183,N_3951);
and U4409 (N_4409,N_3990,N_3734);
or U4410 (N_4410,N_3616,N_3768);
nor U4411 (N_4411,N_4030,N_3783);
or U4412 (N_4412,N_3811,N_4055);
or U4413 (N_4413,N_4027,N_4001);
xnor U4414 (N_4414,N_3897,N_3830);
and U4415 (N_4415,N_4117,N_3677);
nor U4416 (N_4416,N_4036,N_4145);
nor U4417 (N_4417,N_3986,N_3662);
xor U4418 (N_4418,N_4060,N_3604);
nand U4419 (N_4419,N_3858,N_4147);
nand U4420 (N_4420,N_4163,N_3742);
xor U4421 (N_4421,N_3748,N_3936);
or U4422 (N_4422,N_4128,N_4014);
nor U4423 (N_4423,N_3889,N_3658);
nand U4424 (N_4424,N_4042,N_3640);
or U4425 (N_4425,N_3771,N_3600);
or U4426 (N_4426,N_3980,N_3614);
or U4427 (N_4427,N_3987,N_3916);
or U4428 (N_4428,N_4024,N_3705);
nand U4429 (N_4429,N_3619,N_3621);
xnor U4430 (N_4430,N_3890,N_3781);
xor U4431 (N_4431,N_3795,N_3657);
and U4432 (N_4432,N_3834,N_3969);
or U4433 (N_4433,N_4041,N_4105);
and U4434 (N_4434,N_3840,N_3846);
nor U4435 (N_4435,N_4124,N_4025);
nand U4436 (N_4436,N_4053,N_3685);
xor U4437 (N_4437,N_3672,N_4175);
and U4438 (N_4438,N_3983,N_3809);
xor U4439 (N_4439,N_4011,N_3862);
or U4440 (N_4440,N_3694,N_3904);
xnor U4441 (N_4441,N_4177,N_3865);
xor U4442 (N_4442,N_3913,N_3929);
xor U4443 (N_4443,N_4166,N_3959);
nor U4444 (N_4444,N_4112,N_4132);
xnor U4445 (N_4445,N_4171,N_3996);
xor U4446 (N_4446,N_3741,N_3747);
nand U4447 (N_4447,N_3847,N_4070);
xor U4448 (N_4448,N_4021,N_4184);
nor U4449 (N_4449,N_4137,N_3688);
nand U4450 (N_4450,N_3788,N_3638);
and U4451 (N_4451,N_3724,N_4181);
xor U4452 (N_4452,N_4119,N_3661);
or U4453 (N_4453,N_4194,N_3753);
xor U4454 (N_4454,N_3780,N_4048);
or U4455 (N_4455,N_4074,N_3610);
or U4456 (N_4456,N_4040,N_3955);
and U4457 (N_4457,N_4152,N_4096);
nand U4458 (N_4458,N_3687,N_3910);
nand U4459 (N_4459,N_3875,N_4004);
xnor U4460 (N_4460,N_4085,N_3720);
and U4461 (N_4461,N_3879,N_3769);
nand U4462 (N_4462,N_3666,N_4156);
nand U4463 (N_4463,N_4043,N_4121);
xor U4464 (N_4464,N_3624,N_3917);
nor U4465 (N_4465,N_4188,N_4199);
xnor U4466 (N_4466,N_3934,N_3745);
and U4467 (N_4467,N_3787,N_3998);
xnor U4468 (N_4468,N_3945,N_4080);
nor U4469 (N_4469,N_4100,N_3952);
xor U4470 (N_4470,N_3868,N_3860);
and U4471 (N_4471,N_3855,N_3698);
nor U4472 (N_4472,N_3615,N_4029);
nor U4473 (N_4473,N_3824,N_3723);
nor U4474 (N_4474,N_3633,N_4138);
nand U4475 (N_4475,N_3964,N_3777);
and U4476 (N_4476,N_4066,N_3785);
xnor U4477 (N_4477,N_4075,N_4092);
nand U4478 (N_4478,N_3957,N_3866);
or U4479 (N_4479,N_3796,N_4172);
or U4480 (N_4480,N_3861,N_4088);
nor U4481 (N_4481,N_3628,N_4174);
or U4482 (N_4482,N_3974,N_3857);
nor U4483 (N_4483,N_3849,N_3984);
xor U4484 (N_4484,N_3691,N_4078);
nand U4485 (N_4485,N_3979,N_3675);
xor U4486 (N_4486,N_3738,N_3892);
or U4487 (N_4487,N_3627,N_4015);
and U4488 (N_4488,N_3758,N_4135);
xnor U4489 (N_4489,N_3961,N_3710);
and U4490 (N_4490,N_4148,N_3656);
or U4491 (N_4491,N_3634,N_3739);
nand U4492 (N_4492,N_4071,N_4049);
nand U4493 (N_4493,N_3648,N_3649);
xor U4494 (N_4494,N_3774,N_4094);
and U4495 (N_4495,N_3911,N_4165);
nor U4496 (N_4496,N_3715,N_4031);
or U4497 (N_4497,N_3693,N_4130);
and U4498 (N_4498,N_3797,N_3808);
or U4499 (N_4499,N_4173,N_4018);
or U4500 (N_4500,N_3786,N_3989);
nand U4501 (N_4501,N_3908,N_3633);
xnor U4502 (N_4502,N_3858,N_3774);
and U4503 (N_4503,N_3803,N_4176);
xor U4504 (N_4504,N_3768,N_3877);
nand U4505 (N_4505,N_4133,N_4151);
or U4506 (N_4506,N_4100,N_3735);
nand U4507 (N_4507,N_3891,N_3928);
nor U4508 (N_4508,N_4129,N_3632);
xor U4509 (N_4509,N_3830,N_3963);
xor U4510 (N_4510,N_3913,N_3937);
nor U4511 (N_4511,N_3718,N_4067);
xnor U4512 (N_4512,N_3982,N_4169);
xor U4513 (N_4513,N_3748,N_3672);
and U4514 (N_4514,N_4022,N_4036);
nor U4515 (N_4515,N_3915,N_3711);
xor U4516 (N_4516,N_3752,N_3724);
and U4517 (N_4517,N_4106,N_3928);
nand U4518 (N_4518,N_3666,N_4189);
or U4519 (N_4519,N_4125,N_4196);
or U4520 (N_4520,N_3747,N_3863);
nor U4521 (N_4521,N_4142,N_4101);
xor U4522 (N_4522,N_3659,N_3800);
xor U4523 (N_4523,N_4006,N_4047);
nor U4524 (N_4524,N_3720,N_3956);
or U4525 (N_4525,N_3778,N_3754);
xnor U4526 (N_4526,N_3657,N_3726);
nor U4527 (N_4527,N_3700,N_3840);
nor U4528 (N_4528,N_3944,N_3866);
nor U4529 (N_4529,N_4168,N_3979);
or U4530 (N_4530,N_3829,N_4192);
nor U4531 (N_4531,N_3636,N_3609);
nand U4532 (N_4532,N_4012,N_3848);
xor U4533 (N_4533,N_4159,N_3680);
and U4534 (N_4534,N_3937,N_3741);
nor U4535 (N_4535,N_4055,N_3620);
and U4536 (N_4536,N_3661,N_4149);
nor U4537 (N_4537,N_4004,N_4094);
nand U4538 (N_4538,N_3778,N_3918);
nor U4539 (N_4539,N_3807,N_3837);
nand U4540 (N_4540,N_3782,N_3796);
xnor U4541 (N_4541,N_4002,N_3663);
xor U4542 (N_4542,N_3966,N_4151);
nor U4543 (N_4543,N_3937,N_4053);
nand U4544 (N_4544,N_3999,N_3987);
and U4545 (N_4545,N_4146,N_3995);
xor U4546 (N_4546,N_3681,N_3896);
xnor U4547 (N_4547,N_3733,N_3995);
nand U4548 (N_4548,N_4074,N_3784);
or U4549 (N_4549,N_4155,N_3626);
nor U4550 (N_4550,N_4165,N_3825);
nand U4551 (N_4551,N_4049,N_3872);
and U4552 (N_4552,N_3680,N_3779);
or U4553 (N_4553,N_3949,N_4176);
and U4554 (N_4554,N_4087,N_4027);
or U4555 (N_4555,N_3903,N_3821);
or U4556 (N_4556,N_4113,N_3949);
and U4557 (N_4557,N_4152,N_4026);
xor U4558 (N_4558,N_3710,N_3683);
nand U4559 (N_4559,N_3952,N_3938);
xnor U4560 (N_4560,N_3720,N_4173);
or U4561 (N_4561,N_3832,N_3606);
and U4562 (N_4562,N_3620,N_3980);
xor U4563 (N_4563,N_3665,N_4086);
and U4564 (N_4564,N_4121,N_3768);
nor U4565 (N_4565,N_3700,N_3923);
or U4566 (N_4566,N_3703,N_4120);
and U4567 (N_4567,N_3798,N_3736);
nor U4568 (N_4568,N_4090,N_3797);
nor U4569 (N_4569,N_3733,N_3991);
and U4570 (N_4570,N_4085,N_3924);
nand U4571 (N_4571,N_4063,N_4105);
nor U4572 (N_4572,N_3801,N_3958);
nand U4573 (N_4573,N_3797,N_4172);
and U4574 (N_4574,N_3841,N_4117);
xor U4575 (N_4575,N_3631,N_3969);
xor U4576 (N_4576,N_3980,N_3833);
or U4577 (N_4577,N_3681,N_4152);
nand U4578 (N_4578,N_3898,N_3672);
and U4579 (N_4579,N_3877,N_3961);
xor U4580 (N_4580,N_3962,N_4058);
or U4581 (N_4581,N_3814,N_3717);
and U4582 (N_4582,N_4164,N_3648);
and U4583 (N_4583,N_4048,N_4194);
or U4584 (N_4584,N_3612,N_4059);
nand U4585 (N_4585,N_3830,N_4169);
xnor U4586 (N_4586,N_3933,N_3773);
or U4587 (N_4587,N_3726,N_3663);
nand U4588 (N_4588,N_4184,N_4055);
nor U4589 (N_4589,N_3837,N_4184);
nand U4590 (N_4590,N_3773,N_3627);
and U4591 (N_4591,N_3749,N_3793);
or U4592 (N_4592,N_4027,N_4144);
nand U4593 (N_4593,N_3835,N_3621);
or U4594 (N_4594,N_3769,N_4113);
or U4595 (N_4595,N_4182,N_3823);
nor U4596 (N_4596,N_3754,N_3895);
and U4597 (N_4597,N_4184,N_4095);
or U4598 (N_4598,N_4076,N_4064);
and U4599 (N_4599,N_4147,N_4189);
xor U4600 (N_4600,N_3799,N_3912);
and U4601 (N_4601,N_4078,N_4011);
nand U4602 (N_4602,N_4149,N_3810);
or U4603 (N_4603,N_4014,N_3741);
or U4604 (N_4604,N_4150,N_3861);
nand U4605 (N_4605,N_3886,N_3619);
xor U4606 (N_4606,N_3818,N_4186);
xnor U4607 (N_4607,N_4175,N_3938);
xnor U4608 (N_4608,N_3995,N_4124);
nor U4609 (N_4609,N_3888,N_4057);
and U4610 (N_4610,N_3638,N_3686);
or U4611 (N_4611,N_4065,N_3963);
xor U4612 (N_4612,N_3891,N_3805);
nor U4613 (N_4613,N_3600,N_3859);
xnor U4614 (N_4614,N_3611,N_3776);
nor U4615 (N_4615,N_3810,N_3654);
xnor U4616 (N_4616,N_3801,N_3763);
or U4617 (N_4617,N_4010,N_3948);
nand U4618 (N_4618,N_3812,N_3705);
nand U4619 (N_4619,N_3868,N_3600);
and U4620 (N_4620,N_4159,N_3854);
or U4621 (N_4621,N_3701,N_4090);
nand U4622 (N_4622,N_4143,N_3790);
nor U4623 (N_4623,N_3691,N_3891);
xnor U4624 (N_4624,N_4016,N_3719);
nand U4625 (N_4625,N_4091,N_3774);
and U4626 (N_4626,N_3670,N_4044);
nor U4627 (N_4627,N_4094,N_4077);
nand U4628 (N_4628,N_4016,N_3972);
nor U4629 (N_4629,N_3729,N_3919);
or U4630 (N_4630,N_3742,N_3644);
nand U4631 (N_4631,N_3634,N_3610);
and U4632 (N_4632,N_4109,N_4055);
xnor U4633 (N_4633,N_3902,N_3785);
or U4634 (N_4634,N_3837,N_4107);
xnor U4635 (N_4635,N_3946,N_4154);
or U4636 (N_4636,N_3960,N_4186);
xnor U4637 (N_4637,N_3724,N_3989);
xnor U4638 (N_4638,N_4197,N_4086);
and U4639 (N_4639,N_3737,N_3715);
nand U4640 (N_4640,N_3990,N_3673);
nor U4641 (N_4641,N_3613,N_3885);
xor U4642 (N_4642,N_3782,N_4026);
and U4643 (N_4643,N_3698,N_3931);
nor U4644 (N_4644,N_3822,N_3801);
and U4645 (N_4645,N_3714,N_4126);
xnor U4646 (N_4646,N_3797,N_4143);
nor U4647 (N_4647,N_4180,N_3674);
nor U4648 (N_4648,N_4127,N_4148);
or U4649 (N_4649,N_3965,N_4127);
nor U4650 (N_4650,N_3991,N_3926);
nand U4651 (N_4651,N_3926,N_3846);
nand U4652 (N_4652,N_3942,N_4196);
nand U4653 (N_4653,N_3982,N_4082);
nand U4654 (N_4654,N_3806,N_3923);
nand U4655 (N_4655,N_3664,N_3974);
xnor U4656 (N_4656,N_4120,N_4064);
nand U4657 (N_4657,N_4163,N_4193);
and U4658 (N_4658,N_4126,N_3826);
or U4659 (N_4659,N_3694,N_3680);
xor U4660 (N_4660,N_3743,N_4025);
or U4661 (N_4661,N_3712,N_3958);
and U4662 (N_4662,N_3856,N_3680);
and U4663 (N_4663,N_3927,N_4125);
or U4664 (N_4664,N_4000,N_3892);
and U4665 (N_4665,N_4061,N_4017);
nand U4666 (N_4666,N_3809,N_4161);
or U4667 (N_4667,N_3860,N_3736);
and U4668 (N_4668,N_3759,N_3696);
or U4669 (N_4669,N_3906,N_3600);
or U4670 (N_4670,N_3944,N_4169);
nor U4671 (N_4671,N_4172,N_3621);
and U4672 (N_4672,N_4151,N_4127);
nand U4673 (N_4673,N_3900,N_3935);
nand U4674 (N_4674,N_4145,N_4198);
nor U4675 (N_4675,N_4195,N_4156);
or U4676 (N_4676,N_3941,N_4059);
and U4677 (N_4677,N_3789,N_3892);
nand U4678 (N_4678,N_3697,N_3636);
nor U4679 (N_4679,N_3789,N_3969);
nand U4680 (N_4680,N_3977,N_4035);
and U4681 (N_4681,N_3964,N_3897);
nor U4682 (N_4682,N_4176,N_4114);
and U4683 (N_4683,N_3959,N_3993);
nor U4684 (N_4684,N_4042,N_3919);
and U4685 (N_4685,N_4128,N_3969);
and U4686 (N_4686,N_4061,N_3666);
and U4687 (N_4687,N_4028,N_3792);
nand U4688 (N_4688,N_4138,N_3843);
nor U4689 (N_4689,N_3860,N_3843);
xor U4690 (N_4690,N_4109,N_4165);
nand U4691 (N_4691,N_4050,N_3839);
or U4692 (N_4692,N_3785,N_3700);
nor U4693 (N_4693,N_3997,N_3828);
and U4694 (N_4694,N_3861,N_3999);
xor U4695 (N_4695,N_4107,N_4154);
nor U4696 (N_4696,N_3610,N_4039);
xor U4697 (N_4697,N_3913,N_3889);
or U4698 (N_4698,N_4087,N_4179);
nor U4699 (N_4699,N_4076,N_3677);
and U4700 (N_4700,N_3626,N_3917);
nor U4701 (N_4701,N_4007,N_3830);
and U4702 (N_4702,N_3827,N_3999);
nor U4703 (N_4703,N_3633,N_3787);
or U4704 (N_4704,N_4059,N_3883);
and U4705 (N_4705,N_3622,N_4062);
nand U4706 (N_4706,N_3642,N_4073);
or U4707 (N_4707,N_4167,N_3619);
nor U4708 (N_4708,N_4095,N_3697);
xor U4709 (N_4709,N_3611,N_4195);
nor U4710 (N_4710,N_4024,N_4107);
nor U4711 (N_4711,N_4011,N_4158);
nand U4712 (N_4712,N_3691,N_3813);
and U4713 (N_4713,N_3807,N_3736);
or U4714 (N_4714,N_3666,N_3645);
xor U4715 (N_4715,N_3980,N_3827);
or U4716 (N_4716,N_3677,N_3970);
and U4717 (N_4717,N_4155,N_3867);
nor U4718 (N_4718,N_3615,N_4079);
xnor U4719 (N_4719,N_4107,N_4195);
or U4720 (N_4720,N_4162,N_3899);
nor U4721 (N_4721,N_4190,N_3968);
or U4722 (N_4722,N_3871,N_3905);
and U4723 (N_4723,N_3799,N_4010);
xnor U4724 (N_4724,N_3771,N_3817);
and U4725 (N_4725,N_3641,N_3693);
xor U4726 (N_4726,N_3817,N_3736);
xor U4727 (N_4727,N_4095,N_4018);
nor U4728 (N_4728,N_3918,N_3744);
and U4729 (N_4729,N_3647,N_4001);
and U4730 (N_4730,N_3603,N_3771);
nand U4731 (N_4731,N_3844,N_3622);
nand U4732 (N_4732,N_3750,N_3766);
nor U4733 (N_4733,N_4018,N_4056);
and U4734 (N_4734,N_3779,N_3934);
nand U4735 (N_4735,N_3684,N_3975);
xor U4736 (N_4736,N_3705,N_4149);
and U4737 (N_4737,N_3653,N_4156);
nand U4738 (N_4738,N_3644,N_3948);
xor U4739 (N_4739,N_3864,N_3773);
nand U4740 (N_4740,N_4069,N_3914);
xnor U4741 (N_4741,N_3739,N_4174);
nor U4742 (N_4742,N_4118,N_4101);
xnor U4743 (N_4743,N_3998,N_3757);
and U4744 (N_4744,N_3907,N_3600);
and U4745 (N_4745,N_3941,N_3875);
nor U4746 (N_4746,N_3893,N_3746);
nand U4747 (N_4747,N_3991,N_3614);
xnor U4748 (N_4748,N_3952,N_3892);
xor U4749 (N_4749,N_4070,N_3863);
xnor U4750 (N_4750,N_3876,N_3803);
xor U4751 (N_4751,N_3894,N_3791);
xnor U4752 (N_4752,N_3724,N_3924);
nor U4753 (N_4753,N_4183,N_3628);
nor U4754 (N_4754,N_3807,N_4167);
nor U4755 (N_4755,N_4074,N_3754);
nand U4756 (N_4756,N_4199,N_4117);
or U4757 (N_4757,N_4025,N_3865);
and U4758 (N_4758,N_3938,N_3783);
nor U4759 (N_4759,N_4135,N_4195);
nand U4760 (N_4760,N_4112,N_3756);
and U4761 (N_4761,N_3996,N_4119);
and U4762 (N_4762,N_4020,N_3732);
nand U4763 (N_4763,N_3722,N_4128);
or U4764 (N_4764,N_4158,N_4081);
xnor U4765 (N_4765,N_4184,N_3884);
xor U4766 (N_4766,N_3734,N_4114);
or U4767 (N_4767,N_3686,N_4049);
nor U4768 (N_4768,N_4122,N_4040);
xor U4769 (N_4769,N_4001,N_3759);
nand U4770 (N_4770,N_3805,N_3702);
xnor U4771 (N_4771,N_3982,N_4049);
nand U4772 (N_4772,N_4108,N_3904);
xor U4773 (N_4773,N_3998,N_3823);
nor U4774 (N_4774,N_3850,N_3990);
nor U4775 (N_4775,N_3886,N_3943);
nor U4776 (N_4776,N_4096,N_3996);
xor U4777 (N_4777,N_4195,N_4040);
or U4778 (N_4778,N_3614,N_4144);
nand U4779 (N_4779,N_3692,N_3816);
nand U4780 (N_4780,N_3842,N_3970);
nor U4781 (N_4781,N_4009,N_3987);
nor U4782 (N_4782,N_4069,N_4098);
nand U4783 (N_4783,N_3970,N_4078);
nor U4784 (N_4784,N_3771,N_3769);
and U4785 (N_4785,N_3959,N_4093);
and U4786 (N_4786,N_3890,N_3790);
nand U4787 (N_4787,N_3977,N_3852);
or U4788 (N_4788,N_3793,N_3769);
nor U4789 (N_4789,N_4053,N_3844);
or U4790 (N_4790,N_4077,N_3841);
nand U4791 (N_4791,N_3856,N_3835);
and U4792 (N_4792,N_4186,N_4157);
or U4793 (N_4793,N_3937,N_3891);
xor U4794 (N_4794,N_3647,N_4075);
and U4795 (N_4795,N_3830,N_3619);
nand U4796 (N_4796,N_3772,N_3600);
nor U4797 (N_4797,N_3765,N_3608);
xor U4798 (N_4798,N_3953,N_3617);
or U4799 (N_4799,N_3783,N_3723);
xor U4800 (N_4800,N_4279,N_4309);
xnor U4801 (N_4801,N_4650,N_4718);
nand U4802 (N_4802,N_4202,N_4621);
xnor U4803 (N_4803,N_4648,N_4504);
nand U4804 (N_4804,N_4401,N_4752);
xnor U4805 (N_4805,N_4280,N_4766);
and U4806 (N_4806,N_4339,N_4210);
and U4807 (N_4807,N_4751,N_4735);
xnor U4808 (N_4808,N_4509,N_4461);
and U4809 (N_4809,N_4653,N_4326);
and U4810 (N_4810,N_4422,N_4585);
nand U4811 (N_4811,N_4741,N_4278);
or U4812 (N_4812,N_4612,N_4328);
or U4813 (N_4813,N_4680,N_4486);
and U4814 (N_4814,N_4216,N_4563);
nand U4815 (N_4815,N_4400,N_4286);
or U4816 (N_4816,N_4255,N_4379);
or U4817 (N_4817,N_4620,N_4626);
xnor U4818 (N_4818,N_4652,N_4430);
or U4819 (N_4819,N_4588,N_4781);
or U4820 (N_4820,N_4685,N_4742);
nor U4821 (N_4821,N_4533,N_4463);
or U4822 (N_4822,N_4224,N_4789);
nor U4823 (N_4823,N_4432,N_4450);
nor U4824 (N_4824,N_4493,N_4262);
xnor U4825 (N_4825,N_4406,N_4731);
and U4826 (N_4826,N_4420,N_4715);
nor U4827 (N_4827,N_4475,N_4234);
and U4828 (N_4828,N_4675,N_4549);
nand U4829 (N_4829,N_4700,N_4543);
or U4830 (N_4830,N_4765,N_4415);
nor U4831 (N_4831,N_4477,N_4634);
or U4832 (N_4832,N_4394,N_4538);
and U4833 (N_4833,N_4215,N_4448);
xor U4834 (N_4834,N_4753,N_4227);
and U4835 (N_4835,N_4343,N_4598);
xor U4836 (N_4836,N_4433,N_4297);
and U4837 (N_4837,N_4602,N_4269);
or U4838 (N_4838,N_4410,N_4305);
or U4839 (N_4839,N_4520,N_4673);
xnor U4840 (N_4840,N_4387,N_4720);
xor U4841 (N_4841,N_4637,N_4694);
nand U4842 (N_4842,N_4405,N_4689);
nor U4843 (N_4843,N_4787,N_4294);
or U4844 (N_4844,N_4638,N_4383);
nor U4845 (N_4845,N_4431,N_4528);
or U4846 (N_4846,N_4225,N_4726);
and U4847 (N_4847,N_4325,N_4606);
nand U4848 (N_4848,N_4214,N_4756);
nand U4849 (N_4849,N_4738,N_4500);
xnor U4850 (N_4850,N_4745,N_4688);
and U4851 (N_4851,N_4311,N_4341);
nor U4852 (N_4852,N_4396,N_4728);
xor U4853 (N_4853,N_4777,N_4594);
nor U4854 (N_4854,N_4284,N_4764);
and U4855 (N_4855,N_4783,N_4390);
nand U4856 (N_4856,N_4784,N_4357);
nand U4857 (N_4857,N_4571,N_4527);
nor U4858 (N_4858,N_4668,N_4270);
nor U4859 (N_4859,N_4623,N_4749);
nand U4860 (N_4860,N_4220,N_4366);
nor U4861 (N_4861,N_4545,N_4393);
nand U4862 (N_4862,N_4265,N_4659);
xor U4863 (N_4863,N_4734,N_4456);
xnor U4864 (N_4864,N_4324,N_4243);
nand U4865 (N_4865,N_4367,N_4320);
and U4866 (N_4866,N_4567,N_4536);
or U4867 (N_4867,N_4636,N_4656);
nand U4868 (N_4868,N_4247,N_4595);
or U4869 (N_4869,N_4544,N_4285);
or U4870 (N_4870,N_4746,N_4701);
and U4871 (N_4871,N_4307,N_4521);
nor U4872 (N_4872,N_4739,N_4678);
nor U4873 (N_4873,N_4798,N_4615);
nand U4874 (N_4874,N_4449,N_4359);
xor U4875 (N_4875,N_4403,N_4258);
xnor U4876 (N_4876,N_4522,N_4407);
nand U4877 (N_4877,N_4773,N_4750);
nand U4878 (N_4878,N_4691,N_4348);
and U4879 (N_4879,N_4427,N_4568);
nor U4880 (N_4880,N_4235,N_4722);
and U4881 (N_4881,N_4645,N_4441);
or U4882 (N_4882,N_4369,N_4736);
or U4883 (N_4883,N_4529,N_4295);
xor U4884 (N_4884,N_4426,N_4221);
nor U4885 (N_4885,N_4290,N_4414);
and U4886 (N_4886,N_4708,N_4622);
or U4887 (N_4887,N_4667,N_4537);
and U4888 (N_4888,N_4345,N_4797);
xor U4889 (N_4889,N_4206,N_4373);
or U4890 (N_4890,N_4336,N_4785);
and U4891 (N_4891,N_4608,N_4245);
or U4892 (N_4892,N_4548,N_4550);
xor U4893 (N_4893,N_4768,N_4240);
nand U4894 (N_4894,N_4368,N_4635);
or U4895 (N_4895,N_4329,N_4213);
nand U4896 (N_4896,N_4729,N_4799);
xnor U4897 (N_4897,N_4593,N_4763);
and U4898 (N_4898,N_4535,N_4464);
xor U4899 (N_4899,N_4758,N_4724);
nand U4900 (N_4900,N_4695,N_4706);
nand U4901 (N_4901,N_4398,N_4259);
or U4902 (N_4902,N_4481,N_4459);
xnor U4903 (N_4903,N_4384,N_4484);
nand U4904 (N_4904,N_4551,N_4266);
xor U4905 (N_4905,N_4570,N_4374);
nor U4906 (N_4906,N_4762,N_4555);
nor U4907 (N_4907,N_4219,N_4346);
xnor U4908 (N_4908,N_4358,N_4488);
and U4909 (N_4909,N_4730,N_4434);
nand U4910 (N_4910,N_4767,N_4302);
or U4911 (N_4911,N_4237,N_4462);
and U4912 (N_4912,N_4238,N_4508);
or U4913 (N_4913,N_4273,N_4375);
xnor U4914 (N_4914,N_4204,N_4596);
and U4915 (N_4915,N_4479,N_4209);
nor U4916 (N_4916,N_4319,N_4289);
xnor U4917 (N_4917,N_4465,N_4246);
or U4918 (N_4918,N_4625,N_4457);
and U4919 (N_4919,N_4447,N_4361);
and U4920 (N_4920,N_4419,N_4487);
or U4921 (N_4921,N_4292,N_4712);
nand U4922 (N_4922,N_4709,N_4669);
xor U4923 (N_4923,N_4452,N_4697);
and U4924 (N_4924,N_4253,N_4228);
xor U4925 (N_4925,N_4574,N_4658);
nand U4926 (N_4926,N_4282,N_4629);
nand U4927 (N_4927,N_4350,N_4200);
or U4928 (N_4928,N_4268,N_4435);
nand U4929 (N_4929,N_4424,N_4304);
and U4930 (N_4930,N_4370,N_4761);
or U4931 (N_4931,N_4378,N_4467);
xnor U4932 (N_4932,N_4710,N_4205);
xnor U4933 (N_4933,N_4381,N_4428);
and U4934 (N_4934,N_4480,N_4364);
xor U4935 (N_4935,N_4413,N_4445);
or U4936 (N_4936,N_4496,N_4315);
nor U4937 (N_4937,N_4317,N_4578);
nand U4938 (N_4938,N_4416,N_4252);
nor U4939 (N_4939,N_4639,N_4561);
nand U4940 (N_4940,N_4316,N_4587);
or U4941 (N_4941,N_4386,N_4231);
xor U4942 (N_4942,N_4296,N_4776);
or U4943 (N_4943,N_4498,N_4542);
nor U4944 (N_4944,N_4573,N_4466);
nand U4945 (N_4945,N_4786,N_4793);
xor U4946 (N_4946,N_4313,N_4349);
nand U4947 (N_4947,N_4331,N_4380);
and U4948 (N_4948,N_4553,N_4288);
and U4949 (N_4949,N_4663,N_4458);
nor U4950 (N_4950,N_4705,N_4468);
or U4951 (N_4951,N_4512,N_4287);
xnor U4952 (N_4952,N_4372,N_4589);
xnor U4953 (N_4953,N_4355,N_4790);
xnor U4954 (N_4954,N_4641,N_4775);
nand U4955 (N_4955,N_4211,N_4795);
nand U4956 (N_4956,N_4444,N_4779);
nand U4957 (N_4957,N_4633,N_4614);
xnor U4958 (N_4958,N_4392,N_4566);
and U4959 (N_4959,N_4356,N_4554);
and U4960 (N_4960,N_4397,N_4769);
nor U4961 (N_4961,N_4671,N_4308);
and U4962 (N_4962,N_4619,N_4597);
and U4963 (N_4963,N_4478,N_4681);
xor U4964 (N_4964,N_4660,N_4770);
or U4965 (N_4965,N_4409,N_4298);
and U4966 (N_4966,N_4476,N_4686);
nand U4967 (N_4967,N_4404,N_4274);
nand U4968 (N_4968,N_4226,N_4333);
nor U4969 (N_4969,N_4399,N_4515);
nand U4970 (N_4970,N_4702,N_4260);
nand U4971 (N_4971,N_4352,N_4283);
and U4972 (N_4972,N_4519,N_4611);
nand U4973 (N_4973,N_4382,N_4291);
or U4974 (N_4974,N_4569,N_4248);
and U4975 (N_4975,N_4312,N_4759);
nor U4976 (N_4976,N_4794,N_4523);
nor U4977 (N_4977,N_4354,N_4510);
xor U4978 (N_4978,N_4744,N_4613);
and U4979 (N_4979,N_4796,N_4684);
nand U4980 (N_4980,N_4251,N_4719);
and U4981 (N_4981,N_4275,N_4539);
xnor U4982 (N_4982,N_4272,N_4417);
nor U4983 (N_4983,N_4203,N_4664);
and U4984 (N_4984,N_4778,N_4644);
and U4985 (N_4985,N_4552,N_4492);
and U4986 (N_4986,N_4471,N_4497);
nand U4987 (N_4987,N_4208,N_4782);
or U4988 (N_4988,N_4474,N_4682);
nor U4989 (N_4989,N_4690,N_4727);
nand U4990 (N_4990,N_4732,N_4717);
and U4991 (N_4991,N_4322,N_4711);
xnor U4992 (N_4992,N_4412,N_4647);
xor U4993 (N_4993,N_4624,N_4342);
or U4994 (N_4994,N_4323,N_4276);
and U4995 (N_4995,N_4757,N_4666);
nor U4996 (N_4996,N_4513,N_4692);
or U4997 (N_4997,N_4217,N_4391);
xnor U4998 (N_4998,N_4580,N_4310);
nand U4999 (N_4999,N_4353,N_4299);
or U5000 (N_5000,N_4229,N_4725);
or U5001 (N_5001,N_4698,N_4618);
and U5002 (N_5002,N_4429,N_4242);
nand U5003 (N_5003,N_4581,N_4610);
or U5004 (N_5004,N_4603,N_4395);
or U5005 (N_5005,N_4438,N_4491);
nand U5006 (N_5006,N_4338,N_4212);
or U5007 (N_5007,N_4687,N_4747);
nand U5008 (N_5008,N_4505,N_4703);
and U5009 (N_5009,N_4628,N_4455);
or U5010 (N_5010,N_4303,N_4483);
or U5011 (N_5011,N_4517,N_4640);
nor U5012 (N_5012,N_4301,N_4774);
nor U5013 (N_5013,N_4408,N_4207);
nor U5014 (N_5014,N_4489,N_4525);
xor U5015 (N_5015,N_4642,N_4627);
nor U5016 (N_5016,N_4446,N_4314);
nand U5017 (N_5017,N_4583,N_4503);
and U5018 (N_5018,N_4534,N_4236);
and U5019 (N_5019,N_4418,N_4733);
and U5020 (N_5020,N_4707,N_4263);
nand U5021 (N_5021,N_4609,N_4559);
or U5022 (N_5022,N_4264,N_4363);
nand U5023 (N_5023,N_4599,N_4340);
nor U5024 (N_5024,N_4791,N_4755);
and U5025 (N_5025,N_4485,N_4201);
nor U5026 (N_5026,N_4531,N_4526);
nor U5027 (N_5027,N_4584,N_4546);
xor U5028 (N_5028,N_4670,N_4389);
nor U5029 (N_5029,N_4677,N_4601);
or U5030 (N_5030,N_4257,N_4655);
xnor U5031 (N_5031,N_4713,N_4532);
or U5032 (N_5032,N_4502,N_4579);
nor U5033 (N_5033,N_4222,N_4524);
nor U5034 (N_5034,N_4743,N_4771);
xnor U5035 (N_5035,N_4335,N_4649);
nor U5036 (N_5036,N_4575,N_4560);
or U5037 (N_5037,N_4607,N_4230);
nor U5038 (N_5038,N_4425,N_4556);
nor U5039 (N_5039,N_4516,N_4239);
or U5040 (N_5040,N_4267,N_4740);
and U5041 (N_5041,N_4494,N_4693);
nor U5042 (N_5042,N_4388,N_4250);
or U5043 (N_5043,N_4439,N_4699);
or U5044 (N_5044,N_4723,N_4646);
and U5045 (N_5045,N_4318,N_4351);
nor U5046 (N_5046,N_4721,N_4617);
and U5047 (N_5047,N_4662,N_4281);
nor U5048 (N_5048,N_4440,N_4792);
and U5049 (N_5049,N_4592,N_4442);
xnor U5050 (N_5050,N_4233,N_4514);
nor U5051 (N_5051,N_4540,N_4218);
or U5052 (N_5052,N_4760,N_4306);
and U5053 (N_5053,N_4518,N_4344);
or U5054 (N_5054,N_4541,N_4605);
nand U5055 (N_5055,N_4632,N_4511);
xnor U5056 (N_5056,N_4557,N_4737);
nor U5057 (N_5057,N_4716,N_4443);
nand U5058 (N_5058,N_4547,N_4437);
nand U5059 (N_5059,N_4436,N_4321);
nor U5060 (N_5060,N_4454,N_4271);
nand U5061 (N_5061,N_4565,N_4347);
nand U5062 (N_5062,N_4254,N_4327);
nand U5063 (N_5063,N_4423,N_4714);
nand U5064 (N_5064,N_4582,N_4261);
and U5065 (N_5065,N_4704,N_4572);
nand U5066 (N_5066,N_4564,N_4754);
nor U5067 (N_5067,N_4577,N_4654);
and U5068 (N_5068,N_4495,N_4600);
nor U5069 (N_5069,N_4469,N_4558);
or U5070 (N_5070,N_4576,N_4360);
nor U5071 (N_5071,N_4453,N_4661);
or U5072 (N_5072,N_4586,N_4371);
nor U5073 (N_5073,N_4672,N_4665);
and U5074 (N_5074,N_4507,N_4402);
nor U5075 (N_5075,N_4332,N_4562);
nand U5076 (N_5076,N_4676,N_4780);
nor U5077 (N_5077,N_4696,N_4385);
nor U5078 (N_5078,N_4683,N_4470);
or U5079 (N_5079,N_4365,N_4772);
nand U5080 (N_5080,N_4482,N_4460);
or U5081 (N_5081,N_4501,N_4490);
and U5082 (N_5082,N_4591,N_4300);
xnor U5083 (N_5083,N_4277,N_4330);
xor U5084 (N_5084,N_4337,N_4376);
nand U5085 (N_5085,N_4377,N_4451);
nand U5086 (N_5086,N_4643,N_4472);
nand U5087 (N_5087,N_4421,N_4657);
nor U5088 (N_5088,N_4232,N_4334);
or U5089 (N_5089,N_4244,N_4499);
nor U5090 (N_5090,N_4473,N_4241);
nor U5091 (N_5091,N_4590,N_4506);
nand U5092 (N_5092,N_4362,N_4616);
nand U5093 (N_5093,N_4530,N_4631);
or U5094 (N_5094,N_4256,N_4411);
nand U5095 (N_5095,N_4679,N_4788);
or U5096 (N_5096,N_4249,N_4223);
xnor U5097 (N_5097,N_4748,N_4604);
and U5098 (N_5098,N_4293,N_4630);
nor U5099 (N_5099,N_4674,N_4651);
xnor U5100 (N_5100,N_4631,N_4541);
xnor U5101 (N_5101,N_4591,N_4214);
nor U5102 (N_5102,N_4785,N_4569);
and U5103 (N_5103,N_4394,N_4717);
xor U5104 (N_5104,N_4474,N_4376);
nand U5105 (N_5105,N_4432,N_4354);
xnor U5106 (N_5106,N_4456,N_4717);
xor U5107 (N_5107,N_4596,N_4484);
or U5108 (N_5108,N_4448,N_4452);
nand U5109 (N_5109,N_4660,N_4488);
nor U5110 (N_5110,N_4588,N_4714);
and U5111 (N_5111,N_4599,N_4715);
nand U5112 (N_5112,N_4350,N_4731);
or U5113 (N_5113,N_4313,N_4307);
nor U5114 (N_5114,N_4688,N_4242);
or U5115 (N_5115,N_4771,N_4796);
nor U5116 (N_5116,N_4520,N_4206);
and U5117 (N_5117,N_4342,N_4766);
nor U5118 (N_5118,N_4647,N_4566);
xor U5119 (N_5119,N_4556,N_4353);
or U5120 (N_5120,N_4488,N_4653);
nand U5121 (N_5121,N_4792,N_4475);
and U5122 (N_5122,N_4743,N_4752);
xor U5123 (N_5123,N_4612,N_4521);
nand U5124 (N_5124,N_4471,N_4677);
or U5125 (N_5125,N_4765,N_4244);
xor U5126 (N_5126,N_4480,N_4319);
xor U5127 (N_5127,N_4772,N_4775);
nand U5128 (N_5128,N_4455,N_4403);
nor U5129 (N_5129,N_4255,N_4665);
xnor U5130 (N_5130,N_4477,N_4799);
nor U5131 (N_5131,N_4445,N_4240);
or U5132 (N_5132,N_4483,N_4357);
xnor U5133 (N_5133,N_4246,N_4790);
or U5134 (N_5134,N_4510,N_4593);
nor U5135 (N_5135,N_4225,N_4341);
nand U5136 (N_5136,N_4694,N_4609);
xor U5137 (N_5137,N_4478,N_4777);
nand U5138 (N_5138,N_4556,N_4215);
and U5139 (N_5139,N_4783,N_4404);
nand U5140 (N_5140,N_4690,N_4787);
and U5141 (N_5141,N_4773,N_4644);
xnor U5142 (N_5142,N_4577,N_4618);
and U5143 (N_5143,N_4640,N_4255);
or U5144 (N_5144,N_4445,N_4516);
nor U5145 (N_5145,N_4433,N_4626);
xnor U5146 (N_5146,N_4479,N_4312);
nand U5147 (N_5147,N_4263,N_4625);
nand U5148 (N_5148,N_4468,N_4216);
nor U5149 (N_5149,N_4304,N_4314);
xnor U5150 (N_5150,N_4496,N_4564);
and U5151 (N_5151,N_4616,N_4435);
nand U5152 (N_5152,N_4327,N_4500);
and U5153 (N_5153,N_4651,N_4724);
nor U5154 (N_5154,N_4211,N_4432);
xnor U5155 (N_5155,N_4420,N_4643);
and U5156 (N_5156,N_4543,N_4237);
and U5157 (N_5157,N_4527,N_4260);
or U5158 (N_5158,N_4315,N_4799);
nor U5159 (N_5159,N_4681,N_4761);
or U5160 (N_5160,N_4402,N_4701);
and U5161 (N_5161,N_4542,N_4283);
xor U5162 (N_5162,N_4680,N_4404);
xnor U5163 (N_5163,N_4755,N_4541);
xor U5164 (N_5164,N_4278,N_4426);
and U5165 (N_5165,N_4675,N_4661);
nor U5166 (N_5166,N_4718,N_4604);
and U5167 (N_5167,N_4292,N_4720);
nor U5168 (N_5168,N_4222,N_4587);
nand U5169 (N_5169,N_4708,N_4661);
nand U5170 (N_5170,N_4678,N_4597);
or U5171 (N_5171,N_4667,N_4787);
nand U5172 (N_5172,N_4748,N_4785);
and U5173 (N_5173,N_4615,N_4355);
xor U5174 (N_5174,N_4701,N_4489);
or U5175 (N_5175,N_4751,N_4295);
nor U5176 (N_5176,N_4435,N_4492);
or U5177 (N_5177,N_4396,N_4549);
and U5178 (N_5178,N_4417,N_4573);
and U5179 (N_5179,N_4659,N_4371);
and U5180 (N_5180,N_4716,N_4266);
nand U5181 (N_5181,N_4659,N_4738);
nor U5182 (N_5182,N_4787,N_4389);
and U5183 (N_5183,N_4424,N_4573);
xnor U5184 (N_5184,N_4780,N_4274);
and U5185 (N_5185,N_4699,N_4504);
xor U5186 (N_5186,N_4792,N_4246);
xnor U5187 (N_5187,N_4521,N_4596);
and U5188 (N_5188,N_4342,N_4353);
nand U5189 (N_5189,N_4533,N_4468);
or U5190 (N_5190,N_4697,N_4207);
or U5191 (N_5191,N_4601,N_4691);
or U5192 (N_5192,N_4595,N_4529);
or U5193 (N_5193,N_4473,N_4644);
and U5194 (N_5194,N_4537,N_4627);
and U5195 (N_5195,N_4593,N_4282);
or U5196 (N_5196,N_4394,N_4248);
or U5197 (N_5197,N_4528,N_4607);
and U5198 (N_5198,N_4526,N_4239);
and U5199 (N_5199,N_4448,N_4648);
nand U5200 (N_5200,N_4482,N_4779);
nand U5201 (N_5201,N_4535,N_4644);
and U5202 (N_5202,N_4783,N_4277);
nand U5203 (N_5203,N_4771,N_4720);
or U5204 (N_5204,N_4504,N_4289);
nand U5205 (N_5205,N_4681,N_4783);
xor U5206 (N_5206,N_4540,N_4272);
nand U5207 (N_5207,N_4251,N_4417);
nor U5208 (N_5208,N_4343,N_4427);
nand U5209 (N_5209,N_4267,N_4289);
nor U5210 (N_5210,N_4266,N_4201);
or U5211 (N_5211,N_4692,N_4724);
nand U5212 (N_5212,N_4333,N_4373);
nand U5213 (N_5213,N_4404,N_4689);
and U5214 (N_5214,N_4754,N_4676);
xnor U5215 (N_5215,N_4578,N_4592);
or U5216 (N_5216,N_4746,N_4616);
nor U5217 (N_5217,N_4662,N_4544);
or U5218 (N_5218,N_4608,N_4267);
nor U5219 (N_5219,N_4796,N_4517);
nor U5220 (N_5220,N_4645,N_4205);
xnor U5221 (N_5221,N_4748,N_4249);
or U5222 (N_5222,N_4522,N_4640);
nand U5223 (N_5223,N_4602,N_4542);
or U5224 (N_5224,N_4290,N_4426);
or U5225 (N_5225,N_4781,N_4210);
nand U5226 (N_5226,N_4261,N_4725);
or U5227 (N_5227,N_4578,N_4292);
xnor U5228 (N_5228,N_4484,N_4752);
xor U5229 (N_5229,N_4414,N_4636);
nand U5230 (N_5230,N_4219,N_4447);
nand U5231 (N_5231,N_4782,N_4452);
or U5232 (N_5232,N_4760,N_4511);
or U5233 (N_5233,N_4643,N_4261);
nand U5234 (N_5234,N_4285,N_4771);
nand U5235 (N_5235,N_4656,N_4513);
and U5236 (N_5236,N_4316,N_4239);
nand U5237 (N_5237,N_4225,N_4314);
or U5238 (N_5238,N_4225,N_4310);
xor U5239 (N_5239,N_4294,N_4313);
nand U5240 (N_5240,N_4361,N_4262);
xor U5241 (N_5241,N_4608,N_4369);
and U5242 (N_5242,N_4202,N_4224);
nand U5243 (N_5243,N_4791,N_4482);
nand U5244 (N_5244,N_4225,N_4604);
xor U5245 (N_5245,N_4336,N_4373);
and U5246 (N_5246,N_4281,N_4384);
xor U5247 (N_5247,N_4438,N_4270);
and U5248 (N_5248,N_4748,N_4275);
and U5249 (N_5249,N_4230,N_4382);
xnor U5250 (N_5250,N_4701,N_4218);
nand U5251 (N_5251,N_4734,N_4588);
or U5252 (N_5252,N_4394,N_4609);
nand U5253 (N_5253,N_4379,N_4294);
xnor U5254 (N_5254,N_4362,N_4757);
xor U5255 (N_5255,N_4600,N_4774);
nand U5256 (N_5256,N_4495,N_4219);
xor U5257 (N_5257,N_4704,N_4787);
xor U5258 (N_5258,N_4265,N_4381);
or U5259 (N_5259,N_4647,N_4619);
or U5260 (N_5260,N_4521,N_4785);
and U5261 (N_5261,N_4646,N_4352);
or U5262 (N_5262,N_4220,N_4431);
and U5263 (N_5263,N_4249,N_4282);
xnor U5264 (N_5264,N_4203,N_4267);
or U5265 (N_5265,N_4201,N_4789);
or U5266 (N_5266,N_4364,N_4388);
or U5267 (N_5267,N_4438,N_4237);
or U5268 (N_5268,N_4212,N_4697);
xnor U5269 (N_5269,N_4337,N_4449);
nand U5270 (N_5270,N_4413,N_4609);
nand U5271 (N_5271,N_4302,N_4563);
xor U5272 (N_5272,N_4486,N_4421);
nor U5273 (N_5273,N_4297,N_4422);
xnor U5274 (N_5274,N_4270,N_4699);
nand U5275 (N_5275,N_4202,N_4397);
nand U5276 (N_5276,N_4624,N_4383);
nor U5277 (N_5277,N_4390,N_4428);
nand U5278 (N_5278,N_4243,N_4380);
and U5279 (N_5279,N_4779,N_4703);
xnor U5280 (N_5280,N_4290,N_4501);
xor U5281 (N_5281,N_4690,N_4219);
nand U5282 (N_5282,N_4279,N_4669);
nor U5283 (N_5283,N_4684,N_4608);
nor U5284 (N_5284,N_4705,N_4335);
nor U5285 (N_5285,N_4748,N_4799);
nand U5286 (N_5286,N_4439,N_4352);
nand U5287 (N_5287,N_4757,N_4780);
nor U5288 (N_5288,N_4752,N_4200);
nand U5289 (N_5289,N_4787,N_4345);
and U5290 (N_5290,N_4629,N_4373);
or U5291 (N_5291,N_4681,N_4685);
xor U5292 (N_5292,N_4249,N_4698);
or U5293 (N_5293,N_4571,N_4602);
and U5294 (N_5294,N_4214,N_4715);
and U5295 (N_5295,N_4242,N_4797);
nor U5296 (N_5296,N_4335,N_4467);
or U5297 (N_5297,N_4448,N_4795);
or U5298 (N_5298,N_4256,N_4429);
or U5299 (N_5299,N_4548,N_4589);
xor U5300 (N_5300,N_4759,N_4265);
or U5301 (N_5301,N_4632,N_4464);
nand U5302 (N_5302,N_4791,N_4685);
xor U5303 (N_5303,N_4487,N_4370);
xor U5304 (N_5304,N_4655,N_4404);
nor U5305 (N_5305,N_4685,N_4339);
and U5306 (N_5306,N_4301,N_4413);
xor U5307 (N_5307,N_4503,N_4337);
xor U5308 (N_5308,N_4788,N_4644);
nor U5309 (N_5309,N_4514,N_4269);
nor U5310 (N_5310,N_4720,N_4390);
or U5311 (N_5311,N_4734,N_4610);
or U5312 (N_5312,N_4784,N_4427);
nand U5313 (N_5313,N_4644,N_4736);
or U5314 (N_5314,N_4724,N_4763);
or U5315 (N_5315,N_4737,N_4499);
and U5316 (N_5316,N_4259,N_4677);
nor U5317 (N_5317,N_4258,N_4777);
nand U5318 (N_5318,N_4457,N_4202);
or U5319 (N_5319,N_4226,N_4774);
nor U5320 (N_5320,N_4400,N_4649);
and U5321 (N_5321,N_4614,N_4242);
or U5322 (N_5322,N_4448,N_4532);
nor U5323 (N_5323,N_4285,N_4237);
nand U5324 (N_5324,N_4715,N_4274);
xor U5325 (N_5325,N_4669,N_4490);
or U5326 (N_5326,N_4723,N_4478);
nand U5327 (N_5327,N_4780,N_4512);
nand U5328 (N_5328,N_4461,N_4587);
and U5329 (N_5329,N_4799,N_4619);
xor U5330 (N_5330,N_4613,N_4722);
nor U5331 (N_5331,N_4711,N_4662);
and U5332 (N_5332,N_4411,N_4651);
nor U5333 (N_5333,N_4381,N_4592);
nor U5334 (N_5334,N_4349,N_4440);
nor U5335 (N_5335,N_4260,N_4567);
nor U5336 (N_5336,N_4708,N_4651);
and U5337 (N_5337,N_4534,N_4417);
nand U5338 (N_5338,N_4661,N_4491);
nor U5339 (N_5339,N_4458,N_4240);
nand U5340 (N_5340,N_4407,N_4630);
or U5341 (N_5341,N_4459,N_4299);
nor U5342 (N_5342,N_4787,N_4768);
xnor U5343 (N_5343,N_4608,N_4510);
nor U5344 (N_5344,N_4263,N_4508);
or U5345 (N_5345,N_4520,N_4562);
nand U5346 (N_5346,N_4237,N_4559);
and U5347 (N_5347,N_4633,N_4455);
xnor U5348 (N_5348,N_4228,N_4464);
and U5349 (N_5349,N_4383,N_4516);
or U5350 (N_5350,N_4791,N_4528);
nor U5351 (N_5351,N_4503,N_4609);
or U5352 (N_5352,N_4707,N_4231);
nor U5353 (N_5353,N_4451,N_4244);
xnor U5354 (N_5354,N_4662,N_4218);
or U5355 (N_5355,N_4598,N_4424);
xor U5356 (N_5356,N_4281,N_4372);
nand U5357 (N_5357,N_4620,N_4444);
nor U5358 (N_5358,N_4331,N_4644);
xnor U5359 (N_5359,N_4546,N_4706);
and U5360 (N_5360,N_4381,N_4602);
nor U5361 (N_5361,N_4575,N_4640);
xor U5362 (N_5362,N_4726,N_4347);
nor U5363 (N_5363,N_4540,N_4365);
nor U5364 (N_5364,N_4484,N_4574);
nor U5365 (N_5365,N_4419,N_4682);
nand U5366 (N_5366,N_4407,N_4378);
or U5367 (N_5367,N_4550,N_4362);
and U5368 (N_5368,N_4709,N_4742);
nand U5369 (N_5369,N_4387,N_4763);
nand U5370 (N_5370,N_4627,N_4625);
nand U5371 (N_5371,N_4432,N_4740);
nand U5372 (N_5372,N_4413,N_4268);
nand U5373 (N_5373,N_4682,N_4486);
and U5374 (N_5374,N_4571,N_4700);
xnor U5375 (N_5375,N_4215,N_4311);
nand U5376 (N_5376,N_4294,N_4364);
or U5377 (N_5377,N_4613,N_4575);
and U5378 (N_5378,N_4748,N_4466);
or U5379 (N_5379,N_4202,N_4483);
nor U5380 (N_5380,N_4495,N_4443);
and U5381 (N_5381,N_4355,N_4391);
nand U5382 (N_5382,N_4211,N_4646);
and U5383 (N_5383,N_4791,N_4660);
nor U5384 (N_5384,N_4652,N_4658);
nand U5385 (N_5385,N_4585,N_4738);
nor U5386 (N_5386,N_4736,N_4625);
or U5387 (N_5387,N_4306,N_4225);
nand U5388 (N_5388,N_4732,N_4378);
nand U5389 (N_5389,N_4566,N_4347);
xnor U5390 (N_5390,N_4269,N_4455);
or U5391 (N_5391,N_4417,N_4569);
nor U5392 (N_5392,N_4282,N_4745);
nand U5393 (N_5393,N_4244,N_4531);
nand U5394 (N_5394,N_4330,N_4761);
or U5395 (N_5395,N_4661,N_4442);
nand U5396 (N_5396,N_4227,N_4358);
xor U5397 (N_5397,N_4464,N_4246);
nor U5398 (N_5398,N_4747,N_4507);
xnor U5399 (N_5399,N_4544,N_4565);
xnor U5400 (N_5400,N_5164,N_5137);
nand U5401 (N_5401,N_4890,N_5303);
and U5402 (N_5402,N_5255,N_5286);
or U5403 (N_5403,N_5041,N_5182);
nor U5404 (N_5404,N_5150,N_5357);
nand U5405 (N_5405,N_4977,N_4997);
or U5406 (N_5406,N_5399,N_4892);
and U5407 (N_5407,N_4947,N_4983);
and U5408 (N_5408,N_5084,N_4802);
xnor U5409 (N_5409,N_4812,N_5094);
nand U5410 (N_5410,N_5344,N_5025);
nor U5411 (N_5411,N_5024,N_4881);
or U5412 (N_5412,N_4882,N_4841);
nor U5413 (N_5413,N_4928,N_5038);
or U5414 (N_5414,N_4984,N_4819);
or U5415 (N_5415,N_5224,N_4808);
or U5416 (N_5416,N_4973,N_5086);
nand U5417 (N_5417,N_5238,N_4945);
nand U5418 (N_5418,N_4969,N_5358);
xor U5419 (N_5419,N_4979,N_4873);
xor U5420 (N_5420,N_4927,N_4909);
nand U5421 (N_5421,N_4889,N_4865);
and U5422 (N_5422,N_4985,N_4807);
or U5423 (N_5423,N_5370,N_5047);
and U5424 (N_5424,N_4870,N_5010);
nand U5425 (N_5425,N_4834,N_5079);
or U5426 (N_5426,N_5222,N_4916);
xor U5427 (N_5427,N_4987,N_5181);
nor U5428 (N_5428,N_5269,N_5193);
nand U5429 (N_5429,N_5307,N_5132);
or U5430 (N_5430,N_5336,N_4906);
nand U5431 (N_5431,N_4915,N_5302);
and U5432 (N_5432,N_4829,N_5191);
nand U5433 (N_5433,N_5005,N_4930);
xor U5434 (N_5434,N_4817,N_5173);
nor U5435 (N_5435,N_5329,N_5020);
or U5436 (N_5436,N_5163,N_5019);
or U5437 (N_5437,N_5346,N_5216);
nor U5438 (N_5438,N_5258,N_5264);
nand U5439 (N_5439,N_5376,N_5184);
xor U5440 (N_5440,N_4815,N_4978);
xor U5441 (N_5441,N_5069,N_5284);
and U5442 (N_5442,N_5312,N_5231);
and U5443 (N_5443,N_4942,N_5070);
nor U5444 (N_5444,N_4920,N_4867);
or U5445 (N_5445,N_4929,N_5085);
nand U5446 (N_5446,N_5138,N_5285);
nand U5447 (N_5447,N_5052,N_5305);
or U5448 (N_5448,N_4963,N_5168);
or U5449 (N_5449,N_5075,N_5165);
nand U5450 (N_5450,N_4883,N_5237);
nand U5451 (N_5451,N_5128,N_5140);
nand U5452 (N_5452,N_5001,N_5213);
or U5453 (N_5453,N_5333,N_5327);
xnor U5454 (N_5454,N_5023,N_5392);
and U5455 (N_5455,N_5338,N_4858);
or U5456 (N_5456,N_5283,N_5246);
and U5457 (N_5457,N_4833,N_4980);
nand U5458 (N_5458,N_5321,N_5372);
and U5459 (N_5459,N_5233,N_5197);
and U5460 (N_5460,N_5162,N_4849);
nand U5461 (N_5461,N_5027,N_4901);
xnor U5462 (N_5462,N_4863,N_4925);
nand U5463 (N_5463,N_5136,N_4908);
and U5464 (N_5464,N_5248,N_5391);
or U5465 (N_5465,N_5190,N_5249);
xnor U5466 (N_5466,N_5202,N_5268);
or U5467 (N_5467,N_5373,N_5330);
xor U5468 (N_5468,N_5118,N_5334);
or U5469 (N_5469,N_4962,N_4917);
and U5470 (N_5470,N_4886,N_5029);
nand U5471 (N_5471,N_4918,N_4827);
and U5472 (N_5472,N_5218,N_5090);
and U5473 (N_5473,N_4838,N_5206);
and U5474 (N_5474,N_4960,N_5187);
or U5475 (N_5475,N_5091,N_5261);
nor U5476 (N_5476,N_5002,N_5033);
xor U5477 (N_5477,N_4888,N_5148);
nor U5478 (N_5478,N_4988,N_4931);
nor U5479 (N_5479,N_5201,N_5272);
xnor U5480 (N_5480,N_4955,N_5217);
nand U5481 (N_5481,N_5214,N_5039);
xor U5482 (N_5482,N_5388,N_5382);
nand U5483 (N_5483,N_5262,N_5080);
nor U5484 (N_5484,N_5100,N_4999);
xnor U5485 (N_5485,N_5227,N_5176);
and U5486 (N_5486,N_4975,N_5104);
nor U5487 (N_5487,N_5098,N_4823);
and U5488 (N_5488,N_5229,N_5082);
nor U5489 (N_5489,N_5050,N_5016);
or U5490 (N_5490,N_4990,N_5095);
and U5491 (N_5491,N_5194,N_4934);
and U5492 (N_5492,N_5320,N_4933);
xor U5493 (N_5493,N_5185,N_5043);
xor U5494 (N_5494,N_5287,N_5223);
nor U5495 (N_5495,N_5351,N_4900);
xnor U5496 (N_5496,N_5092,N_5073);
or U5497 (N_5497,N_5298,N_5053);
xnor U5498 (N_5498,N_5105,N_5278);
or U5499 (N_5499,N_5276,N_5308);
nand U5500 (N_5500,N_4899,N_5282);
nor U5501 (N_5501,N_5143,N_4904);
and U5502 (N_5502,N_5319,N_4828);
nand U5503 (N_5503,N_5241,N_5364);
or U5504 (N_5504,N_5309,N_4830);
nand U5505 (N_5505,N_4831,N_4861);
nand U5506 (N_5506,N_4837,N_4851);
nand U5507 (N_5507,N_4844,N_4958);
nor U5508 (N_5508,N_5365,N_5074);
xor U5509 (N_5509,N_5167,N_5042);
xnor U5510 (N_5510,N_5022,N_5290);
or U5511 (N_5511,N_4832,N_5062);
nor U5512 (N_5512,N_4898,N_4843);
and U5513 (N_5513,N_5247,N_5355);
nor U5514 (N_5514,N_4804,N_4821);
or U5515 (N_5515,N_4891,N_5297);
or U5516 (N_5516,N_5242,N_5048);
nand U5517 (N_5517,N_4913,N_5310);
xnor U5518 (N_5518,N_5109,N_4856);
nor U5519 (N_5519,N_5347,N_5386);
xnor U5520 (N_5520,N_5230,N_5196);
and U5521 (N_5521,N_5076,N_5175);
and U5522 (N_5522,N_5004,N_5266);
nor U5523 (N_5523,N_5125,N_4943);
nand U5524 (N_5524,N_4970,N_5153);
and U5525 (N_5525,N_5063,N_4974);
nor U5526 (N_5526,N_4869,N_4826);
xor U5527 (N_5527,N_4825,N_4910);
nor U5528 (N_5528,N_4806,N_4902);
or U5529 (N_5529,N_5099,N_4941);
nand U5530 (N_5530,N_5198,N_4814);
xnor U5531 (N_5531,N_4952,N_5381);
nor U5532 (N_5532,N_5061,N_5359);
or U5533 (N_5533,N_5055,N_5172);
nand U5534 (N_5534,N_4995,N_5131);
nor U5535 (N_5535,N_5385,N_5263);
nor U5536 (N_5536,N_5383,N_5369);
nor U5537 (N_5537,N_5178,N_5211);
or U5538 (N_5538,N_5316,N_5368);
and U5539 (N_5539,N_5295,N_5339);
and U5540 (N_5540,N_5111,N_4998);
nand U5541 (N_5541,N_4846,N_5127);
or U5542 (N_5542,N_5067,N_5236);
xnor U5543 (N_5543,N_4874,N_5018);
nor U5544 (N_5544,N_5122,N_4848);
xnor U5545 (N_5545,N_5380,N_5256);
nand U5546 (N_5546,N_4946,N_5171);
or U5547 (N_5547,N_5113,N_5395);
nor U5548 (N_5548,N_4961,N_5155);
nand U5549 (N_5549,N_5366,N_4967);
or U5550 (N_5550,N_4938,N_4847);
nor U5551 (N_5551,N_5342,N_4996);
xnor U5552 (N_5552,N_5151,N_5396);
xor U5553 (N_5553,N_4816,N_4923);
xnor U5554 (N_5554,N_5232,N_5126);
xor U5555 (N_5555,N_4852,N_5296);
or U5556 (N_5556,N_4809,N_5013);
or U5557 (N_5557,N_5387,N_5116);
nor U5558 (N_5558,N_4877,N_5301);
and U5559 (N_5559,N_5174,N_4839);
and U5560 (N_5560,N_5253,N_5007);
xor U5561 (N_5561,N_5087,N_5354);
xor U5562 (N_5562,N_5051,N_5186);
or U5563 (N_5563,N_4884,N_5271);
or U5564 (N_5564,N_5081,N_5158);
nor U5565 (N_5565,N_4879,N_5257);
nor U5566 (N_5566,N_5000,N_5345);
or U5567 (N_5567,N_4878,N_5112);
nor U5568 (N_5568,N_5322,N_4949);
and U5569 (N_5569,N_5147,N_5270);
xor U5570 (N_5570,N_5328,N_5349);
xnor U5571 (N_5571,N_5096,N_5183);
nor U5572 (N_5572,N_5362,N_5389);
and U5573 (N_5573,N_4818,N_5350);
or U5574 (N_5574,N_5108,N_4911);
or U5575 (N_5575,N_5259,N_5252);
or U5576 (N_5576,N_5279,N_5315);
or U5577 (N_5577,N_4991,N_4944);
nand U5578 (N_5578,N_5059,N_5011);
and U5579 (N_5579,N_5275,N_5093);
or U5580 (N_5580,N_4803,N_4805);
or U5581 (N_5581,N_5306,N_5244);
nand U5582 (N_5582,N_4859,N_5220);
xnor U5583 (N_5583,N_5277,N_5121);
xnor U5584 (N_5584,N_5142,N_5144);
xor U5585 (N_5585,N_4820,N_5367);
and U5586 (N_5586,N_5037,N_5267);
xnor U5587 (N_5587,N_4914,N_5304);
or U5588 (N_5588,N_4835,N_5245);
or U5589 (N_5589,N_5145,N_4850);
or U5590 (N_5590,N_5021,N_5243);
xor U5591 (N_5591,N_5215,N_5102);
nand U5592 (N_5592,N_5117,N_5146);
xnor U5593 (N_5593,N_4857,N_5293);
and U5594 (N_5594,N_4811,N_5068);
nor U5595 (N_5595,N_5156,N_5032);
and U5596 (N_5596,N_4971,N_4964);
nor U5597 (N_5597,N_4921,N_4871);
nand U5598 (N_5598,N_5377,N_4982);
nand U5599 (N_5599,N_4897,N_5205);
xor U5600 (N_5600,N_5239,N_5049);
xnor U5601 (N_5601,N_5323,N_5265);
and U5602 (N_5602,N_5030,N_5324);
xnor U5603 (N_5603,N_5341,N_5340);
xnor U5604 (N_5604,N_5135,N_5159);
and U5605 (N_5605,N_4959,N_4994);
nand U5606 (N_5606,N_5240,N_4905);
xor U5607 (N_5607,N_5326,N_5129);
and U5608 (N_5608,N_4954,N_4822);
nor U5609 (N_5609,N_4932,N_4924);
xnor U5610 (N_5610,N_5363,N_5189);
or U5611 (N_5611,N_5212,N_5060);
xor U5612 (N_5612,N_5360,N_5228);
nand U5613 (N_5613,N_5393,N_5361);
nor U5614 (N_5614,N_4939,N_5057);
and U5615 (N_5615,N_5120,N_4972);
nand U5616 (N_5616,N_5078,N_5035);
nand U5617 (N_5617,N_5065,N_5300);
nor U5618 (N_5618,N_5169,N_4935);
and U5619 (N_5619,N_5101,N_5331);
nor U5620 (N_5620,N_5210,N_5274);
nand U5621 (N_5621,N_5292,N_4845);
nand U5622 (N_5622,N_5337,N_4922);
and U5623 (N_5623,N_4801,N_4855);
or U5624 (N_5624,N_5335,N_5015);
nand U5625 (N_5625,N_5254,N_5040);
xnor U5626 (N_5626,N_5054,N_4800);
nand U5627 (N_5627,N_4894,N_5260);
nor U5628 (N_5628,N_5179,N_5317);
xnor U5629 (N_5629,N_4862,N_5160);
nand U5630 (N_5630,N_5072,N_4986);
nor U5631 (N_5631,N_5398,N_5012);
and U5632 (N_5632,N_5281,N_4810);
nor U5633 (N_5633,N_4981,N_5152);
xnor U5634 (N_5634,N_5314,N_5234);
or U5635 (N_5635,N_5291,N_4836);
xor U5636 (N_5636,N_5299,N_5115);
and U5637 (N_5637,N_5313,N_5288);
or U5638 (N_5638,N_4864,N_4948);
nand U5639 (N_5639,N_4957,N_5199);
nand U5640 (N_5640,N_4937,N_4893);
or U5641 (N_5641,N_4993,N_5195);
nand U5642 (N_5642,N_5226,N_5353);
nor U5643 (N_5643,N_5371,N_5332);
nor U5644 (N_5644,N_4842,N_4919);
nor U5645 (N_5645,N_5207,N_5235);
and U5646 (N_5646,N_5154,N_4936);
and U5647 (N_5647,N_5008,N_5034);
and U5648 (N_5648,N_5204,N_4840);
and U5649 (N_5649,N_5384,N_5134);
nor U5650 (N_5650,N_5325,N_5044);
and U5651 (N_5651,N_4875,N_4876);
nor U5652 (N_5652,N_5273,N_5046);
or U5653 (N_5653,N_5119,N_5009);
or U5654 (N_5654,N_4885,N_5141);
nor U5655 (N_5655,N_5083,N_4940);
and U5656 (N_5656,N_5106,N_4976);
nor U5657 (N_5657,N_5375,N_5026);
xor U5658 (N_5658,N_5394,N_5103);
nor U5659 (N_5659,N_4950,N_5225);
nand U5660 (N_5660,N_5177,N_4824);
and U5661 (N_5661,N_5378,N_4912);
and U5662 (N_5662,N_4880,N_5056);
and U5663 (N_5663,N_5149,N_5114);
nand U5664 (N_5664,N_4872,N_5157);
nor U5665 (N_5665,N_5251,N_5088);
and U5666 (N_5666,N_5028,N_5110);
nand U5667 (N_5667,N_5180,N_5188);
and U5668 (N_5668,N_5170,N_4896);
nor U5669 (N_5669,N_5123,N_5036);
nor U5670 (N_5670,N_5097,N_4866);
and U5671 (N_5671,N_4853,N_5066);
nand U5672 (N_5672,N_4903,N_5077);
and U5673 (N_5673,N_4895,N_4953);
xor U5674 (N_5674,N_5071,N_5130);
nand U5675 (N_5675,N_5014,N_5250);
nor U5676 (N_5676,N_5139,N_4966);
or U5677 (N_5677,N_5374,N_4965);
or U5678 (N_5678,N_5352,N_4813);
or U5679 (N_5679,N_4887,N_4868);
nand U5680 (N_5680,N_5219,N_5356);
nor U5681 (N_5681,N_4968,N_4951);
xor U5682 (N_5682,N_5318,N_5208);
nand U5683 (N_5683,N_5280,N_5200);
nor U5684 (N_5684,N_5133,N_5031);
nand U5685 (N_5685,N_5397,N_5064);
nand U5686 (N_5686,N_4989,N_5006);
nor U5687 (N_5687,N_5124,N_5003);
nand U5688 (N_5688,N_5192,N_5089);
nor U5689 (N_5689,N_4907,N_5045);
and U5690 (N_5690,N_5058,N_5166);
or U5691 (N_5691,N_5294,N_4860);
nor U5692 (N_5692,N_5161,N_5289);
or U5693 (N_5693,N_5379,N_5343);
nor U5694 (N_5694,N_4956,N_5107);
nand U5695 (N_5695,N_5311,N_4854);
nand U5696 (N_5696,N_5390,N_4992);
and U5697 (N_5697,N_5221,N_5203);
or U5698 (N_5698,N_5348,N_5017);
and U5699 (N_5699,N_4926,N_5209);
xnor U5700 (N_5700,N_4874,N_5342);
or U5701 (N_5701,N_4941,N_5109);
or U5702 (N_5702,N_5143,N_5197);
xor U5703 (N_5703,N_5298,N_5363);
nor U5704 (N_5704,N_5093,N_4825);
xor U5705 (N_5705,N_5041,N_5263);
and U5706 (N_5706,N_5181,N_5365);
or U5707 (N_5707,N_4906,N_4918);
xor U5708 (N_5708,N_4880,N_5321);
and U5709 (N_5709,N_4878,N_5305);
nand U5710 (N_5710,N_5067,N_5202);
or U5711 (N_5711,N_5391,N_5179);
nand U5712 (N_5712,N_4826,N_5054);
nand U5713 (N_5713,N_5368,N_5204);
and U5714 (N_5714,N_5251,N_4861);
nor U5715 (N_5715,N_5377,N_5001);
nor U5716 (N_5716,N_5362,N_4879);
xnor U5717 (N_5717,N_4932,N_5258);
nor U5718 (N_5718,N_4812,N_4989);
and U5719 (N_5719,N_4926,N_4974);
nor U5720 (N_5720,N_5287,N_5332);
nand U5721 (N_5721,N_5165,N_4883);
and U5722 (N_5722,N_5055,N_5284);
nor U5723 (N_5723,N_5034,N_5012);
nor U5724 (N_5724,N_5328,N_5322);
and U5725 (N_5725,N_5056,N_5102);
nand U5726 (N_5726,N_5341,N_5257);
nor U5727 (N_5727,N_5004,N_5391);
nand U5728 (N_5728,N_5387,N_4874);
nand U5729 (N_5729,N_4850,N_5169);
nor U5730 (N_5730,N_5019,N_5198);
or U5731 (N_5731,N_4838,N_4887);
or U5732 (N_5732,N_5001,N_4964);
and U5733 (N_5733,N_5246,N_4806);
nor U5734 (N_5734,N_5078,N_4911);
nand U5735 (N_5735,N_4835,N_4841);
nand U5736 (N_5736,N_4816,N_5010);
or U5737 (N_5737,N_5027,N_5165);
and U5738 (N_5738,N_5380,N_5385);
and U5739 (N_5739,N_5359,N_4881);
or U5740 (N_5740,N_5077,N_5226);
and U5741 (N_5741,N_4988,N_5331);
nor U5742 (N_5742,N_4976,N_5205);
xor U5743 (N_5743,N_4972,N_5246);
xor U5744 (N_5744,N_5106,N_5141);
or U5745 (N_5745,N_4876,N_5058);
or U5746 (N_5746,N_5333,N_5375);
nand U5747 (N_5747,N_4806,N_4803);
xnor U5748 (N_5748,N_4994,N_5054);
or U5749 (N_5749,N_5180,N_5121);
nor U5750 (N_5750,N_5227,N_5335);
xnor U5751 (N_5751,N_4968,N_4833);
nor U5752 (N_5752,N_4817,N_5205);
nor U5753 (N_5753,N_4983,N_4878);
and U5754 (N_5754,N_4909,N_5397);
nor U5755 (N_5755,N_4947,N_5301);
and U5756 (N_5756,N_5161,N_5230);
or U5757 (N_5757,N_4847,N_4851);
and U5758 (N_5758,N_5139,N_5262);
or U5759 (N_5759,N_4845,N_5040);
or U5760 (N_5760,N_4906,N_5236);
or U5761 (N_5761,N_5030,N_5202);
or U5762 (N_5762,N_4818,N_5222);
and U5763 (N_5763,N_5375,N_5264);
or U5764 (N_5764,N_4985,N_5053);
xor U5765 (N_5765,N_5285,N_5286);
and U5766 (N_5766,N_5145,N_5092);
xnor U5767 (N_5767,N_5119,N_5262);
nand U5768 (N_5768,N_5274,N_5341);
nor U5769 (N_5769,N_4971,N_5083);
xor U5770 (N_5770,N_5295,N_5228);
nand U5771 (N_5771,N_5256,N_5103);
xnor U5772 (N_5772,N_5299,N_5001);
xor U5773 (N_5773,N_5173,N_5147);
nor U5774 (N_5774,N_4809,N_5226);
or U5775 (N_5775,N_5116,N_5179);
and U5776 (N_5776,N_5252,N_5018);
nor U5777 (N_5777,N_4802,N_4845);
and U5778 (N_5778,N_4949,N_5126);
or U5779 (N_5779,N_5334,N_5360);
nor U5780 (N_5780,N_4916,N_5074);
or U5781 (N_5781,N_4868,N_5322);
or U5782 (N_5782,N_5303,N_4872);
and U5783 (N_5783,N_4839,N_5242);
xor U5784 (N_5784,N_5014,N_5055);
nand U5785 (N_5785,N_4885,N_4883);
and U5786 (N_5786,N_5345,N_5246);
and U5787 (N_5787,N_5156,N_4952);
nand U5788 (N_5788,N_5349,N_5306);
xor U5789 (N_5789,N_5009,N_5300);
xnor U5790 (N_5790,N_4816,N_5171);
nor U5791 (N_5791,N_5318,N_5091);
xor U5792 (N_5792,N_5239,N_5127);
or U5793 (N_5793,N_5291,N_4828);
or U5794 (N_5794,N_5036,N_5276);
xnor U5795 (N_5795,N_5006,N_5165);
nor U5796 (N_5796,N_4913,N_5091);
or U5797 (N_5797,N_5359,N_4901);
nor U5798 (N_5798,N_4998,N_5135);
or U5799 (N_5799,N_5276,N_5110);
or U5800 (N_5800,N_4800,N_5258);
nor U5801 (N_5801,N_5117,N_5113);
or U5802 (N_5802,N_5305,N_5357);
nor U5803 (N_5803,N_5098,N_5167);
and U5804 (N_5804,N_5249,N_4948);
nand U5805 (N_5805,N_5019,N_5099);
or U5806 (N_5806,N_4840,N_4916);
nor U5807 (N_5807,N_5234,N_5170);
and U5808 (N_5808,N_4895,N_5264);
nand U5809 (N_5809,N_5228,N_5282);
xor U5810 (N_5810,N_4988,N_4830);
xnor U5811 (N_5811,N_5017,N_5371);
nor U5812 (N_5812,N_4949,N_5275);
nor U5813 (N_5813,N_5087,N_4983);
and U5814 (N_5814,N_4955,N_4978);
nor U5815 (N_5815,N_5243,N_4844);
nor U5816 (N_5816,N_5348,N_5102);
xor U5817 (N_5817,N_5384,N_4863);
nor U5818 (N_5818,N_5250,N_5237);
nor U5819 (N_5819,N_4826,N_5208);
nor U5820 (N_5820,N_4809,N_4986);
nand U5821 (N_5821,N_4821,N_5354);
and U5822 (N_5822,N_5355,N_5269);
nor U5823 (N_5823,N_5367,N_5119);
or U5824 (N_5824,N_4808,N_4976);
or U5825 (N_5825,N_5340,N_5280);
nor U5826 (N_5826,N_4978,N_5218);
or U5827 (N_5827,N_4837,N_4932);
nor U5828 (N_5828,N_4960,N_5282);
and U5829 (N_5829,N_5085,N_4802);
nand U5830 (N_5830,N_5124,N_5055);
nand U5831 (N_5831,N_5227,N_5368);
nor U5832 (N_5832,N_5268,N_5212);
nand U5833 (N_5833,N_5065,N_5136);
nor U5834 (N_5834,N_4903,N_5299);
nor U5835 (N_5835,N_5338,N_5187);
nor U5836 (N_5836,N_4828,N_5052);
or U5837 (N_5837,N_5249,N_5377);
or U5838 (N_5838,N_4904,N_4971);
nand U5839 (N_5839,N_5104,N_5248);
nor U5840 (N_5840,N_5355,N_5315);
nor U5841 (N_5841,N_5152,N_5014);
xnor U5842 (N_5842,N_4866,N_5081);
and U5843 (N_5843,N_4974,N_5025);
and U5844 (N_5844,N_5369,N_4817);
xnor U5845 (N_5845,N_5136,N_5070);
nor U5846 (N_5846,N_5240,N_4890);
or U5847 (N_5847,N_5173,N_5010);
nor U5848 (N_5848,N_5363,N_4885);
xnor U5849 (N_5849,N_5245,N_5014);
nor U5850 (N_5850,N_4998,N_5040);
nor U5851 (N_5851,N_5114,N_5069);
and U5852 (N_5852,N_4918,N_5128);
or U5853 (N_5853,N_5270,N_5018);
nor U5854 (N_5854,N_5203,N_5199);
or U5855 (N_5855,N_5359,N_5069);
nor U5856 (N_5856,N_4837,N_5250);
nand U5857 (N_5857,N_5228,N_5141);
xnor U5858 (N_5858,N_5022,N_5138);
or U5859 (N_5859,N_5237,N_4981);
nand U5860 (N_5860,N_5305,N_5200);
nor U5861 (N_5861,N_5182,N_5019);
nor U5862 (N_5862,N_4975,N_5256);
xnor U5863 (N_5863,N_5158,N_5146);
or U5864 (N_5864,N_4946,N_4950);
and U5865 (N_5865,N_4902,N_4979);
nor U5866 (N_5866,N_4946,N_5324);
or U5867 (N_5867,N_4830,N_4845);
nor U5868 (N_5868,N_5030,N_4842);
xor U5869 (N_5869,N_4999,N_5342);
or U5870 (N_5870,N_5200,N_5050);
or U5871 (N_5871,N_5283,N_4817);
or U5872 (N_5872,N_5281,N_5137);
or U5873 (N_5873,N_5050,N_5240);
or U5874 (N_5874,N_4805,N_4821);
and U5875 (N_5875,N_5262,N_5315);
nor U5876 (N_5876,N_5058,N_5349);
nand U5877 (N_5877,N_4986,N_4893);
xor U5878 (N_5878,N_5150,N_5385);
and U5879 (N_5879,N_5254,N_4800);
xor U5880 (N_5880,N_5308,N_4997);
or U5881 (N_5881,N_4857,N_5315);
nor U5882 (N_5882,N_5135,N_5072);
or U5883 (N_5883,N_4985,N_5159);
and U5884 (N_5884,N_4819,N_5281);
or U5885 (N_5885,N_5174,N_5071);
or U5886 (N_5886,N_5328,N_5286);
or U5887 (N_5887,N_5291,N_5313);
or U5888 (N_5888,N_5077,N_4824);
xnor U5889 (N_5889,N_5288,N_5207);
and U5890 (N_5890,N_4920,N_4925);
nor U5891 (N_5891,N_4977,N_5113);
and U5892 (N_5892,N_5315,N_4850);
nor U5893 (N_5893,N_4877,N_5376);
nand U5894 (N_5894,N_4944,N_5152);
nor U5895 (N_5895,N_5097,N_5059);
and U5896 (N_5896,N_5362,N_4885);
and U5897 (N_5897,N_5328,N_5316);
nand U5898 (N_5898,N_5305,N_5100);
nand U5899 (N_5899,N_5014,N_5101);
or U5900 (N_5900,N_4920,N_5267);
or U5901 (N_5901,N_5001,N_5310);
nor U5902 (N_5902,N_5207,N_4810);
or U5903 (N_5903,N_4929,N_5357);
xor U5904 (N_5904,N_5305,N_5067);
nor U5905 (N_5905,N_5189,N_4802);
nor U5906 (N_5906,N_5256,N_4820);
or U5907 (N_5907,N_5321,N_4824);
nand U5908 (N_5908,N_5344,N_5292);
nand U5909 (N_5909,N_5179,N_4800);
xnor U5910 (N_5910,N_4950,N_4884);
or U5911 (N_5911,N_4924,N_5343);
nand U5912 (N_5912,N_5269,N_4860);
or U5913 (N_5913,N_4863,N_4902);
and U5914 (N_5914,N_4945,N_5289);
xnor U5915 (N_5915,N_5221,N_5202);
xnor U5916 (N_5916,N_5156,N_5142);
and U5917 (N_5917,N_5009,N_5187);
nor U5918 (N_5918,N_5308,N_4986);
or U5919 (N_5919,N_5131,N_5091);
and U5920 (N_5920,N_5336,N_4975);
and U5921 (N_5921,N_5062,N_5115);
nand U5922 (N_5922,N_4997,N_5236);
or U5923 (N_5923,N_4965,N_4845);
nand U5924 (N_5924,N_4919,N_5205);
nor U5925 (N_5925,N_5272,N_4842);
or U5926 (N_5926,N_4827,N_4962);
or U5927 (N_5927,N_4952,N_4884);
and U5928 (N_5928,N_5223,N_4803);
nor U5929 (N_5929,N_5347,N_4980);
and U5930 (N_5930,N_5367,N_5007);
nand U5931 (N_5931,N_4963,N_5005);
nand U5932 (N_5932,N_5116,N_5046);
xor U5933 (N_5933,N_5012,N_5294);
nand U5934 (N_5934,N_5214,N_5383);
or U5935 (N_5935,N_5159,N_5371);
nor U5936 (N_5936,N_5336,N_5348);
and U5937 (N_5937,N_5113,N_4939);
or U5938 (N_5938,N_4995,N_4926);
nor U5939 (N_5939,N_5104,N_4990);
or U5940 (N_5940,N_5295,N_5112);
or U5941 (N_5941,N_5043,N_5351);
nor U5942 (N_5942,N_5172,N_4954);
and U5943 (N_5943,N_5204,N_5105);
or U5944 (N_5944,N_5248,N_4933);
nor U5945 (N_5945,N_5318,N_4887);
or U5946 (N_5946,N_4925,N_5160);
and U5947 (N_5947,N_4801,N_4923);
nand U5948 (N_5948,N_5396,N_5010);
xor U5949 (N_5949,N_5363,N_5260);
or U5950 (N_5950,N_5081,N_5345);
or U5951 (N_5951,N_5165,N_4814);
or U5952 (N_5952,N_4916,N_5138);
nand U5953 (N_5953,N_5312,N_4902);
xnor U5954 (N_5954,N_5220,N_5236);
nor U5955 (N_5955,N_5171,N_5243);
nand U5956 (N_5956,N_5050,N_5241);
nor U5957 (N_5957,N_4926,N_5255);
and U5958 (N_5958,N_4906,N_5269);
or U5959 (N_5959,N_5374,N_5179);
nand U5960 (N_5960,N_5212,N_5084);
and U5961 (N_5961,N_5303,N_5123);
and U5962 (N_5962,N_4922,N_4866);
or U5963 (N_5963,N_5258,N_5004);
or U5964 (N_5964,N_4891,N_5304);
or U5965 (N_5965,N_5243,N_4826);
and U5966 (N_5966,N_4889,N_4883);
nand U5967 (N_5967,N_5178,N_4873);
nor U5968 (N_5968,N_4987,N_5287);
and U5969 (N_5969,N_4858,N_5025);
or U5970 (N_5970,N_5070,N_4827);
nand U5971 (N_5971,N_5119,N_5079);
or U5972 (N_5972,N_4984,N_5221);
or U5973 (N_5973,N_5211,N_4908);
nor U5974 (N_5974,N_5133,N_5282);
xnor U5975 (N_5975,N_5157,N_4963);
xnor U5976 (N_5976,N_4999,N_5366);
and U5977 (N_5977,N_5264,N_5149);
nand U5978 (N_5978,N_4825,N_5142);
or U5979 (N_5979,N_5063,N_5150);
xor U5980 (N_5980,N_5108,N_5046);
and U5981 (N_5981,N_4963,N_5001);
and U5982 (N_5982,N_5292,N_5374);
nor U5983 (N_5983,N_4824,N_4863);
or U5984 (N_5984,N_5156,N_4998);
nand U5985 (N_5985,N_5212,N_5047);
xnor U5986 (N_5986,N_5034,N_5030);
and U5987 (N_5987,N_5065,N_4866);
nand U5988 (N_5988,N_4855,N_5008);
and U5989 (N_5989,N_5038,N_5138);
or U5990 (N_5990,N_4921,N_5328);
and U5991 (N_5991,N_5182,N_5275);
nor U5992 (N_5992,N_4990,N_4865);
or U5993 (N_5993,N_5391,N_4979);
nand U5994 (N_5994,N_5141,N_4968);
nor U5995 (N_5995,N_5299,N_5005);
or U5996 (N_5996,N_5181,N_4913);
and U5997 (N_5997,N_5021,N_5304);
xnor U5998 (N_5998,N_5148,N_4902);
and U5999 (N_5999,N_4807,N_5365);
xor U6000 (N_6000,N_5425,N_5551);
xnor U6001 (N_6001,N_5833,N_5951);
xnor U6002 (N_6002,N_5504,N_5430);
and U6003 (N_6003,N_5666,N_5723);
nand U6004 (N_6004,N_5634,N_5885);
and U6005 (N_6005,N_5645,N_5429);
xnor U6006 (N_6006,N_5703,N_5438);
or U6007 (N_6007,N_5537,N_5939);
or U6008 (N_6008,N_5948,N_5995);
xor U6009 (N_6009,N_5536,N_5938);
nor U6010 (N_6010,N_5636,N_5888);
and U6011 (N_6011,N_5497,N_5968);
or U6012 (N_6012,N_5731,N_5820);
and U6013 (N_6013,N_5729,N_5979);
nor U6014 (N_6014,N_5475,N_5664);
xor U6015 (N_6015,N_5500,N_5622);
nand U6016 (N_6016,N_5456,N_5806);
nor U6017 (N_6017,N_5836,N_5866);
nor U6018 (N_6018,N_5424,N_5800);
xnor U6019 (N_6019,N_5419,N_5615);
nand U6020 (N_6020,N_5743,N_5693);
nand U6021 (N_6021,N_5522,N_5597);
nand U6022 (N_6022,N_5762,N_5576);
and U6023 (N_6023,N_5665,N_5802);
and U6024 (N_6024,N_5959,N_5520);
xor U6025 (N_6025,N_5416,N_5683);
xor U6026 (N_6026,N_5514,N_5450);
or U6027 (N_6027,N_5752,N_5541);
nor U6028 (N_6028,N_5728,N_5978);
xnor U6029 (N_6029,N_5909,N_5851);
or U6030 (N_6030,N_5489,N_5878);
and U6031 (N_6031,N_5630,N_5805);
and U6032 (N_6032,N_5473,N_5761);
nor U6033 (N_6033,N_5692,N_5527);
and U6034 (N_6034,N_5760,N_5765);
xnor U6035 (N_6035,N_5563,N_5400);
nor U6036 (N_6036,N_5508,N_5492);
and U6037 (N_6037,N_5737,N_5980);
nor U6038 (N_6038,N_5436,N_5816);
and U6039 (N_6039,N_5782,N_5523);
and U6040 (N_6040,N_5710,N_5553);
nor U6041 (N_6041,N_5480,N_5907);
xnor U6042 (N_6042,N_5697,N_5864);
xnor U6043 (N_6043,N_5644,N_5470);
or U6044 (N_6044,N_5577,N_5656);
and U6045 (N_6045,N_5617,N_5845);
and U6046 (N_6046,N_5621,N_5844);
nor U6047 (N_6047,N_5659,N_5635);
nor U6048 (N_6048,N_5969,N_5768);
and U6049 (N_6049,N_5991,N_5705);
nand U6050 (N_6050,N_5602,N_5785);
and U6051 (N_6051,N_5799,N_5435);
nor U6052 (N_6052,N_5838,N_5603);
or U6053 (N_6053,N_5414,N_5794);
xnor U6054 (N_6054,N_5755,N_5401);
nand U6055 (N_6055,N_5774,N_5673);
nor U6056 (N_6056,N_5789,N_5787);
xor U6057 (N_6057,N_5931,N_5559);
nand U6058 (N_6058,N_5839,N_5449);
xor U6059 (N_6059,N_5646,N_5674);
xor U6060 (N_6060,N_5834,N_5680);
nand U6061 (N_6061,N_5894,N_5406);
xnor U6062 (N_6062,N_5596,N_5957);
nand U6063 (N_6063,N_5733,N_5854);
xor U6064 (N_6064,N_5681,N_5601);
nor U6065 (N_6065,N_5605,N_5546);
nor U6066 (N_6066,N_5405,N_5444);
xnor U6067 (N_6067,N_5792,N_5496);
nand U6068 (N_6068,N_5403,N_5465);
or U6069 (N_6069,N_5462,N_5619);
or U6070 (N_6070,N_5547,N_5498);
or U6071 (N_6071,N_5455,N_5640);
nand U6072 (N_6072,N_5418,N_5686);
nand U6073 (N_6073,N_5947,N_5638);
and U6074 (N_6074,N_5706,N_5722);
and U6075 (N_6075,N_5687,N_5675);
or U6076 (N_6076,N_5540,N_5671);
and U6077 (N_6077,N_5562,N_5891);
nor U6078 (N_6078,N_5786,N_5572);
or U6079 (N_6079,N_5519,N_5698);
and U6080 (N_6080,N_5433,N_5753);
and U6081 (N_6081,N_5738,N_5837);
nand U6082 (N_6082,N_5846,N_5431);
and U6083 (N_6083,N_5502,N_5653);
nand U6084 (N_6084,N_5442,N_5767);
and U6085 (N_6085,N_5936,N_5955);
xor U6086 (N_6086,N_5925,N_5823);
nand U6087 (N_6087,N_5975,N_5428);
or U6088 (N_6088,N_5921,N_5443);
and U6089 (N_6089,N_5727,N_5411);
nor U6090 (N_6090,N_5953,N_5808);
and U6091 (N_6091,N_5495,N_5629);
and U6092 (N_6092,N_5460,N_5631);
nor U6093 (N_6093,N_5626,N_5696);
nor U6094 (N_6094,N_5604,N_5790);
nor U6095 (N_6095,N_5591,N_5668);
and U6096 (N_6096,N_5814,N_5889);
nand U6097 (N_6097,N_5771,N_5825);
nor U6098 (N_6098,N_5924,N_5875);
and U6099 (N_6099,N_5459,N_5482);
nand U6100 (N_6100,N_5734,N_5478);
nor U6101 (N_6101,N_5472,N_5565);
nor U6102 (N_6102,N_5560,N_5558);
nand U6103 (N_6103,N_5486,N_5454);
or U6104 (N_6104,N_5960,N_5943);
or U6105 (N_6105,N_5999,N_5840);
and U6106 (N_6106,N_5775,N_5507);
or U6107 (N_6107,N_5667,N_5881);
nor U6108 (N_6108,N_5702,N_5783);
and U6109 (N_6109,N_5655,N_5561);
nand U6110 (N_6110,N_5898,N_5842);
xnor U6111 (N_6111,N_5873,N_5926);
and U6112 (N_6112,N_5677,N_5518);
or U6113 (N_6113,N_5609,N_5652);
or U6114 (N_6114,N_5554,N_5803);
or U6115 (N_6115,N_5874,N_5528);
and U6116 (N_6116,N_5896,N_5773);
and U6117 (N_6117,N_5918,N_5440);
nand U6118 (N_6118,N_5707,N_5699);
nand U6119 (N_6119,N_5920,N_5872);
and U6120 (N_6120,N_5643,N_5749);
nand U6121 (N_6121,N_5479,N_5410);
nor U6122 (N_6122,N_5451,N_5915);
nand U6123 (N_6123,N_5510,N_5982);
xnor U6124 (N_6124,N_5530,N_5592);
and U6125 (N_6125,N_5932,N_5748);
or U6126 (N_6126,N_5902,N_5973);
or U6127 (N_6127,N_5946,N_5858);
nor U6128 (N_6128,N_5746,N_5556);
nor U6129 (N_6129,N_5817,N_5917);
or U6130 (N_6130,N_5550,N_5952);
nor U6131 (N_6131,N_5735,N_5777);
nor U6132 (N_6132,N_5684,N_5564);
or U6133 (N_6133,N_5649,N_5719);
nor U6134 (N_6134,N_5614,N_5750);
or U6135 (N_6135,N_5937,N_5966);
and U6136 (N_6136,N_5543,N_5670);
xnor U6137 (N_6137,N_5608,N_5648);
nand U6138 (N_6138,N_5704,N_5852);
xor U6139 (N_6139,N_5720,N_5815);
and U6140 (N_6140,N_5654,N_5911);
nand U6141 (N_6141,N_5914,N_5869);
xnor U6142 (N_6142,N_5461,N_5521);
nor U6143 (N_6143,N_5439,N_5579);
or U6144 (N_6144,N_5819,N_5574);
nand U6145 (N_6145,N_5716,N_5611);
and U6146 (N_6146,N_5493,N_5474);
nor U6147 (N_6147,N_5594,N_5853);
and U6148 (N_6148,N_5784,N_5632);
or U6149 (N_6149,N_5669,N_5534);
xnor U6150 (N_6150,N_5580,N_5679);
or U6151 (N_6151,N_5744,N_5883);
or U6152 (N_6152,N_5730,N_5930);
nand U6153 (N_6153,N_5432,N_5905);
xnor U6154 (N_6154,N_5445,N_5971);
nor U6155 (N_6155,N_5595,N_5721);
or U6156 (N_6156,N_5695,N_5962);
nor U6157 (N_6157,N_5447,N_5647);
xnor U6158 (N_6158,N_5402,N_5548);
nand U6159 (N_6159,N_5877,N_5818);
xor U6160 (N_6160,N_5779,N_5426);
or U6161 (N_6161,N_5657,N_5996);
nand U6162 (N_6162,N_5587,N_5468);
xor U6163 (N_6163,N_5711,N_5639);
and U6164 (N_6164,N_5778,N_5860);
nand U6165 (N_6165,N_5830,N_5857);
nor U6166 (N_6166,N_5490,N_5529);
or U6167 (N_6167,N_5987,N_5689);
xor U6168 (N_6168,N_5812,N_5484);
and U6169 (N_6169,N_5855,N_5974);
and U6170 (N_6170,N_5847,N_5581);
or U6171 (N_6171,N_5567,N_5584);
and U6172 (N_6172,N_5678,N_5694);
nand U6173 (N_6173,N_5663,N_5828);
and U6174 (N_6174,N_5944,N_5506);
nand U6175 (N_6175,N_5709,N_5856);
nand U6176 (N_6176,N_5566,N_5739);
or U6177 (N_6177,N_5763,N_5415);
nand U6178 (N_6178,N_5813,N_5998);
nor U6179 (N_6179,N_5713,N_5977);
nand U6180 (N_6180,N_5916,N_5637);
nand U6181 (N_6181,N_5868,N_5607);
xor U6182 (N_6182,N_5967,N_5427);
nor U6183 (N_6183,N_5688,N_5796);
xor U6184 (N_6184,N_5661,N_5824);
nor U6185 (N_6185,N_5535,N_5981);
xnor U6186 (N_6186,N_5690,N_5954);
nand U6187 (N_6187,N_5811,N_5420);
nor U6188 (N_6188,N_5897,N_5821);
nor U6189 (N_6189,N_5516,N_5745);
and U6190 (N_6190,N_5985,N_5476);
or U6191 (N_6191,N_5423,N_5965);
and U6192 (N_6192,N_5448,N_5512);
or U6193 (N_6193,N_5776,N_5807);
and U6194 (N_6194,N_5539,N_5606);
xor U6195 (N_6195,N_5732,N_5826);
xor U6196 (N_6196,N_5549,N_5757);
or U6197 (N_6197,N_5984,N_5452);
nand U6198 (N_6198,N_5513,N_5804);
or U6199 (N_6199,N_5437,N_5725);
xnor U6200 (N_6200,N_5742,N_5988);
xor U6201 (N_6201,N_5741,N_5612);
xnor U6202 (N_6202,N_5588,N_5571);
or U6203 (N_6203,N_5515,N_5867);
nand U6204 (N_6204,N_5458,N_5582);
or U6205 (N_6205,N_5660,N_5600);
and U6206 (N_6206,N_5469,N_5624);
or U6207 (N_6207,N_5511,N_5958);
xor U6208 (N_6208,N_5487,N_5485);
nand U6209 (N_6209,N_5747,N_5471);
and U6210 (N_6210,N_5569,N_5770);
and U6211 (N_6211,N_5503,N_5434);
or U6212 (N_6212,N_5633,N_5895);
or U6213 (N_6213,N_5583,N_5578);
nand U6214 (N_6214,N_5526,N_5740);
or U6215 (N_6215,N_5751,N_5797);
and U6216 (N_6216,N_5850,N_5422);
xnor U6217 (N_6217,N_5708,N_5533);
nor U6218 (N_6218,N_5993,N_5417);
xor U6219 (N_6219,N_5772,N_5464);
and U6220 (N_6220,N_5650,N_5809);
xor U6221 (N_6221,N_5788,N_5963);
or U6222 (N_6222,N_5682,N_5618);
nand U6223 (N_6223,N_5552,N_5901);
nor U6224 (N_6224,N_5651,N_5590);
nor U6225 (N_6225,N_5736,N_5863);
and U6226 (N_6226,N_5766,N_5832);
or U6227 (N_6227,N_5893,N_5919);
or U6228 (N_6228,N_5467,N_5940);
nor U6229 (N_6229,N_5672,N_5892);
nand U6230 (N_6230,N_5827,N_5463);
nand U6231 (N_6231,N_5625,N_5499);
xnor U6232 (N_6232,N_5585,N_5570);
and U6233 (N_6233,N_5421,N_5509);
nor U6234 (N_6234,N_5876,N_5532);
nor U6235 (N_6235,N_5859,N_5829);
or U6236 (N_6236,N_5997,N_5404);
nor U6237 (N_6237,N_5861,N_5906);
or U6238 (N_6238,N_5505,N_5976);
and U6239 (N_6239,N_5593,N_5620);
and U6240 (N_6240,N_5642,N_5409);
and U6241 (N_6241,N_5555,N_5890);
xor U6242 (N_6242,N_5950,N_5457);
and U6243 (N_6243,N_5589,N_5483);
and U6244 (N_6244,N_5949,N_5575);
nor U6245 (N_6245,N_5942,N_5408);
nand U6246 (N_6246,N_5862,N_5481);
and U6247 (N_6247,N_5964,N_5913);
and U6248 (N_6248,N_5758,N_5544);
and U6249 (N_6249,N_5972,N_5904);
xnor U6250 (N_6250,N_5441,N_5627);
nor U6251 (N_6251,N_5880,N_5494);
nand U6252 (N_6252,N_5488,N_5798);
and U6253 (N_6253,N_5517,N_5992);
nor U6254 (N_6254,N_5871,N_5849);
xor U6255 (N_6255,N_5835,N_5886);
nand U6256 (N_6256,N_5412,N_5870);
xnor U6257 (N_6257,N_5879,N_5717);
or U6258 (N_6258,N_5754,N_5793);
nor U6259 (N_6259,N_5781,N_5928);
nand U6260 (N_6260,N_5910,N_5882);
nor U6261 (N_6261,N_5941,N_5961);
and U6262 (N_6262,N_5714,N_5922);
and U6263 (N_6263,N_5613,N_5477);
nor U6264 (N_6264,N_5945,N_5685);
nor U6265 (N_6265,N_5446,N_5676);
nand U6266 (N_6266,N_5769,N_5843);
or U6267 (N_6267,N_5887,N_5933);
nor U6268 (N_6268,N_5641,N_5822);
xor U6269 (N_6269,N_5935,N_5691);
or U6270 (N_6270,N_5568,N_5501);
or U6271 (N_6271,N_5923,N_5970);
or U6272 (N_6272,N_5801,N_5759);
nor U6273 (N_6273,N_5929,N_5542);
or U6274 (N_6274,N_5756,N_5701);
nor U6275 (N_6275,N_5616,N_5712);
or U6276 (N_6276,N_5662,N_5715);
nor U6277 (N_6277,N_5831,N_5524);
nor U6278 (N_6278,N_5903,N_5628);
or U6279 (N_6279,N_5453,N_5810);
and U6280 (N_6280,N_5956,N_5764);
nor U6281 (N_6281,N_5599,N_5586);
and U6282 (N_6282,N_5658,N_5538);
nand U6283 (N_6283,N_5718,N_5573);
or U6284 (N_6284,N_5990,N_5623);
nor U6285 (N_6285,N_5525,N_5989);
or U6286 (N_6286,N_5927,N_5610);
nand U6287 (N_6287,N_5884,N_5466);
nand U6288 (N_6288,N_5531,N_5491);
xnor U6289 (N_6289,N_5994,N_5900);
and U6290 (N_6290,N_5865,N_5724);
nor U6291 (N_6291,N_5986,N_5899);
or U6292 (N_6292,N_5908,N_5413);
nor U6293 (N_6293,N_5780,N_5545);
or U6294 (N_6294,N_5557,N_5841);
xor U6295 (N_6295,N_5791,N_5700);
nand U6296 (N_6296,N_5407,N_5848);
nand U6297 (N_6297,N_5912,N_5934);
xnor U6298 (N_6298,N_5726,N_5598);
nand U6299 (N_6299,N_5795,N_5983);
xor U6300 (N_6300,N_5859,N_5675);
xor U6301 (N_6301,N_5739,N_5644);
or U6302 (N_6302,N_5545,N_5446);
nor U6303 (N_6303,N_5737,N_5667);
nand U6304 (N_6304,N_5765,N_5892);
xor U6305 (N_6305,N_5466,N_5888);
nand U6306 (N_6306,N_5407,N_5663);
nor U6307 (N_6307,N_5686,N_5874);
or U6308 (N_6308,N_5991,N_5673);
or U6309 (N_6309,N_5463,N_5560);
nor U6310 (N_6310,N_5722,N_5446);
nor U6311 (N_6311,N_5553,N_5525);
and U6312 (N_6312,N_5884,N_5885);
or U6313 (N_6313,N_5757,N_5985);
xnor U6314 (N_6314,N_5746,N_5653);
or U6315 (N_6315,N_5712,N_5476);
and U6316 (N_6316,N_5626,N_5723);
and U6317 (N_6317,N_5852,N_5967);
nor U6318 (N_6318,N_5672,N_5573);
and U6319 (N_6319,N_5714,N_5904);
xor U6320 (N_6320,N_5647,N_5646);
nand U6321 (N_6321,N_5749,N_5896);
or U6322 (N_6322,N_5660,N_5702);
and U6323 (N_6323,N_5765,N_5440);
xor U6324 (N_6324,N_5803,N_5912);
or U6325 (N_6325,N_5478,N_5675);
nor U6326 (N_6326,N_5464,N_5993);
nand U6327 (N_6327,N_5419,N_5989);
and U6328 (N_6328,N_5609,N_5700);
nor U6329 (N_6329,N_5954,N_5605);
nor U6330 (N_6330,N_5602,N_5452);
or U6331 (N_6331,N_5526,N_5601);
nor U6332 (N_6332,N_5489,N_5879);
xor U6333 (N_6333,N_5609,N_5552);
xor U6334 (N_6334,N_5993,N_5906);
xnor U6335 (N_6335,N_5712,N_5582);
and U6336 (N_6336,N_5415,N_5765);
nor U6337 (N_6337,N_5551,N_5642);
xor U6338 (N_6338,N_5597,N_5430);
or U6339 (N_6339,N_5769,N_5781);
or U6340 (N_6340,N_5541,N_5929);
xor U6341 (N_6341,N_5932,N_5910);
nand U6342 (N_6342,N_5730,N_5632);
and U6343 (N_6343,N_5493,N_5745);
xnor U6344 (N_6344,N_5501,N_5444);
nand U6345 (N_6345,N_5811,N_5867);
nor U6346 (N_6346,N_5591,N_5606);
nor U6347 (N_6347,N_5986,N_5794);
nand U6348 (N_6348,N_5890,N_5813);
nor U6349 (N_6349,N_5724,N_5552);
and U6350 (N_6350,N_5539,N_5607);
xor U6351 (N_6351,N_5985,N_5758);
xnor U6352 (N_6352,N_5694,N_5817);
and U6353 (N_6353,N_5793,N_5557);
or U6354 (N_6354,N_5960,N_5687);
nand U6355 (N_6355,N_5884,N_5986);
or U6356 (N_6356,N_5948,N_5778);
nand U6357 (N_6357,N_5576,N_5402);
nand U6358 (N_6358,N_5649,N_5562);
nor U6359 (N_6359,N_5623,N_5677);
or U6360 (N_6360,N_5994,N_5682);
and U6361 (N_6361,N_5928,N_5440);
xor U6362 (N_6362,N_5876,N_5874);
nand U6363 (N_6363,N_5782,N_5462);
and U6364 (N_6364,N_5693,N_5415);
xor U6365 (N_6365,N_5613,N_5948);
or U6366 (N_6366,N_5848,N_5717);
and U6367 (N_6367,N_5710,N_5451);
nand U6368 (N_6368,N_5806,N_5966);
or U6369 (N_6369,N_5823,N_5955);
nand U6370 (N_6370,N_5449,N_5662);
and U6371 (N_6371,N_5787,N_5841);
nor U6372 (N_6372,N_5439,N_5810);
nor U6373 (N_6373,N_5540,N_5537);
nand U6374 (N_6374,N_5992,N_5589);
and U6375 (N_6375,N_5657,N_5560);
xnor U6376 (N_6376,N_5991,N_5893);
nor U6377 (N_6377,N_5496,N_5552);
and U6378 (N_6378,N_5412,N_5687);
and U6379 (N_6379,N_5459,N_5752);
and U6380 (N_6380,N_5821,N_5900);
and U6381 (N_6381,N_5810,N_5538);
or U6382 (N_6382,N_5813,N_5489);
and U6383 (N_6383,N_5525,N_5988);
nor U6384 (N_6384,N_5788,N_5797);
and U6385 (N_6385,N_5490,N_5740);
or U6386 (N_6386,N_5949,N_5633);
and U6387 (N_6387,N_5936,N_5854);
xnor U6388 (N_6388,N_5903,N_5591);
or U6389 (N_6389,N_5447,N_5710);
or U6390 (N_6390,N_5800,N_5877);
or U6391 (N_6391,N_5501,N_5749);
and U6392 (N_6392,N_5864,N_5705);
nor U6393 (N_6393,N_5673,N_5401);
nor U6394 (N_6394,N_5997,N_5688);
nand U6395 (N_6395,N_5668,N_5452);
nand U6396 (N_6396,N_5436,N_5475);
or U6397 (N_6397,N_5997,N_5435);
nor U6398 (N_6398,N_5743,N_5760);
or U6399 (N_6399,N_5578,N_5635);
nor U6400 (N_6400,N_5999,N_5643);
and U6401 (N_6401,N_5427,N_5573);
and U6402 (N_6402,N_5603,N_5429);
nand U6403 (N_6403,N_5624,N_5656);
and U6404 (N_6404,N_5675,N_5481);
nor U6405 (N_6405,N_5570,N_5899);
and U6406 (N_6406,N_5411,N_5459);
nor U6407 (N_6407,N_5967,N_5556);
or U6408 (N_6408,N_5654,N_5533);
xor U6409 (N_6409,N_5698,N_5646);
or U6410 (N_6410,N_5940,N_5814);
xnor U6411 (N_6411,N_5428,N_5584);
or U6412 (N_6412,N_5588,N_5617);
nor U6413 (N_6413,N_5464,N_5793);
and U6414 (N_6414,N_5476,N_5428);
or U6415 (N_6415,N_5724,N_5912);
xnor U6416 (N_6416,N_5623,N_5885);
nand U6417 (N_6417,N_5698,N_5678);
nor U6418 (N_6418,N_5826,N_5658);
and U6419 (N_6419,N_5987,N_5630);
nor U6420 (N_6420,N_5464,N_5614);
or U6421 (N_6421,N_5758,N_5790);
or U6422 (N_6422,N_5401,N_5626);
nand U6423 (N_6423,N_5995,N_5965);
nor U6424 (N_6424,N_5951,N_5821);
nor U6425 (N_6425,N_5915,N_5415);
nand U6426 (N_6426,N_5807,N_5820);
nor U6427 (N_6427,N_5444,N_5660);
nand U6428 (N_6428,N_5906,N_5970);
nor U6429 (N_6429,N_5424,N_5616);
xor U6430 (N_6430,N_5894,N_5581);
and U6431 (N_6431,N_5539,N_5428);
xnor U6432 (N_6432,N_5509,N_5561);
nand U6433 (N_6433,N_5728,N_5740);
xnor U6434 (N_6434,N_5514,N_5410);
or U6435 (N_6435,N_5629,N_5848);
nor U6436 (N_6436,N_5814,N_5599);
and U6437 (N_6437,N_5723,N_5980);
or U6438 (N_6438,N_5753,N_5873);
xor U6439 (N_6439,N_5593,N_5653);
and U6440 (N_6440,N_5596,N_5793);
and U6441 (N_6441,N_5420,N_5497);
or U6442 (N_6442,N_5807,N_5404);
or U6443 (N_6443,N_5906,N_5524);
nand U6444 (N_6444,N_5691,N_5838);
xor U6445 (N_6445,N_5734,N_5899);
xnor U6446 (N_6446,N_5581,N_5418);
or U6447 (N_6447,N_5749,N_5797);
xnor U6448 (N_6448,N_5813,N_5567);
and U6449 (N_6449,N_5407,N_5519);
xor U6450 (N_6450,N_5929,N_5728);
and U6451 (N_6451,N_5620,N_5815);
and U6452 (N_6452,N_5407,N_5601);
nor U6453 (N_6453,N_5771,N_5618);
nand U6454 (N_6454,N_5695,N_5421);
and U6455 (N_6455,N_5802,N_5772);
nor U6456 (N_6456,N_5988,N_5699);
and U6457 (N_6457,N_5893,N_5627);
or U6458 (N_6458,N_5956,N_5930);
xnor U6459 (N_6459,N_5935,N_5416);
or U6460 (N_6460,N_5720,N_5761);
nand U6461 (N_6461,N_5909,N_5533);
nor U6462 (N_6462,N_5929,N_5455);
nand U6463 (N_6463,N_5816,N_5595);
nor U6464 (N_6464,N_5435,N_5753);
nand U6465 (N_6465,N_5801,N_5502);
or U6466 (N_6466,N_5945,N_5452);
and U6467 (N_6467,N_5537,N_5476);
or U6468 (N_6468,N_5997,N_5750);
and U6469 (N_6469,N_5474,N_5480);
nor U6470 (N_6470,N_5912,N_5676);
nand U6471 (N_6471,N_5888,N_5508);
and U6472 (N_6472,N_5954,N_5784);
nor U6473 (N_6473,N_5915,N_5400);
and U6474 (N_6474,N_5522,N_5420);
or U6475 (N_6475,N_5829,N_5574);
xor U6476 (N_6476,N_5630,N_5875);
xor U6477 (N_6477,N_5480,N_5559);
xor U6478 (N_6478,N_5627,N_5870);
and U6479 (N_6479,N_5413,N_5741);
nor U6480 (N_6480,N_5646,N_5904);
and U6481 (N_6481,N_5514,N_5714);
xor U6482 (N_6482,N_5711,N_5977);
nor U6483 (N_6483,N_5708,N_5438);
or U6484 (N_6484,N_5462,N_5888);
nor U6485 (N_6485,N_5724,N_5992);
nand U6486 (N_6486,N_5719,N_5937);
and U6487 (N_6487,N_5667,N_5796);
xor U6488 (N_6488,N_5600,N_5412);
nor U6489 (N_6489,N_5923,N_5963);
and U6490 (N_6490,N_5487,N_5515);
xnor U6491 (N_6491,N_5499,N_5426);
nor U6492 (N_6492,N_5946,N_5859);
and U6493 (N_6493,N_5770,N_5652);
and U6494 (N_6494,N_5656,N_5798);
nand U6495 (N_6495,N_5407,N_5936);
nand U6496 (N_6496,N_5493,N_5717);
nor U6497 (N_6497,N_5495,N_5509);
nor U6498 (N_6498,N_5918,N_5454);
or U6499 (N_6499,N_5491,N_5850);
or U6500 (N_6500,N_5401,N_5470);
xnor U6501 (N_6501,N_5824,N_5648);
and U6502 (N_6502,N_5971,N_5821);
and U6503 (N_6503,N_5458,N_5566);
or U6504 (N_6504,N_5654,N_5989);
and U6505 (N_6505,N_5878,N_5873);
nor U6506 (N_6506,N_5649,N_5591);
nor U6507 (N_6507,N_5683,N_5877);
nand U6508 (N_6508,N_5785,N_5839);
xnor U6509 (N_6509,N_5426,N_5643);
nor U6510 (N_6510,N_5438,N_5613);
and U6511 (N_6511,N_5756,N_5487);
nor U6512 (N_6512,N_5546,N_5986);
nor U6513 (N_6513,N_5587,N_5950);
nor U6514 (N_6514,N_5637,N_5608);
nor U6515 (N_6515,N_5488,N_5653);
xor U6516 (N_6516,N_5882,N_5477);
xnor U6517 (N_6517,N_5636,N_5631);
or U6518 (N_6518,N_5643,N_5452);
or U6519 (N_6519,N_5949,N_5803);
or U6520 (N_6520,N_5817,N_5801);
nor U6521 (N_6521,N_5809,N_5942);
and U6522 (N_6522,N_5768,N_5939);
nand U6523 (N_6523,N_5544,N_5677);
xor U6524 (N_6524,N_5834,N_5996);
and U6525 (N_6525,N_5812,N_5646);
xnor U6526 (N_6526,N_5956,N_5576);
nand U6527 (N_6527,N_5526,N_5481);
and U6528 (N_6528,N_5561,N_5931);
or U6529 (N_6529,N_5581,N_5804);
nand U6530 (N_6530,N_5432,N_5419);
or U6531 (N_6531,N_5777,N_5637);
xor U6532 (N_6532,N_5857,N_5686);
nor U6533 (N_6533,N_5650,N_5618);
nand U6534 (N_6534,N_5458,N_5522);
nand U6535 (N_6535,N_5465,N_5738);
nor U6536 (N_6536,N_5585,N_5979);
and U6537 (N_6537,N_5912,N_5837);
or U6538 (N_6538,N_5944,N_5659);
or U6539 (N_6539,N_5503,N_5766);
nor U6540 (N_6540,N_5782,N_5596);
nor U6541 (N_6541,N_5943,N_5656);
nand U6542 (N_6542,N_5967,N_5746);
or U6543 (N_6543,N_5411,N_5430);
or U6544 (N_6544,N_5712,N_5966);
or U6545 (N_6545,N_5573,N_5945);
xor U6546 (N_6546,N_5719,N_5409);
nor U6547 (N_6547,N_5654,N_5487);
xnor U6548 (N_6548,N_5496,N_5426);
or U6549 (N_6549,N_5763,N_5880);
xor U6550 (N_6550,N_5637,N_5954);
or U6551 (N_6551,N_5605,N_5517);
and U6552 (N_6552,N_5500,N_5437);
nand U6553 (N_6553,N_5692,N_5686);
and U6554 (N_6554,N_5939,N_5633);
xnor U6555 (N_6555,N_5554,N_5740);
nor U6556 (N_6556,N_5834,N_5403);
nor U6557 (N_6557,N_5741,N_5742);
and U6558 (N_6558,N_5708,N_5981);
or U6559 (N_6559,N_5604,N_5427);
or U6560 (N_6560,N_5973,N_5429);
and U6561 (N_6561,N_5833,N_5994);
and U6562 (N_6562,N_5662,N_5736);
nand U6563 (N_6563,N_5710,N_5681);
nor U6564 (N_6564,N_5508,N_5820);
or U6565 (N_6565,N_5873,N_5590);
or U6566 (N_6566,N_5890,N_5962);
xor U6567 (N_6567,N_5603,N_5749);
and U6568 (N_6568,N_5875,N_5794);
or U6569 (N_6569,N_5962,N_5582);
xor U6570 (N_6570,N_5643,N_5404);
nand U6571 (N_6571,N_5965,N_5533);
nor U6572 (N_6572,N_5862,N_5509);
nand U6573 (N_6573,N_5757,N_5638);
nor U6574 (N_6574,N_5811,N_5682);
or U6575 (N_6575,N_5711,N_5998);
nand U6576 (N_6576,N_5502,N_5602);
or U6577 (N_6577,N_5561,N_5927);
nand U6578 (N_6578,N_5596,N_5632);
and U6579 (N_6579,N_5761,N_5834);
nand U6580 (N_6580,N_5650,N_5775);
nor U6581 (N_6581,N_5803,N_5500);
and U6582 (N_6582,N_5779,N_5998);
or U6583 (N_6583,N_5840,N_5912);
nand U6584 (N_6584,N_5670,N_5974);
or U6585 (N_6585,N_5531,N_5974);
and U6586 (N_6586,N_5947,N_5400);
or U6587 (N_6587,N_5782,N_5962);
xnor U6588 (N_6588,N_5694,N_5436);
or U6589 (N_6589,N_5803,N_5625);
nor U6590 (N_6590,N_5462,N_5802);
xnor U6591 (N_6591,N_5807,N_5969);
or U6592 (N_6592,N_5959,N_5745);
or U6593 (N_6593,N_5853,N_5989);
xor U6594 (N_6594,N_5418,N_5950);
nor U6595 (N_6595,N_5401,N_5865);
nand U6596 (N_6596,N_5735,N_5504);
or U6597 (N_6597,N_5525,N_5435);
nand U6598 (N_6598,N_5666,N_5928);
or U6599 (N_6599,N_5455,N_5578);
and U6600 (N_6600,N_6372,N_6255);
or U6601 (N_6601,N_6067,N_6021);
nand U6602 (N_6602,N_6541,N_6418);
nor U6603 (N_6603,N_6078,N_6026);
nor U6604 (N_6604,N_6037,N_6044);
xnor U6605 (N_6605,N_6579,N_6390);
nand U6606 (N_6606,N_6226,N_6259);
nor U6607 (N_6607,N_6353,N_6109);
nor U6608 (N_6608,N_6128,N_6229);
or U6609 (N_6609,N_6370,N_6360);
nand U6610 (N_6610,N_6264,N_6542);
nor U6611 (N_6611,N_6003,N_6237);
nand U6612 (N_6612,N_6130,N_6586);
nor U6613 (N_6613,N_6272,N_6295);
nor U6614 (N_6614,N_6136,N_6431);
or U6615 (N_6615,N_6450,N_6197);
and U6616 (N_6616,N_6001,N_6269);
and U6617 (N_6617,N_6350,N_6207);
xor U6618 (N_6618,N_6564,N_6482);
or U6619 (N_6619,N_6270,N_6010);
nor U6620 (N_6620,N_6235,N_6315);
and U6621 (N_6621,N_6420,N_6498);
nand U6622 (N_6622,N_6361,N_6287);
nor U6623 (N_6623,N_6545,N_6250);
xnor U6624 (N_6624,N_6494,N_6112);
nand U6625 (N_6625,N_6313,N_6457);
nand U6626 (N_6626,N_6331,N_6203);
and U6627 (N_6627,N_6210,N_6345);
nand U6628 (N_6628,N_6260,N_6336);
nor U6629 (N_6629,N_6154,N_6521);
nand U6630 (N_6630,N_6267,N_6576);
and U6631 (N_6631,N_6583,N_6507);
xor U6632 (N_6632,N_6181,N_6569);
xnor U6633 (N_6633,N_6174,N_6536);
xnor U6634 (N_6634,N_6043,N_6311);
nand U6635 (N_6635,N_6359,N_6594);
nand U6636 (N_6636,N_6164,N_6399);
nand U6637 (N_6637,N_6469,N_6434);
xnor U6638 (N_6638,N_6428,N_6484);
and U6639 (N_6639,N_6571,N_6157);
xor U6640 (N_6640,N_6135,N_6076);
nand U6641 (N_6641,N_6139,N_6306);
or U6642 (N_6642,N_6387,N_6349);
or U6643 (N_6643,N_6371,N_6286);
nor U6644 (N_6644,N_6265,N_6432);
nand U6645 (N_6645,N_6563,N_6517);
xor U6646 (N_6646,N_6351,N_6334);
nor U6647 (N_6647,N_6053,N_6453);
xor U6648 (N_6648,N_6276,N_6329);
or U6649 (N_6649,N_6111,N_6554);
nand U6650 (N_6650,N_6014,N_6256);
or U6651 (N_6651,N_6445,N_6557);
nor U6652 (N_6652,N_6142,N_6346);
or U6653 (N_6653,N_6598,N_6296);
and U6654 (N_6654,N_6467,N_6121);
nand U6655 (N_6655,N_6558,N_6385);
and U6656 (N_6656,N_6447,N_6289);
nor U6657 (N_6657,N_6592,N_6438);
or U6658 (N_6658,N_6580,N_6298);
and U6659 (N_6659,N_6200,N_6188);
and U6660 (N_6660,N_6034,N_6326);
or U6661 (N_6661,N_6282,N_6032);
nor U6662 (N_6662,N_6096,N_6468);
or U6663 (N_6663,N_6082,N_6147);
or U6664 (N_6664,N_6068,N_6332);
or U6665 (N_6665,N_6597,N_6069);
or U6666 (N_6666,N_6514,N_6429);
or U6667 (N_6667,N_6187,N_6570);
xnor U6668 (N_6668,N_6045,N_6040);
and U6669 (N_6669,N_6333,N_6340);
and U6670 (N_6670,N_6347,N_6481);
nand U6671 (N_6671,N_6411,N_6539);
or U6672 (N_6672,N_6522,N_6222);
nor U6673 (N_6673,N_6488,N_6195);
xor U6674 (N_6674,N_6101,N_6051);
or U6675 (N_6675,N_6392,N_6129);
nand U6676 (N_6676,N_6253,N_6492);
nor U6677 (N_6677,N_6449,N_6378);
or U6678 (N_6678,N_6283,N_6320);
nand U6679 (N_6679,N_6537,N_6466);
or U6680 (N_6680,N_6066,N_6202);
nand U6681 (N_6681,N_6508,N_6419);
xor U6682 (N_6682,N_6025,N_6527);
xnor U6683 (N_6683,N_6506,N_6070);
nand U6684 (N_6684,N_6451,N_6532);
or U6685 (N_6685,N_6132,N_6007);
nand U6686 (N_6686,N_6413,N_6116);
xnor U6687 (N_6687,N_6303,N_6131);
and U6688 (N_6688,N_6491,N_6213);
xor U6689 (N_6689,N_6100,N_6504);
xor U6690 (N_6690,N_6525,N_6127);
nor U6691 (N_6691,N_6156,N_6047);
nand U6692 (N_6692,N_6145,N_6487);
nand U6693 (N_6693,N_6178,N_6416);
nand U6694 (N_6694,N_6430,N_6016);
nand U6695 (N_6695,N_6182,N_6180);
xor U6696 (N_6696,N_6550,N_6089);
nor U6697 (N_6697,N_6081,N_6031);
nor U6698 (N_6698,N_6389,N_6301);
nand U6699 (N_6699,N_6042,N_6379);
nor U6700 (N_6700,N_6117,N_6470);
nor U6701 (N_6701,N_6199,N_6437);
and U6702 (N_6702,N_6423,N_6348);
and U6703 (N_6703,N_6510,N_6330);
xor U6704 (N_6704,N_6176,N_6046);
xnor U6705 (N_6705,N_6052,N_6146);
or U6706 (N_6706,N_6473,N_6593);
xnor U6707 (N_6707,N_6056,N_6412);
nor U6708 (N_6708,N_6551,N_6155);
xor U6709 (N_6709,N_6489,N_6408);
nor U6710 (N_6710,N_6054,N_6012);
nand U6711 (N_6711,N_6024,N_6472);
xor U6712 (N_6712,N_6533,N_6123);
or U6713 (N_6713,N_6198,N_6574);
nand U6714 (N_6714,N_6582,N_6020);
xnor U6715 (N_6715,N_6038,N_6595);
or U6716 (N_6716,N_6041,N_6236);
or U6717 (N_6717,N_6452,N_6059);
or U6718 (N_6718,N_6573,N_6144);
and U6719 (N_6719,N_6183,N_6138);
or U6720 (N_6720,N_6072,N_6165);
and U6721 (N_6721,N_6538,N_6327);
nor U6722 (N_6722,N_6141,N_6261);
or U6723 (N_6723,N_6175,N_6065);
or U6724 (N_6724,N_6302,N_6454);
nand U6725 (N_6725,N_6036,N_6160);
nor U6726 (N_6726,N_6446,N_6271);
or U6727 (N_6727,N_6425,N_6441);
or U6728 (N_6728,N_6247,N_6075);
and U6729 (N_6729,N_6562,N_6559);
and U6730 (N_6730,N_6575,N_6108);
nand U6731 (N_6731,N_6529,N_6325);
and U6732 (N_6732,N_6279,N_6581);
nand U6733 (N_6733,N_6495,N_6169);
nor U6734 (N_6734,N_6113,N_6401);
nor U6735 (N_6735,N_6208,N_6342);
or U6736 (N_6736,N_6212,N_6262);
or U6737 (N_6737,N_6364,N_6376);
nand U6738 (N_6738,N_6022,N_6166);
nor U6739 (N_6739,N_6167,N_6304);
and U6740 (N_6740,N_6149,N_6480);
xnor U6741 (N_6741,N_6162,N_6086);
or U6742 (N_6742,N_6458,N_6377);
nor U6743 (N_6743,N_6115,N_6502);
nor U6744 (N_6744,N_6388,N_6292);
and U6745 (N_6745,N_6414,N_6344);
or U6746 (N_6746,N_6382,N_6561);
and U6747 (N_6747,N_6114,N_6019);
xnor U6748 (N_6748,N_6515,N_6191);
and U6749 (N_6749,N_6552,N_6319);
or U6750 (N_6750,N_6201,N_6050);
xnor U6751 (N_6751,N_6493,N_6299);
nand U6752 (N_6752,N_6588,N_6355);
nor U6753 (N_6753,N_6280,N_6524);
xnor U6754 (N_6754,N_6476,N_6104);
or U6755 (N_6755,N_6530,N_6206);
or U6756 (N_6756,N_6546,N_6341);
and U6757 (N_6757,N_6005,N_6009);
nand U6758 (N_6758,N_6184,N_6268);
and U6759 (N_6759,N_6540,N_6547);
nand U6760 (N_6760,N_6107,N_6097);
xnor U6761 (N_6761,N_6211,N_6214);
and U6762 (N_6762,N_6231,N_6073);
or U6763 (N_6763,N_6193,N_6153);
nor U6764 (N_6764,N_6479,N_6396);
or U6765 (N_6765,N_6244,N_6589);
nand U6766 (N_6766,N_6219,N_6252);
or U6767 (N_6767,N_6105,N_6460);
and U6768 (N_6768,N_6405,N_6368);
nor U6769 (N_6769,N_6426,N_6061);
nor U6770 (N_6770,N_6230,N_6170);
and U6771 (N_6771,N_6316,N_6238);
and U6772 (N_6772,N_6465,N_6087);
or U6773 (N_6773,N_6375,N_6587);
and U6774 (N_6774,N_6281,N_6088);
nand U6775 (N_6775,N_6173,N_6543);
xnor U6776 (N_6776,N_6463,N_6343);
or U6777 (N_6777,N_6209,N_6158);
nor U6778 (N_6778,N_6442,N_6098);
and U6779 (N_6779,N_6596,N_6185);
nor U6780 (N_6780,N_6404,N_6433);
or U6781 (N_6781,N_6400,N_6365);
or U6782 (N_6782,N_6094,N_6080);
nor U6783 (N_6783,N_6216,N_6106);
xor U6784 (N_6784,N_6233,N_6528);
and U6785 (N_6785,N_6444,N_6566);
nor U6786 (N_6786,N_6555,N_6074);
and U6787 (N_6787,N_6018,N_6324);
and U6788 (N_6788,N_6239,N_6513);
and U6789 (N_6789,N_6168,N_6039);
nand U6790 (N_6790,N_6058,N_6410);
nand U6791 (N_6791,N_6358,N_6556);
nand U6792 (N_6792,N_6464,N_6189);
xnor U6793 (N_6793,N_6085,N_6186);
xnor U6794 (N_6794,N_6049,N_6227);
and U6795 (N_6795,N_6028,N_6534);
nand U6796 (N_6796,N_6338,N_6439);
nand U6797 (N_6797,N_6224,N_6249);
nor U6798 (N_6798,N_6383,N_6461);
xor U6799 (N_6799,N_6159,N_6505);
nor U6800 (N_6800,N_6143,N_6099);
nand U6801 (N_6801,N_6373,N_6415);
nor U6802 (N_6802,N_6218,N_6055);
and U6803 (N_6803,N_6228,N_6307);
nand U6804 (N_6804,N_6485,N_6578);
and U6805 (N_6805,N_6321,N_6590);
nand U6806 (N_6806,N_6374,N_6119);
xnor U6807 (N_6807,N_6223,N_6459);
or U6808 (N_6808,N_6384,N_6516);
xor U6809 (N_6809,N_6477,N_6294);
and U6810 (N_6810,N_6490,N_6064);
or U6811 (N_6811,N_6124,N_6462);
nand U6812 (N_6812,N_6352,N_6150);
xnor U6813 (N_6813,N_6328,N_6291);
nand U6814 (N_6814,N_6284,N_6548);
nand U6815 (N_6815,N_6406,N_6394);
and U6816 (N_6816,N_6565,N_6512);
xnor U6817 (N_6817,N_6486,N_6234);
xnor U6818 (N_6818,N_6205,N_6062);
or U6819 (N_6819,N_6093,N_6277);
nor U6820 (N_6820,N_6323,N_6478);
nor U6821 (N_6821,N_6572,N_6436);
nand U6822 (N_6822,N_6134,N_6083);
xor U6823 (N_6823,N_6310,N_6553);
nand U6824 (N_6824,N_6273,N_6474);
or U6825 (N_6825,N_6091,N_6000);
xnor U6826 (N_6826,N_6519,N_6397);
nor U6827 (N_6827,N_6435,N_6584);
or U6828 (N_6828,N_6403,N_6544);
and U6829 (N_6829,N_6006,N_6503);
xnor U6830 (N_6830,N_6071,N_6190);
and U6831 (N_6831,N_6560,N_6278);
nor U6832 (N_6832,N_6497,N_6290);
nand U6833 (N_6833,N_6318,N_6140);
and U6834 (N_6834,N_6363,N_6386);
xor U6835 (N_6835,N_6013,N_6285);
or U6836 (N_6836,N_6163,N_6221);
nor U6837 (N_6837,N_6004,N_6518);
or U6838 (N_6838,N_6297,N_6422);
or U6839 (N_6839,N_6526,N_6398);
xor U6840 (N_6840,N_6317,N_6417);
xnor U6841 (N_6841,N_6152,N_6500);
and U6842 (N_6842,N_6029,N_6585);
nor U6843 (N_6843,N_6090,N_6103);
or U6844 (N_6844,N_6015,N_6079);
nand U6845 (N_6845,N_6232,N_6240);
nand U6846 (N_6846,N_6033,N_6151);
nor U6847 (N_6847,N_6300,N_6366);
nor U6848 (N_6848,N_6274,N_6393);
nand U6849 (N_6849,N_6030,N_6194);
nand U6850 (N_6850,N_6266,N_6568);
nand U6851 (N_6851,N_6275,N_6309);
or U6852 (N_6852,N_6204,N_6288);
and U6853 (N_6853,N_6196,N_6443);
or U6854 (N_6854,N_6248,N_6337);
nor U6855 (N_6855,N_6395,N_6263);
nor U6856 (N_6856,N_6567,N_6241);
nand U6857 (N_6857,N_6314,N_6023);
or U6858 (N_6858,N_6357,N_6060);
nor U6859 (N_6859,N_6137,N_6354);
and U6860 (N_6860,N_6120,N_6535);
and U6861 (N_6861,N_6424,N_6448);
and U6862 (N_6862,N_6483,N_6225);
nor U6863 (N_6863,N_6475,N_6501);
xor U6864 (N_6864,N_6254,N_6499);
nor U6865 (N_6865,N_6092,N_6496);
or U6866 (N_6866,N_6381,N_6391);
nand U6867 (N_6867,N_6027,N_6148);
xor U6868 (N_6868,N_6246,N_6293);
or U6869 (N_6869,N_6102,N_6171);
xor U6870 (N_6870,N_6011,N_6511);
or U6871 (N_6871,N_6220,N_6577);
xnor U6872 (N_6872,N_6356,N_6427);
or U6873 (N_6873,N_6217,N_6380);
nor U6874 (N_6874,N_6367,N_6531);
nor U6875 (N_6875,N_6455,N_6599);
xor U6876 (N_6876,N_6245,N_6339);
nand U6877 (N_6877,N_6549,N_6509);
xor U6878 (N_6878,N_6161,N_6118);
xor U6879 (N_6879,N_6095,N_6057);
nor U6880 (N_6880,N_6308,N_6456);
nand U6881 (N_6881,N_6305,N_6242);
and U6882 (N_6882,N_6407,N_6257);
xor U6883 (N_6883,N_6179,N_6335);
nand U6884 (N_6884,N_6048,N_6063);
nand U6885 (N_6885,N_6122,N_6312);
nor U6886 (N_6886,N_6421,N_6322);
xor U6887 (N_6887,N_6215,N_6402);
or U6888 (N_6888,N_6520,N_6258);
and U6889 (N_6889,N_6251,N_6409);
xnor U6890 (N_6890,N_6172,N_6471);
nand U6891 (N_6891,N_6125,N_6133);
nand U6892 (N_6892,N_6369,N_6591);
and U6893 (N_6893,N_6440,N_6077);
nand U6894 (N_6894,N_6002,N_6110);
and U6895 (N_6895,N_6177,N_6126);
and U6896 (N_6896,N_6243,N_6362);
and U6897 (N_6897,N_6523,N_6008);
nor U6898 (N_6898,N_6192,N_6035);
nand U6899 (N_6899,N_6084,N_6017);
nand U6900 (N_6900,N_6051,N_6507);
and U6901 (N_6901,N_6444,N_6397);
and U6902 (N_6902,N_6275,N_6269);
or U6903 (N_6903,N_6061,N_6374);
nor U6904 (N_6904,N_6033,N_6506);
nand U6905 (N_6905,N_6158,N_6276);
nand U6906 (N_6906,N_6001,N_6055);
nand U6907 (N_6907,N_6550,N_6561);
or U6908 (N_6908,N_6044,N_6323);
or U6909 (N_6909,N_6401,N_6042);
nand U6910 (N_6910,N_6507,N_6578);
and U6911 (N_6911,N_6263,N_6108);
nor U6912 (N_6912,N_6517,N_6091);
or U6913 (N_6913,N_6530,N_6545);
nand U6914 (N_6914,N_6004,N_6143);
nor U6915 (N_6915,N_6145,N_6576);
xor U6916 (N_6916,N_6150,N_6198);
xor U6917 (N_6917,N_6050,N_6241);
or U6918 (N_6918,N_6530,N_6137);
xnor U6919 (N_6919,N_6409,N_6271);
or U6920 (N_6920,N_6553,N_6112);
or U6921 (N_6921,N_6319,N_6401);
nor U6922 (N_6922,N_6274,N_6169);
xor U6923 (N_6923,N_6006,N_6578);
and U6924 (N_6924,N_6390,N_6111);
nor U6925 (N_6925,N_6408,N_6447);
and U6926 (N_6926,N_6130,N_6251);
and U6927 (N_6927,N_6580,N_6567);
or U6928 (N_6928,N_6303,N_6099);
nor U6929 (N_6929,N_6376,N_6375);
nand U6930 (N_6930,N_6252,N_6286);
or U6931 (N_6931,N_6014,N_6445);
or U6932 (N_6932,N_6340,N_6025);
nand U6933 (N_6933,N_6503,N_6046);
nand U6934 (N_6934,N_6447,N_6094);
xor U6935 (N_6935,N_6457,N_6168);
and U6936 (N_6936,N_6265,N_6460);
and U6937 (N_6937,N_6183,N_6392);
nand U6938 (N_6938,N_6441,N_6431);
or U6939 (N_6939,N_6107,N_6068);
or U6940 (N_6940,N_6196,N_6556);
or U6941 (N_6941,N_6306,N_6243);
nor U6942 (N_6942,N_6027,N_6086);
or U6943 (N_6943,N_6592,N_6316);
xor U6944 (N_6944,N_6518,N_6163);
or U6945 (N_6945,N_6551,N_6170);
nor U6946 (N_6946,N_6213,N_6377);
nand U6947 (N_6947,N_6065,N_6445);
nand U6948 (N_6948,N_6436,N_6079);
nand U6949 (N_6949,N_6489,N_6044);
nand U6950 (N_6950,N_6201,N_6091);
or U6951 (N_6951,N_6589,N_6322);
nand U6952 (N_6952,N_6305,N_6517);
or U6953 (N_6953,N_6070,N_6578);
xnor U6954 (N_6954,N_6427,N_6132);
nand U6955 (N_6955,N_6105,N_6599);
nand U6956 (N_6956,N_6297,N_6061);
xor U6957 (N_6957,N_6593,N_6346);
and U6958 (N_6958,N_6495,N_6462);
and U6959 (N_6959,N_6025,N_6405);
nor U6960 (N_6960,N_6431,N_6021);
nand U6961 (N_6961,N_6204,N_6044);
xor U6962 (N_6962,N_6570,N_6539);
xnor U6963 (N_6963,N_6394,N_6148);
or U6964 (N_6964,N_6309,N_6553);
or U6965 (N_6965,N_6484,N_6220);
and U6966 (N_6966,N_6567,N_6193);
nor U6967 (N_6967,N_6169,N_6582);
or U6968 (N_6968,N_6417,N_6255);
or U6969 (N_6969,N_6458,N_6539);
or U6970 (N_6970,N_6250,N_6079);
and U6971 (N_6971,N_6492,N_6553);
and U6972 (N_6972,N_6014,N_6324);
or U6973 (N_6973,N_6598,N_6474);
and U6974 (N_6974,N_6329,N_6003);
or U6975 (N_6975,N_6403,N_6107);
nor U6976 (N_6976,N_6427,N_6443);
and U6977 (N_6977,N_6243,N_6056);
nand U6978 (N_6978,N_6427,N_6174);
and U6979 (N_6979,N_6082,N_6275);
or U6980 (N_6980,N_6225,N_6338);
or U6981 (N_6981,N_6500,N_6494);
xor U6982 (N_6982,N_6081,N_6319);
xor U6983 (N_6983,N_6008,N_6128);
xor U6984 (N_6984,N_6446,N_6033);
or U6985 (N_6985,N_6286,N_6076);
nand U6986 (N_6986,N_6029,N_6382);
nor U6987 (N_6987,N_6277,N_6052);
or U6988 (N_6988,N_6563,N_6241);
or U6989 (N_6989,N_6194,N_6186);
xor U6990 (N_6990,N_6441,N_6188);
nand U6991 (N_6991,N_6586,N_6541);
nor U6992 (N_6992,N_6308,N_6026);
nand U6993 (N_6993,N_6443,N_6402);
and U6994 (N_6994,N_6009,N_6446);
or U6995 (N_6995,N_6302,N_6070);
or U6996 (N_6996,N_6069,N_6076);
xor U6997 (N_6997,N_6228,N_6001);
or U6998 (N_6998,N_6362,N_6128);
xnor U6999 (N_6999,N_6533,N_6004);
xnor U7000 (N_7000,N_6538,N_6037);
nand U7001 (N_7001,N_6196,N_6314);
nand U7002 (N_7002,N_6551,N_6068);
or U7003 (N_7003,N_6131,N_6180);
and U7004 (N_7004,N_6002,N_6584);
nor U7005 (N_7005,N_6406,N_6155);
nor U7006 (N_7006,N_6165,N_6499);
xnor U7007 (N_7007,N_6583,N_6111);
or U7008 (N_7008,N_6233,N_6088);
xor U7009 (N_7009,N_6019,N_6409);
nand U7010 (N_7010,N_6055,N_6284);
nand U7011 (N_7011,N_6410,N_6477);
xnor U7012 (N_7012,N_6478,N_6068);
and U7013 (N_7013,N_6164,N_6239);
nor U7014 (N_7014,N_6076,N_6445);
or U7015 (N_7015,N_6375,N_6231);
nor U7016 (N_7016,N_6440,N_6524);
xnor U7017 (N_7017,N_6106,N_6067);
nor U7018 (N_7018,N_6347,N_6325);
or U7019 (N_7019,N_6411,N_6433);
and U7020 (N_7020,N_6452,N_6289);
nand U7021 (N_7021,N_6503,N_6231);
nand U7022 (N_7022,N_6406,N_6366);
and U7023 (N_7023,N_6432,N_6426);
or U7024 (N_7024,N_6182,N_6480);
nand U7025 (N_7025,N_6433,N_6362);
nor U7026 (N_7026,N_6572,N_6338);
nand U7027 (N_7027,N_6393,N_6001);
and U7028 (N_7028,N_6344,N_6033);
nand U7029 (N_7029,N_6104,N_6397);
and U7030 (N_7030,N_6177,N_6373);
nor U7031 (N_7031,N_6470,N_6360);
or U7032 (N_7032,N_6013,N_6359);
xnor U7033 (N_7033,N_6163,N_6169);
or U7034 (N_7034,N_6030,N_6193);
xor U7035 (N_7035,N_6579,N_6389);
xnor U7036 (N_7036,N_6049,N_6434);
nand U7037 (N_7037,N_6137,N_6182);
xnor U7038 (N_7038,N_6362,N_6164);
nor U7039 (N_7039,N_6564,N_6477);
xnor U7040 (N_7040,N_6211,N_6277);
xor U7041 (N_7041,N_6067,N_6547);
nand U7042 (N_7042,N_6254,N_6093);
and U7043 (N_7043,N_6382,N_6318);
xor U7044 (N_7044,N_6336,N_6394);
nand U7045 (N_7045,N_6341,N_6096);
or U7046 (N_7046,N_6492,N_6165);
nor U7047 (N_7047,N_6042,N_6163);
or U7048 (N_7048,N_6447,N_6100);
xnor U7049 (N_7049,N_6151,N_6011);
nor U7050 (N_7050,N_6529,N_6032);
and U7051 (N_7051,N_6405,N_6581);
and U7052 (N_7052,N_6273,N_6400);
and U7053 (N_7053,N_6132,N_6224);
or U7054 (N_7054,N_6262,N_6476);
and U7055 (N_7055,N_6157,N_6016);
xor U7056 (N_7056,N_6027,N_6152);
or U7057 (N_7057,N_6544,N_6033);
and U7058 (N_7058,N_6140,N_6477);
or U7059 (N_7059,N_6531,N_6236);
or U7060 (N_7060,N_6401,N_6131);
nor U7061 (N_7061,N_6056,N_6312);
xor U7062 (N_7062,N_6518,N_6175);
and U7063 (N_7063,N_6127,N_6189);
and U7064 (N_7064,N_6453,N_6170);
nor U7065 (N_7065,N_6439,N_6421);
nand U7066 (N_7066,N_6132,N_6293);
nand U7067 (N_7067,N_6490,N_6107);
or U7068 (N_7068,N_6366,N_6599);
nand U7069 (N_7069,N_6330,N_6413);
or U7070 (N_7070,N_6213,N_6293);
nor U7071 (N_7071,N_6370,N_6331);
and U7072 (N_7072,N_6106,N_6179);
xnor U7073 (N_7073,N_6214,N_6436);
or U7074 (N_7074,N_6297,N_6353);
or U7075 (N_7075,N_6345,N_6056);
nor U7076 (N_7076,N_6588,N_6076);
nor U7077 (N_7077,N_6097,N_6333);
xor U7078 (N_7078,N_6304,N_6102);
and U7079 (N_7079,N_6564,N_6066);
xnor U7080 (N_7080,N_6545,N_6291);
and U7081 (N_7081,N_6479,N_6061);
nand U7082 (N_7082,N_6531,N_6002);
or U7083 (N_7083,N_6312,N_6404);
and U7084 (N_7084,N_6529,N_6152);
nand U7085 (N_7085,N_6168,N_6173);
nor U7086 (N_7086,N_6373,N_6016);
nand U7087 (N_7087,N_6308,N_6000);
or U7088 (N_7088,N_6246,N_6533);
nand U7089 (N_7089,N_6267,N_6120);
nor U7090 (N_7090,N_6501,N_6077);
nand U7091 (N_7091,N_6434,N_6134);
nor U7092 (N_7092,N_6265,N_6464);
xor U7093 (N_7093,N_6318,N_6055);
or U7094 (N_7094,N_6599,N_6462);
xnor U7095 (N_7095,N_6023,N_6523);
xnor U7096 (N_7096,N_6165,N_6156);
and U7097 (N_7097,N_6579,N_6386);
or U7098 (N_7098,N_6111,N_6096);
and U7099 (N_7099,N_6541,N_6158);
xnor U7100 (N_7100,N_6261,N_6012);
nor U7101 (N_7101,N_6195,N_6385);
nor U7102 (N_7102,N_6440,N_6320);
or U7103 (N_7103,N_6419,N_6207);
xor U7104 (N_7104,N_6189,N_6495);
or U7105 (N_7105,N_6017,N_6410);
xor U7106 (N_7106,N_6215,N_6092);
and U7107 (N_7107,N_6563,N_6393);
xnor U7108 (N_7108,N_6571,N_6047);
xnor U7109 (N_7109,N_6080,N_6085);
xor U7110 (N_7110,N_6415,N_6571);
xnor U7111 (N_7111,N_6383,N_6525);
or U7112 (N_7112,N_6550,N_6449);
nor U7113 (N_7113,N_6097,N_6564);
nor U7114 (N_7114,N_6063,N_6068);
xnor U7115 (N_7115,N_6284,N_6040);
nor U7116 (N_7116,N_6099,N_6095);
and U7117 (N_7117,N_6495,N_6226);
nor U7118 (N_7118,N_6241,N_6110);
or U7119 (N_7119,N_6067,N_6040);
nand U7120 (N_7120,N_6526,N_6490);
nor U7121 (N_7121,N_6517,N_6076);
nor U7122 (N_7122,N_6375,N_6046);
and U7123 (N_7123,N_6113,N_6013);
xnor U7124 (N_7124,N_6453,N_6213);
nor U7125 (N_7125,N_6490,N_6528);
nand U7126 (N_7126,N_6039,N_6121);
nand U7127 (N_7127,N_6179,N_6508);
xor U7128 (N_7128,N_6178,N_6153);
nor U7129 (N_7129,N_6451,N_6173);
xor U7130 (N_7130,N_6472,N_6195);
nand U7131 (N_7131,N_6575,N_6559);
xnor U7132 (N_7132,N_6387,N_6260);
nor U7133 (N_7133,N_6550,N_6521);
xnor U7134 (N_7134,N_6549,N_6170);
nand U7135 (N_7135,N_6528,N_6026);
nand U7136 (N_7136,N_6429,N_6058);
nand U7137 (N_7137,N_6058,N_6407);
nand U7138 (N_7138,N_6590,N_6224);
nor U7139 (N_7139,N_6287,N_6276);
nor U7140 (N_7140,N_6226,N_6167);
and U7141 (N_7141,N_6025,N_6546);
and U7142 (N_7142,N_6564,N_6227);
nand U7143 (N_7143,N_6116,N_6069);
xnor U7144 (N_7144,N_6391,N_6280);
or U7145 (N_7145,N_6597,N_6403);
nand U7146 (N_7146,N_6437,N_6136);
nand U7147 (N_7147,N_6247,N_6285);
or U7148 (N_7148,N_6104,N_6535);
xor U7149 (N_7149,N_6484,N_6117);
nand U7150 (N_7150,N_6437,N_6078);
xnor U7151 (N_7151,N_6244,N_6327);
nor U7152 (N_7152,N_6594,N_6518);
or U7153 (N_7153,N_6045,N_6500);
or U7154 (N_7154,N_6376,N_6468);
or U7155 (N_7155,N_6554,N_6198);
or U7156 (N_7156,N_6541,N_6019);
and U7157 (N_7157,N_6327,N_6361);
and U7158 (N_7158,N_6010,N_6103);
xnor U7159 (N_7159,N_6495,N_6301);
nor U7160 (N_7160,N_6104,N_6213);
or U7161 (N_7161,N_6523,N_6152);
nand U7162 (N_7162,N_6100,N_6360);
or U7163 (N_7163,N_6413,N_6227);
or U7164 (N_7164,N_6590,N_6016);
nand U7165 (N_7165,N_6305,N_6218);
xor U7166 (N_7166,N_6148,N_6125);
nor U7167 (N_7167,N_6312,N_6053);
nand U7168 (N_7168,N_6305,N_6450);
and U7169 (N_7169,N_6203,N_6320);
nand U7170 (N_7170,N_6072,N_6048);
and U7171 (N_7171,N_6163,N_6296);
nand U7172 (N_7172,N_6202,N_6417);
nand U7173 (N_7173,N_6572,N_6349);
xnor U7174 (N_7174,N_6448,N_6199);
nand U7175 (N_7175,N_6067,N_6519);
and U7176 (N_7176,N_6467,N_6329);
nor U7177 (N_7177,N_6141,N_6122);
and U7178 (N_7178,N_6422,N_6184);
and U7179 (N_7179,N_6507,N_6130);
nand U7180 (N_7180,N_6456,N_6413);
nand U7181 (N_7181,N_6402,N_6563);
nor U7182 (N_7182,N_6093,N_6365);
nor U7183 (N_7183,N_6459,N_6115);
xor U7184 (N_7184,N_6294,N_6058);
nor U7185 (N_7185,N_6228,N_6072);
nor U7186 (N_7186,N_6114,N_6546);
or U7187 (N_7187,N_6380,N_6336);
nand U7188 (N_7188,N_6093,N_6210);
nor U7189 (N_7189,N_6154,N_6013);
or U7190 (N_7190,N_6157,N_6290);
and U7191 (N_7191,N_6468,N_6467);
xnor U7192 (N_7192,N_6287,N_6505);
and U7193 (N_7193,N_6303,N_6336);
xor U7194 (N_7194,N_6209,N_6516);
and U7195 (N_7195,N_6545,N_6492);
nand U7196 (N_7196,N_6391,N_6555);
xnor U7197 (N_7197,N_6328,N_6177);
nor U7198 (N_7198,N_6249,N_6446);
xor U7199 (N_7199,N_6012,N_6219);
nand U7200 (N_7200,N_6946,N_7045);
nor U7201 (N_7201,N_7028,N_6862);
or U7202 (N_7202,N_7163,N_6774);
nand U7203 (N_7203,N_6863,N_6827);
nor U7204 (N_7204,N_6758,N_7162);
and U7205 (N_7205,N_6711,N_6934);
nor U7206 (N_7206,N_6983,N_6633);
nor U7207 (N_7207,N_6620,N_6852);
nor U7208 (N_7208,N_6709,N_7038);
and U7209 (N_7209,N_6676,N_7123);
nor U7210 (N_7210,N_7059,N_7104);
nand U7211 (N_7211,N_7047,N_6624);
nor U7212 (N_7212,N_7125,N_6692);
and U7213 (N_7213,N_7141,N_6656);
nand U7214 (N_7214,N_6646,N_6634);
xnor U7215 (N_7215,N_6981,N_6700);
nand U7216 (N_7216,N_6749,N_6641);
and U7217 (N_7217,N_6752,N_7121);
nor U7218 (N_7218,N_7090,N_6955);
nand U7219 (N_7219,N_7084,N_7132);
nand U7220 (N_7220,N_7102,N_6608);
and U7221 (N_7221,N_6887,N_7051);
xor U7222 (N_7222,N_6655,N_7099);
nand U7223 (N_7223,N_6777,N_7057);
or U7224 (N_7224,N_6923,N_6738);
xor U7225 (N_7225,N_7067,N_7020);
nor U7226 (N_7226,N_6773,N_7147);
or U7227 (N_7227,N_6844,N_6786);
or U7228 (N_7228,N_6917,N_6623);
and U7229 (N_7229,N_6720,N_6658);
or U7230 (N_7230,N_7170,N_6654);
nand U7231 (N_7231,N_6684,N_7120);
nor U7232 (N_7232,N_7189,N_6898);
nor U7233 (N_7233,N_6739,N_6632);
xor U7234 (N_7234,N_6732,N_6926);
and U7235 (N_7235,N_6896,N_6978);
nor U7236 (N_7236,N_7027,N_6859);
xor U7237 (N_7237,N_6878,N_6638);
or U7238 (N_7238,N_6816,N_7004);
xnor U7239 (N_7239,N_6838,N_7173);
xnor U7240 (N_7240,N_6733,N_7142);
or U7241 (N_7241,N_6699,N_7043);
and U7242 (N_7242,N_7075,N_6947);
and U7243 (N_7243,N_6682,N_7136);
and U7244 (N_7244,N_6802,N_6919);
or U7245 (N_7245,N_7165,N_7191);
nand U7246 (N_7246,N_6832,N_7088);
or U7247 (N_7247,N_6845,N_6997);
or U7248 (N_7248,N_6937,N_6693);
nor U7249 (N_7249,N_7113,N_7093);
and U7250 (N_7250,N_6856,N_6755);
nor U7251 (N_7251,N_7100,N_6621);
or U7252 (N_7252,N_6822,N_6872);
xor U7253 (N_7253,N_6931,N_7145);
xor U7254 (N_7254,N_7195,N_6695);
xnor U7255 (N_7255,N_6913,N_6730);
or U7256 (N_7256,N_7111,N_6979);
nor U7257 (N_7257,N_6938,N_7155);
or U7258 (N_7258,N_7172,N_6835);
or U7259 (N_7259,N_6980,N_6817);
xnor U7260 (N_7260,N_6971,N_7044);
or U7261 (N_7261,N_6957,N_7101);
xor U7262 (N_7262,N_6890,N_7112);
xnor U7263 (N_7263,N_7107,N_7146);
nand U7264 (N_7264,N_6895,N_7109);
xor U7265 (N_7265,N_7082,N_6820);
nor U7266 (N_7266,N_7074,N_6814);
and U7267 (N_7267,N_7159,N_6953);
nand U7268 (N_7268,N_7114,N_6746);
nor U7269 (N_7269,N_6678,N_6653);
nand U7270 (N_7270,N_6831,N_6799);
nor U7271 (N_7271,N_7068,N_6761);
and U7272 (N_7272,N_6804,N_6977);
and U7273 (N_7273,N_6716,N_6668);
and U7274 (N_7274,N_6609,N_7106);
and U7275 (N_7275,N_6771,N_6905);
xor U7276 (N_7276,N_7143,N_7181);
nor U7277 (N_7277,N_6885,N_6741);
xnor U7278 (N_7278,N_6629,N_6750);
xor U7279 (N_7279,N_7009,N_7193);
nand U7280 (N_7280,N_6706,N_7118);
or U7281 (N_7281,N_7160,N_6687);
and U7282 (N_7282,N_6839,N_7087);
nand U7283 (N_7283,N_6944,N_6973);
or U7284 (N_7284,N_6858,N_6778);
and U7285 (N_7285,N_6652,N_6787);
or U7286 (N_7286,N_6677,N_6604);
xnor U7287 (N_7287,N_7052,N_7169);
xnor U7288 (N_7288,N_6651,N_6949);
or U7289 (N_7289,N_7115,N_7000);
or U7290 (N_7290,N_6707,N_6660);
nor U7291 (N_7291,N_7003,N_6736);
and U7292 (N_7292,N_6690,N_6779);
and U7293 (N_7293,N_6769,N_6941);
nor U7294 (N_7294,N_6861,N_6866);
nor U7295 (N_7295,N_6968,N_6994);
or U7296 (N_7296,N_6962,N_6970);
nor U7297 (N_7297,N_6770,N_7072);
and U7298 (N_7298,N_6921,N_6734);
nand U7299 (N_7299,N_7137,N_6826);
nor U7300 (N_7300,N_6795,N_6959);
nor U7301 (N_7301,N_7103,N_7190);
xnor U7302 (N_7302,N_6728,N_7161);
nand U7303 (N_7303,N_6891,N_7133);
and U7304 (N_7304,N_6754,N_6909);
or U7305 (N_7305,N_6837,N_7025);
or U7306 (N_7306,N_6631,N_7058);
nand U7307 (N_7307,N_6600,N_7148);
or U7308 (N_7308,N_6672,N_6897);
and U7309 (N_7309,N_7151,N_6607);
xor U7310 (N_7310,N_6829,N_7174);
and U7311 (N_7311,N_7022,N_7012);
and U7312 (N_7312,N_6875,N_7157);
and U7313 (N_7313,N_7117,N_6922);
and U7314 (N_7314,N_6836,N_7071);
or U7315 (N_7315,N_7154,N_6616);
and U7316 (N_7316,N_6650,N_7122);
and U7317 (N_7317,N_6849,N_7186);
nand U7318 (N_7318,N_6731,N_6904);
xor U7319 (N_7319,N_6911,N_7036);
or U7320 (N_7320,N_6993,N_6663);
and U7321 (N_7321,N_6960,N_6988);
nand U7322 (N_7322,N_6865,N_6803);
xor U7323 (N_7323,N_6943,N_6847);
nor U7324 (N_7324,N_6703,N_6864);
nand U7325 (N_7325,N_6880,N_6869);
nand U7326 (N_7326,N_7158,N_6918);
or U7327 (N_7327,N_6940,N_6712);
nand U7328 (N_7328,N_7001,N_6791);
nor U7329 (N_7329,N_6906,N_7076);
nand U7330 (N_7330,N_6657,N_7080);
xnor U7331 (N_7331,N_6942,N_6644);
and U7332 (N_7332,N_6744,N_7180);
nand U7333 (N_7333,N_6810,N_7070);
nand U7334 (N_7334,N_7124,N_6742);
nand U7335 (N_7335,N_6694,N_7056);
xnor U7336 (N_7336,N_6722,N_6920);
or U7337 (N_7337,N_6763,N_7199);
or U7338 (N_7338,N_7039,N_7185);
nor U7339 (N_7339,N_6721,N_6789);
or U7340 (N_7340,N_7017,N_7183);
xnor U7341 (N_7341,N_7184,N_7086);
or U7342 (N_7342,N_6902,N_7131);
nor U7343 (N_7343,N_7006,N_6719);
nand U7344 (N_7344,N_6606,N_6662);
nor U7345 (N_7345,N_6637,N_6884);
and U7346 (N_7346,N_6757,N_6765);
xor U7347 (N_7347,N_7105,N_6785);
or U7348 (N_7348,N_7062,N_6661);
nor U7349 (N_7349,N_7040,N_6797);
or U7350 (N_7350,N_7171,N_6982);
nand U7351 (N_7351,N_6882,N_6740);
and U7352 (N_7352,N_6818,N_6669);
and U7353 (N_7353,N_6975,N_6648);
nand U7354 (N_7354,N_7061,N_6883);
xnor U7355 (N_7355,N_7066,N_6627);
or U7356 (N_7356,N_6821,N_6927);
nand U7357 (N_7357,N_6998,N_6685);
or U7358 (N_7358,N_6751,N_6974);
xor U7359 (N_7359,N_6670,N_6965);
nor U7360 (N_7360,N_7008,N_6612);
nor U7361 (N_7361,N_6850,N_7015);
or U7362 (N_7362,N_7069,N_6893);
nor U7363 (N_7363,N_6701,N_6747);
and U7364 (N_7364,N_6870,N_6647);
nand U7365 (N_7365,N_6665,N_7188);
or U7366 (N_7366,N_6686,N_6729);
or U7367 (N_7367,N_6928,N_7144);
nor U7368 (N_7368,N_6914,N_7127);
and U7369 (N_7369,N_7194,N_7005);
nor U7370 (N_7370,N_6659,N_7098);
nand U7371 (N_7371,N_6886,N_7096);
or U7372 (N_7372,N_7153,N_6824);
xnor U7373 (N_7373,N_7033,N_7023);
or U7374 (N_7374,N_6881,N_6915);
nand U7375 (N_7375,N_6945,N_6848);
or U7376 (N_7376,N_6679,N_7149);
nor U7377 (N_7377,N_6907,N_7034);
and U7378 (N_7378,N_6666,N_6900);
nor U7379 (N_7379,N_7156,N_6833);
nand U7380 (N_7380,N_6996,N_7197);
and U7381 (N_7381,N_6995,N_6723);
or U7382 (N_7382,N_6625,N_6782);
and U7383 (N_7383,N_6759,N_6892);
nor U7384 (N_7384,N_6984,N_7007);
nand U7385 (N_7385,N_6807,N_7150);
or U7386 (N_7386,N_7063,N_6801);
xnor U7387 (N_7387,N_7091,N_6614);
and U7388 (N_7388,N_7094,N_7013);
or U7389 (N_7389,N_7073,N_6969);
and U7390 (N_7390,N_6640,N_6748);
and U7391 (N_7391,N_6718,N_7192);
and U7392 (N_7392,N_7175,N_6708);
nand U7393 (N_7393,N_7018,N_6991);
nand U7394 (N_7394,N_6874,N_6674);
or U7395 (N_7395,N_6813,N_6717);
xnor U7396 (N_7396,N_6626,N_6756);
nand U7397 (N_7397,N_7178,N_6780);
and U7398 (N_7398,N_6854,N_6675);
or U7399 (N_7399,N_6841,N_6617);
xnor U7400 (N_7400,N_6930,N_6846);
nor U7401 (N_7401,N_6806,N_6793);
nand U7402 (N_7402,N_6691,N_7064);
or U7403 (N_7403,N_7032,N_6743);
and U7404 (N_7404,N_6794,N_6636);
or U7405 (N_7405,N_6696,N_7060);
xnor U7406 (N_7406,N_6689,N_7026);
nor U7407 (N_7407,N_6908,N_6933);
nor U7408 (N_7408,N_6956,N_6815);
xnor U7409 (N_7409,N_6857,N_7077);
or U7410 (N_7410,N_6727,N_6783);
or U7411 (N_7411,N_6760,N_7139);
nor U7412 (N_7412,N_6924,N_6990);
nand U7413 (N_7413,N_7029,N_6985);
or U7414 (N_7414,N_6705,N_7152);
xor U7415 (N_7415,N_7024,N_7042);
and U7416 (N_7416,N_7092,N_6868);
nand U7417 (N_7417,N_6936,N_7048);
nor U7418 (N_7418,N_7010,N_6992);
xor U7419 (N_7419,N_6715,N_6673);
xor U7420 (N_7420,N_6961,N_6999);
and U7421 (N_7421,N_7083,N_6951);
nand U7422 (N_7422,N_6966,N_7097);
xnor U7423 (N_7423,N_6828,N_6967);
nand U7424 (N_7424,N_6776,N_6639);
or U7425 (N_7425,N_7110,N_7081);
and U7426 (N_7426,N_6851,N_6910);
and U7427 (N_7427,N_6950,N_6681);
xnor U7428 (N_7428,N_6618,N_6989);
xor U7429 (N_7429,N_7079,N_6688);
and U7430 (N_7430,N_7016,N_6860);
nand U7431 (N_7431,N_7164,N_7095);
nand U7432 (N_7432,N_6808,N_6610);
or U7433 (N_7433,N_6710,N_6903);
nor U7434 (N_7434,N_6683,N_6843);
or U7435 (N_7435,N_6671,N_6842);
nor U7436 (N_7436,N_6876,N_6792);
nand U7437 (N_7437,N_6735,N_7054);
and U7438 (N_7438,N_6935,N_6830);
or U7439 (N_7439,N_6901,N_6867);
nor U7440 (N_7440,N_7166,N_7053);
and U7441 (N_7441,N_7130,N_6798);
and U7442 (N_7442,N_6963,N_7196);
nor U7443 (N_7443,N_6645,N_6805);
nor U7444 (N_7444,N_7135,N_7065);
nor U7445 (N_7445,N_6768,N_7014);
xor U7446 (N_7446,N_6800,N_7176);
and U7447 (N_7447,N_6766,N_6745);
or U7448 (N_7448,N_7041,N_6767);
nor U7449 (N_7449,N_6879,N_6615);
nor U7450 (N_7450,N_7168,N_6812);
or U7451 (N_7451,N_7019,N_6958);
nor U7452 (N_7452,N_6784,N_6916);
or U7453 (N_7453,N_6811,N_6976);
or U7454 (N_7454,N_7085,N_6772);
or U7455 (N_7455,N_6954,N_6899);
and U7456 (N_7456,N_7108,N_6932);
and U7457 (N_7457,N_7179,N_7129);
and U7458 (N_7458,N_7030,N_6877);
and U7459 (N_7459,N_7035,N_6964);
nor U7460 (N_7460,N_6764,N_6698);
nand U7461 (N_7461,N_7177,N_6889);
and U7462 (N_7462,N_6667,N_6605);
nor U7463 (N_7463,N_7167,N_7128);
nor U7464 (N_7464,N_6725,N_6601);
xnor U7465 (N_7465,N_6834,N_6788);
xnor U7466 (N_7466,N_6713,N_7138);
and U7467 (N_7467,N_7049,N_6929);
xnor U7468 (N_7468,N_6737,N_7046);
and U7469 (N_7469,N_6888,N_6664);
or U7470 (N_7470,N_6628,N_6611);
nand U7471 (N_7471,N_6855,N_6972);
and U7472 (N_7472,N_6622,N_6819);
or U7473 (N_7473,N_6613,N_6726);
nand U7474 (N_7474,N_6986,N_7037);
xor U7475 (N_7475,N_6823,N_6714);
nand U7476 (N_7476,N_6952,N_7126);
and U7477 (N_7477,N_7011,N_6948);
or U7478 (N_7478,N_7002,N_7140);
xor U7479 (N_7479,N_6649,N_6894);
and U7480 (N_7480,N_7078,N_6602);
nand U7481 (N_7481,N_6825,N_6724);
xnor U7482 (N_7482,N_6809,N_6987);
and U7483 (N_7483,N_6642,N_6912);
nor U7484 (N_7484,N_6925,N_6704);
nor U7485 (N_7485,N_7134,N_6939);
xor U7486 (N_7486,N_6702,N_6775);
xor U7487 (N_7487,N_6680,N_7187);
nor U7488 (N_7488,N_6790,N_7116);
nor U7489 (N_7489,N_6762,N_7089);
or U7490 (N_7490,N_6840,N_6753);
nand U7491 (N_7491,N_7055,N_6796);
and U7492 (N_7492,N_7198,N_6873);
nor U7493 (N_7493,N_6619,N_7050);
and U7494 (N_7494,N_6853,N_7182);
and U7495 (N_7495,N_6643,N_7021);
nand U7496 (N_7496,N_6635,N_7031);
or U7497 (N_7497,N_6630,N_6871);
nor U7498 (N_7498,N_6697,N_6781);
nor U7499 (N_7499,N_7119,N_6603);
xor U7500 (N_7500,N_7000,N_7175);
nand U7501 (N_7501,N_6888,N_6615);
and U7502 (N_7502,N_7079,N_6683);
xor U7503 (N_7503,N_6782,N_6793);
and U7504 (N_7504,N_7129,N_7144);
nor U7505 (N_7505,N_7138,N_6927);
nand U7506 (N_7506,N_7026,N_6869);
and U7507 (N_7507,N_7014,N_6790);
nor U7508 (N_7508,N_6806,N_6624);
and U7509 (N_7509,N_6611,N_6982);
nor U7510 (N_7510,N_7088,N_7096);
nand U7511 (N_7511,N_7131,N_6712);
nor U7512 (N_7512,N_6874,N_6602);
nor U7513 (N_7513,N_6998,N_6646);
and U7514 (N_7514,N_6763,N_6983);
xor U7515 (N_7515,N_6608,N_6943);
or U7516 (N_7516,N_6843,N_7147);
nor U7517 (N_7517,N_7118,N_6635);
or U7518 (N_7518,N_6959,N_7058);
nand U7519 (N_7519,N_6612,N_7186);
nor U7520 (N_7520,N_6780,N_6737);
nor U7521 (N_7521,N_7103,N_7044);
nand U7522 (N_7522,N_7130,N_6762);
and U7523 (N_7523,N_7040,N_7128);
nor U7524 (N_7524,N_6798,N_7025);
nand U7525 (N_7525,N_6758,N_6805);
xnor U7526 (N_7526,N_6922,N_6908);
or U7527 (N_7527,N_7146,N_6698);
and U7528 (N_7528,N_6697,N_7010);
or U7529 (N_7529,N_6704,N_6710);
nand U7530 (N_7530,N_6739,N_6761);
nor U7531 (N_7531,N_6815,N_7049);
nor U7532 (N_7532,N_6804,N_6648);
nor U7533 (N_7533,N_6648,N_6990);
nor U7534 (N_7534,N_6819,N_6817);
xnor U7535 (N_7535,N_6943,N_6780);
xor U7536 (N_7536,N_7071,N_6816);
nand U7537 (N_7537,N_6636,N_6660);
xnor U7538 (N_7538,N_6993,N_6858);
nor U7539 (N_7539,N_7170,N_6812);
xor U7540 (N_7540,N_6812,N_6850);
xnor U7541 (N_7541,N_6945,N_6685);
nand U7542 (N_7542,N_7016,N_6661);
xor U7543 (N_7543,N_6809,N_6835);
xnor U7544 (N_7544,N_7101,N_6888);
xnor U7545 (N_7545,N_6839,N_6658);
xnor U7546 (N_7546,N_6743,N_6807);
xor U7547 (N_7547,N_6863,N_7162);
or U7548 (N_7548,N_6988,N_7128);
nand U7549 (N_7549,N_6751,N_6989);
nand U7550 (N_7550,N_6758,N_6795);
xnor U7551 (N_7551,N_7156,N_7165);
or U7552 (N_7552,N_6981,N_6661);
nand U7553 (N_7553,N_6709,N_6877);
xor U7554 (N_7554,N_6883,N_6618);
or U7555 (N_7555,N_7179,N_6725);
or U7556 (N_7556,N_7152,N_7029);
or U7557 (N_7557,N_6925,N_6897);
nand U7558 (N_7558,N_6625,N_7071);
and U7559 (N_7559,N_6877,N_6820);
nand U7560 (N_7560,N_7166,N_6961);
nand U7561 (N_7561,N_6943,N_7061);
or U7562 (N_7562,N_6744,N_6691);
or U7563 (N_7563,N_6809,N_7166);
and U7564 (N_7564,N_6620,N_7192);
nand U7565 (N_7565,N_6927,N_6754);
nor U7566 (N_7566,N_7172,N_6759);
and U7567 (N_7567,N_6783,N_7044);
xnor U7568 (N_7568,N_6688,N_6678);
xor U7569 (N_7569,N_6960,N_6727);
and U7570 (N_7570,N_7066,N_6962);
nor U7571 (N_7571,N_7026,N_6832);
or U7572 (N_7572,N_7138,N_7154);
and U7573 (N_7573,N_6837,N_7077);
xnor U7574 (N_7574,N_6769,N_6609);
xnor U7575 (N_7575,N_6601,N_7041);
nor U7576 (N_7576,N_7134,N_6897);
xor U7577 (N_7577,N_6746,N_6650);
and U7578 (N_7578,N_6824,N_6657);
nor U7579 (N_7579,N_6875,N_6907);
nand U7580 (N_7580,N_7144,N_6995);
or U7581 (N_7581,N_6871,N_7160);
xnor U7582 (N_7582,N_6771,N_7091);
nand U7583 (N_7583,N_7067,N_6761);
xor U7584 (N_7584,N_6811,N_6924);
nand U7585 (N_7585,N_6711,N_7194);
xnor U7586 (N_7586,N_7173,N_6942);
xor U7587 (N_7587,N_6781,N_6821);
xnor U7588 (N_7588,N_7119,N_6609);
and U7589 (N_7589,N_6660,N_7009);
and U7590 (N_7590,N_7094,N_6670);
nand U7591 (N_7591,N_6783,N_6717);
and U7592 (N_7592,N_7144,N_6827);
nor U7593 (N_7593,N_7173,N_6705);
and U7594 (N_7594,N_6992,N_6733);
xnor U7595 (N_7595,N_6706,N_7023);
nor U7596 (N_7596,N_6769,N_6974);
or U7597 (N_7597,N_6950,N_7002);
or U7598 (N_7598,N_6775,N_7194);
nor U7599 (N_7599,N_7176,N_6872);
xnor U7600 (N_7600,N_6970,N_6915);
and U7601 (N_7601,N_6969,N_6774);
xnor U7602 (N_7602,N_7186,N_7136);
nand U7603 (N_7603,N_6684,N_7008);
or U7604 (N_7604,N_6835,N_6816);
and U7605 (N_7605,N_6768,N_6712);
and U7606 (N_7606,N_6736,N_7155);
nor U7607 (N_7607,N_6830,N_7122);
xor U7608 (N_7608,N_7095,N_7160);
nor U7609 (N_7609,N_6641,N_7144);
nor U7610 (N_7610,N_6696,N_7166);
nor U7611 (N_7611,N_7038,N_6917);
and U7612 (N_7612,N_6744,N_7032);
nand U7613 (N_7613,N_7142,N_6935);
or U7614 (N_7614,N_7068,N_6888);
or U7615 (N_7615,N_6934,N_6918);
nor U7616 (N_7616,N_6971,N_7001);
and U7617 (N_7617,N_7096,N_6870);
nand U7618 (N_7618,N_6936,N_6736);
xnor U7619 (N_7619,N_6862,N_6607);
nand U7620 (N_7620,N_6972,N_6734);
nand U7621 (N_7621,N_6882,N_6635);
or U7622 (N_7622,N_7083,N_6910);
xnor U7623 (N_7623,N_7066,N_6899);
nor U7624 (N_7624,N_6601,N_6754);
nand U7625 (N_7625,N_6797,N_7114);
nand U7626 (N_7626,N_6600,N_7079);
or U7627 (N_7627,N_6998,N_7160);
nor U7628 (N_7628,N_7055,N_6768);
or U7629 (N_7629,N_6603,N_6766);
xnor U7630 (N_7630,N_7084,N_6915);
or U7631 (N_7631,N_6658,N_6641);
and U7632 (N_7632,N_6794,N_6802);
and U7633 (N_7633,N_6887,N_6774);
and U7634 (N_7634,N_6878,N_6837);
nand U7635 (N_7635,N_7053,N_7057);
and U7636 (N_7636,N_6609,N_6910);
and U7637 (N_7637,N_7071,N_6910);
and U7638 (N_7638,N_6742,N_7165);
and U7639 (N_7639,N_6994,N_6758);
nor U7640 (N_7640,N_7063,N_7018);
nor U7641 (N_7641,N_6947,N_7054);
nor U7642 (N_7642,N_7088,N_6869);
and U7643 (N_7643,N_6926,N_7168);
or U7644 (N_7644,N_6680,N_6709);
nand U7645 (N_7645,N_6953,N_6797);
nand U7646 (N_7646,N_6710,N_6717);
or U7647 (N_7647,N_6769,N_7108);
xor U7648 (N_7648,N_6911,N_6820);
nor U7649 (N_7649,N_6777,N_6789);
and U7650 (N_7650,N_6883,N_6915);
and U7651 (N_7651,N_6741,N_6839);
and U7652 (N_7652,N_6965,N_7145);
xor U7653 (N_7653,N_7101,N_7184);
nor U7654 (N_7654,N_6877,N_7055);
and U7655 (N_7655,N_6987,N_6803);
nand U7656 (N_7656,N_6902,N_6975);
xnor U7657 (N_7657,N_7196,N_6863);
nand U7658 (N_7658,N_6905,N_6946);
nand U7659 (N_7659,N_6728,N_7091);
xnor U7660 (N_7660,N_6820,N_6928);
or U7661 (N_7661,N_7036,N_6817);
and U7662 (N_7662,N_6905,N_6779);
or U7663 (N_7663,N_6809,N_7115);
or U7664 (N_7664,N_7143,N_6754);
xnor U7665 (N_7665,N_7144,N_7176);
nor U7666 (N_7666,N_6857,N_6626);
nor U7667 (N_7667,N_7107,N_7135);
or U7668 (N_7668,N_7129,N_7147);
nor U7669 (N_7669,N_6860,N_7188);
nor U7670 (N_7670,N_7032,N_6796);
and U7671 (N_7671,N_6941,N_7057);
or U7672 (N_7672,N_6780,N_6776);
xnor U7673 (N_7673,N_7064,N_7101);
and U7674 (N_7674,N_6725,N_7129);
nand U7675 (N_7675,N_7059,N_6834);
or U7676 (N_7676,N_6730,N_6626);
nand U7677 (N_7677,N_7087,N_6708);
nor U7678 (N_7678,N_6949,N_6759);
or U7679 (N_7679,N_6802,N_7064);
nand U7680 (N_7680,N_7024,N_7119);
nand U7681 (N_7681,N_6846,N_6619);
nor U7682 (N_7682,N_6844,N_6706);
nand U7683 (N_7683,N_6768,N_6667);
xor U7684 (N_7684,N_7017,N_6904);
nand U7685 (N_7685,N_7020,N_6693);
and U7686 (N_7686,N_7170,N_7011);
or U7687 (N_7687,N_6958,N_7028);
or U7688 (N_7688,N_6925,N_6968);
nor U7689 (N_7689,N_6862,N_6681);
nor U7690 (N_7690,N_6724,N_6668);
or U7691 (N_7691,N_7055,N_6939);
nand U7692 (N_7692,N_7195,N_6972);
nor U7693 (N_7693,N_7160,N_7023);
nand U7694 (N_7694,N_6651,N_6728);
nand U7695 (N_7695,N_6935,N_6901);
nand U7696 (N_7696,N_7034,N_6814);
nand U7697 (N_7697,N_6984,N_7015);
nand U7698 (N_7698,N_7008,N_7176);
xnor U7699 (N_7699,N_7164,N_7009);
nand U7700 (N_7700,N_6969,N_7032);
xor U7701 (N_7701,N_7141,N_6688);
xnor U7702 (N_7702,N_7146,N_6874);
nor U7703 (N_7703,N_6774,N_6709);
xor U7704 (N_7704,N_6960,N_6638);
nand U7705 (N_7705,N_6613,N_7160);
nor U7706 (N_7706,N_6768,N_6943);
or U7707 (N_7707,N_6692,N_7128);
nand U7708 (N_7708,N_7061,N_6789);
nand U7709 (N_7709,N_6968,N_7097);
nor U7710 (N_7710,N_6798,N_6728);
nor U7711 (N_7711,N_6732,N_6655);
nand U7712 (N_7712,N_6946,N_6760);
nand U7713 (N_7713,N_6806,N_6803);
xor U7714 (N_7714,N_7169,N_6759);
or U7715 (N_7715,N_6821,N_6848);
or U7716 (N_7716,N_7198,N_6686);
and U7717 (N_7717,N_6983,N_6909);
or U7718 (N_7718,N_6885,N_7070);
nand U7719 (N_7719,N_7143,N_6824);
nor U7720 (N_7720,N_6911,N_6761);
and U7721 (N_7721,N_7035,N_6723);
xnor U7722 (N_7722,N_7098,N_7171);
or U7723 (N_7723,N_6906,N_7149);
and U7724 (N_7724,N_6991,N_6847);
or U7725 (N_7725,N_7001,N_7168);
nand U7726 (N_7726,N_6931,N_7047);
and U7727 (N_7727,N_6832,N_6984);
nand U7728 (N_7728,N_6733,N_7086);
nand U7729 (N_7729,N_6927,N_7106);
xnor U7730 (N_7730,N_7004,N_7127);
nor U7731 (N_7731,N_7128,N_6848);
or U7732 (N_7732,N_6603,N_6858);
and U7733 (N_7733,N_7089,N_6784);
nand U7734 (N_7734,N_7155,N_7102);
nand U7735 (N_7735,N_6606,N_6962);
xor U7736 (N_7736,N_6697,N_7050);
nand U7737 (N_7737,N_7182,N_6947);
and U7738 (N_7738,N_6838,N_7154);
and U7739 (N_7739,N_6864,N_6902);
and U7740 (N_7740,N_7000,N_6997);
xnor U7741 (N_7741,N_6626,N_6742);
and U7742 (N_7742,N_6855,N_6672);
and U7743 (N_7743,N_6882,N_6692);
or U7744 (N_7744,N_6826,N_7177);
nand U7745 (N_7745,N_6896,N_6957);
and U7746 (N_7746,N_7037,N_7023);
nand U7747 (N_7747,N_6874,N_6620);
and U7748 (N_7748,N_6868,N_7198);
and U7749 (N_7749,N_6866,N_6821);
and U7750 (N_7750,N_7101,N_7162);
nand U7751 (N_7751,N_6810,N_6729);
nand U7752 (N_7752,N_6729,N_7050);
nor U7753 (N_7753,N_6725,N_6776);
nand U7754 (N_7754,N_7168,N_6868);
nor U7755 (N_7755,N_6675,N_7072);
nand U7756 (N_7756,N_7023,N_7125);
nor U7757 (N_7757,N_6848,N_6704);
and U7758 (N_7758,N_6754,N_6738);
xnor U7759 (N_7759,N_6929,N_6897);
nor U7760 (N_7760,N_6971,N_6712);
or U7761 (N_7761,N_6935,N_6728);
or U7762 (N_7762,N_6837,N_6841);
or U7763 (N_7763,N_7104,N_6646);
or U7764 (N_7764,N_7035,N_6865);
xnor U7765 (N_7765,N_6946,N_6636);
xnor U7766 (N_7766,N_7002,N_7059);
nand U7767 (N_7767,N_6754,N_6939);
nor U7768 (N_7768,N_7079,N_6691);
and U7769 (N_7769,N_7011,N_6929);
nand U7770 (N_7770,N_7057,N_6897);
nor U7771 (N_7771,N_6687,N_6766);
and U7772 (N_7772,N_6687,N_6665);
or U7773 (N_7773,N_6938,N_6664);
xnor U7774 (N_7774,N_6975,N_7004);
or U7775 (N_7775,N_7192,N_6762);
nand U7776 (N_7776,N_6760,N_7186);
and U7777 (N_7777,N_6925,N_6774);
or U7778 (N_7778,N_6876,N_6886);
nand U7779 (N_7779,N_6955,N_7193);
xor U7780 (N_7780,N_6970,N_6877);
xnor U7781 (N_7781,N_6927,N_6988);
and U7782 (N_7782,N_6667,N_6780);
or U7783 (N_7783,N_6913,N_7169);
xnor U7784 (N_7784,N_7140,N_6999);
or U7785 (N_7785,N_7128,N_6844);
or U7786 (N_7786,N_6688,N_6735);
nor U7787 (N_7787,N_6888,N_6617);
nand U7788 (N_7788,N_6765,N_6734);
nand U7789 (N_7789,N_7023,N_6720);
or U7790 (N_7790,N_6990,N_6882);
nand U7791 (N_7791,N_7152,N_6601);
xnor U7792 (N_7792,N_6985,N_6669);
xnor U7793 (N_7793,N_6960,N_6806);
nand U7794 (N_7794,N_6628,N_6723);
xor U7795 (N_7795,N_7020,N_7132);
xor U7796 (N_7796,N_6799,N_7050);
nand U7797 (N_7797,N_6755,N_7042);
nor U7798 (N_7798,N_6943,N_6868);
and U7799 (N_7799,N_6648,N_6876);
and U7800 (N_7800,N_7782,N_7335);
and U7801 (N_7801,N_7688,N_7684);
nor U7802 (N_7802,N_7741,N_7443);
nor U7803 (N_7803,N_7796,N_7632);
nor U7804 (N_7804,N_7547,N_7300);
or U7805 (N_7805,N_7543,N_7601);
or U7806 (N_7806,N_7572,N_7452);
nor U7807 (N_7807,N_7683,N_7240);
or U7808 (N_7808,N_7320,N_7783);
or U7809 (N_7809,N_7234,N_7721);
nand U7810 (N_7810,N_7231,N_7448);
nand U7811 (N_7811,N_7607,N_7315);
xnor U7812 (N_7812,N_7505,N_7723);
nand U7813 (N_7813,N_7730,N_7344);
or U7814 (N_7814,N_7449,N_7359);
nor U7815 (N_7815,N_7690,N_7617);
and U7816 (N_7816,N_7209,N_7576);
and U7817 (N_7817,N_7790,N_7524);
and U7818 (N_7818,N_7337,N_7250);
nand U7819 (N_7819,N_7507,N_7373);
nand U7820 (N_7820,N_7674,N_7385);
nor U7821 (N_7821,N_7597,N_7454);
nor U7822 (N_7822,N_7622,N_7546);
nor U7823 (N_7823,N_7791,N_7598);
nor U7824 (N_7824,N_7716,N_7357);
xor U7825 (N_7825,N_7729,N_7327);
and U7826 (N_7826,N_7522,N_7257);
and U7827 (N_7827,N_7540,N_7680);
nand U7828 (N_7828,N_7478,N_7466);
or U7829 (N_7829,N_7290,N_7686);
nand U7830 (N_7830,N_7301,N_7429);
and U7831 (N_7831,N_7370,N_7244);
nand U7832 (N_7832,N_7289,N_7776);
or U7833 (N_7833,N_7433,N_7494);
nor U7834 (N_7834,N_7313,N_7465);
nand U7835 (N_7835,N_7308,N_7423);
or U7836 (N_7836,N_7795,N_7797);
xnor U7837 (N_7837,N_7718,N_7724);
nand U7838 (N_7838,N_7519,N_7446);
or U7839 (N_7839,N_7275,N_7487);
xnor U7840 (N_7840,N_7331,N_7656);
nor U7841 (N_7841,N_7734,N_7554);
and U7842 (N_7842,N_7752,N_7355);
xor U7843 (N_7843,N_7468,N_7295);
xnor U7844 (N_7844,N_7419,N_7412);
nand U7845 (N_7845,N_7657,N_7658);
nor U7846 (N_7846,N_7411,N_7521);
xor U7847 (N_7847,N_7604,N_7709);
xnor U7848 (N_7848,N_7529,N_7259);
nand U7849 (N_7849,N_7489,N_7365);
nand U7850 (N_7850,N_7341,N_7261);
nand U7851 (N_7851,N_7215,N_7749);
nand U7852 (N_7852,N_7418,N_7799);
nand U7853 (N_7853,N_7390,N_7508);
or U7854 (N_7854,N_7386,N_7611);
xnor U7855 (N_7855,N_7348,N_7303);
or U7856 (N_7856,N_7515,N_7474);
and U7857 (N_7857,N_7410,N_7606);
nand U7858 (N_7858,N_7281,N_7538);
or U7859 (N_7859,N_7777,N_7774);
xor U7860 (N_7860,N_7694,N_7445);
or U7861 (N_7861,N_7273,N_7773);
or U7862 (N_7862,N_7541,N_7556);
or U7863 (N_7863,N_7728,N_7230);
xnor U7864 (N_7864,N_7582,N_7316);
nand U7865 (N_7865,N_7266,N_7485);
or U7866 (N_7866,N_7772,N_7246);
xor U7867 (N_7867,N_7587,N_7623);
or U7868 (N_7868,N_7428,N_7398);
and U7869 (N_7869,N_7283,N_7490);
or U7870 (N_7870,N_7374,N_7340);
nand U7871 (N_7871,N_7416,N_7731);
nand U7872 (N_7872,N_7450,N_7531);
or U7873 (N_7873,N_7545,N_7533);
nand U7874 (N_7874,N_7462,N_7691);
or U7875 (N_7875,N_7479,N_7424);
nand U7876 (N_7876,N_7210,N_7251);
nand U7877 (N_7877,N_7594,N_7548);
nor U7878 (N_7878,N_7375,N_7253);
or U7879 (N_7879,N_7417,N_7558);
nor U7880 (N_7880,N_7422,N_7229);
or U7881 (N_7881,N_7496,N_7669);
xor U7882 (N_7882,N_7233,N_7382);
xnor U7883 (N_7883,N_7368,N_7406);
and U7884 (N_7884,N_7612,N_7653);
or U7885 (N_7885,N_7595,N_7740);
nand U7886 (N_7886,N_7467,N_7338);
or U7887 (N_7887,N_7279,N_7397);
xor U7888 (N_7888,N_7792,N_7704);
nand U7889 (N_7889,N_7277,N_7322);
xor U7890 (N_7890,N_7225,N_7343);
xor U7891 (N_7891,N_7592,N_7330);
nand U7892 (N_7892,N_7769,N_7352);
nand U7893 (N_7893,N_7564,N_7329);
and U7894 (N_7894,N_7747,N_7732);
and U7895 (N_7895,N_7224,N_7756);
xor U7896 (N_7896,N_7642,N_7274);
and U7897 (N_7897,N_7380,N_7270);
and U7898 (N_7898,N_7719,N_7254);
nand U7899 (N_7899,N_7506,N_7414);
or U7900 (N_7900,N_7463,N_7255);
and U7901 (N_7901,N_7248,N_7460);
xor U7902 (N_7902,N_7237,N_7648);
nor U7903 (N_7903,N_7523,N_7408);
nand U7904 (N_7904,N_7761,N_7659);
or U7905 (N_7905,N_7513,N_7206);
nor U7906 (N_7906,N_7318,N_7407);
nand U7907 (N_7907,N_7364,N_7638);
or U7908 (N_7908,N_7498,N_7590);
or U7909 (N_7909,N_7349,N_7635);
nor U7910 (N_7910,N_7326,N_7561);
xnor U7911 (N_7911,N_7625,N_7511);
nor U7912 (N_7912,N_7204,N_7325);
xnor U7913 (N_7913,N_7744,N_7285);
and U7914 (N_7914,N_7353,N_7333);
nor U7915 (N_7915,N_7312,N_7654);
xnor U7916 (N_7916,N_7586,N_7346);
or U7917 (N_7917,N_7559,N_7366);
xor U7918 (N_7918,N_7563,N_7299);
nand U7919 (N_7919,N_7581,N_7557);
or U7920 (N_7920,N_7770,N_7593);
or U7921 (N_7921,N_7778,N_7666);
nand U7922 (N_7922,N_7512,N_7608);
xnor U7923 (N_7923,N_7514,N_7534);
nor U7924 (N_7924,N_7766,N_7748);
nand U7925 (N_7925,N_7535,N_7311);
nor U7926 (N_7926,N_7702,N_7631);
nor U7927 (N_7927,N_7323,N_7453);
nand U7928 (N_7928,N_7425,N_7268);
xor U7929 (N_7929,N_7575,N_7413);
xnor U7930 (N_7930,N_7614,N_7710);
nor U7931 (N_7931,N_7367,N_7305);
nand U7932 (N_7932,N_7616,N_7354);
nor U7933 (N_7933,N_7220,N_7495);
and U7934 (N_7934,N_7228,N_7222);
and U7935 (N_7935,N_7660,N_7288);
nand U7936 (N_7936,N_7457,N_7409);
or U7937 (N_7937,N_7542,N_7434);
and U7938 (N_7938,N_7497,N_7400);
nor U7939 (N_7939,N_7464,N_7726);
or U7940 (N_7940,N_7389,N_7698);
or U7941 (N_7941,N_7663,N_7361);
xnor U7942 (N_7942,N_7664,N_7238);
xnor U7943 (N_7943,N_7665,N_7739);
nor U7944 (N_7944,N_7202,N_7319);
nor U7945 (N_7945,N_7712,N_7271);
and U7946 (N_7946,N_7420,N_7763);
xnor U7947 (N_7947,N_7570,N_7603);
xor U7948 (N_7948,N_7336,N_7342);
and U7949 (N_7949,N_7550,N_7351);
nor U7950 (N_7950,N_7526,N_7219);
nor U7951 (N_7951,N_7636,N_7471);
nor U7952 (N_7952,N_7596,N_7458);
nor U7953 (N_7953,N_7626,N_7713);
or U7954 (N_7954,N_7404,N_7633);
or U7955 (N_7955,N_7286,N_7201);
nor U7956 (N_7956,N_7759,N_7501);
nand U7957 (N_7957,N_7272,N_7527);
xor U7958 (N_7958,N_7641,N_7758);
xnor U7959 (N_7959,N_7269,N_7309);
xnor U7960 (N_7960,N_7383,N_7403);
xnor U7961 (N_7961,N_7306,N_7571);
and U7962 (N_7962,N_7530,N_7589);
xnor U7963 (N_7963,N_7214,N_7245);
or U7964 (N_7964,N_7249,N_7562);
nor U7965 (N_7965,N_7481,N_7753);
or U7966 (N_7966,N_7236,N_7304);
and U7967 (N_7967,N_7788,N_7700);
xor U7968 (N_7968,N_7701,N_7263);
nand U7969 (N_7969,N_7282,N_7668);
nor U7970 (N_7970,N_7447,N_7476);
nor U7971 (N_7971,N_7256,N_7401);
nand U7972 (N_7972,N_7332,N_7339);
or U7973 (N_7973,N_7738,N_7262);
or U7974 (N_7974,N_7678,N_7284);
nand U7975 (N_7975,N_7567,N_7402);
nand U7976 (N_7976,N_7395,N_7786);
or U7977 (N_7977,N_7544,N_7399);
nand U7978 (N_7978,N_7552,N_7579);
nand U7979 (N_7979,N_7280,N_7627);
nor U7980 (N_7980,N_7583,N_7207);
nor U7981 (N_7981,N_7693,N_7297);
and U7982 (N_7982,N_7265,N_7314);
xnor U7983 (N_7983,N_7681,N_7588);
nor U7984 (N_7984,N_7293,N_7500);
or U7985 (N_7985,N_7672,N_7662);
and U7986 (N_7986,N_7682,N_7358);
xor U7987 (N_7987,N_7405,N_7208);
or U7988 (N_7988,N_7427,N_7624);
nand U7989 (N_7989,N_7287,N_7580);
or U7990 (N_7990,N_7430,N_7647);
nor U7991 (N_7991,N_7363,N_7298);
nor U7992 (N_7992,N_7620,N_7421);
nor U7993 (N_7993,N_7517,N_7321);
and U7994 (N_7994,N_7651,N_7599);
or U7995 (N_7995,N_7733,N_7509);
and U7996 (N_7996,N_7762,N_7745);
and U7997 (N_7997,N_7569,N_7644);
and U7998 (N_7998,N_7372,N_7650);
nand U7999 (N_7999,N_7394,N_7211);
nor U8000 (N_8000,N_7798,N_7675);
or U8001 (N_8001,N_7605,N_7396);
and U8002 (N_8002,N_7520,N_7439);
or U8003 (N_8003,N_7577,N_7317);
and U8004 (N_8004,N_7735,N_7661);
xor U8005 (N_8005,N_7767,N_7568);
and U8006 (N_8006,N_7736,N_7781);
xor U8007 (N_8007,N_7573,N_7760);
nand U8008 (N_8008,N_7722,N_7223);
and U8009 (N_8009,N_7765,N_7221);
nand U8010 (N_8010,N_7676,N_7768);
xnor U8011 (N_8011,N_7241,N_7750);
xor U8012 (N_8012,N_7388,N_7461);
nor U8013 (N_8013,N_7387,N_7585);
or U8014 (N_8014,N_7706,N_7737);
nor U8015 (N_8015,N_7560,N_7673);
and U8016 (N_8016,N_7708,N_7278);
and U8017 (N_8017,N_7431,N_7324);
nor U8018 (N_8018,N_7294,N_7473);
xnor U8019 (N_8019,N_7714,N_7291);
nor U8020 (N_8020,N_7685,N_7391);
nor U8021 (N_8021,N_7536,N_7493);
xor U8022 (N_8022,N_7757,N_7785);
nor U8023 (N_8023,N_7630,N_7574);
or U8024 (N_8024,N_7213,N_7393);
nand U8025 (N_8025,N_7591,N_7426);
nor U8026 (N_8026,N_7252,N_7720);
or U8027 (N_8027,N_7565,N_7356);
and U8028 (N_8028,N_7646,N_7742);
and U8029 (N_8029,N_7216,N_7384);
and U8030 (N_8030,N_7537,N_7743);
and U8031 (N_8031,N_7687,N_7755);
nor U8032 (N_8032,N_7670,N_7692);
or U8033 (N_8033,N_7584,N_7551);
and U8034 (N_8034,N_7444,N_7243);
or U8035 (N_8035,N_7634,N_7618);
or U8036 (N_8036,N_7609,N_7499);
xnor U8037 (N_8037,N_7532,N_7566);
nand U8038 (N_8038,N_7455,N_7267);
xnor U8039 (N_8039,N_7707,N_7480);
xor U8040 (N_8040,N_7486,N_7754);
or U8041 (N_8041,N_7475,N_7711);
nor U8042 (N_8042,N_7516,N_7307);
nor U8043 (N_8043,N_7264,N_7725);
nor U8044 (N_8044,N_7751,N_7226);
xnor U8045 (N_8045,N_7203,N_7677);
or U8046 (N_8046,N_7779,N_7470);
and U8047 (N_8047,N_7371,N_7483);
nand U8048 (N_8048,N_7696,N_7775);
and U8049 (N_8049,N_7381,N_7328);
and U8050 (N_8050,N_7610,N_7679);
nor U8051 (N_8051,N_7459,N_7469);
xor U8052 (N_8052,N_7440,N_7518);
nand U8053 (N_8053,N_7671,N_7784);
or U8054 (N_8054,N_7771,N_7697);
nand U8055 (N_8055,N_7345,N_7602);
nand U8056 (N_8056,N_7510,N_7296);
nand U8057 (N_8057,N_7482,N_7491);
nor U8058 (N_8058,N_7437,N_7689);
xnor U8059 (N_8059,N_7637,N_7362);
nor U8060 (N_8060,N_7212,N_7360);
xnor U8061 (N_8061,N_7699,N_7379);
or U8062 (N_8062,N_7787,N_7695);
nor U8063 (N_8063,N_7715,N_7432);
or U8064 (N_8064,N_7705,N_7621);
nand U8065 (N_8065,N_7350,N_7369);
and U8066 (N_8066,N_7539,N_7528);
nand U8067 (N_8067,N_7347,N_7438);
and U8068 (N_8068,N_7488,N_7292);
nor U8069 (N_8069,N_7502,N_7628);
and U8070 (N_8070,N_7525,N_7477);
xnor U8071 (N_8071,N_7615,N_7789);
and U8072 (N_8072,N_7232,N_7764);
or U8073 (N_8073,N_7793,N_7639);
xnor U8074 (N_8074,N_7441,N_7794);
and U8075 (N_8075,N_7578,N_7504);
xnor U8076 (N_8076,N_7456,N_7451);
and U8077 (N_8077,N_7376,N_7217);
or U8078 (N_8078,N_7242,N_7727);
xor U8079 (N_8079,N_7235,N_7436);
and U8080 (N_8080,N_7649,N_7442);
nand U8081 (N_8081,N_7205,N_7549);
xor U8082 (N_8082,N_7613,N_7310);
and U8083 (N_8083,N_7746,N_7484);
xor U8084 (N_8084,N_7655,N_7247);
xor U8085 (N_8085,N_7645,N_7703);
nor U8086 (N_8086,N_7555,N_7652);
or U8087 (N_8087,N_7200,N_7492);
xnor U8088 (N_8088,N_7640,N_7227);
nor U8089 (N_8089,N_7415,N_7334);
xor U8090 (N_8090,N_7378,N_7553);
xor U8091 (N_8091,N_7260,N_7667);
nand U8092 (N_8092,N_7218,N_7629);
or U8093 (N_8093,N_7377,N_7600);
nand U8094 (N_8094,N_7239,N_7503);
nand U8095 (N_8095,N_7435,N_7717);
or U8096 (N_8096,N_7258,N_7643);
nor U8097 (N_8097,N_7392,N_7619);
and U8098 (N_8098,N_7780,N_7302);
or U8099 (N_8099,N_7276,N_7472);
xnor U8100 (N_8100,N_7490,N_7499);
nand U8101 (N_8101,N_7588,N_7750);
nor U8102 (N_8102,N_7515,N_7292);
and U8103 (N_8103,N_7539,N_7761);
and U8104 (N_8104,N_7366,N_7444);
or U8105 (N_8105,N_7344,N_7238);
nand U8106 (N_8106,N_7769,N_7496);
xnor U8107 (N_8107,N_7366,N_7485);
nand U8108 (N_8108,N_7491,N_7289);
nand U8109 (N_8109,N_7573,N_7747);
or U8110 (N_8110,N_7539,N_7317);
xor U8111 (N_8111,N_7324,N_7277);
xor U8112 (N_8112,N_7568,N_7279);
nor U8113 (N_8113,N_7474,N_7333);
nor U8114 (N_8114,N_7344,N_7777);
or U8115 (N_8115,N_7569,N_7595);
nor U8116 (N_8116,N_7562,N_7544);
nor U8117 (N_8117,N_7279,N_7444);
nor U8118 (N_8118,N_7792,N_7730);
or U8119 (N_8119,N_7575,N_7338);
xor U8120 (N_8120,N_7334,N_7530);
nor U8121 (N_8121,N_7688,N_7308);
and U8122 (N_8122,N_7698,N_7678);
or U8123 (N_8123,N_7609,N_7745);
nand U8124 (N_8124,N_7308,N_7700);
xnor U8125 (N_8125,N_7271,N_7644);
or U8126 (N_8126,N_7287,N_7206);
nand U8127 (N_8127,N_7313,N_7523);
or U8128 (N_8128,N_7453,N_7359);
or U8129 (N_8129,N_7532,N_7689);
and U8130 (N_8130,N_7588,N_7615);
or U8131 (N_8131,N_7634,N_7310);
nand U8132 (N_8132,N_7533,N_7675);
nand U8133 (N_8133,N_7241,N_7479);
nand U8134 (N_8134,N_7391,N_7471);
or U8135 (N_8135,N_7507,N_7311);
nand U8136 (N_8136,N_7469,N_7518);
or U8137 (N_8137,N_7401,N_7267);
xnor U8138 (N_8138,N_7393,N_7369);
and U8139 (N_8139,N_7250,N_7762);
nor U8140 (N_8140,N_7752,N_7313);
and U8141 (N_8141,N_7628,N_7500);
nand U8142 (N_8142,N_7437,N_7682);
or U8143 (N_8143,N_7593,N_7647);
and U8144 (N_8144,N_7490,N_7445);
or U8145 (N_8145,N_7514,N_7576);
or U8146 (N_8146,N_7459,N_7683);
nand U8147 (N_8147,N_7781,N_7734);
nand U8148 (N_8148,N_7741,N_7785);
xor U8149 (N_8149,N_7217,N_7462);
and U8150 (N_8150,N_7236,N_7614);
and U8151 (N_8151,N_7459,N_7707);
or U8152 (N_8152,N_7761,N_7358);
or U8153 (N_8153,N_7693,N_7405);
or U8154 (N_8154,N_7269,N_7239);
xor U8155 (N_8155,N_7641,N_7684);
nand U8156 (N_8156,N_7344,N_7733);
nor U8157 (N_8157,N_7531,N_7594);
nand U8158 (N_8158,N_7393,N_7455);
or U8159 (N_8159,N_7717,N_7654);
nor U8160 (N_8160,N_7782,N_7308);
and U8161 (N_8161,N_7374,N_7317);
nand U8162 (N_8162,N_7279,N_7609);
xnor U8163 (N_8163,N_7247,N_7639);
nor U8164 (N_8164,N_7498,N_7274);
nand U8165 (N_8165,N_7515,N_7424);
and U8166 (N_8166,N_7716,N_7309);
nand U8167 (N_8167,N_7489,N_7582);
xor U8168 (N_8168,N_7755,N_7416);
and U8169 (N_8169,N_7670,N_7571);
nor U8170 (N_8170,N_7499,N_7219);
and U8171 (N_8171,N_7635,N_7650);
nor U8172 (N_8172,N_7656,N_7618);
and U8173 (N_8173,N_7553,N_7694);
nor U8174 (N_8174,N_7406,N_7674);
or U8175 (N_8175,N_7764,N_7257);
nand U8176 (N_8176,N_7345,N_7228);
and U8177 (N_8177,N_7517,N_7490);
and U8178 (N_8178,N_7606,N_7387);
nor U8179 (N_8179,N_7590,N_7645);
nand U8180 (N_8180,N_7300,N_7228);
or U8181 (N_8181,N_7649,N_7566);
or U8182 (N_8182,N_7317,N_7566);
or U8183 (N_8183,N_7716,N_7744);
nand U8184 (N_8184,N_7279,N_7483);
and U8185 (N_8185,N_7742,N_7595);
and U8186 (N_8186,N_7585,N_7568);
or U8187 (N_8187,N_7661,N_7704);
nand U8188 (N_8188,N_7612,N_7415);
and U8189 (N_8189,N_7488,N_7654);
or U8190 (N_8190,N_7546,N_7611);
nor U8191 (N_8191,N_7377,N_7508);
and U8192 (N_8192,N_7219,N_7677);
or U8193 (N_8193,N_7570,N_7656);
xnor U8194 (N_8194,N_7703,N_7291);
xor U8195 (N_8195,N_7447,N_7599);
nor U8196 (N_8196,N_7246,N_7650);
xnor U8197 (N_8197,N_7667,N_7520);
nand U8198 (N_8198,N_7261,N_7626);
nor U8199 (N_8199,N_7475,N_7346);
or U8200 (N_8200,N_7326,N_7316);
xor U8201 (N_8201,N_7326,N_7422);
nand U8202 (N_8202,N_7240,N_7667);
and U8203 (N_8203,N_7530,N_7577);
xnor U8204 (N_8204,N_7665,N_7572);
or U8205 (N_8205,N_7749,N_7707);
or U8206 (N_8206,N_7576,N_7604);
or U8207 (N_8207,N_7388,N_7483);
xor U8208 (N_8208,N_7618,N_7725);
and U8209 (N_8209,N_7784,N_7485);
or U8210 (N_8210,N_7720,N_7787);
xor U8211 (N_8211,N_7779,N_7657);
or U8212 (N_8212,N_7444,N_7340);
nor U8213 (N_8213,N_7224,N_7795);
xnor U8214 (N_8214,N_7434,N_7697);
and U8215 (N_8215,N_7229,N_7260);
xor U8216 (N_8216,N_7727,N_7411);
nor U8217 (N_8217,N_7414,N_7781);
and U8218 (N_8218,N_7672,N_7569);
nand U8219 (N_8219,N_7738,N_7614);
nor U8220 (N_8220,N_7569,N_7682);
and U8221 (N_8221,N_7517,N_7678);
nor U8222 (N_8222,N_7253,N_7369);
xor U8223 (N_8223,N_7293,N_7607);
nor U8224 (N_8224,N_7527,N_7287);
nand U8225 (N_8225,N_7719,N_7708);
xnor U8226 (N_8226,N_7412,N_7561);
and U8227 (N_8227,N_7481,N_7639);
or U8228 (N_8228,N_7629,N_7306);
nand U8229 (N_8229,N_7635,N_7771);
nand U8230 (N_8230,N_7706,N_7566);
xor U8231 (N_8231,N_7419,N_7292);
and U8232 (N_8232,N_7216,N_7354);
or U8233 (N_8233,N_7751,N_7502);
nand U8234 (N_8234,N_7227,N_7410);
or U8235 (N_8235,N_7470,N_7491);
nand U8236 (N_8236,N_7307,N_7601);
or U8237 (N_8237,N_7751,N_7478);
nand U8238 (N_8238,N_7685,N_7735);
xnor U8239 (N_8239,N_7541,N_7544);
and U8240 (N_8240,N_7210,N_7516);
nor U8241 (N_8241,N_7319,N_7415);
xor U8242 (N_8242,N_7640,N_7447);
and U8243 (N_8243,N_7239,N_7433);
xor U8244 (N_8244,N_7563,N_7425);
or U8245 (N_8245,N_7347,N_7569);
and U8246 (N_8246,N_7745,N_7260);
nand U8247 (N_8247,N_7205,N_7500);
nor U8248 (N_8248,N_7390,N_7425);
or U8249 (N_8249,N_7598,N_7582);
nand U8250 (N_8250,N_7714,N_7752);
xnor U8251 (N_8251,N_7586,N_7534);
or U8252 (N_8252,N_7290,N_7731);
nand U8253 (N_8253,N_7718,N_7614);
xnor U8254 (N_8254,N_7272,N_7784);
or U8255 (N_8255,N_7689,N_7413);
xor U8256 (N_8256,N_7533,N_7654);
nand U8257 (N_8257,N_7608,N_7497);
nor U8258 (N_8258,N_7467,N_7431);
xnor U8259 (N_8259,N_7325,N_7377);
xor U8260 (N_8260,N_7639,N_7383);
or U8261 (N_8261,N_7401,N_7502);
nor U8262 (N_8262,N_7263,N_7406);
nor U8263 (N_8263,N_7781,N_7660);
and U8264 (N_8264,N_7467,N_7208);
or U8265 (N_8265,N_7466,N_7775);
xnor U8266 (N_8266,N_7770,N_7612);
nor U8267 (N_8267,N_7549,N_7287);
nor U8268 (N_8268,N_7593,N_7600);
nor U8269 (N_8269,N_7739,N_7275);
nand U8270 (N_8270,N_7252,N_7573);
nand U8271 (N_8271,N_7662,N_7339);
or U8272 (N_8272,N_7792,N_7437);
and U8273 (N_8273,N_7512,N_7690);
or U8274 (N_8274,N_7414,N_7769);
xor U8275 (N_8275,N_7426,N_7267);
nor U8276 (N_8276,N_7667,N_7301);
and U8277 (N_8277,N_7583,N_7251);
nor U8278 (N_8278,N_7731,N_7792);
and U8279 (N_8279,N_7456,N_7655);
nor U8280 (N_8280,N_7615,N_7336);
and U8281 (N_8281,N_7754,N_7759);
nor U8282 (N_8282,N_7459,N_7672);
nor U8283 (N_8283,N_7749,N_7254);
nand U8284 (N_8284,N_7390,N_7474);
nand U8285 (N_8285,N_7387,N_7351);
xnor U8286 (N_8286,N_7500,N_7606);
xnor U8287 (N_8287,N_7775,N_7268);
nor U8288 (N_8288,N_7572,N_7549);
nand U8289 (N_8289,N_7248,N_7264);
xnor U8290 (N_8290,N_7534,N_7652);
nand U8291 (N_8291,N_7786,N_7694);
or U8292 (N_8292,N_7640,N_7726);
nor U8293 (N_8293,N_7550,N_7545);
or U8294 (N_8294,N_7711,N_7626);
nor U8295 (N_8295,N_7753,N_7605);
nand U8296 (N_8296,N_7227,N_7583);
nor U8297 (N_8297,N_7577,N_7588);
and U8298 (N_8298,N_7788,N_7704);
and U8299 (N_8299,N_7515,N_7730);
nand U8300 (N_8300,N_7747,N_7324);
or U8301 (N_8301,N_7547,N_7200);
xor U8302 (N_8302,N_7348,N_7781);
or U8303 (N_8303,N_7486,N_7593);
and U8304 (N_8304,N_7509,N_7701);
and U8305 (N_8305,N_7207,N_7681);
nand U8306 (N_8306,N_7783,N_7765);
xor U8307 (N_8307,N_7344,N_7401);
or U8308 (N_8308,N_7237,N_7460);
nor U8309 (N_8309,N_7752,N_7574);
xor U8310 (N_8310,N_7615,N_7651);
xnor U8311 (N_8311,N_7631,N_7380);
nand U8312 (N_8312,N_7654,N_7283);
nand U8313 (N_8313,N_7258,N_7440);
nand U8314 (N_8314,N_7502,N_7763);
and U8315 (N_8315,N_7236,N_7605);
and U8316 (N_8316,N_7442,N_7325);
and U8317 (N_8317,N_7368,N_7447);
nand U8318 (N_8318,N_7204,N_7558);
nor U8319 (N_8319,N_7280,N_7459);
nor U8320 (N_8320,N_7315,N_7277);
and U8321 (N_8321,N_7508,N_7701);
and U8322 (N_8322,N_7512,N_7437);
xor U8323 (N_8323,N_7443,N_7614);
and U8324 (N_8324,N_7343,N_7743);
nand U8325 (N_8325,N_7296,N_7578);
or U8326 (N_8326,N_7261,N_7455);
and U8327 (N_8327,N_7563,N_7770);
or U8328 (N_8328,N_7300,N_7330);
xor U8329 (N_8329,N_7210,N_7460);
nor U8330 (N_8330,N_7290,N_7568);
and U8331 (N_8331,N_7707,N_7383);
nand U8332 (N_8332,N_7437,N_7370);
or U8333 (N_8333,N_7518,N_7496);
nor U8334 (N_8334,N_7584,N_7718);
nand U8335 (N_8335,N_7200,N_7607);
and U8336 (N_8336,N_7689,N_7702);
xnor U8337 (N_8337,N_7277,N_7406);
xor U8338 (N_8338,N_7666,N_7598);
nor U8339 (N_8339,N_7760,N_7484);
and U8340 (N_8340,N_7522,N_7383);
nor U8341 (N_8341,N_7472,N_7700);
or U8342 (N_8342,N_7312,N_7672);
nand U8343 (N_8343,N_7574,N_7511);
or U8344 (N_8344,N_7704,N_7470);
or U8345 (N_8345,N_7286,N_7271);
or U8346 (N_8346,N_7387,N_7509);
nand U8347 (N_8347,N_7793,N_7707);
xnor U8348 (N_8348,N_7617,N_7738);
nor U8349 (N_8349,N_7265,N_7690);
nor U8350 (N_8350,N_7577,N_7517);
or U8351 (N_8351,N_7541,N_7405);
xnor U8352 (N_8352,N_7463,N_7263);
and U8353 (N_8353,N_7559,N_7208);
nand U8354 (N_8354,N_7506,N_7542);
nor U8355 (N_8355,N_7557,N_7207);
and U8356 (N_8356,N_7717,N_7302);
nor U8357 (N_8357,N_7276,N_7575);
nor U8358 (N_8358,N_7699,N_7580);
xnor U8359 (N_8359,N_7496,N_7214);
xnor U8360 (N_8360,N_7789,N_7555);
nor U8361 (N_8361,N_7395,N_7663);
nor U8362 (N_8362,N_7301,N_7729);
xor U8363 (N_8363,N_7484,N_7260);
nor U8364 (N_8364,N_7639,N_7384);
or U8365 (N_8365,N_7202,N_7246);
or U8366 (N_8366,N_7631,N_7755);
nor U8367 (N_8367,N_7402,N_7356);
nand U8368 (N_8368,N_7545,N_7558);
or U8369 (N_8369,N_7632,N_7526);
nand U8370 (N_8370,N_7217,N_7387);
or U8371 (N_8371,N_7611,N_7435);
or U8372 (N_8372,N_7413,N_7374);
nor U8373 (N_8373,N_7385,N_7735);
and U8374 (N_8374,N_7700,N_7200);
xnor U8375 (N_8375,N_7299,N_7465);
or U8376 (N_8376,N_7577,N_7644);
or U8377 (N_8377,N_7355,N_7766);
nand U8378 (N_8378,N_7323,N_7762);
and U8379 (N_8379,N_7731,N_7288);
xnor U8380 (N_8380,N_7250,N_7572);
nand U8381 (N_8381,N_7732,N_7408);
and U8382 (N_8382,N_7331,N_7796);
and U8383 (N_8383,N_7684,N_7313);
nor U8384 (N_8384,N_7291,N_7305);
nor U8385 (N_8385,N_7530,N_7249);
nand U8386 (N_8386,N_7664,N_7574);
and U8387 (N_8387,N_7506,N_7710);
or U8388 (N_8388,N_7377,N_7661);
nor U8389 (N_8389,N_7318,N_7530);
nand U8390 (N_8390,N_7639,N_7553);
nand U8391 (N_8391,N_7794,N_7235);
nand U8392 (N_8392,N_7453,N_7289);
nand U8393 (N_8393,N_7625,N_7562);
xor U8394 (N_8394,N_7263,N_7547);
xnor U8395 (N_8395,N_7665,N_7292);
nand U8396 (N_8396,N_7528,N_7231);
nor U8397 (N_8397,N_7613,N_7700);
or U8398 (N_8398,N_7223,N_7218);
xor U8399 (N_8399,N_7474,N_7585);
and U8400 (N_8400,N_8028,N_8049);
and U8401 (N_8401,N_8352,N_7905);
or U8402 (N_8402,N_8086,N_7856);
nand U8403 (N_8403,N_7802,N_8017);
nor U8404 (N_8404,N_7849,N_8335);
nor U8405 (N_8405,N_8253,N_8209);
or U8406 (N_8406,N_7911,N_8260);
nor U8407 (N_8407,N_8298,N_8362);
xnor U8408 (N_8408,N_8398,N_8125);
or U8409 (N_8409,N_8081,N_8007);
nor U8410 (N_8410,N_8337,N_8107);
or U8411 (N_8411,N_7800,N_7917);
xnor U8412 (N_8412,N_8350,N_7862);
and U8413 (N_8413,N_8376,N_8185);
xor U8414 (N_8414,N_8382,N_8392);
xnor U8415 (N_8415,N_7968,N_7861);
xnor U8416 (N_8416,N_7847,N_8122);
xnor U8417 (N_8417,N_8277,N_7959);
xnor U8418 (N_8418,N_8315,N_8189);
or U8419 (N_8419,N_8041,N_7907);
or U8420 (N_8420,N_7990,N_8039);
nand U8421 (N_8421,N_8083,N_8345);
nor U8422 (N_8422,N_8073,N_8267);
and U8423 (N_8423,N_8326,N_7895);
xnor U8424 (N_8424,N_8372,N_8265);
and U8425 (N_8425,N_7936,N_8332);
or U8426 (N_8426,N_8232,N_8109);
and U8427 (N_8427,N_8201,N_8274);
and U8428 (N_8428,N_7947,N_7900);
nor U8429 (N_8429,N_8011,N_8047);
xor U8430 (N_8430,N_8286,N_8261);
nand U8431 (N_8431,N_8129,N_8155);
xnor U8432 (N_8432,N_8099,N_8355);
or U8433 (N_8433,N_7814,N_8138);
and U8434 (N_8434,N_8124,N_8116);
xor U8435 (N_8435,N_8238,N_8323);
and U8436 (N_8436,N_7840,N_7854);
and U8437 (N_8437,N_8066,N_7932);
xor U8438 (N_8438,N_7954,N_7839);
xnor U8439 (N_8439,N_7801,N_8187);
and U8440 (N_8440,N_8271,N_7992);
xor U8441 (N_8441,N_8018,N_8316);
or U8442 (N_8442,N_8077,N_8084);
nor U8443 (N_8443,N_8289,N_8374);
nand U8444 (N_8444,N_7989,N_8210);
nor U8445 (N_8445,N_8024,N_8164);
nand U8446 (N_8446,N_7898,N_8059);
or U8447 (N_8447,N_8222,N_8309);
nor U8448 (N_8448,N_7916,N_8218);
xnor U8449 (N_8449,N_7904,N_7995);
or U8450 (N_8450,N_8297,N_7808);
xnor U8451 (N_8451,N_8281,N_7979);
nor U8452 (N_8452,N_8159,N_8091);
nor U8453 (N_8453,N_7891,N_8108);
nor U8454 (N_8454,N_8212,N_8148);
nand U8455 (N_8455,N_8399,N_8031);
nor U8456 (N_8456,N_7957,N_8019);
and U8457 (N_8457,N_7881,N_7953);
nor U8458 (N_8458,N_7883,N_8249);
or U8459 (N_8459,N_7841,N_8293);
xnor U8460 (N_8460,N_8360,N_8319);
xor U8461 (N_8461,N_7944,N_7882);
or U8462 (N_8462,N_7805,N_8068);
or U8463 (N_8463,N_8368,N_8135);
or U8464 (N_8464,N_8283,N_8342);
xnor U8465 (N_8465,N_8063,N_7829);
nand U8466 (N_8466,N_8176,N_7817);
or U8467 (N_8467,N_8141,N_8112);
nor U8468 (N_8468,N_8291,N_8026);
nand U8469 (N_8469,N_7828,N_8065);
nand U8470 (N_8470,N_8178,N_7923);
and U8471 (N_8471,N_8013,N_8095);
or U8472 (N_8472,N_7945,N_8167);
nand U8473 (N_8473,N_7937,N_7943);
nand U8474 (N_8474,N_8002,N_8223);
nand U8475 (N_8475,N_8036,N_8321);
nor U8476 (N_8476,N_8113,N_7848);
nor U8477 (N_8477,N_8053,N_8211);
nand U8478 (N_8478,N_7999,N_8353);
xnor U8479 (N_8479,N_7921,N_8179);
nor U8480 (N_8480,N_8142,N_7868);
nand U8481 (N_8481,N_7876,N_8246);
xor U8482 (N_8482,N_7869,N_8397);
nand U8483 (N_8483,N_7842,N_8133);
or U8484 (N_8484,N_8177,N_8328);
xnor U8485 (N_8485,N_7967,N_8240);
or U8486 (N_8486,N_8393,N_8106);
or U8487 (N_8487,N_7858,N_7844);
nor U8488 (N_8488,N_7815,N_8366);
nand U8489 (N_8489,N_8154,N_7867);
nand U8490 (N_8490,N_8225,N_8126);
nand U8491 (N_8491,N_8237,N_8361);
and U8492 (N_8492,N_7822,N_8330);
nor U8493 (N_8493,N_8388,N_8371);
nand U8494 (N_8494,N_7894,N_8186);
and U8495 (N_8495,N_8358,N_7860);
or U8496 (N_8496,N_8322,N_8224);
nand U8497 (N_8497,N_8386,N_7933);
or U8498 (N_8498,N_8035,N_8389);
or U8499 (N_8499,N_8151,N_8247);
or U8500 (N_8500,N_8137,N_8061);
xor U8501 (N_8501,N_8001,N_8020);
xnor U8502 (N_8502,N_8296,N_8005);
xnor U8503 (N_8503,N_8391,N_8021);
nand U8504 (N_8504,N_8268,N_7925);
or U8505 (N_8505,N_8115,N_7927);
nor U8506 (N_8506,N_8182,N_7913);
nor U8507 (N_8507,N_8236,N_8085);
nand U8508 (N_8508,N_7922,N_7972);
nand U8509 (N_8509,N_8288,N_8255);
xor U8510 (N_8510,N_8040,N_8314);
or U8511 (N_8511,N_8134,N_8384);
or U8512 (N_8512,N_7806,N_7807);
or U8513 (N_8513,N_8147,N_8029);
and U8514 (N_8514,N_8207,N_8287);
or U8515 (N_8515,N_7816,N_8079);
nor U8516 (N_8516,N_8320,N_8146);
xnor U8517 (N_8517,N_8044,N_7978);
xor U8518 (N_8518,N_8336,N_8143);
nand U8519 (N_8519,N_8217,N_8279);
and U8520 (N_8520,N_8284,N_7950);
or U8521 (N_8521,N_8269,N_8311);
or U8522 (N_8522,N_8308,N_8022);
xor U8523 (N_8523,N_8048,N_7819);
and U8524 (N_8524,N_8248,N_7884);
nor U8525 (N_8525,N_8299,N_7892);
xor U8526 (N_8526,N_7930,N_8145);
nor U8527 (N_8527,N_7998,N_8227);
or U8528 (N_8528,N_8183,N_7902);
or U8529 (N_8529,N_8060,N_8363);
and U8530 (N_8530,N_7935,N_8136);
or U8531 (N_8531,N_7912,N_8057);
and U8532 (N_8532,N_8329,N_8160);
nor U8533 (N_8533,N_8027,N_8094);
xnor U8534 (N_8534,N_7973,N_8233);
or U8535 (N_8535,N_8144,N_8303);
nor U8536 (N_8536,N_8307,N_8132);
xor U8537 (N_8537,N_8226,N_8276);
xor U8538 (N_8538,N_8102,N_8254);
or U8539 (N_8539,N_7827,N_8295);
and U8540 (N_8540,N_8317,N_7880);
and U8541 (N_8541,N_7981,N_8009);
xnor U8542 (N_8542,N_8300,N_8341);
nand U8543 (N_8543,N_8064,N_8069);
nand U8544 (N_8544,N_8357,N_8356);
xor U8545 (N_8545,N_8275,N_8175);
xnor U8546 (N_8546,N_7803,N_8032);
and U8547 (N_8547,N_7871,N_8266);
and U8548 (N_8548,N_8256,N_8121);
nand U8549 (N_8549,N_8184,N_8383);
and U8550 (N_8550,N_8093,N_8340);
nand U8551 (N_8551,N_8367,N_7924);
and U8552 (N_8552,N_7926,N_7908);
and U8553 (N_8553,N_8070,N_7890);
nand U8554 (N_8554,N_7826,N_7929);
xnor U8555 (N_8555,N_8200,N_7952);
and U8556 (N_8556,N_7928,N_8195);
nor U8557 (N_8557,N_7966,N_8369);
xnor U8558 (N_8558,N_8394,N_8103);
and U8559 (N_8559,N_8072,N_8023);
xor U8560 (N_8560,N_8202,N_8174);
nand U8561 (N_8561,N_8098,N_8313);
xor U8562 (N_8562,N_8150,N_7846);
nand U8563 (N_8563,N_8364,N_7938);
nand U8564 (N_8564,N_7879,N_8385);
nor U8565 (N_8565,N_8338,N_8205);
xor U8566 (N_8566,N_8170,N_8278);
nand U8567 (N_8567,N_8131,N_8243);
nand U8568 (N_8568,N_8231,N_8310);
or U8569 (N_8569,N_8280,N_8348);
nand U8570 (N_8570,N_8140,N_8118);
or U8571 (N_8571,N_8343,N_8123);
and U8572 (N_8572,N_7980,N_8215);
nor U8573 (N_8573,N_8191,N_7853);
and U8574 (N_8574,N_7857,N_8046);
or U8575 (N_8575,N_8339,N_8169);
xnor U8576 (N_8576,N_8192,N_7996);
xnor U8577 (N_8577,N_8324,N_7956);
or U8578 (N_8578,N_7920,N_7971);
or U8579 (N_8579,N_7811,N_8318);
and U8580 (N_8580,N_7825,N_7866);
or U8581 (N_8581,N_8062,N_7875);
and U8582 (N_8582,N_7974,N_7948);
nand U8583 (N_8583,N_7977,N_7885);
nor U8584 (N_8584,N_7993,N_7969);
xor U8585 (N_8585,N_7909,N_7813);
xnor U8586 (N_8586,N_8188,N_8025);
nor U8587 (N_8587,N_7940,N_8156);
xnor U8588 (N_8588,N_7960,N_8263);
xnor U8589 (N_8589,N_8334,N_8333);
nand U8590 (N_8590,N_7804,N_7835);
nand U8591 (N_8591,N_8104,N_8043);
and U8592 (N_8592,N_8216,N_7919);
and U8593 (N_8593,N_8219,N_7834);
xor U8594 (N_8594,N_8220,N_8290);
nand U8595 (N_8595,N_7991,N_7837);
nand U8596 (N_8596,N_8050,N_7851);
nand U8597 (N_8597,N_8301,N_7889);
nand U8598 (N_8598,N_8306,N_7832);
xnor U8599 (N_8599,N_8387,N_8370);
nor U8600 (N_8600,N_8239,N_8245);
and U8601 (N_8601,N_7863,N_7855);
nand U8602 (N_8602,N_7962,N_8197);
nand U8603 (N_8603,N_7961,N_7838);
or U8604 (N_8604,N_8285,N_8228);
nor U8605 (N_8605,N_8259,N_8365);
and U8606 (N_8606,N_7965,N_8230);
xor U8607 (N_8607,N_8080,N_7914);
and U8608 (N_8608,N_7931,N_8344);
nor U8609 (N_8609,N_7850,N_7918);
xnor U8610 (N_8610,N_7988,N_8194);
nand U8611 (N_8611,N_7903,N_7946);
and U8612 (N_8612,N_7963,N_8252);
nor U8613 (N_8613,N_8139,N_7864);
nand U8614 (N_8614,N_8128,N_8257);
or U8615 (N_8615,N_7983,N_8075);
nor U8616 (N_8616,N_8105,N_8078);
or U8617 (N_8617,N_8006,N_7821);
xnor U8618 (N_8618,N_8234,N_8327);
nor U8619 (N_8619,N_7865,N_8012);
nand U8620 (N_8620,N_8058,N_8166);
xor U8621 (N_8621,N_8258,N_8294);
and U8622 (N_8622,N_7810,N_8395);
nor U8623 (N_8623,N_8067,N_8042);
nor U8624 (N_8624,N_8096,N_8008);
or U8625 (N_8625,N_7859,N_8302);
and U8626 (N_8626,N_8242,N_8162);
xnor U8627 (N_8627,N_8264,N_8052);
nand U8628 (N_8628,N_8037,N_8172);
nand U8629 (N_8629,N_8054,N_7888);
xor U8630 (N_8630,N_8130,N_7887);
nor U8631 (N_8631,N_8325,N_8203);
nor U8632 (N_8632,N_8071,N_8359);
xnor U8633 (N_8633,N_7823,N_8181);
nand U8634 (N_8634,N_8347,N_8171);
xor U8635 (N_8635,N_8196,N_8190);
and U8636 (N_8636,N_8045,N_8272);
xor U8637 (N_8637,N_8375,N_7976);
or U8638 (N_8638,N_8076,N_8173);
and U8639 (N_8639,N_8331,N_8250);
xnor U8640 (N_8640,N_8030,N_7886);
and U8641 (N_8641,N_8282,N_7870);
and U8642 (N_8642,N_8111,N_8101);
and U8643 (N_8643,N_8152,N_8114);
nand U8644 (N_8644,N_7955,N_7893);
nor U8645 (N_8645,N_7897,N_7899);
xor U8646 (N_8646,N_7836,N_8204);
or U8647 (N_8647,N_8090,N_7941);
xnor U8648 (N_8648,N_8119,N_7997);
and U8649 (N_8649,N_7951,N_8056);
nor U8650 (N_8650,N_7964,N_8016);
or U8651 (N_8651,N_8379,N_8206);
xor U8652 (N_8652,N_7824,N_8380);
or U8653 (N_8653,N_8377,N_8244);
xnor U8654 (N_8654,N_7949,N_7843);
nor U8655 (N_8655,N_8055,N_7831);
xnor U8656 (N_8656,N_7833,N_8213);
xnor U8657 (N_8657,N_8346,N_7873);
nand U8658 (N_8658,N_8168,N_7910);
or U8659 (N_8659,N_8161,N_8003);
xor U8660 (N_8660,N_8014,N_8292);
and U8661 (N_8661,N_7896,N_8088);
nand U8662 (N_8662,N_8082,N_8312);
nor U8663 (N_8663,N_8251,N_8373);
or U8664 (N_8664,N_8229,N_8000);
nand U8665 (N_8665,N_8097,N_8198);
xnor U8666 (N_8666,N_7818,N_7812);
and U8667 (N_8667,N_8034,N_8165);
xor U8668 (N_8668,N_8208,N_8193);
nand U8669 (N_8669,N_8305,N_7915);
nor U8670 (N_8670,N_7906,N_8153);
nor U8671 (N_8671,N_7830,N_8149);
and U8672 (N_8672,N_8235,N_8087);
xor U8673 (N_8673,N_8396,N_8273);
nand U8674 (N_8674,N_7994,N_8120);
nand U8675 (N_8675,N_8110,N_7942);
nor U8676 (N_8676,N_8038,N_8051);
and U8677 (N_8677,N_7986,N_8033);
and U8678 (N_8678,N_8354,N_8378);
nand U8679 (N_8679,N_8199,N_7984);
nand U8680 (N_8680,N_8074,N_7958);
nand U8681 (N_8681,N_8262,N_7901);
and U8682 (N_8682,N_8089,N_8004);
or U8683 (N_8683,N_7975,N_8241);
and U8684 (N_8684,N_8270,N_8349);
xor U8685 (N_8685,N_7872,N_7987);
and U8686 (N_8686,N_7970,N_7874);
or U8687 (N_8687,N_7939,N_8221);
and U8688 (N_8688,N_8214,N_8010);
xnor U8689 (N_8689,N_8351,N_7820);
nor U8690 (N_8690,N_7809,N_8163);
nand U8691 (N_8691,N_8381,N_7852);
xnor U8692 (N_8692,N_8180,N_8304);
nor U8693 (N_8693,N_7934,N_8092);
nor U8694 (N_8694,N_7845,N_8117);
or U8695 (N_8695,N_8015,N_8100);
xor U8696 (N_8696,N_8157,N_7877);
nand U8697 (N_8697,N_8127,N_7985);
nand U8698 (N_8698,N_8390,N_7982);
xor U8699 (N_8699,N_7878,N_8158);
xnor U8700 (N_8700,N_7956,N_7948);
xnor U8701 (N_8701,N_8010,N_8345);
and U8702 (N_8702,N_8283,N_8325);
nor U8703 (N_8703,N_7805,N_7963);
or U8704 (N_8704,N_8310,N_8204);
or U8705 (N_8705,N_7981,N_8232);
and U8706 (N_8706,N_8116,N_8210);
or U8707 (N_8707,N_7856,N_8226);
nor U8708 (N_8708,N_7898,N_8030);
and U8709 (N_8709,N_8107,N_8004);
and U8710 (N_8710,N_8046,N_8292);
nand U8711 (N_8711,N_8116,N_8384);
or U8712 (N_8712,N_8376,N_8307);
and U8713 (N_8713,N_8129,N_7920);
or U8714 (N_8714,N_8334,N_8354);
and U8715 (N_8715,N_7937,N_7920);
nor U8716 (N_8716,N_7888,N_8207);
nor U8717 (N_8717,N_8230,N_7864);
nand U8718 (N_8718,N_7879,N_8308);
or U8719 (N_8719,N_8334,N_8266);
xnor U8720 (N_8720,N_8336,N_7900);
nor U8721 (N_8721,N_7980,N_8312);
and U8722 (N_8722,N_7828,N_7814);
nor U8723 (N_8723,N_8244,N_8115);
xor U8724 (N_8724,N_8026,N_8010);
xnor U8725 (N_8725,N_8027,N_7968);
xor U8726 (N_8726,N_8109,N_8152);
or U8727 (N_8727,N_7892,N_8377);
nor U8728 (N_8728,N_8190,N_7887);
and U8729 (N_8729,N_7813,N_8105);
xnor U8730 (N_8730,N_8150,N_8357);
nor U8731 (N_8731,N_8030,N_8194);
xor U8732 (N_8732,N_8341,N_7933);
and U8733 (N_8733,N_8073,N_7964);
nand U8734 (N_8734,N_8356,N_8135);
xnor U8735 (N_8735,N_7856,N_8301);
or U8736 (N_8736,N_7948,N_8294);
nand U8737 (N_8737,N_8067,N_7910);
or U8738 (N_8738,N_7815,N_7865);
and U8739 (N_8739,N_7852,N_8129);
nand U8740 (N_8740,N_7822,N_8215);
nand U8741 (N_8741,N_7839,N_8394);
nand U8742 (N_8742,N_8383,N_7877);
nand U8743 (N_8743,N_8014,N_8004);
and U8744 (N_8744,N_7838,N_8376);
nand U8745 (N_8745,N_8160,N_8089);
xor U8746 (N_8746,N_8282,N_8243);
nand U8747 (N_8747,N_8342,N_8288);
nand U8748 (N_8748,N_7920,N_8031);
xor U8749 (N_8749,N_8165,N_7832);
or U8750 (N_8750,N_8041,N_8355);
nor U8751 (N_8751,N_8019,N_8080);
and U8752 (N_8752,N_8189,N_8384);
nor U8753 (N_8753,N_7811,N_8160);
or U8754 (N_8754,N_8074,N_7947);
xor U8755 (N_8755,N_8394,N_7837);
nand U8756 (N_8756,N_8335,N_7892);
nor U8757 (N_8757,N_7805,N_8123);
and U8758 (N_8758,N_8358,N_7909);
and U8759 (N_8759,N_8005,N_8143);
nor U8760 (N_8760,N_8193,N_8026);
and U8761 (N_8761,N_8378,N_8267);
and U8762 (N_8762,N_7944,N_8218);
or U8763 (N_8763,N_8222,N_8326);
nor U8764 (N_8764,N_8078,N_8357);
and U8765 (N_8765,N_8335,N_7805);
nor U8766 (N_8766,N_7983,N_8328);
xor U8767 (N_8767,N_7955,N_7823);
nor U8768 (N_8768,N_8362,N_7821);
nor U8769 (N_8769,N_8173,N_7814);
nand U8770 (N_8770,N_8190,N_7906);
xnor U8771 (N_8771,N_7836,N_7950);
nor U8772 (N_8772,N_7961,N_7907);
xor U8773 (N_8773,N_7808,N_8040);
nand U8774 (N_8774,N_8051,N_8028);
and U8775 (N_8775,N_7951,N_8231);
nand U8776 (N_8776,N_8297,N_8180);
or U8777 (N_8777,N_8329,N_7943);
nor U8778 (N_8778,N_8099,N_8297);
nor U8779 (N_8779,N_7978,N_8070);
and U8780 (N_8780,N_8028,N_8107);
xor U8781 (N_8781,N_7880,N_8174);
nand U8782 (N_8782,N_8353,N_8106);
xnor U8783 (N_8783,N_8305,N_7807);
nor U8784 (N_8784,N_8393,N_8179);
nor U8785 (N_8785,N_7822,N_8135);
and U8786 (N_8786,N_8124,N_7807);
or U8787 (N_8787,N_8161,N_7949);
and U8788 (N_8788,N_8081,N_8234);
nor U8789 (N_8789,N_8152,N_8313);
or U8790 (N_8790,N_7871,N_7852);
nor U8791 (N_8791,N_8267,N_8033);
or U8792 (N_8792,N_8176,N_7833);
nor U8793 (N_8793,N_7982,N_8259);
xor U8794 (N_8794,N_8139,N_8294);
xor U8795 (N_8795,N_8295,N_7900);
nor U8796 (N_8796,N_8172,N_8208);
nor U8797 (N_8797,N_7998,N_7893);
and U8798 (N_8798,N_8206,N_8383);
and U8799 (N_8799,N_7843,N_7892);
nand U8800 (N_8800,N_8080,N_8242);
nor U8801 (N_8801,N_8260,N_8028);
or U8802 (N_8802,N_8046,N_8247);
xor U8803 (N_8803,N_8260,N_7862);
or U8804 (N_8804,N_8006,N_8119);
nand U8805 (N_8805,N_8121,N_8376);
or U8806 (N_8806,N_8136,N_8205);
nor U8807 (N_8807,N_8364,N_8081);
xnor U8808 (N_8808,N_8115,N_7960);
nand U8809 (N_8809,N_8150,N_8240);
xor U8810 (N_8810,N_8380,N_8229);
or U8811 (N_8811,N_8161,N_8347);
nor U8812 (N_8812,N_8314,N_8146);
and U8813 (N_8813,N_8324,N_8394);
nand U8814 (N_8814,N_8394,N_7997);
xor U8815 (N_8815,N_7932,N_7942);
xor U8816 (N_8816,N_8107,N_7932);
nor U8817 (N_8817,N_7980,N_8060);
nand U8818 (N_8818,N_8294,N_8264);
and U8819 (N_8819,N_8392,N_8343);
nor U8820 (N_8820,N_8362,N_8080);
nand U8821 (N_8821,N_8230,N_8164);
xnor U8822 (N_8822,N_8100,N_7865);
and U8823 (N_8823,N_8040,N_8294);
nand U8824 (N_8824,N_8167,N_8130);
nor U8825 (N_8825,N_7800,N_7971);
nand U8826 (N_8826,N_8128,N_8112);
or U8827 (N_8827,N_8230,N_8070);
or U8828 (N_8828,N_7814,N_8209);
nand U8829 (N_8829,N_8169,N_8137);
xor U8830 (N_8830,N_7845,N_7973);
or U8831 (N_8831,N_7889,N_7920);
nand U8832 (N_8832,N_8193,N_7983);
or U8833 (N_8833,N_8052,N_8001);
or U8834 (N_8834,N_7954,N_8280);
nand U8835 (N_8835,N_8084,N_8024);
and U8836 (N_8836,N_8395,N_8138);
and U8837 (N_8837,N_8142,N_7851);
nand U8838 (N_8838,N_8255,N_7913);
nand U8839 (N_8839,N_8148,N_8337);
and U8840 (N_8840,N_8145,N_8046);
nand U8841 (N_8841,N_8063,N_7967);
xor U8842 (N_8842,N_7871,N_8019);
nor U8843 (N_8843,N_8311,N_8068);
and U8844 (N_8844,N_8194,N_8383);
xnor U8845 (N_8845,N_8073,N_8276);
nand U8846 (N_8846,N_7836,N_8005);
and U8847 (N_8847,N_8230,N_7875);
nand U8848 (N_8848,N_8063,N_8290);
xor U8849 (N_8849,N_7990,N_8382);
nor U8850 (N_8850,N_8185,N_8348);
xor U8851 (N_8851,N_8268,N_7808);
and U8852 (N_8852,N_8044,N_8205);
and U8853 (N_8853,N_8151,N_8164);
or U8854 (N_8854,N_8307,N_8036);
nor U8855 (N_8855,N_8217,N_7918);
nand U8856 (N_8856,N_8155,N_8361);
nor U8857 (N_8857,N_7852,N_7942);
and U8858 (N_8858,N_8163,N_7939);
and U8859 (N_8859,N_7984,N_8376);
and U8860 (N_8860,N_7964,N_8263);
xor U8861 (N_8861,N_7921,N_7815);
nand U8862 (N_8862,N_7941,N_7809);
xor U8863 (N_8863,N_8283,N_8049);
nand U8864 (N_8864,N_8304,N_7827);
or U8865 (N_8865,N_8261,N_7890);
and U8866 (N_8866,N_8116,N_7920);
xnor U8867 (N_8867,N_8189,N_8129);
nand U8868 (N_8868,N_8015,N_8240);
nand U8869 (N_8869,N_8342,N_8068);
xnor U8870 (N_8870,N_7857,N_8140);
xor U8871 (N_8871,N_7854,N_8232);
or U8872 (N_8872,N_8141,N_8062);
xnor U8873 (N_8873,N_8352,N_8295);
and U8874 (N_8874,N_8002,N_8011);
and U8875 (N_8875,N_7908,N_8321);
nor U8876 (N_8876,N_8289,N_8054);
xor U8877 (N_8877,N_8144,N_8152);
or U8878 (N_8878,N_8343,N_7898);
or U8879 (N_8879,N_7886,N_8107);
xor U8880 (N_8880,N_7800,N_8208);
xor U8881 (N_8881,N_8261,N_8042);
nand U8882 (N_8882,N_8213,N_8125);
nor U8883 (N_8883,N_8033,N_8283);
xor U8884 (N_8884,N_8024,N_7967);
nand U8885 (N_8885,N_8387,N_8385);
or U8886 (N_8886,N_8118,N_8211);
nand U8887 (N_8887,N_8132,N_8085);
nor U8888 (N_8888,N_8193,N_8233);
or U8889 (N_8889,N_8223,N_7817);
xnor U8890 (N_8890,N_8235,N_8096);
nor U8891 (N_8891,N_8138,N_8394);
or U8892 (N_8892,N_7908,N_7841);
nand U8893 (N_8893,N_8287,N_8336);
xnor U8894 (N_8894,N_8390,N_8392);
or U8895 (N_8895,N_8071,N_7879);
nand U8896 (N_8896,N_8312,N_7810);
xnor U8897 (N_8897,N_7854,N_8066);
nor U8898 (N_8898,N_7887,N_7976);
nand U8899 (N_8899,N_8060,N_8381);
nor U8900 (N_8900,N_8343,N_8055);
xnor U8901 (N_8901,N_7884,N_8377);
nand U8902 (N_8902,N_7924,N_7884);
xor U8903 (N_8903,N_8057,N_8394);
and U8904 (N_8904,N_8152,N_8362);
or U8905 (N_8905,N_7960,N_8387);
or U8906 (N_8906,N_7994,N_8279);
and U8907 (N_8907,N_8102,N_7928);
or U8908 (N_8908,N_8244,N_7911);
nor U8909 (N_8909,N_8070,N_7828);
xnor U8910 (N_8910,N_8371,N_7844);
nor U8911 (N_8911,N_7984,N_7913);
or U8912 (N_8912,N_8352,N_7829);
nand U8913 (N_8913,N_7903,N_7857);
and U8914 (N_8914,N_7925,N_7893);
or U8915 (N_8915,N_7981,N_8209);
nor U8916 (N_8916,N_8092,N_8108);
nand U8917 (N_8917,N_8274,N_8260);
or U8918 (N_8918,N_8213,N_7936);
xor U8919 (N_8919,N_7949,N_7817);
and U8920 (N_8920,N_8159,N_8178);
and U8921 (N_8921,N_8133,N_8039);
or U8922 (N_8922,N_8229,N_7939);
nand U8923 (N_8923,N_8393,N_7834);
xor U8924 (N_8924,N_8365,N_8033);
and U8925 (N_8925,N_7938,N_8291);
nor U8926 (N_8926,N_7886,N_7919);
or U8927 (N_8927,N_8321,N_8275);
xor U8928 (N_8928,N_7993,N_8232);
or U8929 (N_8929,N_7839,N_8264);
nor U8930 (N_8930,N_8348,N_7845);
xor U8931 (N_8931,N_8014,N_8010);
or U8932 (N_8932,N_8397,N_8262);
xor U8933 (N_8933,N_8236,N_8271);
and U8934 (N_8934,N_8297,N_7999);
and U8935 (N_8935,N_8358,N_8324);
and U8936 (N_8936,N_8148,N_8162);
and U8937 (N_8937,N_8109,N_8126);
nand U8938 (N_8938,N_8047,N_8069);
xor U8939 (N_8939,N_8141,N_8330);
and U8940 (N_8940,N_8299,N_8358);
nor U8941 (N_8941,N_8325,N_8290);
nand U8942 (N_8942,N_8377,N_8136);
or U8943 (N_8943,N_8122,N_7879);
nor U8944 (N_8944,N_7846,N_8217);
xnor U8945 (N_8945,N_8030,N_7865);
nor U8946 (N_8946,N_8001,N_8080);
or U8947 (N_8947,N_8326,N_8216);
or U8948 (N_8948,N_8087,N_8234);
and U8949 (N_8949,N_8221,N_8031);
nand U8950 (N_8950,N_8253,N_8308);
xnor U8951 (N_8951,N_7835,N_8339);
or U8952 (N_8952,N_7862,N_7874);
and U8953 (N_8953,N_8228,N_8284);
and U8954 (N_8954,N_8250,N_7905);
nor U8955 (N_8955,N_8247,N_7908);
nor U8956 (N_8956,N_7991,N_8241);
and U8957 (N_8957,N_7951,N_7874);
xnor U8958 (N_8958,N_8344,N_8216);
and U8959 (N_8959,N_8182,N_7935);
and U8960 (N_8960,N_7834,N_8283);
xor U8961 (N_8961,N_8176,N_7950);
or U8962 (N_8962,N_8000,N_8240);
xor U8963 (N_8963,N_8056,N_7962);
xor U8964 (N_8964,N_8147,N_8324);
xnor U8965 (N_8965,N_8145,N_7862);
nand U8966 (N_8966,N_8354,N_8194);
xnor U8967 (N_8967,N_7868,N_8064);
and U8968 (N_8968,N_8268,N_8173);
and U8969 (N_8969,N_8232,N_7875);
or U8970 (N_8970,N_7898,N_8370);
and U8971 (N_8971,N_8312,N_8067);
nor U8972 (N_8972,N_7840,N_8284);
nand U8973 (N_8973,N_7915,N_8196);
xnor U8974 (N_8974,N_8214,N_8371);
nor U8975 (N_8975,N_8370,N_7963);
nor U8976 (N_8976,N_7890,N_8227);
xor U8977 (N_8977,N_8146,N_8285);
xnor U8978 (N_8978,N_7975,N_8385);
or U8979 (N_8979,N_7915,N_8084);
or U8980 (N_8980,N_8259,N_8346);
or U8981 (N_8981,N_7965,N_7998);
or U8982 (N_8982,N_8295,N_8392);
nor U8983 (N_8983,N_7818,N_8389);
and U8984 (N_8984,N_7879,N_7993);
xor U8985 (N_8985,N_8378,N_7995);
nand U8986 (N_8986,N_7956,N_8263);
and U8987 (N_8987,N_8195,N_7957);
and U8988 (N_8988,N_8095,N_8219);
or U8989 (N_8989,N_8217,N_8339);
or U8990 (N_8990,N_7911,N_8066);
or U8991 (N_8991,N_8124,N_8009);
nor U8992 (N_8992,N_8158,N_8141);
xnor U8993 (N_8993,N_8377,N_8180);
nor U8994 (N_8994,N_8223,N_7811);
and U8995 (N_8995,N_8085,N_8398);
or U8996 (N_8996,N_8316,N_8268);
nor U8997 (N_8997,N_8011,N_7943);
or U8998 (N_8998,N_8315,N_8113);
nand U8999 (N_8999,N_8040,N_7922);
nor U9000 (N_9000,N_8532,N_8546);
xnor U9001 (N_9001,N_8442,N_8571);
or U9002 (N_9002,N_8488,N_8435);
and U9003 (N_9003,N_8632,N_8906);
xor U9004 (N_9004,N_8612,N_8425);
xnor U9005 (N_9005,N_8477,N_8835);
nor U9006 (N_9006,N_8625,N_8930);
nor U9007 (N_9007,N_8826,N_8588);
nand U9008 (N_9008,N_8815,N_8418);
xnor U9009 (N_9009,N_8499,N_8963);
nor U9010 (N_9010,N_8730,N_8807);
nor U9011 (N_9011,N_8973,N_8735);
nor U9012 (N_9012,N_8829,N_8616);
nor U9013 (N_9013,N_8522,N_8479);
nor U9014 (N_9014,N_8689,N_8832);
nand U9015 (N_9015,N_8683,N_8590);
nor U9016 (N_9016,N_8657,N_8461);
and U9017 (N_9017,N_8905,N_8605);
or U9018 (N_9018,N_8794,N_8959);
nor U9019 (N_9019,N_8989,N_8961);
nand U9020 (N_9020,N_8766,N_8878);
xnor U9021 (N_9021,N_8814,N_8551);
and U9022 (N_9022,N_8548,N_8437);
xor U9023 (N_9023,N_8604,N_8646);
xor U9024 (N_9024,N_8473,N_8898);
and U9025 (N_9025,N_8462,N_8861);
or U9026 (N_9026,N_8642,N_8708);
and U9027 (N_9027,N_8534,N_8446);
and U9028 (N_9028,N_8744,N_8500);
or U9029 (N_9029,N_8860,N_8764);
nand U9030 (N_9030,N_8851,N_8609);
xnor U9031 (N_9031,N_8809,N_8748);
nor U9032 (N_9032,N_8990,N_8909);
or U9033 (N_9033,N_8677,N_8515);
nand U9034 (N_9034,N_8722,N_8570);
and U9035 (N_9035,N_8638,N_8673);
or U9036 (N_9036,N_8426,N_8767);
xor U9037 (N_9037,N_8793,N_8816);
xnor U9038 (N_9038,N_8402,N_8541);
xnor U9039 (N_9039,N_8576,N_8664);
and U9040 (N_9040,N_8801,N_8684);
nand U9041 (N_9041,N_8456,N_8536);
nor U9042 (N_9042,N_8650,N_8624);
nand U9043 (N_9043,N_8655,N_8465);
xor U9044 (N_9044,N_8406,N_8769);
nor U9045 (N_9045,N_8804,N_8935);
nor U9046 (N_9046,N_8928,N_8792);
or U9047 (N_9047,N_8439,N_8666);
and U9048 (N_9048,N_8892,N_8981);
xor U9049 (N_9049,N_8692,N_8954);
xor U9050 (N_9050,N_8450,N_8608);
or U9051 (N_9051,N_8503,N_8926);
nor U9052 (N_9052,N_8466,N_8485);
xor U9053 (N_9053,N_8760,N_8552);
nor U9054 (N_9054,N_8537,N_8510);
and U9055 (N_9055,N_8951,N_8988);
xnor U9056 (N_9056,N_8824,N_8920);
nand U9057 (N_9057,N_8888,N_8698);
or U9058 (N_9058,N_8429,N_8980);
nand U9059 (N_9059,N_8753,N_8413);
nand U9060 (N_9060,N_8563,N_8535);
xnor U9061 (N_9061,N_8583,N_8617);
or U9062 (N_9062,N_8797,N_8978);
nand U9063 (N_9063,N_8498,N_8452);
nand U9064 (N_9064,N_8490,N_8607);
and U9065 (N_9065,N_8676,N_8433);
or U9066 (N_9066,N_8436,N_8484);
nor U9067 (N_9067,N_8560,N_8717);
or U9068 (N_9068,N_8780,N_8486);
nand U9069 (N_9069,N_8886,N_8525);
nor U9070 (N_9070,N_8697,N_8471);
and U9071 (N_9071,N_8595,N_8953);
and U9072 (N_9072,N_8745,N_8724);
nor U9073 (N_9073,N_8983,N_8428);
xnor U9074 (N_9074,N_8416,N_8995);
nand U9075 (N_9075,N_8977,N_8845);
and U9076 (N_9076,N_8573,N_8670);
or U9077 (N_9077,N_8514,N_8755);
xnor U9078 (N_9078,N_8825,N_8787);
nor U9079 (N_9079,N_8915,N_8687);
nand U9080 (N_9080,N_8774,N_8979);
nand U9081 (N_9081,N_8672,N_8727);
nand U9082 (N_9082,N_8876,N_8508);
xor U9083 (N_9083,N_8476,N_8518);
nor U9084 (N_9084,N_8715,N_8934);
nand U9085 (N_9085,N_8858,N_8564);
nor U9086 (N_9086,N_8709,N_8547);
nand U9087 (N_9087,N_8771,N_8946);
and U9088 (N_9088,N_8740,N_8529);
nand U9089 (N_9089,N_8736,N_8719);
nor U9090 (N_9090,N_8955,N_8495);
or U9091 (N_9091,N_8584,N_8778);
nand U9092 (N_9092,N_8966,N_8555);
xor U9093 (N_9093,N_8678,N_8985);
or U9094 (N_9094,N_8480,N_8649);
xor U9095 (N_9095,N_8893,N_8663);
nand U9096 (N_9096,N_8732,N_8516);
xor U9097 (N_9097,N_8455,N_8422);
nor U9098 (N_9098,N_8941,N_8540);
xnor U9099 (N_9099,N_8854,N_8613);
or U9100 (N_9100,N_8901,N_8621);
and U9101 (N_9101,N_8531,N_8772);
nand U9102 (N_9102,N_8943,N_8820);
and U9103 (N_9103,N_8556,N_8836);
and U9104 (N_9104,N_8526,N_8773);
nor U9105 (N_9105,N_8883,N_8958);
or U9106 (N_9106,N_8833,N_8937);
nor U9107 (N_9107,N_8568,N_8759);
xnor U9108 (N_9108,N_8700,N_8743);
xor U9109 (N_9109,N_8411,N_8770);
nand U9110 (N_9110,N_8523,N_8630);
and U9111 (N_9111,N_8427,N_8862);
or U9112 (N_9112,N_8999,N_8566);
or U9113 (N_9113,N_8817,N_8492);
xnor U9114 (N_9114,N_8972,N_8493);
and U9115 (N_9115,N_8931,N_8574);
nand U9116 (N_9116,N_8749,N_8636);
nand U9117 (N_9117,N_8579,N_8661);
or U9118 (N_9118,N_8970,N_8502);
nand U9119 (N_9119,N_8557,N_8856);
xor U9120 (N_9120,N_8589,N_8762);
and U9121 (N_9121,N_8631,N_8713);
nor U9122 (N_9122,N_8728,N_8671);
nand U9123 (N_9123,N_8783,N_8553);
xnor U9124 (N_9124,N_8731,N_8877);
or U9125 (N_9125,N_8790,N_8592);
nor U9126 (N_9126,N_8599,N_8795);
xnor U9127 (N_9127,N_8582,N_8469);
nor U9128 (N_9128,N_8738,N_8847);
or U9129 (N_9129,N_8414,N_8751);
and U9130 (N_9130,N_8662,N_8850);
and U9131 (N_9131,N_8975,N_8470);
or U9132 (N_9132,N_8761,N_8707);
nor U9133 (N_9133,N_8887,N_8725);
nand U9134 (N_9134,N_8947,N_8453);
xor U9135 (N_9135,N_8869,N_8782);
and U9136 (N_9136,N_8705,N_8902);
nor U9137 (N_9137,N_8412,N_8859);
nand U9138 (N_9138,N_8458,N_8781);
xor U9139 (N_9139,N_8944,N_8994);
and U9140 (N_9140,N_8965,N_8679);
xnor U9141 (N_9141,N_8581,N_8597);
nor U9142 (N_9142,N_8596,N_8936);
nand U9143 (N_9143,N_8550,N_8483);
nand U9144 (N_9144,N_8496,N_8565);
and U9145 (N_9145,N_8948,N_8842);
xor U9146 (N_9146,N_8474,N_8885);
xor U9147 (N_9147,N_8441,N_8976);
nand U9148 (N_9148,N_8921,N_8598);
and U9149 (N_9149,N_8415,N_8643);
xnor U9150 (N_9150,N_8424,N_8665);
and U9151 (N_9151,N_8688,N_8704);
or U9152 (N_9152,N_8494,N_8680);
and U9153 (N_9153,N_8559,N_8695);
and U9154 (N_9154,N_8945,N_8964);
or U9155 (N_9155,N_8667,N_8996);
nor U9156 (N_9156,N_8949,N_8932);
nor U9157 (N_9157,N_8528,N_8606);
nand U9158 (N_9158,N_8897,N_8784);
and U9159 (N_9159,N_8669,N_8530);
xor U9160 (N_9160,N_8501,N_8660);
and U9161 (N_9161,N_8940,N_8626);
xor U9162 (N_9162,N_8635,N_8448);
or U9163 (N_9163,N_8591,N_8992);
nand U9164 (N_9164,N_8711,N_8871);
or U9165 (N_9165,N_8813,N_8545);
nand U9166 (N_9166,N_8524,N_8870);
or U9167 (N_9167,N_8447,N_8777);
or U9168 (N_9168,N_8974,N_8923);
nand U9169 (N_9169,N_8925,N_8723);
nand U9170 (N_9170,N_8916,N_8853);
nand U9171 (N_9171,N_8800,N_8648);
or U9172 (N_9172,N_8637,N_8475);
and U9173 (N_9173,N_8880,N_8873);
nor U9174 (N_9174,N_8913,N_8747);
nand U9175 (N_9175,N_8575,N_8789);
or U9176 (N_9176,N_8417,N_8865);
or U9177 (N_9177,N_8868,N_8844);
or U9178 (N_9178,N_8806,N_8910);
nor U9179 (N_9179,N_8758,N_8796);
xor U9180 (N_9180,N_8400,N_8714);
or U9181 (N_9181,N_8968,N_8681);
nor U9182 (N_9182,N_8997,N_8544);
nor U9183 (N_9183,N_8984,N_8504);
or U9184 (N_9184,N_8757,N_8918);
xor U9185 (N_9185,N_8633,N_8879);
xnor U9186 (N_9186,N_8481,N_8939);
or U9187 (N_9187,N_8721,N_8701);
or U9188 (N_9188,N_8752,N_8419);
nand U9189 (N_9189,N_8423,N_8520);
nand U9190 (N_9190,N_8691,N_8644);
xor U9191 (N_9191,N_8699,N_8962);
or U9192 (N_9192,N_8942,N_8432);
and U9193 (N_9193,N_8924,N_8952);
nand U9194 (N_9194,N_8658,N_8956);
or U9195 (N_9195,N_8614,N_8449);
nor U9196 (N_9196,N_8487,N_8726);
nand U9197 (N_9197,N_8686,N_8497);
or U9198 (N_9198,N_8933,N_8899);
nor U9199 (N_9199,N_8750,N_8656);
xnor U9200 (N_9200,N_8907,N_8776);
and U9201 (N_9201,N_8830,N_8640);
nor U9202 (N_9202,N_8538,N_8706);
nor U9203 (N_9203,N_8875,N_8652);
xor U9204 (N_9204,N_8690,N_8653);
and U9205 (N_9205,N_8615,N_8857);
nor U9206 (N_9206,N_8603,N_8840);
nor U9207 (N_9207,N_8443,N_8622);
nand U9208 (N_9208,N_8867,N_8927);
or U9209 (N_9209,N_8512,N_8950);
xor U9210 (N_9210,N_8505,N_8912);
nor U9211 (N_9211,N_8601,N_8779);
nand U9212 (N_9212,N_8693,N_8872);
nand U9213 (N_9213,N_8982,N_8506);
and U9214 (N_9214,N_8756,N_8710);
or U9215 (N_9215,N_8403,N_8929);
nor U9216 (N_9216,N_8464,N_8517);
or U9217 (N_9217,N_8737,N_8874);
nand U9218 (N_9218,N_8408,N_8482);
nand U9219 (N_9219,N_8729,N_8908);
xnor U9220 (N_9220,N_8647,N_8957);
and U9221 (N_9221,N_8986,N_8739);
xor U9222 (N_9222,N_8866,N_8472);
nor U9223 (N_9223,N_8821,N_8884);
or U9224 (N_9224,N_8463,N_8562);
xor U9225 (N_9225,N_8991,N_8572);
and U9226 (N_9226,N_8651,N_8919);
or U9227 (N_9227,N_8914,N_8827);
nor U9228 (N_9228,N_8768,N_8539);
nand U9229 (N_9229,N_8716,N_8900);
nor U9230 (N_9230,N_8467,N_8685);
nor U9231 (N_9231,N_8491,N_8839);
nand U9232 (N_9232,N_8527,N_8468);
or U9233 (N_9233,N_8533,N_8519);
or U9234 (N_9234,N_8846,N_8430);
and U9235 (N_9235,N_8855,N_8803);
nand U9236 (N_9236,N_8788,N_8863);
and U9237 (N_9237,N_8746,N_8712);
and U9238 (N_9238,N_8852,N_8754);
xor U9239 (N_9239,N_8401,N_8922);
and U9240 (N_9240,N_8421,N_8405);
xor U9241 (N_9241,N_8993,N_8831);
nor U9242 (N_9242,N_8967,N_8882);
nor U9243 (N_9243,N_8460,N_8577);
or U9244 (N_9244,N_8513,N_8620);
nand U9245 (N_9245,N_8849,N_8542);
xor U9246 (N_9246,N_8785,N_8628);
nand U9247 (N_9247,N_8805,N_8811);
xnor U9248 (N_9248,N_8521,N_8627);
nand U9249 (N_9249,N_8702,N_8509);
nor U9250 (N_9250,N_8610,N_8654);
xor U9251 (N_9251,N_8798,N_8420);
and U9252 (N_9252,N_8763,N_8511);
and U9253 (N_9253,N_8543,N_8822);
xor U9254 (N_9254,N_8799,N_8602);
nor U9255 (N_9255,N_8791,N_8634);
xor U9256 (N_9256,N_8587,N_8765);
nor U9257 (N_9257,N_8434,N_8600);
nand U9258 (N_9258,N_8733,N_8734);
xor U9259 (N_9259,N_8478,N_8404);
and U9260 (N_9260,N_8969,N_8549);
nor U9261 (N_9261,N_8457,N_8742);
xnor U9262 (N_9262,N_8489,N_8623);
and U9263 (N_9263,N_8558,N_8645);
and U9264 (N_9264,N_8819,N_8694);
or U9265 (N_9265,N_8911,N_8554);
or U9266 (N_9266,N_8881,N_8864);
nor U9267 (N_9267,N_8838,N_8834);
nand U9268 (N_9268,N_8889,N_8903);
and U9269 (N_9269,N_8438,N_8917);
nor U9270 (N_9270,N_8444,N_8775);
nand U9271 (N_9271,N_8998,N_8585);
nor U9272 (N_9272,N_8431,N_8703);
xor U9273 (N_9273,N_8823,N_8629);
and U9274 (N_9274,N_8802,N_8682);
and U9275 (N_9275,N_8741,N_8812);
nor U9276 (N_9276,N_8561,N_8810);
nor U9277 (N_9277,N_8459,N_8674);
or U9278 (N_9278,N_8454,N_8619);
and U9279 (N_9279,N_8593,N_8569);
xnor U9280 (N_9280,N_8639,N_8938);
and U9281 (N_9281,N_8507,N_8837);
and U9282 (N_9282,N_8843,N_8578);
xnor U9283 (N_9283,N_8904,N_8718);
nand U9284 (N_9284,N_8567,N_8828);
nand U9285 (N_9285,N_8818,N_8987);
or U9286 (N_9286,N_8786,N_8407);
nor U9287 (N_9287,N_8960,N_8440);
xor U9288 (N_9288,N_8586,N_8594);
nor U9289 (N_9289,N_8410,N_8720);
xor U9290 (N_9290,N_8891,N_8971);
nor U9291 (N_9291,N_8580,N_8696);
xor U9292 (N_9292,N_8841,N_8451);
or U9293 (N_9293,N_8894,N_8896);
nor U9294 (N_9294,N_8611,N_8659);
xnor U9295 (N_9295,N_8409,N_8668);
nand U9296 (N_9296,N_8848,N_8675);
or U9297 (N_9297,N_8445,N_8808);
nor U9298 (N_9298,N_8890,N_8641);
nor U9299 (N_9299,N_8618,N_8895);
nor U9300 (N_9300,N_8686,N_8805);
nand U9301 (N_9301,N_8617,N_8667);
nand U9302 (N_9302,N_8645,N_8995);
nand U9303 (N_9303,N_8568,N_8496);
nand U9304 (N_9304,N_8483,N_8515);
xor U9305 (N_9305,N_8479,N_8764);
and U9306 (N_9306,N_8485,N_8651);
nand U9307 (N_9307,N_8970,N_8721);
nor U9308 (N_9308,N_8977,N_8937);
and U9309 (N_9309,N_8614,N_8991);
nand U9310 (N_9310,N_8912,N_8737);
and U9311 (N_9311,N_8609,N_8440);
nor U9312 (N_9312,N_8795,N_8955);
nor U9313 (N_9313,N_8504,N_8555);
xor U9314 (N_9314,N_8813,N_8948);
or U9315 (N_9315,N_8783,N_8551);
nor U9316 (N_9316,N_8861,N_8585);
nand U9317 (N_9317,N_8676,N_8688);
nor U9318 (N_9318,N_8931,N_8635);
xnor U9319 (N_9319,N_8472,N_8988);
or U9320 (N_9320,N_8854,N_8563);
nand U9321 (N_9321,N_8635,N_8411);
and U9322 (N_9322,N_8676,N_8847);
nand U9323 (N_9323,N_8954,N_8739);
or U9324 (N_9324,N_8846,N_8999);
or U9325 (N_9325,N_8491,N_8727);
nor U9326 (N_9326,N_8584,N_8601);
nand U9327 (N_9327,N_8702,N_8954);
or U9328 (N_9328,N_8998,N_8779);
nor U9329 (N_9329,N_8965,N_8528);
nor U9330 (N_9330,N_8794,N_8934);
or U9331 (N_9331,N_8573,N_8434);
nor U9332 (N_9332,N_8578,N_8979);
and U9333 (N_9333,N_8875,N_8768);
nand U9334 (N_9334,N_8996,N_8934);
or U9335 (N_9335,N_8929,N_8863);
nand U9336 (N_9336,N_8583,N_8516);
and U9337 (N_9337,N_8641,N_8428);
nor U9338 (N_9338,N_8560,N_8666);
nand U9339 (N_9339,N_8534,N_8641);
and U9340 (N_9340,N_8705,N_8410);
or U9341 (N_9341,N_8473,N_8436);
and U9342 (N_9342,N_8604,N_8920);
nor U9343 (N_9343,N_8756,N_8989);
and U9344 (N_9344,N_8511,N_8412);
nand U9345 (N_9345,N_8408,N_8452);
xnor U9346 (N_9346,N_8705,N_8889);
and U9347 (N_9347,N_8522,N_8448);
nor U9348 (N_9348,N_8623,N_8795);
or U9349 (N_9349,N_8716,N_8579);
nor U9350 (N_9350,N_8557,N_8603);
nand U9351 (N_9351,N_8441,N_8516);
nand U9352 (N_9352,N_8708,N_8502);
and U9353 (N_9353,N_8825,N_8896);
and U9354 (N_9354,N_8504,N_8798);
xnor U9355 (N_9355,N_8837,N_8411);
nor U9356 (N_9356,N_8452,N_8728);
nand U9357 (N_9357,N_8931,N_8893);
nor U9358 (N_9358,N_8795,N_8908);
nand U9359 (N_9359,N_8956,N_8784);
nor U9360 (N_9360,N_8635,N_8531);
or U9361 (N_9361,N_8451,N_8514);
nor U9362 (N_9362,N_8407,N_8657);
nor U9363 (N_9363,N_8637,N_8724);
or U9364 (N_9364,N_8679,N_8865);
nor U9365 (N_9365,N_8780,N_8429);
nand U9366 (N_9366,N_8989,N_8649);
nand U9367 (N_9367,N_8874,N_8978);
or U9368 (N_9368,N_8582,N_8875);
and U9369 (N_9369,N_8748,N_8672);
nor U9370 (N_9370,N_8984,N_8465);
xnor U9371 (N_9371,N_8633,N_8887);
nor U9372 (N_9372,N_8562,N_8428);
and U9373 (N_9373,N_8710,N_8727);
or U9374 (N_9374,N_8578,N_8569);
xor U9375 (N_9375,N_8863,N_8473);
and U9376 (N_9376,N_8614,N_8915);
or U9377 (N_9377,N_8567,N_8470);
nor U9378 (N_9378,N_8992,N_8457);
or U9379 (N_9379,N_8405,N_8435);
or U9380 (N_9380,N_8994,N_8886);
nand U9381 (N_9381,N_8539,N_8658);
or U9382 (N_9382,N_8983,N_8840);
and U9383 (N_9383,N_8469,N_8848);
and U9384 (N_9384,N_8924,N_8697);
nand U9385 (N_9385,N_8741,N_8636);
and U9386 (N_9386,N_8446,N_8513);
and U9387 (N_9387,N_8985,N_8755);
nor U9388 (N_9388,N_8454,N_8880);
and U9389 (N_9389,N_8536,N_8448);
nand U9390 (N_9390,N_8907,N_8515);
xor U9391 (N_9391,N_8415,N_8512);
or U9392 (N_9392,N_8429,N_8884);
and U9393 (N_9393,N_8437,N_8776);
xor U9394 (N_9394,N_8990,N_8531);
nand U9395 (N_9395,N_8756,N_8800);
or U9396 (N_9396,N_8795,N_8778);
nand U9397 (N_9397,N_8803,N_8563);
nand U9398 (N_9398,N_8810,N_8548);
and U9399 (N_9399,N_8550,N_8646);
and U9400 (N_9400,N_8870,N_8832);
xnor U9401 (N_9401,N_8442,N_8416);
and U9402 (N_9402,N_8865,N_8496);
xor U9403 (N_9403,N_8685,N_8783);
and U9404 (N_9404,N_8757,N_8574);
nand U9405 (N_9405,N_8706,N_8557);
and U9406 (N_9406,N_8451,N_8733);
and U9407 (N_9407,N_8908,N_8941);
or U9408 (N_9408,N_8974,N_8588);
xor U9409 (N_9409,N_8490,N_8569);
and U9410 (N_9410,N_8769,N_8404);
xor U9411 (N_9411,N_8460,N_8744);
or U9412 (N_9412,N_8527,N_8542);
nand U9413 (N_9413,N_8466,N_8642);
nor U9414 (N_9414,N_8578,N_8614);
xnor U9415 (N_9415,N_8623,N_8453);
nand U9416 (N_9416,N_8957,N_8699);
nand U9417 (N_9417,N_8901,N_8726);
xor U9418 (N_9418,N_8715,N_8846);
xnor U9419 (N_9419,N_8758,N_8753);
nor U9420 (N_9420,N_8637,N_8694);
xor U9421 (N_9421,N_8906,N_8950);
nand U9422 (N_9422,N_8930,N_8638);
xor U9423 (N_9423,N_8947,N_8553);
nor U9424 (N_9424,N_8803,N_8760);
nand U9425 (N_9425,N_8903,N_8450);
xor U9426 (N_9426,N_8552,N_8410);
or U9427 (N_9427,N_8433,N_8680);
nand U9428 (N_9428,N_8725,N_8690);
nand U9429 (N_9429,N_8996,N_8498);
or U9430 (N_9430,N_8753,N_8865);
nand U9431 (N_9431,N_8470,N_8658);
nor U9432 (N_9432,N_8991,N_8659);
nand U9433 (N_9433,N_8638,N_8460);
and U9434 (N_9434,N_8866,N_8910);
or U9435 (N_9435,N_8431,N_8548);
or U9436 (N_9436,N_8959,N_8676);
nor U9437 (N_9437,N_8809,N_8594);
nand U9438 (N_9438,N_8962,N_8970);
nand U9439 (N_9439,N_8810,N_8824);
or U9440 (N_9440,N_8749,N_8457);
nor U9441 (N_9441,N_8500,N_8945);
nor U9442 (N_9442,N_8498,N_8594);
or U9443 (N_9443,N_8545,N_8423);
nor U9444 (N_9444,N_8643,N_8623);
or U9445 (N_9445,N_8492,N_8749);
nand U9446 (N_9446,N_8614,N_8928);
nand U9447 (N_9447,N_8873,N_8941);
xnor U9448 (N_9448,N_8536,N_8463);
and U9449 (N_9449,N_8900,N_8842);
nor U9450 (N_9450,N_8762,N_8668);
nand U9451 (N_9451,N_8601,N_8900);
nand U9452 (N_9452,N_8571,N_8930);
nand U9453 (N_9453,N_8869,N_8867);
nor U9454 (N_9454,N_8639,N_8778);
xnor U9455 (N_9455,N_8851,N_8415);
nor U9456 (N_9456,N_8614,N_8751);
and U9457 (N_9457,N_8430,N_8473);
nor U9458 (N_9458,N_8675,N_8600);
nor U9459 (N_9459,N_8517,N_8890);
or U9460 (N_9460,N_8647,N_8780);
or U9461 (N_9461,N_8500,N_8859);
or U9462 (N_9462,N_8941,N_8944);
or U9463 (N_9463,N_8670,N_8798);
nand U9464 (N_9464,N_8763,N_8925);
or U9465 (N_9465,N_8747,N_8965);
nand U9466 (N_9466,N_8498,N_8984);
or U9467 (N_9467,N_8642,N_8490);
xnor U9468 (N_9468,N_8694,N_8533);
nor U9469 (N_9469,N_8863,N_8793);
nand U9470 (N_9470,N_8446,N_8716);
xor U9471 (N_9471,N_8920,N_8955);
xnor U9472 (N_9472,N_8670,N_8501);
xor U9473 (N_9473,N_8938,N_8582);
nor U9474 (N_9474,N_8853,N_8522);
nand U9475 (N_9475,N_8431,N_8669);
or U9476 (N_9476,N_8797,N_8696);
or U9477 (N_9477,N_8645,N_8832);
and U9478 (N_9478,N_8629,N_8574);
nor U9479 (N_9479,N_8844,N_8803);
xnor U9480 (N_9480,N_8476,N_8683);
xnor U9481 (N_9481,N_8709,N_8725);
nand U9482 (N_9482,N_8777,N_8762);
nand U9483 (N_9483,N_8551,N_8561);
xor U9484 (N_9484,N_8542,N_8887);
nand U9485 (N_9485,N_8775,N_8642);
xor U9486 (N_9486,N_8429,N_8500);
xor U9487 (N_9487,N_8780,N_8456);
nor U9488 (N_9488,N_8637,N_8877);
nor U9489 (N_9489,N_8477,N_8847);
and U9490 (N_9490,N_8939,N_8828);
xnor U9491 (N_9491,N_8758,N_8628);
nor U9492 (N_9492,N_8644,N_8559);
nand U9493 (N_9493,N_8735,N_8402);
nand U9494 (N_9494,N_8766,N_8521);
nand U9495 (N_9495,N_8626,N_8854);
xnor U9496 (N_9496,N_8515,N_8918);
and U9497 (N_9497,N_8927,N_8841);
or U9498 (N_9498,N_8701,N_8832);
or U9499 (N_9499,N_8523,N_8547);
xor U9500 (N_9500,N_8754,N_8522);
or U9501 (N_9501,N_8426,N_8529);
and U9502 (N_9502,N_8980,N_8851);
nand U9503 (N_9503,N_8840,N_8513);
or U9504 (N_9504,N_8867,N_8800);
and U9505 (N_9505,N_8469,N_8591);
nand U9506 (N_9506,N_8864,N_8654);
nor U9507 (N_9507,N_8732,N_8512);
nand U9508 (N_9508,N_8452,N_8532);
and U9509 (N_9509,N_8456,N_8777);
or U9510 (N_9510,N_8743,N_8678);
nor U9511 (N_9511,N_8486,N_8734);
nand U9512 (N_9512,N_8715,N_8873);
nand U9513 (N_9513,N_8753,N_8959);
or U9514 (N_9514,N_8782,N_8933);
nor U9515 (N_9515,N_8507,N_8468);
xor U9516 (N_9516,N_8742,N_8462);
or U9517 (N_9517,N_8912,N_8805);
and U9518 (N_9518,N_8680,N_8576);
nor U9519 (N_9519,N_8793,N_8627);
xor U9520 (N_9520,N_8506,N_8622);
xnor U9521 (N_9521,N_8635,N_8499);
nor U9522 (N_9522,N_8713,N_8824);
and U9523 (N_9523,N_8606,N_8889);
or U9524 (N_9524,N_8627,N_8613);
and U9525 (N_9525,N_8663,N_8961);
or U9526 (N_9526,N_8628,N_8903);
and U9527 (N_9527,N_8406,N_8635);
nand U9528 (N_9528,N_8575,N_8401);
or U9529 (N_9529,N_8808,N_8553);
nor U9530 (N_9530,N_8940,N_8779);
nand U9531 (N_9531,N_8489,N_8673);
or U9532 (N_9532,N_8972,N_8907);
nor U9533 (N_9533,N_8591,N_8758);
or U9534 (N_9534,N_8522,N_8492);
nor U9535 (N_9535,N_8539,N_8619);
or U9536 (N_9536,N_8727,N_8685);
nand U9537 (N_9537,N_8525,N_8943);
nand U9538 (N_9538,N_8786,N_8806);
or U9539 (N_9539,N_8779,N_8944);
nor U9540 (N_9540,N_8518,N_8975);
or U9541 (N_9541,N_8952,N_8418);
nand U9542 (N_9542,N_8940,N_8965);
nand U9543 (N_9543,N_8866,N_8502);
xnor U9544 (N_9544,N_8548,N_8711);
nor U9545 (N_9545,N_8816,N_8548);
xor U9546 (N_9546,N_8755,N_8867);
and U9547 (N_9547,N_8461,N_8744);
xnor U9548 (N_9548,N_8977,N_8870);
and U9549 (N_9549,N_8554,N_8888);
xnor U9550 (N_9550,N_8831,N_8589);
nor U9551 (N_9551,N_8740,N_8926);
or U9552 (N_9552,N_8426,N_8473);
and U9553 (N_9553,N_8442,N_8455);
nand U9554 (N_9554,N_8662,N_8417);
and U9555 (N_9555,N_8527,N_8936);
or U9556 (N_9556,N_8538,N_8691);
and U9557 (N_9557,N_8755,N_8722);
xor U9558 (N_9558,N_8765,N_8792);
xnor U9559 (N_9559,N_8632,N_8502);
nand U9560 (N_9560,N_8909,N_8882);
nor U9561 (N_9561,N_8684,N_8751);
or U9562 (N_9562,N_8847,N_8732);
or U9563 (N_9563,N_8978,N_8435);
and U9564 (N_9564,N_8468,N_8939);
nor U9565 (N_9565,N_8806,N_8606);
or U9566 (N_9566,N_8952,N_8953);
nand U9567 (N_9567,N_8827,N_8531);
nor U9568 (N_9568,N_8895,N_8590);
nand U9569 (N_9569,N_8769,N_8909);
nand U9570 (N_9570,N_8843,N_8486);
xnor U9571 (N_9571,N_8400,N_8818);
xnor U9572 (N_9572,N_8539,N_8678);
and U9573 (N_9573,N_8505,N_8615);
or U9574 (N_9574,N_8905,N_8440);
xnor U9575 (N_9575,N_8530,N_8915);
xnor U9576 (N_9576,N_8957,N_8708);
nor U9577 (N_9577,N_8984,N_8649);
or U9578 (N_9578,N_8502,N_8843);
nor U9579 (N_9579,N_8412,N_8818);
nand U9580 (N_9580,N_8585,N_8689);
xor U9581 (N_9581,N_8946,N_8754);
or U9582 (N_9582,N_8409,N_8708);
and U9583 (N_9583,N_8879,N_8728);
nor U9584 (N_9584,N_8669,N_8443);
or U9585 (N_9585,N_8470,N_8527);
or U9586 (N_9586,N_8698,N_8514);
nor U9587 (N_9587,N_8418,N_8944);
or U9588 (N_9588,N_8700,N_8522);
xor U9589 (N_9589,N_8902,N_8718);
nand U9590 (N_9590,N_8935,N_8444);
xnor U9591 (N_9591,N_8504,N_8459);
or U9592 (N_9592,N_8971,N_8402);
nand U9593 (N_9593,N_8529,N_8448);
xor U9594 (N_9594,N_8586,N_8931);
nand U9595 (N_9595,N_8775,N_8565);
nand U9596 (N_9596,N_8613,N_8941);
xnor U9597 (N_9597,N_8627,N_8581);
nor U9598 (N_9598,N_8435,N_8610);
and U9599 (N_9599,N_8752,N_8965);
xnor U9600 (N_9600,N_9337,N_9253);
xnor U9601 (N_9601,N_9343,N_9131);
nand U9602 (N_9602,N_9298,N_9536);
nor U9603 (N_9603,N_9501,N_9290);
and U9604 (N_9604,N_9202,N_9389);
xor U9605 (N_9605,N_9418,N_9005);
nor U9606 (N_9606,N_9361,N_9270);
xnor U9607 (N_9607,N_9106,N_9488);
xor U9608 (N_9608,N_9257,N_9365);
or U9609 (N_9609,N_9357,N_9232);
and U9610 (N_9610,N_9380,N_9109);
and U9611 (N_9611,N_9024,N_9540);
nor U9612 (N_9612,N_9555,N_9471);
xnor U9613 (N_9613,N_9146,N_9420);
nand U9614 (N_9614,N_9514,N_9563);
xor U9615 (N_9615,N_9165,N_9414);
and U9616 (N_9616,N_9523,N_9020);
and U9617 (N_9617,N_9546,N_9276);
xnor U9618 (N_9618,N_9396,N_9511);
xor U9619 (N_9619,N_9537,N_9338);
nand U9620 (N_9620,N_9522,N_9599);
nor U9621 (N_9621,N_9325,N_9272);
and U9622 (N_9622,N_9056,N_9311);
and U9623 (N_9623,N_9271,N_9332);
or U9624 (N_9624,N_9558,N_9138);
nor U9625 (N_9625,N_9330,N_9196);
nand U9626 (N_9626,N_9499,N_9076);
nor U9627 (N_9627,N_9370,N_9044);
nor U9628 (N_9628,N_9513,N_9541);
nor U9629 (N_9629,N_9309,N_9548);
and U9630 (N_9630,N_9463,N_9022);
nand U9631 (N_9631,N_9391,N_9144);
nor U9632 (N_9632,N_9326,N_9207);
and U9633 (N_9633,N_9063,N_9034);
nor U9634 (N_9634,N_9426,N_9170);
nor U9635 (N_9635,N_9121,N_9268);
nand U9636 (N_9636,N_9572,N_9503);
or U9637 (N_9637,N_9139,N_9344);
nor U9638 (N_9638,N_9000,N_9545);
nand U9639 (N_9639,N_9397,N_9490);
nor U9640 (N_9640,N_9130,N_9367);
xor U9641 (N_9641,N_9115,N_9028);
xnor U9642 (N_9642,N_9183,N_9596);
nor U9643 (N_9643,N_9035,N_9073);
nand U9644 (N_9644,N_9440,N_9421);
nor U9645 (N_9645,N_9052,N_9096);
or U9646 (N_9646,N_9314,N_9235);
xnor U9647 (N_9647,N_9571,N_9327);
nand U9648 (N_9648,N_9319,N_9510);
xor U9649 (N_9649,N_9295,N_9013);
nand U9650 (N_9650,N_9439,N_9104);
or U9651 (N_9651,N_9316,N_9410);
and U9652 (N_9652,N_9495,N_9456);
xnor U9653 (N_9653,N_9529,N_9582);
and U9654 (N_9654,N_9533,N_9059);
or U9655 (N_9655,N_9526,N_9559);
nor U9656 (N_9656,N_9105,N_9349);
nand U9657 (N_9657,N_9366,N_9486);
and U9658 (N_9658,N_9348,N_9262);
nor U9659 (N_9659,N_9473,N_9247);
nand U9660 (N_9660,N_9408,N_9031);
xnor U9661 (N_9661,N_9378,N_9094);
nor U9662 (N_9662,N_9551,N_9335);
nand U9663 (N_9663,N_9097,N_9212);
xor U9664 (N_9664,N_9099,N_9467);
nand U9665 (N_9665,N_9149,N_9432);
xnor U9666 (N_9666,N_9532,N_9275);
nand U9667 (N_9667,N_9350,N_9014);
or U9668 (N_9668,N_9032,N_9218);
nor U9669 (N_9669,N_9515,N_9573);
or U9670 (N_9670,N_9591,N_9304);
and U9671 (N_9671,N_9435,N_9554);
or U9672 (N_9672,N_9012,N_9113);
or U9673 (N_9673,N_9407,N_9140);
and U9674 (N_9674,N_9285,N_9217);
nand U9675 (N_9675,N_9557,N_9565);
nand U9676 (N_9676,N_9084,N_9172);
or U9677 (N_9677,N_9322,N_9036);
xnor U9678 (N_9678,N_9588,N_9147);
or U9679 (N_9679,N_9225,N_9100);
or U9680 (N_9680,N_9011,N_9382);
nand U9681 (N_9681,N_9334,N_9254);
and U9682 (N_9682,N_9021,N_9354);
nor U9683 (N_9683,N_9249,N_9284);
and U9684 (N_9684,N_9064,N_9449);
and U9685 (N_9685,N_9162,N_9019);
or U9686 (N_9686,N_9491,N_9240);
nor U9687 (N_9687,N_9143,N_9219);
and U9688 (N_9688,N_9328,N_9200);
or U9689 (N_9689,N_9244,N_9209);
xor U9690 (N_9690,N_9347,N_9107);
nand U9691 (N_9691,N_9164,N_9241);
nor U9692 (N_9692,N_9524,N_9252);
nor U9693 (N_9693,N_9310,N_9306);
xor U9694 (N_9694,N_9087,N_9137);
xor U9695 (N_9695,N_9505,N_9233);
xnor U9696 (N_9696,N_9261,N_9160);
nand U9697 (N_9697,N_9267,N_9208);
nor U9698 (N_9698,N_9058,N_9531);
and U9699 (N_9699,N_9430,N_9075);
xor U9700 (N_9700,N_9043,N_9114);
nor U9701 (N_9701,N_9446,N_9188);
or U9702 (N_9702,N_9040,N_9485);
and U9703 (N_9703,N_9050,N_9145);
nor U9704 (N_9704,N_9383,N_9458);
or U9705 (N_9705,N_9251,N_9385);
and U9706 (N_9706,N_9083,N_9069);
or U9707 (N_9707,N_9323,N_9238);
or U9708 (N_9708,N_9193,N_9198);
and U9709 (N_9709,N_9124,N_9102);
nand U9710 (N_9710,N_9008,N_9568);
xor U9711 (N_9711,N_9215,N_9269);
nor U9712 (N_9712,N_9226,N_9376);
nor U9713 (N_9713,N_9530,N_9108);
or U9714 (N_9714,N_9369,N_9561);
and U9715 (N_9715,N_9082,N_9179);
nor U9716 (N_9716,N_9589,N_9002);
nor U9717 (N_9717,N_9060,N_9372);
and U9718 (N_9718,N_9228,N_9199);
nor U9719 (N_9719,N_9182,N_9534);
nand U9720 (N_9720,N_9091,N_9175);
xor U9721 (N_9721,N_9417,N_9462);
nand U9722 (N_9722,N_9161,N_9007);
nor U9723 (N_9723,N_9273,N_9393);
and U9724 (N_9724,N_9441,N_9363);
and U9725 (N_9725,N_9569,N_9041);
xnor U9726 (N_9726,N_9299,N_9203);
xor U9727 (N_9727,N_9025,N_9313);
nand U9728 (N_9728,N_9519,N_9255);
xor U9729 (N_9729,N_9263,N_9436);
nor U9730 (N_9730,N_9142,N_9427);
xnor U9731 (N_9731,N_9029,N_9566);
nand U9732 (N_9732,N_9174,N_9506);
xnor U9733 (N_9733,N_9429,N_9570);
and U9734 (N_9734,N_9477,N_9468);
nand U9735 (N_9735,N_9312,N_9101);
nand U9736 (N_9736,N_9460,N_9250);
xnor U9737 (N_9737,N_9197,N_9184);
nor U9738 (N_9738,N_9543,N_9339);
nor U9739 (N_9739,N_9006,N_9289);
nor U9740 (N_9740,N_9438,N_9521);
or U9741 (N_9741,N_9583,N_9067);
xnor U9742 (N_9742,N_9317,N_9151);
nor U9743 (N_9743,N_9388,N_9333);
or U9744 (N_9744,N_9489,N_9281);
and U9745 (N_9745,N_9592,N_9051);
or U9746 (N_9746,N_9454,N_9258);
or U9747 (N_9747,N_9359,N_9504);
nand U9748 (N_9748,N_9552,N_9210);
nand U9749 (N_9749,N_9528,N_9079);
nor U9750 (N_9750,N_9345,N_9448);
xnor U9751 (N_9751,N_9077,N_9057);
xor U9752 (N_9752,N_9221,N_9033);
xnor U9753 (N_9753,N_9411,N_9336);
nand U9754 (N_9754,N_9178,N_9443);
xor U9755 (N_9755,N_9214,N_9211);
xor U9756 (N_9756,N_9466,N_9472);
xnor U9757 (N_9757,N_9593,N_9116);
nor U9758 (N_9758,N_9265,N_9132);
xnor U9759 (N_9759,N_9315,N_9562);
nand U9760 (N_9760,N_9416,N_9401);
and U9761 (N_9761,N_9527,N_9459);
nand U9762 (N_9762,N_9597,N_9483);
nor U9763 (N_9763,N_9474,N_9260);
and U9764 (N_9764,N_9027,N_9498);
nor U9765 (N_9765,N_9098,N_9293);
xnor U9766 (N_9766,N_9213,N_9457);
and U9767 (N_9767,N_9296,N_9015);
and U9768 (N_9768,N_9078,N_9291);
nand U9769 (N_9769,N_9577,N_9154);
and U9770 (N_9770,N_9404,N_9119);
or U9771 (N_9771,N_9090,N_9227);
or U9772 (N_9772,N_9173,N_9358);
or U9773 (N_9773,N_9246,N_9346);
nor U9774 (N_9774,N_9297,N_9039);
xnor U9775 (N_9775,N_9062,N_9123);
or U9776 (N_9776,N_9351,N_9392);
nor U9777 (N_9777,N_9074,N_9018);
or U9778 (N_9778,N_9379,N_9305);
nor U9779 (N_9779,N_9243,N_9395);
or U9780 (N_9780,N_9017,N_9576);
nor U9781 (N_9781,N_9331,N_9470);
or U9782 (N_9782,N_9434,N_9171);
or U9783 (N_9783,N_9229,N_9095);
or U9784 (N_9784,N_9371,N_9181);
xnor U9785 (N_9785,N_9356,N_9259);
xnor U9786 (N_9786,N_9512,N_9085);
nand U9787 (N_9787,N_9423,N_9482);
nand U9788 (N_9788,N_9386,N_9177);
xnor U9789 (N_9789,N_9387,N_9176);
or U9790 (N_9790,N_9152,N_9186);
nor U9791 (N_9791,N_9070,N_9341);
xnor U9792 (N_9792,N_9413,N_9180);
nand U9793 (N_9793,N_9318,N_9053);
or U9794 (N_9794,N_9080,N_9167);
and U9795 (N_9795,N_9484,N_9567);
xor U9796 (N_9796,N_9009,N_9578);
and U9797 (N_9797,N_9072,N_9564);
xnor U9798 (N_9798,N_9442,N_9437);
or U9799 (N_9799,N_9403,N_9539);
or U9800 (N_9800,N_9308,N_9419);
or U9801 (N_9801,N_9103,N_9425);
and U9802 (N_9802,N_9450,N_9465);
nor U9803 (N_9803,N_9294,N_9508);
and U9804 (N_9804,N_9239,N_9481);
nand U9805 (N_9805,N_9594,N_9518);
nand U9806 (N_9806,N_9093,N_9377);
or U9807 (N_9807,N_9185,N_9163);
xor U9808 (N_9808,N_9237,N_9402);
nand U9809 (N_9809,N_9242,N_9047);
nand U9810 (N_9810,N_9223,N_9081);
or U9811 (N_9811,N_9201,N_9560);
xor U9812 (N_9812,N_9128,N_9464);
xnor U9813 (N_9813,N_9493,N_9042);
and U9814 (N_9814,N_9355,N_9360);
or U9815 (N_9815,N_9065,N_9480);
xor U9816 (N_9816,N_9122,N_9579);
nand U9817 (N_9817,N_9517,N_9340);
and U9818 (N_9818,N_9342,N_9234);
nand U9819 (N_9819,N_9150,N_9157);
or U9820 (N_9820,N_9544,N_9469);
nand U9821 (N_9821,N_9245,N_9502);
xor U9822 (N_9822,N_9368,N_9061);
nor U9823 (N_9823,N_9045,N_9478);
nor U9824 (N_9824,N_9492,N_9542);
and U9825 (N_9825,N_9230,N_9324);
nor U9826 (N_9826,N_9054,N_9415);
and U9827 (N_9827,N_9153,N_9155);
and U9828 (N_9828,N_9046,N_9278);
or U9829 (N_9829,N_9399,N_9026);
nor U9830 (N_9830,N_9086,N_9169);
or U9831 (N_9831,N_9134,N_9274);
xnor U9832 (N_9832,N_9487,N_9409);
and U9833 (N_9833,N_9390,N_9364);
xor U9834 (N_9834,N_9166,N_9520);
nand U9835 (N_9835,N_9126,N_9190);
nor U9836 (N_9836,N_9037,N_9538);
xor U9837 (N_9837,N_9156,N_9136);
or U9838 (N_9838,N_9374,N_9148);
and U9839 (N_9839,N_9194,N_9509);
and U9840 (N_9840,N_9447,N_9373);
and U9841 (N_9841,N_9353,N_9248);
nand U9842 (N_9842,N_9224,N_9352);
xnor U9843 (N_9843,N_9277,N_9112);
and U9844 (N_9844,N_9329,N_9475);
nor U9845 (N_9845,N_9586,N_9236);
xnor U9846 (N_9846,N_9129,N_9575);
nand U9847 (N_9847,N_9159,N_9206);
nand U9848 (N_9848,N_9071,N_9191);
nand U9849 (N_9849,N_9118,N_9433);
nand U9850 (N_9850,N_9204,N_9452);
or U9851 (N_9851,N_9038,N_9550);
nand U9852 (N_9852,N_9205,N_9282);
nor U9853 (N_9853,N_9444,N_9496);
and U9854 (N_9854,N_9590,N_9535);
xnor U9855 (N_9855,N_9494,N_9189);
nor U9856 (N_9856,N_9320,N_9216);
xnor U9857 (N_9857,N_9451,N_9406);
nor U9858 (N_9858,N_9135,N_9453);
nor U9859 (N_9859,N_9362,N_9553);
nor U9860 (N_9860,N_9595,N_9580);
or U9861 (N_9861,N_9141,N_9110);
xor U9862 (N_9862,N_9287,N_9003);
and U9863 (N_9863,N_9394,N_9168);
nor U9864 (N_9864,N_9120,N_9497);
nand U9865 (N_9865,N_9111,N_9030);
and U9866 (N_9866,N_9516,N_9461);
nand U9867 (N_9867,N_9133,N_9187);
or U9868 (N_9868,N_9422,N_9092);
xnor U9869 (N_9869,N_9405,N_9375);
xor U9870 (N_9870,N_9195,N_9585);
nor U9871 (N_9871,N_9001,N_9088);
and U9872 (N_9872,N_9279,N_9424);
or U9873 (N_9873,N_9384,N_9547);
nand U9874 (N_9874,N_9431,N_9004);
nor U9875 (N_9875,N_9256,N_9192);
xnor U9876 (N_9876,N_9412,N_9303);
nand U9877 (N_9877,N_9302,N_9549);
nor U9878 (N_9878,N_9264,N_9055);
or U9879 (N_9879,N_9381,N_9584);
xnor U9880 (N_9880,N_9556,N_9301);
xnor U9881 (N_9881,N_9048,N_9598);
xor U9882 (N_9882,N_9127,N_9125);
or U9883 (N_9883,N_9068,N_9266);
nor U9884 (N_9884,N_9300,N_9016);
xor U9885 (N_9885,N_9574,N_9398);
nand U9886 (N_9886,N_9222,N_9479);
and U9887 (N_9887,N_9089,N_9220);
nor U9888 (N_9888,N_9117,N_9307);
and U9889 (N_9889,N_9283,N_9525);
xnor U9890 (N_9890,N_9321,N_9500);
or U9891 (N_9891,N_9010,N_9476);
nor U9892 (N_9892,N_9455,N_9023);
xnor U9893 (N_9893,N_9049,N_9428);
or U9894 (N_9894,N_9400,N_9066);
nor U9895 (N_9895,N_9445,N_9158);
nand U9896 (N_9896,N_9231,N_9581);
or U9897 (N_9897,N_9280,N_9286);
or U9898 (N_9898,N_9292,N_9587);
and U9899 (N_9899,N_9507,N_9288);
nand U9900 (N_9900,N_9523,N_9422);
nand U9901 (N_9901,N_9053,N_9057);
or U9902 (N_9902,N_9062,N_9178);
and U9903 (N_9903,N_9234,N_9291);
nand U9904 (N_9904,N_9369,N_9298);
xor U9905 (N_9905,N_9486,N_9062);
nand U9906 (N_9906,N_9019,N_9390);
xor U9907 (N_9907,N_9330,N_9277);
nand U9908 (N_9908,N_9219,N_9120);
or U9909 (N_9909,N_9249,N_9044);
nand U9910 (N_9910,N_9372,N_9023);
nand U9911 (N_9911,N_9294,N_9250);
nor U9912 (N_9912,N_9085,N_9303);
nor U9913 (N_9913,N_9440,N_9054);
xor U9914 (N_9914,N_9299,N_9499);
nand U9915 (N_9915,N_9471,N_9469);
nand U9916 (N_9916,N_9437,N_9114);
nor U9917 (N_9917,N_9096,N_9583);
xnor U9918 (N_9918,N_9398,N_9353);
and U9919 (N_9919,N_9590,N_9207);
xor U9920 (N_9920,N_9039,N_9384);
nand U9921 (N_9921,N_9471,N_9474);
nor U9922 (N_9922,N_9504,N_9448);
and U9923 (N_9923,N_9032,N_9120);
nor U9924 (N_9924,N_9372,N_9343);
nor U9925 (N_9925,N_9449,N_9415);
xnor U9926 (N_9926,N_9480,N_9418);
and U9927 (N_9927,N_9123,N_9265);
nand U9928 (N_9928,N_9584,N_9339);
xnor U9929 (N_9929,N_9452,N_9064);
nor U9930 (N_9930,N_9380,N_9377);
xnor U9931 (N_9931,N_9449,N_9424);
nand U9932 (N_9932,N_9303,N_9160);
and U9933 (N_9933,N_9536,N_9154);
xor U9934 (N_9934,N_9513,N_9251);
or U9935 (N_9935,N_9453,N_9391);
and U9936 (N_9936,N_9366,N_9438);
xor U9937 (N_9937,N_9008,N_9535);
nand U9938 (N_9938,N_9206,N_9142);
and U9939 (N_9939,N_9092,N_9220);
nor U9940 (N_9940,N_9108,N_9437);
xnor U9941 (N_9941,N_9148,N_9294);
or U9942 (N_9942,N_9114,N_9536);
nor U9943 (N_9943,N_9431,N_9533);
nor U9944 (N_9944,N_9060,N_9220);
xor U9945 (N_9945,N_9361,N_9124);
xnor U9946 (N_9946,N_9063,N_9425);
nand U9947 (N_9947,N_9192,N_9357);
nor U9948 (N_9948,N_9189,N_9599);
nand U9949 (N_9949,N_9401,N_9146);
and U9950 (N_9950,N_9126,N_9463);
nand U9951 (N_9951,N_9371,N_9155);
nand U9952 (N_9952,N_9446,N_9245);
xnor U9953 (N_9953,N_9134,N_9484);
and U9954 (N_9954,N_9030,N_9523);
nor U9955 (N_9955,N_9359,N_9116);
nor U9956 (N_9956,N_9277,N_9430);
or U9957 (N_9957,N_9529,N_9301);
nor U9958 (N_9958,N_9017,N_9127);
nand U9959 (N_9959,N_9165,N_9153);
nand U9960 (N_9960,N_9049,N_9493);
xnor U9961 (N_9961,N_9571,N_9013);
or U9962 (N_9962,N_9271,N_9411);
or U9963 (N_9963,N_9333,N_9592);
xnor U9964 (N_9964,N_9195,N_9086);
or U9965 (N_9965,N_9434,N_9329);
xnor U9966 (N_9966,N_9376,N_9036);
nor U9967 (N_9967,N_9426,N_9160);
nand U9968 (N_9968,N_9344,N_9076);
and U9969 (N_9969,N_9527,N_9200);
and U9970 (N_9970,N_9036,N_9070);
and U9971 (N_9971,N_9442,N_9452);
xor U9972 (N_9972,N_9163,N_9062);
or U9973 (N_9973,N_9399,N_9438);
nand U9974 (N_9974,N_9226,N_9037);
xnor U9975 (N_9975,N_9517,N_9547);
or U9976 (N_9976,N_9241,N_9442);
and U9977 (N_9977,N_9072,N_9399);
nand U9978 (N_9978,N_9018,N_9145);
or U9979 (N_9979,N_9027,N_9279);
nand U9980 (N_9980,N_9220,N_9059);
and U9981 (N_9981,N_9446,N_9047);
nor U9982 (N_9982,N_9350,N_9194);
nor U9983 (N_9983,N_9517,N_9001);
nand U9984 (N_9984,N_9198,N_9523);
nand U9985 (N_9985,N_9014,N_9391);
or U9986 (N_9986,N_9500,N_9113);
nor U9987 (N_9987,N_9006,N_9287);
xnor U9988 (N_9988,N_9587,N_9165);
and U9989 (N_9989,N_9381,N_9391);
nand U9990 (N_9990,N_9122,N_9511);
or U9991 (N_9991,N_9586,N_9057);
and U9992 (N_9992,N_9207,N_9187);
xnor U9993 (N_9993,N_9244,N_9518);
xnor U9994 (N_9994,N_9041,N_9511);
and U9995 (N_9995,N_9331,N_9111);
xnor U9996 (N_9996,N_9099,N_9415);
and U9997 (N_9997,N_9391,N_9465);
nor U9998 (N_9998,N_9121,N_9122);
and U9999 (N_9999,N_9211,N_9234);
xnor U10000 (N_10000,N_9437,N_9434);
nor U10001 (N_10001,N_9438,N_9147);
nor U10002 (N_10002,N_9345,N_9027);
or U10003 (N_10003,N_9109,N_9181);
or U10004 (N_10004,N_9549,N_9559);
nor U10005 (N_10005,N_9288,N_9089);
xor U10006 (N_10006,N_9044,N_9234);
nor U10007 (N_10007,N_9482,N_9046);
nor U10008 (N_10008,N_9453,N_9002);
and U10009 (N_10009,N_9592,N_9202);
xnor U10010 (N_10010,N_9525,N_9256);
xnor U10011 (N_10011,N_9153,N_9186);
nor U10012 (N_10012,N_9481,N_9385);
nor U10013 (N_10013,N_9478,N_9205);
and U10014 (N_10014,N_9083,N_9461);
or U10015 (N_10015,N_9374,N_9426);
xnor U10016 (N_10016,N_9441,N_9405);
xnor U10017 (N_10017,N_9432,N_9435);
nor U10018 (N_10018,N_9461,N_9310);
or U10019 (N_10019,N_9439,N_9249);
nand U10020 (N_10020,N_9509,N_9116);
and U10021 (N_10021,N_9018,N_9517);
nand U10022 (N_10022,N_9289,N_9552);
and U10023 (N_10023,N_9529,N_9230);
and U10024 (N_10024,N_9218,N_9042);
or U10025 (N_10025,N_9447,N_9254);
nand U10026 (N_10026,N_9152,N_9269);
nor U10027 (N_10027,N_9212,N_9262);
xor U10028 (N_10028,N_9290,N_9039);
nor U10029 (N_10029,N_9134,N_9182);
xnor U10030 (N_10030,N_9510,N_9307);
xor U10031 (N_10031,N_9408,N_9517);
and U10032 (N_10032,N_9163,N_9259);
nor U10033 (N_10033,N_9574,N_9284);
xnor U10034 (N_10034,N_9343,N_9593);
and U10035 (N_10035,N_9111,N_9492);
nor U10036 (N_10036,N_9545,N_9172);
xnor U10037 (N_10037,N_9236,N_9095);
or U10038 (N_10038,N_9475,N_9594);
and U10039 (N_10039,N_9168,N_9553);
xnor U10040 (N_10040,N_9580,N_9318);
nor U10041 (N_10041,N_9198,N_9389);
nor U10042 (N_10042,N_9082,N_9509);
xnor U10043 (N_10043,N_9019,N_9067);
nor U10044 (N_10044,N_9327,N_9012);
xor U10045 (N_10045,N_9107,N_9054);
nand U10046 (N_10046,N_9075,N_9373);
and U10047 (N_10047,N_9071,N_9061);
xor U10048 (N_10048,N_9309,N_9532);
or U10049 (N_10049,N_9300,N_9289);
xnor U10050 (N_10050,N_9136,N_9442);
and U10051 (N_10051,N_9563,N_9505);
and U10052 (N_10052,N_9127,N_9174);
nor U10053 (N_10053,N_9234,N_9391);
xor U10054 (N_10054,N_9470,N_9153);
nand U10055 (N_10055,N_9194,N_9084);
xor U10056 (N_10056,N_9035,N_9283);
or U10057 (N_10057,N_9326,N_9194);
xnor U10058 (N_10058,N_9213,N_9210);
nor U10059 (N_10059,N_9293,N_9560);
and U10060 (N_10060,N_9261,N_9213);
nor U10061 (N_10061,N_9479,N_9048);
nand U10062 (N_10062,N_9093,N_9115);
or U10063 (N_10063,N_9553,N_9269);
and U10064 (N_10064,N_9094,N_9374);
xnor U10065 (N_10065,N_9515,N_9510);
nand U10066 (N_10066,N_9277,N_9015);
nand U10067 (N_10067,N_9570,N_9074);
nor U10068 (N_10068,N_9203,N_9514);
nor U10069 (N_10069,N_9266,N_9205);
nor U10070 (N_10070,N_9099,N_9566);
xor U10071 (N_10071,N_9195,N_9005);
nor U10072 (N_10072,N_9517,N_9360);
nor U10073 (N_10073,N_9306,N_9579);
or U10074 (N_10074,N_9433,N_9342);
nand U10075 (N_10075,N_9533,N_9033);
nor U10076 (N_10076,N_9093,N_9185);
or U10077 (N_10077,N_9437,N_9372);
and U10078 (N_10078,N_9495,N_9598);
xnor U10079 (N_10079,N_9574,N_9467);
and U10080 (N_10080,N_9400,N_9487);
xnor U10081 (N_10081,N_9105,N_9411);
xor U10082 (N_10082,N_9155,N_9559);
nor U10083 (N_10083,N_9026,N_9502);
and U10084 (N_10084,N_9440,N_9324);
or U10085 (N_10085,N_9236,N_9185);
nand U10086 (N_10086,N_9564,N_9293);
nor U10087 (N_10087,N_9583,N_9445);
nor U10088 (N_10088,N_9234,N_9217);
or U10089 (N_10089,N_9062,N_9128);
nand U10090 (N_10090,N_9400,N_9172);
or U10091 (N_10091,N_9389,N_9571);
or U10092 (N_10092,N_9061,N_9002);
or U10093 (N_10093,N_9347,N_9542);
xor U10094 (N_10094,N_9264,N_9312);
or U10095 (N_10095,N_9232,N_9277);
nor U10096 (N_10096,N_9238,N_9372);
nor U10097 (N_10097,N_9180,N_9201);
and U10098 (N_10098,N_9133,N_9399);
or U10099 (N_10099,N_9083,N_9381);
nor U10100 (N_10100,N_9219,N_9401);
xnor U10101 (N_10101,N_9551,N_9254);
xnor U10102 (N_10102,N_9297,N_9198);
and U10103 (N_10103,N_9557,N_9141);
xnor U10104 (N_10104,N_9151,N_9472);
nor U10105 (N_10105,N_9279,N_9453);
xor U10106 (N_10106,N_9223,N_9029);
xnor U10107 (N_10107,N_9215,N_9478);
nor U10108 (N_10108,N_9498,N_9439);
xor U10109 (N_10109,N_9413,N_9358);
nor U10110 (N_10110,N_9437,N_9452);
nor U10111 (N_10111,N_9067,N_9057);
xor U10112 (N_10112,N_9002,N_9149);
and U10113 (N_10113,N_9546,N_9016);
xor U10114 (N_10114,N_9132,N_9164);
xnor U10115 (N_10115,N_9255,N_9304);
and U10116 (N_10116,N_9305,N_9119);
and U10117 (N_10117,N_9439,N_9140);
nor U10118 (N_10118,N_9368,N_9350);
or U10119 (N_10119,N_9082,N_9348);
xor U10120 (N_10120,N_9584,N_9061);
nand U10121 (N_10121,N_9495,N_9205);
nand U10122 (N_10122,N_9351,N_9192);
nand U10123 (N_10123,N_9159,N_9591);
and U10124 (N_10124,N_9164,N_9415);
nand U10125 (N_10125,N_9056,N_9341);
or U10126 (N_10126,N_9057,N_9437);
nor U10127 (N_10127,N_9374,N_9361);
and U10128 (N_10128,N_9081,N_9405);
and U10129 (N_10129,N_9181,N_9575);
nor U10130 (N_10130,N_9592,N_9392);
and U10131 (N_10131,N_9517,N_9060);
or U10132 (N_10132,N_9268,N_9133);
and U10133 (N_10133,N_9334,N_9058);
xnor U10134 (N_10134,N_9486,N_9042);
xnor U10135 (N_10135,N_9242,N_9542);
nand U10136 (N_10136,N_9191,N_9366);
or U10137 (N_10137,N_9142,N_9384);
nor U10138 (N_10138,N_9194,N_9046);
nor U10139 (N_10139,N_9573,N_9285);
xor U10140 (N_10140,N_9228,N_9361);
nor U10141 (N_10141,N_9503,N_9148);
xor U10142 (N_10142,N_9582,N_9577);
nand U10143 (N_10143,N_9513,N_9473);
nand U10144 (N_10144,N_9241,N_9251);
or U10145 (N_10145,N_9143,N_9064);
or U10146 (N_10146,N_9434,N_9380);
xnor U10147 (N_10147,N_9253,N_9226);
or U10148 (N_10148,N_9366,N_9004);
or U10149 (N_10149,N_9173,N_9050);
xor U10150 (N_10150,N_9169,N_9031);
nand U10151 (N_10151,N_9343,N_9578);
or U10152 (N_10152,N_9053,N_9121);
and U10153 (N_10153,N_9561,N_9495);
nor U10154 (N_10154,N_9009,N_9325);
and U10155 (N_10155,N_9094,N_9182);
or U10156 (N_10156,N_9573,N_9047);
or U10157 (N_10157,N_9378,N_9079);
or U10158 (N_10158,N_9355,N_9321);
xor U10159 (N_10159,N_9340,N_9344);
or U10160 (N_10160,N_9557,N_9352);
or U10161 (N_10161,N_9080,N_9234);
xor U10162 (N_10162,N_9215,N_9381);
and U10163 (N_10163,N_9529,N_9463);
or U10164 (N_10164,N_9248,N_9295);
nor U10165 (N_10165,N_9410,N_9034);
nand U10166 (N_10166,N_9430,N_9312);
or U10167 (N_10167,N_9290,N_9338);
and U10168 (N_10168,N_9449,N_9167);
or U10169 (N_10169,N_9036,N_9502);
and U10170 (N_10170,N_9568,N_9291);
nor U10171 (N_10171,N_9551,N_9574);
xnor U10172 (N_10172,N_9470,N_9571);
and U10173 (N_10173,N_9174,N_9293);
nor U10174 (N_10174,N_9154,N_9503);
nand U10175 (N_10175,N_9226,N_9173);
nor U10176 (N_10176,N_9378,N_9397);
or U10177 (N_10177,N_9362,N_9058);
xnor U10178 (N_10178,N_9416,N_9034);
nor U10179 (N_10179,N_9065,N_9013);
and U10180 (N_10180,N_9483,N_9027);
xnor U10181 (N_10181,N_9210,N_9435);
or U10182 (N_10182,N_9054,N_9434);
and U10183 (N_10183,N_9182,N_9081);
nor U10184 (N_10184,N_9480,N_9024);
and U10185 (N_10185,N_9379,N_9081);
and U10186 (N_10186,N_9025,N_9042);
nor U10187 (N_10187,N_9507,N_9137);
nand U10188 (N_10188,N_9150,N_9102);
xnor U10189 (N_10189,N_9368,N_9565);
xnor U10190 (N_10190,N_9152,N_9572);
nand U10191 (N_10191,N_9220,N_9140);
xnor U10192 (N_10192,N_9425,N_9130);
xnor U10193 (N_10193,N_9383,N_9389);
nor U10194 (N_10194,N_9066,N_9471);
nor U10195 (N_10195,N_9021,N_9476);
nor U10196 (N_10196,N_9225,N_9485);
nor U10197 (N_10197,N_9061,N_9370);
xnor U10198 (N_10198,N_9594,N_9490);
and U10199 (N_10199,N_9376,N_9000);
nand U10200 (N_10200,N_9795,N_9952);
or U10201 (N_10201,N_9891,N_10062);
or U10202 (N_10202,N_9782,N_9611);
nand U10203 (N_10203,N_10188,N_9883);
nand U10204 (N_10204,N_9990,N_10146);
nor U10205 (N_10205,N_10114,N_9756);
and U10206 (N_10206,N_10177,N_9815);
and U10207 (N_10207,N_10125,N_9750);
nand U10208 (N_10208,N_9961,N_9651);
nor U10209 (N_10209,N_9881,N_9767);
and U10210 (N_10210,N_9775,N_9863);
nor U10211 (N_10211,N_10159,N_10142);
and U10212 (N_10212,N_9793,N_9777);
nand U10213 (N_10213,N_9758,N_9989);
nand U10214 (N_10214,N_9853,N_9824);
or U10215 (N_10215,N_10123,N_9983);
and U10216 (N_10216,N_10175,N_9980);
and U10217 (N_10217,N_9702,N_10106);
xnor U10218 (N_10218,N_10046,N_9601);
or U10219 (N_10219,N_10100,N_9647);
nand U10220 (N_10220,N_10086,N_9972);
nand U10221 (N_10221,N_9716,N_9920);
and U10222 (N_10222,N_10149,N_9654);
xnor U10223 (N_10223,N_9762,N_9948);
nand U10224 (N_10224,N_9909,N_9728);
nand U10225 (N_10225,N_9783,N_9910);
and U10226 (N_10226,N_9691,N_9818);
and U10227 (N_10227,N_9944,N_9878);
and U10228 (N_10228,N_9698,N_10119);
or U10229 (N_10229,N_9773,N_9638);
or U10230 (N_10230,N_9760,N_10191);
nor U10231 (N_10231,N_9641,N_9988);
nor U10232 (N_10232,N_9688,N_10048);
nor U10233 (N_10233,N_9656,N_9757);
and U10234 (N_10234,N_9998,N_9974);
xor U10235 (N_10235,N_10002,N_9821);
or U10236 (N_10236,N_9840,N_9721);
and U10237 (N_10237,N_9867,N_10044);
and U10238 (N_10238,N_10129,N_9659);
or U10239 (N_10239,N_9904,N_9907);
xnor U10240 (N_10240,N_9649,N_9704);
nand U10241 (N_10241,N_9623,N_9754);
or U10242 (N_10242,N_9785,N_9849);
and U10243 (N_10243,N_9732,N_9660);
xnor U10244 (N_10244,N_9938,N_9928);
or U10245 (N_10245,N_9960,N_9671);
and U10246 (N_10246,N_10045,N_9986);
nand U10247 (N_10247,N_9994,N_9788);
nand U10248 (N_10248,N_9666,N_10032);
or U10249 (N_10249,N_10053,N_9642);
and U10250 (N_10250,N_9876,N_9893);
and U10251 (N_10251,N_9792,N_9820);
or U10252 (N_10252,N_10172,N_9977);
nor U10253 (N_10253,N_9620,N_9720);
and U10254 (N_10254,N_10051,N_10012);
nor U10255 (N_10255,N_9799,N_10094);
xnor U10256 (N_10256,N_10179,N_9913);
or U10257 (N_10257,N_9607,N_10133);
nor U10258 (N_10258,N_10000,N_9838);
or U10259 (N_10259,N_9852,N_10026);
or U10260 (N_10260,N_9796,N_9610);
and U10261 (N_10261,N_9812,N_9939);
nand U10262 (N_10262,N_9662,N_10145);
and U10263 (N_10263,N_10084,N_9618);
xnor U10264 (N_10264,N_10090,N_9632);
nor U10265 (N_10265,N_9900,N_9930);
or U10266 (N_10266,N_9786,N_9709);
nand U10267 (N_10267,N_10047,N_9832);
nor U10268 (N_10268,N_9860,N_9755);
nor U10269 (N_10269,N_9609,N_9707);
and U10270 (N_10270,N_10015,N_10108);
xnor U10271 (N_10271,N_9926,N_10006);
nor U10272 (N_10272,N_10088,N_9615);
and U10273 (N_10273,N_10120,N_9740);
and U10274 (N_10274,N_9810,N_9946);
xor U10275 (N_10275,N_9997,N_10140);
nor U10276 (N_10276,N_9700,N_9637);
nand U10277 (N_10277,N_9759,N_9970);
or U10278 (N_10278,N_9646,N_10096);
nand U10279 (N_10279,N_9809,N_10166);
xnor U10280 (N_10280,N_10139,N_10054);
xor U10281 (N_10281,N_9669,N_9639);
nand U10282 (N_10282,N_9922,N_10071);
or U10283 (N_10283,N_9828,N_9882);
and U10284 (N_10284,N_10132,N_9635);
and U10285 (N_10285,N_10173,N_9789);
or U10286 (N_10286,N_9914,N_9872);
and U10287 (N_10287,N_9667,N_10031);
xor U10288 (N_10288,N_10025,N_9801);
nand U10289 (N_10289,N_10131,N_10092);
and U10290 (N_10290,N_9836,N_9866);
nor U10291 (N_10291,N_10034,N_10095);
nand U10292 (N_10292,N_10136,N_9606);
nor U10293 (N_10293,N_10137,N_9778);
and U10294 (N_10294,N_9825,N_9644);
or U10295 (N_10295,N_10013,N_10043);
nor U10296 (N_10296,N_10164,N_10082);
and U10297 (N_10297,N_10112,N_9627);
nor U10298 (N_10298,N_9906,N_10028);
nor U10299 (N_10299,N_10102,N_10056);
and U10300 (N_10300,N_9945,N_10041);
nor U10301 (N_10301,N_9678,N_9886);
nand U10302 (N_10302,N_9874,N_10030);
or U10303 (N_10303,N_9991,N_9676);
xor U10304 (N_10304,N_10004,N_10192);
nor U10305 (N_10305,N_10184,N_9854);
and U10306 (N_10306,N_9631,N_10049);
nand U10307 (N_10307,N_10079,N_10040);
nor U10308 (N_10308,N_9898,N_10196);
nand U10309 (N_10309,N_9803,N_10117);
nor U10310 (N_10310,N_10021,N_10099);
xor U10311 (N_10311,N_9680,N_10087);
and U10312 (N_10312,N_10148,N_9625);
or U10313 (N_10313,N_10039,N_9889);
nand U10314 (N_10314,N_10147,N_10181);
nor U10315 (N_10315,N_9665,N_9743);
nand U10316 (N_10316,N_9770,N_9830);
and U10317 (N_10317,N_10174,N_9748);
and U10318 (N_10318,N_10063,N_9684);
nand U10319 (N_10319,N_9817,N_9925);
or U10320 (N_10320,N_10070,N_9912);
nor U10321 (N_10321,N_9902,N_9957);
or U10322 (N_10322,N_10135,N_9738);
nand U10323 (N_10323,N_10073,N_10198);
xor U10324 (N_10324,N_10016,N_9622);
xnor U10325 (N_10325,N_9776,N_9981);
nand U10326 (N_10326,N_9718,N_10093);
xnor U10327 (N_10327,N_10029,N_9640);
xnor U10328 (N_10328,N_9741,N_9712);
nand U10329 (N_10329,N_10190,N_9927);
xor U10330 (N_10330,N_10182,N_9822);
or U10331 (N_10331,N_10023,N_10115);
nand U10332 (N_10332,N_10162,N_9703);
xor U10333 (N_10333,N_9630,N_9616);
or U10334 (N_10334,N_9650,N_9950);
or U10335 (N_10335,N_10124,N_9917);
xnor U10336 (N_10336,N_10078,N_10017);
xnor U10337 (N_10337,N_9865,N_9655);
xnor U10338 (N_10338,N_9781,N_9947);
nand U10339 (N_10339,N_9870,N_9608);
or U10340 (N_10340,N_9805,N_10022);
and U10341 (N_10341,N_10060,N_9965);
xnor U10342 (N_10342,N_10199,N_9962);
nor U10343 (N_10343,N_9600,N_10169);
nor U10344 (N_10344,N_9919,N_9784);
nor U10345 (N_10345,N_10141,N_9675);
nor U10346 (N_10346,N_9621,N_9847);
and U10347 (N_10347,N_9887,N_10130);
nor U10348 (N_10348,N_9713,N_9976);
nand U10349 (N_10349,N_9674,N_10197);
nor U10350 (N_10350,N_10144,N_10186);
xnor U10351 (N_10351,N_9835,N_10008);
nor U10352 (N_10352,N_10121,N_9686);
nor U10353 (N_10353,N_10165,N_9672);
and U10354 (N_10354,N_10083,N_10076);
nand U10355 (N_10355,N_10055,N_9956);
nand U10356 (N_10356,N_9987,N_9831);
xor U10357 (N_10357,N_10009,N_9843);
and U10358 (N_10358,N_9636,N_9966);
nand U10359 (N_10359,N_9745,N_10097);
nand U10360 (N_10360,N_10042,N_9816);
or U10361 (N_10361,N_9619,N_9747);
xnor U10362 (N_10362,N_9855,N_9690);
xnor U10363 (N_10363,N_9829,N_9873);
xor U10364 (N_10364,N_9984,N_9779);
xor U10365 (N_10365,N_10089,N_10080);
or U10366 (N_10366,N_10143,N_10003);
and U10367 (N_10367,N_9614,N_9746);
nand U10368 (N_10368,N_9908,N_9934);
nor U10369 (N_10369,N_9694,N_10085);
or U10370 (N_10370,N_9645,N_9879);
xnor U10371 (N_10371,N_9868,N_9715);
nand U10372 (N_10372,N_10038,N_9888);
xnor U10373 (N_10373,N_10058,N_9624);
or U10374 (N_10374,N_10187,N_9683);
and U10375 (N_10375,N_9733,N_9911);
nand U10376 (N_10376,N_9725,N_10110);
or U10377 (N_10377,N_9711,N_9869);
nand U10378 (N_10378,N_10153,N_9985);
xnor U10379 (N_10379,N_10011,N_9895);
or U10380 (N_10380,N_9969,N_10195);
or U10381 (N_10381,N_9996,N_9931);
or U10382 (N_10382,N_9661,N_9769);
or U10383 (N_10383,N_9749,N_10194);
nor U10384 (N_10384,N_9679,N_10036);
nor U10385 (N_10385,N_9916,N_9664);
and U10386 (N_10386,N_9811,N_9681);
nor U10387 (N_10387,N_9658,N_9932);
nand U10388 (N_10388,N_9670,N_10077);
nand U10389 (N_10389,N_9871,N_9626);
xor U10390 (N_10390,N_9864,N_10067);
nand U10391 (N_10391,N_9790,N_9768);
or U10392 (N_10392,N_9942,N_9673);
xnor U10393 (N_10393,N_10193,N_9992);
and U10394 (N_10394,N_9940,N_9894);
nand U10395 (N_10395,N_9604,N_9924);
nand U10396 (N_10396,N_9612,N_9742);
nand U10397 (N_10397,N_9951,N_9851);
and U10398 (N_10398,N_10007,N_9826);
xnor U10399 (N_10399,N_10134,N_9633);
nor U10400 (N_10400,N_9719,N_10001);
or U10401 (N_10401,N_9813,N_9959);
or U10402 (N_10402,N_10163,N_9724);
nor U10403 (N_10403,N_9978,N_9763);
and U10404 (N_10404,N_10118,N_9697);
nand U10405 (N_10405,N_9794,N_10010);
nand U10406 (N_10406,N_9696,N_10167);
or U10407 (N_10407,N_9628,N_9735);
and U10408 (N_10408,N_9936,N_9933);
xnor U10409 (N_10409,N_10154,N_9791);
and U10410 (N_10410,N_10052,N_9905);
nand U10411 (N_10411,N_9850,N_10066);
nand U10412 (N_10412,N_9753,N_10035);
or U10413 (N_10413,N_10059,N_9689);
and U10414 (N_10414,N_9915,N_9995);
and U10415 (N_10415,N_10061,N_10156);
nor U10416 (N_10416,N_9848,N_10098);
xnor U10417 (N_10417,N_10104,N_10158);
nand U10418 (N_10418,N_10005,N_9761);
nor U10419 (N_10419,N_9653,N_9964);
and U10420 (N_10420,N_10014,N_9744);
nor U10421 (N_10421,N_9892,N_9844);
or U10422 (N_10422,N_10151,N_10127);
and U10423 (N_10423,N_9634,N_9752);
nor U10424 (N_10424,N_9837,N_9901);
and U10425 (N_10425,N_9982,N_10107);
nand U10426 (N_10426,N_9841,N_9780);
or U10427 (N_10427,N_9935,N_10128);
xnor U10428 (N_10428,N_9884,N_9975);
xnor U10429 (N_10429,N_9899,N_9877);
xor U10430 (N_10430,N_10018,N_9802);
or U10431 (N_10431,N_10122,N_9714);
and U10432 (N_10432,N_9856,N_10138);
nor U10433 (N_10433,N_10074,N_10075);
xnor U10434 (N_10434,N_9629,N_9923);
or U10435 (N_10435,N_9723,N_10157);
or U10436 (N_10436,N_9765,N_9705);
nand U10437 (N_10437,N_10091,N_9706);
or U10438 (N_10438,N_9834,N_9833);
nor U10439 (N_10439,N_10103,N_9823);
nand U10440 (N_10440,N_10176,N_9875);
xor U10441 (N_10441,N_9973,N_9668);
nor U10442 (N_10442,N_9652,N_9727);
xor U10443 (N_10443,N_9929,N_9839);
nor U10444 (N_10444,N_9695,N_9682);
and U10445 (N_10445,N_9979,N_9993);
nor U10446 (N_10446,N_10081,N_9722);
or U10447 (N_10447,N_9657,N_9842);
xor U10448 (N_10448,N_9739,N_9726);
xnor U10449 (N_10449,N_9808,N_10033);
and U10450 (N_10450,N_9766,N_10160);
nand U10451 (N_10451,N_10178,N_9804);
nor U10452 (N_10452,N_9717,N_9699);
nand U10453 (N_10453,N_10069,N_9953);
and U10454 (N_10454,N_9737,N_9858);
and U10455 (N_10455,N_10024,N_9603);
nor U10456 (N_10456,N_9800,N_9774);
nand U10457 (N_10457,N_10183,N_9955);
xor U10458 (N_10458,N_10101,N_9814);
xnor U10459 (N_10459,N_10020,N_9918);
and U10460 (N_10460,N_9797,N_9859);
or U10461 (N_10461,N_9613,N_10170);
xnor U10462 (N_10462,N_9734,N_10185);
xor U10463 (N_10463,N_9963,N_10150);
and U10464 (N_10464,N_9798,N_9643);
or U10465 (N_10465,N_9617,N_9819);
nor U10466 (N_10466,N_10068,N_10152);
or U10467 (N_10467,N_9954,N_10161);
xnor U10468 (N_10468,N_9949,N_9663);
xnor U10469 (N_10469,N_10057,N_9648);
xor U10470 (N_10470,N_9885,N_9880);
nand U10471 (N_10471,N_10189,N_9941);
and U10472 (N_10472,N_10050,N_9827);
or U10473 (N_10473,N_9692,N_9701);
xnor U10474 (N_10474,N_9729,N_10180);
xor U10475 (N_10475,N_10109,N_9903);
nor U10476 (N_10476,N_10155,N_10126);
nand U10477 (N_10477,N_10064,N_10027);
or U10478 (N_10478,N_9710,N_9846);
nor U10479 (N_10479,N_9771,N_10019);
or U10480 (N_10480,N_10111,N_9677);
and U10481 (N_10481,N_9687,N_9685);
or U10482 (N_10482,N_9857,N_9772);
nand U10483 (N_10483,N_9845,N_10171);
nand U10484 (N_10484,N_9730,N_10113);
and U10485 (N_10485,N_9787,N_9751);
and U10486 (N_10486,N_9861,N_9605);
nor U10487 (N_10487,N_9708,N_10105);
or U10488 (N_10488,N_9896,N_9736);
nand U10489 (N_10489,N_10072,N_9999);
nor U10490 (N_10490,N_9807,N_9968);
and U10491 (N_10491,N_9943,N_9967);
or U10492 (N_10492,N_10168,N_9862);
nor U10493 (N_10493,N_9693,N_9937);
or U10494 (N_10494,N_9890,N_10065);
nor U10495 (N_10495,N_9921,N_10116);
nor U10496 (N_10496,N_10037,N_9602);
xor U10497 (N_10497,N_9958,N_9897);
or U10498 (N_10498,N_9971,N_9806);
nor U10499 (N_10499,N_9764,N_9731);
xor U10500 (N_10500,N_9884,N_9626);
xor U10501 (N_10501,N_9900,N_9926);
nand U10502 (N_10502,N_9637,N_9931);
or U10503 (N_10503,N_10027,N_10014);
nor U10504 (N_10504,N_9914,N_9958);
and U10505 (N_10505,N_9923,N_10086);
and U10506 (N_10506,N_9612,N_9784);
and U10507 (N_10507,N_9673,N_9775);
nand U10508 (N_10508,N_9675,N_9714);
and U10509 (N_10509,N_9861,N_9702);
nor U10510 (N_10510,N_9759,N_9706);
or U10511 (N_10511,N_9975,N_9861);
xor U10512 (N_10512,N_10092,N_9969);
nand U10513 (N_10513,N_9636,N_9702);
nand U10514 (N_10514,N_10014,N_9900);
and U10515 (N_10515,N_9716,N_10122);
or U10516 (N_10516,N_10181,N_9720);
xnor U10517 (N_10517,N_10134,N_9910);
nand U10518 (N_10518,N_9779,N_9727);
nand U10519 (N_10519,N_10163,N_10008);
and U10520 (N_10520,N_9676,N_9684);
or U10521 (N_10521,N_9901,N_9667);
or U10522 (N_10522,N_9968,N_9820);
xor U10523 (N_10523,N_10052,N_9903);
and U10524 (N_10524,N_10034,N_9692);
nand U10525 (N_10525,N_10175,N_9826);
xor U10526 (N_10526,N_9851,N_9811);
and U10527 (N_10527,N_9767,N_9616);
and U10528 (N_10528,N_9867,N_10143);
nor U10529 (N_10529,N_9906,N_9807);
and U10530 (N_10530,N_9834,N_10138);
xnor U10531 (N_10531,N_9865,N_9906);
xor U10532 (N_10532,N_9921,N_9959);
xor U10533 (N_10533,N_9815,N_9862);
nand U10534 (N_10534,N_9919,N_10157);
and U10535 (N_10535,N_10176,N_9755);
xnor U10536 (N_10536,N_10036,N_9806);
nand U10537 (N_10537,N_10112,N_9779);
xnor U10538 (N_10538,N_10196,N_9752);
nand U10539 (N_10539,N_9890,N_9749);
xnor U10540 (N_10540,N_10025,N_9634);
or U10541 (N_10541,N_10124,N_10126);
nor U10542 (N_10542,N_10054,N_9851);
nor U10543 (N_10543,N_10017,N_10083);
and U10544 (N_10544,N_9909,N_9643);
nand U10545 (N_10545,N_9705,N_9857);
nor U10546 (N_10546,N_9601,N_9785);
and U10547 (N_10547,N_9820,N_10172);
xor U10548 (N_10548,N_10167,N_10073);
and U10549 (N_10549,N_10069,N_9998);
and U10550 (N_10550,N_9946,N_9734);
xnor U10551 (N_10551,N_9881,N_9922);
nand U10552 (N_10552,N_9759,N_9860);
nor U10553 (N_10553,N_9769,N_9876);
or U10554 (N_10554,N_10191,N_9825);
nor U10555 (N_10555,N_9936,N_9761);
xnor U10556 (N_10556,N_9730,N_10131);
or U10557 (N_10557,N_9728,N_9755);
xor U10558 (N_10558,N_9902,N_10088);
xor U10559 (N_10559,N_9719,N_10188);
or U10560 (N_10560,N_10137,N_9954);
or U10561 (N_10561,N_9774,N_10120);
nand U10562 (N_10562,N_9823,N_9732);
and U10563 (N_10563,N_10096,N_10084);
nor U10564 (N_10564,N_9984,N_9750);
xnor U10565 (N_10565,N_10194,N_9932);
nor U10566 (N_10566,N_9974,N_10041);
xor U10567 (N_10567,N_10079,N_10139);
nand U10568 (N_10568,N_9789,N_10094);
or U10569 (N_10569,N_10016,N_9651);
nor U10570 (N_10570,N_9906,N_10108);
or U10571 (N_10571,N_9849,N_9679);
or U10572 (N_10572,N_10157,N_10076);
and U10573 (N_10573,N_9627,N_9666);
and U10574 (N_10574,N_9728,N_10038);
or U10575 (N_10575,N_9948,N_10027);
nand U10576 (N_10576,N_10171,N_10157);
nand U10577 (N_10577,N_10048,N_10172);
xor U10578 (N_10578,N_9699,N_9645);
xor U10579 (N_10579,N_9795,N_9724);
nor U10580 (N_10580,N_9754,N_10199);
or U10581 (N_10581,N_9611,N_9665);
xor U10582 (N_10582,N_10114,N_9889);
and U10583 (N_10583,N_9807,N_9761);
or U10584 (N_10584,N_10038,N_9842);
nand U10585 (N_10585,N_9813,N_9690);
and U10586 (N_10586,N_9750,N_9872);
nand U10587 (N_10587,N_9753,N_10023);
and U10588 (N_10588,N_9616,N_9951);
nor U10589 (N_10589,N_9978,N_9631);
nand U10590 (N_10590,N_10169,N_10138);
nor U10591 (N_10591,N_9722,N_9996);
xor U10592 (N_10592,N_9927,N_10198);
and U10593 (N_10593,N_9919,N_9636);
and U10594 (N_10594,N_9683,N_9815);
nor U10595 (N_10595,N_9941,N_9860);
xor U10596 (N_10596,N_10159,N_9826);
and U10597 (N_10597,N_9820,N_9898);
and U10598 (N_10598,N_9868,N_10147);
nor U10599 (N_10599,N_9636,N_9811);
nand U10600 (N_10600,N_9651,N_9917);
and U10601 (N_10601,N_9966,N_9870);
and U10602 (N_10602,N_9842,N_9749);
and U10603 (N_10603,N_9668,N_10118);
nand U10604 (N_10604,N_9605,N_10018);
nor U10605 (N_10605,N_9929,N_9942);
nor U10606 (N_10606,N_9847,N_10115);
nor U10607 (N_10607,N_9813,N_9930);
and U10608 (N_10608,N_9977,N_9895);
or U10609 (N_10609,N_9830,N_9737);
nand U10610 (N_10610,N_9628,N_10020);
nor U10611 (N_10611,N_9939,N_9865);
and U10612 (N_10612,N_9819,N_9935);
nand U10613 (N_10613,N_9890,N_10026);
nand U10614 (N_10614,N_9729,N_9980);
nand U10615 (N_10615,N_10048,N_9778);
nor U10616 (N_10616,N_9657,N_9646);
nand U10617 (N_10617,N_10012,N_9810);
or U10618 (N_10618,N_9941,N_10099);
nor U10619 (N_10619,N_9808,N_9988);
and U10620 (N_10620,N_9961,N_9908);
nand U10621 (N_10621,N_9680,N_10103);
or U10622 (N_10622,N_9749,N_9946);
and U10623 (N_10623,N_9638,N_9929);
xor U10624 (N_10624,N_9996,N_10008);
or U10625 (N_10625,N_9889,N_10016);
or U10626 (N_10626,N_10066,N_10005);
xor U10627 (N_10627,N_9711,N_9736);
nor U10628 (N_10628,N_10140,N_9616);
xnor U10629 (N_10629,N_9636,N_9876);
nand U10630 (N_10630,N_9700,N_10168);
and U10631 (N_10631,N_10101,N_9653);
or U10632 (N_10632,N_9874,N_9869);
nor U10633 (N_10633,N_9959,N_9782);
or U10634 (N_10634,N_9857,N_9815);
and U10635 (N_10635,N_9774,N_9738);
xnor U10636 (N_10636,N_9972,N_9678);
or U10637 (N_10637,N_9787,N_9948);
and U10638 (N_10638,N_9963,N_9714);
nand U10639 (N_10639,N_9710,N_9662);
and U10640 (N_10640,N_9762,N_9725);
nand U10641 (N_10641,N_9707,N_9657);
nor U10642 (N_10642,N_10046,N_9656);
or U10643 (N_10643,N_10008,N_9791);
or U10644 (N_10644,N_10153,N_9830);
or U10645 (N_10645,N_10041,N_9709);
nor U10646 (N_10646,N_9702,N_10180);
nor U10647 (N_10647,N_9782,N_10033);
and U10648 (N_10648,N_9787,N_9989);
nor U10649 (N_10649,N_10158,N_9913);
nor U10650 (N_10650,N_9982,N_9950);
xor U10651 (N_10651,N_9732,N_9752);
xnor U10652 (N_10652,N_9681,N_10164);
xnor U10653 (N_10653,N_9682,N_9750);
nand U10654 (N_10654,N_9777,N_9609);
and U10655 (N_10655,N_9749,N_10132);
nor U10656 (N_10656,N_10000,N_9707);
nor U10657 (N_10657,N_9708,N_9926);
nor U10658 (N_10658,N_9797,N_9854);
or U10659 (N_10659,N_10192,N_10145);
nand U10660 (N_10660,N_9703,N_9959);
nand U10661 (N_10661,N_9771,N_9625);
or U10662 (N_10662,N_10152,N_9879);
or U10663 (N_10663,N_9921,N_9894);
or U10664 (N_10664,N_9870,N_9650);
nor U10665 (N_10665,N_9767,N_9914);
and U10666 (N_10666,N_9657,N_10038);
nor U10667 (N_10667,N_10169,N_9837);
nor U10668 (N_10668,N_9740,N_9913);
nor U10669 (N_10669,N_10027,N_10142);
nand U10670 (N_10670,N_10051,N_9896);
nor U10671 (N_10671,N_9898,N_10140);
nand U10672 (N_10672,N_10050,N_9722);
nor U10673 (N_10673,N_10059,N_9718);
and U10674 (N_10674,N_9722,N_9652);
or U10675 (N_10675,N_9984,N_9626);
or U10676 (N_10676,N_10081,N_9627);
xnor U10677 (N_10677,N_10141,N_9927);
nand U10678 (N_10678,N_9978,N_10083);
or U10679 (N_10679,N_9645,N_9947);
nand U10680 (N_10680,N_9912,N_9862);
nand U10681 (N_10681,N_9723,N_9982);
xnor U10682 (N_10682,N_10090,N_9879);
or U10683 (N_10683,N_9867,N_9663);
nand U10684 (N_10684,N_9968,N_9642);
nor U10685 (N_10685,N_9663,N_10149);
nand U10686 (N_10686,N_9666,N_9863);
and U10687 (N_10687,N_9761,N_10084);
xnor U10688 (N_10688,N_9973,N_10001);
and U10689 (N_10689,N_10120,N_9871);
nor U10690 (N_10690,N_9661,N_10099);
nand U10691 (N_10691,N_9629,N_9699);
and U10692 (N_10692,N_9908,N_9781);
and U10693 (N_10693,N_9750,N_9711);
or U10694 (N_10694,N_9603,N_9695);
or U10695 (N_10695,N_10002,N_10025);
nand U10696 (N_10696,N_10000,N_9984);
xnor U10697 (N_10697,N_10118,N_9852);
nor U10698 (N_10698,N_9798,N_9971);
nand U10699 (N_10699,N_9965,N_10098);
nor U10700 (N_10700,N_9955,N_9694);
nor U10701 (N_10701,N_9789,N_9777);
nand U10702 (N_10702,N_10039,N_9633);
and U10703 (N_10703,N_9779,N_9746);
nand U10704 (N_10704,N_9731,N_9707);
or U10705 (N_10705,N_10090,N_9718);
or U10706 (N_10706,N_9724,N_9711);
xor U10707 (N_10707,N_9762,N_9870);
nand U10708 (N_10708,N_10187,N_9946);
nor U10709 (N_10709,N_9750,N_9855);
nor U10710 (N_10710,N_10074,N_9849);
or U10711 (N_10711,N_9949,N_9657);
nand U10712 (N_10712,N_10083,N_9613);
nor U10713 (N_10713,N_9600,N_9878);
xor U10714 (N_10714,N_10081,N_9900);
nor U10715 (N_10715,N_10099,N_9634);
or U10716 (N_10716,N_10033,N_10072);
xnor U10717 (N_10717,N_9634,N_9867);
nand U10718 (N_10718,N_9671,N_9807);
nand U10719 (N_10719,N_9778,N_10069);
nor U10720 (N_10720,N_9602,N_9774);
nor U10721 (N_10721,N_9848,N_9623);
nand U10722 (N_10722,N_10002,N_9889);
nand U10723 (N_10723,N_9691,N_9662);
nand U10724 (N_10724,N_9615,N_10015);
nor U10725 (N_10725,N_10185,N_9743);
nor U10726 (N_10726,N_9998,N_10144);
xor U10727 (N_10727,N_10053,N_10186);
nand U10728 (N_10728,N_9729,N_10057);
xor U10729 (N_10729,N_10156,N_10144);
or U10730 (N_10730,N_10106,N_9785);
and U10731 (N_10731,N_9602,N_9868);
or U10732 (N_10732,N_10188,N_9748);
xnor U10733 (N_10733,N_9697,N_10099);
and U10734 (N_10734,N_9871,N_10096);
xnor U10735 (N_10735,N_9940,N_9764);
xnor U10736 (N_10736,N_9927,N_9906);
xor U10737 (N_10737,N_9636,N_9646);
xnor U10738 (N_10738,N_9646,N_9967);
and U10739 (N_10739,N_9876,N_9895);
nand U10740 (N_10740,N_9932,N_9742);
and U10741 (N_10741,N_9911,N_10061);
or U10742 (N_10742,N_9778,N_9697);
or U10743 (N_10743,N_9610,N_10015);
nand U10744 (N_10744,N_9917,N_9684);
or U10745 (N_10745,N_10027,N_9702);
nor U10746 (N_10746,N_9662,N_9939);
or U10747 (N_10747,N_9962,N_9776);
nor U10748 (N_10748,N_9686,N_10130);
or U10749 (N_10749,N_10085,N_9936);
or U10750 (N_10750,N_9666,N_10183);
nand U10751 (N_10751,N_9619,N_10017);
or U10752 (N_10752,N_10124,N_9791);
nand U10753 (N_10753,N_10109,N_9704);
and U10754 (N_10754,N_9841,N_10122);
and U10755 (N_10755,N_9984,N_10174);
xor U10756 (N_10756,N_10127,N_10149);
nor U10757 (N_10757,N_10043,N_9947);
nand U10758 (N_10758,N_10114,N_10036);
nand U10759 (N_10759,N_9793,N_9718);
nand U10760 (N_10760,N_9761,N_9876);
or U10761 (N_10761,N_9736,N_10159);
or U10762 (N_10762,N_9770,N_10077);
or U10763 (N_10763,N_10032,N_10035);
or U10764 (N_10764,N_10138,N_9867);
nand U10765 (N_10765,N_10045,N_9931);
and U10766 (N_10766,N_10135,N_10057);
and U10767 (N_10767,N_10153,N_10050);
xnor U10768 (N_10768,N_9856,N_9957);
nand U10769 (N_10769,N_10084,N_9963);
and U10770 (N_10770,N_9767,N_9975);
nor U10771 (N_10771,N_10164,N_10195);
xor U10772 (N_10772,N_9761,N_10190);
and U10773 (N_10773,N_9840,N_9679);
xor U10774 (N_10774,N_9862,N_10133);
nor U10775 (N_10775,N_9745,N_10194);
and U10776 (N_10776,N_9791,N_9857);
nand U10777 (N_10777,N_9789,N_9733);
and U10778 (N_10778,N_9628,N_10116);
and U10779 (N_10779,N_10028,N_10141);
xnor U10780 (N_10780,N_9745,N_9690);
or U10781 (N_10781,N_10041,N_9652);
nand U10782 (N_10782,N_10009,N_10064);
nand U10783 (N_10783,N_9722,N_9761);
nor U10784 (N_10784,N_9979,N_9654);
xor U10785 (N_10785,N_9879,N_9857);
xor U10786 (N_10786,N_9861,N_9780);
nand U10787 (N_10787,N_10195,N_9738);
or U10788 (N_10788,N_9693,N_9876);
or U10789 (N_10789,N_10157,N_9921);
nor U10790 (N_10790,N_9690,N_9789);
xor U10791 (N_10791,N_10025,N_10170);
nand U10792 (N_10792,N_9942,N_9932);
or U10793 (N_10793,N_10118,N_10008);
and U10794 (N_10794,N_9952,N_9754);
xor U10795 (N_10795,N_10005,N_9898);
xor U10796 (N_10796,N_9945,N_10094);
and U10797 (N_10797,N_10126,N_9780);
and U10798 (N_10798,N_10075,N_9956);
nor U10799 (N_10799,N_9725,N_9917);
and U10800 (N_10800,N_10350,N_10451);
and U10801 (N_10801,N_10556,N_10440);
and U10802 (N_10802,N_10318,N_10676);
nor U10803 (N_10803,N_10373,N_10678);
xor U10804 (N_10804,N_10494,N_10763);
nor U10805 (N_10805,N_10206,N_10796);
or U10806 (N_10806,N_10308,N_10477);
and U10807 (N_10807,N_10755,N_10201);
xnor U10808 (N_10808,N_10718,N_10468);
and U10809 (N_10809,N_10250,N_10534);
or U10810 (N_10810,N_10307,N_10243);
nor U10811 (N_10811,N_10341,N_10479);
or U10812 (N_10812,N_10405,N_10654);
xor U10813 (N_10813,N_10359,N_10649);
and U10814 (N_10814,N_10524,N_10708);
and U10815 (N_10815,N_10411,N_10400);
and U10816 (N_10816,N_10358,N_10490);
xor U10817 (N_10817,N_10784,N_10563);
or U10818 (N_10818,N_10404,N_10203);
and U10819 (N_10819,N_10735,N_10728);
nand U10820 (N_10820,N_10785,N_10261);
nand U10821 (N_10821,N_10329,N_10268);
and U10822 (N_10822,N_10255,N_10566);
and U10823 (N_10823,N_10464,N_10497);
or U10824 (N_10824,N_10576,N_10586);
or U10825 (N_10825,N_10284,N_10366);
nand U10826 (N_10826,N_10377,N_10661);
or U10827 (N_10827,N_10722,N_10474);
and U10828 (N_10828,N_10221,N_10651);
nand U10829 (N_10829,N_10275,N_10627);
xor U10830 (N_10830,N_10500,N_10395);
nor U10831 (N_10831,N_10344,N_10484);
and U10832 (N_10832,N_10752,N_10634);
or U10833 (N_10833,N_10239,N_10273);
nor U10834 (N_10834,N_10629,N_10548);
nand U10835 (N_10835,N_10657,N_10636);
nor U10836 (N_10836,N_10381,N_10449);
nor U10837 (N_10837,N_10697,N_10444);
nor U10838 (N_10838,N_10711,N_10383);
nor U10839 (N_10839,N_10232,N_10443);
or U10840 (N_10840,N_10648,N_10496);
nand U10841 (N_10841,N_10541,N_10675);
or U10842 (N_10842,N_10592,N_10355);
xor U10843 (N_10843,N_10633,N_10776);
and U10844 (N_10844,N_10367,N_10594);
and U10845 (N_10845,N_10683,N_10709);
or U10846 (N_10846,N_10288,N_10672);
nor U10847 (N_10847,N_10253,N_10228);
and U10848 (N_10848,N_10768,N_10260);
xnor U10849 (N_10849,N_10388,N_10567);
nor U10850 (N_10850,N_10605,N_10336);
nand U10851 (N_10851,N_10271,N_10274);
nand U10852 (N_10852,N_10608,N_10364);
and U10853 (N_10853,N_10237,N_10356);
and U10854 (N_10854,N_10354,N_10481);
nand U10855 (N_10855,N_10701,N_10674);
or U10856 (N_10856,N_10795,N_10687);
and U10857 (N_10857,N_10655,N_10475);
or U10858 (N_10858,N_10458,N_10517);
or U10859 (N_10859,N_10345,N_10418);
nor U10860 (N_10860,N_10281,N_10276);
or U10861 (N_10861,N_10278,N_10339);
nand U10862 (N_10862,N_10585,N_10421);
or U10863 (N_10863,N_10300,N_10348);
or U10864 (N_10864,N_10736,N_10615);
nor U10865 (N_10865,N_10721,N_10542);
nor U10866 (N_10866,N_10272,N_10422);
or U10867 (N_10867,N_10425,N_10466);
nand U10868 (N_10868,N_10287,N_10782);
nand U10869 (N_10869,N_10595,N_10311);
xnor U10870 (N_10870,N_10323,N_10489);
xnor U10871 (N_10871,N_10771,N_10414);
xnor U10872 (N_10872,N_10705,N_10387);
and U10873 (N_10873,N_10673,N_10378);
nand U10874 (N_10874,N_10719,N_10445);
and U10875 (N_10875,N_10682,N_10390);
xor U10876 (N_10876,N_10505,N_10270);
xor U10877 (N_10877,N_10770,N_10393);
or U10878 (N_10878,N_10342,N_10266);
xnor U10879 (N_10879,N_10251,N_10320);
nand U10880 (N_10880,N_10453,N_10392);
or U10881 (N_10881,N_10580,N_10536);
and U10882 (N_10882,N_10787,N_10551);
or U10883 (N_10883,N_10745,N_10360);
and U10884 (N_10884,N_10603,N_10562);
and U10885 (N_10885,N_10365,N_10666);
nand U10886 (N_10886,N_10290,N_10423);
nor U10887 (N_10887,N_10609,N_10315);
xnor U10888 (N_10888,N_10503,N_10502);
xnor U10889 (N_10889,N_10783,N_10470);
nor U10890 (N_10890,N_10498,N_10463);
nor U10891 (N_10891,N_10408,N_10547);
nand U10892 (N_10892,N_10611,N_10428);
or U10893 (N_10893,N_10429,N_10321);
and U10894 (N_10894,N_10733,N_10616);
or U10895 (N_10895,N_10600,N_10431);
nor U10896 (N_10896,N_10406,N_10205);
xnor U10897 (N_10897,N_10244,N_10695);
nor U10898 (N_10898,N_10349,N_10249);
or U10899 (N_10899,N_10679,N_10762);
nor U10900 (N_10900,N_10375,N_10434);
nor U10901 (N_10901,N_10412,N_10297);
and U10902 (N_10902,N_10696,N_10769);
nor U10903 (N_10903,N_10773,N_10658);
or U10904 (N_10904,N_10749,N_10650);
and U10905 (N_10905,N_10508,N_10637);
xor U10906 (N_10906,N_10545,N_10647);
and U10907 (N_10907,N_10372,N_10664);
nor U10908 (N_10908,N_10732,N_10645);
nand U10909 (N_10909,N_10471,N_10461);
xor U10910 (N_10910,N_10706,N_10472);
nand U10911 (N_10911,N_10280,N_10361);
and U10912 (N_10912,N_10277,N_10368);
or U10913 (N_10913,N_10791,N_10671);
or U10914 (N_10914,N_10699,N_10382);
and U10915 (N_10915,N_10402,N_10564);
nand U10916 (N_10916,N_10779,N_10513);
and U10917 (N_10917,N_10766,N_10691);
and U10918 (N_10918,N_10240,N_10758);
xnor U10919 (N_10919,N_10501,N_10415);
nand U10920 (N_10920,N_10764,N_10371);
xnor U10921 (N_10921,N_10242,N_10426);
and U10922 (N_10922,N_10519,N_10606);
and U10923 (N_10923,N_10739,N_10639);
nand U10924 (N_10924,N_10570,N_10238);
nand U10925 (N_10925,N_10430,N_10495);
or U10926 (N_10926,N_10293,N_10690);
nand U10927 (N_10927,N_10312,N_10235);
nor U10928 (N_10928,N_10553,N_10224);
nor U10929 (N_10929,N_10557,N_10227);
nor U10930 (N_10930,N_10401,N_10598);
or U10931 (N_10931,N_10642,N_10202);
or U10932 (N_10932,N_10700,N_10760);
nor U10933 (N_10933,N_10712,N_10630);
nand U10934 (N_10934,N_10663,N_10427);
or U10935 (N_10935,N_10537,N_10473);
xor U10936 (N_10936,N_10767,N_10511);
and U10937 (N_10937,N_10579,N_10209);
xor U10938 (N_10938,N_10236,N_10295);
and U10939 (N_10939,N_10741,N_10535);
xor U10940 (N_10940,N_10680,N_10743);
and U10941 (N_10941,N_10447,N_10689);
or U10942 (N_10942,N_10759,N_10327);
xnor U10943 (N_10943,N_10554,N_10317);
nand U10944 (N_10944,N_10413,N_10338);
nand U10945 (N_10945,N_10593,N_10510);
xor U10946 (N_10946,N_10573,N_10283);
nand U10947 (N_10947,N_10219,N_10248);
xor U10948 (N_10948,N_10226,N_10581);
nand U10949 (N_10949,N_10319,N_10407);
xnor U10950 (N_10950,N_10460,N_10643);
nor U10951 (N_10951,N_10313,N_10296);
xnor U10952 (N_10952,N_10459,N_10644);
nor U10953 (N_10953,N_10265,N_10222);
xor U10954 (N_10954,N_10362,N_10589);
nor U10955 (N_10955,N_10493,N_10399);
xor U10956 (N_10956,N_10525,N_10761);
or U10957 (N_10957,N_10750,N_10546);
xor U10958 (N_10958,N_10625,N_10246);
or U10959 (N_10959,N_10544,N_10638);
xor U10960 (N_10960,N_10754,N_10702);
nor U10961 (N_10961,N_10619,N_10436);
nor U10962 (N_10962,N_10374,N_10488);
and U10963 (N_10963,N_10204,N_10716);
nor U10964 (N_10964,N_10569,N_10578);
nor U10965 (N_10965,N_10397,N_10291);
or U10966 (N_10966,N_10439,N_10515);
nor U10967 (N_10967,N_10379,N_10279);
nor U10968 (N_10968,N_10725,N_10538);
nor U10969 (N_10969,N_10624,N_10765);
or U10970 (N_10970,N_10455,N_10792);
and U10971 (N_10971,N_10301,N_10607);
nor U10972 (N_10972,N_10211,N_10499);
and U10973 (N_10973,N_10668,N_10631);
xnor U10974 (N_10974,N_10245,N_10324);
nor U10975 (N_10975,N_10568,N_10748);
nor U10976 (N_10976,N_10335,N_10516);
and U10977 (N_10977,N_10207,N_10480);
nand U10978 (N_10978,N_10467,N_10487);
or U10979 (N_10979,N_10234,N_10386);
nor U10980 (N_10980,N_10730,N_10376);
or U10981 (N_10981,N_10522,N_10703);
xnor U10982 (N_10982,N_10457,N_10756);
and U10983 (N_10983,N_10230,N_10714);
nand U10984 (N_10984,N_10604,N_10332);
and U10985 (N_10985,N_10417,N_10640);
nand U10986 (N_10986,N_10757,N_10707);
nor U10987 (N_10987,N_10737,N_10613);
or U10988 (N_10988,N_10628,N_10257);
nor U10989 (N_10989,N_10208,N_10521);
and U10990 (N_10990,N_10740,N_10662);
nand U10991 (N_10991,N_10384,N_10282);
and U10992 (N_10992,N_10292,N_10575);
and U10993 (N_10993,N_10433,N_10231);
and U10994 (N_10994,N_10316,N_10491);
nand U10995 (N_10995,N_10256,N_10591);
and U10996 (N_10996,N_10210,N_10688);
and U10997 (N_10997,N_10326,N_10778);
nand U10998 (N_10998,N_10622,N_10482);
or U10999 (N_10999,N_10533,N_10247);
and U11000 (N_11000,N_10396,N_10596);
xnor U11001 (N_11001,N_10310,N_10555);
nand U11002 (N_11002,N_10322,N_10420);
or U11003 (N_11003,N_10529,N_10303);
nand U11004 (N_11004,N_10610,N_10602);
nor U11005 (N_11005,N_10797,N_10789);
or U11006 (N_11006,N_10478,N_10217);
and U11007 (N_11007,N_10777,N_10469);
and U11008 (N_11008,N_10262,N_10685);
and U11009 (N_11009,N_10485,N_10693);
and U11010 (N_11010,N_10456,N_10552);
nor U11011 (N_11011,N_10794,N_10419);
or U11012 (N_11012,N_10370,N_10220);
and U11013 (N_11013,N_10462,N_10684);
nor U11014 (N_11014,N_10223,N_10744);
nand U11015 (N_11015,N_10790,N_10465);
or U11016 (N_11016,N_10723,N_10286);
and U11017 (N_11017,N_10530,N_10799);
xor U11018 (N_11018,N_10669,N_10729);
nand U11019 (N_11019,N_10670,N_10786);
or U11020 (N_11020,N_10528,N_10410);
and U11021 (N_11021,N_10442,N_10233);
nand U11022 (N_11022,N_10263,N_10632);
and U11023 (N_11023,N_10539,N_10333);
or U11024 (N_11024,N_10652,N_10352);
and U11025 (N_11025,N_10656,N_10599);
nand U11026 (N_11026,N_10572,N_10588);
nand U11027 (N_11027,N_10518,N_10438);
xor U11028 (N_11028,N_10492,N_10351);
xnor U11029 (N_11029,N_10681,N_10294);
xor U11030 (N_11030,N_10686,N_10582);
nor U11031 (N_11031,N_10617,N_10724);
xor U11032 (N_11032,N_10738,N_10446);
nand U11033 (N_11033,N_10450,N_10483);
xor U11034 (N_11034,N_10774,N_10549);
or U11035 (N_11035,N_10357,N_10571);
or U11036 (N_11036,N_10403,N_10710);
nor U11037 (N_11037,N_10330,N_10646);
xnor U11038 (N_11038,N_10612,N_10432);
or U11039 (N_11039,N_10583,N_10660);
nor U11040 (N_11040,N_10309,N_10742);
or U11041 (N_11041,N_10259,N_10254);
and U11042 (N_11042,N_10452,N_10213);
xor U11043 (N_11043,N_10340,N_10653);
nor U11044 (N_11044,N_10531,N_10731);
nor U11045 (N_11045,N_10424,N_10574);
and U11046 (N_11046,N_10512,N_10713);
nor U11047 (N_11047,N_10264,N_10526);
nand U11048 (N_11048,N_10550,N_10398);
nor U11049 (N_11049,N_10314,N_10698);
nand U11050 (N_11050,N_10577,N_10258);
or U11051 (N_11051,N_10726,N_10346);
nand U11052 (N_11052,N_10734,N_10793);
and U11053 (N_11053,N_10641,N_10561);
nand U11054 (N_11054,N_10218,N_10704);
and U11055 (N_11055,N_10241,N_10601);
xor U11056 (N_11056,N_10380,N_10781);
nor U11057 (N_11057,N_10635,N_10788);
xor U11058 (N_11058,N_10775,N_10394);
xor U11059 (N_11059,N_10559,N_10665);
or U11060 (N_11060,N_10597,N_10618);
nand U11061 (N_11061,N_10435,N_10298);
nand U11062 (N_11062,N_10385,N_10780);
and U11063 (N_11063,N_10343,N_10506);
or U11064 (N_11064,N_10289,N_10565);
nand U11065 (N_11065,N_10353,N_10299);
or U11066 (N_11066,N_10751,N_10389);
xor U11067 (N_11067,N_10523,N_10325);
or U11068 (N_11068,N_10659,N_10747);
xnor U11069 (N_11069,N_10626,N_10363);
nand U11070 (N_11070,N_10304,N_10614);
nand U11071 (N_11071,N_10532,N_10328);
nand U11072 (N_11072,N_10448,N_10269);
nand U11073 (N_11073,N_10543,N_10391);
or U11074 (N_11074,N_10558,N_10677);
nor U11075 (N_11075,N_10216,N_10798);
xnor U11076 (N_11076,N_10212,N_10305);
or U11077 (N_11077,N_10302,N_10667);
nand U11078 (N_11078,N_10331,N_10509);
and U11079 (N_11079,N_10337,N_10520);
and U11080 (N_11080,N_10441,N_10409);
xnor U11081 (N_11081,N_10486,N_10504);
xnor U11082 (N_11082,N_10590,N_10623);
and U11083 (N_11083,N_10334,N_10692);
nor U11084 (N_11084,N_10587,N_10514);
or U11085 (N_11085,N_10560,N_10437);
xor U11086 (N_11086,N_10267,N_10200);
xnor U11087 (N_11087,N_10285,N_10476);
xor U11088 (N_11088,N_10772,N_10369);
nor U11089 (N_11089,N_10527,N_10717);
or U11090 (N_11090,N_10252,N_10225);
xor U11091 (N_11091,N_10584,N_10229);
xor U11092 (N_11092,N_10620,N_10540);
nor U11093 (N_11093,N_10621,N_10416);
nand U11094 (N_11094,N_10746,N_10720);
and U11095 (N_11095,N_10715,N_10507);
xnor U11096 (N_11096,N_10454,N_10347);
xor U11097 (N_11097,N_10215,N_10214);
and U11098 (N_11098,N_10753,N_10694);
nor U11099 (N_11099,N_10727,N_10306);
nor U11100 (N_11100,N_10742,N_10641);
xor U11101 (N_11101,N_10673,N_10716);
xnor U11102 (N_11102,N_10620,N_10665);
xnor U11103 (N_11103,N_10381,N_10583);
and U11104 (N_11104,N_10725,N_10569);
xnor U11105 (N_11105,N_10388,N_10780);
or U11106 (N_11106,N_10462,N_10731);
nor U11107 (N_11107,N_10453,N_10506);
or U11108 (N_11108,N_10647,N_10555);
nand U11109 (N_11109,N_10591,N_10682);
nand U11110 (N_11110,N_10629,N_10617);
nor U11111 (N_11111,N_10338,N_10500);
nand U11112 (N_11112,N_10549,N_10300);
nor U11113 (N_11113,N_10549,N_10521);
xnor U11114 (N_11114,N_10651,N_10383);
and U11115 (N_11115,N_10756,N_10718);
or U11116 (N_11116,N_10768,N_10504);
xnor U11117 (N_11117,N_10574,N_10578);
or U11118 (N_11118,N_10281,N_10598);
nor U11119 (N_11119,N_10730,N_10617);
nor U11120 (N_11120,N_10298,N_10687);
nor U11121 (N_11121,N_10777,N_10740);
and U11122 (N_11122,N_10486,N_10218);
nand U11123 (N_11123,N_10325,N_10318);
xnor U11124 (N_11124,N_10526,N_10202);
nand U11125 (N_11125,N_10243,N_10345);
or U11126 (N_11126,N_10567,N_10437);
and U11127 (N_11127,N_10348,N_10211);
and U11128 (N_11128,N_10414,N_10318);
xnor U11129 (N_11129,N_10291,N_10243);
or U11130 (N_11130,N_10680,N_10634);
nand U11131 (N_11131,N_10262,N_10702);
nor U11132 (N_11132,N_10398,N_10582);
nand U11133 (N_11133,N_10618,N_10304);
or U11134 (N_11134,N_10768,N_10331);
xnor U11135 (N_11135,N_10226,N_10603);
or U11136 (N_11136,N_10546,N_10284);
xnor U11137 (N_11137,N_10486,N_10401);
or U11138 (N_11138,N_10582,N_10716);
and U11139 (N_11139,N_10659,N_10605);
nor U11140 (N_11140,N_10421,N_10259);
or U11141 (N_11141,N_10314,N_10425);
and U11142 (N_11142,N_10780,N_10319);
or U11143 (N_11143,N_10756,N_10234);
nor U11144 (N_11144,N_10248,N_10353);
nor U11145 (N_11145,N_10527,N_10458);
or U11146 (N_11146,N_10246,N_10431);
nand U11147 (N_11147,N_10295,N_10314);
and U11148 (N_11148,N_10671,N_10704);
nor U11149 (N_11149,N_10453,N_10489);
or U11150 (N_11150,N_10267,N_10730);
nor U11151 (N_11151,N_10471,N_10238);
nand U11152 (N_11152,N_10574,N_10289);
nand U11153 (N_11153,N_10367,N_10778);
nor U11154 (N_11154,N_10305,N_10459);
nor U11155 (N_11155,N_10539,N_10719);
nor U11156 (N_11156,N_10649,N_10791);
xor U11157 (N_11157,N_10420,N_10447);
or U11158 (N_11158,N_10274,N_10777);
and U11159 (N_11159,N_10729,N_10291);
nand U11160 (N_11160,N_10751,N_10231);
or U11161 (N_11161,N_10377,N_10748);
and U11162 (N_11162,N_10397,N_10384);
or U11163 (N_11163,N_10378,N_10660);
xor U11164 (N_11164,N_10511,N_10758);
or U11165 (N_11165,N_10222,N_10518);
nand U11166 (N_11166,N_10711,N_10685);
xnor U11167 (N_11167,N_10690,N_10699);
nand U11168 (N_11168,N_10422,N_10271);
nand U11169 (N_11169,N_10549,N_10348);
nand U11170 (N_11170,N_10397,N_10324);
or U11171 (N_11171,N_10317,N_10662);
nand U11172 (N_11172,N_10625,N_10498);
or U11173 (N_11173,N_10416,N_10615);
or U11174 (N_11174,N_10758,N_10489);
xor U11175 (N_11175,N_10311,N_10346);
xor U11176 (N_11176,N_10200,N_10691);
nand U11177 (N_11177,N_10268,N_10512);
and U11178 (N_11178,N_10749,N_10698);
and U11179 (N_11179,N_10720,N_10540);
xor U11180 (N_11180,N_10526,N_10688);
nor U11181 (N_11181,N_10477,N_10648);
or U11182 (N_11182,N_10382,N_10593);
xor U11183 (N_11183,N_10557,N_10221);
xnor U11184 (N_11184,N_10675,N_10762);
nor U11185 (N_11185,N_10338,N_10347);
nor U11186 (N_11186,N_10481,N_10217);
nand U11187 (N_11187,N_10756,N_10726);
and U11188 (N_11188,N_10582,N_10545);
or U11189 (N_11189,N_10788,N_10705);
and U11190 (N_11190,N_10227,N_10686);
xor U11191 (N_11191,N_10766,N_10523);
or U11192 (N_11192,N_10425,N_10418);
xor U11193 (N_11193,N_10343,N_10720);
xor U11194 (N_11194,N_10242,N_10559);
or U11195 (N_11195,N_10295,N_10673);
and U11196 (N_11196,N_10410,N_10214);
and U11197 (N_11197,N_10448,N_10205);
xnor U11198 (N_11198,N_10418,N_10268);
or U11199 (N_11199,N_10542,N_10404);
and U11200 (N_11200,N_10307,N_10627);
and U11201 (N_11201,N_10211,N_10343);
xor U11202 (N_11202,N_10249,N_10255);
or U11203 (N_11203,N_10703,N_10455);
nor U11204 (N_11204,N_10317,N_10316);
nor U11205 (N_11205,N_10231,N_10465);
and U11206 (N_11206,N_10705,N_10440);
nor U11207 (N_11207,N_10648,N_10374);
xnor U11208 (N_11208,N_10490,N_10709);
or U11209 (N_11209,N_10228,N_10608);
nand U11210 (N_11210,N_10461,N_10770);
or U11211 (N_11211,N_10422,N_10424);
nand U11212 (N_11212,N_10220,N_10506);
nor U11213 (N_11213,N_10556,N_10523);
or U11214 (N_11214,N_10422,N_10516);
and U11215 (N_11215,N_10388,N_10492);
nor U11216 (N_11216,N_10290,N_10621);
or U11217 (N_11217,N_10608,N_10740);
nand U11218 (N_11218,N_10790,N_10231);
nand U11219 (N_11219,N_10281,N_10774);
and U11220 (N_11220,N_10691,N_10679);
xnor U11221 (N_11221,N_10775,N_10789);
xor U11222 (N_11222,N_10238,N_10671);
xor U11223 (N_11223,N_10224,N_10483);
xnor U11224 (N_11224,N_10340,N_10496);
nand U11225 (N_11225,N_10351,N_10313);
nand U11226 (N_11226,N_10588,N_10695);
nand U11227 (N_11227,N_10450,N_10383);
xor U11228 (N_11228,N_10411,N_10586);
nor U11229 (N_11229,N_10761,N_10285);
xor U11230 (N_11230,N_10324,N_10517);
and U11231 (N_11231,N_10612,N_10352);
xor U11232 (N_11232,N_10504,N_10446);
xnor U11233 (N_11233,N_10724,N_10613);
nand U11234 (N_11234,N_10462,N_10719);
xnor U11235 (N_11235,N_10361,N_10246);
nand U11236 (N_11236,N_10796,N_10584);
nand U11237 (N_11237,N_10685,N_10634);
nand U11238 (N_11238,N_10495,N_10374);
and U11239 (N_11239,N_10614,N_10265);
nand U11240 (N_11240,N_10443,N_10449);
nor U11241 (N_11241,N_10474,N_10259);
or U11242 (N_11242,N_10799,N_10753);
nor U11243 (N_11243,N_10687,N_10203);
nand U11244 (N_11244,N_10704,N_10394);
xor U11245 (N_11245,N_10451,N_10237);
or U11246 (N_11246,N_10786,N_10220);
xnor U11247 (N_11247,N_10788,N_10341);
and U11248 (N_11248,N_10320,N_10476);
nand U11249 (N_11249,N_10235,N_10233);
xnor U11250 (N_11250,N_10250,N_10768);
nand U11251 (N_11251,N_10545,N_10725);
nor U11252 (N_11252,N_10392,N_10576);
and U11253 (N_11253,N_10433,N_10233);
nor U11254 (N_11254,N_10533,N_10571);
xor U11255 (N_11255,N_10562,N_10769);
or U11256 (N_11256,N_10681,N_10421);
or U11257 (N_11257,N_10613,N_10473);
or U11258 (N_11258,N_10201,N_10591);
and U11259 (N_11259,N_10623,N_10491);
nand U11260 (N_11260,N_10744,N_10562);
nand U11261 (N_11261,N_10395,N_10470);
nand U11262 (N_11262,N_10778,N_10659);
xnor U11263 (N_11263,N_10230,N_10622);
nand U11264 (N_11264,N_10738,N_10212);
nand U11265 (N_11265,N_10355,N_10413);
nand U11266 (N_11266,N_10418,N_10581);
nor U11267 (N_11267,N_10450,N_10507);
nand U11268 (N_11268,N_10446,N_10290);
xor U11269 (N_11269,N_10451,N_10301);
nand U11270 (N_11270,N_10206,N_10758);
or U11271 (N_11271,N_10675,N_10784);
nor U11272 (N_11272,N_10228,N_10567);
or U11273 (N_11273,N_10229,N_10200);
xor U11274 (N_11274,N_10279,N_10342);
or U11275 (N_11275,N_10473,N_10729);
nand U11276 (N_11276,N_10619,N_10657);
nor U11277 (N_11277,N_10206,N_10391);
and U11278 (N_11278,N_10452,N_10477);
and U11279 (N_11279,N_10294,N_10607);
and U11280 (N_11280,N_10569,N_10348);
and U11281 (N_11281,N_10672,N_10323);
nor U11282 (N_11282,N_10398,N_10713);
nor U11283 (N_11283,N_10381,N_10529);
nor U11284 (N_11284,N_10339,N_10212);
or U11285 (N_11285,N_10227,N_10669);
nand U11286 (N_11286,N_10228,N_10346);
nand U11287 (N_11287,N_10548,N_10200);
or U11288 (N_11288,N_10217,N_10302);
xnor U11289 (N_11289,N_10337,N_10629);
xor U11290 (N_11290,N_10748,N_10623);
and U11291 (N_11291,N_10611,N_10704);
and U11292 (N_11292,N_10622,N_10633);
nor U11293 (N_11293,N_10270,N_10409);
nand U11294 (N_11294,N_10356,N_10268);
or U11295 (N_11295,N_10231,N_10438);
nor U11296 (N_11296,N_10362,N_10757);
xor U11297 (N_11297,N_10762,N_10367);
xor U11298 (N_11298,N_10432,N_10481);
nor U11299 (N_11299,N_10776,N_10600);
nand U11300 (N_11300,N_10242,N_10533);
or U11301 (N_11301,N_10439,N_10653);
nand U11302 (N_11302,N_10743,N_10560);
xor U11303 (N_11303,N_10728,N_10201);
or U11304 (N_11304,N_10281,N_10451);
nor U11305 (N_11305,N_10283,N_10687);
nand U11306 (N_11306,N_10302,N_10202);
nand U11307 (N_11307,N_10747,N_10602);
and U11308 (N_11308,N_10622,N_10397);
nor U11309 (N_11309,N_10395,N_10672);
and U11310 (N_11310,N_10502,N_10467);
or U11311 (N_11311,N_10543,N_10442);
nor U11312 (N_11312,N_10477,N_10615);
nor U11313 (N_11313,N_10537,N_10654);
xnor U11314 (N_11314,N_10279,N_10280);
nor U11315 (N_11315,N_10539,N_10771);
or U11316 (N_11316,N_10234,N_10703);
nor U11317 (N_11317,N_10227,N_10460);
and U11318 (N_11318,N_10702,N_10799);
nand U11319 (N_11319,N_10672,N_10482);
xnor U11320 (N_11320,N_10369,N_10327);
and U11321 (N_11321,N_10780,N_10296);
and U11322 (N_11322,N_10495,N_10652);
or U11323 (N_11323,N_10443,N_10363);
xnor U11324 (N_11324,N_10409,N_10775);
and U11325 (N_11325,N_10524,N_10597);
nor U11326 (N_11326,N_10231,N_10607);
nand U11327 (N_11327,N_10684,N_10288);
and U11328 (N_11328,N_10211,N_10342);
or U11329 (N_11329,N_10420,N_10564);
nor U11330 (N_11330,N_10673,N_10209);
and U11331 (N_11331,N_10643,N_10323);
or U11332 (N_11332,N_10413,N_10741);
or U11333 (N_11333,N_10667,N_10777);
nor U11334 (N_11334,N_10282,N_10298);
xnor U11335 (N_11335,N_10529,N_10799);
xor U11336 (N_11336,N_10200,N_10499);
xnor U11337 (N_11337,N_10305,N_10373);
nor U11338 (N_11338,N_10617,N_10329);
xnor U11339 (N_11339,N_10701,N_10599);
xnor U11340 (N_11340,N_10715,N_10595);
nand U11341 (N_11341,N_10204,N_10762);
nand U11342 (N_11342,N_10492,N_10289);
xor U11343 (N_11343,N_10749,N_10329);
nand U11344 (N_11344,N_10333,N_10403);
nand U11345 (N_11345,N_10202,N_10732);
or U11346 (N_11346,N_10239,N_10300);
or U11347 (N_11347,N_10477,N_10482);
xnor U11348 (N_11348,N_10575,N_10345);
or U11349 (N_11349,N_10756,N_10344);
xor U11350 (N_11350,N_10592,N_10476);
and U11351 (N_11351,N_10493,N_10792);
nor U11352 (N_11352,N_10262,N_10460);
or U11353 (N_11353,N_10347,N_10274);
and U11354 (N_11354,N_10301,N_10629);
nor U11355 (N_11355,N_10266,N_10586);
xor U11356 (N_11356,N_10797,N_10383);
xor U11357 (N_11357,N_10297,N_10377);
xnor U11358 (N_11358,N_10317,N_10345);
xor U11359 (N_11359,N_10299,N_10236);
xnor U11360 (N_11360,N_10437,N_10358);
nand U11361 (N_11361,N_10403,N_10534);
nand U11362 (N_11362,N_10253,N_10433);
xor U11363 (N_11363,N_10218,N_10530);
or U11364 (N_11364,N_10536,N_10389);
or U11365 (N_11365,N_10226,N_10562);
nor U11366 (N_11366,N_10438,N_10230);
nand U11367 (N_11367,N_10745,N_10266);
or U11368 (N_11368,N_10493,N_10774);
nor U11369 (N_11369,N_10607,N_10282);
nand U11370 (N_11370,N_10246,N_10451);
nand U11371 (N_11371,N_10785,N_10254);
or U11372 (N_11372,N_10682,N_10339);
or U11373 (N_11373,N_10704,N_10788);
or U11374 (N_11374,N_10784,N_10553);
nor U11375 (N_11375,N_10749,N_10516);
nor U11376 (N_11376,N_10698,N_10553);
and U11377 (N_11377,N_10228,N_10380);
nor U11378 (N_11378,N_10571,N_10697);
nand U11379 (N_11379,N_10503,N_10455);
xor U11380 (N_11380,N_10701,N_10606);
and U11381 (N_11381,N_10559,N_10315);
or U11382 (N_11382,N_10274,N_10212);
or U11383 (N_11383,N_10620,N_10390);
and U11384 (N_11384,N_10257,N_10631);
and U11385 (N_11385,N_10458,N_10521);
and U11386 (N_11386,N_10798,N_10532);
or U11387 (N_11387,N_10308,N_10221);
xnor U11388 (N_11388,N_10451,N_10738);
nand U11389 (N_11389,N_10450,N_10421);
nor U11390 (N_11390,N_10548,N_10584);
and U11391 (N_11391,N_10553,N_10517);
nand U11392 (N_11392,N_10591,N_10476);
nand U11393 (N_11393,N_10756,N_10482);
xnor U11394 (N_11394,N_10510,N_10480);
nor U11395 (N_11395,N_10756,N_10620);
nand U11396 (N_11396,N_10207,N_10227);
nor U11397 (N_11397,N_10442,N_10507);
and U11398 (N_11398,N_10720,N_10527);
and U11399 (N_11399,N_10345,N_10283);
and U11400 (N_11400,N_10818,N_11160);
or U11401 (N_11401,N_11170,N_11175);
and U11402 (N_11402,N_10858,N_11308);
xor U11403 (N_11403,N_11314,N_11343);
nand U11404 (N_11404,N_11390,N_10868);
nand U11405 (N_11405,N_11145,N_10938);
and U11406 (N_11406,N_11178,N_11211);
and U11407 (N_11407,N_11080,N_11251);
and U11408 (N_11408,N_10966,N_11374);
xnor U11409 (N_11409,N_10974,N_11011);
xnor U11410 (N_11410,N_10863,N_11187);
or U11411 (N_11411,N_11033,N_11064);
xnor U11412 (N_11412,N_10809,N_11154);
and U11413 (N_11413,N_11017,N_10881);
xnor U11414 (N_11414,N_10888,N_11009);
xor U11415 (N_11415,N_10836,N_10939);
nand U11416 (N_11416,N_10835,N_10906);
or U11417 (N_11417,N_11373,N_11140);
and U11418 (N_11418,N_11347,N_10903);
nor U11419 (N_11419,N_11333,N_11079);
or U11420 (N_11420,N_10909,N_10821);
nand U11421 (N_11421,N_11227,N_11172);
or U11422 (N_11422,N_11038,N_10981);
nor U11423 (N_11423,N_11281,N_10896);
nand U11424 (N_11424,N_11209,N_10986);
or U11425 (N_11425,N_11327,N_10875);
and U11426 (N_11426,N_11032,N_10829);
nor U11427 (N_11427,N_11118,N_11087);
xor U11428 (N_11428,N_10982,N_11036);
nor U11429 (N_11429,N_11357,N_10990);
and U11430 (N_11430,N_11286,N_11103);
and U11431 (N_11431,N_11122,N_10940);
nor U11432 (N_11432,N_11385,N_11290);
xor U11433 (N_11433,N_11034,N_10915);
or U11434 (N_11434,N_11142,N_11173);
nand U11435 (N_11435,N_10843,N_11271);
xor U11436 (N_11436,N_10877,N_11295);
or U11437 (N_11437,N_10947,N_11367);
or U11438 (N_11438,N_11049,N_10894);
and U11439 (N_11439,N_11188,N_11361);
and U11440 (N_11440,N_11375,N_11312);
nand U11441 (N_11441,N_11383,N_11394);
or U11442 (N_11442,N_10871,N_11307);
and U11443 (N_11443,N_10866,N_10907);
or U11444 (N_11444,N_10804,N_11255);
nor U11445 (N_11445,N_11092,N_11129);
nor U11446 (N_11446,N_10897,N_10997);
nor U11447 (N_11447,N_11042,N_11245);
xor U11448 (N_11448,N_10993,N_10834);
or U11449 (N_11449,N_11197,N_10910);
xor U11450 (N_11450,N_11063,N_10820);
and U11451 (N_11451,N_10919,N_11168);
nand U11452 (N_11452,N_10950,N_11313);
and U11453 (N_11453,N_11039,N_11167);
nand U11454 (N_11454,N_11370,N_11297);
nor U11455 (N_11455,N_10912,N_10878);
nor U11456 (N_11456,N_10840,N_11289);
xor U11457 (N_11457,N_11349,N_11005);
nand U11458 (N_11458,N_11330,N_10850);
or U11459 (N_11459,N_11382,N_11350);
or U11460 (N_11460,N_11056,N_11391);
and U11461 (N_11461,N_11176,N_10864);
nand U11462 (N_11462,N_11166,N_10819);
nor U11463 (N_11463,N_10892,N_10839);
or U11464 (N_11464,N_11224,N_11083);
or U11465 (N_11465,N_11284,N_11228);
nand U11466 (N_11466,N_11257,N_11134);
xor U11467 (N_11467,N_11318,N_11196);
nor U11468 (N_11468,N_11287,N_11293);
and U11469 (N_11469,N_11029,N_11316);
nand U11470 (N_11470,N_11086,N_10830);
nor U11471 (N_11471,N_10833,N_10854);
nor U11472 (N_11472,N_11202,N_11301);
xor U11473 (N_11473,N_11315,N_10806);
nor U11474 (N_11474,N_10817,N_11192);
nor U11475 (N_11475,N_11095,N_10926);
xnor U11476 (N_11476,N_11232,N_11085);
and U11477 (N_11477,N_10846,N_11244);
xnor U11478 (N_11478,N_11008,N_11282);
or U11479 (N_11479,N_11221,N_11354);
or U11480 (N_11480,N_10998,N_11112);
xor U11481 (N_11481,N_11276,N_10802);
or U11482 (N_11482,N_11148,N_11078);
and U11483 (N_11483,N_11003,N_11352);
xor U11484 (N_11484,N_11236,N_10822);
or U11485 (N_11485,N_10923,N_11132);
nand U11486 (N_11486,N_11046,N_11096);
or U11487 (N_11487,N_10949,N_10925);
and U11488 (N_11488,N_11061,N_11066);
nand U11489 (N_11489,N_11323,N_11261);
and U11490 (N_11490,N_11194,N_11351);
nor U11491 (N_11491,N_11217,N_11065);
nor U11492 (N_11492,N_11212,N_11262);
xor U11493 (N_11493,N_11143,N_11163);
or U11494 (N_11494,N_10955,N_11097);
and U11495 (N_11495,N_11067,N_10898);
nor U11496 (N_11496,N_10911,N_10967);
xnor U11497 (N_11497,N_10985,N_11291);
xnor U11498 (N_11498,N_11213,N_11107);
nor U11499 (N_11499,N_11277,N_11119);
nand U11500 (N_11500,N_11075,N_10831);
or U11501 (N_11501,N_10913,N_10825);
nand U11502 (N_11502,N_10952,N_11060);
xnor U11503 (N_11503,N_10893,N_11157);
xor U11504 (N_11504,N_10922,N_11115);
nor U11505 (N_11505,N_11283,N_11309);
and U11506 (N_11506,N_11372,N_11052);
or U11507 (N_11507,N_11089,N_11210);
nand U11508 (N_11508,N_10953,N_11111);
nand U11509 (N_11509,N_10928,N_11376);
nand U11510 (N_11510,N_11044,N_10989);
nor U11511 (N_11511,N_10828,N_11048);
nand U11512 (N_11512,N_11246,N_10921);
xor U11513 (N_11513,N_10951,N_11346);
nand U11514 (N_11514,N_11072,N_11189);
nor U11515 (N_11515,N_11105,N_10874);
or U11516 (N_11516,N_11389,N_11356);
nand U11517 (N_11517,N_11090,N_11322);
and U11518 (N_11518,N_11340,N_10927);
nor U11519 (N_11519,N_11319,N_11031);
and U11520 (N_11520,N_10957,N_11137);
or U11521 (N_11521,N_11128,N_11222);
nand U11522 (N_11522,N_11300,N_11071);
nand U11523 (N_11523,N_10869,N_11264);
and U11524 (N_11524,N_11151,N_11205);
xor U11525 (N_11525,N_10841,N_11139);
nor U11526 (N_11526,N_11216,N_11328);
nand U11527 (N_11527,N_11133,N_11303);
xnor U11528 (N_11528,N_10931,N_10815);
nor U11529 (N_11529,N_11358,N_10900);
or U11530 (N_11530,N_10899,N_10977);
xor U11531 (N_11531,N_11062,N_11219);
nor U11532 (N_11532,N_10917,N_11325);
and U11533 (N_11533,N_10852,N_11237);
xnor U11534 (N_11534,N_10976,N_11004);
or U11535 (N_11535,N_10845,N_11195);
or U11536 (N_11536,N_10860,N_11165);
and U11537 (N_11537,N_11368,N_11113);
nor U11538 (N_11538,N_11344,N_10849);
nand U11539 (N_11539,N_11225,N_11399);
xor U11540 (N_11540,N_11100,N_10884);
xnor U11541 (N_11541,N_11338,N_10891);
nor U11542 (N_11542,N_11392,N_10969);
or U11543 (N_11543,N_10961,N_10945);
nor U11544 (N_11544,N_10859,N_11233);
xnor U11545 (N_11545,N_11028,N_11256);
nor U11546 (N_11546,N_11109,N_10879);
nor U11547 (N_11547,N_11135,N_11158);
or U11548 (N_11548,N_11020,N_11114);
xor U11549 (N_11549,N_10811,N_11248);
nor U11550 (N_11550,N_10870,N_11006);
nand U11551 (N_11551,N_11305,N_11288);
nand U11552 (N_11552,N_11377,N_11126);
or U11553 (N_11553,N_11339,N_10942);
and U11554 (N_11554,N_11332,N_11279);
or U11555 (N_11555,N_11334,N_10873);
xor U11556 (N_11556,N_11002,N_11050);
nand U11557 (N_11557,N_10812,N_11164);
and U11558 (N_11558,N_11384,N_10880);
nand U11559 (N_11559,N_11018,N_11070);
and U11560 (N_11560,N_11169,N_11059);
or U11561 (N_11561,N_11296,N_11342);
xor U11562 (N_11562,N_11030,N_11182);
and U11563 (N_11563,N_10803,N_10968);
nand U11564 (N_11564,N_10895,N_11191);
xor U11565 (N_11565,N_11231,N_11155);
and U11566 (N_11566,N_11241,N_11088);
and U11567 (N_11567,N_11058,N_11311);
nand U11568 (N_11568,N_11206,N_11269);
or U11569 (N_11569,N_11335,N_10960);
xnor U11570 (N_11570,N_10837,N_11180);
and U11571 (N_11571,N_11381,N_11320);
xnor U11572 (N_11572,N_11144,N_10994);
or U11573 (N_11573,N_11324,N_11161);
nor U11574 (N_11574,N_10827,N_11068);
and U11575 (N_11575,N_11185,N_11117);
nor U11576 (N_11576,N_11130,N_10962);
nor U11577 (N_11577,N_11215,N_11190);
or U11578 (N_11578,N_11304,N_10887);
or U11579 (N_11579,N_11380,N_10935);
nand U11580 (N_11580,N_11016,N_10980);
or U11581 (N_11581,N_11146,N_10885);
or U11582 (N_11582,N_11278,N_11076);
nor U11583 (N_11583,N_11024,N_10901);
and U11584 (N_11584,N_11014,N_10999);
nor U11585 (N_11585,N_10857,N_11104);
and U11586 (N_11586,N_10978,N_11198);
and U11587 (N_11587,N_11243,N_11345);
xnor U11588 (N_11588,N_10958,N_10936);
nor U11589 (N_11589,N_11027,N_11055);
nand U11590 (N_11590,N_11041,N_11274);
nand U11591 (N_11591,N_10838,N_10832);
and U11592 (N_11592,N_11127,N_11378);
nand U11593 (N_11593,N_11084,N_11081);
and U11594 (N_11594,N_11331,N_11116);
or U11595 (N_11595,N_11341,N_11159);
nand U11596 (N_11596,N_11193,N_11379);
and U11597 (N_11597,N_10855,N_11238);
or U11598 (N_11598,N_11201,N_10972);
or U11599 (N_11599,N_11292,N_11214);
nor U11600 (N_11600,N_10941,N_11102);
or U11601 (N_11601,N_11149,N_11294);
nor U11602 (N_11602,N_11247,N_11268);
and U11603 (N_11603,N_11397,N_11153);
nor U11604 (N_11604,N_11037,N_10975);
nor U11605 (N_11605,N_10933,N_11199);
xor U11606 (N_11606,N_11120,N_10971);
nand U11607 (N_11607,N_11235,N_11125);
or U11608 (N_11608,N_10853,N_10883);
or U11609 (N_11609,N_11051,N_11147);
nor U11610 (N_11610,N_11364,N_10956);
and U11611 (N_11611,N_11043,N_11174);
or U11612 (N_11612,N_10805,N_10861);
or U11613 (N_11613,N_10916,N_11093);
xnor U11614 (N_11614,N_11138,N_10842);
nor U11615 (N_11615,N_10867,N_10929);
nand U11616 (N_11616,N_11074,N_11353);
xor U11617 (N_11617,N_11156,N_10808);
xnor U11618 (N_11618,N_10800,N_10844);
xnor U11619 (N_11619,N_11280,N_11208);
nor U11620 (N_11620,N_11181,N_11259);
nand U11621 (N_11621,N_10991,N_11365);
and U11622 (N_11622,N_10959,N_11183);
nand U11623 (N_11623,N_11150,N_11249);
or U11624 (N_11624,N_10816,N_10904);
xor U11625 (N_11625,N_11393,N_11023);
or U11626 (N_11626,N_11371,N_10872);
and U11627 (N_11627,N_11220,N_11203);
or U11628 (N_11628,N_11310,N_10865);
or U11629 (N_11629,N_11360,N_11223);
xnor U11630 (N_11630,N_11329,N_11131);
nor U11631 (N_11631,N_10946,N_11053);
and U11632 (N_11632,N_11123,N_11226);
or U11633 (N_11633,N_11298,N_10914);
xnor U11634 (N_11634,N_11021,N_11326);
nor U11635 (N_11635,N_11204,N_10813);
nor U11636 (N_11636,N_11270,N_10847);
or U11637 (N_11637,N_11252,N_10807);
and U11638 (N_11638,N_11045,N_11040);
and U11639 (N_11639,N_10924,N_11250);
nor U11640 (N_11640,N_11124,N_11101);
nor U11641 (N_11641,N_11366,N_11054);
xnor U11642 (N_11642,N_11362,N_11355);
and U11643 (N_11643,N_10973,N_11395);
or U11644 (N_11644,N_11207,N_11110);
or U11645 (N_11645,N_11077,N_10992);
and U11646 (N_11646,N_11302,N_11082);
xnor U11647 (N_11647,N_10905,N_10902);
nand U11648 (N_11648,N_11108,N_10930);
or U11649 (N_11649,N_11121,N_11069);
or U11650 (N_11650,N_10983,N_11022);
nor U11651 (N_11651,N_11386,N_11398);
xnor U11652 (N_11652,N_11171,N_11057);
nor U11653 (N_11653,N_11010,N_10944);
nand U11654 (N_11654,N_10882,N_10848);
and U11655 (N_11655,N_10890,N_11336);
xor U11656 (N_11656,N_11007,N_10943);
nor U11657 (N_11657,N_10954,N_11177);
xor U11658 (N_11658,N_10876,N_11200);
nand U11659 (N_11659,N_11000,N_11019);
nand U11660 (N_11660,N_11267,N_11186);
nor U11661 (N_11661,N_10801,N_11015);
xnor U11662 (N_11662,N_11136,N_11317);
xor U11663 (N_11663,N_10814,N_10826);
nor U11664 (N_11664,N_10823,N_11234);
nor U11665 (N_11665,N_11073,N_10862);
xor U11666 (N_11666,N_10984,N_10908);
and U11667 (N_11667,N_11242,N_11275);
nor U11668 (N_11668,N_10824,N_11162);
xor U11669 (N_11669,N_10934,N_11263);
nor U11670 (N_11670,N_10979,N_11285);
nand U11671 (N_11671,N_10988,N_11012);
xnor U11672 (N_11672,N_11240,N_10995);
xor U11673 (N_11673,N_11091,N_11260);
nand U11674 (N_11674,N_11230,N_10920);
nor U11675 (N_11675,N_11359,N_11369);
nor U11676 (N_11676,N_10918,N_11179);
xor U11677 (N_11677,N_11026,N_11348);
xor U11678 (N_11678,N_11001,N_11025);
nand U11679 (N_11679,N_10932,N_11098);
and U11680 (N_11680,N_10996,N_11099);
and U11681 (N_11681,N_11306,N_11035);
xnor U11682 (N_11682,N_11047,N_10948);
xnor U11683 (N_11683,N_11321,N_10963);
nor U11684 (N_11684,N_11272,N_11094);
xnor U11685 (N_11685,N_11265,N_11337);
or U11686 (N_11686,N_11184,N_10964);
xor U11687 (N_11687,N_11273,N_10987);
or U11688 (N_11688,N_11299,N_11387);
and U11689 (N_11689,N_10889,N_10886);
nand U11690 (N_11690,N_11363,N_11396);
and U11691 (N_11691,N_11106,N_11253);
xnor U11692 (N_11692,N_10851,N_11254);
xnor U11693 (N_11693,N_10937,N_10965);
or U11694 (N_11694,N_10810,N_11258);
or U11695 (N_11695,N_11013,N_11141);
or U11696 (N_11696,N_10856,N_11152);
and U11697 (N_11697,N_11388,N_11229);
nor U11698 (N_11698,N_11239,N_10970);
xor U11699 (N_11699,N_11218,N_11266);
nand U11700 (N_11700,N_10981,N_11186);
xor U11701 (N_11701,N_11154,N_11136);
nor U11702 (N_11702,N_11396,N_11171);
xnor U11703 (N_11703,N_11244,N_10956);
nor U11704 (N_11704,N_10915,N_11067);
or U11705 (N_11705,N_11045,N_11115);
xor U11706 (N_11706,N_10813,N_11071);
and U11707 (N_11707,N_11327,N_10800);
or U11708 (N_11708,N_11012,N_11013);
nor U11709 (N_11709,N_11050,N_10933);
and U11710 (N_11710,N_10836,N_10849);
xnor U11711 (N_11711,N_10969,N_11174);
xnor U11712 (N_11712,N_10924,N_10899);
or U11713 (N_11713,N_11064,N_10982);
nand U11714 (N_11714,N_11315,N_11053);
nand U11715 (N_11715,N_10950,N_11355);
xnor U11716 (N_11716,N_10893,N_11195);
xor U11717 (N_11717,N_11176,N_11031);
nor U11718 (N_11718,N_10921,N_11062);
and U11719 (N_11719,N_10926,N_10871);
or U11720 (N_11720,N_11206,N_11385);
xnor U11721 (N_11721,N_10935,N_11255);
xnor U11722 (N_11722,N_11279,N_11238);
and U11723 (N_11723,N_11344,N_10882);
or U11724 (N_11724,N_11217,N_11120);
or U11725 (N_11725,N_10985,N_11072);
xor U11726 (N_11726,N_11009,N_11371);
xnor U11727 (N_11727,N_10986,N_10894);
nor U11728 (N_11728,N_11320,N_10835);
or U11729 (N_11729,N_11184,N_10959);
nand U11730 (N_11730,N_11239,N_10814);
nor U11731 (N_11731,N_11003,N_10858);
nand U11732 (N_11732,N_11175,N_11187);
xor U11733 (N_11733,N_10814,N_11270);
or U11734 (N_11734,N_11216,N_10932);
nor U11735 (N_11735,N_11068,N_10900);
xor U11736 (N_11736,N_11141,N_10814);
xor U11737 (N_11737,N_11344,N_11281);
nand U11738 (N_11738,N_11381,N_10912);
nand U11739 (N_11739,N_10848,N_11009);
nand U11740 (N_11740,N_11166,N_11191);
and U11741 (N_11741,N_10859,N_10840);
xnor U11742 (N_11742,N_10808,N_11307);
xnor U11743 (N_11743,N_11319,N_10805);
nor U11744 (N_11744,N_10947,N_10859);
or U11745 (N_11745,N_10820,N_10960);
or U11746 (N_11746,N_11353,N_11159);
or U11747 (N_11747,N_11390,N_11054);
nand U11748 (N_11748,N_11372,N_11253);
or U11749 (N_11749,N_11263,N_10906);
nor U11750 (N_11750,N_11383,N_11075);
nor U11751 (N_11751,N_11240,N_10906);
nor U11752 (N_11752,N_10911,N_11203);
nor U11753 (N_11753,N_11257,N_10911);
xnor U11754 (N_11754,N_11378,N_11019);
or U11755 (N_11755,N_10851,N_10828);
xor U11756 (N_11756,N_11339,N_11074);
nor U11757 (N_11757,N_11048,N_11246);
or U11758 (N_11758,N_11008,N_10835);
xnor U11759 (N_11759,N_11312,N_10927);
nand U11760 (N_11760,N_11246,N_11336);
xor U11761 (N_11761,N_11066,N_11324);
nand U11762 (N_11762,N_11051,N_10881);
xor U11763 (N_11763,N_10909,N_11121);
and U11764 (N_11764,N_11127,N_11121);
nor U11765 (N_11765,N_11346,N_10996);
nand U11766 (N_11766,N_11233,N_11385);
xnor U11767 (N_11767,N_11291,N_11044);
and U11768 (N_11768,N_11010,N_11096);
and U11769 (N_11769,N_11338,N_11089);
and U11770 (N_11770,N_11186,N_11098);
nand U11771 (N_11771,N_11351,N_11134);
nand U11772 (N_11772,N_10852,N_10989);
or U11773 (N_11773,N_11175,N_11096);
xor U11774 (N_11774,N_11314,N_11268);
nand U11775 (N_11775,N_11347,N_10890);
nand U11776 (N_11776,N_11046,N_11390);
xor U11777 (N_11777,N_11236,N_11359);
and U11778 (N_11778,N_10977,N_11184);
nor U11779 (N_11779,N_11393,N_10923);
and U11780 (N_11780,N_11276,N_11250);
xnor U11781 (N_11781,N_10804,N_11233);
nor U11782 (N_11782,N_10875,N_10842);
nor U11783 (N_11783,N_11143,N_11273);
xnor U11784 (N_11784,N_11202,N_11005);
or U11785 (N_11785,N_10998,N_11392);
xnor U11786 (N_11786,N_10998,N_11379);
or U11787 (N_11787,N_11264,N_10940);
xor U11788 (N_11788,N_10978,N_11361);
xor U11789 (N_11789,N_11043,N_11222);
nand U11790 (N_11790,N_10921,N_10811);
nand U11791 (N_11791,N_10969,N_11034);
and U11792 (N_11792,N_11180,N_11391);
or U11793 (N_11793,N_11389,N_11068);
nand U11794 (N_11794,N_11283,N_11247);
nor U11795 (N_11795,N_10869,N_10881);
or U11796 (N_11796,N_11242,N_11328);
nor U11797 (N_11797,N_10955,N_11189);
xnor U11798 (N_11798,N_11143,N_11042);
and U11799 (N_11799,N_11037,N_11066);
nor U11800 (N_11800,N_11377,N_11390);
nor U11801 (N_11801,N_11386,N_11381);
and U11802 (N_11802,N_11026,N_11111);
or U11803 (N_11803,N_10934,N_11318);
xor U11804 (N_11804,N_11295,N_10931);
nor U11805 (N_11805,N_10912,N_11266);
nor U11806 (N_11806,N_10998,N_10969);
or U11807 (N_11807,N_10947,N_11106);
and U11808 (N_11808,N_10965,N_11312);
and U11809 (N_11809,N_11050,N_11028);
or U11810 (N_11810,N_10895,N_11216);
or U11811 (N_11811,N_11148,N_10805);
xnor U11812 (N_11812,N_11354,N_11012);
and U11813 (N_11813,N_11059,N_11139);
and U11814 (N_11814,N_11369,N_11378);
or U11815 (N_11815,N_10866,N_10898);
and U11816 (N_11816,N_11127,N_11115);
and U11817 (N_11817,N_11397,N_11308);
xor U11818 (N_11818,N_10916,N_10887);
nor U11819 (N_11819,N_10822,N_11246);
nor U11820 (N_11820,N_11020,N_11211);
xor U11821 (N_11821,N_10980,N_11356);
or U11822 (N_11822,N_10963,N_11302);
or U11823 (N_11823,N_11239,N_10957);
nor U11824 (N_11824,N_11076,N_11061);
xor U11825 (N_11825,N_11144,N_11159);
nand U11826 (N_11826,N_11070,N_11060);
nand U11827 (N_11827,N_11196,N_11035);
nor U11828 (N_11828,N_11391,N_10921);
xnor U11829 (N_11829,N_11398,N_11371);
nor U11830 (N_11830,N_10854,N_11322);
and U11831 (N_11831,N_10961,N_11169);
nor U11832 (N_11832,N_11116,N_11100);
nor U11833 (N_11833,N_11002,N_11064);
nor U11834 (N_11834,N_11026,N_10800);
nand U11835 (N_11835,N_11312,N_11284);
xor U11836 (N_11836,N_11390,N_11283);
nor U11837 (N_11837,N_11097,N_11214);
and U11838 (N_11838,N_10978,N_11312);
xnor U11839 (N_11839,N_11078,N_11311);
and U11840 (N_11840,N_11366,N_11337);
nor U11841 (N_11841,N_11159,N_11265);
and U11842 (N_11842,N_11276,N_11068);
nand U11843 (N_11843,N_10988,N_11148);
xor U11844 (N_11844,N_10855,N_11391);
and U11845 (N_11845,N_11147,N_11354);
or U11846 (N_11846,N_11340,N_11156);
nand U11847 (N_11847,N_11070,N_11206);
xor U11848 (N_11848,N_11004,N_11133);
nor U11849 (N_11849,N_11240,N_11368);
and U11850 (N_11850,N_10940,N_11035);
nor U11851 (N_11851,N_11299,N_10938);
xor U11852 (N_11852,N_10914,N_11212);
nor U11853 (N_11853,N_10860,N_11267);
xnor U11854 (N_11854,N_11100,N_11200);
nand U11855 (N_11855,N_10943,N_10937);
and U11856 (N_11856,N_10996,N_11328);
or U11857 (N_11857,N_11332,N_11340);
and U11858 (N_11858,N_11213,N_10981);
or U11859 (N_11859,N_10876,N_11279);
nor U11860 (N_11860,N_11269,N_11239);
and U11861 (N_11861,N_11042,N_11292);
xnor U11862 (N_11862,N_10895,N_11274);
nand U11863 (N_11863,N_11250,N_11121);
nor U11864 (N_11864,N_11250,N_10813);
and U11865 (N_11865,N_10940,N_10828);
nand U11866 (N_11866,N_11052,N_11038);
nor U11867 (N_11867,N_10833,N_10999);
or U11868 (N_11868,N_11397,N_11181);
nand U11869 (N_11869,N_10823,N_11193);
or U11870 (N_11870,N_10949,N_11020);
and U11871 (N_11871,N_11303,N_11135);
or U11872 (N_11872,N_10854,N_11261);
nand U11873 (N_11873,N_11037,N_11322);
or U11874 (N_11874,N_11297,N_11258);
nor U11875 (N_11875,N_11106,N_10908);
or U11876 (N_11876,N_11287,N_11005);
or U11877 (N_11877,N_10931,N_11191);
and U11878 (N_11878,N_11233,N_10964);
or U11879 (N_11879,N_11314,N_11397);
or U11880 (N_11880,N_11033,N_11186);
nor U11881 (N_11881,N_11194,N_11255);
nand U11882 (N_11882,N_10813,N_11221);
nor U11883 (N_11883,N_10966,N_10866);
nand U11884 (N_11884,N_11233,N_10950);
and U11885 (N_11885,N_11000,N_10845);
nor U11886 (N_11886,N_11225,N_11289);
nand U11887 (N_11887,N_11236,N_10848);
and U11888 (N_11888,N_10943,N_11277);
or U11889 (N_11889,N_11388,N_10955);
xor U11890 (N_11890,N_11118,N_10950);
or U11891 (N_11891,N_11174,N_11350);
and U11892 (N_11892,N_10822,N_10839);
xor U11893 (N_11893,N_11050,N_11285);
or U11894 (N_11894,N_10999,N_11338);
or U11895 (N_11895,N_11225,N_11246);
or U11896 (N_11896,N_11046,N_10910);
and U11897 (N_11897,N_10907,N_11366);
nor U11898 (N_11898,N_10958,N_10814);
or U11899 (N_11899,N_11128,N_11151);
or U11900 (N_11900,N_10994,N_10884);
nand U11901 (N_11901,N_11330,N_10901);
nor U11902 (N_11902,N_10875,N_11096);
nand U11903 (N_11903,N_10873,N_11391);
xor U11904 (N_11904,N_10948,N_11085);
nor U11905 (N_11905,N_11261,N_10941);
and U11906 (N_11906,N_11320,N_11074);
xor U11907 (N_11907,N_11021,N_10887);
or U11908 (N_11908,N_10855,N_11369);
nand U11909 (N_11909,N_11374,N_10810);
xor U11910 (N_11910,N_10851,N_11172);
nand U11911 (N_11911,N_10907,N_10956);
nand U11912 (N_11912,N_11337,N_10879);
nor U11913 (N_11913,N_11159,N_10856);
xor U11914 (N_11914,N_11286,N_10921);
nor U11915 (N_11915,N_11226,N_11262);
or U11916 (N_11916,N_11184,N_11068);
nor U11917 (N_11917,N_11393,N_10998);
xnor U11918 (N_11918,N_10820,N_11218);
xnor U11919 (N_11919,N_11022,N_10956);
or U11920 (N_11920,N_10933,N_11346);
and U11921 (N_11921,N_10804,N_11043);
nand U11922 (N_11922,N_10966,N_11126);
nor U11923 (N_11923,N_11301,N_11091);
xor U11924 (N_11924,N_11219,N_10954);
xnor U11925 (N_11925,N_10904,N_10981);
nor U11926 (N_11926,N_10996,N_11189);
or U11927 (N_11927,N_11050,N_10914);
or U11928 (N_11928,N_10877,N_11112);
nand U11929 (N_11929,N_10861,N_10895);
nor U11930 (N_11930,N_11035,N_10903);
nand U11931 (N_11931,N_11216,N_10863);
xor U11932 (N_11932,N_11285,N_11310);
xnor U11933 (N_11933,N_11007,N_10802);
or U11934 (N_11934,N_11127,N_10901);
or U11935 (N_11935,N_11061,N_11108);
xor U11936 (N_11936,N_10863,N_11314);
or U11937 (N_11937,N_10933,N_11242);
nand U11938 (N_11938,N_11272,N_11348);
nor U11939 (N_11939,N_11042,N_11302);
nor U11940 (N_11940,N_11130,N_11191);
nor U11941 (N_11941,N_11101,N_11266);
xor U11942 (N_11942,N_11328,N_11383);
or U11943 (N_11943,N_11048,N_11241);
xnor U11944 (N_11944,N_10897,N_10991);
or U11945 (N_11945,N_11271,N_11215);
or U11946 (N_11946,N_11300,N_11137);
xor U11947 (N_11947,N_11244,N_11182);
nor U11948 (N_11948,N_11278,N_11137);
and U11949 (N_11949,N_11132,N_11321);
and U11950 (N_11950,N_11196,N_11301);
nand U11951 (N_11951,N_11038,N_10832);
xor U11952 (N_11952,N_11001,N_11252);
nor U11953 (N_11953,N_10862,N_11360);
or U11954 (N_11954,N_11204,N_11034);
and U11955 (N_11955,N_11032,N_11054);
nor U11956 (N_11956,N_11302,N_11333);
nor U11957 (N_11957,N_11054,N_11289);
nor U11958 (N_11958,N_11252,N_11297);
or U11959 (N_11959,N_10969,N_11036);
nand U11960 (N_11960,N_11156,N_10854);
and U11961 (N_11961,N_11179,N_11066);
and U11962 (N_11962,N_11272,N_11064);
nand U11963 (N_11963,N_11024,N_11278);
xor U11964 (N_11964,N_10810,N_11247);
and U11965 (N_11965,N_11187,N_11272);
nor U11966 (N_11966,N_11272,N_11246);
nor U11967 (N_11967,N_11072,N_10856);
and U11968 (N_11968,N_11069,N_11160);
or U11969 (N_11969,N_11081,N_11383);
nor U11970 (N_11970,N_11020,N_11335);
xor U11971 (N_11971,N_11356,N_11323);
xnor U11972 (N_11972,N_11008,N_11348);
or U11973 (N_11973,N_11377,N_11205);
nor U11974 (N_11974,N_11284,N_11250);
nand U11975 (N_11975,N_10842,N_11154);
nand U11976 (N_11976,N_11383,N_11094);
or U11977 (N_11977,N_10811,N_10833);
or U11978 (N_11978,N_10995,N_11388);
and U11979 (N_11979,N_10934,N_10846);
or U11980 (N_11980,N_11093,N_11392);
nor U11981 (N_11981,N_11314,N_11310);
nand U11982 (N_11982,N_10865,N_11002);
or U11983 (N_11983,N_11042,N_10976);
or U11984 (N_11984,N_11143,N_11360);
and U11985 (N_11985,N_10986,N_11030);
nand U11986 (N_11986,N_11070,N_11323);
xor U11987 (N_11987,N_10959,N_10932);
and U11988 (N_11988,N_11323,N_11104);
nor U11989 (N_11989,N_11397,N_11273);
and U11990 (N_11990,N_10802,N_11177);
or U11991 (N_11991,N_10904,N_11027);
xnor U11992 (N_11992,N_11006,N_10996);
nor U11993 (N_11993,N_11066,N_11088);
nor U11994 (N_11994,N_11208,N_10835);
nor U11995 (N_11995,N_10883,N_10937);
xnor U11996 (N_11996,N_11280,N_11185);
xnor U11997 (N_11997,N_11253,N_10945);
nor U11998 (N_11998,N_11312,N_10888);
nand U11999 (N_11999,N_11175,N_10935);
nand U12000 (N_12000,N_11908,N_11711);
or U12001 (N_12001,N_11572,N_11527);
nand U12002 (N_12002,N_11708,N_11904);
nor U12003 (N_12003,N_11858,N_11604);
nor U12004 (N_12004,N_11629,N_11437);
or U12005 (N_12005,N_11988,N_11412);
nand U12006 (N_12006,N_11656,N_11570);
and U12007 (N_12007,N_11466,N_11718);
or U12008 (N_12008,N_11468,N_11712);
nor U12009 (N_12009,N_11594,N_11431);
nor U12010 (N_12010,N_11804,N_11725);
nand U12011 (N_12011,N_11498,N_11567);
xnor U12012 (N_12012,N_11770,N_11910);
nand U12013 (N_12013,N_11701,N_11839);
nand U12014 (N_12014,N_11899,N_11669);
xnor U12015 (N_12015,N_11496,N_11798);
xor U12016 (N_12016,N_11430,N_11873);
nand U12017 (N_12017,N_11891,N_11447);
or U12018 (N_12018,N_11513,N_11483);
and U12019 (N_12019,N_11451,N_11813);
or U12020 (N_12020,N_11864,N_11994);
xnor U12021 (N_12021,N_11687,N_11933);
nor U12022 (N_12022,N_11485,N_11550);
nand U12023 (N_12023,N_11674,N_11805);
xor U12024 (N_12024,N_11928,N_11775);
nand U12025 (N_12025,N_11519,N_11759);
xor U12026 (N_12026,N_11621,N_11965);
nor U12027 (N_12027,N_11489,N_11683);
xnor U12028 (N_12028,N_11408,N_11426);
or U12029 (N_12029,N_11405,N_11411);
xnor U12030 (N_12030,N_11709,N_11760);
nand U12031 (N_12031,N_11542,N_11727);
nand U12032 (N_12032,N_11852,N_11884);
or U12033 (N_12033,N_11860,N_11638);
and U12034 (N_12034,N_11942,N_11750);
and U12035 (N_12035,N_11761,N_11639);
or U12036 (N_12036,N_11467,N_11738);
and U12037 (N_12037,N_11609,N_11866);
and U12038 (N_12038,N_11953,N_11577);
nand U12039 (N_12039,N_11991,N_11957);
nand U12040 (N_12040,N_11603,N_11934);
and U12041 (N_12041,N_11459,N_11917);
xor U12042 (N_12042,N_11778,N_11903);
and U12043 (N_12043,N_11777,N_11555);
and U12044 (N_12044,N_11890,N_11861);
nor U12045 (N_12045,N_11710,N_11837);
xnor U12046 (N_12046,N_11673,N_11438);
nor U12047 (N_12047,N_11829,N_11754);
xor U12048 (N_12048,N_11600,N_11435);
and U12049 (N_12049,N_11509,N_11532);
and U12050 (N_12050,N_11416,N_11882);
xor U12051 (N_12051,N_11569,N_11992);
nor U12052 (N_12052,N_11444,N_11493);
xnor U12053 (N_12053,N_11644,N_11900);
nor U12054 (N_12054,N_11661,N_11596);
or U12055 (N_12055,N_11633,N_11460);
and U12056 (N_12056,N_11767,N_11529);
or U12057 (N_12057,N_11658,N_11838);
xnor U12058 (N_12058,N_11453,N_11476);
nand U12059 (N_12059,N_11440,N_11537);
or U12060 (N_12060,N_11722,N_11625);
nand U12061 (N_12061,N_11848,N_11528);
nand U12062 (N_12062,N_11840,N_11828);
xnor U12063 (N_12063,N_11671,N_11901);
nand U12064 (N_12064,N_11441,N_11788);
xor U12065 (N_12065,N_11794,N_11772);
or U12066 (N_12066,N_11583,N_11993);
or U12067 (N_12067,N_11650,N_11574);
and U12068 (N_12068,N_11739,N_11575);
nand U12069 (N_12069,N_11931,N_11691);
nand U12070 (N_12070,N_11472,N_11700);
and U12071 (N_12071,N_11636,N_11565);
xnor U12072 (N_12072,N_11892,N_11606);
nand U12073 (N_12073,N_11497,N_11886);
and U12074 (N_12074,N_11870,N_11659);
or U12075 (N_12075,N_11960,N_11543);
and U12076 (N_12076,N_11921,N_11424);
nor U12077 (N_12077,N_11803,N_11611);
or U12078 (N_12078,N_11915,N_11959);
xnor U12079 (N_12079,N_11789,N_11961);
nor U12080 (N_12080,N_11998,N_11679);
xor U12081 (N_12081,N_11952,N_11896);
nand U12082 (N_12082,N_11932,N_11702);
nor U12083 (N_12083,N_11927,N_11446);
nand U12084 (N_12084,N_11913,N_11732);
nand U12085 (N_12085,N_11449,N_11587);
or U12086 (N_12086,N_11560,N_11844);
nor U12087 (N_12087,N_11589,N_11597);
xnor U12088 (N_12088,N_11799,N_11598);
nor U12089 (N_12089,N_11938,N_11480);
xor U12090 (N_12090,N_11943,N_11949);
or U12091 (N_12091,N_11919,N_11699);
or U12092 (N_12092,N_11554,N_11643);
nand U12093 (N_12093,N_11403,N_11514);
nand U12094 (N_12094,N_11568,N_11746);
and U12095 (N_12095,N_11432,N_11925);
nand U12096 (N_12096,N_11595,N_11734);
xnor U12097 (N_12097,N_11862,N_11946);
xor U12098 (N_12098,N_11558,N_11563);
and U12099 (N_12099,N_11400,N_11623);
or U12100 (N_12100,N_11456,N_11628);
or U12101 (N_12101,N_11676,N_11976);
nand U12102 (N_12102,N_11856,N_11627);
nor U12103 (N_12103,N_11795,N_11473);
and U12104 (N_12104,N_11404,N_11835);
nand U12105 (N_12105,N_11546,N_11423);
nand U12106 (N_12106,N_11420,N_11657);
or U12107 (N_12107,N_11757,N_11985);
nor U12108 (N_12108,N_11747,N_11979);
xnor U12109 (N_12109,N_11463,N_11635);
and U12110 (N_12110,N_11601,N_11487);
nor U12111 (N_12111,N_11830,N_11731);
nand U12112 (N_12112,N_11531,N_11954);
or U12113 (N_12113,N_11667,N_11849);
xnor U12114 (N_12114,N_11479,N_11749);
or U12115 (N_12115,N_11439,N_11501);
nor U12116 (N_12116,N_11461,N_11854);
xor U12117 (N_12117,N_11980,N_11434);
xnor U12118 (N_12118,N_11974,N_11963);
xnor U12119 (N_12119,N_11783,N_11678);
nand U12120 (N_12120,N_11719,N_11822);
or U12121 (N_12121,N_11736,N_11881);
nand U12122 (N_12122,N_11713,N_11755);
nor U12123 (N_12123,N_11771,N_11724);
nor U12124 (N_12124,N_11551,N_11492);
or U12125 (N_12125,N_11816,N_11445);
xor U12126 (N_12126,N_11966,N_11521);
or U12127 (N_12127,N_11672,N_11526);
nand U12128 (N_12128,N_11720,N_11859);
xnor U12129 (N_12129,N_11885,N_11879);
xor U12130 (N_12130,N_11666,N_11682);
or U12131 (N_12131,N_11926,N_11616);
or U12132 (N_12132,N_11969,N_11688);
xnor U12133 (N_12133,N_11455,N_11471);
or U12134 (N_12134,N_11645,N_11704);
nand U12135 (N_12135,N_11626,N_11902);
xor U12136 (N_12136,N_11842,N_11436);
nor U12137 (N_12137,N_11477,N_11721);
nor U12138 (N_12138,N_11580,N_11401);
or U12139 (N_12139,N_11681,N_11996);
xor U12140 (N_12140,N_11951,N_11787);
and U12141 (N_12141,N_11553,N_11448);
and U12142 (N_12142,N_11922,N_11695);
or U12143 (N_12143,N_11808,N_11630);
nand U12144 (N_12144,N_11614,N_11971);
or U12145 (N_12145,N_11562,N_11923);
nand U12146 (N_12146,N_11751,N_11769);
or U12147 (N_12147,N_11581,N_11450);
and U12148 (N_12148,N_11579,N_11647);
xnor U12149 (N_12149,N_11642,N_11832);
xor U12150 (N_12150,N_11615,N_11774);
and U12151 (N_12151,N_11402,N_11648);
and U12152 (N_12152,N_11525,N_11482);
nor U12153 (N_12153,N_11566,N_11536);
or U12154 (N_12154,N_11465,N_11433);
nand U12155 (N_12155,N_11584,N_11768);
xor U12156 (N_12156,N_11586,N_11429);
nor U12157 (N_12157,N_11425,N_11680);
nand U12158 (N_12158,N_11895,N_11940);
nand U12159 (N_12159,N_11977,N_11517);
nor U12160 (N_12160,N_11894,N_11811);
and U12161 (N_12161,N_11409,N_11817);
and U12162 (N_12162,N_11833,N_11786);
nand U12163 (N_12163,N_11415,N_11847);
nand U12164 (N_12164,N_11573,N_11462);
and U12165 (N_12165,N_11726,N_11765);
nand U12166 (N_12166,N_11978,N_11756);
nand U12167 (N_12167,N_11876,N_11693);
nand U12168 (N_12168,N_11481,N_11790);
or U12169 (N_12169,N_11729,N_11905);
xnor U12170 (N_12170,N_11836,N_11652);
nand U12171 (N_12171,N_11685,N_11883);
and U12172 (N_12172,N_11875,N_11524);
or U12173 (N_12173,N_11945,N_11488);
and U12174 (N_12174,N_11970,N_11571);
and U12175 (N_12175,N_11662,N_11855);
and U12176 (N_12176,N_11898,N_11793);
and U12177 (N_12177,N_11893,N_11619);
or U12178 (N_12178,N_11559,N_11897);
nand U12179 (N_12179,N_11541,N_11490);
nor U12180 (N_12180,N_11421,N_11937);
nand U12181 (N_12181,N_11631,N_11742);
xnor U12182 (N_12182,N_11510,N_11780);
nand U12183 (N_12183,N_11730,N_11723);
and U12184 (N_12184,N_11944,N_11810);
and U12185 (N_12185,N_11801,N_11707);
and U12186 (N_12186,N_11776,N_11624);
or U12187 (N_12187,N_11458,N_11964);
or U12188 (N_12188,N_11582,N_11474);
xnor U12189 (N_12189,N_11651,N_11622);
nor U12190 (N_12190,N_11936,N_11867);
and U12191 (N_12191,N_11637,N_11846);
or U12192 (N_12192,N_11956,N_11831);
or U12193 (N_12193,N_11728,N_11989);
nor U12194 (N_12194,N_11958,N_11869);
nor U12195 (N_12195,N_11857,N_11911);
and U12196 (N_12196,N_11706,N_11602);
and U12197 (N_12197,N_11987,N_11690);
or U12198 (N_12198,N_11552,N_11877);
xor U12199 (N_12199,N_11735,N_11698);
xor U12200 (N_12200,N_11807,N_11797);
nand U12201 (N_12201,N_11853,N_11781);
or U12202 (N_12202,N_11578,N_11743);
nand U12203 (N_12203,N_11752,N_11535);
nor U12204 (N_12204,N_11533,N_11605);
and U12205 (N_12205,N_11914,N_11689);
nand U12206 (N_12206,N_11538,N_11684);
or U12207 (N_12207,N_11834,N_11796);
xnor U12208 (N_12208,N_11784,N_11613);
xnor U12209 (N_12209,N_11585,N_11806);
nor U12210 (N_12210,N_11668,N_11556);
xnor U12211 (N_12211,N_11507,N_11443);
nor U12212 (N_12212,N_11791,N_11410);
nand U12213 (N_12213,N_11664,N_11428);
nor U12214 (N_12214,N_11871,N_11414);
or U12215 (N_12215,N_11417,N_11851);
and U12216 (N_12216,N_11740,N_11995);
nand U12217 (N_12217,N_11544,N_11545);
xor U12218 (N_12218,N_11715,N_11815);
nor U12219 (N_12219,N_11955,N_11654);
xor U12220 (N_12220,N_11686,N_11618);
nor U12221 (N_12221,N_11504,N_11494);
xnor U12222 (N_12222,N_11522,N_11475);
or U12223 (N_12223,N_11520,N_11863);
xor U12224 (N_12224,N_11696,N_11406);
xnor U12225 (N_12225,N_11705,N_11653);
or U12226 (N_12226,N_11564,N_11744);
nor U12227 (N_12227,N_11549,N_11868);
xnor U12228 (N_12228,N_11649,N_11590);
nor U12229 (N_12229,N_11454,N_11665);
or U12230 (N_12230,N_11986,N_11469);
nor U12231 (N_12231,N_11766,N_11427);
xor U12232 (N_12232,N_11418,N_11792);
nor U12233 (N_12233,N_11948,N_11534);
or U12234 (N_12234,N_11655,N_11984);
or U12235 (N_12235,N_11924,N_11413);
xor U12236 (N_12236,N_11753,N_11763);
xor U12237 (N_12237,N_11845,N_11610);
nor U12238 (N_12238,N_11677,N_11640);
nor U12239 (N_12239,N_11997,N_11697);
nor U12240 (N_12240,N_11782,N_11714);
nand U12241 (N_12241,N_11576,N_11820);
nand U12242 (N_12242,N_11470,N_11916);
nand U12243 (N_12243,N_11508,N_11814);
and U12244 (N_12244,N_11983,N_11975);
or U12245 (N_12245,N_11495,N_11512);
or U12246 (N_12246,N_11748,N_11692);
nand U12247 (N_12247,N_11548,N_11634);
nor U12248 (N_12248,N_11872,N_11675);
xor U12249 (N_12249,N_11982,N_11620);
nor U12250 (N_12250,N_11663,N_11502);
xor U12251 (N_12251,N_11999,N_11407);
nor U12252 (N_12252,N_11741,N_11646);
and U12253 (N_12253,N_11515,N_11809);
or U12254 (N_12254,N_11608,N_11823);
nand U12255 (N_12255,N_11530,N_11561);
nor U12256 (N_12256,N_11825,N_11499);
and U12257 (N_12257,N_11972,N_11632);
xnor U12258 (N_12258,N_11930,N_11500);
and U12259 (N_12259,N_11906,N_11733);
nand U12260 (N_12260,N_11464,N_11506);
and U12261 (N_12261,N_11660,N_11967);
or U12262 (N_12262,N_11929,N_11800);
xnor U12263 (N_12263,N_11779,N_11422);
nand U12264 (N_12264,N_11540,N_11821);
nor U12265 (N_12265,N_11592,N_11593);
and U12266 (N_12266,N_11617,N_11457);
xnor U12267 (N_12267,N_11612,N_11880);
and U12268 (N_12268,N_11516,N_11865);
nand U12269 (N_12269,N_11827,N_11511);
and U12270 (N_12270,N_11703,N_11950);
nand U12271 (N_12271,N_11981,N_11850);
xnor U12272 (N_12272,N_11641,N_11442);
nor U12273 (N_12273,N_11947,N_11826);
and U12274 (N_12274,N_11888,N_11419);
and U12275 (N_12275,N_11670,N_11452);
or U12276 (N_12276,N_11716,N_11737);
nor U12277 (N_12277,N_11599,N_11874);
nand U12278 (N_12278,N_11841,N_11962);
nor U12279 (N_12279,N_11591,N_11758);
and U12280 (N_12280,N_11478,N_11843);
nand U12281 (N_12281,N_11785,N_11818);
or U12282 (N_12282,N_11762,N_11503);
or U12283 (N_12283,N_11745,N_11973);
or U12284 (N_12284,N_11935,N_11920);
xor U12285 (N_12285,N_11518,N_11918);
or U12286 (N_12286,N_11812,N_11773);
xor U12287 (N_12287,N_11547,N_11484);
and U12288 (N_12288,N_11968,N_11939);
nand U12289 (N_12289,N_11909,N_11557);
nand U12290 (N_12290,N_11824,N_11694);
or U12291 (N_12291,N_11887,N_11941);
nor U12292 (N_12292,N_11491,N_11607);
or U12293 (N_12293,N_11802,N_11588);
nor U12294 (N_12294,N_11764,N_11819);
and U12295 (N_12295,N_11486,N_11505);
or U12296 (N_12296,N_11539,N_11717);
and U12297 (N_12297,N_11990,N_11878);
or U12298 (N_12298,N_11912,N_11889);
or U12299 (N_12299,N_11523,N_11907);
nor U12300 (N_12300,N_11777,N_11978);
nor U12301 (N_12301,N_11479,N_11697);
nand U12302 (N_12302,N_11517,N_11590);
xor U12303 (N_12303,N_11905,N_11833);
nor U12304 (N_12304,N_11765,N_11937);
and U12305 (N_12305,N_11512,N_11755);
and U12306 (N_12306,N_11708,N_11541);
or U12307 (N_12307,N_11589,N_11461);
nor U12308 (N_12308,N_11785,N_11852);
nand U12309 (N_12309,N_11708,N_11432);
xor U12310 (N_12310,N_11896,N_11556);
or U12311 (N_12311,N_11454,N_11947);
and U12312 (N_12312,N_11819,N_11672);
nand U12313 (N_12313,N_11793,N_11968);
nor U12314 (N_12314,N_11751,N_11890);
nor U12315 (N_12315,N_11719,N_11911);
or U12316 (N_12316,N_11883,N_11627);
nand U12317 (N_12317,N_11608,N_11716);
or U12318 (N_12318,N_11414,N_11565);
nand U12319 (N_12319,N_11419,N_11590);
nand U12320 (N_12320,N_11533,N_11862);
nand U12321 (N_12321,N_11593,N_11999);
xnor U12322 (N_12322,N_11849,N_11983);
nor U12323 (N_12323,N_11607,N_11490);
or U12324 (N_12324,N_11551,N_11642);
or U12325 (N_12325,N_11644,N_11713);
nand U12326 (N_12326,N_11492,N_11885);
xor U12327 (N_12327,N_11582,N_11408);
or U12328 (N_12328,N_11556,N_11948);
nor U12329 (N_12329,N_11580,N_11532);
xor U12330 (N_12330,N_11563,N_11452);
or U12331 (N_12331,N_11809,N_11517);
xor U12332 (N_12332,N_11443,N_11817);
and U12333 (N_12333,N_11669,N_11914);
nand U12334 (N_12334,N_11732,N_11876);
and U12335 (N_12335,N_11454,N_11970);
or U12336 (N_12336,N_11666,N_11943);
xor U12337 (N_12337,N_11666,N_11676);
and U12338 (N_12338,N_11713,N_11665);
and U12339 (N_12339,N_11415,N_11776);
xor U12340 (N_12340,N_11506,N_11891);
xor U12341 (N_12341,N_11511,N_11589);
and U12342 (N_12342,N_11472,N_11810);
and U12343 (N_12343,N_11771,N_11943);
xor U12344 (N_12344,N_11807,N_11982);
or U12345 (N_12345,N_11855,N_11484);
or U12346 (N_12346,N_11992,N_11528);
and U12347 (N_12347,N_11447,N_11603);
and U12348 (N_12348,N_11715,N_11433);
xor U12349 (N_12349,N_11433,N_11425);
xor U12350 (N_12350,N_11896,N_11898);
nor U12351 (N_12351,N_11879,N_11892);
xor U12352 (N_12352,N_11748,N_11706);
nand U12353 (N_12353,N_11659,N_11700);
nor U12354 (N_12354,N_11726,N_11459);
or U12355 (N_12355,N_11939,N_11696);
nand U12356 (N_12356,N_11812,N_11984);
nor U12357 (N_12357,N_11826,N_11964);
nor U12358 (N_12358,N_11511,N_11629);
xor U12359 (N_12359,N_11939,N_11512);
or U12360 (N_12360,N_11737,N_11455);
nand U12361 (N_12361,N_11780,N_11508);
xor U12362 (N_12362,N_11875,N_11572);
and U12363 (N_12363,N_11938,N_11562);
xnor U12364 (N_12364,N_11731,N_11646);
nand U12365 (N_12365,N_11966,N_11649);
nand U12366 (N_12366,N_11556,N_11743);
nand U12367 (N_12367,N_11804,N_11568);
or U12368 (N_12368,N_11482,N_11838);
nor U12369 (N_12369,N_11776,N_11866);
nand U12370 (N_12370,N_11822,N_11547);
nor U12371 (N_12371,N_11541,N_11470);
xnor U12372 (N_12372,N_11734,N_11798);
and U12373 (N_12373,N_11944,N_11855);
nor U12374 (N_12374,N_11543,N_11657);
or U12375 (N_12375,N_11785,N_11961);
xor U12376 (N_12376,N_11590,N_11705);
nand U12377 (N_12377,N_11693,N_11691);
and U12378 (N_12378,N_11798,N_11441);
and U12379 (N_12379,N_11530,N_11413);
nor U12380 (N_12380,N_11957,N_11477);
nor U12381 (N_12381,N_11406,N_11871);
and U12382 (N_12382,N_11773,N_11886);
xnor U12383 (N_12383,N_11509,N_11843);
xor U12384 (N_12384,N_11550,N_11556);
and U12385 (N_12385,N_11946,N_11978);
xnor U12386 (N_12386,N_11605,N_11513);
nand U12387 (N_12387,N_11533,N_11568);
xor U12388 (N_12388,N_11848,N_11503);
xor U12389 (N_12389,N_11556,N_11806);
nand U12390 (N_12390,N_11817,N_11927);
nor U12391 (N_12391,N_11854,N_11874);
or U12392 (N_12392,N_11972,N_11535);
or U12393 (N_12393,N_11708,N_11682);
xor U12394 (N_12394,N_11678,N_11931);
nor U12395 (N_12395,N_11647,N_11728);
xor U12396 (N_12396,N_11707,N_11443);
and U12397 (N_12397,N_11708,N_11849);
xnor U12398 (N_12398,N_11586,N_11605);
xnor U12399 (N_12399,N_11677,N_11580);
or U12400 (N_12400,N_11677,N_11654);
nor U12401 (N_12401,N_11952,N_11746);
xnor U12402 (N_12402,N_11896,N_11451);
nand U12403 (N_12403,N_11545,N_11952);
nor U12404 (N_12404,N_11406,N_11815);
xnor U12405 (N_12405,N_11759,N_11979);
and U12406 (N_12406,N_11426,N_11467);
and U12407 (N_12407,N_11515,N_11622);
nand U12408 (N_12408,N_11721,N_11750);
and U12409 (N_12409,N_11591,N_11645);
nor U12410 (N_12410,N_11588,N_11857);
nor U12411 (N_12411,N_11973,N_11439);
xnor U12412 (N_12412,N_11604,N_11939);
and U12413 (N_12413,N_11875,N_11943);
and U12414 (N_12414,N_11940,N_11804);
xor U12415 (N_12415,N_11576,N_11818);
xnor U12416 (N_12416,N_11466,N_11637);
nand U12417 (N_12417,N_11576,N_11759);
nand U12418 (N_12418,N_11702,N_11884);
or U12419 (N_12419,N_11671,N_11626);
xnor U12420 (N_12420,N_11502,N_11924);
and U12421 (N_12421,N_11476,N_11677);
xor U12422 (N_12422,N_11896,N_11525);
xnor U12423 (N_12423,N_11476,N_11857);
and U12424 (N_12424,N_11585,N_11944);
xor U12425 (N_12425,N_11554,N_11516);
and U12426 (N_12426,N_11877,N_11529);
and U12427 (N_12427,N_11980,N_11862);
xor U12428 (N_12428,N_11482,N_11728);
nor U12429 (N_12429,N_11856,N_11913);
or U12430 (N_12430,N_11746,N_11700);
and U12431 (N_12431,N_11586,N_11866);
xor U12432 (N_12432,N_11536,N_11412);
nor U12433 (N_12433,N_11598,N_11513);
and U12434 (N_12434,N_11630,N_11524);
nand U12435 (N_12435,N_11795,N_11792);
xor U12436 (N_12436,N_11530,N_11865);
nor U12437 (N_12437,N_11585,N_11413);
nand U12438 (N_12438,N_11700,N_11478);
and U12439 (N_12439,N_11634,N_11741);
nor U12440 (N_12440,N_11935,N_11455);
and U12441 (N_12441,N_11905,N_11480);
xor U12442 (N_12442,N_11790,N_11806);
and U12443 (N_12443,N_11769,N_11616);
xnor U12444 (N_12444,N_11763,N_11625);
and U12445 (N_12445,N_11499,N_11701);
or U12446 (N_12446,N_11629,N_11950);
nor U12447 (N_12447,N_11518,N_11488);
xor U12448 (N_12448,N_11922,N_11874);
and U12449 (N_12449,N_11523,N_11980);
xnor U12450 (N_12450,N_11519,N_11718);
or U12451 (N_12451,N_11822,N_11949);
and U12452 (N_12452,N_11618,N_11748);
nor U12453 (N_12453,N_11589,N_11569);
nand U12454 (N_12454,N_11775,N_11710);
xor U12455 (N_12455,N_11685,N_11755);
nor U12456 (N_12456,N_11710,N_11751);
or U12457 (N_12457,N_11499,N_11736);
nand U12458 (N_12458,N_11681,N_11837);
nand U12459 (N_12459,N_11977,N_11982);
xor U12460 (N_12460,N_11414,N_11614);
nor U12461 (N_12461,N_11992,N_11959);
or U12462 (N_12462,N_11887,N_11615);
xnor U12463 (N_12463,N_11871,N_11822);
or U12464 (N_12464,N_11976,N_11856);
nor U12465 (N_12465,N_11717,N_11594);
and U12466 (N_12466,N_11487,N_11742);
or U12467 (N_12467,N_11957,N_11567);
nand U12468 (N_12468,N_11726,N_11403);
nor U12469 (N_12469,N_11916,N_11679);
and U12470 (N_12470,N_11427,N_11919);
nor U12471 (N_12471,N_11627,N_11683);
or U12472 (N_12472,N_11957,N_11728);
xnor U12473 (N_12473,N_11804,N_11780);
nor U12474 (N_12474,N_11818,N_11919);
or U12475 (N_12475,N_11741,N_11424);
nor U12476 (N_12476,N_11478,N_11544);
xor U12477 (N_12477,N_11933,N_11928);
xnor U12478 (N_12478,N_11582,N_11889);
or U12479 (N_12479,N_11429,N_11441);
and U12480 (N_12480,N_11976,N_11885);
xor U12481 (N_12481,N_11981,N_11995);
and U12482 (N_12482,N_11711,N_11915);
nand U12483 (N_12483,N_11498,N_11767);
xnor U12484 (N_12484,N_11595,N_11646);
nor U12485 (N_12485,N_11449,N_11758);
nand U12486 (N_12486,N_11435,N_11533);
and U12487 (N_12487,N_11873,N_11459);
and U12488 (N_12488,N_11506,N_11995);
and U12489 (N_12489,N_11664,N_11405);
or U12490 (N_12490,N_11509,N_11452);
xnor U12491 (N_12491,N_11828,N_11936);
nor U12492 (N_12492,N_11688,N_11746);
and U12493 (N_12493,N_11926,N_11619);
nand U12494 (N_12494,N_11649,N_11753);
nand U12495 (N_12495,N_11402,N_11730);
nand U12496 (N_12496,N_11804,N_11420);
nand U12497 (N_12497,N_11915,N_11431);
or U12498 (N_12498,N_11517,N_11431);
nor U12499 (N_12499,N_11929,N_11633);
xor U12500 (N_12500,N_11928,N_11676);
or U12501 (N_12501,N_11474,N_11728);
or U12502 (N_12502,N_11538,N_11466);
nor U12503 (N_12503,N_11745,N_11859);
and U12504 (N_12504,N_11436,N_11908);
and U12505 (N_12505,N_11893,N_11980);
xor U12506 (N_12506,N_11597,N_11822);
nor U12507 (N_12507,N_11555,N_11963);
xnor U12508 (N_12508,N_11518,N_11894);
nand U12509 (N_12509,N_11721,N_11665);
nor U12510 (N_12510,N_11608,N_11402);
xor U12511 (N_12511,N_11973,N_11724);
or U12512 (N_12512,N_11635,N_11743);
nand U12513 (N_12513,N_11760,N_11603);
nor U12514 (N_12514,N_11581,N_11792);
or U12515 (N_12515,N_11969,N_11474);
nand U12516 (N_12516,N_11550,N_11521);
or U12517 (N_12517,N_11644,N_11856);
nand U12518 (N_12518,N_11671,N_11600);
or U12519 (N_12519,N_11689,N_11637);
xnor U12520 (N_12520,N_11525,N_11444);
nand U12521 (N_12521,N_11904,N_11618);
and U12522 (N_12522,N_11718,N_11907);
and U12523 (N_12523,N_11721,N_11983);
nand U12524 (N_12524,N_11797,N_11620);
nand U12525 (N_12525,N_11712,N_11719);
and U12526 (N_12526,N_11555,N_11489);
or U12527 (N_12527,N_11720,N_11576);
and U12528 (N_12528,N_11448,N_11403);
nor U12529 (N_12529,N_11495,N_11910);
or U12530 (N_12530,N_11920,N_11419);
or U12531 (N_12531,N_11780,N_11813);
or U12532 (N_12532,N_11846,N_11428);
nand U12533 (N_12533,N_11637,N_11523);
nand U12534 (N_12534,N_11919,N_11831);
nor U12535 (N_12535,N_11695,N_11572);
nand U12536 (N_12536,N_11968,N_11739);
nor U12537 (N_12537,N_11591,N_11913);
xnor U12538 (N_12538,N_11963,N_11783);
and U12539 (N_12539,N_11748,N_11862);
xor U12540 (N_12540,N_11758,N_11691);
xnor U12541 (N_12541,N_11972,N_11850);
nand U12542 (N_12542,N_11993,N_11940);
nor U12543 (N_12543,N_11416,N_11680);
nor U12544 (N_12544,N_11588,N_11410);
nand U12545 (N_12545,N_11559,N_11503);
nor U12546 (N_12546,N_11601,N_11534);
nand U12547 (N_12547,N_11960,N_11499);
nor U12548 (N_12548,N_11983,N_11959);
nand U12549 (N_12549,N_11504,N_11986);
or U12550 (N_12550,N_11593,N_11451);
or U12551 (N_12551,N_11993,N_11644);
nand U12552 (N_12552,N_11837,N_11993);
or U12553 (N_12553,N_11799,N_11533);
nand U12554 (N_12554,N_11655,N_11888);
nand U12555 (N_12555,N_11672,N_11844);
or U12556 (N_12556,N_11667,N_11656);
xor U12557 (N_12557,N_11806,N_11953);
and U12558 (N_12558,N_11440,N_11761);
xor U12559 (N_12559,N_11810,N_11637);
and U12560 (N_12560,N_11962,N_11770);
and U12561 (N_12561,N_11713,N_11721);
nand U12562 (N_12562,N_11906,N_11504);
nor U12563 (N_12563,N_11851,N_11791);
xor U12564 (N_12564,N_11775,N_11528);
or U12565 (N_12565,N_11438,N_11563);
nand U12566 (N_12566,N_11685,N_11448);
nand U12567 (N_12567,N_11409,N_11954);
and U12568 (N_12568,N_11616,N_11491);
nand U12569 (N_12569,N_11672,N_11889);
or U12570 (N_12570,N_11836,N_11978);
nand U12571 (N_12571,N_11685,N_11834);
nor U12572 (N_12572,N_11413,N_11692);
xnor U12573 (N_12573,N_11444,N_11556);
xnor U12574 (N_12574,N_11580,N_11486);
xnor U12575 (N_12575,N_11468,N_11706);
nand U12576 (N_12576,N_11815,N_11994);
xor U12577 (N_12577,N_11792,N_11957);
xnor U12578 (N_12578,N_11542,N_11776);
nand U12579 (N_12579,N_11833,N_11872);
nand U12580 (N_12580,N_11763,N_11550);
or U12581 (N_12581,N_11866,N_11891);
nand U12582 (N_12582,N_11510,N_11913);
nor U12583 (N_12583,N_11802,N_11875);
nor U12584 (N_12584,N_11946,N_11417);
and U12585 (N_12585,N_11936,N_11582);
or U12586 (N_12586,N_11444,N_11544);
xnor U12587 (N_12587,N_11486,N_11701);
nand U12588 (N_12588,N_11426,N_11839);
xor U12589 (N_12589,N_11964,N_11647);
nor U12590 (N_12590,N_11543,N_11688);
nor U12591 (N_12591,N_11865,N_11998);
or U12592 (N_12592,N_11468,N_11787);
and U12593 (N_12593,N_11939,N_11480);
nor U12594 (N_12594,N_11560,N_11922);
xnor U12595 (N_12595,N_11446,N_11617);
and U12596 (N_12596,N_11715,N_11809);
nor U12597 (N_12597,N_11474,N_11909);
and U12598 (N_12598,N_11530,N_11982);
nand U12599 (N_12599,N_11750,N_11578);
or U12600 (N_12600,N_12576,N_12478);
nor U12601 (N_12601,N_12514,N_12445);
nand U12602 (N_12602,N_12570,N_12199);
xor U12603 (N_12603,N_12437,N_12475);
xnor U12604 (N_12604,N_12196,N_12515);
and U12605 (N_12605,N_12556,N_12581);
nor U12606 (N_12606,N_12489,N_12592);
and U12607 (N_12607,N_12200,N_12119);
and U12608 (N_12608,N_12415,N_12062);
and U12609 (N_12609,N_12168,N_12153);
nor U12610 (N_12610,N_12346,N_12539);
and U12611 (N_12611,N_12281,N_12438);
nand U12612 (N_12612,N_12145,N_12340);
xnor U12613 (N_12613,N_12543,N_12375);
or U12614 (N_12614,N_12076,N_12257);
or U12615 (N_12615,N_12560,N_12042);
nor U12616 (N_12616,N_12597,N_12063);
nand U12617 (N_12617,N_12580,N_12313);
xnor U12618 (N_12618,N_12315,N_12506);
nand U12619 (N_12619,N_12216,N_12289);
nand U12620 (N_12620,N_12084,N_12279);
xnor U12621 (N_12621,N_12277,N_12136);
xnor U12622 (N_12622,N_12057,N_12227);
nand U12623 (N_12623,N_12088,N_12558);
nand U12624 (N_12624,N_12518,N_12473);
or U12625 (N_12625,N_12362,N_12274);
and U12626 (N_12626,N_12266,N_12567);
and U12627 (N_12627,N_12228,N_12588);
nand U12628 (N_12628,N_12085,N_12432);
and U12629 (N_12629,N_12133,N_12115);
or U12630 (N_12630,N_12511,N_12190);
or U12631 (N_12631,N_12400,N_12010);
or U12632 (N_12632,N_12409,N_12155);
nor U12633 (N_12633,N_12165,N_12380);
nor U12634 (N_12634,N_12564,N_12156);
nor U12635 (N_12635,N_12268,N_12512);
xnor U12636 (N_12636,N_12272,N_12218);
xor U12637 (N_12637,N_12466,N_12083);
nand U12638 (N_12638,N_12307,N_12540);
nor U12639 (N_12639,N_12278,N_12056);
or U12640 (N_12640,N_12534,N_12080);
and U12641 (N_12641,N_12286,N_12126);
xnor U12642 (N_12642,N_12501,N_12535);
nor U12643 (N_12643,N_12565,N_12276);
or U12644 (N_12644,N_12548,N_12325);
or U12645 (N_12645,N_12127,N_12214);
xnor U12646 (N_12646,N_12033,N_12555);
xnor U12647 (N_12647,N_12270,N_12064);
and U12648 (N_12648,N_12249,N_12171);
xnor U12649 (N_12649,N_12446,N_12338);
and U12650 (N_12650,N_12184,N_12179);
or U12651 (N_12651,N_12436,N_12566);
xor U12652 (N_12652,N_12455,N_12053);
nand U12653 (N_12653,N_12385,N_12383);
nand U12654 (N_12654,N_12141,N_12202);
or U12655 (N_12655,N_12001,N_12364);
or U12656 (N_12656,N_12073,N_12495);
xnor U12657 (N_12657,N_12284,N_12020);
nand U12658 (N_12658,N_12476,N_12132);
nand U12659 (N_12659,N_12028,N_12187);
nor U12660 (N_12660,N_12203,N_12186);
xor U12661 (N_12661,N_12298,N_12331);
xnor U12662 (N_12662,N_12386,N_12144);
nor U12663 (N_12663,N_12069,N_12549);
and U12664 (N_12664,N_12061,N_12074);
and U12665 (N_12665,N_12529,N_12522);
and U12666 (N_12666,N_12381,N_12269);
xor U12667 (N_12667,N_12154,N_12584);
and U12668 (N_12668,N_12009,N_12220);
or U12669 (N_12669,N_12356,N_12414);
or U12670 (N_12670,N_12508,N_12265);
and U12671 (N_12671,N_12367,N_12273);
nor U12672 (N_12672,N_12547,N_12305);
nor U12673 (N_12673,N_12398,N_12113);
nand U12674 (N_12674,N_12431,N_12236);
nand U12675 (N_12675,N_12123,N_12102);
and U12676 (N_12676,N_12421,N_12246);
xor U12677 (N_12677,N_12324,N_12538);
and U12678 (N_12678,N_12497,N_12354);
or U12679 (N_12679,N_12129,N_12034);
and U12680 (N_12680,N_12321,N_12388);
or U12681 (N_12681,N_12244,N_12271);
and U12682 (N_12682,N_12092,N_12389);
or U12683 (N_12683,N_12553,N_12222);
nand U12684 (N_12684,N_12103,N_12152);
nand U12685 (N_12685,N_12349,N_12245);
and U12686 (N_12686,N_12086,N_12045);
nor U12687 (N_12687,N_12376,N_12348);
nor U12688 (N_12688,N_12173,N_12079);
or U12689 (N_12689,N_12505,N_12259);
xor U12690 (N_12690,N_12365,N_12101);
xor U12691 (N_12691,N_12328,N_12330);
or U12692 (N_12692,N_12430,N_12509);
xnor U12693 (N_12693,N_12206,N_12453);
nand U12694 (N_12694,N_12402,N_12451);
nor U12695 (N_12695,N_12462,N_12551);
xor U12696 (N_12696,N_12254,N_12146);
nor U12697 (N_12697,N_12049,N_12358);
or U12698 (N_12698,N_12089,N_12311);
nor U12699 (N_12699,N_12366,N_12219);
nor U12700 (N_12700,N_12379,N_12377);
and U12701 (N_12701,N_12066,N_12517);
nor U12702 (N_12702,N_12541,N_12559);
xnor U12703 (N_12703,N_12308,N_12104);
or U12704 (N_12704,N_12019,N_12160);
and U12705 (N_12705,N_12468,N_12111);
and U12706 (N_12706,N_12295,N_12467);
xnor U12707 (N_12707,N_12006,N_12137);
or U12708 (N_12708,N_12312,N_12590);
nor U12709 (N_12709,N_12485,N_12335);
nor U12710 (N_12710,N_12327,N_12230);
or U12711 (N_12711,N_12240,N_12166);
nand U12712 (N_12712,N_12239,N_12121);
nor U12713 (N_12713,N_12122,N_12371);
xnor U12714 (N_12714,N_12003,N_12068);
and U12715 (N_12715,N_12435,N_12359);
or U12716 (N_12716,N_12285,N_12428);
xor U12717 (N_12717,N_12233,N_12208);
nor U12718 (N_12718,N_12169,N_12194);
nor U12719 (N_12719,N_12460,N_12051);
or U12720 (N_12720,N_12545,N_12180);
nand U12721 (N_12721,N_12118,N_12296);
or U12722 (N_12722,N_12162,N_12442);
nor U12723 (N_12723,N_12036,N_12072);
or U12724 (N_12724,N_12091,N_12472);
nand U12725 (N_12725,N_12316,N_12484);
nand U12726 (N_12726,N_12352,N_12177);
and U12727 (N_12727,N_12164,N_12302);
nand U12728 (N_12728,N_12411,N_12158);
nand U12729 (N_12729,N_12382,N_12077);
and U12730 (N_12730,N_12050,N_12107);
and U12731 (N_12731,N_12557,N_12023);
and U12732 (N_12732,N_12572,N_12544);
xnor U12733 (N_12733,N_12192,N_12004);
or U12734 (N_12734,N_12212,N_12013);
xor U12735 (N_12735,N_12052,N_12550);
nor U12736 (N_12736,N_12563,N_12135);
and U12737 (N_12737,N_12444,N_12441);
nand U12738 (N_12738,N_12439,N_12403);
nor U12739 (N_12739,N_12314,N_12114);
nand U12740 (N_12740,N_12070,N_12320);
or U12741 (N_12741,N_12189,N_12465);
nand U12742 (N_12742,N_12372,N_12456);
nor U12743 (N_12743,N_12542,N_12591);
or U12744 (N_12744,N_12291,N_12474);
and U12745 (N_12745,N_12578,N_12554);
xor U12746 (N_12746,N_12443,N_12067);
nand U12747 (N_12747,N_12477,N_12207);
or U12748 (N_12748,N_12260,N_12215);
xor U12749 (N_12749,N_12420,N_12015);
nand U12750 (N_12750,N_12205,N_12329);
or U12751 (N_12751,N_12392,N_12157);
xnor U12752 (N_12752,N_12434,N_12536);
nand U12753 (N_12753,N_12110,N_12232);
or U12754 (N_12754,N_12450,N_12098);
nand U12755 (N_12755,N_12297,N_12594);
xor U12756 (N_12756,N_12410,N_12502);
nand U12757 (N_12757,N_12520,N_12575);
and U12758 (N_12758,N_12097,N_12041);
or U12759 (N_12759,N_12256,N_12226);
nor U12760 (N_12760,N_12470,N_12336);
and U12761 (N_12761,N_12503,N_12482);
nor U12762 (N_12762,N_12191,N_12014);
nor U12763 (N_12763,N_12176,N_12280);
xor U12764 (N_12764,N_12494,N_12391);
or U12765 (N_12765,N_12306,N_12526);
nor U12766 (N_12766,N_12011,N_12483);
nor U12767 (N_12767,N_12387,N_12243);
xnor U12768 (N_12768,N_12109,N_12587);
nor U12769 (N_12769,N_12188,N_12290);
and U12770 (N_12770,N_12140,N_12027);
nand U12771 (N_12771,N_12310,N_12530);
nand U12772 (N_12772,N_12163,N_12283);
or U12773 (N_12773,N_12419,N_12369);
nand U12774 (N_12774,N_12447,N_12363);
and U12775 (N_12775,N_12234,N_12337);
xnor U12776 (N_12776,N_12007,N_12504);
or U12777 (N_12777,N_12424,N_12026);
nor U12778 (N_12778,N_12397,N_12131);
nor U12779 (N_12779,N_12585,N_12116);
or U12780 (N_12780,N_12275,N_12598);
nor U12781 (N_12781,N_12595,N_12174);
nand U12782 (N_12782,N_12039,N_12108);
nor U12783 (N_12783,N_12481,N_12082);
nor U12784 (N_12784,N_12422,N_12251);
nand U12785 (N_12785,N_12303,N_12405);
and U12786 (N_12786,N_12000,N_12055);
or U12787 (N_12787,N_12525,N_12416);
or U12788 (N_12788,N_12147,N_12360);
xor U12789 (N_12789,N_12406,N_12537);
xnor U12790 (N_12790,N_12461,N_12343);
nand U12791 (N_12791,N_12008,N_12464);
xor U12792 (N_12792,N_12573,N_12571);
nor U12793 (N_12793,N_12071,N_12247);
or U12794 (N_12794,N_12440,N_12326);
nand U12795 (N_12795,N_12095,N_12081);
nor U12796 (N_12796,N_12596,N_12025);
nor U12797 (N_12797,N_12225,N_12459);
nor U12798 (N_12798,N_12150,N_12087);
and U12799 (N_12799,N_12401,N_12117);
or U12800 (N_12800,N_12396,N_12344);
xnor U12801 (N_12801,N_12035,N_12394);
nor U12802 (N_12802,N_12390,N_12238);
nand U12803 (N_12803,N_12599,N_12263);
xnor U12804 (N_12804,N_12323,N_12350);
and U12805 (N_12805,N_12458,N_12574);
xnor U12806 (N_12806,N_12499,N_12353);
and U12807 (N_12807,N_12378,N_12005);
or U12808 (N_12808,N_12427,N_12112);
nor U12809 (N_12809,N_12094,N_12048);
nor U12810 (N_12810,N_12407,N_12317);
and U12811 (N_12811,N_12037,N_12490);
nand U12812 (N_12812,N_12075,N_12292);
xnor U12813 (N_12813,N_12524,N_12469);
and U12814 (N_12814,N_12301,N_12583);
nor U12815 (N_12815,N_12167,N_12017);
and U12816 (N_12816,N_12425,N_12347);
or U12817 (N_12817,N_12496,N_12204);
or U12818 (N_12818,N_12498,N_12488);
and U12819 (N_12819,N_12139,N_12471);
and U12820 (N_12820,N_12217,N_12134);
and U12821 (N_12821,N_12492,N_12175);
nand U12822 (N_12822,N_12293,N_12357);
or U12823 (N_12823,N_12031,N_12252);
xor U12824 (N_12824,N_12149,N_12448);
nand U12825 (N_12825,N_12513,N_12493);
or U12826 (N_12826,N_12142,N_12449);
or U12827 (N_12827,N_12510,N_12429);
xnor U12828 (N_12828,N_12183,N_12237);
nand U12829 (N_12829,N_12355,N_12374);
or U12830 (N_12830,N_12333,N_12030);
nor U12831 (N_12831,N_12248,N_12213);
xor U12832 (N_12832,N_12258,N_12589);
and U12833 (N_12833,N_12527,N_12128);
and U12834 (N_12834,N_12253,N_12546);
or U12835 (N_12835,N_12143,N_12264);
nand U12836 (N_12836,N_12224,N_12148);
or U12837 (N_12837,N_12267,N_12582);
and U12838 (N_12838,N_12255,N_12457);
and U12839 (N_12839,N_12193,N_12408);
or U12840 (N_12840,N_12361,N_12568);
nand U12841 (N_12841,N_12046,N_12022);
nand U12842 (N_12842,N_12021,N_12016);
xnor U12843 (N_12843,N_12454,N_12185);
and U12844 (N_12844,N_12404,N_12294);
xor U12845 (N_12845,N_12059,N_12433);
nand U12846 (N_12846,N_12309,N_12210);
or U12847 (N_12847,N_12373,N_12012);
or U12848 (N_12848,N_12507,N_12491);
or U12849 (N_12849,N_12029,N_12231);
nand U12850 (N_12850,N_12384,N_12304);
xnor U12851 (N_12851,N_12463,N_12120);
nand U12852 (N_12852,N_12368,N_12322);
or U12853 (N_12853,N_12500,N_12197);
nand U12854 (N_12854,N_12332,N_12531);
nand U12855 (N_12855,N_12521,N_12209);
and U12856 (N_12856,N_12593,N_12172);
xor U12857 (N_12857,N_12261,N_12486);
nor U12858 (N_12858,N_12479,N_12334);
xor U12859 (N_12859,N_12318,N_12130);
and U12860 (N_12860,N_12198,N_12452);
and U12861 (N_12861,N_12201,N_12351);
xnor U12862 (N_12862,N_12093,N_12096);
xnor U12863 (N_12863,N_12282,N_12523);
or U12864 (N_12864,N_12287,N_12242);
and U12865 (N_12865,N_12412,N_12299);
or U12866 (N_12866,N_12182,N_12105);
nor U12867 (N_12867,N_12229,N_12032);
nand U12868 (N_12868,N_12533,N_12040);
or U12869 (N_12869,N_12178,N_12345);
nor U12870 (N_12870,N_12519,N_12043);
nand U12871 (N_12871,N_12342,N_12399);
nand U12872 (N_12872,N_12516,N_12561);
or U12873 (N_12873,N_12223,N_12002);
nand U12874 (N_12874,N_12562,N_12370);
nand U12875 (N_12875,N_12138,N_12339);
xor U12876 (N_12876,N_12417,N_12235);
nand U12877 (N_12877,N_12181,N_12159);
nor U12878 (N_12878,N_12319,N_12480);
nand U12879 (N_12879,N_12024,N_12221);
or U12880 (N_12880,N_12125,N_12241);
xor U12881 (N_12881,N_12099,N_12426);
or U12882 (N_12882,N_12552,N_12393);
xnor U12883 (N_12883,N_12395,N_12528);
or U12884 (N_12884,N_12487,N_12018);
or U12885 (N_12885,N_12586,N_12418);
nand U12886 (N_12886,N_12065,N_12577);
and U12887 (N_12887,N_12195,N_12151);
nand U12888 (N_12888,N_12047,N_12060);
nor U12889 (N_12889,N_12090,N_12423);
and U12890 (N_12890,N_12579,N_12211);
or U12891 (N_12891,N_12161,N_12262);
and U12892 (N_12892,N_12532,N_12250);
nand U12893 (N_12893,N_12413,N_12044);
nor U12894 (N_12894,N_12078,N_12038);
or U12895 (N_12895,N_12100,N_12341);
or U12896 (N_12896,N_12106,N_12569);
nand U12897 (N_12897,N_12058,N_12124);
nand U12898 (N_12898,N_12288,N_12170);
xor U12899 (N_12899,N_12054,N_12300);
or U12900 (N_12900,N_12040,N_12067);
nor U12901 (N_12901,N_12493,N_12379);
nor U12902 (N_12902,N_12183,N_12081);
or U12903 (N_12903,N_12258,N_12517);
xnor U12904 (N_12904,N_12343,N_12191);
nand U12905 (N_12905,N_12164,N_12521);
nor U12906 (N_12906,N_12306,N_12444);
nand U12907 (N_12907,N_12506,N_12529);
and U12908 (N_12908,N_12441,N_12427);
nand U12909 (N_12909,N_12506,N_12076);
or U12910 (N_12910,N_12231,N_12408);
or U12911 (N_12911,N_12485,N_12358);
or U12912 (N_12912,N_12587,N_12195);
nand U12913 (N_12913,N_12086,N_12207);
nand U12914 (N_12914,N_12411,N_12357);
xnor U12915 (N_12915,N_12529,N_12163);
nand U12916 (N_12916,N_12586,N_12217);
xor U12917 (N_12917,N_12336,N_12012);
and U12918 (N_12918,N_12539,N_12281);
and U12919 (N_12919,N_12189,N_12367);
and U12920 (N_12920,N_12111,N_12559);
nand U12921 (N_12921,N_12490,N_12260);
nor U12922 (N_12922,N_12342,N_12327);
and U12923 (N_12923,N_12060,N_12595);
and U12924 (N_12924,N_12019,N_12331);
xor U12925 (N_12925,N_12123,N_12254);
xor U12926 (N_12926,N_12545,N_12352);
nand U12927 (N_12927,N_12383,N_12495);
xnor U12928 (N_12928,N_12363,N_12451);
nand U12929 (N_12929,N_12422,N_12180);
and U12930 (N_12930,N_12509,N_12362);
nand U12931 (N_12931,N_12598,N_12362);
and U12932 (N_12932,N_12226,N_12483);
nand U12933 (N_12933,N_12223,N_12275);
nor U12934 (N_12934,N_12133,N_12300);
or U12935 (N_12935,N_12324,N_12166);
and U12936 (N_12936,N_12087,N_12142);
xor U12937 (N_12937,N_12524,N_12539);
or U12938 (N_12938,N_12592,N_12234);
nor U12939 (N_12939,N_12135,N_12518);
or U12940 (N_12940,N_12104,N_12595);
nand U12941 (N_12941,N_12010,N_12149);
nor U12942 (N_12942,N_12053,N_12344);
or U12943 (N_12943,N_12235,N_12126);
nor U12944 (N_12944,N_12384,N_12556);
and U12945 (N_12945,N_12115,N_12552);
and U12946 (N_12946,N_12514,N_12107);
xnor U12947 (N_12947,N_12306,N_12500);
or U12948 (N_12948,N_12150,N_12047);
xor U12949 (N_12949,N_12433,N_12328);
nor U12950 (N_12950,N_12526,N_12434);
nand U12951 (N_12951,N_12185,N_12573);
or U12952 (N_12952,N_12035,N_12057);
and U12953 (N_12953,N_12526,N_12254);
or U12954 (N_12954,N_12496,N_12306);
nor U12955 (N_12955,N_12158,N_12489);
and U12956 (N_12956,N_12236,N_12343);
xnor U12957 (N_12957,N_12063,N_12544);
nor U12958 (N_12958,N_12490,N_12007);
nand U12959 (N_12959,N_12364,N_12580);
and U12960 (N_12960,N_12537,N_12333);
nand U12961 (N_12961,N_12230,N_12006);
nor U12962 (N_12962,N_12523,N_12078);
nand U12963 (N_12963,N_12166,N_12287);
and U12964 (N_12964,N_12298,N_12143);
or U12965 (N_12965,N_12192,N_12223);
and U12966 (N_12966,N_12274,N_12176);
nand U12967 (N_12967,N_12557,N_12510);
and U12968 (N_12968,N_12370,N_12114);
or U12969 (N_12969,N_12252,N_12554);
and U12970 (N_12970,N_12332,N_12021);
and U12971 (N_12971,N_12071,N_12548);
and U12972 (N_12972,N_12231,N_12198);
xor U12973 (N_12973,N_12002,N_12403);
and U12974 (N_12974,N_12075,N_12125);
and U12975 (N_12975,N_12234,N_12588);
nand U12976 (N_12976,N_12203,N_12200);
nand U12977 (N_12977,N_12395,N_12125);
nor U12978 (N_12978,N_12012,N_12142);
nor U12979 (N_12979,N_12494,N_12362);
nand U12980 (N_12980,N_12166,N_12159);
or U12981 (N_12981,N_12348,N_12049);
xor U12982 (N_12982,N_12155,N_12229);
nor U12983 (N_12983,N_12548,N_12133);
or U12984 (N_12984,N_12267,N_12257);
nor U12985 (N_12985,N_12493,N_12343);
or U12986 (N_12986,N_12548,N_12599);
and U12987 (N_12987,N_12233,N_12543);
or U12988 (N_12988,N_12397,N_12088);
nand U12989 (N_12989,N_12431,N_12408);
nand U12990 (N_12990,N_12009,N_12555);
xnor U12991 (N_12991,N_12553,N_12484);
and U12992 (N_12992,N_12599,N_12083);
or U12993 (N_12993,N_12242,N_12486);
nor U12994 (N_12994,N_12169,N_12344);
nor U12995 (N_12995,N_12550,N_12139);
nor U12996 (N_12996,N_12308,N_12085);
xor U12997 (N_12997,N_12214,N_12004);
and U12998 (N_12998,N_12581,N_12246);
or U12999 (N_12999,N_12270,N_12186);
and U13000 (N_13000,N_12377,N_12439);
nand U13001 (N_13001,N_12130,N_12274);
nor U13002 (N_13002,N_12294,N_12156);
nand U13003 (N_13003,N_12371,N_12096);
nand U13004 (N_13004,N_12132,N_12243);
nor U13005 (N_13005,N_12551,N_12039);
and U13006 (N_13006,N_12459,N_12399);
or U13007 (N_13007,N_12112,N_12014);
or U13008 (N_13008,N_12059,N_12142);
nor U13009 (N_13009,N_12082,N_12168);
xor U13010 (N_13010,N_12044,N_12578);
xnor U13011 (N_13011,N_12182,N_12581);
and U13012 (N_13012,N_12309,N_12308);
nor U13013 (N_13013,N_12415,N_12149);
nor U13014 (N_13014,N_12002,N_12517);
nand U13015 (N_13015,N_12191,N_12292);
xnor U13016 (N_13016,N_12343,N_12323);
xor U13017 (N_13017,N_12207,N_12043);
xnor U13018 (N_13018,N_12220,N_12135);
xnor U13019 (N_13019,N_12079,N_12278);
xor U13020 (N_13020,N_12486,N_12034);
or U13021 (N_13021,N_12481,N_12561);
or U13022 (N_13022,N_12219,N_12113);
xor U13023 (N_13023,N_12115,N_12081);
xor U13024 (N_13024,N_12389,N_12297);
xor U13025 (N_13025,N_12129,N_12472);
nor U13026 (N_13026,N_12266,N_12004);
nor U13027 (N_13027,N_12445,N_12048);
or U13028 (N_13028,N_12322,N_12165);
xor U13029 (N_13029,N_12261,N_12125);
xnor U13030 (N_13030,N_12078,N_12037);
or U13031 (N_13031,N_12319,N_12565);
nor U13032 (N_13032,N_12558,N_12036);
nor U13033 (N_13033,N_12117,N_12350);
nand U13034 (N_13034,N_12129,N_12596);
xnor U13035 (N_13035,N_12001,N_12461);
xor U13036 (N_13036,N_12518,N_12272);
nand U13037 (N_13037,N_12055,N_12017);
or U13038 (N_13038,N_12055,N_12251);
or U13039 (N_13039,N_12306,N_12107);
and U13040 (N_13040,N_12534,N_12360);
nand U13041 (N_13041,N_12059,N_12015);
nor U13042 (N_13042,N_12183,N_12115);
nand U13043 (N_13043,N_12269,N_12103);
or U13044 (N_13044,N_12469,N_12532);
nand U13045 (N_13045,N_12585,N_12192);
nand U13046 (N_13046,N_12122,N_12564);
or U13047 (N_13047,N_12000,N_12187);
nand U13048 (N_13048,N_12246,N_12210);
nand U13049 (N_13049,N_12355,N_12001);
or U13050 (N_13050,N_12549,N_12187);
or U13051 (N_13051,N_12018,N_12517);
and U13052 (N_13052,N_12215,N_12012);
nand U13053 (N_13053,N_12583,N_12148);
and U13054 (N_13054,N_12490,N_12221);
or U13055 (N_13055,N_12203,N_12404);
or U13056 (N_13056,N_12055,N_12597);
nand U13057 (N_13057,N_12503,N_12362);
and U13058 (N_13058,N_12519,N_12419);
or U13059 (N_13059,N_12481,N_12105);
nor U13060 (N_13060,N_12330,N_12282);
nand U13061 (N_13061,N_12594,N_12313);
or U13062 (N_13062,N_12036,N_12209);
xnor U13063 (N_13063,N_12493,N_12235);
nand U13064 (N_13064,N_12391,N_12027);
and U13065 (N_13065,N_12376,N_12469);
nand U13066 (N_13066,N_12581,N_12267);
nor U13067 (N_13067,N_12481,N_12559);
xnor U13068 (N_13068,N_12207,N_12572);
nor U13069 (N_13069,N_12249,N_12343);
or U13070 (N_13070,N_12312,N_12477);
xor U13071 (N_13071,N_12287,N_12229);
nor U13072 (N_13072,N_12440,N_12385);
nand U13073 (N_13073,N_12477,N_12304);
or U13074 (N_13074,N_12304,N_12543);
and U13075 (N_13075,N_12238,N_12573);
nor U13076 (N_13076,N_12178,N_12513);
nor U13077 (N_13077,N_12225,N_12060);
and U13078 (N_13078,N_12579,N_12535);
nor U13079 (N_13079,N_12049,N_12352);
or U13080 (N_13080,N_12450,N_12067);
xnor U13081 (N_13081,N_12058,N_12513);
and U13082 (N_13082,N_12524,N_12591);
nor U13083 (N_13083,N_12004,N_12233);
or U13084 (N_13084,N_12035,N_12127);
and U13085 (N_13085,N_12383,N_12197);
nand U13086 (N_13086,N_12524,N_12131);
nor U13087 (N_13087,N_12151,N_12285);
nor U13088 (N_13088,N_12044,N_12109);
nand U13089 (N_13089,N_12291,N_12577);
nand U13090 (N_13090,N_12341,N_12329);
or U13091 (N_13091,N_12273,N_12513);
and U13092 (N_13092,N_12478,N_12218);
and U13093 (N_13093,N_12362,N_12129);
xnor U13094 (N_13094,N_12025,N_12484);
xnor U13095 (N_13095,N_12070,N_12528);
and U13096 (N_13096,N_12597,N_12117);
xnor U13097 (N_13097,N_12100,N_12284);
xor U13098 (N_13098,N_12523,N_12516);
xor U13099 (N_13099,N_12075,N_12448);
nand U13100 (N_13100,N_12559,N_12178);
xnor U13101 (N_13101,N_12502,N_12014);
nor U13102 (N_13102,N_12217,N_12107);
and U13103 (N_13103,N_12430,N_12528);
nand U13104 (N_13104,N_12599,N_12492);
xor U13105 (N_13105,N_12538,N_12142);
and U13106 (N_13106,N_12053,N_12596);
nor U13107 (N_13107,N_12494,N_12081);
nor U13108 (N_13108,N_12109,N_12383);
and U13109 (N_13109,N_12345,N_12504);
or U13110 (N_13110,N_12218,N_12081);
nand U13111 (N_13111,N_12377,N_12285);
or U13112 (N_13112,N_12551,N_12294);
or U13113 (N_13113,N_12531,N_12243);
xnor U13114 (N_13114,N_12376,N_12033);
nor U13115 (N_13115,N_12294,N_12313);
nor U13116 (N_13116,N_12081,N_12370);
nor U13117 (N_13117,N_12002,N_12053);
nor U13118 (N_13118,N_12074,N_12459);
xor U13119 (N_13119,N_12032,N_12556);
xnor U13120 (N_13120,N_12169,N_12594);
or U13121 (N_13121,N_12095,N_12039);
nor U13122 (N_13122,N_12040,N_12559);
and U13123 (N_13123,N_12150,N_12149);
or U13124 (N_13124,N_12095,N_12177);
nor U13125 (N_13125,N_12315,N_12565);
nor U13126 (N_13126,N_12183,N_12460);
nor U13127 (N_13127,N_12375,N_12482);
nand U13128 (N_13128,N_12234,N_12100);
nand U13129 (N_13129,N_12479,N_12406);
nand U13130 (N_13130,N_12036,N_12134);
xnor U13131 (N_13131,N_12089,N_12335);
nor U13132 (N_13132,N_12319,N_12582);
nand U13133 (N_13133,N_12297,N_12457);
or U13134 (N_13134,N_12023,N_12402);
nand U13135 (N_13135,N_12332,N_12100);
and U13136 (N_13136,N_12348,N_12240);
or U13137 (N_13137,N_12001,N_12029);
or U13138 (N_13138,N_12245,N_12041);
and U13139 (N_13139,N_12190,N_12157);
nor U13140 (N_13140,N_12276,N_12045);
nor U13141 (N_13141,N_12249,N_12188);
and U13142 (N_13142,N_12268,N_12248);
or U13143 (N_13143,N_12004,N_12141);
or U13144 (N_13144,N_12089,N_12111);
nand U13145 (N_13145,N_12032,N_12402);
and U13146 (N_13146,N_12165,N_12437);
nand U13147 (N_13147,N_12461,N_12437);
nand U13148 (N_13148,N_12196,N_12119);
xor U13149 (N_13149,N_12417,N_12592);
xor U13150 (N_13150,N_12164,N_12341);
or U13151 (N_13151,N_12208,N_12278);
xnor U13152 (N_13152,N_12018,N_12260);
nor U13153 (N_13153,N_12468,N_12013);
nand U13154 (N_13154,N_12175,N_12120);
xnor U13155 (N_13155,N_12175,N_12201);
nor U13156 (N_13156,N_12004,N_12577);
or U13157 (N_13157,N_12284,N_12012);
nand U13158 (N_13158,N_12498,N_12092);
nand U13159 (N_13159,N_12152,N_12422);
and U13160 (N_13160,N_12108,N_12488);
xor U13161 (N_13161,N_12250,N_12500);
nor U13162 (N_13162,N_12016,N_12022);
nor U13163 (N_13163,N_12544,N_12488);
xor U13164 (N_13164,N_12180,N_12218);
nand U13165 (N_13165,N_12298,N_12018);
xnor U13166 (N_13166,N_12322,N_12234);
and U13167 (N_13167,N_12064,N_12191);
nand U13168 (N_13168,N_12380,N_12189);
nor U13169 (N_13169,N_12483,N_12036);
or U13170 (N_13170,N_12455,N_12542);
or U13171 (N_13171,N_12177,N_12396);
and U13172 (N_13172,N_12026,N_12333);
xnor U13173 (N_13173,N_12110,N_12087);
or U13174 (N_13174,N_12084,N_12507);
and U13175 (N_13175,N_12423,N_12508);
xnor U13176 (N_13176,N_12462,N_12250);
nand U13177 (N_13177,N_12101,N_12335);
or U13178 (N_13178,N_12220,N_12274);
or U13179 (N_13179,N_12281,N_12566);
and U13180 (N_13180,N_12570,N_12015);
and U13181 (N_13181,N_12035,N_12182);
and U13182 (N_13182,N_12549,N_12470);
nand U13183 (N_13183,N_12261,N_12219);
and U13184 (N_13184,N_12398,N_12432);
nor U13185 (N_13185,N_12001,N_12586);
xor U13186 (N_13186,N_12159,N_12201);
nor U13187 (N_13187,N_12511,N_12501);
xor U13188 (N_13188,N_12004,N_12213);
nor U13189 (N_13189,N_12414,N_12107);
nand U13190 (N_13190,N_12440,N_12330);
nand U13191 (N_13191,N_12375,N_12342);
xnor U13192 (N_13192,N_12577,N_12468);
nor U13193 (N_13193,N_12466,N_12366);
or U13194 (N_13194,N_12436,N_12393);
xor U13195 (N_13195,N_12438,N_12421);
nand U13196 (N_13196,N_12552,N_12190);
nor U13197 (N_13197,N_12111,N_12535);
or U13198 (N_13198,N_12386,N_12547);
nand U13199 (N_13199,N_12013,N_12430);
nor U13200 (N_13200,N_12624,N_12783);
xnor U13201 (N_13201,N_12675,N_12886);
nand U13202 (N_13202,N_13028,N_12643);
or U13203 (N_13203,N_12664,N_12666);
nand U13204 (N_13204,N_13167,N_12665);
nor U13205 (N_13205,N_12977,N_12797);
nand U13206 (N_13206,N_12689,N_12895);
nand U13207 (N_13207,N_13160,N_12924);
nand U13208 (N_13208,N_12639,N_12874);
and U13209 (N_13209,N_13018,N_13199);
or U13210 (N_13210,N_13020,N_12626);
or U13211 (N_13211,N_13008,N_12962);
nand U13212 (N_13212,N_13176,N_12775);
nor U13213 (N_13213,N_12949,N_12673);
nor U13214 (N_13214,N_13090,N_13050);
or U13215 (N_13215,N_12873,N_13148);
nand U13216 (N_13216,N_12835,N_12700);
nor U13217 (N_13217,N_12885,N_12697);
and U13218 (N_13218,N_12632,N_13197);
and U13219 (N_13219,N_12703,N_12820);
nor U13220 (N_13220,N_12779,N_12988);
or U13221 (N_13221,N_12630,N_13045);
or U13222 (N_13222,N_12945,N_12832);
xor U13223 (N_13223,N_13052,N_12781);
or U13224 (N_13224,N_12684,N_13185);
xnor U13225 (N_13225,N_12996,N_13125);
xnor U13226 (N_13226,N_12909,N_12602);
or U13227 (N_13227,N_12829,N_13066);
nand U13228 (N_13228,N_13130,N_13123);
nor U13229 (N_13229,N_12989,N_13055);
and U13230 (N_13230,N_13117,N_12894);
xnor U13231 (N_13231,N_13101,N_12869);
nand U13232 (N_13232,N_13108,N_13021);
nand U13233 (N_13233,N_13150,N_13189);
or U13234 (N_13234,N_12899,N_12991);
xnor U13235 (N_13235,N_13048,N_13103);
or U13236 (N_13236,N_12870,N_13057);
or U13237 (N_13237,N_12745,N_13182);
and U13238 (N_13238,N_13105,N_12738);
xnor U13239 (N_13239,N_12857,N_12970);
xnor U13240 (N_13240,N_12711,N_12735);
xnor U13241 (N_13241,N_12682,N_13067);
nand U13242 (N_13242,N_12640,N_12696);
xor U13243 (N_13243,N_12645,N_12903);
nand U13244 (N_13244,N_12985,N_12938);
xor U13245 (N_13245,N_12678,N_13064);
or U13246 (N_13246,N_12880,N_13091);
or U13247 (N_13247,N_12720,N_13035);
nor U13248 (N_13248,N_12633,N_13120);
nand U13249 (N_13249,N_12758,N_13177);
and U13250 (N_13250,N_12651,N_12688);
nand U13251 (N_13251,N_13168,N_12919);
nor U13252 (N_13252,N_13071,N_13163);
nor U13253 (N_13253,N_13190,N_13136);
nor U13254 (N_13254,N_12957,N_12722);
nand U13255 (N_13255,N_12963,N_12744);
and U13256 (N_13256,N_13157,N_12943);
xnor U13257 (N_13257,N_12809,N_13068);
nand U13258 (N_13258,N_12824,N_13063);
nand U13259 (N_13259,N_13142,N_12853);
or U13260 (N_13260,N_12828,N_12601);
or U13261 (N_13261,N_13011,N_12992);
and U13262 (N_13262,N_12661,N_12997);
xnor U13263 (N_13263,N_12913,N_12763);
or U13264 (N_13264,N_12891,N_13037);
and U13265 (N_13265,N_12721,N_13043);
xor U13266 (N_13266,N_13039,N_12770);
and U13267 (N_13267,N_12803,N_12768);
nor U13268 (N_13268,N_12612,N_12852);
and U13269 (N_13269,N_12851,N_13187);
xor U13270 (N_13270,N_12685,N_12608);
or U13271 (N_13271,N_12847,N_12769);
and U13272 (N_13272,N_12937,N_12946);
nor U13273 (N_13273,N_12817,N_12707);
or U13274 (N_13274,N_12975,N_13022);
nand U13275 (N_13275,N_12955,N_12887);
or U13276 (N_13276,N_12756,N_12843);
nor U13277 (N_13277,N_13001,N_12863);
nand U13278 (N_13278,N_13088,N_13026);
or U13279 (N_13279,N_12858,N_12905);
and U13280 (N_13280,N_12623,N_12849);
xor U13281 (N_13281,N_13155,N_12939);
xnor U13282 (N_13282,N_13195,N_12927);
nor U13283 (N_13283,N_12680,N_13181);
xnor U13284 (N_13284,N_13113,N_13129);
xor U13285 (N_13285,N_12699,N_12944);
nand U13286 (N_13286,N_12833,N_12622);
and U13287 (N_13287,N_13072,N_13191);
nor U13288 (N_13288,N_12967,N_12830);
nand U13289 (N_13289,N_12751,N_12733);
nand U13290 (N_13290,N_12686,N_12875);
or U13291 (N_13291,N_12649,N_12998);
or U13292 (N_13292,N_12627,N_12710);
or U13293 (N_13293,N_12951,N_13070);
nand U13294 (N_13294,N_12877,N_12774);
xnor U13295 (N_13295,N_13034,N_13134);
and U13296 (N_13296,N_13078,N_12636);
xnor U13297 (N_13297,N_12979,N_13042);
xnor U13298 (N_13298,N_12901,N_12804);
or U13299 (N_13299,N_13178,N_13075);
nand U13300 (N_13300,N_13016,N_12719);
nor U13301 (N_13301,N_13077,N_12658);
and U13302 (N_13302,N_12637,N_12753);
and U13303 (N_13303,N_12671,N_13116);
xor U13304 (N_13304,N_12819,N_12629);
xnor U13305 (N_13305,N_13127,N_13100);
nor U13306 (N_13306,N_12916,N_12872);
or U13307 (N_13307,N_13061,N_12790);
nor U13308 (N_13308,N_13076,N_12978);
nor U13309 (N_13309,N_12906,N_12915);
and U13310 (N_13310,N_12952,N_12902);
xor U13311 (N_13311,N_12926,N_12865);
nor U13312 (N_13312,N_12812,N_13121);
nor U13313 (N_13313,N_12876,N_12948);
nand U13314 (N_13314,N_12907,N_13166);
and U13315 (N_13315,N_12814,N_13053);
or U13316 (N_13316,N_13193,N_13014);
or U13317 (N_13317,N_12652,N_12785);
or U13318 (N_13318,N_12752,N_13173);
nor U13319 (N_13319,N_13186,N_13084);
nand U13320 (N_13320,N_13031,N_12610);
or U13321 (N_13321,N_12815,N_12780);
xnor U13322 (N_13322,N_12904,N_12844);
and U13323 (N_13323,N_13004,N_12917);
and U13324 (N_13324,N_13161,N_13169);
or U13325 (N_13325,N_12846,N_13165);
and U13326 (N_13326,N_12896,N_12972);
or U13327 (N_13327,N_13183,N_12777);
nand U13328 (N_13328,N_12766,N_12914);
or U13329 (N_13329,N_12648,N_13119);
nor U13330 (N_13330,N_13089,N_13162);
and U13331 (N_13331,N_13097,N_13102);
xnor U13332 (N_13332,N_12806,N_13056);
and U13333 (N_13333,N_12642,N_13051);
and U13334 (N_13334,N_12826,N_13188);
and U13335 (N_13335,N_12701,N_13128);
xor U13336 (N_13336,N_12940,N_12726);
nor U13337 (N_13337,N_13096,N_13094);
nand U13338 (N_13338,N_12981,N_13025);
or U13339 (N_13339,N_12741,N_12838);
or U13340 (N_13340,N_12805,N_12708);
xnor U13341 (N_13341,N_12653,N_12793);
and U13342 (N_13342,N_13083,N_12947);
xnor U13343 (N_13343,N_12897,N_12757);
nand U13344 (N_13344,N_12728,N_13138);
xor U13345 (N_13345,N_12729,N_12739);
or U13346 (N_13346,N_12882,N_13159);
nor U13347 (N_13347,N_13062,N_12725);
nand U13348 (N_13348,N_13137,N_12736);
and U13349 (N_13349,N_13087,N_12811);
or U13350 (N_13350,N_13118,N_13005);
xor U13351 (N_13351,N_12836,N_12717);
nand U13352 (N_13352,N_12816,N_12754);
nand U13353 (N_13353,N_12966,N_12922);
or U13354 (N_13354,N_12848,N_12615);
xor U13355 (N_13355,N_12784,N_13184);
nor U13356 (N_13356,N_12614,N_12990);
and U13357 (N_13357,N_13093,N_12714);
or U13358 (N_13358,N_13000,N_12954);
nand U13359 (N_13359,N_12950,N_12831);
nand U13360 (N_13360,N_12823,N_12737);
or U13361 (N_13361,N_13106,N_13111);
or U13362 (N_13362,N_13192,N_13170);
or U13363 (N_13363,N_12698,N_13143);
nor U13364 (N_13364,N_12837,N_12931);
nand U13365 (N_13365,N_12867,N_12965);
xnor U13366 (N_13366,N_12794,N_13012);
or U13367 (N_13367,N_12659,N_12799);
xor U13368 (N_13368,N_13131,N_12859);
nor U13369 (N_13369,N_12881,N_12702);
xnor U13370 (N_13370,N_12605,N_12968);
nor U13371 (N_13371,N_13036,N_12760);
nand U13372 (N_13372,N_13158,N_12980);
and U13373 (N_13373,N_12868,N_13074);
xor U13374 (N_13374,N_12713,N_12692);
or U13375 (N_13375,N_13114,N_12613);
xnor U13376 (N_13376,N_13041,N_12618);
nor U13377 (N_13377,N_12861,N_12617);
or U13378 (N_13378,N_12860,N_12842);
nor U13379 (N_13379,N_13086,N_12734);
nor U13380 (N_13380,N_12864,N_13098);
nor U13381 (N_13381,N_12893,N_12724);
nor U13382 (N_13382,N_13149,N_12767);
or U13383 (N_13383,N_13141,N_12929);
nor U13384 (N_13384,N_12941,N_12986);
and U13385 (N_13385,N_13135,N_13017);
or U13386 (N_13386,N_12670,N_12772);
and U13387 (N_13387,N_12663,N_12961);
nand U13388 (N_13388,N_12727,N_12856);
xor U13389 (N_13389,N_12789,N_12732);
xnor U13390 (N_13390,N_13095,N_12810);
xnor U13391 (N_13391,N_12807,N_12956);
xnor U13392 (N_13392,N_12890,N_12813);
nand U13393 (N_13393,N_12761,N_12934);
nand U13394 (N_13394,N_12620,N_12616);
xnor U13395 (N_13395,N_13110,N_13099);
nor U13396 (N_13396,N_13019,N_12987);
nor U13397 (N_13397,N_12668,N_12973);
xor U13398 (N_13398,N_12958,N_12695);
nor U13399 (N_13399,N_12604,N_12969);
nor U13400 (N_13400,N_12788,N_12834);
nor U13401 (N_13401,N_12884,N_13081);
nor U13402 (N_13402,N_12638,N_13082);
or U13403 (N_13403,N_13024,N_13171);
or U13404 (N_13404,N_12776,N_13079);
or U13405 (N_13405,N_12839,N_13196);
nand U13406 (N_13406,N_12762,N_12621);
nand U13407 (N_13407,N_12693,N_12995);
xnor U13408 (N_13408,N_12748,N_12764);
or U13409 (N_13409,N_12676,N_12889);
nor U13410 (N_13410,N_13151,N_13049);
or U13411 (N_13411,N_12959,N_12999);
and U13412 (N_13412,N_12641,N_13174);
nand U13413 (N_13413,N_12694,N_12964);
nand U13414 (N_13414,N_12912,N_13133);
xor U13415 (N_13415,N_13030,N_12821);
and U13416 (N_13416,N_12827,N_12611);
or U13417 (N_13417,N_13115,N_12681);
and U13418 (N_13418,N_12647,N_12953);
xnor U13419 (N_13419,N_12960,N_12749);
xor U13420 (N_13420,N_13013,N_12936);
nand U13421 (N_13421,N_12845,N_12984);
nor U13422 (N_13422,N_12606,N_13126);
or U13423 (N_13423,N_12609,N_12921);
and U13424 (N_13424,N_12778,N_13069);
and U13425 (N_13425,N_12866,N_12910);
nor U13426 (N_13426,N_13059,N_12660);
nand U13427 (N_13427,N_13060,N_13107);
xor U13428 (N_13428,N_12712,N_12669);
xnor U13429 (N_13429,N_13154,N_13085);
nor U13430 (N_13430,N_13145,N_13146);
nand U13431 (N_13431,N_13175,N_12918);
or U13432 (N_13432,N_13179,N_12715);
nor U13433 (N_13433,N_13033,N_12787);
or U13434 (N_13434,N_12705,N_12709);
nor U13435 (N_13435,N_12878,N_13080);
nor U13436 (N_13436,N_12600,N_12855);
nand U13437 (N_13437,N_12607,N_12801);
nand U13438 (N_13438,N_12656,N_12840);
and U13439 (N_13439,N_12932,N_12928);
and U13440 (N_13440,N_13194,N_12750);
or U13441 (N_13441,N_12976,N_12730);
nand U13442 (N_13442,N_12971,N_13023);
or U13443 (N_13443,N_13002,N_12646);
and U13444 (N_13444,N_13032,N_12898);
or U13445 (N_13445,N_12796,N_12672);
and U13446 (N_13446,N_12631,N_13152);
nand U13447 (N_13447,N_13003,N_12743);
xor U13448 (N_13448,N_12759,N_12900);
nand U13449 (N_13449,N_13038,N_12718);
and U13450 (N_13450,N_12786,N_12818);
or U13451 (N_13451,N_13164,N_13065);
nand U13452 (N_13452,N_12841,N_12771);
nand U13453 (N_13453,N_12691,N_12795);
xor U13454 (N_13454,N_13172,N_12603);
xor U13455 (N_13455,N_12747,N_12782);
nand U13456 (N_13456,N_13147,N_12644);
nand U13457 (N_13457,N_13104,N_12683);
nand U13458 (N_13458,N_12862,N_12908);
nor U13459 (N_13459,N_12679,N_13006);
nand U13460 (N_13460,N_12723,N_13144);
xor U13461 (N_13461,N_12704,N_13015);
nand U13462 (N_13462,N_13139,N_12755);
nor U13463 (N_13463,N_13047,N_12930);
nor U13464 (N_13464,N_12808,N_12993);
and U13465 (N_13465,N_13122,N_12706);
nand U13466 (N_13466,N_12740,N_12650);
nor U13467 (N_13467,N_13027,N_12925);
or U13468 (N_13468,N_12742,N_12635);
xor U13469 (N_13469,N_13044,N_12667);
xor U13470 (N_13470,N_13007,N_13040);
xor U13471 (N_13471,N_12765,N_13073);
or U13472 (N_13472,N_12674,N_13112);
and U13473 (N_13473,N_12920,N_12942);
or U13474 (N_13474,N_13046,N_13058);
and U13475 (N_13475,N_12791,N_12687);
nor U13476 (N_13476,N_12994,N_12690);
nor U13477 (N_13477,N_12822,N_13198);
nand U13478 (N_13478,N_12892,N_12677);
nand U13479 (N_13479,N_13132,N_12974);
and U13480 (N_13480,N_13156,N_13029);
nor U13481 (N_13481,N_13009,N_12628);
or U13482 (N_13482,N_12655,N_12731);
or U13483 (N_13483,N_13054,N_12850);
nand U13484 (N_13484,N_12657,N_13109);
nand U13485 (N_13485,N_12933,N_12888);
xnor U13486 (N_13486,N_12923,N_13010);
and U13487 (N_13487,N_12619,N_12800);
and U13488 (N_13488,N_12716,N_12983);
or U13489 (N_13489,N_12911,N_12879);
nand U13490 (N_13490,N_12883,N_12802);
or U13491 (N_13491,N_12982,N_12798);
nand U13492 (N_13492,N_12746,N_12662);
and U13493 (N_13493,N_13092,N_12935);
nor U13494 (N_13494,N_12634,N_12871);
nand U13495 (N_13495,N_12825,N_12792);
and U13496 (N_13496,N_12773,N_12854);
or U13497 (N_13497,N_13124,N_13180);
or U13498 (N_13498,N_12625,N_12654);
or U13499 (N_13499,N_13153,N_13140);
nor U13500 (N_13500,N_13187,N_13082);
nor U13501 (N_13501,N_12972,N_12727);
xor U13502 (N_13502,N_12729,N_12918);
nand U13503 (N_13503,N_12704,N_13113);
and U13504 (N_13504,N_13123,N_12916);
nor U13505 (N_13505,N_12832,N_12606);
nand U13506 (N_13506,N_13132,N_12666);
nor U13507 (N_13507,N_13158,N_12890);
nand U13508 (N_13508,N_12826,N_12841);
or U13509 (N_13509,N_12896,N_13028);
xnor U13510 (N_13510,N_12683,N_12779);
nor U13511 (N_13511,N_12627,N_12605);
or U13512 (N_13512,N_12886,N_13166);
nor U13513 (N_13513,N_12761,N_12893);
nor U13514 (N_13514,N_12749,N_12698);
nor U13515 (N_13515,N_12892,N_12807);
and U13516 (N_13516,N_13045,N_12949);
nand U13517 (N_13517,N_12898,N_13124);
or U13518 (N_13518,N_12713,N_12960);
nor U13519 (N_13519,N_13021,N_12762);
or U13520 (N_13520,N_12887,N_13066);
xor U13521 (N_13521,N_13140,N_12936);
nand U13522 (N_13522,N_12687,N_12720);
and U13523 (N_13523,N_12977,N_13146);
and U13524 (N_13524,N_13123,N_12911);
nand U13525 (N_13525,N_12713,N_12685);
and U13526 (N_13526,N_12872,N_12818);
xnor U13527 (N_13527,N_12883,N_12669);
and U13528 (N_13528,N_12678,N_12847);
nor U13529 (N_13529,N_12628,N_12838);
or U13530 (N_13530,N_13000,N_12784);
nand U13531 (N_13531,N_13057,N_12714);
nor U13532 (N_13532,N_12920,N_12617);
nor U13533 (N_13533,N_13140,N_12797);
or U13534 (N_13534,N_12641,N_12853);
nor U13535 (N_13535,N_13012,N_12876);
or U13536 (N_13536,N_12738,N_13097);
nor U13537 (N_13537,N_12991,N_12973);
xor U13538 (N_13538,N_12643,N_12919);
nor U13539 (N_13539,N_13048,N_13110);
xor U13540 (N_13540,N_12611,N_13002);
or U13541 (N_13541,N_12979,N_12948);
nand U13542 (N_13542,N_13076,N_12847);
or U13543 (N_13543,N_12931,N_12750);
or U13544 (N_13544,N_12781,N_13089);
or U13545 (N_13545,N_12920,N_13035);
xnor U13546 (N_13546,N_12991,N_12789);
and U13547 (N_13547,N_12633,N_13189);
nor U13548 (N_13548,N_12628,N_12859);
nor U13549 (N_13549,N_12799,N_12838);
nand U13550 (N_13550,N_13101,N_13164);
nor U13551 (N_13551,N_12793,N_12868);
xnor U13552 (N_13552,N_12762,N_12771);
nor U13553 (N_13553,N_12922,N_12973);
or U13554 (N_13554,N_12954,N_12641);
and U13555 (N_13555,N_13039,N_12915);
nand U13556 (N_13556,N_13076,N_13159);
or U13557 (N_13557,N_13074,N_12742);
nor U13558 (N_13558,N_13010,N_12656);
and U13559 (N_13559,N_12742,N_12912);
and U13560 (N_13560,N_12690,N_12738);
or U13561 (N_13561,N_12896,N_13048);
nand U13562 (N_13562,N_12938,N_13157);
nand U13563 (N_13563,N_12707,N_13107);
or U13564 (N_13564,N_13062,N_13174);
and U13565 (N_13565,N_12996,N_13166);
nand U13566 (N_13566,N_13142,N_12653);
and U13567 (N_13567,N_12776,N_12878);
or U13568 (N_13568,N_13196,N_12677);
nand U13569 (N_13569,N_13079,N_12844);
and U13570 (N_13570,N_12772,N_12948);
nor U13571 (N_13571,N_12946,N_13074);
xnor U13572 (N_13572,N_13177,N_12980);
xor U13573 (N_13573,N_12943,N_12619);
or U13574 (N_13574,N_12953,N_13129);
and U13575 (N_13575,N_12663,N_12784);
nor U13576 (N_13576,N_12603,N_12807);
or U13577 (N_13577,N_13178,N_12966);
and U13578 (N_13578,N_12938,N_13020);
or U13579 (N_13579,N_12752,N_12836);
xnor U13580 (N_13580,N_13139,N_12961);
or U13581 (N_13581,N_13041,N_13198);
nor U13582 (N_13582,N_12972,N_12946);
and U13583 (N_13583,N_13159,N_12774);
xnor U13584 (N_13584,N_12763,N_12667);
xor U13585 (N_13585,N_12912,N_12947);
nand U13586 (N_13586,N_13011,N_13166);
xor U13587 (N_13587,N_12700,N_12622);
or U13588 (N_13588,N_13032,N_12989);
and U13589 (N_13589,N_13054,N_12683);
nor U13590 (N_13590,N_13144,N_12623);
nor U13591 (N_13591,N_12781,N_12805);
or U13592 (N_13592,N_12875,N_13095);
nor U13593 (N_13593,N_12764,N_13060);
nor U13594 (N_13594,N_12663,N_13174);
nand U13595 (N_13595,N_12720,N_12809);
and U13596 (N_13596,N_12944,N_12701);
nor U13597 (N_13597,N_13035,N_12682);
nor U13598 (N_13598,N_12977,N_12871);
or U13599 (N_13599,N_12997,N_12742);
nor U13600 (N_13600,N_13187,N_12992);
xnor U13601 (N_13601,N_13186,N_12628);
xnor U13602 (N_13602,N_12722,N_12647);
xor U13603 (N_13603,N_12748,N_12870);
or U13604 (N_13604,N_13177,N_12765);
xor U13605 (N_13605,N_12731,N_12810);
or U13606 (N_13606,N_12777,N_13075);
xnor U13607 (N_13607,N_12805,N_13183);
nor U13608 (N_13608,N_13023,N_13145);
xor U13609 (N_13609,N_13190,N_13106);
and U13610 (N_13610,N_13067,N_12721);
xor U13611 (N_13611,N_13179,N_12872);
and U13612 (N_13612,N_12846,N_13029);
and U13613 (N_13613,N_13087,N_12820);
xnor U13614 (N_13614,N_12983,N_13180);
xnor U13615 (N_13615,N_12969,N_13185);
xnor U13616 (N_13616,N_12953,N_12792);
nor U13617 (N_13617,N_13172,N_12746);
and U13618 (N_13618,N_12670,N_12863);
or U13619 (N_13619,N_12782,N_12862);
or U13620 (N_13620,N_13006,N_13088);
nor U13621 (N_13621,N_12648,N_12964);
and U13622 (N_13622,N_13150,N_13080);
or U13623 (N_13623,N_12979,N_13091);
nand U13624 (N_13624,N_13058,N_12905);
nand U13625 (N_13625,N_13151,N_12831);
nor U13626 (N_13626,N_13022,N_12789);
xnor U13627 (N_13627,N_12629,N_12719);
xor U13628 (N_13628,N_12879,N_12651);
nor U13629 (N_13629,N_12764,N_13012);
and U13630 (N_13630,N_12785,N_12776);
xor U13631 (N_13631,N_12665,N_12872);
xor U13632 (N_13632,N_12752,N_12936);
nand U13633 (N_13633,N_13080,N_12635);
nor U13634 (N_13634,N_13070,N_12772);
or U13635 (N_13635,N_12841,N_13101);
xor U13636 (N_13636,N_12880,N_12726);
nand U13637 (N_13637,N_12875,N_12991);
nor U13638 (N_13638,N_12991,N_12841);
xnor U13639 (N_13639,N_12847,N_12832);
nand U13640 (N_13640,N_12622,N_13068);
or U13641 (N_13641,N_13031,N_12749);
xor U13642 (N_13642,N_12838,N_13009);
nand U13643 (N_13643,N_13041,N_12924);
and U13644 (N_13644,N_13006,N_13159);
and U13645 (N_13645,N_12751,N_12634);
nor U13646 (N_13646,N_12803,N_12663);
nand U13647 (N_13647,N_12796,N_13158);
or U13648 (N_13648,N_13032,N_12823);
nand U13649 (N_13649,N_12622,N_13055);
and U13650 (N_13650,N_12964,N_12971);
or U13651 (N_13651,N_12866,N_13065);
and U13652 (N_13652,N_12780,N_12854);
nor U13653 (N_13653,N_13130,N_13027);
nor U13654 (N_13654,N_12681,N_12685);
xnor U13655 (N_13655,N_12625,N_12704);
xor U13656 (N_13656,N_12995,N_13116);
nand U13657 (N_13657,N_13024,N_12611);
nor U13658 (N_13658,N_12826,N_12956);
xor U13659 (N_13659,N_13070,N_13092);
or U13660 (N_13660,N_12763,N_12754);
nand U13661 (N_13661,N_13064,N_12625);
nor U13662 (N_13662,N_12686,N_13063);
nand U13663 (N_13663,N_13043,N_13081);
xnor U13664 (N_13664,N_13064,N_13097);
nand U13665 (N_13665,N_12931,N_12955);
or U13666 (N_13666,N_13100,N_12979);
or U13667 (N_13667,N_12817,N_12813);
xor U13668 (N_13668,N_13109,N_12651);
or U13669 (N_13669,N_12792,N_12846);
nor U13670 (N_13670,N_12797,N_12942);
or U13671 (N_13671,N_13011,N_12935);
nand U13672 (N_13672,N_12942,N_12683);
and U13673 (N_13673,N_12891,N_12757);
xnor U13674 (N_13674,N_12827,N_13073);
xnor U13675 (N_13675,N_12760,N_12919);
xor U13676 (N_13676,N_12724,N_13126);
nand U13677 (N_13677,N_12895,N_12901);
xor U13678 (N_13678,N_12603,N_12783);
xor U13679 (N_13679,N_12905,N_12902);
and U13680 (N_13680,N_13154,N_13174);
nand U13681 (N_13681,N_13053,N_12774);
nand U13682 (N_13682,N_12726,N_12902);
and U13683 (N_13683,N_13011,N_13035);
xor U13684 (N_13684,N_12938,N_12615);
nor U13685 (N_13685,N_13099,N_13184);
nor U13686 (N_13686,N_13065,N_12975);
nand U13687 (N_13687,N_12863,N_13192);
xor U13688 (N_13688,N_13036,N_13115);
nand U13689 (N_13689,N_13166,N_12993);
nor U13690 (N_13690,N_12754,N_13039);
nand U13691 (N_13691,N_12612,N_13050);
nor U13692 (N_13692,N_12749,N_12670);
xnor U13693 (N_13693,N_12637,N_13113);
or U13694 (N_13694,N_12836,N_12901);
or U13695 (N_13695,N_13004,N_12765);
nand U13696 (N_13696,N_12844,N_12863);
nand U13697 (N_13697,N_12687,N_12834);
nand U13698 (N_13698,N_12736,N_12965);
xor U13699 (N_13699,N_12706,N_13173);
nor U13700 (N_13700,N_12651,N_12647);
or U13701 (N_13701,N_13069,N_12917);
and U13702 (N_13702,N_13071,N_12734);
nor U13703 (N_13703,N_13012,N_12606);
nor U13704 (N_13704,N_12868,N_13043);
nand U13705 (N_13705,N_12927,N_12640);
or U13706 (N_13706,N_12682,N_13078);
and U13707 (N_13707,N_12808,N_12634);
or U13708 (N_13708,N_12719,N_12922);
and U13709 (N_13709,N_12728,N_13081);
xor U13710 (N_13710,N_12785,N_12806);
nand U13711 (N_13711,N_12756,N_12830);
or U13712 (N_13712,N_13122,N_13105);
xnor U13713 (N_13713,N_12667,N_13198);
nand U13714 (N_13714,N_13048,N_12846);
xnor U13715 (N_13715,N_12865,N_13134);
xnor U13716 (N_13716,N_12728,N_12601);
xor U13717 (N_13717,N_13000,N_12624);
nand U13718 (N_13718,N_13190,N_12653);
or U13719 (N_13719,N_13137,N_13124);
or U13720 (N_13720,N_13146,N_13034);
xnor U13721 (N_13721,N_12624,N_13145);
or U13722 (N_13722,N_13000,N_12732);
xor U13723 (N_13723,N_12773,N_12631);
nand U13724 (N_13724,N_12761,N_12750);
nand U13725 (N_13725,N_12924,N_13012);
nor U13726 (N_13726,N_12984,N_13179);
xor U13727 (N_13727,N_12964,N_12935);
or U13728 (N_13728,N_12794,N_13047);
nor U13729 (N_13729,N_13019,N_12959);
and U13730 (N_13730,N_13051,N_13014);
and U13731 (N_13731,N_13000,N_13120);
nor U13732 (N_13732,N_12633,N_12649);
nor U13733 (N_13733,N_13106,N_13069);
and U13734 (N_13734,N_12697,N_13189);
and U13735 (N_13735,N_12795,N_12881);
nand U13736 (N_13736,N_12925,N_12624);
nor U13737 (N_13737,N_12719,N_13035);
and U13738 (N_13738,N_13061,N_12791);
nand U13739 (N_13739,N_13025,N_12741);
and U13740 (N_13740,N_12749,N_12707);
xor U13741 (N_13741,N_12934,N_12854);
and U13742 (N_13742,N_12684,N_12828);
nor U13743 (N_13743,N_13127,N_13085);
nor U13744 (N_13744,N_13178,N_12606);
or U13745 (N_13745,N_12616,N_12830);
xor U13746 (N_13746,N_12961,N_12845);
and U13747 (N_13747,N_12917,N_12940);
and U13748 (N_13748,N_12734,N_13072);
and U13749 (N_13749,N_13017,N_13124);
or U13750 (N_13750,N_12936,N_12738);
nand U13751 (N_13751,N_12845,N_12792);
xnor U13752 (N_13752,N_12978,N_12968);
or U13753 (N_13753,N_12755,N_12805);
or U13754 (N_13754,N_12633,N_12904);
nor U13755 (N_13755,N_13099,N_12899);
and U13756 (N_13756,N_12770,N_12628);
or U13757 (N_13757,N_12936,N_12962);
and U13758 (N_13758,N_12885,N_12928);
xnor U13759 (N_13759,N_12762,N_13055);
and U13760 (N_13760,N_12715,N_12977);
nor U13761 (N_13761,N_12763,N_12792);
xor U13762 (N_13762,N_13022,N_13140);
nand U13763 (N_13763,N_12904,N_12921);
nor U13764 (N_13764,N_12884,N_12778);
xor U13765 (N_13765,N_13172,N_12696);
nor U13766 (N_13766,N_12759,N_12996);
or U13767 (N_13767,N_12676,N_12862);
and U13768 (N_13768,N_12699,N_13128);
xor U13769 (N_13769,N_12792,N_12890);
xnor U13770 (N_13770,N_13068,N_12699);
and U13771 (N_13771,N_12909,N_12888);
nor U13772 (N_13772,N_12603,N_13012);
nor U13773 (N_13773,N_12975,N_12681);
nand U13774 (N_13774,N_13054,N_12919);
xnor U13775 (N_13775,N_13190,N_12980);
or U13776 (N_13776,N_12884,N_12761);
nor U13777 (N_13777,N_13189,N_12602);
nor U13778 (N_13778,N_13129,N_13066);
nand U13779 (N_13779,N_12849,N_12853);
nor U13780 (N_13780,N_12940,N_12875);
nand U13781 (N_13781,N_12758,N_12772);
xor U13782 (N_13782,N_13112,N_13122);
or U13783 (N_13783,N_12898,N_13136);
nor U13784 (N_13784,N_13113,N_12676);
or U13785 (N_13785,N_12822,N_13013);
nand U13786 (N_13786,N_13125,N_13106);
or U13787 (N_13787,N_12793,N_12734);
nor U13788 (N_13788,N_12752,N_13017);
or U13789 (N_13789,N_12705,N_12719);
and U13790 (N_13790,N_12600,N_12928);
and U13791 (N_13791,N_12972,N_12629);
nand U13792 (N_13792,N_12916,N_13134);
and U13793 (N_13793,N_12931,N_12724);
nor U13794 (N_13794,N_12756,N_13020);
xnor U13795 (N_13795,N_12790,N_12914);
nor U13796 (N_13796,N_13161,N_13048);
and U13797 (N_13797,N_13075,N_12683);
xnor U13798 (N_13798,N_12905,N_12768);
or U13799 (N_13799,N_12823,N_12695);
or U13800 (N_13800,N_13705,N_13309);
xnor U13801 (N_13801,N_13283,N_13277);
nand U13802 (N_13802,N_13677,N_13399);
and U13803 (N_13803,N_13753,N_13560);
or U13804 (N_13804,N_13248,N_13365);
nor U13805 (N_13805,N_13566,N_13527);
nand U13806 (N_13806,N_13534,N_13230);
nand U13807 (N_13807,N_13554,N_13784);
and U13808 (N_13808,N_13726,N_13440);
nand U13809 (N_13809,N_13639,N_13235);
or U13810 (N_13810,N_13561,N_13655);
nand U13811 (N_13811,N_13492,N_13624);
nand U13812 (N_13812,N_13654,N_13638);
nor U13813 (N_13813,N_13468,N_13535);
xor U13814 (N_13814,N_13204,N_13388);
nand U13815 (N_13815,N_13360,N_13270);
or U13816 (N_13816,N_13519,N_13251);
nand U13817 (N_13817,N_13316,N_13289);
nand U13818 (N_13818,N_13462,N_13770);
or U13819 (N_13819,N_13608,N_13245);
nor U13820 (N_13820,N_13651,N_13595);
and U13821 (N_13821,N_13584,N_13363);
nand U13822 (N_13822,N_13573,N_13418);
nor U13823 (N_13823,N_13280,N_13215);
or U13824 (N_13824,N_13750,N_13776);
and U13825 (N_13825,N_13577,N_13713);
nor U13826 (N_13826,N_13323,N_13611);
xnor U13827 (N_13827,N_13241,N_13400);
nor U13828 (N_13828,N_13236,N_13412);
or U13829 (N_13829,N_13751,N_13794);
and U13830 (N_13830,N_13565,N_13327);
nor U13831 (N_13831,N_13684,N_13614);
and U13832 (N_13832,N_13719,N_13646);
nor U13833 (N_13833,N_13539,N_13580);
or U13834 (N_13834,N_13797,N_13723);
and U13835 (N_13835,N_13508,N_13387);
nand U13836 (N_13836,N_13778,N_13475);
and U13837 (N_13837,N_13469,N_13210);
nand U13838 (N_13838,N_13626,N_13273);
xnor U13839 (N_13839,N_13775,N_13504);
and U13840 (N_13840,N_13663,N_13421);
nand U13841 (N_13841,N_13693,N_13308);
and U13842 (N_13842,N_13579,N_13582);
xor U13843 (N_13843,N_13473,N_13450);
or U13844 (N_13844,N_13333,N_13668);
xor U13845 (N_13845,N_13556,N_13786);
nand U13846 (N_13846,N_13292,N_13716);
and U13847 (N_13847,N_13567,N_13518);
or U13848 (N_13848,N_13446,N_13372);
nand U13849 (N_13849,N_13540,N_13672);
nor U13850 (N_13850,N_13356,N_13417);
nand U13851 (N_13851,N_13671,N_13375);
xor U13852 (N_13852,N_13366,N_13521);
or U13853 (N_13853,N_13601,N_13688);
or U13854 (N_13854,N_13649,N_13261);
and U13855 (N_13855,N_13774,N_13335);
xnor U13856 (N_13856,N_13736,N_13414);
xnor U13857 (N_13857,N_13634,N_13267);
nand U13858 (N_13858,N_13437,N_13558);
and U13859 (N_13859,N_13741,N_13279);
xor U13860 (N_13860,N_13765,N_13218);
nand U13861 (N_13861,N_13409,N_13721);
nor U13862 (N_13862,N_13536,N_13590);
or U13863 (N_13863,N_13661,N_13201);
xnor U13864 (N_13864,N_13644,N_13452);
or U13865 (N_13865,N_13460,N_13274);
or U13866 (N_13866,N_13255,N_13404);
xnor U13867 (N_13867,N_13799,N_13773);
nand U13868 (N_13868,N_13520,N_13530);
nand U13869 (N_13869,N_13317,N_13334);
nand U13870 (N_13870,N_13740,N_13710);
xor U13871 (N_13871,N_13711,N_13636);
nor U13872 (N_13872,N_13435,N_13547);
and U13873 (N_13873,N_13406,N_13275);
nand U13874 (N_13874,N_13328,N_13393);
nand U13875 (N_13875,N_13653,N_13569);
or U13876 (N_13876,N_13550,N_13780);
nand U13877 (N_13877,N_13712,N_13208);
nor U13878 (N_13878,N_13304,N_13262);
or U13879 (N_13879,N_13330,N_13629);
and U13880 (N_13880,N_13214,N_13747);
nor U13881 (N_13881,N_13260,N_13227);
nand U13882 (N_13882,N_13683,N_13633);
nand U13883 (N_13883,N_13345,N_13500);
nor U13884 (N_13884,N_13616,N_13477);
nor U13885 (N_13885,N_13532,N_13493);
or U13886 (N_13886,N_13687,N_13746);
xnor U13887 (N_13887,N_13359,N_13542);
nand U13888 (N_13888,N_13732,N_13762);
nor U13889 (N_13889,N_13464,N_13715);
xnor U13890 (N_13890,N_13312,N_13311);
nand U13891 (N_13891,N_13205,N_13457);
xor U13892 (N_13892,N_13470,N_13781);
xnor U13893 (N_13893,N_13463,N_13298);
nand U13894 (N_13894,N_13242,N_13574);
nand U13895 (N_13895,N_13465,N_13511);
xnor U13896 (N_13896,N_13707,N_13202);
or U13897 (N_13897,N_13771,N_13240);
and U13898 (N_13898,N_13395,N_13622);
nand U13899 (N_13899,N_13225,N_13433);
nand U13900 (N_13900,N_13216,N_13320);
xnor U13901 (N_13901,N_13618,N_13660);
xor U13902 (N_13902,N_13386,N_13353);
and U13903 (N_13903,N_13695,N_13401);
and U13904 (N_13904,N_13376,N_13318);
or U13905 (N_13905,N_13594,N_13607);
nand U13906 (N_13906,N_13438,N_13495);
xnor U13907 (N_13907,N_13276,N_13354);
nor U13908 (N_13908,N_13664,N_13228);
nand U13909 (N_13909,N_13620,N_13343);
nand U13910 (N_13910,N_13602,N_13777);
and U13911 (N_13911,N_13459,N_13627);
nor U13912 (N_13912,N_13220,N_13296);
nand U13913 (N_13913,N_13321,N_13581);
nand U13914 (N_13914,N_13796,N_13458);
and U13915 (N_13915,N_13538,N_13717);
nor U13916 (N_13916,N_13411,N_13691);
or U13917 (N_13917,N_13754,N_13206);
xor U13918 (N_13918,N_13377,N_13436);
or U13919 (N_13919,N_13301,N_13730);
nor U13920 (N_13920,N_13515,N_13787);
nand U13921 (N_13921,N_13416,N_13449);
or U13922 (N_13922,N_13385,N_13383);
nand U13923 (N_13923,N_13244,N_13355);
xnor U13924 (N_13924,N_13246,N_13571);
nor U13925 (N_13925,N_13722,N_13669);
nor U13926 (N_13926,N_13505,N_13362);
and U13927 (N_13927,N_13430,N_13336);
or U13928 (N_13928,N_13352,N_13200);
xnor U13929 (N_13929,N_13303,N_13643);
nor U13930 (N_13930,N_13474,N_13631);
nor U13931 (N_13931,N_13657,N_13325);
or U13932 (N_13932,N_13517,N_13297);
or U13933 (N_13933,N_13662,N_13718);
nor U13934 (N_13934,N_13613,N_13403);
or U13935 (N_13935,N_13541,N_13442);
and U13936 (N_13936,N_13307,N_13757);
nand U13937 (N_13937,N_13300,N_13338);
nor U13938 (N_13938,N_13247,N_13702);
nand U13939 (N_13939,N_13642,N_13548);
nor U13940 (N_13940,N_13394,N_13609);
and U13941 (N_13941,N_13331,N_13391);
and U13942 (N_13942,N_13456,N_13488);
xor U13943 (N_13943,N_13531,N_13699);
xnor U13944 (N_13944,N_13454,N_13523);
nand U13945 (N_13945,N_13689,N_13340);
nand U13946 (N_13946,N_13670,N_13769);
xor U13947 (N_13947,N_13641,N_13525);
nor U13948 (N_13948,N_13708,N_13397);
or U13949 (N_13949,N_13549,N_13698);
and U13950 (N_13950,N_13645,N_13380);
nor U13951 (N_13951,N_13291,N_13322);
and U13952 (N_13952,N_13252,N_13258);
and U13953 (N_13953,N_13374,N_13281);
and U13954 (N_13954,N_13486,N_13351);
or U13955 (N_13955,N_13489,N_13451);
nor U13956 (N_13956,N_13337,N_13587);
or U13957 (N_13957,N_13231,N_13288);
nor U13958 (N_13958,N_13428,N_13226);
and U13959 (N_13959,N_13499,N_13603);
nand U13960 (N_13960,N_13744,N_13329);
nand U13961 (N_13961,N_13528,N_13219);
and U13962 (N_13962,N_13564,N_13572);
nand U13963 (N_13963,N_13426,N_13332);
nor U13964 (N_13964,N_13379,N_13271);
and U13965 (N_13965,N_13768,N_13447);
nand U13966 (N_13966,N_13686,N_13295);
and U13967 (N_13967,N_13546,N_13315);
and U13968 (N_13968,N_13306,N_13632);
nor U13969 (N_13969,N_13739,N_13339);
xnor U13970 (N_13970,N_13358,N_13563);
nor U13971 (N_13971,N_13445,N_13405);
nor U13972 (N_13972,N_13479,N_13265);
and U13973 (N_13973,N_13795,N_13585);
and U13974 (N_13974,N_13290,N_13466);
nor U13975 (N_13975,N_13763,N_13779);
xor U13976 (N_13976,N_13256,N_13396);
xnor U13977 (N_13977,N_13667,N_13413);
and U13978 (N_13978,N_13203,N_13434);
nand U13979 (N_13979,N_13368,N_13207);
and U13980 (N_13980,N_13497,N_13788);
or U13981 (N_13981,N_13266,N_13250);
or U13982 (N_13982,N_13524,N_13791);
nand U13983 (N_13983,N_13217,N_13415);
nand U13984 (N_13984,N_13709,N_13487);
xor U13985 (N_13985,N_13692,N_13344);
and U13986 (N_13986,N_13269,N_13483);
and U13987 (N_13987,N_13249,N_13658);
xnor U13988 (N_13988,N_13496,N_13761);
xnor U13989 (N_13989,N_13238,N_13284);
or U13990 (N_13990,N_13706,N_13568);
nand U13991 (N_13991,N_13342,N_13237);
nand U13992 (N_13992,N_13424,N_13472);
nor U13993 (N_13993,N_13259,N_13685);
or U13994 (N_13994,N_13738,N_13697);
nand U13995 (N_13995,N_13509,N_13526);
or U13996 (N_13996,N_13610,N_13724);
nand U13997 (N_13997,N_13224,N_13543);
nand U13998 (N_13998,N_13615,N_13731);
xnor U13999 (N_13999,N_13482,N_13302);
xnor U14000 (N_14000,N_13232,N_13478);
xor U14001 (N_14001,N_13586,N_13367);
and U14002 (N_14002,N_13756,N_13348);
or U14003 (N_14003,N_13503,N_13326);
or U14004 (N_14004,N_13553,N_13420);
xnor U14005 (N_14005,N_13467,N_13234);
xnor U14006 (N_14006,N_13617,N_13597);
nand U14007 (N_14007,N_13551,N_13696);
nor U14008 (N_14008,N_13264,N_13282);
or U14009 (N_14009,N_13516,N_13453);
xor U14010 (N_14010,N_13253,N_13263);
and U14011 (N_14011,N_13305,N_13294);
or U14012 (N_14012,N_13425,N_13213);
nand U14013 (N_14013,N_13490,N_13647);
nand U14014 (N_14014,N_13537,N_13714);
nor U14015 (N_14015,N_13512,N_13346);
xor U14016 (N_14016,N_13557,N_13254);
nand U14017 (N_14017,N_13212,N_13369);
xnor U14018 (N_14018,N_13211,N_13443);
xor U14019 (N_14019,N_13507,N_13690);
and U14020 (N_14020,N_13792,N_13432);
and U14021 (N_14021,N_13364,N_13748);
nor U14022 (N_14022,N_13485,N_13233);
and U14023 (N_14023,N_13370,N_13349);
and U14024 (N_14024,N_13628,N_13498);
or U14025 (N_14025,N_13268,N_13675);
or U14026 (N_14026,N_13737,N_13593);
or U14027 (N_14027,N_13239,N_13625);
nor U14028 (N_14028,N_13665,N_13619);
nor U14029 (N_14029,N_13431,N_13529);
or U14030 (N_14030,N_13604,N_13576);
and U14031 (N_14031,N_13510,N_13745);
and U14032 (N_14032,N_13589,N_13640);
nor U14033 (N_14033,N_13514,N_13559);
nor U14034 (N_14034,N_13314,N_13389);
nand U14035 (N_14035,N_13357,N_13407);
nand U14036 (N_14036,N_13680,N_13600);
nor U14037 (N_14037,N_13533,N_13727);
and U14038 (N_14038,N_13286,N_13378);
nand U14039 (N_14039,N_13361,N_13729);
nor U14040 (N_14040,N_13703,N_13229);
nand U14041 (N_14041,N_13402,N_13381);
xor U14042 (N_14042,N_13444,N_13598);
nor U14043 (N_14043,N_13513,N_13630);
and U14044 (N_14044,N_13701,N_13341);
nand U14045 (N_14045,N_13410,N_13742);
xor U14046 (N_14046,N_13764,N_13461);
xnor U14047 (N_14047,N_13222,N_13656);
xnor U14048 (N_14048,N_13790,N_13423);
xor U14049 (N_14049,N_13676,N_13319);
xor U14050 (N_14050,N_13674,N_13783);
and U14051 (N_14051,N_13599,N_13789);
nor U14052 (N_14052,N_13350,N_13591);
nand U14053 (N_14053,N_13544,N_13371);
xnor U14054 (N_14054,N_13455,N_13429);
or U14055 (N_14055,N_13398,N_13382);
nand U14056 (N_14056,N_13725,N_13390);
nand U14057 (N_14057,N_13313,N_13782);
nand U14058 (N_14058,N_13439,N_13592);
nand U14059 (N_14059,N_13502,N_13749);
nor U14060 (N_14060,N_13257,N_13506);
or U14061 (N_14061,N_13720,N_13700);
nor U14062 (N_14062,N_13635,N_13678);
nand U14063 (N_14063,N_13481,N_13223);
or U14064 (N_14064,N_13659,N_13755);
nand U14065 (N_14065,N_13491,N_13612);
nor U14066 (N_14066,N_13694,N_13552);
nand U14067 (N_14067,N_13772,N_13422);
or U14068 (N_14068,N_13570,N_13759);
and U14069 (N_14069,N_13441,N_13373);
and U14070 (N_14070,N_13785,N_13652);
xor U14071 (N_14071,N_13743,N_13209);
nand U14072 (N_14072,N_13679,N_13347);
xor U14073 (N_14073,N_13522,N_13596);
xor U14074 (N_14074,N_13583,N_13704);
or U14075 (N_14075,N_13793,N_13650);
and U14076 (N_14076,N_13758,N_13767);
and U14077 (N_14077,N_13578,N_13494);
nand U14078 (N_14078,N_13588,N_13621);
and U14079 (N_14079,N_13471,N_13666);
nand U14080 (N_14080,N_13293,N_13310);
xor U14081 (N_14081,N_13448,N_13728);
nand U14082 (N_14082,N_13766,N_13484);
and U14083 (N_14083,N_13476,N_13734);
or U14084 (N_14084,N_13606,N_13555);
nand U14085 (N_14085,N_13278,N_13673);
xnor U14086 (N_14086,N_13324,N_13798);
and U14087 (N_14087,N_13501,N_13427);
nand U14088 (N_14088,N_13733,N_13752);
nand U14089 (N_14089,N_13480,N_13419);
xnor U14090 (N_14090,N_13562,N_13681);
nor U14091 (N_14091,N_13287,N_13299);
nand U14092 (N_14092,N_13575,N_13605);
nand U14093 (N_14093,N_13285,N_13221);
xnor U14094 (N_14094,N_13384,N_13760);
or U14095 (N_14095,N_13272,N_13392);
and U14096 (N_14096,N_13623,N_13408);
nand U14097 (N_14097,N_13682,N_13243);
nor U14098 (N_14098,N_13648,N_13735);
xnor U14099 (N_14099,N_13545,N_13637);
nand U14100 (N_14100,N_13654,N_13425);
xnor U14101 (N_14101,N_13630,N_13473);
nor U14102 (N_14102,N_13666,N_13654);
or U14103 (N_14103,N_13469,N_13457);
xnor U14104 (N_14104,N_13285,N_13683);
or U14105 (N_14105,N_13258,N_13645);
xor U14106 (N_14106,N_13426,N_13699);
and U14107 (N_14107,N_13798,N_13533);
and U14108 (N_14108,N_13436,N_13321);
xnor U14109 (N_14109,N_13559,N_13284);
and U14110 (N_14110,N_13653,N_13265);
nand U14111 (N_14111,N_13450,N_13214);
and U14112 (N_14112,N_13466,N_13688);
nor U14113 (N_14113,N_13651,N_13492);
nor U14114 (N_14114,N_13650,N_13284);
or U14115 (N_14115,N_13679,N_13668);
nand U14116 (N_14116,N_13478,N_13270);
nor U14117 (N_14117,N_13679,N_13426);
nor U14118 (N_14118,N_13498,N_13418);
nand U14119 (N_14119,N_13281,N_13298);
nand U14120 (N_14120,N_13741,N_13523);
nor U14121 (N_14121,N_13775,N_13241);
or U14122 (N_14122,N_13617,N_13560);
and U14123 (N_14123,N_13674,N_13639);
and U14124 (N_14124,N_13554,N_13687);
and U14125 (N_14125,N_13344,N_13467);
or U14126 (N_14126,N_13715,N_13568);
nand U14127 (N_14127,N_13243,N_13770);
nor U14128 (N_14128,N_13766,N_13660);
nand U14129 (N_14129,N_13200,N_13632);
and U14130 (N_14130,N_13768,N_13361);
xnor U14131 (N_14131,N_13574,N_13380);
xor U14132 (N_14132,N_13450,N_13218);
nand U14133 (N_14133,N_13735,N_13333);
or U14134 (N_14134,N_13294,N_13763);
nor U14135 (N_14135,N_13644,N_13353);
nor U14136 (N_14136,N_13671,N_13332);
or U14137 (N_14137,N_13498,N_13340);
nor U14138 (N_14138,N_13606,N_13684);
nand U14139 (N_14139,N_13357,N_13216);
nor U14140 (N_14140,N_13732,N_13320);
or U14141 (N_14141,N_13632,N_13784);
nor U14142 (N_14142,N_13439,N_13696);
or U14143 (N_14143,N_13231,N_13420);
or U14144 (N_14144,N_13474,N_13326);
xor U14145 (N_14145,N_13231,N_13421);
or U14146 (N_14146,N_13409,N_13512);
nand U14147 (N_14147,N_13524,N_13269);
nand U14148 (N_14148,N_13726,N_13529);
and U14149 (N_14149,N_13235,N_13567);
and U14150 (N_14150,N_13594,N_13307);
and U14151 (N_14151,N_13520,N_13441);
xnor U14152 (N_14152,N_13280,N_13383);
nand U14153 (N_14153,N_13729,N_13373);
nor U14154 (N_14154,N_13692,N_13572);
or U14155 (N_14155,N_13784,N_13316);
nand U14156 (N_14156,N_13519,N_13293);
and U14157 (N_14157,N_13205,N_13676);
nand U14158 (N_14158,N_13498,N_13274);
or U14159 (N_14159,N_13274,N_13390);
nand U14160 (N_14160,N_13765,N_13251);
nor U14161 (N_14161,N_13416,N_13548);
and U14162 (N_14162,N_13572,N_13710);
or U14163 (N_14163,N_13706,N_13304);
nand U14164 (N_14164,N_13489,N_13764);
nand U14165 (N_14165,N_13459,N_13461);
xnor U14166 (N_14166,N_13723,N_13799);
and U14167 (N_14167,N_13517,N_13732);
or U14168 (N_14168,N_13456,N_13444);
or U14169 (N_14169,N_13475,N_13638);
or U14170 (N_14170,N_13649,N_13659);
xnor U14171 (N_14171,N_13308,N_13513);
and U14172 (N_14172,N_13759,N_13519);
nand U14173 (N_14173,N_13271,N_13233);
and U14174 (N_14174,N_13623,N_13274);
xor U14175 (N_14175,N_13276,N_13501);
xnor U14176 (N_14176,N_13269,N_13503);
or U14177 (N_14177,N_13352,N_13398);
or U14178 (N_14178,N_13785,N_13513);
and U14179 (N_14179,N_13321,N_13294);
and U14180 (N_14180,N_13380,N_13253);
nor U14181 (N_14181,N_13426,N_13763);
and U14182 (N_14182,N_13420,N_13338);
or U14183 (N_14183,N_13392,N_13778);
or U14184 (N_14184,N_13223,N_13710);
nor U14185 (N_14185,N_13392,N_13234);
or U14186 (N_14186,N_13535,N_13366);
xor U14187 (N_14187,N_13449,N_13474);
or U14188 (N_14188,N_13797,N_13574);
xnor U14189 (N_14189,N_13347,N_13589);
or U14190 (N_14190,N_13546,N_13305);
xor U14191 (N_14191,N_13688,N_13308);
and U14192 (N_14192,N_13573,N_13734);
nand U14193 (N_14193,N_13604,N_13209);
nor U14194 (N_14194,N_13526,N_13335);
xor U14195 (N_14195,N_13688,N_13787);
xor U14196 (N_14196,N_13718,N_13436);
nor U14197 (N_14197,N_13344,N_13715);
and U14198 (N_14198,N_13696,N_13781);
nor U14199 (N_14199,N_13445,N_13212);
nand U14200 (N_14200,N_13782,N_13607);
or U14201 (N_14201,N_13503,N_13532);
or U14202 (N_14202,N_13588,N_13494);
xor U14203 (N_14203,N_13739,N_13480);
nand U14204 (N_14204,N_13266,N_13344);
nand U14205 (N_14205,N_13541,N_13792);
nand U14206 (N_14206,N_13535,N_13753);
xor U14207 (N_14207,N_13688,N_13653);
or U14208 (N_14208,N_13680,N_13339);
nor U14209 (N_14209,N_13331,N_13211);
xnor U14210 (N_14210,N_13738,N_13210);
or U14211 (N_14211,N_13580,N_13599);
and U14212 (N_14212,N_13690,N_13365);
nor U14213 (N_14213,N_13684,N_13753);
nor U14214 (N_14214,N_13436,N_13598);
nor U14215 (N_14215,N_13591,N_13631);
and U14216 (N_14216,N_13548,N_13472);
nand U14217 (N_14217,N_13566,N_13445);
nand U14218 (N_14218,N_13519,N_13522);
and U14219 (N_14219,N_13399,N_13492);
xnor U14220 (N_14220,N_13558,N_13790);
nor U14221 (N_14221,N_13594,N_13500);
and U14222 (N_14222,N_13530,N_13483);
xnor U14223 (N_14223,N_13796,N_13264);
xnor U14224 (N_14224,N_13588,N_13204);
and U14225 (N_14225,N_13792,N_13276);
and U14226 (N_14226,N_13710,N_13743);
and U14227 (N_14227,N_13367,N_13273);
and U14228 (N_14228,N_13706,N_13779);
nor U14229 (N_14229,N_13599,N_13654);
nor U14230 (N_14230,N_13665,N_13264);
xor U14231 (N_14231,N_13681,N_13658);
and U14232 (N_14232,N_13266,N_13667);
or U14233 (N_14233,N_13266,N_13545);
or U14234 (N_14234,N_13337,N_13673);
and U14235 (N_14235,N_13565,N_13654);
and U14236 (N_14236,N_13737,N_13284);
xor U14237 (N_14237,N_13394,N_13307);
nand U14238 (N_14238,N_13584,N_13254);
nor U14239 (N_14239,N_13661,N_13628);
or U14240 (N_14240,N_13574,N_13581);
nor U14241 (N_14241,N_13415,N_13583);
and U14242 (N_14242,N_13407,N_13527);
nor U14243 (N_14243,N_13234,N_13351);
xor U14244 (N_14244,N_13606,N_13599);
or U14245 (N_14245,N_13632,N_13564);
nor U14246 (N_14246,N_13364,N_13660);
nor U14247 (N_14247,N_13394,N_13516);
xor U14248 (N_14248,N_13674,N_13325);
xor U14249 (N_14249,N_13605,N_13676);
or U14250 (N_14250,N_13611,N_13441);
nand U14251 (N_14251,N_13342,N_13694);
nand U14252 (N_14252,N_13383,N_13585);
nand U14253 (N_14253,N_13534,N_13789);
nand U14254 (N_14254,N_13650,N_13436);
nand U14255 (N_14255,N_13361,N_13451);
xnor U14256 (N_14256,N_13312,N_13423);
or U14257 (N_14257,N_13771,N_13633);
nor U14258 (N_14258,N_13457,N_13353);
nor U14259 (N_14259,N_13689,N_13649);
xnor U14260 (N_14260,N_13342,N_13532);
nand U14261 (N_14261,N_13309,N_13431);
and U14262 (N_14262,N_13652,N_13778);
or U14263 (N_14263,N_13272,N_13660);
nor U14264 (N_14264,N_13549,N_13472);
and U14265 (N_14265,N_13770,N_13793);
xnor U14266 (N_14266,N_13566,N_13424);
or U14267 (N_14267,N_13369,N_13375);
xnor U14268 (N_14268,N_13632,N_13390);
or U14269 (N_14269,N_13519,N_13643);
and U14270 (N_14270,N_13430,N_13333);
and U14271 (N_14271,N_13398,N_13775);
xor U14272 (N_14272,N_13481,N_13391);
xor U14273 (N_14273,N_13646,N_13597);
and U14274 (N_14274,N_13548,N_13454);
nor U14275 (N_14275,N_13719,N_13216);
nand U14276 (N_14276,N_13335,N_13307);
xor U14277 (N_14277,N_13288,N_13239);
nor U14278 (N_14278,N_13311,N_13591);
xnor U14279 (N_14279,N_13264,N_13767);
and U14280 (N_14280,N_13419,N_13637);
and U14281 (N_14281,N_13258,N_13281);
and U14282 (N_14282,N_13316,N_13619);
and U14283 (N_14283,N_13307,N_13265);
nand U14284 (N_14284,N_13324,N_13265);
nor U14285 (N_14285,N_13740,N_13358);
and U14286 (N_14286,N_13620,N_13610);
and U14287 (N_14287,N_13768,N_13628);
and U14288 (N_14288,N_13463,N_13317);
or U14289 (N_14289,N_13686,N_13732);
nand U14290 (N_14290,N_13364,N_13245);
or U14291 (N_14291,N_13437,N_13608);
nand U14292 (N_14292,N_13382,N_13574);
nand U14293 (N_14293,N_13348,N_13770);
or U14294 (N_14294,N_13725,N_13735);
nor U14295 (N_14295,N_13367,N_13316);
nor U14296 (N_14296,N_13311,N_13671);
nand U14297 (N_14297,N_13552,N_13233);
nand U14298 (N_14298,N_13283,N_13426);
or U14299 (N_14299,N_13495,N_13561);
xor U14300 (N_14300,N_13682,N_13358);
or U14301 (N_14301,N_13773,N_13787);
nor U14302 (N_14302,N_13581,N_13713);
or U14303 (N_14303,N_13423,N_13484);
nand U14304 (N_14304,N_13696,N_13518);
and U14305 (N_14305,N_13249,N_13342);
xnor U14306 (N_14306,N_13376,N_13395);
or U14307 (N_14307,N_13619,N_13627);
nand U14308 (N_14308,N_13343,N_13281);
nor U14309 (N_14309,N_13525,N_13322);
nor U14310 (N_14310,N_13260,N_13514);
nand U14311 (N_14311,N_13333,N_13297);
xnor U14312 (N_14312,N_13202,N_13729);
and U14313 (N_14313,N_13242,N_13221);
xnor U14314 (N_14314,N_13697,N_13427);
nor U14315 (N_14315,N_13733,N_13692);
nor U14316 (N_14316,N_13729,N_13431);
and U14317 (N_14317,N_13727,N_13415);
xor U14318 (N_14318,N_13295,N_13471);
and U14319 (N_14319,N_13726,N_13703);
and U14320 (N_14320,N_13373,N_13390);
nor U14321 (N_14321,N_13461,N_13455);
or U14322 (N_14322,N_13625,N_13271);
or U14323 (N_14323,N_13453,N_13243);
xor U14324 (N_14324,N_13636,N_13610);
or U14325 (N_14325,N_13757,N_13471);
xnor U14326 (N_14326,N_13547,N_13799);
and U14327 (N_14327,N_13799,N_13618);
nand U14328 (N_14328,N_13720,N_13224);
or U14329 (N_14329,N_13465,N_13567);
xnor U14330 (N_14330,N_13448,N_13472);
and U14331 (N_14331,N_13698,N_13354);
xor U14332 (N_14332,N_13509,N_13685);
nand U14333 (N_14333,N_13519,N_13612);
nand U14334 (N_14334,N_13463,N_13758);
or U14335 (N_14335,N_13630,N_13452);
nand U14336 (N_14336,N_13688,N_13712);
and U14337 (N_14337,N_13753,N_13776);
nor U14338 (N_14338,N_13407,N_13247);
or U14339 (N_14339,N_13794,N_13428);
nor U14340 (N_14340,N_13458,N_13450);
or U14341 (N_14341,N_13500,N_13235);
nor U14342 (N_14342,N_13523,N_13266);
xnor U14343 (N_14343,N_13283,N_13754);
xor U14344 (N_14344,N_13617,N_13653);
nor U14345 (N_14345,N_13772,N_13673);
nor U14346 (N_14346,N_13408,N_13378);
nor U14347 (N_14347,N_13621,N_13228);
xnor U14348 (N_14348,N_13662,N_13719);
xnor U14349 (N_14349,N_13549,N_13577);
nand U14350 (N_14350,N_13289,N_13673);
and U14351 (N_14351,N_13539,N_13630);
nor U14352 (N_14352,N_13446,N_13766);
and U14353 (N_14353,N_13518,N_13391);
xor U14354 (N_14354,N_13283,N_13556);
or U14355 (N_14355,N_13702,N_13648);
and U14356 (N_14356,N_13456,N_13794);
xnor U14357 (N_14357,N_13239,N_13356);
xor U14358 (N_14358,N_13275,N_13578);
nor U14359 (N_14359,N_13684,N_13499);
xor U14360 (N_14360,N_13488,N_13638);
nor U14361 (N_14361,N_13554,N_13470);
or U14362 (N_14362,N_13341,N_13475);
nor U14363 (N_14363,N_13417,N_13522);
nor U14364 (N_14364,N_13380,N_13349);
xnor U14365 (N_14365,N_13260,N_13472);
and U14366 (N_14366,N_13738,N_13569);
xnor U14367 (N_14367,N_13289,N_13371);
nand U14368 (N_14368,N_13319,N_13430);
nor U14369 (N_14369,N_13329,N_13712);
or U14370 (N_14370,N_13737,N_13312);
and U14371 (N_14371,N_13485,N_13559);
and U14372 (N_14372,N_13503,N_13595);
and U14373 (N_14373,N_13532,N_13370);
nand U14374 (N_14374,N_13400,N_13726);
and U14375 (N_14375,N_13447,N_13608);
nand U14376 (N_14376,N_13627,N_13456);
and U14377 (N_14377,N_13438,N_13511);
nor U14378 (N_14378,N_13722,N_13421);
and U14379 (N_14379,N_13685,N_13511);
xor U14380 (N_14380,N_13638,N_13771);
or U14381 (N_14381,N_13364,N_13445);
nand U14382 (N_14382,N_13439,N_13341);
nor U14383 (N_14383,N_13722,N_13523);
nor U14384 (N_14384,N_13396,N_13355);
or U14385 (N_14385,N_13362,N_13733);
nor U14386 (N_14386,N_13319,N_13236);
or U14387 (N_14387,N_13694,N_13630);
nor U14388 (N_14388,N_13624,N_13217);
nand U14389 (N_14389,N_13717,N_13356);
nand U14390 (N_14390,N_13259,N_13749);
or U14391 (N_14391,N_13456,N_13475);
nand U14392 (N_14392,N_13629,N_13699);
and U14393 (N_14393,N_13421,N_13716);
xor U14394 (N_14394,N_13562,N_13447);
nand U14395 (N_14395,N_13588,N_13275);
nor U14396 (N_14396,N_13641,N_13459);
or U14397 (N_14397,N_13227,N_13419);
and U14398 (N_14398,N_13220,N_13323);
xor U14399 (N_14399,N_13231,N_13485);
or U14400 (N_14400,N_14283,N_13984);
nor U14401 (N_14401,N_14331,N_14355);
and U14402 (N_14402,N_13973,N_14307);
or U14403 (N_14403,N_13906,N_13961);
and U14404 (N_14404,N_14090,N_14238);
nand U14405 (N_14405,N_14374,N_13941);
or U14406 (N_14406,N_13917,N_14073);
or U14407 (N_14407,N_14266,N_13985);
nor U14408 (N_14408,N_14182,N_14080);
xor U14409 (N_14409,N_14148,N_14013);
nor U14410 (N_14410,N_14152,N_14246);
nor U14411 (N_14411,N_14033,N_14378);
xor U14412 (N_14412,N_13820,N_14149);
xor U14413 (N_14413,N_13910,N_14397);
xnor U14414 (N_14414,N_14293,N_14213);
and U14415 (N_14415,N_13949,N_14169);
nand U14416 (N_14416,N_13840,N_13905);
xnor U14417 (N_14417,N_14196,N_13998);
and U14418 (N_14418,N_14019,N_14278);
nor U14419 (N_14419,N_14223,N_14018);
nor U14420 (N_14420,N_13940,N_14275);
xor U14421 (N_14421,N_14204,N_13821);
or U14422 (N_14422,N_13945,N_13921);
nor U14423 (N_14423,N_14039,N_14093);
xnor U14424 (N_14424,N_13895,N_14072);
xnor U14425 (N_14425,N_14021,N_14024);
nor U14426 (N_14426,N_13926,N_14311);
nand U14427 (N_14427,N_14134,N_14390);
nand U14428 (N_14428,N_14023,N_13878);
or U14429 (N_14429,N_14343,N_13986);
or U14430 (N_14430,N_14012,N_14339);
xnor U14431 (N_14431,N_14187,N_13849);
and U14432 (N_14432,N_14146,N_13946);
and U14433 (N_14433,N_14245,N_14167);
nand U14434 (N_14434,N_14208,N_14360);
xor U14435 (N_14435,N_13831,N_14124);
nor U14436 (N_14436,N_14011,N_13979);
or U14437 (N_14437,N_13992,N_14352);
xor U14438 (N_14438,N_14359,N_13935);
nor U14439 (N_14439,N_13835,N_14086);
nor U14440 (N_14440,N_14338,N_14209);
nand U14441 (N_14441,N_14108,N_13823);
or U14442 (N_14442,N_14285,N_14040);
or U14443 (N_14443,N_13809,N_14372);
nor U14444 (N_14444,N_14261,N_14370);
nor U14445 (N_14445,N_14294,N_14098);
xor U14446 (N_14446,N_14003,N_13960);
nand U14447 (N_14447,N_13892,N_14353);
nor U14448 (N_14448,N_14198,N_13863);
xnor U14449 (N_14449,N_14303,N_13942);
nand U14450 (N_14450,N_14308,N_13964);
nand U14451 (N_14451,N_14221,N_13890);
or U14452 (N_14452,N_14186,N_14113);
nand U14453 (N_14453,N_14335,N_14350);
nor U14454 (N_14454,N_14361,N_14314);
xor U14455 (N_14455,N_13933,N_14006);
and U14456 (N_14456,N_13885,N_13834);
or U14457 (N_14457,N_14328,N_13853);
xnor U14458 (N_14458,N_14380,N_14357);
nor U14459 (N_14459,N_14399,N_13841);
or U14460 (N_14460,N_14009,N_13873);
xor U14461 (N_14461,N_13925,N_14016);
nor U14462 (N_14462,N_14337,N_14202);
and U14463 (N_14463,N_13909,N_13970);
nor U14464 (N_14464,N_14005,N_13819);
or U14465 (N_14465,N_14385,N_13958);
nor U14466 (N_14466,N_14274,N_14387);
or U14467 (N_14467,N_14068,N_14162);
and U14468 (N_14468,N_14103,N_13860);
xnor U14469 (N_14469,N_14161,N_14048);
nand U14470 (N_14470,N_14156,N_13988);
or U14471 (N_14471,N_13957,N_14346);
nand U14472 (N_14472,N_14194,N_14078);
nand U14473 (N_14473,N_14295,N_13865);
xor U14474 (N_14474,N_14392,N_13805);
and U14475 (N_14475,N_14030,N_14114);
xor U14476 (N_14476,N_14118,N_14287);
and U14477 (N_14477,N_14371,N_13887);
nand U14478 (N_14478,N_14061,N_14244);
and U14479 (N_14479,N_13978,N_14174);
xnor U14480 (N_14480,N_14166,N_14193);
and U14481 (N_14481,N_14304,N_14233);
xnor U14482 (N_14482,N_14249,N_14368);
nand U14483 (N_14483,N_13822,N_14047);
nand U14484 (N_14484,N_14289,N_14083);
or U14485 (N_14485,N_14165,N_14127);
nor U14486 (N_14486,N_14321,N_13882);
or U14487 (N_14487,N_14237,N_14260);
nor U14488 (N_14488,N_14345,N_14111);
nor U14489 (N_14489,N_14248,N_14173);
and U14490 (N_14490,N_14032,N_14170);
and U14491 (N_14491,N_14325,N_14354);
and U14492 (N_14492,N_14376,N_14130);
nor U14493 (N_14493,N_14207,N_13826);
xor U14494 (N_14494,N_14183,N_14117);
xnor U14495 (N_14495,N_13918,N_13971);
xnor U14496 (N_14496,N_14153,N_13923);
and U14497 (N_14497,N_13824,N_14126);
xor U14498 (N_14498,N_14190,N_14042);
and U14499 (N_14499,N_13886,N_14200);
xnor U14500 (N_14500,N_14389,N_14089);
nor U14501 (N_14501,N_14097,N_14375);
or U14502 (N_14502,N_13943,N_14273);
and U14503 (N_14503,N_14116,N_13884);
and U14504 (N_14504,N_14020,N_14091);
or U14505 (N_14505,N_13838,N_14230);
nand U14506 (N_14506,N_13876,N_14188);
or U14507 (N_14507,N_14057,N_14300);
or U14508 (N_14508,N_13847,N_13851);
and U14509 (N_14509,N_14277,N_14034);
xor U14510 (N_14510,N_14205,N_13829);
nand U14511 (N_14511,N_13915,N_14365);
nor U14512 (N_14512,N_13830,N_14071);
xor U14513 (N_14513,N_14171,N_14324);
xor U14514 (N_14514,N_14143,N_13811);
and U14515 (N_14515,N_14065,N_13939);
xnor U14516 (N_14516,N_14029,N_14004);
nor U14517 (N_14517,N_14235,N_13994);
nand U14518 (N_14518,N_13952,N_13974);
and U14519 (N_14519,N_14382,N_13810);
or U14520 (N_14520,N_14059,N_13833);
or U14521 (N_14521,N_13968,N_14128);
nor U14522 (N_14522,N_14053,N_13862);
nand U14523 (N_14523,N_14122,N_14251);
nand U14524 (N_14524,N_14177,N_14210);
xor U14525 (N_14525,N_14102,N_14329);
xnor U14526 (N_14526,N_14082,N_14270);
nor U14527 (N_14527,N_14322,N_14120);
nor U14528 (N_14528,N_14280,N_13959);
xor U14529 (N_14529,N_14369,N_14227);
nor U14530 (N_14530,N_14229,N_14211);
xnor U14531 (N_14531,N_14381,N_13813);
nor U14532 (N_14532,N_14250,N_14144);
nand U14533 (N_14533,N_14074,N_14041);
or U14534 (N_14534,N_13936,N_13894);
xnor U14535 (N_14535,N_14301,N_14298);
nand U14536 (N_14536,N_13897,N_14031);
nor U14537 (N_14537,N_14388,N_14394);
nand U14538 (N_14538,N_14069,N_13857);
nor U14539 (N_14539,N_14362,N_14231);
nand U14540 (N_14540,N_13907,N_14131);
nand U14541 (N_14541,N_14062,N_14077);
or U14542 (N_14542,N_14168,N_14136);
and U14543 (N_14543,N_14038,N_14263);
nand U14544 (N_14544,N_14348,N_14220);
or U14545 (N_14545,N_14297,N_14133);
nor U14546 (N_14546,N_13877,N_13914);
nor U14547 (N_14547,N_13870,N_13983);
nand U14548 (N_14548,N_14054,N_13956);
or U14549 (N_14549,N_13927,N_13814);
nor U14550 (N_14550,N_14225,N_14035);
nand U14551 (N_14551,N_14036,N_14224);
nor U14552 (N_14552,N_14290,N_13919);
or U14553 (N_14553,N_14119,N_13975);
or U14554 (N_14554,N_14101,N_14259);
or U14555 (N_14555,N_13896,N_14257);
xnor U14556 (N_14556,N_14140,N_13997);
or U14557 (N_14557,N_14109,N_14395);
and U14558 (N_14558,N_13911,N_14219);
or U14559 (N_14559,N_14125,N_14215);
and U14560 (N_14560,N_14367,N_13981);
nand U14561 (N_14561,N_14067,N_14253);
nand U14562 (N_14562,N_13867,N_14323);
xnor U14563 (N_14563,N_14234,N_14104);
nand U14564 (N_14564,N_13804,N_14037);
xor U14565 (N_14565,N_13965,N_14342);
nor U14566 (N_14566,N_13976,N_13871);
xor U14567 (N_14567,N_13891,N_14272);
and U14568 (N_14568,N_14007,N_14028);
nor U14569 (N_14569,N_14100,N_14099);
nor U14570 (N_14570,N_14154,N_13812);
or U14571 (N_14571,N_14305,N_14141);
nand U14572 (N_14572,N_14159,N_13928);
nand U14573 (N_14573,N_14351,N_14180);
or U14574 (N_14574,N_13913,N_13880);
nand U14575 (N_14575,N_13991,N_13903);
nand U14576 (N_14576,N_13962,N_13980);
nor U14577 (N_14577,N_14066,N_13931);
or U14578 (N_14578,N_14269,N_14265);
nand U14579 (N_14579,N_13845,N_13825);
and U14580 (N_14580,N_13855,N_14236);
or U14581 (N_14581,N_14192,N_14115);
and U14582 (N_14582,N_14060,N_14317);
and U14583 (N_14583,N_14226,N_13874);
and U14584 (N_14584,N_14185,N_13869);
xor U14585 (N_14585,N_14214,N_14002);
xnor U14586 (N_14586,N_13990,N_14129);
and U14587 (N_14587,N_13837,N_14212);
or U14588 (N_14588,N_14046,N_14216);
nand U14589 (N_14589,N_14123,N_14106);
nor U14590 (N_14590,N_13881,N_14096);
xnor U14591 (N_14591,N_14306,N_13859);
xnor U14592 (N_14592,N_13938,N_14377);
nor U14593 (N_14593,N_14001,N_14296);
nor U14594 (N_14594,N_13844,N_14094);
and U14595 (N_14595,N_14396,N_14292);
and U14596 (N_14596,N_14332,N_13889);
nand U14597 (N_14597,N_13948,N_14151);
or U14598 (N_14598,N_14199,N_14302);
and U14599 (N_14599,N_14058,N_14085);
and U14600 (N_14600,N_14049,N_14195);
nand U14601 (N_14601,N_13888,N_14175);
nand U14602 (N_14602,N_13852,N_14178);
or U14603 (N_14603,N_13828,N_13932);
nor U14604 (N_14604,N_14391,N_13817);
and U14605 (N_14605,N_13879,N_14142);
nand U14606 (N_14606,N_14256,N_14055);
nor U14607 (N_14607,N_13920,N_14064);
nand U14608 (N_14608,N_14241,N_13944);
nor U14609 (N_14609,N_13987,N_14027);
and U14610 (N_14610,N_14240,N_14158);
or U14611 (N_14611,N_14313,N_13807);
nand U14612 (N_14612,N_14336,N_14373);
or U14613 (N_14613,N_14135,N_13953);
xnor U14614 (N_14614,N_13848,N_14150);
and U14615 (N_14615,N_14110,N_14184);
nand U14616 (N_14616,N_14267,N_14384);
nand U14617 (N_14617,N_14326,N_13864);
nor U14618 (N_14618,N_14056,N_14330);
and U14619 (N_14619,N_14268,N_13861);
nand U14620 (N_14620,N_14309,N_14201);
nand U14621 (N_14621,N_14264,N_14383);
nand U14622 (N_14622,N_14315,N_13854);
and U14623 (N_14623,N_14333,N_13832);
xnor U14624 (N_14624,N_14087,N_14203);
xnor U14625 (N_14625,N_13868,N_13916);
nor U14626 (N_14626,N_13856,N_13898);
nand U14627 (N_14627,N_14138,N_14132);
or U14628 (N_14628,N_13977,N_13929);
nor U14629 (N_14629,N_14107,N_13866);
nor U14630 (N_14630,N_14393,N_13954);
or U14631 (N_14631,N_14105,N_14147);
and U14632 (N_14632,N_14121,N_14242);
xor U14633 (N_14633,N_14088,N_14398);
or U14634 (N_14634,N_14197,N_14095);
nand U14635 (N_14635,N_14081,N_14164);
xor U14636 (N_14636,N_14084,N_14320);
nor U14637 (N_14637,N_14022,N_14026);
xnor U14638 (N_14638,N_14222,N_13995);
xnor U14639 (N_14639,N_13808,N_13815);
nand U14640 (N_14640,N_14218,N_14243);
nand U14641 (N_14641,N_13904,N_14079);
and U14642 (N_14642,N_14327,N_14163);
nand U14643 (N_14643,N_14176,N_14043);
or U14644 (N_14644,N_13872,N_14310);
and U14645 (N_14645,N_14366,N_14172);
nor U14646 (N_14646,N_13924,N_13893);
and U14647 (N_14647,N_13934,N_14316);
or U14648 (N_14648,N_13963,N_13858);
xnor U14649 (N_14649,N_13803,N_13800);
xor U14650 (N_14650,N_14157,N_14255);
xor U14651 (N_14651,N_14000,N_14341);
and U14652 (N_14652,N_14044,N_13950);
and U14653 (N_14653,N_13818,N_14386);
nand U14654 (N_14654,N_14239,N_14191);
or U14655 (N_14655,N_14045,N_14364);
xnor U14656 (N_14656,N_14189,N_14145);
or U14657 (N_14657,N_14008,N_14075);
nor U14658 (N_14658,N_13883,N_14281);
xnor U14659 (N_14659,N_14291,N_14358);
nand U14660 (N_14660,N_14356,N_13843);
and U14661 (N_14661,N_13827,N_14279);
nor U14662 (N_14662,N_14160,N_13842);
or U14663 (N_14663,N_13955,N_13972);
nand U14664 (N_14664,N_14262,N_14347);
or U14665 (N_14665,N_13969,N_13912);
nand U14666 (N_14666,N_14010,N_14340);
nand U14667 (N_14667,N_13908,N_13839);
or U14668 (N_14668,N_14282,N_14284);
and U14669 (N_14669,N_14252,N_14217);
or U14670 (N_14670,N_14247,N_13937);
nor U14671 (N_14671,N_14139,N_13899);
xor U14672 (N_14672,N_13802,N_13902);
or U14673 (N_14673,N_13966,N_13982);
xnor U14674 (N_14674,N_14112,N_14228);
xor U14675 (N_14675,N_14137,N_14076);
nor U14676 (N_14676,N_14276,N_14232);
nor U14677 (N_14677,N_14179,N_13801);
xor U14678 (N_14678,N_13846,N_14334);
or U14679 (N_14679,N_14318,N_14017);
nand U14680 (N_14680,N_13816,N_14288);
and U14681 (N_14681,N_13806,N_14271);
or U14682 (N_14682,N_14181,N_14051);
nand U14683 (N_14683,N_14258,N_13850);
nand U14684 (N_14684,N_13967,N_13836);
nor U14685 (N_14685,N_13989,N_14092);
or U14686 (N_14686,N_14050,N_14014);
and U14687 (N_14687,N_14025,N_14299);
xor U14688 (N_14688,N_13875,N_13930);
nor U14689 (N_14689,N_14155,N_14286);
and U14690 (N_14690,N_14070,N_13900);
nand U14691 (N_14691,N_13999,N_14344);
xor U14692 (N_14692,N_14379,N_14254);
nor U14693 (N_14693,N_14052,N_13951);
or U14694 (N_14694,N_13922,N_14312);
nand U14695 (N_14695,N_14363,N_14206);
nand U14696 (N_14696,N_13947,N_13901);
or U14697 (N_14697,N_14063,N_14349);
or U14698 (N_14698,N_13993,N_14319);
nand U14699 (N_14699,N_13996,N_14015);
and U14700 (N_14700,N_14197,N_14211);
or U14701 (N_14701,N_14356,N_14362);
or U14702 (N_14702,N_14325,N_14315);
and U14703 (N_14703,N_13985,N_13914);
or U14704 (N_14704,N_14119,N_14332);
and U14705 (N_14705,N_14367,N_13807);
nand U14706 (N_14706,N_14099,N_14063);
or U14707 (N_14707,N_13847,N_14098);
xor U14708 (N_14708,N_13836,N_14101);
nand U14709 (N_14709,N_13970,N_14185);
nor U14710 (N_14710,N_14282,N_13935);
xnor U14711 (N_14711,N_14104,N_14067);
nor U14712 (N_14712,N_13859,N_13856);
nand U14713 (N_14713,N_14320,N_14124);
xor U14714 (N_14714,N_13874,N_14073);
nor U14715 (N_14715,N_13900,N_13912);
and U14716 (N_14716,N_13990,N_13874);
xnor U14717 (N_14717,N_14354,N_14087);
nor U14718 (N_14718,N_14034,N_13960);
nor U14719 (N_14719,N_14259,N_13902);
nor U14720 (N_14720,N_14078,N_14140);
nand U14721 (N_14721,N_13942,N_13828);
and U14722 (N_14722,N_14303,N_13880);
or U14723 (N_14723,N_14397,N_14262);
or U14724 (N_14724,N_14285,N_14102);
and U14725 (N_14725,N_13923,N_14338);
and U14726 (N_14726,N_14147,N_14035);
xor U14727 (N_14727,N_13904,N_13946);
nand U14728 (N_14728,N_13866,N_14292);
and U14729 (N_14729,N_14102,N_13841);
and U14730 (N_14730,N_14391,N_14108);
and U14731 (N_14731,N_14116,N_14321);
or U14732 (N_14732,N_13807,N_14031);
and U14733 (N_14733,N_14236,N_13939);
or U14734 (N_14734,N_14260,N_14054);
and U14735 (N_14735,N_14389,N_14295);
or U14736 (N_14736,N_13939,N_13969);
or U14737 (N_14737,N_14180,N_13922);
nor U14738 (N_14738,N_13995,N_14230);
and U14739 (N_14739,N_14354,N_13817);
nor U14740 (N_14740,N_13862,N_13803);
or U14741 (N_14741,N_14378,N_14139);
xnor U14742 (N_14742,N_14139,N_13983);
and U14743 (N_14743,N_14113,N_14065);
or U14744 (N_14744,N_14298,N_14170);
and U14745 (N_14745,N_14399,N_14221);
or U14746 (N_14746,N_14315,N_14259);
nand U14747 (N_14747,N_14130,N_14000);
nor U14748 (N_14748,N_14304,N_14046);
xnor U14749 (N_14749,N_13840,N_13996);
xor U14750 (N_14750,N_13904,N_14213);
and U14751 (N_14751,N_14178,N_14237);
and U14752 (N_14752,N_13812,N_14279);
or U14753 (N_14753,N_14341,N_13914);
or U14754 (N_14754,N_13899,N_14315);
and U14755 (N_14755,N_14161,N_14338);
nor U14756 (N_14756,N_13898,N_14192);
or U14757 (N_14757,N_13958,N_13833);
or U14758 (N_14758,N_14199,N_14059);
nor U14759 (N_14759,N_13889,N_13977);
and U14760 (N_14760,N_14162,N_14381);
and U14761 (N_14761,N_14069,N_13934);
or U14762 (N_14762,N_13854,N_14237);
xnor U14763 (N_14763,N_14120,N_14335);
nor U14764 (N_14764,N_14004,N_13933);
and U14765 (N_14765,N_14184,N_14270);
nor U14766 (N_14766,N_14210,N_14385);
nand U14767 (N_14767,N_14369,N_13834);
xnor U14768 (N_14768,N_13930,N_14343);
or U14769 (N_14769,N_14136,N_13982);
xnor U14770 (N_14770,N_13961,N_14283);
xnor U14771 (N_14771,N_13989,N_14199);
nand U14772 (N_14772,N_14100,N_13856);
nor U14773 (N_14773,N_14224,N_14325);
and U14774 (N_14774,N_14383,N_14251);
or U14775 (N_14775,N_14292,N_13902);
xor U14776 (N_14776,N_14257,N_14016);
or U14777 (N_14777,N_13941,N_13871);
nand U14778 (N_14778,N_14170,N_14355);
nor U14779 (N_14779,N_13824,N_13827);
or U14780 (N_14780,N_14101,N_14150);
nor U14781 (N_14781,N_14197,N_14118);
xnor U14782 (N_14782,N_13802,N_14036);
nor U14783 (N_14783,N_13873,N_13978);
nand U14784 (N_14784,N_14309,N_13807);
xnor U14785 (N_14785,N_14177,N_14024);
or U14786 (N_14786,N_13971,N_14008);
and U14787 (N_14787,N_14038,N_14022);
nand U14788 (N_14788,N_13949,N_13875);
or U14789 (N_14789,N_13831,N_13955);
or U14790 (N_14790,N_13926,N_14321);
nand U14791 (N_14791,N_13847,N_14255);
nor U14792 (N_14792,N_14255,N_14231);
and U14793 (N_14793,N_13950,N_14306);
nand U14794 (N_14794,N_13903,N_14079);
nor U14795 (N_14795,N_13999,N_14112);
nor U14796 (N_14796,N_14078,N_14283);
xor U14797 (N_14797,N_14184,N_14135);
or U14798 (N_14798,N_14096,N_13941);
xor U14799 (N_14799,N_14315,N_13953);
nor U14800 (N_14800,N_14105,N_14169);
nand U14801 (N_14801,N_13940,N_14137);
xor U14802 (N_14802,N_14248,N_14165);
xor U14803 (N_14803,N_13923,N_14142);
nand U14804 (N_14804,N_14222,N_14250);
xor U14805 (N_14805,N_14228,N_13883);
and U14806 (N_14806,N_13835,N_13846);
or U14807 (N_14807,N_13827,N_14287);
and U14808 (N_14808,N_13830,N_14130);
or U14809 (N_14809,N_13982,N_14045);
and U14810 (N_14810,N_14106,N_14243);
nand U14811 (N_14811,N_14346,N_14089);
and U14812 (N_14812,N_13901,N_13978);
nand U14813 (N_14813,N_14259,N_14393);
nor U14814 (N_14814,N_14325,N_14189);
nor U14815 (N_14815,N_14139,N_13830);
xor U14816 (N_14816,N_14041,N_14381);
nor U14817 (N_14817,N_14238,N_14025);
xnor U14818 (N_14818,N_14128,N_13923);
or U14819 (N_14819,N_13992,N_14360);
xor U14820 (N_14820,N_14306,N_13913);
and U14821 (N_14821,N_13895,N_14287);
or U14822 (N_14822,N_14032,N_14110);
nor U14823 (N_14823,N_14358,N_13872);
nor U14824 (N_14824,N_13923,N_13881);
xor U14825 (N_14825,N_13949,N_13982);
nand U14826 (N_14826,N_13818,N_14269);
xnor U14827 (N_14827,N_13919,N_14388);
xor U14828 (N_14828,N_14060,N_13818);
or U14829 (N_14829,N_13967,N_14389);
nand U14830 (N_14830,N_14366,N_14151);
nor U14831 (N_14831,N_14071,N_13822);
or U14832 (N_14832,N_14226,N_13880);
and U14833 (N_14833,N_14187,N_14317);
nand U14834 (N_14834,N_13818,N_14204);
or U14835 (N_14835,N_13991,N_14165);
and U14836 (N_14836,N_14217,N_14096);
nand U14837 (N_14837,N_14283,N_14397);
nor U14838 (N_14838,N_14077,N_14211);
and U14839 (N_14839,N_14033,N_13908);
xor U14840 (N_14840,N_13898,N_14277);
nand U14841 (N_14841,N_14039,N_14301);
or U14842 (N_14842,N_14343,N_13947);
xnor U14843 (N_14843,N_13931,N_14266);
xor U14844 (N_14844,N_13970,N_13912);
or U14845 (N_14845,N_14249,N_14282);
and U14846 (N_14846,N_14355,N_13812);
or U14847 (N_14847,N_14381,N_13914);
nand U14848 (N_14848,N_14194,N_14155);
and U14849 (N_14849,N_14304,N_14049);
and U14850 (N_14850,N_14307,N_14215);
nor U14851 (N_14851,N_14355,N_13868);
nand U14852 (N_14852,N_14267,N_13953);
nor U14853 (N_14853,N_14327,N_13918);
or U14854 (N_14854,N_13833,N_14340);
nand U14855 (N_14855,N_13927,N_14365);
nor U14856 (N_14856,N_14358,N_13929);
xnor U14857 (N_14857,N_13915,N_14082);
nor U14858 (N_14858,N_14289,N_14386);
xor U14859 (N_14859,N_14164,N_14193);
nand U14860 (N_14860,N_13802,N_14338);
nand U14861 (N_14861,N_14048,N_14314);
nand U14862 (N_14862,N_13960,N_13973);
or U14863 (N_14863,N_14193,N_13962);
nor U14864 (N_14864,N_13842,N_14295);
nor U14865 (N_14865,N_13837,N_13856);
nand U14866 (N_14866,N_13970,N_14093);
and U14867 (N_14867,N_14076,N_14302);
xor U14868 (N_14868,N_14197,N_13929);
xnor U14869 (N_14869,N_13950,N_13986);
or U14870 (N_14870,N_13839,N_14168);
xor U14871 (N_14871,N_14071,N_14369);
or U14872 (N_14872,N_14155,N_13833);
xnor U14873 (N_14873,N_13907,N_14327);
or U14874 (N_14874,N_13805,N_14285);
and U14875 (N_14875,N_13888,N_13959);
nand U14876 (N_14876,N_13827,N_14237);
xnor U14877 (N_14877,N_14185,N_14215);
xor U14878 (N_14878,N_14356,N_14333);
xnor U14879 (N_14879,N_14011,N_14365);
nand U14880 (N_14880,N_14104,N_14083);
or U14881 (N_14881,N_14136,N_14325);
nor U14882 (N_14882,N_13990,N_14105);
and U14883 (N_14883,N_13992,N_14340);
nand U14884 (N_14884,N_13978,N_14000);
nor U14885 (N_14885,N_13951,N_14112);
nand U14886 (N_14886,N_13855,N_13951);
and U14887 (N_14887,N_14364,N_14329);
nand U14888 (N_14888,N_14228,N_14335);
and U14889 (N_14889,N_14247,N_14296);
and U14890 (N_14890,N_14275,N_14281);
and U14891 (N_14891,N_14160,N_14297);
and U14892 (N_14892,N_14164,N_14361);
nand U14893 (N_14893,N_14330,N_13914);
nand U14894 (N_14894,N_13989,N_14186);
or U14895 (N_14895,N_14200,N_14229);
or U14896 (N_14896,N_14305,N_14284);
nor U14897 (N_14897,N_14032,N_14350);
or U14898 (N_14898,N_13963,N_13827);
and U14899 (N_14899,N_14355,N_14319);
nor U14900 (N_14900,N_14313,N_13952);
nor U14901 (N_14901,N_14387,N_14168);
xnor U14902 (N_14902,N_14142,N_14020);
nor U14903 (N_14903,N_14083,N_13956);
and U14904 (N_14904,N_13906,N_14057);
nand U14905 (N_14905,N_14373,N_13812);
or U14906 (N_14906,N_14345,N_13924);
nor U14907 (N_14907,N_14073,N_13853);
xnor U14908 (N_14908,N_14150,N_14042);
or U14909 (N_14909,N_13983,N_14067);
nor U14910 (N_14910,N_13813,N_13878);
and U14911 (N_14911,N_14006,N_14132);
nand U14912 (N_14912,N_14191,N_14141);
xnor U14913 (N_14913,N_13973,N_14045);
xnor U14914 (N_14914,N_14204,N_13840);
nor U14915 (N_14915,N_14040,N_14153);
nand U14916 (N_14916,N_14389,N_14285);
and U14917 (N_14917,N_14187,N_14394);
or U14918 (N_14918,N_13965,N_14058);
xnor U14919 (N_14919,N_14075,N_13963);
nor U14920 (N_14920,N_14050,N_14143);
nor U14921 (N_14921,N_14152,N_13982);
xor U14922 (N_14922,N_13918,N_14025);
nand U14923 (N_14923,N_13919,N_14188);
and U14924 (N_14924,N_13940,N_14265);
and U14925 (N_14925,N_13972,N_14225);
and U14926 (N_14926,N_14026,N_13943);
or U14927 (N_14927,N_13857,N_14281);
nand U14928 (N_14928,N_13803,N_14224);
nor U14929 (N_14929,N_14109,N_14125);
nor U14930 (N_14930,N_13822,N_14302);
nor U14931 (N_14931,N_14010,N_13852);
xor U14932 (N_14932,N_14316,N_13881);
xor U14933 (N_14933,N_14266,N_14011);
xor U14934 (N_14934,N_14003,N_14148);
xnor U14935 (N_14935,N_14212,N_14384);
or U14936 (N_14936,N_13850,N_14327);
and U14937 (N_14937,N_14280,N_14168);
nand U14938 (N_14938,N_14019,N_14296);
or U14939 (N_14939,N_14201,N_13948);
and U14940 (N_14940,N_13945,N_13973);
xor U14941 (N_14941,N_14293,N_14367);
xor U14942 (N_14942,N_14356,N_14240);
or U14943 (N_14943,N_13841,N_14274);
or U14944 (N_14944,N_14064,N_14166);
or U14945 (N_14945,N_13826,N_13943);
xor U14946 (N_14946,N_13841,N_14208);
and U14947 (N_14947,N_14079,N_14364);
and U14948 (N_14948,N_14265,N_13875);
nand U14949 (N_14949,N_13984,N_13874);
nor U14950 (N_14950,N_14314,N_13808);
and U14951 (N_14951,N_14097,N_14296);
xor U14952 (N_14952,N_14269,N_14290);
xor U14953 (N_14953,N_14226,N_13830);
or U14954 (N_14954,N_13934,N_14389);
or U14955 (N_14955,N_14074,N_14169);
or U14956 (N_14956,N_14090,N_14159);
nor U14957 (N_14957,N_14095,N_13861);
or U14958 (N_14958,N_13939,N_13881);
xor U14959 (N_14959,N_14330,N_13889);
xor U14960 (N_14960,N_13857,N_14264);
and U14961 (N_14961,N_14067,N_14070);
and U14962 (N_14962,N_14307,N_13955);
nor U14963 (N_14963,N_13869,N_14369);
xnor U14964 (N_14964,N_13844,N_14394);
nand U14965 (N_14965,N_14361,N_14349);
or U14966 (N_14966,N_14170,N_14058);
xor U14967 (N_14967,N_14207,N_13987);
and U14968 (N_14968,N_14143,N_13868);
nor U14969 (N_14969,N_14032,N_14057);
nand U14970 (N_14970,N_14350,N_14161);
and U14971 (N_14971,N_13809,N_14221);
xor U14972 (N_14972,N_14083,N_14281);
or U14973 (N_14973,N_14128,N_13842);
xor U14974 (N_14974,N_13894,N_14040);
and U14975 (N_14975,N_14386,N_14096);
nand U14976 (N_14976,N_14376,N_13972);
nand U14977 (N_14977,N_14234,N_14220);
and U14978 (N_14978,N_14395,N_14394);
nor U14979 (N_14979,N_14159,N_14032);
and U14980 (N_14980,N_14158,N_14244);
xor U14981 (N_14981,N_13918,N_13920);
and U14982 (N_14982,N_13858,N_14384);
nand U14983 (N_14983,N_13962,N_14197);
or U14984 (N_14984,N_13849,N_14154);
or U14985 (N_14985,N_13821,N_13842);
or U14986 (N_14986,N_14183,N_13816);
nand U14987 (N_14987,N_14186,N_13941);
or U14988 (N_14988,N_14009,N_13859);
or U14989 (N_14989,N_13958,N_13946);
and U14990 (N_14990,N_14110,N_14018);
and U14991 (N_14991,N_14315,N_14133);
nand U14992 (N_14992,N_14344,N_14255);
xor U14993 (N_14993,N_13944,N_13859);
nand U14994 (N_14994,N_13866,N_14195);
nor U14995 (N_14995,N_13812,N_14295);
or U14996 (N_14996,N_14184,N_14209);
and U14997 (N_14997,N_13808,N_14245);
and U14998 (N_14998,N_14095,N_14377);
or U14999 (N_14999,N_13991,N_14130);
nand U15000 (N_15000,N_14503,N_14913);
nor U15001 (N_15001,N_14853,N_14718);
and U15002 (N_15002,N_14854,N_14589);
or U15003 (N_15003,N_14551,N_14986);
and U15004 (N_15004,N_14792,N_14634);
or U15005 (N_15005,N_14538,N_14964);
nand U15006 (N_15006,N_14424,N_14895);
and U15007 (N_15007,N_14631,N_14745);
nand U15008 (N_15008,N_14507,N_14533);
or U15009 (N_15009,N_14418,N_14476);
xnor U15010 (N_15010,N_14413,N_14782);
and U15011 (N_15011,N_14681,N_14771);
and U15012 (N_15012,N_14547,N_14567);
nor U15013 (N_15013,N_14530,N_14889);
or U15014 (N_15014,N_14412,N_14740);
or U15015 (N_15015,N_14402,N_14788);
nor U15016 (N_15016,N_14861,N_14441);
xnor U15017 (N_15017,N_14756,N_14950);
and U15018 (N_15018,N_14744,N_14723);
xor U15019 (N_15019,N_14687,N_14463);
nand U15020 (N_15020,N_14557,N_14799);
and U15021 (N_15021,N_14961,N_14860);
or U15022 (N_15022,N_14443,N_14856);
or U15023 (N_15023,N_14651,N_14855);
nand U15024 (N_15024,N_14815,N_14935);
and U15025 (N_15025,N_14731,N_14603);
nor U15026 (N_15026,N_14900,N_14978);
nand U15027 (N_15027,N_14863,N_14554);
xnor U15028 (N_15028,N_14695,N_14505);
nand U15029 (N_15029,N_14991,N_14786);
and U15030 (N_15030,N_14619,N_14586);
nor U15031 (N_15031,N_14438,N_14422);
xnor U15032 (N_15032,N_14997,N_14578);
nor U15033 (N_15033,N_14852,N_14597);
xnor U15034 (N_15034,N_14667,N_14694);
xnor U15035 (N_15035,N_14563,N_14436);
nor U15036 (N_15036,N_14657,N_14433);
and U15037 (N_15037,N_14618,N_14529);
or U15038 (N_15038,N_14638,N_14420);
and U15039 (N_15039,N_14918,N_14939);
nand U15040 (N_15040,N_14962,N_14887);
or U15041 (N_15041,N_14437,N_14704);
and U15042 (N_15042,N_14558,N_14481);
nor U15043 (N_15043,N_14548,N_14595);
xnor U15044 (N_15044,N_14838,N_14601);
xnor U15045 (N_15045,N_14905,N_14751);
nand U15046 (N_15046,N_14800,N_14886);
nand U15047 (N_15047,N_14693,N_14980);
nor U15048 (N_15048,N_14791,N_14864);
nor U15049 (N_15049,N_14573,N_14661);
nand U15050 (N_15050,N_14707,N_14931);
or U15051 (N_15051,N_14896,N_14600);
nand U15052 (N_15052,N_14585,N_14545);
or U15053 (N_15053,N_14726,N_14671);
xnor U15054 (N_15054,N_14472,N_14921);
or U15055 (N_15055,N_14881,N_14859);
and U15056 (N_15056,N_14591,N_14793);
and U15057 (N_15057,N_14679,N_14839);
nor U15058 (N_15058,N_14974,N_14449);
or U15059 (N_15059,N_14957,N_14807);
xor U15060 (N_15060,N_14621,N_14665);
and U15061 (N_15061,N_14592,N_14893);
and U15062 (N_15062,N_14453,N_14627);
and U15063 (N_15063,N_14570,N_14459);
or U15064 (N_15064,N_14720,N_14970);
nand U15065 (N_15065,N_14491,N_14952);
xnor U15066 (N_15066,N_14524,N_14717);
nand U15067 (N_15067,N_14611,N_14419);
xor U15068 (N_15068,N_14865,N_14596);
and U15069 (N_15069,N_14408,N_14810);
and U15070 (N_15070,N_14743,N_14902);
xor U15071 (N_15071,N_14527,N_14645);
nand U15072 (N_15072,N_14625,N_14605);
nor U15073 (N_15073,N_14653,N_14663);
nor U15074 (N_15074,N_14564,N_14655);
nand U15075 (N_15075,N_14836,N_14470);
xnor U15076 (N_15076,N_14516,N_14812);
or U15077 (N_15077,N_14517,N_14827);
and U15078 (N_15078,N_14696,N_14892);
or U15079 (N_15079,N_14942,N_14879);
nor U15080 (N_15080,N_14811,N_14832);
nand U15081 (N_15081,N_14672,N_14562);
nand U15082 (N_15082,N_14725,N_14479);
or U15083 (N_15083,N_14849,N_14737);
nor U15084 (N_15084,N_14427,N_14506);
nand U15085 (N_15085,N_14803,N_14561);
and U15086 (N_15086,N_14708,N_14642);
or U15087 (N_15087,N_14835,N_14568);
nand U15088 (N_15088,N_14794,N_14727);
nand U15089 (N_15089,N_14778,N_14712);
nor U15090 (N_15090,N_14483,N_14843);
xor U15091 (N_15091,N_14415,N_14898);
and U15092 (N_15092,N_14641,N_14903);
xor U15093 (N_15093,N_14757,N_14440);
or U15094 (N_15094,N_14569,N_14714);
or U15095 (N_15095,N_14783,N_14465);
nand U15096 (N_15096,N_14456,N_14654);
nand U15097 (N_15097,N_14938,N_14878);
nand U15098 (N_15098,N_14546,N_14508);
xnor U15099 (N_15099,N_14581,N_14457);
and U15100 (N_15100,N_14721,N_14949);
nand U15101 (N_15101,N_14553,N_14475);
nor U15102 (N_15102,N_14846,N_14594);
nand U15103 (N_15103,N_14409,N_14729);
nand U15104 (N_15104,N_14877,N_14790);
and U15105 (N_15105,N_14405,N_14742);
or U15106 (N_15106,N_14588,N_14640);
and U15107 (N_15107,N_14431,N_14749);
xnor U15108 (N_15108,N_14981,N_14784);
or U15109 (N_15109,N_14403,N_14922);
or U15110 (N_15110,N_14710,N_14700);
nor U15111 (N_15111,N_14871,N_14444);
xor U15112 (N_15112,N_14460,N_14531);
and U15113 (N_15113,N_14802,N_14822);
nor U15114 (N_15114,N_14628,N_14658);
nand U15115 (N_15115,N_14761,N_14776);
nand U15116 (N_15116,N_14501,N_14801);
xor U15117 (N_15117,N_14614,N_14495);
nor U15118 (N_15118,N_14764,N_14432);
nor U15119 (N_15119,N_14539,N_14484);
nor U15120 (N_15120,N_14450,N_14883);
and U15121 (N_15121,N_14825,N_14834);
and U15122 (N_15122,N_14713,N_14880);
or U15123 (N_15123,N_14537,N_14647);
or U15124 (N_15124,N_14979,N_14994);
nor U15125 (N_15125,N_14795,N_14798);
xnor U15126 (N_15126,N_14455,N_14682);
and U15127 (N_15127,N_14552,N_14940);
or U15128 (N_15128,N_14987,N_14674);
and U15129 (N_15129,N_14866,N_14650);
xor U15130 (N_15130,N_14623,N_14543);
nand U15131 (N_15131,N_14604,N_14451);
and U15132 (N_15132,N_14519,N_14908);
nand U15133 (N_15133,N_14488,N_14872);
nor U15134 (N_15134,N_14643,N_14504);
xnor U15135 (N_15135,N_14662,N_14929);
nor U15136 (N_15136,N_14609,N_14933);
and U15137 (N_15137,N_14464,N_14728);
and U15138 (N_15138,N_14781,N_14549);
and U15139 (N_15139,N_14703,N_14818);
nor U15140 (N_15140,N_14960,N_14709);
or U15141 (N_15141,N_14789,N_14840);
and U15142 (N_15142,N_14613,N_14577);
or U15143 (N_15143,N_14733,N_14497);
nor U15144 (N_15144,N_14528,N_14458);
nor U15145 (N_15145,N_14705,N_14753);
xor U15146 (N_15146,N_14848,N_14471);
nand U15147 (N_15147,N_14820,N_14411);
or U15148 (N_15148,N_14435,N_14500);
and U15149 (N_15149,N_14817,N_14924);
and U15150 (N_15150,N_14829,N_14862);
nor U15151 (N_15151,N_14758,N_14514);
nor U15152 (N_15152,N_14785,N_14511);
xnor U15153 (N_15153,N_14824,N_14912);
xor U15154 (N_15154,N_14639,N_14899);
xor U15155 (N_15155,N_14697,N_14636);
xor U15156 (N_15156,N_14485,N_14747);
nor U15157 (N_15157,N_14947,N_14869);
nor U15158 (N_15158,N_14915,N_14664);
nand U15159 (N_15159,N_14425,N_14828);
xnor U15160 (N_15160,N_14755,N_14885);
nor U15161 (N_15161,N_14735,N_14423);
and U15162 (N_15162,N_14926,N_14582);
or U15163 (N_15163,N_14620,N_14610);
xor U15164 (N_15164,N_14487,N_14752);
nor U15165 (N_15165,N_14525,N_14909);
and U15166 (N_15166,N_14956,N_14477);
nand U15167 (N_15167,N_14739,N_14617);
nand U15168 (N_15168,N_14668,N_14816);
nor U15169 (N_15169,N_14711,N_14689);
nor U15170 (N_15170,N_14478,N_14722);
or U15171 (N_15171,N_14951,N_14809);
or U15172 (N_15172,N_14576,N_14945);
and U15173 (N_15173,N_14648,N_14917);
and U15174 (N_15174,N_14536,N_14421);
nor U15175 (N_15175,N_14630,N_14906);
and U15176 (N_15176,N_14489,N_14968);
or U15177 (N_15177,N_14482,N_14948);
nand U15178 (N_15178,N_14738,N_14649);
nand U15179 (N_15179,N_14890,N_14719);
and U15180 (N_15180,N_14990,N_14923);
nand U15181 (N_15181,N_14996,N_14426);
nor U15182 (N_15182,N_14414,N_14873);
and U15183 (N_15183,N_14959,N_14901);
and U15184 (N_15184,N_14540,N_14897);
nor U15185 (N_15185,N_14676,N_14767);
or U15186 (N_15186,N_14870,N_14686);
and U15187 (N_15187,N_14925,N_14891);
and U15188 (N_15188,N_14644,N_14876);
nor U15189 (N_15189,N_14646,N_14982);
or U15190 (N_15190,N_14407,N_14599);
nand U15191 (N_15191,N_14404,N_14919);
nand U15192 (N_15192,N_14928,N_14984);
xnor U15193 (N_15193,N_14606,N_14448);
xnor U15194 (N_15194,N_14760,N_14401);
or U15195 (N_15195,N_14916,N_14842);
and U15196 (N_15196,N_14583,N_14715);
or U15197 (N_15197,N_14584,N_14833);
nor U15198 (N_15198,N_14821,N_14512);
xnor U15199 (N_15199,N_14868,N_14565);
nor U15200 (N_15200,N_14635,N_14963);
nor U15201 (N_15201,N_14805,N_14773);
nand U15202 (N_15202,N_14754,N_14999);
xor U15203 (N_15203,N_14851,N_14943);
nor U15204 (N_15204,N_14995,N_14607);
or U15205 (N_15205,N_14777,N_14701);
nand U15206 (N_15206,N_14845,N_14509);
or U15207 (N_15207,N_14468,N_14779);
nand U15208 (N_15208,N_14461,N_14541);
and U15209 (N_15209,N_14660,N_14823);
or U15210 (N_15210,N_14480,N_14692);
and U15211 (N_15211,N_14847,N_14493);
nor U15212 (N_15212,N_14965,N_14542);
nand U15213 (N_15213,N_14574,N_14699);
or U15214 (N_15214,N_14882,N_14615);
xor U15215 (N_15215,N_14819,N_14904);
xor U15216 (N_15216,N_14944,N_14813);
nand U15217 (N_15217,N_14598,N_14804);
and U15218 (N_15218,N_14410,N_14958);
xnor U15219 (N_15219,N_14555,N_14732);
nand U15220 (N_15220,N_14808,N_14972);
and U15221 (N_15221,N_14983,N_14560);
or U15222 (N_15222,N_14602,N_14550);
nand U15223 (N_15223,N_14520,N_14766);
xnor U15224 (N_15224,N_14989,N_14417);
or U15225 (N_15225,N_14772,N_14927);
and U15226 (N_15226,N_14806,N_14690);
nand U15227 (N_15227,N_14685,N_14748);
xnor U15228 (N_15228,N_14666,N_14988);
and U15229 (N_15229,N_14716,N_14656);
xor U15230 (N_15230,N_14741,N_14490);
or U15231 (N_15231,N_14434,N_14706);
xor U15232 (N_15232,N_14797,N_14734);
xnor U15233 (N_15233,N_14499,N_14626);
xor U15234 (N_15234,N_14932,N_14494);
nor U15235 (N_15235,N_14850,N_14775);
and U15236 (N_15236,N_14442,N_14774);
and U15237 (N_15237,N_14616,N_14580);
xor U15238 (N_15238,N_14910,N_14867);
xnor U15239 (N_15239,N_14452,N_14612);
xor U15240 (N_15240,N_14724,N_14759);
or U15241 (N_15241,N_14518,N_14780);
nor U15242 (N_15242,N_14429,N_14914);
nand U15243 (N_15243,N_14966,N_14954);
xnor U15244 (N_15244,N_14985,N_14688);
or U15245 (N_15245,N_14571,N_14765);
nor U15246 (N_15246,N_14579,N_14526);
or U15247 (N_15247,N_14502,N_14416);
and U15248 (N_15248,N_14447,N_14894);
xor U15249 (N_15249,N_14521,N_14572);
and U15250 (N_15250,N_14969,N_14515);
and U15251 (N_15251,N_14467,N_14454);
or U15252 (N_15252,N_14763,N_14953);
nand U15253 (N_15253,N_14474,N_14633);
or U15254 (N_15254,N_14532,N_14875);
xnor U15255 (N_15255,N_14566,N_14769);
and U15256 (N_15256,N_14973,N_14770);
nor U15257 (N_15257,N_14683,N_14466);
or U15258 (N_15258,N_14858,N_14907);
or U15259 (N_15259,N_14977,N_14670);
xor U15260 (N_15260,N_14993,N_14608);
nand U15261 (N_15261,N_14637,N_14691);
nor U15262 (N_15262,N_14837,N_14787);
xnor U15263 (N_15263,N_14874,N_14675);
xor U15264 (N_15264,N_14857,N_14469);
xnor U15265 (N_15265,N_14746,N_14677);
nand U15266 (N_15266,N_14522,N_14702);
nor U15267 (N_15267,N_14523,N_14439);
and U15268 (N_15268,N_14678,N_14445);
nand U15269 (N_15269,N_14462,N_14534);
and U15270 (N_15270,N_14652,N_14629);
xor U15271 (N_15271,N_14684,N_14473);
nand U15272 (N_15272,N_14830,N_14698);
and U15273 (N_15273,N_14934,N_14510);
nand U15274 (N_15274,N_14998,N_14673);
nor U15275 (N_15275,N_14911,N_14730);
xor U15276 (N_15276,N_14920,N_14400);
nor U15277 (N_15277,N_14768,N_14680);
or U15278 (N_15278,N_14750,N_14622);
nand U15279 (N_15279,N_14992,N_14593);
and U15280 (N_15280,N_14888,N_14575);
nor U15281 (N_15281,N_14446,N_14967);
xor U15282 (N_15282,N_14796,N_14513);
nand U15283 (N_15283,N_14669,N_14971);
and U15284 (N_15284,N_14632,N_14936);
xnor U15285 (N_15285,N_14535,N_14976);
and U15286 (N_15286,N_14762,N_14486);
xnor U15287 (N_15287,N_14937,N_14406);
or U15288 (N_15288,N_14624,N_14559);
nand U15289 (N_15289,N_14659,N_14955);
nor U15290 (N_15290,N_14428,N_14930);
nand U15291 (N_15291,N_14430,N_14496);
nor U15292 (N_15292,N_14975,N_14826);
nor U15293 (N_15293,N_14884,N_14590);
and U15294 (N_15294,N_14736,N_14498);
xnor U15295 (N_15295,N_14492,N_14814);
or U15296 (N_15296,N_14841,N_14556);
and U15297 (N_15297,N_14587,N_14946);
xor U15298 (N_15298,N_14844,N_14544);
and U15299 (N_15299,N_14941,N_14831);
and U15300 (N_15300,N_14568,N_14574);
xnor U15301 (N_15301,N_14894,N_14872);
or U15302 (N_15302,N_14614,N_14586);
xor U15303 (N_15303,N_14739,N_14563);
nand U15304 (N_15304,N_14424,N_14891);
and U15305 (N_15305,N_14884,N_14582);
or U15306 (N_15306,N_14963,N_14685);
and U15307 (N_15307,N_14625,N_14561);
and U15308 (N_15308,N_14623,N_14533);
xnor U15309 (N_15309,N_14841,N_14570);
and U15310 (N_15310,N_14875,N_14996);
nor U15311 (N_15311,N_14548,N_14539);
and U15312 (N_15312,N_14985,N_14837);
and U15313 (N_15313,N_14855,N_14929);
nand U15314 (N_15314,N_14540,N_14498);
nor U15315 (N_15315,N_14874,N_14875);
nor U15316 (N_15316,N_14500,N_14720);
or U15317 (N_15317,N_14758,N_14487);
nor U15318 (N_15318,N_14818,N_14855);
xnor U15319 (N_15319,N_14936,N_14780);
nor U15320 (N_15320,N_14622,N_14451);
and U15321 (N_15321,N_14837,N_14968);
or U15322 (N_15322,N_14673,N_14418);
nand U15323 (N_15323,N_14969,N_14681);
or U15324 (N_15324,N_14657,N_14628);
nand U15325 (N_15325,N_14882,N_14659);
and U15326 (N_15326,N_14820,N_14572);
nor U15327 (N_15327,N_14865,N_14485);
nor U15328 (N_15328,N_14477,N_14987);
nor U15329 (N_15329,N_14416,N_14965);
nand U15330 (N_15330,N_14871,N_14778);
nor U15331 (N_15331,N_14540,N_14425);
and U15332 (N_15332,N_14910,N_14606);
xnor U15333 (N_15333,N_14900,N_14994);
nand U15334 (N_15334,N_14792,N_14755);
or U15335 (N_15335,N_14720,N_14939);
nand U15336 (N_15336,N_14802,N_14947);
and U15337 (N_15337,N_14767,N_14558);
and U15338 (N_15338,N_14945,N_14949);
nand U15339 (N_15339,N_14598,N_14903);
or U15340 (N_15340,N_14508,N_14847);
nor U15341 (N_15341,N_14550,N_14783);
and U15342 (N_15342,N_14858,N_14604);
or U15343 (N_15343,N_14656,N_14904);
or U15344 (N_15344,N_14438,N_14949);
xor U15345 (N_15345,N_14462,N_14729);
nand U15346 (N_15346,N_14448,N_14656);
or U15347 (N_15347,N_14569,N_14462);
nor U15348 (N_15348,N_14532,N_14425);
nand U15349 (N_15349,N_14615,N_14699);
or U15350 (N_15350,N_14664,N_14672);
or U15351 (N_15351,N_14635,N_14717);
xor U15352 (N_15352,N_14917,N_14634);
and U15353 (N_15353,N_14460,N_14789);
or U15354 (N_15354,N_14633,N_14982);
or U15355 (N_15355,N_14764,N_14518);
nand U15356 (N_15356,N_14480,N_14850);
xnor U15357 (N_15357,N_14642,N_14521);
nand U15358 (N_15358,N_14975,N_14588);
nand U15359 (N_15359,N_14472,N_14538);
or U15360 (N_15360,N_14643,N_14606);
or U15361 (N_15361,N_14786,N_14648);
nand U15362 (N_15362,N_14870,N_14614);
xor U15363 (N_15363,N_14546,N_14640);
nor U15364 (N_15364,N_14734,N_14761);
nor U15365 (N_15365,N_14632,N_14768);
nand U15366 (N_15366,N_14625,N_14731);
nand U15367 (N_15367,N_14644,N_14488);
xnor U15368 (N_15368,N_14980,N_14773);
nor U15369 (N_15369,N_14887,N_14837);
xor U15370 (N_15370,N_14876,N_14889);
or U15371 (N_15371,N_14506,N_14546);
and U15372 (N_15372,N_14692,N_14472);
or U15373 (N_15373,N_14575,N_14413);
nor U15374 (N_15374,N_14744,N_14512);
xnor U15375 (N_15375,N_14871,N_14530);
nor U15376 (N_15376,N_14589,N_14812);
or U15377 (N_15377,N_14697,N_14542);
and U15378 (N_15378,N_14765,N_14659);
xor U15379 (N_15379,N_14757,N_14944);
or U15380 (N_15380,N_14931,N_14930);
xor U15381 (N_15381,N_14947,N_14936);
xnor U15382 (N_15382,N_14916,N_14946);
nand U15383 (N_15383,N_14578,N_14632);
nand U15384 (N_15384,N_14647,N_14994);
and U15385 (N_15385,N_14692,N_14995);
nor U15386 (N_15386,N_14865,N_14694);
and U15387 (N_15387,N_14713,N_14714);
nor U15388 (N_15388,N_14792,N_14782);
or U15389 (N_15389,N_14858,N_14964);
or U15390 (N_15390,N_14517,N_14672);
nand U15391 (N_15391,N_14433,N_14639);
or U15392 (N_15392,N_14405,N_14664);
and U15393 (N_15393,N_14592,N_14694);
or U15394 (N_15394,N_14890,N_14969);
and U15395 (N_15395,N_14490,N_14709);
xor U15396 (N_15396,N_14479,N_14403);
xor U15397 (N_15397,N_14876,N_14815);
xor U15398 (N_15398,N_14972,N_14747);
nand U15399 (N_15399,N_14494,N_14874);
nand U15400 (N_15400,N_14552,N_14448);
or U15401 (N_15401,N_14696,N_14869);
and U15402 (N_15402,N_14500,N_14793);
xor U15403 (N_15403,N_14513,N_14759);
and U15404 (N_15404,N_14514,N_14868);
xor U15405 (N_15405,N_14953,N_14444);
xor U15406 (N_15406,N_14865,N_14461);
xnor U15407 (N_15407,N_14533,N_14845);
nand U15408 (N_15408,N_14599,N_14503);
nor U15409 (N_15409,N_14444,N_14412);
nand U15410 (N_15410,N_14882,N_14750);
or U15411 (N_15411,N_14850,N_14801);
nand U15412 (N_15412,N_14547,N_14934);
nand U15413 (N_15413,N_14836,N_14888);
and U15414 (N_15414,N_14412,N_14646);
xor U15415 (N_15415,N_14716,N_14937);
xnor U15416 (N_15416,N_14982,N_14892);
or U15417 (N_15417,N_14607,N_14614);
nand U15418 (N_15418,N_14826,N_14756);
nand U15419 (N_15419,N_14858,N_14937);
or U15420 (N_15420,N_14533,N_14620);
or U15421 (N_15421,N_14751,N_14608);
or U15422 (N_15422,N_14496,N_14877);
and U15423 (N_15423,N_14523,N_14716);
xor U15424 (N_15424,N_14697,N_14454);
xor U15425 (N_15425,N_14473,N_14467);
and U15426 (N_15426,N_14699,N_14483);
nor U15427 (N_15427,N_14871,N_14797);
and U15428 (N_15428,N_14499,N_14432);
or U15429 (N_15429,N_14921,N_14654);
and U15430 (N_15430,N_14534,N_14514);
xor U15431 (N_15431,N_14602,N_14816);
or U15432 (N_15432,N_14710,N_14757);
and U15433 (N_15433,N_14468,N_14527);
nor U15434 (N_15434,N_14683,N_14980);
or U15435 (N_15435,N_14758,N_14603);
nand U15436 (N_15436,N_14845,N_14732);
and U15437 (N_15437,N_14534,N_14516);
and U15438 (N_15438,N_14519,N_14433);
nor U15439 (N_15439,N_14606,N_14827);
and U15440 (N_15440,N_14506,N_14753);
xnor U15441 (N_15441,N_14662,N_14409);
or U15442 (N_15442,N_14422,N_14597);
nor U15443 (N_15443,N_14715,N_14617);
nor U15444 (N_15444,N_14485,N_14414);
and U15445 (N_15445,N_14778,N_14646);
nand U15446 (N_15446,N_14466,N_14782);
nand U15447 (N_15447,N_14941,N_14872);
and U15448 (N_15448,N_14675,N_14816);
and U15449 (N_15449,N_14648,N_14635);
nand U15450 (N_15450,N_14438,N_14509);
or U15451 (N_15451,N_14689,N_14826);
xnor U15452 (N_15452,N_14923,N_14882);
and U15453 (N_15453,N_14767,N_14745);
nor U15454 (N_15454,N_14950,N_14662);
nor U15455 (N_15455,N_14856,N_14419);
or U15456 (N_15456,N_14641,N_14652);
nand U15457 (N_15457,N_14448,N_14922);
or U15458 (N_15458,N_14601,N_14686);
or U15459 (N_15459,N_14866,N_14731);
or U15460 (N_15460,N_14519,N_14703);
nor U15461 (N_15461,N_14977,N_14591);
or U15462 (N_15462,N_14584,N_14875);
nor U15463 (N_15463,N_14864,N_14446);
and U15464 (N_15464,N_14484,N_14606);
nand U15465 (N_15465,N_14413,N_14991);
xor U15466 (N_15466,N_14609,N_14798);
xnor U15467 (N_15467,N_14603,N_14838);
and U15468 (N_15468,N_14501,N_14607);
or U15469 (N_15469,N_14424,N_14938);
or U15470 (N_15470,N_14602,N_14673);
xor U15471 (N_15471,N_14426,N_14766);
or U15472 (N_15472,N_14416,N_14634);
nand U15473 (N_15473,N_14985,N_14982);
and U15474 (N_15474,N_14477,N_14770);
nand U15475 (N_15475,N_14743,N_14967);
or U15476 (N_15476,N_14536,N_14526);
xor U15477 (N_15477,N_14934,N_14694);
or U15478 (N_15478,N_14478,N_14801);
and U15479 (N_15479,N_14528,N_14851);
nand U15480 (N_15480,N_14726,N_14649);
nor U15481 (N_15481,N_14848,N_14885);
xor U15482 (N_15482,N_14843,N_14807);
nor U15483 (N_15483,N_14569,N_14633);
xnor U15484 (N_15484,N_14888,N_14778);
xor U15485 (N_15485,N_14891,N_14605);
and U15486 (N_15486,N_14845,N_14750);
and U15487 (N_15487,N_14767,N_14619);
xnor U15488 (N_15488,N_14791,N_14488);
nand U15489 (N_15489,N_14469,N_14533);
nor U15490 (N_15490,N_14891,N_14854);
or U15491 (N_15491,N_14523,N_14648);
and U15492 (N_15492,N_14652,N_14943);
nor U15493 (N_15493,N_14968,N_14766);
xnor U15494 (N_15494,N_14446,N_14744);
nand U15495 (N_15495,N_14512,N_14886);
and U15496 (N_15496,N_14621,N_14739);
xnor U15497 (N_15497,N_14632,N_14764);
nor U15498 (N_15498,N_14892,N_14907);
xnor U15499 (N_15499,N_14567,N_14911);
nand U15500 (N_15500,N_14434,N_14842);
nand U15501 (N_15501,N_14694,N_14852);
nand U15502 (N_15502,N_14830,N_14548);
xnor U15503 (N_15503,N_14405,N_14833);
xor U15504 (N_15504,N_14527,N_14824);
xnor U15505 (N_15505,N_14719,N_14723);
nand U15506 (N_15506,N_14735,N_14508);
nor U15507 (N_15507,N_14562,N_14803);
nand U15508 (N_15508,N_14481,N_14736);
nand U15509 (N_15509,N_14765,N_14608);
or U15510 (N_15510,N_14678,N_14641);
or U15511 (N_15511,N_14614,N_14565);
xnor U15512 (N_15512,N_14715,N_14447);
or U15513 (N_15513,N_14481,N_14490);
and U15514 (N_15514,N_14439,N_14646);
nor U15515 (N_15515,N_14927,N_14445);
nand U15516 (N_15516,N_14450,N_14989);
or U15517 (N_15517,N_14973,N_14504);
nor U15518 (N_15518,N_14758,N_14694);
and U15519 (N_15519,N_14931,N_14850);
or U15520 (N_15520,N_14916,N_14459);
nor U15521 (N_15521,N_14823,N_14863);
xnor U15522 (N_15522,N_14934,N_14845);
xnor U15523 (N_15523,N_14436,N_14994);
and U15524 (N_15524,N_14483,N_14583);
nor U15525 (N_15525,N_14609,N_14863);
xor U15526 (N_15526,N_14558,N_14480);
or U15527 (N_15527,N_14537,N_14559);
and U15528 (N_15528,N_14992,N_14553);
nor U15529 (N_15529,N_14996,N_14847);
nand U15530 (N_15530,N_14497,N_14449);
nor U15531 (N_15531,N_14663,N_14580);
xor U15532 (N_15532,N_14784,N_14980);
xnor U15533 (N_15533,N_14851,N_14940);
or U15534 (N_15534,N_14812,N_14595);
or U15535 (N_15535,N_14563,N_14777);
nand U15536 (N_15536,N_14581,N_14912);
and U15537 (N_15537,N_14569,N_14454);
or U15538 (N_15538,N_14663,N_14924);
or U15539 (N_15539,N_14630,N_14889);
and U15540 (N_15540,N_14893,N_14498);
or U15541 (N_15541,N_14972,N_14936);
nand U15542 (N_15542,N_14710,N_14750);
nand U15543 (N_15543,N_14935,N_14544);
nor U15544 (N_15544,N_14978,N_14729);
xor U15545 (N_15545,N_14916,N_14855);
xor U15546 (N_15546,N_14602,N_14703);
and U15547 (N_15547,N_14514,N_14403);
xnor U15548 (N_15548,N_14993,N_14976);
or U15549 (N_15549,N_14907,N_14903);
or U15550 (N_15550,N_14908,N_14506);
xor U15551 (N_15551,N_14670,N_14489);
nand U15552 (N_15552,N_14686,N_14727);
nor U15553 (N_15553,N_14937,N_14413);
or U15554 (N_15554,N_14707,N_14608);
or U15555 (N_15555,N_14973,N_14700);
and U15556 (N_15556,N_14461,N_14994);
xor U15557 (N_15557,N_14443,N_14890);
or U15558 (N_15558,N_14612,N_14601);
nor U15559 (N_15559,N_14832,N_14956);
or U15560 (N_15560,N_14818,N_14959);
xor U15561 (N_15561,N_14702,N_14461);
xor U15562 (N_15562,N_14470,N_14890);
xnor U15563 (N_15563,N_14757,N_14722);
nor U15564 (N_15564,N_14649,N_14907);
or U15565 (N_15565,N_14787,N_14465);
and U15566 (N_15566,N_14857,N_14773);
xor U15567 (N_15567,N_14634,N_14527);
nand U15568 (N_15568,N_14934,N_14548);
nor U15569 (N_15569,N_14918,N_14468);
and U15570 (N_15570,N_14749,N_14908);
and U15571 (N_15571,N_14684,N_14457);
and U15572 (N_15572,N_14854,N_14839);
and U15573 (N_15573,N_14745,N_14576);
or U15574 (N_15574,N_14480,N_14778);
or U15575 (N_15575,N_14577,N_14943);
and U15576 (N_15576,N_14476,N_14626);
nand U15577 (N_15577,N_14577,N_14456);
nor U15578 (N_15578,N_14504,N_14451);
nor U15579 (N_15579,N_14639,N_14719);
nor U15580 (N_15580,N_14977,N_14590);
xnor U15581 (N_15581,N_14451,N_14616);
or U15582 (N_15582,N_14611,N_14819);
nor U15583 (N_15583,N_14772,N_14834);
nand U15584 (N_15584,N_14894,N_14728);
xnor U15585 (N_15585,N_14813,N_14857);
or U15586 (N_15586,N_14571,N_14542);
and U15587 (N_15587,N_14765,N_14817);
xnor U15588 (N_15588,N_14827,N_14493);
and U15589 (N_15589,N_14798,N_14841);
xnor U15590 (N_15590,N_14857,N_14878);
nor U15591 (N_15591,N_14966,N_14859);
or U15592 (N_15592,N_14554,N_14421);
or U15593 (N_15593,N_14445,N_14585);
nor U15594 (N_15594,N_14862,N_14763);
and U15595 (N_15595,N_14432,N_14745);
xor U15596 (N_15596,N_14779,N_14873);
and U15597 (N_15597,N_14453,N_14483);
nand U15598 (N_15598,N_14715,N_14441);
nor U15599 (N_15599,N_14608,N_14571);
and U15600 (N_15600,N_15373,N_15427);
and U15601 (N_15601,N_15128,N_15514);
nor U15602 (N_15602,N_15038,N_15308);
xor U15603 (N_15603,N_15421,N_15026);
nor U15604 (N_15604,N_15178,N_15077);
nor U15605 (N_15605,N_15585,N_15235);
xnor U15606 (N_15606,N_15206,N_15096);
xnor U15607 (N_15607,N_15299,N_15356);
nor U15608 (N_15608,N_15247,N_15076);
or U15609 (N_15609,N_15036,N_15069);
nand U15610 (N_15610,N_15030,N_15536);
and U15611 (N_15611,N_15365,N_15366);
and U15612 (N_15612,N_15535,N_15326);
nor U15613 (N_15613,N_15542,N_15011);
nand U15614 (N_15614,N_15462,N_15009);
xor U15615 (N_15615,N_15100,N_15199);
and U15616 (N_15616,N_15147,N_15507);
xnor U15617 (N_15617,N_15483,N_15437);
nor U15618 (N_15618,N_15088,N_15598);
or U15619 (N_15619,N_15538,N_15564);
nor U15620 (N_15620,N_15043,N_15496);
and U15621 (N_15621,N_15313,N_15281);
nor U15622 (N_15622,N_15397,N_15590);
nor U15623 (N_15623,N_15052,N_15372);
and U15624 (N_15624,N_15101,N_15423);
nor U15625 (N_15625,N_15544,N_15436);
nor U15626 (N_15626,N_15388,N_15217);
or U15627 (N_15627,N_15249,N_15470);
or U15628 (N_15628,N_15449,N_15228);
nor U15629 (N_15629,N_15552,N_15198);
xor U15630 (N_15630,N_15021,N_15041);
xnor U15631 (N_15631,N_15288,N_15401);
and U15632 (N_15632,N_15229,N_15018);
xor U15633 (N_15633,N_15475,N_15334);
xor U15634 (N_15634,N_15068,N_15195);
nand U15635 (N_15635,N_15551,N_15042);
nor U15636 (N_15636,N_15580,N_15087);
nand U15637 (N_15637,N_15261,N_15255);
nor U15638 (N_15638,N_15520,N_15426);
and U15639 (N_15639,N_15224,N_15553);
or U15640 (N_15640,N_15345,N_15211);
and U15641 (N_15641,N_15588,N_15127);
or U15642 (N_15642,N_15303,N_15025);
nor U15643 (N_15643,N_15435,N_15502);
nor U15644 (N_15644,N_15204,N_15560);
xor U15645 (N_15645,N_15010,N_15444);
nor U15646 (N_15646,N_15186,N_15152);
or U15647 (N_15647,N_15368,N_15486);
xor U15648 (N_15648,N_15484,N_15425);
and U15649 (N_15649,N_15504,N_15503);
and U15650 (N_15650,N_15254,N_15434);
nor U15651 (N_15651,N_15293,N_15012);
nor U15652 (N_15652,N_15364,N_15051);
xnor U15653 (N_15653,N_15192,N_15099);
or U15654 (N_15654,N_15080,N_15294);
nor U15655 (N_15655,N_15278,N_15476);
nor U15656 (N_15656,N_15323,N_15005);
xnor U15657 (N_15657,N_15120,N_15180);
and U15658 (N_15658,N_15457,N_15349);
nor U15659 (N_15659,N_15493,N_15413);
nand U15660 (N_15660,N_15572,N_15311);
and U15661 (N_15661,N_15122,N_15407);
nor U15662 (N_15662,N_15357,N_15557);
nor U15663 (N_15663,N_15379,N_15257);
nand U15664 (N_15664,N_15221,N_15424);
or U15665 (N_15665,N_15074,N_15545);
and U15666 (N_15666,N_15082,N_15156);
or U15667 (N_15667,N_15008,N_15202);
nor U15668 (N_15668,N_15550,N_15078);
nand U15669 (N_15669,N_15050,N_15587);
and U15670 (N_15670,N_15184,N_15153);
and U15671 (N_15671,N_15145,N_15451);
and U15672 (N_15672,N_15328,N_15273);
or U15673 (N_15673,N_15055,N_15512);
nand U15674 (N_15674,N_15213,N_15582);
nor U15675 (N_15675,N_15060,N_15419);
nor U15676 (N_15676,N_15300,N_15515);
xor U15677 (N_15677,N_15044,N_15154);
nor U15678 (N_15678,N_15286,N_15363);
or U15679 (N_15679,N_15280,N_15347);
or U15680 (N_15680,N_15385,N_15464);
xnor U15681 (N_15681,N_15392,N_15494);
nand U15682 (N_15682,N_15239,N_15028);
xnor U15683 (N_15683,N_15495,N_15343);
xnor U15684 (N_15684,N_15162,N_15137);
nor U15685 (N_15685,N_15310,N_15505);
and U15686 (N_15686,N_15595,N_15134);
nor U15687 (N_15687,N_15081,N_15024);
nand U15688 (N_15688,N_15252,N_15523);
and U15689 (N_15689,N_15270,N_15090);
nand U15690 (N_15690,N_15161,N_15117);
nor U15691 (N_15691,N_15139,N_15471);
xor U15692 (N_15692,N_15032,N_15188);
xor U15693 (N_15693,N_15583,N_15375);
nor U15694 (N_15694,N_15467,N_15194);
xor U15695 (N_15695,N_15584,N_15168);
nand U15696 (N_15696,N_15321,N_15091);
or U15697 (N_15697,N_15408,N_15358);
nor U15698 (N_15698,N_15004,N_15193);
nand U15699 (N_15699,N_15561,N_15489);
or U15700 (N_15700,N_15304,N_15348);
and U15701 (N_15701,N_15015,N_15525);
and U15702 (N_15702,N_15260,N_15377);
nor U15703 (N_15703,N_15067,N_15400);
and U15704 (N_15704,N_15001,N_15244);
nor U15705 (N_15705,N_15532,N_15405);
or U15706 (N_15706,N_15465,N_15170);
xnor U15707 (N_15707,N_15558,N_15393);
and U15708 (N_15708,N_15214,N_15146);
nand U15709 (N_15709,N_15573,N_15232);
xor U15710 (N_15710,N_15135,N_15597);
nand U15711 (N_15711,N_15225,N_15121);
or U15712 (N_15712,N_15003,N_15353);
and U15713 (N_15713,N_15374,N_15089);
or U15714 (N_15714,N_15140,N_15342);
nor U15715 (N_15715,N_15445,N_15540);
nand U15716 (N_15716,N_15452,N_15518);
nor U15717 (N_15717,N_15218,N_15528);
or U15718 (N_15718,N_15243,N_15565);
xor U15719 (N_15719,N_15095,N_15291);
nand U15720 (N_15720,N_15238,N_15057);
or U15721 (N_15721,N_15460,N_15468);
nor U15722 (N_15722,N_15322,N_15124);
and U15723 (N_15723,N_15104,N_15509);
or U15724 (N_15724,N_15591,N_15568);
nor U15725 (N_15725,N_15317,N_15559);
xor U15726 (N_15726,N_15242,N_15466);
nor U15727 (N_15727,N_15163,N_15183);
or U15728 (N_15728,N_15566,N_15298);
nor U15729 (N_15729,N_15053,N_15073);
xor U15730 (N_15730,N_15272,N_15223);
or U15731 (N_15731,N_15453,N_15325);
and U15732 (N_15732,N_15338,N_15189);
or U15733 (N_15733,N_15376,N_15555);
xnor U15734 (N_15734,N_15207,N_15306);
xor U15735 (N_15735,N_15118,N_15480);
nand U15736 (N_15736,N_15455,N_15463);
xnor U15737 (N_15737,N_15324,N_15222);
xnor U15738 (N_15738,N_15182,N_15442);
nand U15739 (N_15739,N_15083,N_15138);
and U15740 (N_15740,N_15205,N_15287);
or U15741 (N_15741,N_15058,N_15341);
and U15742 (N_15742,N_15440,N_15332);
or U15743 (N_15743,N_15355,N_15279);
and U15744 (N_15744,N_15266,N_15250);
xor U15745 (N_15745,N_15367,N_15237);
or U15746 (N_15746,N_15383,N_15354);
nor U15747 (N_15747,N_15196,N_15219);
xnor U15748 (N_15748,N_15174,N_15056);
and U15749 (N_15749,N_15581,N_15529);
and U15750 (N_15750,N_15386,N_15190);
nor U15751 (N_15751,N_15599,N_15416);
and U15752 (N_15752,N_15179,N_15592);
and U15753 (N_15753,N_15268,N_15337);
or U15754 (N_15754,N_15409,N_15309);
or U15755 (N_15755,N_15570,N_15215);
xnor U15756 (N_15756,N_15404,N_15234);
or U15757 (N_15757,N_15173,N_15301);
xor U15758 (N_15758,N_15269,N_15062);
nor U15759 (N_15759,N_15399,N_15487);
nand U15760 (N_15760,N_15548,N_15061);
and U15761 (N_15761,N_15418,N_15420);
and U15762 (N_15762,N_15537,N_15458);
nor U15763 (N_15763,N_15048,N_15240);
nor U15764 (N_15764,N_15441,N_15501);
or U15765 (N_15765,N_15481,N_15586);
nand U15766 (N_15766,N_15246,N_15226);
or U15767 (N_15767,N_15267,N_15295);
or U15768 (N_15768,N_15274,N_15506);
or U15769 (N_15769,N_15143,N_15446);
and U15770 (N_15770,N_15072,N_15149);
or U15771 (N_15771,N_15172,N_15265);
nor U15772 (N_15772,N_15316,N_15497);
xor U15773 (N_15773,N_15220,N_15102);
nor U15774 (N_15774,N_15396,N_15554);
nor U15775 (N_15775,N_15181,N_15575);
nor U15776 (N_15776,N_15187,N_15033);
and U15777 (N_15777,N_15567,N_15006);
xnor U15778 (N_15778,N_15394,N_15106);
or U15779 (N_15779,N_15263,N_15539);
nand U15780 (N_15780,N_15283,N_15157);
xnor U15781 (N_15781,N_15105,N_15438);
and U15782 (N_15782,N_15159,N_15439);
nand U15783 (N_15783,N_15327,N_15208);
nand U15784 (N_15784,N_15136,N_15175);
xnor U15785 (N_15785,N_15071,N_15197);
or U15786 (N_15786,N_15177,N_15248);
xor U15787 (N_15787,N_15478,N_15133);
nand U15788 (N_15788,N_15447,N_15417);
or U15789 (N_15789,N_15031,N_15085);
and U15790 (N_15790,N_15473,N_15359);
and U15791 (N_15791,N_15027,N_15201);
nor U15792 (N_15792,N_15569,N_15176);
and U15793 (N_15793,N_15378,N_15155);
or U15794 (N_15794,N_15084,N_15241);
nor U15795 (N_15795,N_15524,N_15513);
or U15796 (N_15796,N_15093,N_15164);
and U15797 (N_15797,N_15526,N_15171);
or U15798 (N_15798,N_15039,N_15414);
nand U15799 (N_15799,N_15271,N_15329);
or U15800 (N_15800,N_15492,N_15549);
xnor U15801 (N_15801,N_15285,N_15191);
nor U15802 (N_15802,N_15395,N_15533);
or U15803 (N_15803,N_15531,N_15126);
xnor U15804 (N_15804,N_15350,N_15256);
or U15805 (N_15805,N_15412,N_15115);
or U15806 (N_15806,N_15461,N_15185);
nor U15807 (N_15807,N_15169,N_15002);
and U15808 (N_15808,N_15109,N_15107);
nor U15809 (N_15809,N_15264,N_15203);
nor U15810 (N_15810,N_15230,N_15362);
xor U15811 (N_15811,N_15258,N_15541);
and U15812 (N_15812,N_15040,N_15499);
and U15813 (N_15813,N_15275,N_15562);
nor U15814 (N_15814,N_15556,N_15474);
xnor U15815 (N_15815,N_15023,N_15488);
nor U15816 (N_15816,N_15116,N_15000);
xnor U15817 (N_15817,N_15029,N_15398);
and U15818 (N_15818,N_15103,N_15119);
nand U15819 (N_15819,N_15064,N_15339);
and U15820 (N_15820,N_15047,N_15251);
nand U15821 (N_15821,N_15129,N_15522);
nor U15822 (N_15822,N_15482,N_15491);
or U15823 (N_15823,N_15530,N_15498);
nand U15824 (N_15824,N_15411,N_15013);
xor U15825 (N_15825,N_15546,N_15380);
and U15826 (N_15826,N_15070,N_15016);
and U15827 (N_15827,N_15390,N_15307);
nand U15828 (N_15828,N_15130,N_15167);
xnor U15829 (N_15829,N_15577,N_15382);
nor U15830 (N_15830,N_15007,N_15144);
or U15831 (N_15831,N_15098,N_15079);
or U15832 (N_15832,N_15576,N_15389);
nor U15833 (N_15833,N_15422,N_15131);
nand U15834 (N_15834,N_15360,N_15333);
or U15835 (N_15835,N_15276,N_15166);
and U15836 (N_15836,N_15305,N_15108);
nor U15837 (N_15837,N_15054,N_15477);
xor U15838 (N_15838,N_15472,N_15142);
nor U15839 (N_15839,N_15563,N_15510);
xnor U15840 (N_15840,N_15508,N_15430);
nand U15841 (N_15841,N_15132,N_15361);
nor U15842 (N_15842,N_15517,N_15296);
or U15843 (N_15843,N_15500,N_15245);
or U15844 (N_15844,N_15037,N_15593);
xor U15845 (N_15845,N_15479,N_15314);
and U15846 (N_15846,N_15469,N_15262);
nor U15847 (N_15847,N_15277,N_15292);
nor U15848 (N_15848,N_15406,N_15335);
nor U15849 (N_15849,N_15151,N_15017);
or U15850 (N_15850,N_15158,N_15113);
nor U15851 (N_15851,N_15485,N_15014);
xnor U15852 (N_15852,N_15216,N_15346);
and U15853 (N_15853,N_15125,N_15547);
xor U15854 (N_15854,N_15236,N_15259);
nand U15855 (N_15855,N_15302,N_15370);
xor U15856 (N_15856,N_15319,N_15290);
xor U15857 (N_15857,N_15297,N_15094);
or U15858 (N_15858,N_15456,N_15336);
or U15859 (N_15859,N_15112,N_15209);
and U15860 (N_15860,N_15391,N_15340);
xor U15861 (N_15861,N_15111,N_15231);
nand U15862 (N_15862,N_15282,N_15433);
xor U15863 (N_15863,N_15429,N_15097);
and U15864 (N_15864,N_15344,N_15450);
nand U15865 (N_15865,N_15046,N_15110);
and U15866 (N_15866,N_15459,N_15233);
or U15867 (N_15867,N_15589,N_15065);
and U15868 (N_15868,N_15020,N_15086);
and U15869 (N_15869,N_15066,N_15511);
and U15870 (N_15870,N_15284,N_15579);
nor U15871 (N_15871,N_15150,N_15351);
and U15872 (N_15872,N_15571,N_15034);
nand U15873 (N_15873,N_15534,N_15200);
nor U15874 (N_15874,N_15403,N_15369);
xnor U15875 (N_15875,N_15160,N_15454);
or U15876 (N_15876,N_15594,N_15432);
or U15877 (N_15877,N_15045,N_15289);
nor U15878 (N_15878,N_15431,N_15596);
nor U15879 (N_15879,N_15165,N_15075);
and U15880 (N_15880,N_15035,N_15519);
or U15881 (N_15881,N_15387,N_15320);
or U15882 (N_15882,N_15448,N_15331);
nor U15883 (N_15883,N_15516,N_15059);
xnor U15884 (N_15884,N_15578,N_15490);
xnor U15885 (N_15885,N_15049,N_15114);
xnor U15886 (N_15886,N_15352,N_15381);
and U15887 (N_15887,N_15212,N_15227);
nand U15888 (N_15888,N_15428,N_15022);
and U15889 (N_15889,N_15330,N_15019);
nand U15890 (N_15890,N_15574,N_15527);
xor U15891 (N_15891,N_15092,N_15371);
xnor U15892 (N_15892,N_15312,N_15402);
nand U15893 (N_15893,N_15410,N_15253);
nor U15894 (N_15894,N_15148,N_15443);
xnor U15895 (N_15895,N_15123,N_15318);
and U15896 (N_15896,N_15543,N_15384);
or U15897 (N_15897,N_15315,N_15210);
nand U15898 (N_15898,N_15063,N_15415);
nor U15899 (N_15899,N_15141,N_15521);
or U15900 (N_15900,N_15119,N_15568);
nor U15901 (N_15901,N_15248,N_15368);
xnor U15902 (N_15902,N_15470,N_15589);
nor U15903 (N_15903,N_15399,N_15206);
xnor U15904 (N_15904,N_15299,N_15413);
nand U15905 (N_15905,N_15561,N_15135);
nand U15906 (N_15906,N_15461,N_15318);
xor U15907 (N_15907,N_15439,N_15381);
xnor U15908 (N_15908,N_15487,N_15531);
nand U15909 (N_15909,N_15279,N_15565);
and U15910 (N_15910,N_15248,N_15323);
and U15911 (N_15911,N_15347,N_15257);
or U15912 (N_15912,N_15402,N_15058);
nand U15913 (N_15913,N_15328,N_15054);
xor U15914 (N_15914,N_15003,N_15263);
and U15915 (N_15915,N_15452,N_15224);
or U15916 (N_15916,N_15509,N_15417);
nor U15917 (N_15917,N_15136,N_15370);
nand U15918 (N_15918,N_15153,N_15359);
or U15919 (N_15919,N_15316,N_15371);
and U15920 (N_15920,N_15240,N_15258);
xor U15921 (N_15921,N_15512,N_15558);
nand U15922 (N_15922,N_15597,N_15569);
xor U15923 (N_15923,N_15445,N_15077);
nand U15924 (N_15924,N_15266,N_15354);
nor U15925 (N_15925,N_15009,N_15598);
nor U15926 (N_15926,N_15424,N_15157);
nor U15927 (N_15927,N_15309,N_15149);
nor U15928 (N_15928,N_15093,N_15075);
nor U15929 (N_15929,N_15536,N_15263);
nor U15930 (N_15930,N_15194,N_15308);
nor U15931 (N_15931,N_15045,N_15278);
nand U15932 (N_15932,N_15499,N_15354);
nand U15933 (N_15933,N_15517,N_15201);
nor U15934 (N_15934,N_15353,N_15568);
xnor U15935 (N_15935,N_15381,N_15263);
xnor U15936 (N_15936,N_15459,N_15311);
nor U15937 (N_15937,N_15088,N_15082);
nor U15938 (N_15938,N_15275,N_15288);
xnor U15939 (N_15939,N_15002,N_15103);
or U15940 (N_15940,N_15247,N_15588);
or U15941 (N_15941,N_15517,N_15306);
xor U15942 (N_15942,N_15454,N_15220);
nor U15943 (N_15943,N_15379,N_15340);
nor U15944 (N_15944,N_15513,N_15581);
nand U15945 (N_15945,N_15226,N_15332);
nand U15946 (N_15946,N_15584,N_15160);
nand U15947 (N_15947,N_15141,N_15221);
nor U15948 (N_15948,N_15388,N_15210);
or U15949 (N_15949,N_15158,N_15565);
nand U15950 (N_15950,N_15312,N_15410);
xnor U15951 (N_15951,N_15385,N_15255);
or U15952 (N_15952,N_15290,N_15360);
nand U15953 (N_15953,N_15413,N_15369);
nor U15954 (N_15954,N_15453,N_15002);
nand U15955 (N_15955,N_15010,N_15185);
xor U15956 (N_15956,N_15548,N_15202);
or U15957 (N_15957,N_15461,N_15383);
nand U15958 (N_15958,N_15006,N_15370);
or U15959 (N_15959,N_15268,N_15328);
xor U15960 (N_15960,N_15490,N_15010);
nor U15961 (N_15961,N_15432,N_15344);
nor U15962 (N_15962,N_15470,N_15017);
xnor U15963 (N_15963,N_15136,N_15358);
and U15964 (N_15964,N_15286,N_15400);
and U15965 (N_15965,N_15261,N_15496);
xor U15966 (N_15966,N_15192,N_15538);
xnor U15967 (N_15967,N_15276,N_15125);
or U15968 (N_15968,N_15539,N_15407);
or U15969 (N_15969,N_15292,N_15031);
xor U15970 (N_15970,N_15319,N_15082);
and U15971 (N_15971,N_15082,N_15413);
or U15972 (N_15972,N_15552,N_15276);
nor U15973 (N_15973,N_15580,N_15108);
or U15974 (N_15974,N_15159,N_15371);
or U15975 (N_15975,N_15162,N_15496);
and U15976 (N_15976,N_15477,N_15363);
and U15977 (N_15977,N_15402,N_15568);
and U15978 (N_15978,N_15066,N_15515);
xor U15979 (N_15979,N_15214,N_15525);
and U15980 (N_15980,N_15566,N_15156);
and U15981 (N_15981,N_15106,N_15436);
and U15982 (N_15982,N_15326,N_15038);
nor U15983 (N_15983,N_15251,N_15550);
and U15984 (N_15984,N_15402,N_15080);
and U15985 (N_15985,N_15151,N_15536);
xor U15986 (N_15986,N_15400,N_15506);
nor U15987 (N_15987,N_15148,N_15540);
nand U15988 (N_15988,N_15536,N_15211);
nand U15989 (N_15989,N_15211,N_15545);
or U15990 (N_15990,N_15565,N_15584);
or U15991 (N_15991,N_15508,N_15493);
nand U15992 (N_15992,N_15112,N_15045);
xnor U15993 (N_15993,N_15176,N_15417);
xnor U15994 (N_15994,N_15361,N_15329);
xor U15995 (N_15995,N_15479,N_15148);
xor U15996 (N_15996,N_15325,N_15527);
and U15997 (N_15997,N_15416,N_15157);
nor U15998 (N_15998,N_15274,N_15332);
and U15999 (N_15999,N_15544,N_15281);
or U16000 (N_16000,N_15199,N_15452);
and U16001 (N_16001,N_15235,N_15445);
nand U16002 (N_16002,N_15289,N_15567);
nor U16003 (N_16003,N_15352,N_15123);
xor U16004 (N_16004,N_15204,N_15215);
or U16005 (N_16005,N_15098,N_15131);
nand U16006 (N_16006,N_15134,N_15143);
nand U16007 (N_16007,N_15502,N_15411);
nor U16008 (N_16008,N_15061,N_15328);
nor U16009 (N_16009,N_15007,N_15062);
or U16010 (N_16010,N_15228,N_15073);
nand U16011 (N_16011,N_15521,N_15286);
or U16012 (N_16012,N_15021,N_15178);
nor U16013 (N_16013,N_15297,N_15405);
nor U16014 (N_16014,N_15427,N_15405);
xor U16015 (N_16015,N_15470,N_15366);
nand U16016 (N_16016,N_15263,N_15574);
and U16017 (N_16017,N_15368,N_15140);
or U16018 (N_16018,N_15533,N_15317);
nand U16019 (N_16019,N_15044,N_15419);
or U16020 (N_16020,N_15257,N_15340);
nand U16021 (N_16021,N_15343,N_15128);
or U16022 (N_16022,N_15412,N_15108);
and U16023 (N_16023,N_15402,N_15041);
nand U16024 (N_16024,N_15405,N_15327);
nor U16025 (N_16025,N_15046,N_15038);
nand U16026 (N_16026,N_15416,N_15577);
or U16027 (N_16027,N_15374,N_15048);
nor U16028 (N_16028,N_15210,N_15466);
and U16029 (N_16029,N_15584,N_15367);
xor U16030 (N_16030,N_15396,N_15155);
nand U16031 (N_16031,N_15570,N_15164);
nor U16032 (N_16032,N_15480,N_15425);
and U16033 (N_16033,N_15182,N_15009);
xnor U16034 (N_16034,N_15325,N_15539);
or U16035 (N_16035,N_15225,N_15367);
nand U16036 (N_16036,N_15524,N_15199);
xnor U16037 (N_16037,N_15430,N_15290);
xnor U16038 (N_16038,N_15015,N_15581);
and U16039 (N_16039,N_15505,N_15525);
xor U16040 (N_16040,N_15592,N_15129);
nand U16041 (N_16041,N_15220,N_15342);
xnor U16042 (N_16042,N_15425,N_15491);
xor U16043 (N_16043,N_15596,N_15440);
and U16044 (N_16044,N_15392,N_15244);
or U16045 (N_16045,N_15477,N_15046);
nor U16046 (N_16046,N_15424,N_15016);
nor U16047 (N_16047,N_15049,N_15336);
nand U16048 (N_16048,N_15413,N_15158);
nor U16049 (N_16049,N_15597,N_15582);
nand U16050 (N_16050,N_15174,N_15159);
nand U16051 (N_16051,N_15075,N_15103);
nor U16052 (N_16052,N_15390,N_15049);
xor U16053 (N_16053,N_15150,N_15125);
xor U16054 (N_16054,N_15272,N_15241);
nand U16055 (N_16055,N_15426,N_15065);
nor U16056 (N_16056,N_15313,N_15330);
or U16057 (N_16057,N_15296,N_15399);
or U16058 (N_16058,N_15439,N_15171);
or U16059 (N_16059,N_15371,N_15023);
and U16060 (N_16060,N_15537,N_15334);
or U16061 (N_16061,N_15021,N_15468);
nand U16062 (N_16062,N_15151,N_15399);
nand U16063 (N_16063,N_15036,N_15511);
or U16064 (N_16064,N_15439,N_15183);
xor U16065 (N_16065,N_15033,N_15412);
nand U16066 (N_16066,N_15021,N_15299);
nor U16067 (N_16067,N_15485,N_15045);
and U16068 (N_16068,N_15566,N_15476);
nand U16069 (N_16069,N_15205,N_15494);
or U16070 (N_16070,N_15459,N_15283);
or U16071 (N_16071,N_15445,N_15495);
xnor U16072 (N_16072,N_15038,N_15305);
xor U16073 (N_16073,N_15049,N_15414);
and U16074 (N_16074,N_15137,N_15249);
xnor U16075 (N_16075,N_15141,N_15212);
nor U16076 (N_16076,N_15079,N_15554);
nand U16077 (N_16077,N_15042,N_15545);
or U16078 (N_16078,N_15395,N_15531);
and U16079 (N_16079,N_15327,N_15129);
nor U16080 (N_16080,N_15079,N_15006);
xnor U16081 (N_16081,N_15217,N_15491);
or U16082 (N_16082,N_15348,N_15472);
or U16083 (N_16083,N_15164,N_15050);
xor U16084 (N_16084,N_15051,N_15512);
nand U16085 (N_16085,N_15199,N_15217);
and U16086 (N_16086,N_15010,N_15256);
or U16087 (N_16087,N_15015,N_15018);
nand U16088 (N_16088,N_15248,N_15277);
xor U16089 (N_16089,N_15157,N_15474);
nor U16090 (N_16090,N_15369,N_15000);
nand U16091 (N_16091,N_15360,N_15209);
nor U16092 (N_16092,N_15484,N_15241);
nor U16093 (N_16093,N_15177,N_15339);
xnor U16094 (N_16094,N_15269,N_15245);
or U16095 (N_16095,N_15325,N_15542);
xnor U16096 (N_16096,N_15308,N_15462);
nor U16097 (N_16097,N_15395,N_15150);
nand U16098 (N_16098,N_15334,N_15042);
and U16099 (N_16099,N_15514,N_15436);
or U16100 (N_16100,N_15466,N_15181);
and U16101 (N_16101,N_15523,N_15365);
nand U16102 (N_16102,N_15485,N_15037);
xor U16103 (N_16103,N_15128,N_15361);
and U16104 (N_16104,N_15044,N_15224);
nand U16105 (N_16105,N_15004,N_15552);
nor U16106 (N_16106,N_15576,N_15271);
and U16107 (N_16107,N_15383,N_15183);
xor U16108 (N_16108,N_15001,N_15584);
or U16109 (N_16109,N_15522,N_15432);
xor U16110 (N_16110,N_15365,N_15250);
and U16111 (N_16111,N_15037,N_15587);
xnor U16112 (N_16112,N_15347,N_15381);
nand U16113 (N_16113,N_15118,N_15244);
and U16114 (N_16114,N_15123,N_15592);
xnor U16115 (N_16115,N_15410,N_15588);
nand U16116 (N_16116,N_15341,N_15106);
and U16117 (N_16117,N_15218,N_15381);
nand U16118 (N_16118,N_15453,N_15590);
and U16119 (N_16119,N_15201,N_15442);
xnor U16120 (N_16120,N_15206,N_15496);
nand U16121 (N_16121,N_15089,N_15108);
or U16122 (N_16122,N_15393,N_15459);
and U16123 (N_16123,N_15051,N_15460);
nor U16124 (N_16124,N_15290,N_15231);
nand U16125 (N_16125,N_15463,N_15568);
or U16126 (N_16126,N_15179,N_15322);
nand U16127 (N_16127,N_15442,N_15033);
or U16128 (N_16128,N_15240,N_15213);
nor U16129 (N_16129,N_15235,N_15326);
xor U16130 (N_16130,N_15073,N_15462);
nor U16131 (N_16131,N_15266,N_15191);
or U16132 (N_16132,N_15521,N_15419);
and U16133 (N_16133,N_15370,N_15221);
and U16134 (N_16134,N_15401,N_15533);
nand U16135 (N_16135,N_15311,N_15533);
nand U16136 (N_16136,N_15128,N_15565);
and U16137 (N_16137,N_15086,N_15128);
xnor U16138 (N_16138,N_15079,N_15154);
and U16139 (N_16139,N_15220,N_15133);
or U16140 (N_16140,N_15016,N_15298);
or U16141 (N_16141,N_15091,N_15320);
or U16142 (N_16142,N_15520,N_15387);
nor U16143 (N_16143,N_15408,N_15442);
and U16144 (N_16144,N_15118,N_15092);
and U16145 (N_16145,N_15408,N_15050);
xor U16146 (N_16146,N_15253,N_15323);
or U16147 (N_16147,N_15144,N_15356);
and U16148 (N_16148,N_15092,N_15511);
nor U16149 (N_16149,N_15581,N_15251);
or U16150 (N_16150,N_15221,N_15272);
xor U16151 (N_16151,N_15162,N_15423);
nand U16152 (N_16152,N_15286,N_15402);
or U16153 (N_16153,N_15215,N_15069);
xnor U16154 (N_16154,N_15281,N_15188);
xnor U16155 (N_16155,N_15446,N_15512);
nor U16156 (N_16156,N_15366,N_15555);
or U16157 (N_16157,N_15220,N_15432);
or U16158 (N_16158,N_15099,N_15079);
nand U16159 (N_16159,N_15076,N_15352);
nand U16160 (N_16160,N_15499,N_15015);
nor U16161 (N_16161,N_15251,N_15166);
or U16162 (N_16162,N_15097,N_15422);
nand U16163 (N_16163,N_15352,N_15264);
nand U16164 (N_16164,N_15238,N_15345);
and U16165 (N_16165,N_15521,N_15575);
nand U16166 (N_16166,N_15201,N_15482);
nand U16167 (N_16167,N_15314,N_15457);
or U16168 (N_16168,N_15453,N_15579);
nor U16169 (N_16169,N_15087,N_15288);
or U16170 (N_16170,N_15125,N_15550);
nand U16171 (N_16171,N_15074,N_15377);
nand U16172 (N_16172,N_15472,N_15478);
nand U16173 (N_16173,N_15250,N_15029);
or U16174 (N_16174,N_15435,N_15278);
or U16175 (N_16175,N_15346,N_15100);
nor U16176 (N_16176,N_15441,N_15017);
nor U16177 (N_16177,N_15517,N_15334);
xor U16178 (N_16178,N_15154,N_15273);
and U16179 (N_16179,N_15597,N_15415);
nand U16180 (N_16180,N_15240,N_15403);
nand U16181 (N_16181,N_15247,N_15325);
and U16182 (N_16182,N_15113,N_15263);
or U16183 (N_16183,N_15574,N_15174);
xnor U16184 (N_16184,N_15273,N_15459);
or U16185 (N_16185,N_15483,N_15348);
nor U16186 (N_16186,N_15062,N_15023);
nand U16187 (N_16187,N_15198,N_15328);
or U16188 (N_16188,N_15016,N_15304);
and U16189 (N_16189,N_15430,N_15240);
nand U16190 (N_16190,N_15540,N_15322);
or U16191 (N_16191,N_15502,N_15074);
and U16192 (N_16192,N_15378,N_15594);
xnor U16193 (N_16193,N_15161,N_15552);
or U16194 (N_16194,N_15477,N_15059);
nor U16195 (N_16195,N_15425,N_15018);
and U16196 (N_16196,N_15166,N_15456);
and U16197 (N_16197,N_15268,N_15013);
and U16198 (N_16198,N_15167,N_15341);
and U16199 (N_16199,N_15584,N_15550);
nand U16200 (N_16200,N_16127,N_15956);
nand U16201 (N_16201,N_15680,N_15681);
or U16202 (N_16202,N_15961,N_15846);
and U16203 (N_16203,N_15606,N_15993);
xnor U16204 (N_16204,N_16069,N_15906);
nor U16205 (N_16205,N_15851,N_15827);
or U16206 (N_16206,N_15860,N_16123);
xor U16207 (N_16207,N_15636,N_15826);
nand U16208 (N_16208,N_15809,N_15647);
nand U16209 (N_16209,N_15706,N_15669);
xor U16210 (N_16210,N_16095,N_16191);
nor U16211 (N_16211,N_16176,N_15867);
or U16212 (N_16212,N_16067,N_15743);
nor U16213 (N_16213,N_15836,N_15666);
nor U16214 (N_16214,N_15810,N_16077);
and U16215 (N_16215,N_15639,N_16143);
nor U16216 (N_16216,N_15813,N_15767);
xnor U16217 (N_16217,N_16179,N_16039);
or U16218 (N_16218,N_15741,N_15861);
nor U16219 (N_16219,N_15764,N_16013);
or U16220 (N_16220,N_15896,N_16126);
nand U16221 (N_16221,N_15736,N_16119);
and U16222 (N_16222,N_16007,N_16034);
or U16223 (N_16223,N_16004,N_15963);
or U16224 (N_16224,N_15693,N_15845);
nor U16225 (N_16225,N_15638,N_15910);
nor U16226 (N_16226,N_15912,N_15942);
nand U16227 (N_16227,N_15795,N_16121);
or U16228 (N_16228,N_16137,N_15624);
xnor U16229 (N_16229,N_15721,N_15978);
xnor U16230 (N_16230,N_15878,N_15713);
and U16231 (N_16231,N_15691,N_16112);
and U16232 (N_16232,N_16037,N_15717);
and U16233 (N_16233,N_16110,N_15848);
and U16234 (N_16234,N_16064,N_15923);
and U16235 (N_16235,N_16146,N_15864);
xnor U16236 (N_16236,N_15931,N_16080);
xor U16237 (N_16237,N_15899,N_16173);
nor U16238 (N_16238,N_15665,N_16133);
xor U16239 (N_16239,N_15729,N_15857);
or U16240 (N_16240,N_15779,N_16047);
nand U16241 (N_16241,N_15742,N_15966);
xnor U16242 (N_16242,N_15811,N_16085);
xnor U16243 (N_16243,N_15799,N_15840);
and U16244 (N_16244,N_16149,N_16076);
nand U16245 (N_16245,N_15780,N_15756);
xnor U16246 (N_16246,N_15866,N_15828);
nor U16247 (N_16247,N_16038,N_15890);
nor U16248 (N_16248,N_15996,N_15618);
or U16249 (N_16249,N_15698,N_16180);
nor U16250 (N_16250,N_15654,N_16078);
or U16251 (N_16251,N_16114,N_15824);
xnor U16252 (N_16252,N_15869,N_16008);
nand U16253 (N_16253,N_15925,N_16079);
and U16254 (N_16254,N_16159,N_16056);
xor U16255 (N_16255,N_16059,N_15834);
xor U16256 (N_16256,N_15648,N_15633);
nor U16257 (N_16257,N_15823,N_15985);
xor U16258 (N_16258,N_15871,N_15865);
or U16259 (N_16259,N_16071,N_15999);
nor U16260 (N_16260,N_16144,N_15979);
and U16261 (N_16261,N_15762,N_15850);
and U16262 (N_16262,N_16031,N_16048);
xnor U16263 (N_16263,N_16167,N_15621);
and U16264 (N_16264,N_15971,N_16141);
or U16265 (N_16265,N_16044,N_15752);
or U16266 (N_16266,N_16014,N_15883);
nor U16267 (N_16267,N_15619,N_15808);
xor U16268 (N_16268,N_16186,N_15992);
and U16269 (N_16269,N_16171,N_15874);
xnor U16270 (N_16270,N_16193,N_15806);
and U16271 (N_16271,N_15714,N_16073);
or U16272 (N_16272,N_16160,N_16156);
or U16273 (N_16273,N_16166,N_15941);
xnor U16274 (N_16274,N_15632,N_16061);
nand U16275 (N_16275,N_15642,N_15924);
and U16276 (N_16276,N_15653,N_15807);
xor U16277 (N_16277,N_15952,N_16089);
nor U16278 (N_16278,N_16084,N_15674);
and U16279 (N_16279,N_15786,N_15991);
nand U16280 (N_16280,N_15782,N_15684);
xor U16281 (N_16281,N_15841,N_15877);
nand U16282 (N_16282,N_16118,N_15640);
or U16283 (N_16283,N_16020,N_15699);
and U16284 (N_16284,N_16041,N_15613);
and U16285 (N_16285,N_15897,N_15607);
nor U16286 (N_16286,N_15611,N_15948);
nor U16287 (N_16287,N_15600,N_16097);
xor U16288 (N_16288,N_16099,N_15820);
nand U16289 (N_16289,N_16122,N_16115);
xor U16290 (N_16290,N_15749,N_15888);
and U16291 (N_16291,N_16055,N_15730);
or U16292 (N_16292,N_15967,N_16053);
nand U16293 (N_16293,N_16125,N_15614);
or U16294 (N_16294,N_15715,N_16030);
and U16295 (N_16295,N_15880,N_15670);
xnor U16296 (N_16296,N_16036,N_15928);
and U16297 (N_16297,N_15946,N_16090);
nand U16298 (N_16298,N_15609,N_16103);
and U16299 (N_16299,N_15832,N_15711);
xnor U16300 (N_16300,N_15605,N_15821);
nor U16301 (N_16301,N_15602,N_16196);
xnor U16302 (N_16302,N_15801,N_15745);
nand U16303 (N_16303,N_16132,N_15672);
nand U16304 (N_16304,N_16063,N_15601);
or U16305 (N_16305,N_15989,N_16134);
xor U16306 (N_16306,N_15737,N_15889);
nand U16307 (N_16307,N_16065,N_15709);
xnor U16308 (N_16308,N_15696,N_15676);
or U16309 (N_16309,N_16022,N_15853);
xnor U16310 (N_16310,N_15833,N_15785);
xnor U16311 (N_16311,N_15759,N_15944);
and U16312 (N_16312,N_16109,N_15689);
nor U16313 (N_16313,N_16023,N_16100);
nor U16314 (N_16314,N_16182,N_15969);
or U16315 (N_16315,N_15917,N_16172);
nor U16316 (N_16316,N_15740,N_16162);
and U16317 (N_16317,N_15754,N_15976);
and U16318 (N_16318,N_15987,N_16165);
nand U16319 (N_16319,N_15977,N_15915);
nor U16320 (N_16320,N_15658,N_15814);
or U16321 (N_16321,N_15708,N_16113);
or U16322 (N_16322,N_15849,N_15817);
and U16323 (N_16323,N_15997,N_15794);
or U16324 (N_16324,N_15879,N_15943);
nor U16325 (N_16325,N_16108,N_15616);
and U16326 (N_16326,N_15651,N_16151);
xnor U16327 (N_16327,N_15755,N_16001);
nor U16328 (N_16328,N_16129,N_16012);
nand U16329 (N_16329,N_15988,N_16117);
and U16330 (N_16330,N_15898,N_15704);
or U16331 (N_16331,N_15758,N_15733);
nand U16332 (N_16332,N_16083,N_15913);
nand U16333 (N_16333,N_16046,N_16028);
or U16334 (N_16334,N_16091,N_15789);
xnor U16335 (N_16335,N_15875,N_16060);
and U16336 (N_16336,N_15830,N_15995);
nand U16337 (N_16337,N_16111,N_16152);
nand U16338 (N_16338,N_16018,N_15902);
nor U16339 (N_16339,N_15784,N_16153);
and U16340 (N_16340,N_15936,N_15885);
xnor U16341 (N_16341,N_15778,N_15723);
nand U16342 (N_16342,N_15679,N_15986);
or U16343 (N_16343,N_16106,N_16158);
nand U16344 (N_16344,N_15703,N_15661);
nand U16345 (N_16345,N_15858,N_15934);
xnor U16346 (N_16346,N_15949,N_16058);
and U16347 (N_16347,N_15712,N_16101);
and U16348 (N_16348,N_16006,N_15731);
and U16349 (N_16349,N_15710,N_15635);
xnor U16350 (N_16350,N_16124,N_15629);
nor U16351 (N_16351,N_15907,N_16054);
or U16352 (N_16352,N_16197,N_16198);
and U16353 (N_16353,N_16016,N_16187);
xnor U16354 (N_16354,N_15604,N_15751);
and U16355 (N_16355,N_16145,N_16000);
or U16356 (N_16356,N_15735,N_15694);
or U16357 (N_16357,N_16026,N_16189);
and U16358 (N_16358,N_16181,N_15677);
and U16359 (N_16359,N_15678,N_15726);
nor U16360 (N_16360,N_15825,N_16105);
xnor U16361 (N_16361,N_15938,N_15771);
nand U16362 (N_16362,N_15775,N_15972);
or U16363 (N_16363,N_15870,N_15620);
or U16364 (N_16364,N_15937,N_15700);
and U16365 (N_16365,N_15660,N_15932);
or U16366 (N_16366,N_15748,N_16025);
nor U16367 (N_16367,N_16051,N_15671);
nand U16368 (N_16368,N_15626,N_15905);
nand U16369 (N_16369,N_15984,N_16042);
nand U16370 (N_16370,N_16147,N_15650);
nand U16371 (N_16371,N_15831,N_15904);
and U16372 (N_16372,N_15772,N_15753);
or U16373 (N_16373,N_15746,N_15876);
xnor U16374 (N_16374,N_16011,N_15707);
nor U16375 (N_16375,N_16081,N_15697);
nand U16376 (N_16376,N_15757,N_16195);
or U16377 (N_16377,N_15854,N_15882);
nor U16378 (N_16378,N_16005,N_16170);
or U16379 (N_16379,N_16094,N_15615);
xnor U16380 (N_16380,N_15732,N_16074);
xnor U16381 (N_16381,N_16049,N_15921);
nor U16382 (N_16382,N_15982,N_16154);
nand U16383 (N_16383,N_15628,N_16168);
nand U16384 (N_16384,N_15900,N_16032);
or U16385 (N_16385,N_16174,N_16027);
and U16386 (N_16386,N_16043,N_15927);
nand U16387 (N_16387,N_15998,N_16130);
nor U16388 (N_16388,N_16092,N_15655);
nor U16389 (N_16389,N_15617,N_15873);
or U16390 (N_16390,N_15686,N_15862);
and U16391 (N_16391,N_15829,N_15702);
nand U16392 (N_16392,N_16093,N_15692);
xnor U16393 (N_16393,N_15816,N_15603);
and U16394 (N_16394,N_16184,N_15662);
and U16395 (N_16395,N_15657,N_15947);
xor U16396 (N_16396,N_16072,N_15940);
or U16397 (N_16397,N_15856,N_15776);
or U16398 (N_16398,N_15981,N_15815);
and U16399 (N_16399,N_16157,N_16029);
xnor U16400 (N_16400,N_15783,N_15768);
nand U16401 (N_16401,N_16135,N_15770);
or U16402 (N_16402,N_15951,N_15855);
or U16403 (N_16403,N_15769,N_16033);
xor U16404 (N_16404,N_16150,N_15818);
or U16405 (N_16405,N_16070,N_16024);
xor U16406 (N_16406,N_15791,N_15634);
nor U16407 (N_16407,N_15796,N_15962);
nor U16408 (N_16408,N_15909,N_15787);
and U16409 (N_16409,N_15922,N_16136);
xnor U16410 (N_16410,N_15652,N_16188);
xnor U16411 (N_16411,N_16102,N_15950);
nor U16412 (N_16412,N_15687,N_15911);
and U16413 (N_16413,N_15837,N_15610);
or U16414 (N_16414,N_15903,N_15819);
nor U16415 (N_16415,N_15872,N_15920);
nor U16416 (N_16416,N_15935,N_16086);
and U16417 (N_16417,N_15690,N_15724);
nand U16418 (N_16418,N_16104,N_16155);
and U16419 (N_16419,N_15804,N_15964);
nand U16420 (N_16420,N_15627,N_15887);
nand U16421 (N_16421,N_15983,N_15631);
or U16422 (N_16422,N_15608,N_15918);
nor U16423 (N_16423,N_16185,N_15641);
xor U16424 (N_16424,N_15894,N_15645);
and U16425 (N_16425,N_15649,N_15750);
nand U16426 (N_16426,N_16003,N_15926);
and U16427 (N_16427,N_15719,N_15908);
xnor U16428 (N_16428,N_15667,N_15842);
nor U16429 (N_16429,N_16139,N_15763);
xor U16430 (N_16430,N_15695,N_16057);
xor U16431 (N_16431,N_15975,N_16098);
and U16432 (N_16432,N_15727,N_15930);
and U16433 (N_16433,N_15958,N_15761);
nand U16434 (N_16434,N_15725,N_16175);
xor U16435 (N_16435,N_15622,N_15675);
and U16436 (N_16436,N_15974,N_15844);
nand U16437 (N_16437,N_15863,N_16192);
nand U16438 (N_16438,N_15859,N_16035);
xnor U16439 (N_16439,N_15980,N_15797);
xor U16440 (N_16440,N_15893,N_16140);
nor U16441 (N_16441,N_15822,N_15777);
or U16442 (N_16442,N_15744,N_15973);
nor U16443 (N_16443,N_15747,N_15919);
and U16444 (N_16444,N_15843,N_16131);
or U16445 (N_16445,N_15728,N_16120);
and U16446 (N_16446,N_15929,N_15664);
nor U16447 (N_16447,N_15773,N_16010);
nor U16448 (N_16448,N_15722,N_16088);
and U16449 (N_16449,N_15960,N_16052);
or U16450 (N_16450,N_15805,N_15895);
nand U16451 (N_16451,N_15734,N_15933);
and U16452 (N_16452,N_16015,N_16082);
nor U16453 (N_16453,N_15838,N_15790);
or U16454 (N_16454,N_15612,N_16190);
nor U16455 (N_16455,N_15798,N_15701);
nand U16456 (N_16456,N_15623,N_15803);
or U16457 (N_16457,N_16138,N_15891);
or U16458 (N_16458,N_15955,N_15868);
or U16459 (N_16459,N_15774,N_15673);
or U16460 (N_16460,N_16148,N_16164);
or U16461 (N_16461,N_16021,N_15884);
nand U16462 (N_16462,N_15901,N_15800);
or U16463 (N_16463,N_15886,N_15739);
nor U16464 (N_16464,N_15760,N_16169);
and U16465 (N_16465,N_15852,N_15953);
xor U16466 (N_16466,N_15847,N_16075);
and U16467 (N_16467,N_15637,N_15765);
nand U16468 (N_16468,N_16183,N_15625);
nand U16469 (N_16469,N_15683,N_15688);
nand U16470 (N_16470,N_15792,N_15685);
or U16471 (N_16471,N_16068,N_15990);
or U16472 (N_16472,N_15957,N_15766);
nand U16473 (N_16473,N_15881,N_15802);
xnor U16474 (N_16474,N_15656,N_16161);
or U16475 (N_16475,N_16045,N_15643);
xor U16476 (N_16476,N_15965,N_16019);
and U16477 (N_16477,N_15720,N_16009);
nand U16478 (N_16478,N_15781,N_16116);
xnor U16479 (N_16479,N_16017,N_16177);
or U16480 (N_16480,N_16142,N_15644);
and U16481 (N_16481,N_15916,N_16040);
or U16482 (N_16482,N_15682,N_15663);
xor U16483 (N_16483,N_15994,N_16107);
nand U16484 (N_16484,N_15705,N_16062);
nor U16485 (N_16485,N_15716,N_16002);
xor U16486 (N_16486,N_16087,N_15954);
nand U16487 (N_16487,N_15630,N_15793);
nor U16488 (N_16488,N_15668,N_15892);
nor U16489 (N_16489,N_16128,N_15914);
nand U16490 (N_16490,N_15812,N_15839);
nor U16491 (N_16491,N_16050,N_15968);
and U16492 (N_16492,N_15718,N_15738);
nand U16493 (N_16493,N_16066,N_16163);
nand U16494 (N_16494,N_16194,N_15646);
or U16495 (N_16495,N_16178,N_15959);
nand U16496 (N_16496,N_15788,N_15945);
or U16497 (N_16497,N_16096,N_16199);
or U16498 (N_16498,N_15659,N_15835);
and U16499 (N_16499,N_15970,N_15939);
nor U16500 (N_16500,N_15929,N_16113);
and U16501 (N_16501,N_15905,N_15632);
xor U16502 (N_16502,N_15946,N_15745);
and U16503 (N_16503,N_15927,N_16053);
or U16504 (N_16504,N_15965,N_15782);
nor U16505 (N_16505,N_15724,N_15973);
and U16506 (N_16506,N_16169,N_15847);
nor U16507 (N_16507,N_15667,N_16136);
nor U16508 (N_16508,N_15649,N_16008);
and U16509 (N_16509,N_15880,N_15822);
xor U16510 (N_16510,N_15706,N_16090);
nand U16511 (N_16511,N_15753,N_16061);
xor U16512 (N_16512,N_15822,N_15904);
nor U16513 (N_16513,N_16178,N_15933);
nand U16514 (N_16514,N_15741,N_15977);
nor U16515 (N_16515,N_15744,N_16146);
nor U16516 (N_16516,N_15924,N_16162);
or U16517 (N_16517,N_15928,N_15845);
xnor U16518 (N_16518,N_15785,N_15784);
and U16519 (N_16519,N_15964,N_16035);
xor U16520 (N_16520,N_15987,N_16027);
xnor U16521 (N_16521,N_15673,N_15845);
and U16522 (N_16522,N_16070,N_15850);
xor U16523 (N_16523,N_15864,N_15636);
or U16524 (N_16524,N_15636,N_15757);
nor U16525 (N_16525,N_16032,N_16018);
xor U16526 (N_16526,N_15812,N_15917);
xnor U16527 (N_16527,N_15707,N_16197);
xor U16528 (N_16528,N_15947,N_16151);
nor U16529 (N_16529,N_16012,N_15785);
xnor U16530 (N_16530,N_15671,N_15926);
and U16531 (N_16531,N_15786,N_16185);
nand U16532 (N_16532,N_16005,N_16064);
and U16533 (N_16533,N_15974,N_16105);
and U16534 (N_16534,N_16124,N_16057);
xor U16535 (N_16535,N_16179,N_15694);
and U16536 (N_16536,N_16164,N_16183);
and U16537 (N_16537,N_16125,N_15970);
or U16538 (N_16538,N_15666,N_16138);
nand U16539 (N_16539,N_15735,N_16074);
xnor U16540 (N_16540,N_15657,N_16168);
or U16541 (N_16541,N_16038,N_15858);
and U16542 (N_16542,N_15668,N_15769);
nor U16543 (N_16543,N_15634,N_15915);
nor U16544 (N_16544,N_15657,N_15986);
nor U16545 (N_16545,N_15985,N_15855);
and U16546 (N_16546,N_15655,N_15895);
xor U16547 (N_16547,N_16161,N_15973);
nor U16548 (N_16548,N_15669,N_15668);
xnor U16549 (N_16549,N_15888,N_15982);
nand U16550 (N_16550,N_16069,N_15800);
and U16551 (N_16551,N_15931,N_15726);
nor U16552 (N_16552,N_15606,N_15961);
or U16553 (N_16553,N_16160,N_15907);
or U16554 (N_16554,N_15865,N_15911);
xnor U16555 (N_16555,N_16044,N_15786);
nor U16556 (N_16556,N_16059,N_16111);
nand U16557 (N_16557,N_15746,N_15899);
nand U16558 (N_16558,N_15786,N_16191);
or U16559 (N_16559,N_15752,N_16125);
xor U16560 (N_16560,N_15905,N_16001);
nand U16561 (N_16561,N_15661,N_16141);
nor U16562 (N_16562,N_15953,N_15704);
or U16563 (N_16563,N_16126,N_16093);
nand U16564 (N_16564,N_15910,N_15926);
nand U16565 (N_16565,N_16026,N_16112);
and U16566 (N_16566,N_16075,N_15631);
or U16567 (N_16567,N_16061,N_15946);
xnor U16568 (N_16568,N_15844,N_16187);
nor U16569 (N_16569,N_16052,N_15945);
nor U16570 (N_16570,N_16049,N_15848);
and U16571 (N_16571,N_16023,N_15822);
and U16572 (N_16572,N_16004,N_15758);
and U16573 (N_16573,N_16173,N_15723);
nand U16574 (N_16574,N_15831,N_15861);
nor U16575 (N_16575,N_15602,N_15766);
nand U16576 (N_16576,N_16038,N_16002);
or U16577 (N_16577,N_15762,N_15790);
xnor U16578 (N_16578,N_15638,N_15925);
xnor U16579 (N_16579,N_16074,N_15872);
and U16580 (N_16580,N_15896,N_15616);
nand U16581 (N_16581,N_16008,N_16122);
nand U16582 (N_16582,N_15726,N_15981);
nor U16583 (N_16583,N_16194,N_16101);
nand U16584 (N_16584,N_15689,N_16134);
or U16585 (N_16585,N_15637,N_15689);
nor U16586 (N_16586,N_15606,N_16055);
or U16587 (N_16587,N_15620,N_15733);
nand U16588 (N_16588,N_15858,N_15762);
nand U16589 (N_16589,N_15734,N_15977);
xor U16590 (N_16590,N_15824,N_15618);
nand U16591 (N_16591,N_16002,N_16065);
or U16592 (N_16592,N_16126,N_15859);
or U16593 (N_16593,N_15630,N_15847);
and U16594 (N_16594,N_16171,N_15905);
or U16595 (N_16595,N_15708,N_15965);
xnor U16596 (N_16596,N_15962,N_15974);
xnor U16597 (N_16597,N_16063,N_15916);
xor U16598 (N_16598,N_15659,N_15828);
or U16599 (N_16599,N_15657,N_15686);
and U16600 (N_16600,N_15718,N_16096);
and U16601 (N_16601,N_15928,N_15630);
nor U16602 (N_16602,N_16194,N_16070);
nand U16603 (N_16603,N_16167,N_15976);
xnor U16604 (N_16604,N_15946,N_16075);
nor U16605 (N_16605,N_16065,N_15988);
xor U16606 (N_16606,N_16167,N_15680);
and U16607 (N_16607,N_16045,N_15977);
and U16608 (N_16608,N_15796,N_15993);
or U16609 (N_16609,N_16015,N_15838);
nand U16610 (N_16610,N_15990,N_15613);
nor U16611 (N_16611,N_15625,N_15982);
xor U16612 (N_16612,N_15773,N_16093);
xor U16613 (N_16613,N_15748,N_16009);
and U16614 (N_16614,N_15922,N_16045);
nor U16615 (N_16615,N_16068,N_15776);
xnor U16616 (N_16616,N_15918,N_15988);
xnor U16617 (N_16617,N_15765,N_16189);
and U16618 (N_16618,N_15640,N_15738);
nor U16619 (N_16619,N_15832,N_16154);
or U16620 (N_16620,N_15715,N_15721);
and U16621 (N_16621,N_15709,N_15983);
nand U16622 (N_16622,N_15848,N_15759);
or U16623 (N_16623,N_15736,N_16174);
xor U16624 (N_16624,N_15875,N_16081);
nor U16625 (N_16625,N_15863,N_15809);
xor U16626 (N_16626,N_16041,N_16164);
xor U16627 (N_16627,N_15936,N_15607);
and U16628 (N_16628,N_15831,N_15616);
nand U16629 (N_16629,N_15719,N_16118);
or U16630 (N_16630,N_16109,N_15725);
nor U16631 (N_16631,N_15958,N_16056);
or U16632 (N_16632,N_15793,N_15600);
and U16633 (N_16633,N_16046,N_15752);
or U16634 (N_16634,N_15975,N_15712);
and U16635 (N_16635,N_16118,N_15738);
and U16636 (N_16636,N_15820,N_16047);
xnor U16637 (N_16637,N_16148,N_15792);
nand U16638 (N_16638,N_15771,N_16003);
and U16639 (N_16639,N_16034,N_15986);
xor U16640 (N_16640,N_15750,N_15948);
nand U16641 (N_16641,N_15610,N_16102);
nor U16642 (N_16642,N_16176,N_15644);
or U16643 (N_16643,N_16130,N_15851);
nor U16644 (N_16644,N_16084,N_16086);
nor U16645 (N_16645,N_16108,N_15936);
or U16646 (N_16646,N_15734,N_15932);
and U16647 (N_16647,N_15626,N_16121);
nand U16648 (N_16648,N_16092,N_15752);
xor U16649 (N_16649,N_15727,N_15933);
nor U16650 (N_16650,N_15738,N_15802);
nand U16651 (N_16651,N_15825,N_16198);
or U16652 (N_16652,N_15832,N_15774);
xnor U16653 (N_16653,N_15707,N_15929);
or U16654 (N_16654,N_16117,N_15807);
xnor U16655 (N_16655,N_16193,N_16064);
nand U16656 (N_16656,N_16112,N_15777);
nor U16657 (N_16657,N_15605,N_16153);
nor U16658 (N_16658,N_16021,N_15654);
xnor U16659 (N_16659,N_15760,N_16124);
nor U16660 (N_16660,N_15820,N_16059);
nor U16661 (N_16661,N_15627,N_16124);
xnor U16662 (N_16662,N_16000,N_15884);
nor U16663 (N_16663,N_15697,N_15991);
nand U16664 (N_16664,N_15601,N_16182);
nand U16665 (N_16665,N_16184,N_16136);
nand U16666 (N_16666,N_15764,N_15972);
nor U16667 (N_16667,N_15696,N_15800);
and U16668 (N_16668,N_15986,N_15701);
nor U16669 (N_16669,N_16197,N_16100);
and U16670 (N_16670,N_16065,N_16051);
or U16671 (N_16671,N_16013,N_15853);
nor U16672 (N_16672,N_15749,N_16194);
xor U16673 (N_16673,N_16157,N_15928);
nor U16674 (N_16674,N_15741,N_15902);
nor U16675 (N_16675,N_15662,N_15986);
or U16676 (N_16676,N_15834,N_16149);
nor U16677 (N_16677,N_15940,N_15934);
nor U16678 (N_16678,N_15630,N_15994);
and U16679 (N_16679,N_15602,N_15638);
and U16680 (N_16680,N_15681,N_16161);
xnor U16681 (N_16681,N_16065,N_15812);
and U16682 (N_16682,N_16152,N_15867);
nand U16683 (N_16683,N_15825,N_15738);
or U16684 (N_16684,N_15793,N_15787);
or U16685 (N_16685,N_15670,N_15920);
nor U16686 (N_16686,N_15868,N_16078);
xor U16687 (N_16687,N_16092,N_15722);
nand U16688 (N_16688,N_16066,N_15944);
nand U16689 (N_16689,N_15692,N_16132);
and U16690 (N_16690,N_16055,N_15722);
or U16691 (N_16691,N_15912,N_15852);
nand U16692 (N_16692,N_15950,N_15956);
and U16693 (N_16693,N_16042,N_16114);
or U16694 (N_16694,N_15638,N_15681);
and U16695 (N_16695,N_16195,N_16120);
nor U16696 (N_16696,N_15969,N_15929);
nor U16697 (N_16697,N_15862,N_16132);
and U16698 (N_16698,N_15789,N_16134);
or U16699 (N_16699,N_16023,N_15652);
nand U16700 (N_16700,N_15756,N_15728);
nand U16701 (N_16701,N_16155,N_15651);
nor U16702 (N_16702,N_15897,N_15885);
xor U16703 (N_16703,N_15823,N_15670);
and U16704 (N_16704,N_16129,N_15928);
nor U16705 (N_16705,N_15892,N_15872);
or U16706 (N_16706,N_15895,N_15947);
nor U16707 (N_16707,N_15855,N_16068);
and U16708 (N_16708,N_16097,N_15691);
nor U16709 (N_16709,N_16169,N_15831);
nor U16710 (N_16710,N_15713,N_15607);
nor U16711 (N_16711,N_15712,N_16008);
and U16712 (N_16712,N_16116,N_15924);
or U16713 (N_16713,N_15682,N_15982);
and U16714 (N_16714,N_16152,N_15941);
or U16715 (N_16715,N_16179,N_15983);
xor U16716 (N_16716,N_15691,N_15707);
nor U16717 (N_16717,N_16088,N_15993);
and U16718 (N_16718,N_15713,N_15997);
or U16719 (N_16719,N_15702,N_15989);
nor U16720 (N_16720,N_15619,N_16198);
and U16721 (N_16721,N_15627,N_16146);
xnor U16722 (N_16722,N_16187,N_15837);
or U16723 (N_16723,N_15853,N_15745);
and U16724 (N_16724,N_15980,N_15636);
or U16725 (N_16725,N_16169,N_16032);
xor U16726 (N_16726,N_16028,N_15837);
nand U16727 (N_16727,N_15683,N_15704);
nand U16728 (N_16728,N_15726,N_15839);
and U16729 (N_16729,N_16044,N_15850);
xor U16730 (N_16730,N_15831,N_16060);
nor U16731 (N_16731,N_15800,N_15982);
nor U16732 (N_16732,N_15683,N_15994);
and U16733 (N_16733,N_16035,N_16088);
or U16734 (N_16734,N_15605,N_15995);
or U16735 (N_16735,N_16121,N_16137);
nor U16736 (N_16736,N_15680,N_16098);
or U16737 (N_16737,N_16187,N_16042);
or U16738 (N_16738,N_15632,N_16150);
or U16739 (N_16739,N_15857,N_15668);
or U16740 (N_16740,N_15947,N_15821);
and U16741 (N_16741,N_15736,N_15916);
or U16742 (N_16742,N_15622,N_15982);
nand U16743 (N_16743,N_15663,N_16136);
nand U16744 (N_16744,N_16100,N_16090);
and U16745 (N_16745,N_16122,N_15817);
nand U16746 (N_16746,N_15655,N_15625);
and U16747 (N_16747,N_15730,N_15706);
nor U16748 (N_16748,N_16180,N_15625);
nand U16749 (N_16749,N_16068,N_15904);
xnor U16750 (N_16750,N_15702,N_16171);
xnor U16751 (N_16751,N_15689,N_15788);
nand U16752 (N_16752,N_16031,N_15740);
xor U16753 (N_16753,N_15623,N_16050);
nand U16754 (N_16754,N_15967,N_16079);
nand U16755 (N_16755,N_15696,N_15995);
xor U16756 (N_16756,N_15901,N_15734);
and U16757 (N_16757,N_15646,N_16062);
xor U16758 (N_16758,N_16088,N_16132);
and U16759 (N_16759,N_15850,N_15968);
and U16760 (N_16760,N_15724,N_15956);
nand U16761 (N_16761,N_16071,N_16078);
xnor U16762 (N_16762,N_16161,N_15639);
nor U16763 (N_16763,N_16025,N_16149);
xor U16764 (N_16764,N_15931,N_15690);
or U16765 (N_16765,N_16049,N_15893);
and U16766 (N_16766,N_15982,N_16162);
nand U16767 (N_16767,N_16103,N_15786);
or U16768 (N_16768,N_15829,N_15610);
nor U16769 (N_16769,N_16112,N_15968);
or U16770 (N_16770,N_15942,N_15772);
and U16771 (N_16771,N_16064,N_15752);
nand U16772 (N_16772,N_15878,N_15789);
nor U16773 (N_16773,N_16100,N_16018);
and U16774 (N_16774,N_16021,N_15886);
nand U16775 (N_16775,N_16170,N_15944);
or U16776 (N_16776,N_15987,N_15803);
nor U16777 (N_16777,N_15955,N_15851);
and U16778 (N_16778,N_15694,N_15839);
nor U16779 (N_16779,N_15776,N_15960);
xor U16780 (N_16780,N_16186,N_15882);
xor U16781 (N_16781,N_15966,N_16178);
xnor U16782 (N_16782,N_15911,N_15859);
nor U16783 (N_16783,N_16061,N_15629);
nor U16784 (N_16784,N_15889,N_16161);
xnor U16785 (N_16785,N_15652,N_15935);
nand U16786 (N_16786,N_15646,N_16182);
nand U16787 (N_16787,N_15657,N_15752);
nand U16788 (N_16788,N_15640,N_15743);
or U16789 (N_16789,N_15889,N_16095);
or U16790 (N_16790,N_16008,N_15865);
nor U16791 (N_16791,N_16141,N_15664);
nand U16792 (N_16792,N_16062,N_15851);
nand U16793 (N_16793,N_15918,N_15920);
xor U16794 (N_16794,N_15664,N_15834);
xor U16795 (N_16795,N_16051,N_15911);
nor U16796 (N_16796,N_15787,N_15658);
nand U16797 (N_16797,N_16045,N_16124);
or U16798 (N_16798,N_15720,N_15949);
nand U16799 (N_16799,N_16127,N_15611);
xor U16800 (N_16800,N_16309,N_16556);
nand U16801 (N_16801,N_16694,N_16224);
nand U16802 (N_16802,N_16447,N_16413);
nand U16803 (N_16803,N_16263,N_16281);
and U16804 (N_16804,N_16215,N_16517);
nor U16805 (N_16805,N_16227,N_16350);
nand U16806 (N_16806,N_16703,N_16418);
and U16807 (N_16807,N_16608,N_16532);
xor U16808 (N_16808,N_16237,N_16654);
and U16809 (N_16809,N_16799,N_16425);
nor U16810 (N_16810,N_16376,N_16226);
and U16811 (N_16811,N_16409,N_16445);
xnor U16812 (N_16812,N_16559,N_16613);
nand U16813 (N_16813,N_16718,N_16455);
xor U16814 (N_16814,N_16500,N_16213);
and U16815 (N_16815,N_16543,N_16744);
nor U16816 (N_16816,N_16553,N_16468);
or U16817 (N_16817,N_16364,N_16444);
nor U16818 (N_16818,N_16489,N_16552);
and U16819 (N_16819,N_16358,N_16763);
nand U16820 (N_16820,N_16235,N_16363);
nor U16821 (N_16821,N_16776,N_16443);
xor U16822 (N_16822,N_16317,N_16473);
or U16823 (N_16823,N_16259,N_16393);
and U16824 (N_16824,N_16360,N_16507);
nor U16825 (N_16825,N_16678,N_16704);
nor U16826 (N_16826,N_16539,N_16380);
nand U16827 (N_16827,N_16382,N_16446);
nor U16828 (N_16828,N_16297,N_16333);
and U16829 (N_16829,N_16492,N_16529);
or U16830 (N_16830,N_16330,N_16672);
xnor U16831 (N_16831,N_16274,N_16467);
xor U16832 (N_16832,N_16684,N_16448);
nand U16833 (N_16833,N_16547,N_16244);
nand U16834 (N_16834,N_16220,N_16412);
and U16835 (N_16835,N_16739,N_16522);
xnor U16836 (N_16836,N_16784,N_16427);
nor U16837 (N_16837,N_16696,N_16479);
nand U16838 (N_16838,N_16276,N_16219);
xnor U16839 (N_16839,N_16581,N_16688);
nand U16840 (N_16840,N_16262,N_16241);
and U16841 (N_16841,N_16301,N_16622);
nor U16842 (N_16842,N_16261,N_16247);
or U16843 (N_16843,N_16214,N_16527);
and U16844 (N_16844,N_16604,N_16668);
xor U16845 (N_16845,N_16757,N_16269);
and U16846 (N_16846,N_16755,N_16795);
or U16847 (N_16847,N_16779,N_16586);
xor U16848 (N_16848,N_16619,N_16599);
and U16849 (N_16849,N_16629,N_16457);
nand U16850 (N_16850,N_16571,N_16416);
or U16851 (N_16851,N_16524,N_16582);
nand U16852 (N_16852,N_16595,N_16521);
nand U16853 (N_16853,N_16496,N_16525);
nand U16854 (N_16854,N_16265,N_16440);
nand U16855 (N_16855,N_16652,N_16614);
xor U16856 (N_16856,N_16284,N_16669);
xor U16857 (N_16857,N_16450,N_16208);
nand U16858 (N_16858,N_16796,N_16502);
xor U16859 (N_16859,N_16501,N_16794);
nor U16860 (N_16860,N_16673,N_16603);
xnor U16861 (N_16861,N_16609,N_16729);
nand U16862 (N_16862,N_16615,N_16740);
xor U16863 (N_16863,N_16697,N_16216);
xor U16864 (N_16864,N_16706,N_16751);
nor U16865 (N_16865,N_16289,N_16712);
or U16866 (N_16866,N_16228,N_16731);
nor U16867 (N_16867,N_16748,N_16365);
xnor U16868 (N_16868,N_16437,N_16592);
xnor U16869 (N_16869,N_16737,N_16632);
and U16870 (N_16870,N_16370,N_16346);
or U16871 (N_16871,N_16415,N_16429);
or U16872 (N_16872,N_16331,N_16223);
and U16873 (N_16873,N_16225,N_16464);
nor U16874 (N_16874,N_16232,N_16465);
nand U16875 (N_16875,N_16480,N_16229);
or U16876 (N_16876,N_16400,N_16371);
and U16877 (N_16877,N_16327,N_16466);
or U16878 (N_16878,N_16620,N_16666);
and U16879 (N_16879,N_16377,N_16659);
xnor U16880 (N_16880,N_16385,N_16563);
or U16881 (N_16881,N_16670,N_16775);
and U16882 (N_16882,N_16639,N_16733);
nor U16883 (N_16883,N_16353,N_16372);
nor U16884 (N_16884,N_16456,N_16637);
nor U16885 (N_16885,N_16329,N_16319);
or U16886 (N_16886,N_16342,N_16352);
xor U16887 (N_16887,N_16252,N_16635);
or U16888 (N_16888,N_16497,N_16407);
nor U16889 (N_16889,N_16575,N_16302);
nand U16890 (N_16890,N_16288,N_16207);
and U16891 (N_16891,N_16630,N_16290);
nor U16892 (N_16892,N_16769,N_16756);
or U16893 (N_16893,N_16222,N_16475);
xnor U16894 (N_16894,N_16246,N_16461);
xnor U16895 (N_16895,N_16405,N_16598);
or U16896 (N_16896,N_16625,N_16686);
nor U16897 (N_16897,N_16515,N_16294);
or U16898 (N_16898,N_16537,N_16633);
or U16899 (N_16899,N_16390,N_16312);
xnor U16900 (N_16900,N_16495,N_16375);
and U16901 (N_16901,N_16588,N_16477);
or U16902 (N_16902,N_16391,N_16727);
nor U16903 (N_16903,N_16260,N_16538);
and U16904 (N_16904,N_16408,N_16218);
or U16905 (N_16905,N_16789,N_16255);
xor U16906 (N_16906,N_16315,N_16430);
or U16907 (N_16907,N_16541,N_16610);
xnor U16908 (N_16908,N_16568,N_16798);
nand U16909 (N_16909,N_16257,N_16531);
nand U16910 (N_16910,N_16422,N_16303);
and U16911 (N_16911,N_16253,N_16745);
or U16912 (N_16912,N_16759,N_16264);
and U16913 (N_16913,N_16387,N_16460);
or U16914 (N_16914,N_16535,N_16411);
nand U16915 (N_16915,N_16518,N_16771);
and U16916 (N_16916,N_16548,N_16643);
or U16917 (N_16917,N_16349,N_16243);
nand U16918 (N_16918,N_16476,N_16392);
nor U16919 (N_16919,N_16549,N_16296);
or U16920 (N_16920,N_16238,N_16627);
nand U16921 (N_16921,N_16750,N_16722);
and U16922 (N_16922,N_16557,N_16396);
nand U16923 (N_16923,N_16277,N_16470);
nor U16924 (N_16924,N_16645,N_16715);
and U16925 (N_16925,N_16641,N_16356);
xor U16926 (N_16926,N_16487,N_16647);
xnor U16927 (N_16927,N_16761,N_16732);
xnor U16928 (N_16928,N_16449,N_16401);
nand U16929 (N_16929,N_16601,N_16359);
nand U16930 (N_16930,N_16690,N_16693);
nand U16931 (N_16931,N_16587,N_16590);
nand U16932 (N_16932,N_16459,N_16323);
nor U16933 (N_16933,N_16683,N_16310);
or U16934 (N_16934,N_16602,N_16767);
nand U16935 (N_16935,N_16245,N_16607);
or U16936 (N_16936,N_16504,N_16511);
or U16937 (N_16937,N_16283,N_16658);
nor U16938 (N_16938,N_16583,N_16488);
nand U16939 (N_16939,N_16250,N_16741);
and U16940 (N_16940,N_16536,N_16716);
nand U16941 (N_16941,N_16728,N_16591);
xnor U16942 (N_16942,N_16505,N_16558);
and U16943 (N_16943,N_16378,N_16562);
and U16944 (N_16944,N_16648,N_16785);
or U16945 (N_16945,N_16691,N_16777);
and U16946 (N_16946,N_16542,N_16702);
nor U16947 (N_16947,N_16597,N_16644);
and U16948 (N_16948,N_16486,N_16206);
nand U16949 (N_16949,N_16221,N_16273);
xor U16950 (N_16950,N_16786,N_16337);
nor U16951 (N_16951,N_16438,N_16793);
and U16952 (N_16952,N_16249,N_16369);
nor U16953 (N_16953,N_16423,N_16490);
or U16954 (N_16954,N_16316,N_16660);
nor U16955 (N_16955,N_16338,N_16394);
and U16956 (N_16956,N_16267,N_16624);
nor U16957 (N_16957,N_16279,N_16334);
nor U16958 (N_16958,N_16421,N_16540);
nand U16959 (N_16959,N_16720,N_16402);
or U16960 (N_16960,N_16388,N_16503);
xor U16961 (N_16961,N_16636,N_16469);
nor U16962 (N_16962,N_16367,N_16574);
or U16963 (N_16963,N_16512,N_16485);
nand U16964 (N_16964,N_16254,N_16424);
or U16965 (N_16965,N_16420,N_16291);
nor U16966 (N_16966,N_16345,N_16239);
xnor U16967 (N_16967,N_16617,N_16406);
nand U16968 (N_16968,N_16471,N_16311);
and U16969 (N_16969,N_16256,N_16593);
and U16970 (N_16970,N_16355,N_16596);
nor U16971 (N_16971,N_16714,N_16640);
and U16972 (N_16972,N_16634,N_16736);
or U16973 (N_16973,N_16546,N_16711);
xor U16974 (N_16974,N_16621,N_16506);
nor U16975 (N_16975,N_16493,N_16236);
and U16976 (N_16976,N_16509,N_16653);
nand U16977 (N_16977,N_16560,N_16677);
nand U16978 (N_16978,N_16611,N_16278);
nor U16979 (N_16979,N_16667,N_16498);
nor U16980 (N_16980,N_16638,N_16764);
or U16981 (N_16981,N_16680,N_16307);
and U16982 (N_16982,N_16395,N_16272);
and U16983 (N_16983,N_16554,N_16211);
xor U16984 (N_16984,N_16730,N_16724);
and U16985 (N_16985,N_16441,N_16682);
nand U16986 (N_16986,N_16758,N_16550);
nor U16987 (N_16987,N_16725,N_16605);
nand U16988 (N_16988,N_16201,N_16293);
xnor U16989 (N_16989,N_16651,N_16780);
nor U16990 (N_16990,N_16580,N_16404);
nand U16991 (N_16991,N_16689,N_16204);
nor U16992 (N_16992,N_16526,N_16205);
nor U16993 (N_16993,N_16735,N_16472);
or U16994 (N_16994,N_16569,N_16564);
nand U16995 (N_16995,N_16344,N_16774);
or U16996 (N_16996,N_16414,N_16499);
xnor U16997 (N_16997,N_16474,N_16510);
or U16998 (N_16998,N_16519,N_16212);
and U16999 (N_16999,N_16631,N_16778);
nand U17000 (N_17000,N_16282,N_16734);
xnor U17001 (N_17001,N_16452,N_16585);
nand U17002 (N_17002,N_16579,N_16671);
nand U17003 (N_17003,N_16544,N_16772);
and U17004 (N_17004,N_16719,N_16626);
and U17005 (N_17005,N_16292,N_16742);
nor U17006 (N_17006,N_16433,N_16687);
or U17007 (N_17007,N_16584,N_16271);
nand U17008 (N_17008,N_16322,N_16484);
nor U17009 (N_17009,N_16379,N_16304);
and U17010 (N_17010,N_16781,N_16721);
or U17011 (N_17011,N_16747,N_16663);
xnor U17012 (N_17012,N_16577,N_16661);
and U17013 (N_17013,N_16523,N_16708);
nand U17014 (N_17014,N_16534,N_16381);
and U17015 (N_17015,N_16746,N_16770);
xnor U17016 (N_17016,N_16508,N_16528);
xor U17017 (N_17017,N_16341,N_16326);
or U17018 (N_17018,N_16578,N_16209);
nor U17019 (N_17019,N_16270,N_16618);
xnor U17020 (N_17020,N_16695,N_16463);
or U17021 (N_17021,N_16399,N_16374);
xor U17022 (N_17022,N_16428,N_16752);
nor U17023 (N_17023,N_16516,N_16646);
nor U17024 (N_17024,N_16328,N_16572);
or U17025 (N_17025,N_16797,N_16234);
xnor U17026 (N_17026,N_16681,N_16373);
nor U17027 (N_17027,N_16649,N_16612);
nand U17028 (N_17028,N_16567,N_16616);
nand U17029 (N_17029,N_16431,N_16545);
nand U17030 (N_17030,N_16332,N_16491);
xnor U17031 (N_17031,N_16231,N_16765);
nor U17032 (N_17032,N_16699,N_16240);
nand U17033 (N_17033,N_16242,N_16287);
and U17034 (N_17034,N_16709,N_16439);
xor U17035 (N_17035,N_16383,N_16674);
xor U17036 (N_17036,N_16664,N_16320);
nor U17037 (N_17037,N_16743,N_16513);
nand U17038 (N_17038,N_16478,N_16707);
nor U17039 (N_17039,N_16436,N_16295);
nand U17040 (N_17040,N_16650,N_16773);
and U17041 (N_17041,N_16749,N_16313);
xor U17042 (N_17042,N_16754,N_16386);
nand U17043 (N_17043,N_16266,N_16268);
and U17044 (N_17044,N_16453,N_16692);
nor U17045 (N_17045,N_16551,N_16665);
and U17046 (N_17046,N_16600,N_16642);
nand U17047 (N_17047,N_16410,N_16366);
xor U17048 (N_17048,N_16606,N_16361);
nand U17049 (N_17049,N_16717,N_16451);
and U17050 (N_17050,N_16657,N_16520);
xor U17051 (N_17051,N_16403,N_16442);
and U17052 (N_17052,N_16766,N_16335);
nand U17053 (N_17053,N_16790,N_16251);
or U17054 (N_17054,N_16482,N_16573);
or U17055 (N_17055,N_16753,N_16594);
xor U17056 (N_17056,N_16308,N_16299);
and U17057 (N_17057,N_16565,N_16306);
or U17058 (N_17058,N_16762,N_16738);
and U17059 (N_17059,N_16589,N_16280);
nor U17060 (N_17060,N_16791,N_16351);
xnor U17061 (N_17061,N_16726,N_16417);
xor U17062 (N_17062,N_16788,N_16655);
xor U17063 (N_17063,N_16555,N_16576);
nand U17064 (N_17064,N_16233,N_16210);
and U17065 (N_17065,N_16248,N_16723);
nor U17066 (N_17066,N_16792,N_16570);
nor U17067 (N_17067,N_16368,N_16389);
nor U17068 (N_17068,N_16700,N_16275);
or U17069 (N_17069,N_16676,N_16783);
or U17070 (N_17070,N_16533,N_16434);
nor U17071 (N_17071,N_16462,N_16398);
nor U17072 (N_17072,N_16494,N_16483);
or U17073 (N_17073,N_16343,N_16432);
and U17074 (N_17074,N_16454,N_16318);
and U17075 (N_17075,N_16514,N_16481);
and U17076 (N_17076,N_16217,N_16656);
or U17077 (N_17077,N_16662,N_16321);
nor U17078 (N_17078,N_16675,N_16384);
nand U17079 (N_17079,N_16679,N_16347);
xor U17080 (N_17080,N_16285,N_16354);
nor U17081 (N_17081,N_16701,N_16348);
xor U17082 (N_17082,N_16768,N_16298);
or U17083 (N_17083,N_16203,N_16357);
and U17084 (N_17084,N_16397,N_16435);
xnor U17085 (N_17085,N_16324,N_16362);
nand U17086 (N_17086,N_16325,N_16258);
nor U17087 (N_17087,N_16426,N_16230);
nor U17088 (N_17088,N_16458,N_16628);
or U17089 (N_17089,N_16340,N_16710);
nor U17090 (N_17090,N_16202,N_16782);
nand U17091 (N_17091,N_16286,N_16305);
or U17092 (N_17092,N_16698,N_16561);
and U17093 (N_17093,N_16339,N_16760);
and U17094 (N_17094,N_16200,N_16566);
nand U17095 (N_17095,N_16336,N_16705);
nand U17096 (N_17096,N_16713,N_16300);
or U17097 (N_17097,N_16530,N_16787);
nor U17098 (N_17098,N_16419,N_16685);
nor U17099 (N_17099,N_16623,N_16314);
nand U17100 (N_17100,N_16539,N_16723);
nand U17101 (N_17101,N_16733,N_16533);
nor U17102 (N_17102,N_16585,N_16460);
xnor U17103 (N_17103,N_16793,N_16412);
and U17104 (N_17104,N_16523,N_16532);
nor U17105 (N_17105,N_16246,N_16572);
nor U17106 (N_17106,N_16272,N_16574);
nor U17107 (N_17107,N_16615,N_16342);
or U17108 (N_17108,N_16261,N_16239);
or U17109 (N_17109,N_16438,N_16716);
nand U17110 (N_17110,N_16509,N_16590);
and U17111 (N_17111,N_16592,N_16474);
nand U17112 (N_17112,N_16491,N_16456);
nor U17113 (N_17113,N_16772,N_16409);
and U17114 (N_17114,N_16537,N_16504);
or U17115 (N_17115,N_16734,N_16202);
xor U17116 (N_17116,N_16687,N_16630);
xor U17117 (N_17117,N_16761,N_16592);
and U17118 (N_17118,N_16312,N_16294);
nor U17119 (N_17119,N_16426,N_16454);
nand U17120 (N_17120,N_16481,N_16303);
and U17121 (N_17121,N_16427,N_16747);
or U17122 (N_17122,N_16570,N_16439);
and U17123 (N_17123,N_16758,N_16234);
and U17124 (N_17124,N_16611,N_16784);
or U17125 (N_17125,N_16543,N_16760);
or U17126 (N_17126,N_16495,N_16291);
xor U17127 (N_17127,N_16216,N_16764);
nor U17128 (N_17128,N_16517,N_16782);
nand U17129 (N_17129,N_16500,N_16241);
and U17130 (N_17130,N_16677,N_16476);
xnor U17131 (N_17131,N_16635,N_16456);
nor U17132 (N_17132,N_16330,N_16455);
nand U17133 (N_17133,N_16784,N_16769);
xor U17134 (N_17134,N_16583,N_16690);
and U17135 (N_17135,N_16640,N_16648);
nor U17136 (N_17136,N_16443,N_16497);
nor U17137 (N_17137,N_16757,N_16332);
nand U17138 (N_17138,N_16480,N_16542);
and U17139 (N_17139,N_16541,N_16218);
nor U17140 (N_17140,N_16504,N_16536);
xor U17141 (N_17141,N_16652,N_16555);
and U17142 (N_17142,N_16755,N_16514);
and U17143 (N_17143,N_16439,N_16223);
xnor U17144 (N_17144,N_16418,N_16617);
xor U17145 (N_17145,N_16534,N_16460);
and U17146 (N_17146,N_16560,N_16429);
and U17147 (N_17147,N_16492,N_16604);
and U17148 (N_17148,N_16216,N_16767);
and U17149 (N_17149,N_16563,N_16402);
nand U17150 (N_17150,N_16255,N_16670);
and U17151 (N_17151,N_16643,N_16327);
xnor U17152 (N_17152,N_16590,N_16508);
and U17153 (N_17153,N_16225,N_16254);
or U17154 (N_17154,N_16718,N_16660);
and U17155 (N_17155,N_16291,N_16451);
and U17156 (N_17156,N_16406,N_16262);
and U17157 (N_17157,N_16619,N_16574);
nand U17158 (N_17158,N_16327,N_16636);
xnor U17159 (N_17159,N_16749,N_16507);
or U17160 (N_17160,N_16727,N_16619);
nand U17161 (N_17161,N_16588,N_16631);
and U17162 (N_17162,N_16695,N_16287);
nor U17163 (N_17163,N_16755,N_16215);
xor U17164 (N_17164,N_16422,N_16730);
or U17165 (N_17165,N_16496,N_16541);
and U17166 (N_17166,N_16796,N_16470);
nor U17167 (N_17167,N_16263,N_16301);
or U17168 (N_17168,N_16244,N_16694);
nand U17169 (N_17169,N_16670,N_16210);
xor U17170 (N_17170,N_16771,N_16241);
nand U17171 (N_17171,N_16509,N_16460);
or U17172 (N_17172,N_16726,N_16399);
xor U17173 (N_17173,N_16387,N_16594);
and U17174 (N_17174,N_16776,N_16722);
or U17175 (N_17175,N_16321,N_16550);
nand U17176 (N_17176,N_16484,N_16631);
or U17177 (N_17177,N_16375,N_16510);
or U17178 (N_17178,N_16495,N_16574);
xor U17179 (N_17179,N_16565,N_16674);
nand U17180 (N_17180,N_16797,N_16551);
or U17181 (N_17181,N_16729,N_16261);
nand U17182 (N_17182,N_16423,N_16594);
xor U17183 (N_17183,N_16764,N_16789);
nor U17184 (N_17184,N_16352,N_16331);
nand U17185 (N_17185,N_16331,N_16548);
nand U17186 (N_17186,N_16568,N_16483);
nor U17187 (N_17187,N_16565,N_16504);
nor U17188 (N_17188,N_16764,N_16531);
xor U17189 (N_17189,N_16568,N_16255);
and U17190 (N_17190,N_16244,N_16480);
nand U17191 (N_17191,N_16758,N_16536);
or U17192 (N_17192,N_16745,N_16697);
nand U17193 (N_17193,N_16297,N_16796);
and U17194 (N_17194,N_16705,N_16285);
and U17195 (N_17195,N_16613,N_16358);
or U17196 (N_17196,N_16452,N_16241);
and U17197 (N_17197,N_16431,N_16373);
nand U17198 (N_17198,N_16744,N_16550);
nor U17199 (N_17199,N_16450,N_16738);
nor U17200 (N_17200,N_16340,N_16506);
and U17201 (N_17201,N_16318,N_16333);
xor U17202 (N_17202,N_16686,N_16706);
nand U17203 (N_17203,N_16453,N_16582);
nand U17204 (N_17204,N_16239,N_16579);
or U17205 (N_17205,N_16768,N_16388);
nor U17206 (N_17206,N_16472,N_16355);
or U17207 (N_17207,N_16627,N_16210);
nand U17208 (N_17208,N_16738,N_16496);
nand U17209 (N_17209,N_16384,N_16657);
or U17210 (N_17210,N_16746,N_16411);
or U17211 (N_17211,N_16717,N_16270);
nand U17212 (N_17212,N_16693,N_16700);
and U17213 (N_17213,N_16476,N_16587);
nand U17214 (N_17214,N_16595,N_16421);
nand U17215 (N_17215,N_16218,N_16324);
nor U17216 (N_17216,N_16775,N_16375);
or U17217 (N_17217,N_16570,N_16378);
or U17218 (N_17218,N_16216,N_16680);
or U17219 (N_17219,N_16516,N_16730);
xor U17220 (N_17220,N_16211,N_16571);
or U17221 (N_17221,N_16489,N_16701);
xnor U17222 (N_17222,N_16544,N_16262);
nand U17223 (N_17223,N_16312,N_16769);
xnor U17224 (N_17224,N_16508,N_16431);
or U17225 (N_17225,N_16718,N_16707);
xnor U17226 (N_17226,N_16639,N_16418);
or U17227 (N_17227,N_16250,N_16764);
and U17228 (N_17228,N_16309,N_16300);
nor U17229 (N_17229,N_16689,N_16466);
xor U17230 (N_17230,N_16263,N_16540);
and U17231 (N_17231,N_16343,N_16639);
nor U17232 (N_17232,N_16639,N_16402);
or U17233 (N_17233,N_16688,N_16237);
and U17234 (N_17234,N_16495,N_16242);
and U17235 (N_17235,N_16538,N_16555);
xor U17236 (N_17236,N_16211,N_16324);
and U17237 (N_17237,N_16371,N_16677);
nand U17238 (N_17238,N_16207,N_16746);
xnor U17239 (N_17239,N_16517,N_16550);
xnor U17240 (N_17240,N_16675,N_16321);
and U17241 (N_17241,N_16265,N_16639);
or U17242 (N_17242,N_16200,N_16622);
nor U17243 (N_17243,N_16712,N_16664);
and U17244 (N_17244,N_16702,N_16392);
and U17245 (N_17245,N_16588,N_16278);
xnor U17246 (N_17246,N_16487,N_16341);
and U17247 (N_17247,N_16787,N_16796);
nor U17248 (N_17248,N_16764,N_16332);
nor U17249 (N_17249,N_16703,N_16577);
and U17250 (N_17250,N_16723,N_16404);
or U17251 (N_17251,N_16323,N_16547);
xor U17252 (N_17252,N_16782,N_16737);
nor U17253 (N_17253,N_16661,N_16628);
or U17254 (N_17254,N_16208,N_16514);
nand U17255 (N_17255,N_16323,N_16559);
nor U17256 (N_17256,N_16788,N_16529);
nand U17257 (N_17257,N_16562,N_16582);
xor U17258 (N_17258,N_16751,N_16709);
nand U17259 (N_17259,N_16696,N_16225);
or U17260 (N_17260,N_16447,N_16661);
and U17261 (N_17261,N_16288,N_16570);
and U17262 (N_17262,N_16536,N_16760);
nand U17263 (N_17263,N_16519,N_16209);
and U17264 (N_17264,N_16491,N_16601);
xor U17265 (N_17265,N_16678,N_16514);
nand U17266 (N_17266,N_16254,N_16516);
or U17267 (N_17267,N_16776,N_16529);
or U17268 (N_17268,N_16279,N_16590);
xnor U17269 (N_17269,N_16647,N_16657);
and U17270 (N_17270,N_16538,N_16295);
nor U17271 (N_17271,N_16330,N_16705);
and U17272 (N_17272,N_16436,N_16569);
or U17273 (N_17273,N_16537,N_16389);
xnor U17274 (N_17274,N_16342,N_16416);
xnor U17275 (N_17275,N_16619,N_16591);
or U17276 (N_17276,N_16285,N_16661);
nor U17277 (N_17277,N_16590,N_16610);
and U17278 (N_17278,N_16203,N_16615);
xnor U17279 (N_17279,N_16616,N_16773);
and U17280 (N_17280,N_16395,N_16226);
or U17281 (N_17281,N_16253,N_16509);
nor U17282 (N_17282,N_16376,N_16338);
and U17283 (N_17283,N_16667,N_16564);
nor U17284 (N_17284,N_16482,N_16326);
xnor U17285 (N_17285,N_16488,N_16310);
nor U17286 (N_17286,N_16420,N_16343);
nor U17287 (N_17287,N_16586,N_16646);
and U17288 (N_17288,N_16685,N_16451);
nand U17289 (N_17289,N_16669,N_16473);
xor U17290 (N_17290,N_16743,N_16220);
xnor U17291 (N_17291,N_16235,N_16234);
nand U17292 (N_17292,N_16212,N_16799);
or U17293 (N_17293,N_16357,N_16623);
nand U17294 (N_17294,N_16314,N_16456);
xnor U17295 (N_17295,N_16393,N_16670);
nand U17296 (N_17296,N_16391,N_16240);
xor U17297 (N_17297,N_16771,N_16314);
or U17298 (N_17298,N_16377,N_16585);
xor U17299 (N_17299,N_16335,N_16290);
nor U17300 (N_17300,N_16375,N_16616);
nand U17301 (N_17301,N_16661,N_16731);
or U17302 (N_17302,N_16751,N_16381);
and U17303 (N_17303,N_16250,N_16644);
nor U17304 (N_17304,N_16356,N_16352);
nor U17305 (N_17305,N_16614,N_16559);
xnor U17306 (N_17306,N_16343,N_16516);
and U17307 (N_17307,N_16578,N_16341);
or U17308 (N_17308,N_16309,N_16784);
or U17309 (N_17309,N_16604,N_16311);
nor U17310 (N_17310,N_16551,N_16341);
nand U17311 (N_17311,N_16513,N_16376);
or U17312 (N_17312,N_16768,N_16359);
and U17313 (N_17313,N_16343,N_16628);
and U17314 (N_17314,N_16445,N_16779);
nor U17315 (N_17315,N_16284,N_16781);
or U17316 (N_17316,N_16401,N_16589);
or U17317 (N_17317,N_16350,N_16432);
or U17318 (N_17318,N_16637,N_16257);
xor U17319 (N_17319,N_16555,N_16397);
xnor U17320 (N_17320,N_16511,N_16609);
nand U17321 (N_17321,N_16407,N_16690);
nor U17322 (N_17322,N_16735,N_16469);
xor U17323 (N_17323,N_16332,N_16431);
nor U17324 (N_17324,N_16525,N_16585);
xnor U17325 (N_17325,N_16618,N_16568);
xor U17326 (N_17326,N_16238,N_16208);
nor U17327 (N_17327,N_16288,N_16418);
or U17328 (N_17328,N_16794,N_16608);
and U17329 (N_17329,N_16486,N_16731);
nor U17330 (N_17330,N_16734,N_16259);
and U17331 (N_17331,N_16353,N_16720);
or U17332 (N_17332,N_16314,N_16201);
nor U17333 (N_17333,N_16466,N_16269);
nand U17334 (N_17334,N_16793,N_16541);
nand U17335 (N_17335,N_16329,N_16692);
and U17336 (N_17336,N_16380,N_16358);
and U17337 (N_17337,N_16235,N_16564);
nor U17338 (N_17338,N_16213,N_16389);
xnor U17339 (N_17339,N_16433,N_16317);
nand U17340 (N_17340,N_16577,N_16532);
xor U17341 (N_17341,N_16412,N_16591);
and U17342 (N_17342,N_16440,N_16780);
nand U17343 (N_17343,N_16654,N_16292);
and U17344 (N_17344,N_16399,N_16259);
and U17345 (N_17345,N_16514,N_16703);
nor U17346 (N_17346,N_16265,N_16204);
or U17347 (N_17347,N_16653,N_16325);
xor U17348 (N_17348,N_16763,N_16313);
nand U17349 (N_17349,N_16722,N_16745);
nand U17350 (N_17350,N_16746,N_16427);
or U17351 (N_17351,N_16669,N_16749);
or U17352 (N_17352,N_16653,N_16797);
nor U17353 (N_17353,N_16750,N_16658);
and U17354 (N_17354,N_16350,N_16729);
and U17355 (N_17355,N_16778,N_16655);
or U17356 (N_17356,N_16661,N_16714);
and U17357 (N_17357,N_16790,N_16260);
nor U17358 (N_17358,N_16671,N_16465);
and U17359 (N_17359,N_16331,N_16457);
or U17360 (N_17360,N_16371,N_16365);
nand U17361 (N_17361,N_16544,N_16694);
xor U17362 (N_17362,N_16560,N_16664);
xor U17363 (N_17363,N_16271,N_16537);
and U17364 (N_17364,N_16399,N_16276);
xnor U17365 (N_17365,N_16657,N_16250);
or U17366 (N_17366,N_16704,N_16322);
and U17367 (N_17367,N_16595,N_16726);
nand U17368 (N_17368,N_16703,N_16727);
nor U17369 (N_17369,N_16499,N_16488);
nor U17370 (N_17370,N_16412,N_16503);
or U17371 (N_17371,N_16313,N_16237);
or U17372 (N_17372,N_16573,N_16369);
nand U17373 (N_17373,N_16588,N_16310);
or U17374 (N_17374,N_16514,N_16237);
and U17375 (N_17375,N_16723,N_16258);
nand U17376 (N_17376,N_16428,N_16728);
and U17377 (N_17377,N_16605,N_16702);
xnor U17378 (N_17378,N_16629,N_16724);
or U17379 (N_17379,N_16640,N_16500);
nor U17380 (N_17380,N_16457,N_16635);
nor U17381 (N_17381,N_16760,N_16785);
or U17382 (N_17382,N_16484,N_16717);
nor U17383 (N_17383,N_16311,N_16310);
nor U17384 (N_17384,N_16633,N_16608);
or U17385 (N_17385,N_16570,N_16572);
or U17386 (N_17386,N_16765,N_16456);
and U17387 (N_17387,N_16316,N_16284);
and U17388 (N_17388,N_16731,N_16570);
nand U17389 (N_17389,N_16438,N_16315);
nand U17390 (N_17390,N_16585,N_16740);
and U17391 (N_17391,N_16359,N_16701);
xor U17392 (N_17392,N_16255,N_16235);
xnor U17393 (N_17393,N_16252,N_16332);
or U17394 (N_17394,N_16340,N_16640);
nand U17395 (N_17395,N_16566,N_16264);
xor U17396 (N_17396,N_16472,N_16554);
nor U17397 (N_17397,N_16698,N_16724);
and U17398 (N_17398,N_16468,N_16665);
and U17399 (N_17399,N_16790,N_16342);
xor U17400 (N_17400,N_17173,N_17109);
nand U17401 (N_17401,N_16980,N_17314);
and U17402 (N_17402,N_16916,N_16908);
nor U17403 (N_17403,N_16923,N_17203);
nor U17404 (N_17404,N_17299,N_17216);
or U17405 (N_17405,N_17289,N_17336);
and U17406 (N_17406,N_17330,N_17030);
xnor U17407 (N_17407,N_17175,N_17176);
nor U17408 (N_17408,N_17154,N_16894);
nand U17409 (N_17409,N_16988,N_17095);
nor U17410 (N_17410,N_16942,N_16833);
xnor U17411 (N_17411,N_17139,N_16843);
nor U17412 (N_17412,N_17145,N_16941);
nor U17413 (N_17413,N_17363,N_16956);
xor U17414 (N_17414,N_17353,N_17241);
nand U17415 (N_17415,N_16837,N_16889);
xnor U17416 (N_17416,N_16861,N_16917);
nand U17417 (N_17417,N_17047,N_17227);
and U17418 (N_17418,N_16817,N_17246);
xnor U17419 (N_17419,N_16966,N_17219);
and U17420 (N_17420,N_17191,N_17107);
nand U17421 (N_17421,N_16830,N_17122);
or U17422 (N_17422,N_17003,N_17206);
or U17423 (N_17423,N_16802,N_17218);
and U17424 (N_17424,N_17288,N_17204);
nor U17425 (N_17425,N_17129,N_16899);
nand U17426 (N_17426,N_17230,N_17036);
nand U17427 (N_17427,N_17275,N_17351);
nand U17428 (N_17428,N_16930,N_17048);
nor U17429 (N_17429,N_16847,N_17022);
nor U17430 (N_17430,N_17044,N_17225);
xor U17431 (N_17431,N_17380,N_17214);
xor U17432 (N_17432,N_16890,N_16807);
xor U17433 (N_17433,N_17012,N_16912);
nor U17434 (N_17434,N_16951,N_17372);
or U17435 (N_17435,N_17252,N_17328);
or U17436 (N_17436,N_17117,N_17237);
nor U17437 (N_17437,N_17053,N_17282);
nand U17438 (N_17438,N_16869,N_17358);
and U17439 (N_17439,N_16971,N_16927);
and U17440 (N_17440,N_16846,N_17050);
xnor U17441 (N_17441,N_16827,N_17256);
nor U17442 (N_17442,N_17049,N_17034);
nand U17443 (N_17443,N_16812,N_16961);
xor U17444 (N_17444,N_17069,N_17066);
or U17445 (N_17445,N_16829,N_16892);
nand U17446 (N_17446,N_16875,N_17322);
and U17447 (N_17447,N_16925,N_17113);
nand U17448 (N_17448,N_17199,N_16937);
or U17449 (N_17449,N_17338,N_17391);
xor U17450 (N_17450,N_17174,N_17323);
nand U17451 (N_17451,N_17248,N_16882);
xnor U17452 (N_17452,N_17133,N_17339);
nor U17453 (N_17453,N_16898,N_16852);
xor U17454 (N_17454,N_16881,N_17132);
xnor U17455 (N_17455,N_16987,N_17192);
xnor U17456 (N_17456,N_16953,N_17040);
xor U17457 (N_17457,N_17002,N_16835);
nand U17458 (N_17458,N_16858,N_17213);
xnor U17459 (N_17459,N_17155,N_16887);
and U17460 (N_17460,N_16945,N_17290);
xor U17461 (N_17461,N_17183,N_17032);
nor U17462 (N_17462,N_17123,N_17131);
nand U17463 (N_17463,N_16909,N_17115);
nor U17464 (N_17464,N_16914,N_17031);
xor U17465 (N_17465,N_17368,N_16960);
nor U17466 (N_17466,N_17148,N_17126);
nor U17467 (N_17467,N_17025,N_16863);
and U17468 (N_17468,N_16883,N_17268);
and U17469 (N_17469,N_17327,N_17217);
nor U17470 (N_17470,N_16986,N_17073);
or U17471 (N_17471,N_17271,N_17325);
xor U17472 (N_17472,N_16848,N_16928);
nor U17473 (N_17473,N_16813,N_17081);
nand U17474 (N_17474,N_16824,N_17096);
and U17475 (N_17475,N_16954,N_16996);
nor U17476 (N_17476,N_16976,N_16910);
and U17477 (N_17477,N_17394,N_17352);
or U17478 (N_17478,N_16845,N_17196);
nand U17479 (N_17479,N_16904,N_17181);
and U17480 (N_17480,N_16943,N_17251);
and U17481 (N_17481,N_17011,N_16839);
and U17482 (N_17482,N_17396,N_17104);
xor U17483 (N_17483,N_17138,N_16809);
or U17484 (N_17484,N_17112,N_17334);
nand U17485 (N_17485,N_16952,N_17153);
or U17486 (N_17486,N_17305,N_16978);
nand U17487 (N_17487,N_16977,N_17395);
xnor U17488 (N_17488,N_17114,N_17057);
xnor U17489 (N_17489,N_16993,N_17361);
or U17490 (N_17490,N_17038,N_17009);
nor U17491 (N_17491,N_17215,N_17267);
nand U17492 (N_17492,N_17228,N_16901);
nand U17493 (N_17493,N_17062,N_17164);
or U17494 (N_17494,N_16880,N_17033);
nand U17495 (N_17495,N_17209,N_17375);
and U17496 (N_17496,N_17234,N_17143);
xor U17497 (N_17497,N_16804,N_16849);
nor U17498 (N_17498,N_17318,N_16879);
nand U17499 (N_17499,N_16860,N_17223);
or U17500 (N_17500,N_17021,N_17356);
or U17501 (N_17501,N_16840,N_16962);
xor U17502 (N_17502,N_17399,N_16844);
or U17503 (N_17503,N_17370,N_17283);
nand U17504 (N_17504,N_16982,N_17151);
nand U17505 (N_17505,N_17158,N_17257);
xor U17506 (N_17506,N_17287,N_17130);
or U17507 (N_17507,N_17024,N_17377);
and U17508 (N_17508,N_17142,N_16874);
nor U17509 (N_17509,N_17125,N_17310);
or U17510 (N_17510,N_17397,N_17018);
xor U17511 (N_17511,N_17160,N_16929);
or U17512 (N_17512,N_17020,N_16876);
xnor U17513 (N_17513,N_17366,N_16877);
and U17514 (N_17514,N_17000,N_17278);
xor U17515 (N_17515,N_17019,N_17297);
nand U17516 (N_17516,N_17205,N_16826);
xor U17517 (N_17517,N_16949,N_17263);
xor U17518 (N_17518,N_17211,N_17393);
nand U17519 (N_17519,N_17269,N_16850);
nor U17520 (N_17520,N_17088,N_16854);
nor U17521 (N_17521,N_17382,N_16832);
and U17522 (N_17522,N_17208,N_17337);
xor U17523 (N_17523,N_17308,N_17277);
or U17524 (N_17524,N_16998,N_16969);
nor U17525 (N_17525,N_17304,N_17182);
or U17526 (N_17526,N_17065,N_17162);
nand U17527 (N_17527,N_16936,N_17159);
nand U17528 (N_17528,N_16800,N_16934);
nand U17529 (N_17529,N_17171,N_17312);
xor U17530 (N_17530,N_17200,N_17245);
nor U17531 (N_17531,N_17367,N_17386);
and U17532 (N_17532,N_17046,N_17015);
or U17533 (N_17533,N_16856,N_17070);
xor U17534 (N_17534,N_17309,N_17371);
nand U17535 (N_17535,N_17313,N_17186);
xnor U17536 (N_17536,N_17167,N_17398);
xnor U17537 (N_17537,N_16965,N_17101);
xor U17538 (N_17538,N_17307,N_16979);
and U17539 (N_17539,N_17381,N_17128);
xor U17540 (N_17540,N_16906,N_16924);
xnor U17541 (N_17541,N_17166,N_17333);
nand U17542 (N_17542,N_17387,N_16926);
xnor U17543 (N_17543,N_17127,N_17179);
xnor U17544 (N_17544,N_16821,N_17284);
or U17545 (N_17545,N_17043,N_17279);
nor U17546 (N_17546,N_17347,N_17094);
or U17547 (N_17547,N_17086,N_17212);
or U17548 (N_17548,N_17332,N_17074);
xnor U17549 (N_17549,N_17235,N_17343);
and U17550 (N_17550,N_17335,N_16918);
xor U17551 (N_17551,N_17004,N_17285);
and U17552 (N_17552,N_17005,N_17311);
and U17553 (N_17553,N_17258,N_17001);
and U17554 (N_17554,N_17222,N_16871);
xor U17555 (N_17555,N_16911,N_17080);
xnor U17556 (N_17556,N_17274,N_16873);
or U17557 (N_17557,N_17346,N_16920);
or U17558 (N_17558,N_17273,N_17071);
nor U17559 (N_17559,N_17354,N_17055);
xnor U17560 (N_17560,N_17303,N_17321);
xor U17561 (N_17561,N_16915,N_16963);
nor U17562 (N_17562,N_17326,N_17253);
nand U17563 (N_17563,N_17184,N_17302);
and U17564 (N_17564,N_16913,N_17374);
xor U17565 (N_17565,N_16985,N_16907);
and U17566 (N_17566,N_17341,N_16872);
or U17567 (N_17567,N_17098,N_16895);
nor U17568 (N_17568,N_17190,N_16975);
xnor U17569 (N_17569,N_17063,N_17238);
nor U17570 (N_17570,N_17232,N_17198);
nor U17571 (N_17571,N_17168,N_16967);
nor U17572 (N_17572,N_17260,N_17102);
xnor U17573 (N_17573,N_17137,N_17188);
or U17574 (N_17574,N_17239,N_17061);
nand U17575 (N_17575,N_17006,N_17250);
and U17576 (N_17576,N_17266,N_16878);
and U17577 (N_17577,N_17270,N_17082);
or U17578 (N_17578,N_17110,N_17317);
or U17579 (N_17579,N_16801,N_17017);
nand U17580 (N_17580,N_17085,N_16931);
nor U17581 (N_17581,N_17056,N_17296);
xor U17582 (N_17582,N_17300,N_16997);
and U17583 (N_17583,N_16818,N_17076);
or U17584 (N_17584,N_16825,N_16888);
or U17585 (N_17585,N_17195,N_16964);
xnor U17586 (N_17586,N_17344,N_17150);
and U17587 (N_17587,N_17345,N_17052);
xnor U17588 (N_17588,N_16959,N_17389);
nor U17589 (N_17589,N_17028,N_17280);
xnor U17590 (N_17590,N_17348,N_16851);
nor U17591 (N_17591,N_17185,N_17116);
nand U17592 (N_17592,N_17390,N_16973);
nor U17593 (N_17593,N_16855,N_17340);
nor U17594 (N_17594,N_16932,N_17255);
nor U17595 (N_17595,N_16838,N_17124);
and U17596 (N_17596,N_17320,N_16947);
xor U17597 (N_17597,N_17329,N_17178);
nand U17598 (N_17598,N_17315,N_17249);
or U17599 (N_17599,N_17058,N_17037);
and U17600 (N_17600,N_17295,N_16950);
or U17601 (N_17601,N_17149,N_17189);
and U17602 (N_17602,N_17265,N_16970);
nand U17603 (N_17603,N_17243,N_17023);
and U17604 (N_17604,N_16865,N_17362);
xnor U17605 (N_17605,N_17226,N_17210);
xor U17606 (N_17606,N_17383,N_17342);
xnor U17607 (N_17607,N_17201,N_17349);
nand U17608 (N_17608,N_17376,N_16811);
and U17609 (N_17609,N_17165,N_17286);
and U17610 (N_17610,N_17016,N_17259);
and U17611 (N_17611,N_17331,N_17077);
xor U17612 (N_17612,N_17156,N_16834);
nand U17613 (N_17613,N_17229,N_16893);
or U17614 (N_17614,N_16944,N_17301);
nor U17615 (N_17615,N_17068,N_17014);
xor U17616 (N_17616,N_16955,N_17097);
nor U17617 (N_17617,N_17294,N_17388);
xor U17618 (N_17618,N_16938,N_17378);
nand U17619 (N_17619,N_16822,N_17029);
nand U17620 (N_17620,N_17293,N_17045);
or U17621 (N_17621,N_16808,N_17254);
nor U17622 (N_17622,N_16995,N_17152);
and U17623 (N_17623,N_17261,N_17091);
nor U17624 (N_17624,N_16919,N_16983);
nor U17625 (N_17625,N_17008,N_16958);
nor U17626 (N_17626,N_16870,N_17197);
nand U17627 (N_17627,N_16922,N_17281);
and U17628 (N_17628,N_16900,N_16841);
or U17629 (N_17629,N_16884,N_17207);
or U17630 (N_17630,N_17316,N_17067);
or U17631 (N_17631,N_17035,N_17141);
or U17632 (N_17632,N_17392,N_17224);
nor U17633 (N_17633,N_17157,N_17100);
xor U17634 (N_17634,N_16828,N_17079);
and U17635 (N_17635,N_17359,N_17276);
nand U17636 (N_17636,N_17108,N_17136);
nor U17637 (N_17637,N_17240,N_17170);
and U17638 (N_17638,N_17144,N_16819);
nor U17639 (N_17639,N_17093,N_16885);
nand U17640 (N_17640,N_17120,N_16836);
nand U17641 (N_17641,N_17172,N_17121);
and U17642 (N_17642,N_17180,N_17291);
nand U17643 (N_17643,N_16989,N_17064);
nor U17644 (N_17644,N_17298,N_17010);
and U17645 (N_17645,N_16815,N_16891);
or U17646 (N_17646,N_16857,N_17357);
or U17647 (N_17647,N_17084,N_17134);
and U17648 (N_17648,N_17054,N_16940);
xor U17649 (N_17649,N_17072,N_16933);
and U17650 (N_17650,N_17272,N_16831);
nand U17651 (N_17651,N_17087,N_17105);
or U17652 (N_17652,N_17364,N_17146);
xnor U17653 (N_17653,N_17119,N_16902);
nand U17654 (N_17654,N_17051,N_16968);
xor U17655 (N_17655,N_16903,N_17194);
xor U17656 (N_17656,N_17089,N_17360);
or U17657 (N_17657,N_17373,N_17220);
or U17658 (N_17658,N_17147,N_17111);
and U17659 (N_17659,N_16896,N_17385);
or U17660 (N_17660,N_16897,N_17161);
nand U17661 (N_17661,N_17027,N_16984);
nand U17662 (N_17662,N_17177,N_17236);
nand U17663 (N_17663,N_17103,N_17306);
or U17664 (N_17664,N_16972,N_16810);
and U17665 (N_17665,N_16905,N_17355);
xnor U17666 (N_17666,N_17193,N_16990);
nor U17667 (N_17667,N_17379,N_17242);
xor U17668 (N_17668,N_16868,N_17233);
nor U17669 (N_17669,N_17135,N_16935);
nand U17670 (N_17670,N_16853,N_17202);
nor U17671 (N_17671,N_17106,N_16999);
nor U17672 (N_17672,N_16994,N_17042);
or U17673 (N_17673,N_16867,N_17350);
and U17674 (N_17674,N_16866,N_17118);
and U17675 (N_17675,N_17092,N_17264);
nor U17676 (N_17676,N_16862,N_17292);
or U17677 (N_17677,N_17221,N_17187);
xnor U17678 (N_17678,N_17384,N_17231);
xor U17679 (N_17679,N_16806,N_16991);
xor U17680 (N_17680,N_16823,N_17140);
or U17681 (N_17681,N_17163,N_16957);
nor U17682 (N_17682,N_17262,N_16939);
nand U17683 (N_17683,N_16803,N_17169);
xnor U17684 (N_17684,N_16992,N_16820);
nand U17685 (N_17685,N_16864,N_17324);
nand U17686 (N_17686,N_17078,N_17075);
nor U17687 (N_17687,N_16946,N_17060);
and U17688 (N_17688,N_16816,N_17365);
nand U17689 (N_17689,N_17026,N_17013);
or U17690 (N_17690,N_17247,N_17099);
or U17691 (N_17691,N_16859,N_17039);
or U17692 (N_17692,N_17090,N_16981);
nor U17693 (N_17693,N_17007,N_16974);
nor U17694 (N_17694,N_17041,N_16948);
nor U17695 (N_17695,N_16886,N_16814);
or U17696 (N_17696,N_17244,N_17083);
or U17697 (N_17697,N_16921,N_17059);
nor U17698 (N_17698,N_17319,N_16842);
xnor U17699 (N_17699,N_17369,N_16805);
nor U17700 (N_17700,N_17145,N_17342);
or U17701 (N_17701,N_16991,N_17292);
nor U17702 (N_17702,N_16997,N_16974);
nand U17703 (N_17703,N_16910,N_17314);
or U17704 (N_17704,N_17301,N_16919);
xnor U17705 (N_17705,N_16864,N_17314);
nand U17706 (N_17706,N_16881,N_16802);
nor U17707 (N_17707,N_17321,N_17152);
or U17708 (N_17708,N_17303,N_17150);
nand U17709 (N_17709,N_17199,N_17138);
or U17710 (N_17710,N_16947,N_17110);
and U17711 (N_17711,N_17304,N_17045);
xor U17712 (N_17712,N_16878,N_17185);
xor U17713 (N_17713,N_17055,N_17140);
or U17714 (N_17714,N_17098,N_16838);
and U17715 (N_17715,N_17131,N_16807);
and U17716 (N_17716,N_17099,N_16953);
or U17717 (N_17717,N_17352,N_17148);
and U17718 (N_17718,N_17122,N_17059);
xor U17719 (N_17719,N_17203,N_17004);
xor U17720 (N_17720,N_17273,N_17048);
and U17721 (N_17721,N_17060,N_16970);
or U17722 (N_17722,N_16845,N_17062);
or U17723 (N_17723,N_16828,N_17151);
xor U17724 (N_17724,N_17284,N_16916);
and U17725 (N_17725,N_16930,N_17360);
nand U17726 (N_17726,N_16919,N_16916);
or U17727 (N_17727,N_16952,N_17314);
nand U17728 (N_17728,N_17070,N_17259);
or U17729 (N_17729,N_16954,N_17150);
nand U17730 (N_17730,N_16862,N_17288);
or U17731 (N_17731,N_17184,N_17383);
nor U17732 (N_17732,N_17348,N_17167);
and U17733 (N_17733,N_17084,N_17357);
xnor U17734 (N_17734,N_17342,N_16940);
nand U17735 (N_17735,N_17090,N_16977);
nand U17736 (N_17736,N_17291,N_17148);
and U17737 (N_17737,N_16900,N_16851);
nor U17738 (N_17738,N_17141,N_17161);
xnor U17739 (N_17739,N_17161,N_16969);
nor U17740 (N_17740,N_17352,N_16805);
nand U17741 (N_17741,N_17173,N_17189);
nand U17742 (N_17742,N_16851,N_17238);
xnor U17743 (N_17743,N_16814,N_17084);
and U17744 (N_17744,N_16962,N_17111);
or U17745 (N_17745,N_17116,N_17395);
nand U17746 (N_17746,N_17161,N_16942);
xor U17747 (N_17747,N_16982,N_16889);
nor U17748 (N_17748,N_17332,N_16992);
nand U17749 (N_17749,N_16831,N_17091);
nand U17750 (N_17750,N_16933,N_16963);
xnor U17751 (N_17751,N_17158,N_17195);
nand U17752 (N_17752,N_16946,N_16982);
xor U17753 (N_17753,N_17055,N_16941);
nor U17754 (N_17754,N_16952,N_16885);
and U17755 (N_17755,N_17161,N_17360);
nand U17756 (N_17756,N_16963,N_17024);
and U17757 (N_17757,N_17250,N_17392);
nor U17758 (N_17758,N_17343,N_17204);
and U17759 (N_17759,N_17146,N_17057);
nor U17760 (N_17760,N_17129,N_16831);
nor U17761 (N_17761,N_16975,N_17362);
nor U17762 (N_17762,N_17198,N_17180);
nand U17763 (N_17763,N_17286,N_17003);
xnor U17764 (N_17764,N_17029,N_17106);
xor U17765 (N_17765,N_17249,N_16966);
or U17766 (N_17766,N_17289,N_16856);
nor U17767 (N_17767,N_17221,N_17210);
nor U17768 (N_17768,N_16862,N_16892);
or U17769 (N_17769,N_17396,N_16878);
nand U17770 (N_17770,N_16962,N_17359);
and U17771 (N_17771,N_16872,N_16907);
nand U17772 (N_17772,N_17112,N_17254);
or U17773 (N_17773,N_17022,N_16949);
nor U17774 (N_17774,N_17109,N_16896);
xnor U17775 (N_17775,N_17342,N_17286);
xor U17776 (N_17776,N_16821,N_17349);
and U17777 (N_17777,N_17277,N_16997);
nor U17778 (N_17778,N_17127,N_17335);
nor U17779 (N_17779,N_17335,N_16888);
or U17780 (N_17780,N_17397,N_17129);
or U17781 (N_17781,N_17051,N_17156);
xnor U17782 (N_17782,N_16978,N_17026);
nand U17783 (N_17783,N_17201,N_17396);
nand U17784 (N_17784,N_17394,N_17350);
nand U17785 (N_17785,N_17338,N_17053);
xnor U17786 (N_17786,N_17012,N_17026);
xor U17787 (N_17787,N_17333,N_16959);
and U17788 (N_17788,N_17038,N_17096);
and U17789 (N_17789,N_16928,N_17212);
or U17790 (N_17790,N_16892,N_16907);
nand U17791 (N_17791,N_17377,N_16867);
or U17792 (N_17792,N_17338,N_17206);
and U17793 (N_17793,N_16892,N_17009);
xor U17794 (N_17794,N_17279,N_16998);
nand U17795 (N_17795,N_17355,N_17246);
and U17796 (N_17796,N_16878,N_16816);
or U17797 (N_17797,N_17169,N_17237);
nand U17798 (N_17798,N_17140,N_17114);
nor U17799 (N_17799,N_17109,N_17273);
and U17800 (N_17800,N_17107,N_17196);
nor U17801 (N_17801,N_17326,N_17020);
xor U17802 (N_17802,N_17085,N_16988);
or U17803 (N_17803,N_16834,N_17095);
and U17804 (N_17804,N_17056,N_17161);
nand U17805 (N_17805,N_17050,N_16930);
nand U17806 (N_17806,N_17234,N_17077);
xor U17807 (N_17807,N_17016,N_17356);
xnor U17808 (N_17808,N_17176,N_17174);
nor U17809 (N_17809,N_17071,N_17183);
and U17810 (N_17810,N_16856,N_16915);
xnor U17811 (N_17811,N_16984,N_16975);
and U17812 (N_17812,N_16808,N_16814);
nand U17813 (N_17813,N_17225,N_17297);
nand U17814 (N_17814,N_17202,N_16967);
or U17815 (N_17815,N_17291,N_17228);
nor U17816 (N_17816,N_17108,N_17291);
and U17817 (N_17817,N_17009,N_16841);
nor U17818 (N_17818,N_16855,N_16983);
and U17819 (N_17819,N_17147,N_16950);
nor U17820 (N_17820,N_16865,N_17076);
and U17821 (N_17821,N_16820,N_16902);
nand U17822 (N_17822,N_17342,N_17076);
nand U17823 (N_17823,N_17162,N_17373);
nand U17824 (N_17824,N_16932,N_17233);
and U17825 (N_17825,N_16989,N_17347);
and U17826 (N_17826,N_17061,N_17165);
nand U17827 (N_17827,N_17344,N_16839);
xnor U17828 (N_17828,N_16839,N_17058);
or U17829 (N_17829,N_16879,N_17241);
nor U17830 (N_17830,N_17392,N_17193);
nor U17831 (N_17831,N_17259,N_16942);
nand U17832 (N_17832,N_17367,N_17124);
nor U17833 (N_17833,N_17043,N_17074);
nor U17834 (N_17834,N_16983,N_17015);
nand U17835 (N_17835,N_17147,N_16802);
xor U17836 (N_17836,N_16809,N_16986);
and U17837 (N_17837,N_17096,N_17023);
xor U17838 (N_17838,N_17084,N_17252);
or U17839 (N_17839,N_16912,N_17209);
and U17840 (N_17840,N_17224,N_17046);
nand U17841 (N_17841,N_16927,N_17379);
xor U17842 (N_17842,N_17131,N_16931);
xnor U17843 (N_17843,N_16848,N_16983);
xnor U17844 (N_17844,N_16833,N_17331);
nand U17845 (N_17845,N_17103,N_17382);
xnor U17846 (N_17846,N_17195,N_17388);
nor U17847 (N_17847,N_17079,N_17376);
nor U17848 (N_17848,N_16859,N_17145);
xor U17849 (N_17849,N_16943,N_17395);
nor U17850 (N_17850,N_16800,N_17300);
and U17851 (N_17851,N_16849,N_17170);
nand U17852 (N_17852,N_16810,N_16873);
or U17853 (N_17853,N_16949,N_17141);
xnor U17854 (N_17854,N_17289,N_17324);
or U17855 (N_17855,N_17105,N_17129);
xnor U17856 (N_17856,N_17108,N_17337);
and U17857 (N_17857,N_16910,N_17008);
nand U17858 (N_17858,N_17389,N_17323);
xnor U17859 (N_17859,N_16899,N_17213);
nand U17860 (N_17860,N_17185,N_16819);
xnor U17861 (N_17861,N_17169,N_17185);
and U17862 (N_17862,N_17154,N_16818);
xnor U17863 (N_17863,N_17224,N_17398);
nand U17864 (N_17864,N_17229,N_16940);
nand U17865 (N_17865,N_17185,N_17191);
or U17866 (N_17866,N_17101,N_17016);
nand U17867 (N_17867,N_17155,N_17324);
xnor U17868 (N_17868,N_17313,N_16982);
or U17869 (N_17869,N_17365,N_17092);
nor U17870 (N_17870,N_16944,N_17300);
nand U17871 (N_17871,N_17250,N_16930);
or U17872 (N_17872,N_17385,N_17250);
nor U17873 (N_17873,N_17344,N_16912);
and U17874 (N_17874,N_17172,N_17131);
xnor U17875 (N_17875,N_17281,N_16966);
nor U17876 (N_17876,N_17286,N_17185);
nand U17877 (N_17877,N_17336,N_17144);
nand U17878 (N_17878,N_17058,N_17253);
and U17879 (N_17879,N_16933,N_17032);
nor U17880 (N_17880,N_16953,N_16967);
nand U17881 (N_17881,N_16845,N_16890);
xnor U17882 (N_17882,N_17134,N_16903);
nand U17883 (N_17883,N_17129,N_16977);
or U17884 (N_17884,N_17012,N_17223);
nor U17885 (N_17885,N_17278,N_17141);
and U17886 (N_17886,N_17252,N_17130);
and U17887 (N_17887,N_17247,N_16941);
nand U17888 (N_17888,N_17038,N_17378);
or U17889 (N_17889,N_17097,N_16843);
nand U17890 (N_17890,N_17100,N_17116);
xor U17891 (N_17891,N_16936,N_17212);
nor U17892 (N_17892,N_17033,N_17055);
or U17893 (N_17893,N_17041,N_17066);
and U17894 (N_17894,N_17377,N_16881);
and U17895 (N_17895,N_17159,N_17055);
xnor U17896 (N_17896,N_17278,N_17338);
nand U17897 (N_17897,N_17290,N_17255);
xnor U17898 (N_17898,N_17240,N_17311);
nor U17899 (N_17899,N_17021,N_16843);
and U17900 (N_17900,N_17057,N_17108);
nor U17901 (N_17901,N_17022,N_16843);
nand U17902 (N_17902,N_16808,N_16816);
nand U17903 (N_17903,N_16859,N_17220);
and U17904 (N_17904,N_17093,N_16906);
nor U17905 (N_17905,N_17306,N_16833);
xnor U17906 (N_17906,N_17220,N_17312);
or U17907 (N_17907,N_17133,N_16902);
nand U17908 (N_17908,N_17136,N_16988);
xnor U17909 (N_17909,N_17021,N_16920);
nand U17910 (N_17910,N_17229,N_17151);
nor U17911 (N_17911,N_17050,N_16811);
or U17912 (N_17912,N_17141,N_17174);
nor U17913 (N_17913,N_17303,N_17183);
and U17914 (N_17914,N_17062,N_16932);
and U17915 (N_17915,N_17220,N_17081);
or U17916 (N_17916,N_17232,N_16893);
or U17917 (N_17917,N_17390,N_17162);
nand U17918 (N_17918,N_17111,N_17286);
and U17919 (N_17919,N_16959,N_16807);
nor U17920 (N_17920,N_16908,N_17314);
nor U17921 (N_17921,N_17222,N_17302);
and U17922 (N_17922,N_16974,N_17390);
nand U17923 (N_17923,N_17091,N_17262);
nor U17924 (N_17924,N_16837,N_16851);
xnor U17925 (N_17925,N_17214,N_17346);
or U17926 (N_17926,N_16842,N_17023);
nand U17927 (N_17927,N_17176,N_17132);
xor U17928 (N_17928,N_17234,N_17121);
or U17929 (N_17929,N_17331,N_17302);
nand U17930 (N_17930,N_16913,N_17165);
and U17931 (N_17931,N_16981,N_16900);
and U17932 (N_17932,N_17133,N_17120);
nor U17933 (N_17933,N_17049,N_17078);
and U17934 (N_17934,N_17267,N_17110);
nand U17935 (N_17935,N_16852,N_17056);
or U17936 (N_17936,N_16984,N_16863);
xnor U17937 (N_17937,N_17176,N_17013);
or U17938 (N_17938,N_16814,N_16810);
xnor U17939 (N_17939,N_16873,N_16930);
and U17940 (N_17940,N_17331,N_16873);
or U17941 (N_17941,N_17103,N_17106);
or U17942 (N_17942,N_16948,N_16917);
and U17943 (N_17943,N_17086,N_17323);
xor U17944 (N_17944,N_17111,N_17165);
nand U17945 (N_17945,N_17116,N_17270);
xnor U17946 (N_17946,N_17170,N_16833);
xor U17947 (N_17947,N_16983,N_17342);
and U17948 (N_17948,N_17047,N_16950);
xor U17949 (N_17949,N_17065,N_17127);
nand U17950 (N_17950,N_16807,N_17290);
or U17951 (N_17951,N_17375,N_16985);
xor U17952 (N_17952,N_17203,N_16985);
nand U17953 (N_17953,N_17345,N_17194);
xor U17954 (N_17954,N_17303,N_16871);
nand U17955 (N_17955,N_17287,N_16827);
nand U17956 (N_17956,N_17368,N_16871);
nor U17957 (N_17957,N_17250,N_16990);
or U17958 (N_17958,N_17280,N_16856);
nor U17959 (N_17959,N_17297,N_17041);
xor U17960 (N_17960,N_17211,N_17370);
or U17961 (N_17961,N_16892,N_17122);
or U17962 (N_17962,N_17396,N_16917);
xor U17963 (N_17963,N_17361,N_16921);
nor U17964 (N_17964,N_16893,N_17231);
nor U17965 (N_17965,N_17023,N_16860);
or U17966 (N_17966,N_16894,N_16917);
and U17967 (N_17967,N_16972,N_17396);
and U17968 (N_17968,N_16945,N_16906);
nand U17969 (N_17969,N_16960,N_17276);
or U17970 (N_17970,N_17061,N_17000);
xor U17971 (N_17971,N_17342,N_16986);
nor U17972 (N_17972,N_17177,N_17161);
and U17973 (N_17973,N_16821,N_16872);
nor U17974 (N_17974,N_17263,N_17198);
and U17975 (N_17975,N_16902,N_17319);
nand U17976 (N_17976,N_17266,N_17310);
or U17977 (N_17977,N_16874,N_16888);
nor U17978 (N_17978,N_17127,N_17310);
or U17979 (N_17979,N_17343,N_16977);
nor U17980 (N_17980,N_17294,N_16903);
nor U17981 (N_17981,N_17352,N_17389);
and U17982 (N_17982,N_17172,N_17343);
or U17983 (N_17983,N_16893,N_16953);
xnor U17984 (N_17984,N_16828,N_17310);
nand U17985 (N_17985,N_17122,N_17380);
nor U17986 (N_17986,N_17079,N_17283);
nand U17987 (N_17987,N_17301,N_16991);
and U17988 (N_17988,N_17147,N_16935);
xnor U17989 (N_17989,N_17255,N_16942);
and U17990 (N_17990,N_16840,N_16843);
nand U17991 (N_17991,N_17057,N_17353);
nand U17992 (N_17992,N_17201,N_16934);
xor U17993 (N_17993,N_16982,N_17383);
and U17994 (N_17994,N_17072,N_17369);
and U17995 (N_17995,N_17060,N_16826);
and U17996 (N_17996,N_17296,N_16943);
or U17997 (N_17997,N_17028,N_17353);
and U17998 (N_17998,N_17234,N_17034);
nand U17999 (N_17999,N_17265,N_17107);
nor U18000 (N_18000,N_17516,N_17507);
nand U18001 (N_18001,N_17476,N_17865);
xnor U18002 (N_18002,N_17475,N_17598);
or U18003 (N_18003,N_17977,N_17410);
nand U18004 (N_18004,N_17624,N_17660);
and U18005 (N_18005,N_17872,N_17726);
and U18006 (N_18006,N_17675,N_17674);
and U18007 (N_18007,N_17453,N_17945);
nand U18008 (N_18008,N_17537,N_17999);
nand U18009 (N_18009,N_17748,N_17727);
nand U18010 (N_18010,N_17502,N_17959);
or U18011 (N_18011,N_17582,N_17577);
nand U18012 (N_18012,N_17928,N_17721);
nor U18013 (N_18013,N_17784,N_17406);
nor U18014 (N_18014,N_17790,N_17432);
and U18015 (N_18015,N_17503,N_17665);
xnor U18016 (N_18016,N_17742,N_17631);
xor U18017 (N_18017,N_17500,N_17749);
nor U18018 (N_18018,N_17964,N_17879);
nand U18019 (N_18019,N_17894,N_17980);
nor U18020 (N_18020,N_17940,N_17454);
and U18021 (N_18021,N_17645,N_17847);
or U18022 (N_18022,N_17765,N_17963);
nor U18023 (N_18023,N_17540,N_17933);
nor U18024 (N_18024,N_17889,N_17524);
nor U18025 (N_18025,N_17857,N_17567);
nand U18026 (N_18026,N_17447,N_17490);
nor U18027 (N_18027,N_17952,N_17725);
nor U18028 (N_18028,N_17689,N_17844);
and U18029 (N_18029,N_17955,N_17758);
and U18030 (N_18030,N_17628,N_17691);
or U18031 (N_18031,N_17702,N_17536);
or U18032 (N_18032,N_17926,N_17442);
and U18033 (N_18033,N_17545,N_17415);
or U18034 (N_18034,N_17534,N_17757);
and U18035 (N_18035,N_17991,N_17616);
nor U18036 (N_18036,N_17734,N_17968);
and U18037 (N_18037,N_17767,N_17431);
and U18038 (N_18038,N_17600,N_17935);
nand U18039 (N_18039,N_17411,N_17547);
nand U18040 (N_18040,N_17508,N_17774);
xor U18041 (N_18041,N_17854,N_17615);
nor U18042 (N_18042,N_17944,N_17730);
nor U18043 (N_18043,N_17992,N_17778);
nand U18044 (N_18044,N_17750,N_17576);
or U18045 (N_18045,N_17412,N_17484);
and U18046 (N_18046,N_17528,N_17904);
and U18047 (N_18047,N_17762,N_17541);
or U18048 (N_18048,N_17895,N_17979);
or U18049 (N_18049,N_17648,N_17661);
or U18050 (N_18050,N_17998,N_17527);
or U18051 (N_18051,N_17829,N_17409);
and U18052 (N_18052,N_17662,N_17563);
xnor U18053 (N_18053,N_17664,N_17960);
nand U18054 (N_18054,N_17638,N_17679);
or U18055 (N_18055,N_17472,N_17728);
and U18056 (N_18056,N_17429,N_17636);
or U18057 (N_18057,N_17569,N_17986);
nor U18058 (N_18058,N_17818,N_17587);
and U18059 (N_18059,N_17592,N_17712);
or U18060 (N_18060,N_17623,N_17705);
nand U18061 (N_18061,N_17698,N_17511);
nor U18062 (N_18062,N_17512,N_17848);
xor U18063 (N_18063,N_17554,N_17753);
xnor U18064 (N_18064,N_17743,N_17850);
nand U18065 (N_18065,N_17449,N_17962);
xnor U18066 (N_18066,N_17918,N_17408);
and U18067 (N_18067,N_17611,N_17708);
nor U18068 (N_18068,N_17416,N_17744);
or U18069 (N_18069,N_17701,N_17514);
xnor U18070 (N_18070,N_17997,N_17806);
nand U18071 (N_18071,N_17450,N_17871);
nand U18072 (N_18072,N_17609,N_17629);
xor U18073 (N_18073,N_17506,N_17639);
nand U18074 (N_18074,N_17875,N_17771);
nand U18075 (N_18075,N_17413,N_17455);
and U18076 (N_18076,N_17703,N_17909);
nand U18077 (N_18077,N_17770,N_17633);
nand U18078 (N_18078,N_17535,N_17751);
xnor U18079 (N_18079,N_17678,N_17626);
or U18080 (N_18080,N_17884,N_17888);
or U18081 (N_18081,N_17988,N_17583);
xnor U18082 (N_18082,N_17612,N_17927);
nor U18083 (N_18083,N_17747,N_17613);
nand U18084 (N_18084,N_17594,N_17797);
nor U18085 (N_18085,N_17863,N_17597);
and U18086 (N_18086,N_17978,N_17816);
and U18087 (N_18087,N_17970,N_17634);
or U18088 (N_18088,N_17627,N_17720);
xor U18089 (N_18089,N_17619,N_17777);
xnor U18090 (N_18090,N_17669,N_17433);
and U18091 (N_18091,N_17448,N_17716);
xnor U18092 (N_18092,N_17779,N_17985);
and U18093 (N_18093,N_17425,N_17699);
nor U18094 (N_18094,N_17976,N_17843);
or U18095 (N_18095,N_17859,N_17658);
and U18096 (N_18096,N_17557,N_17805);
and U18097 (N_18097,N_17568,N_17795);
nand U18098 (N_18098,N_17921,N_17403);
nor U18099 (N_18099,N_17531,N_17407);
nor U18100 (N_18100,N_17562,N_17761);
xnor U18101 (N_18101,N_17853,N_17438);
xnor U18102 (N_18102,N_17915,N_17752);
nor U18103 (N_18103,N_17934,N_17707);
nand U18104 (N_18104,N_17617,N_17656);
or U18105 (N_18105,N_17693,N_17901);
nor U18106 (N_18106,N_17911,N_17719);
nand U18107 (N_18107,N_17841,N_17709);
and U18108 (N_18108,N_17852,N_17836);
nor U18109 (N_18109,N_17437,N_17897);
nor U18110 (N_18110,N_17845,N_17826);
xnor U18111 (N_18111,N_17780,N_17542);
nand U18112 (N_18112,N_17899,N_17929);
or U18113 (N_18113,N_17706,N_17644);
and U18114 (N_18114,N_17427,N_17526);
xnor U18115 (N_18115,N_17519,N_17440);
xnor U18116 (N_18116,N_17724,N_17942);
nand U18117 (N_18117,N_17849,N_17579);
and U18118 (N_18118,N_17653,N_17956);
or U18119 (N_18119,N_17457,N_17912);
nand U18120 (N_18120,N_17768,N_17808);
xnor U18121 (N_18121,N_17493,N_17824);
nor U18122 (N_18122,N_17763,N_17821);
and U18123 (N_18123,N_17870,N_17781);
and U18124 (N_18124,N_17866,N_17441);
and U18125 (N_18125,N_17867,N_17975);
xnor U18126 (N_18126,N_17922,N_17776);
nor U18127 (N_18127,N_17800,N_17681);
nand U18128 (N_18128,N_17489,N_17878);
nor U18129 (N_18129,N_17984,N_17657);
and U18130 (N_18130,N_17801,N_17769);
and U18131 (N_18131,N_17604,N_17682);
nand U18132 (N_18132,N_17522,N_17811);
xor U18133 (N_18133,N_17677,N_17939);
or U18134 (N_18134,N_17649,N_17428);
and U18135 (N_18135,N_17509,N_17903);
xor U18136 (N_18136,N_17467,N_17936);
nand U18137 (N_18137,N_17722,N_17443);
or U18138 (N_18138,N_17814,N_17640);
nor U18139 (N_18139,N_17543,N_17858);
and U18140 (N_18140,N_17614,N_17869);
nor U18141 (N_18141,N_17953,N_17802);
nor U18142 (N_18142,N_17607,N_17840);
or U18143 (N_18143,N_17823,N_17570);
and U18144 (N_18144,N_17710,N_17578);
or U18145 (N_18145,N_17573,N_17856);
xor U18146 (N_18146,N_17704,N_17605);
and U18147 (N_18147,N_17659,N_17813);
nand U18148 (N_18148,N_17591,N_17599);
or U18149 (N_18149,N_17555,N_17670);
and U18150 (N_18150,N_17550,N_17949);
nor U18151 (N_18151,N_17739,N_17561);
nand U18152 (N_18152,N_17825,N_17470);
and U18153 (N_18153,N_17828,N_17737);
nor U18154 (N_18154,N_17917,N_17495);
or U18155 (N_18155,N_17460,N_17520);
nor U18156 (N_18156,N_17958,N_17993);
and U18157 (N_18157,N_17864,N_17954);
or U18158 (N_18158,N_17606,N_17723);
and U18159 (N_18159,N_17401,N_17630);
and U18160 (N_18160,N_17715,N_17652);
nor U18161 (N_18161,N_17835,N_17913);
nand U18162 (N_18162,N_17951,N_17523);
nand U18163 (N_18163,N_17556,N_17434);
nand U18164 (N_18164,N_17581,N_17893);
and U18165 (N_18165,N_17480,N_17946);
and U18166 (N_18166,N_17685,N_17931);
or U18167 (N_18167,N_17435,N_17738);
or U18168 (N_18168,N_17792,N_17812);
xor U18169 (N_18169,N_17880,N_17444);
and U18170 (N_18170,N_17546,N_17566);
nand U18171 (N_18171,N_17994,N_17558);
nand U18172 (N_18172,N_17919,N_17745);
and U18173 (N_18173,N_17876,N_17593);
nand U18174 (N_18174,N_17430,N_17451);
nand U18175 (N_18175,N_17477,N_17683);
nor U18176 (N_18176,N_17474,N_17655);
nand U18177 (N_18177,N_17462,N_17647);
and U18178 (N_18178,N_17972,N_17798);
and U18179 (N_18179,N_17982,N_17833);
xnor U18180 (N_18180,N_17673,N_17422);
nand U18181 (N_18181,N_17908,N_17873);
nand U18182 (N_18182,N_17862,N_17874);
nor U18183 (N_18183,N_17799,N_17552);
nor U18184 (N_18184,N_17646,N_17436);
xor U18185 (N_18185,N_17713,N_17957);
or U18186 (N_18186,N_17608,N_17832);
nor U18187 (N_18187,N_17783,N_17896);
nor U18188 (N_18188,N_17494,N_17941);
nand U18189 (N_18189,N_17654,N_17855);
nor U18190 (N_18190,N_17481,N_17690);
or U18191 (N_18191,N_17900,N_17989);
nand U18192 (N_18192,N_17834,N_17445);
nand U18193 (N_18193,N_17817,N_17610);
nand U18194 (N_18194,N_17948,N_17529);
nand U18195 (N_18195,N_17595,N_17830);
nor U18196 (N_18196,N_17794,N_17544);
and U18197 (N_18197,N_17603,N_17461);
nand U18198 (N_18198,N_17478,N_17589);
nand U18199 (N_18199,N_17414,N_17981);
nand U18200 (N_18200,N_17618,N_17990);
xnor U18201 (N_18201,N_17575,N_17965);
or U18202 (N_18202,N_17505,N_17551);
or U18203 (N_18203,N_17787,N_17882);
nand U18204 (N_18204,N_17565,N_17471);
nand U18205 (N_18205,N_17404,N_17525);
and U18206 (N_18206,N_17861,N_17521);
or U18207 (N_18207,N_17733,N_17424);
and U18208 (N_18208,N_17729,N_17692);
nand U18209 (N_18209,N_17796,N_17786);
or U18210 (N_18210,N_17731,N_17572);
nand U18211 (N_18211,N_17877,N_17559);
xor U18212 (N_18212,N_17684,N_17446);
and U18213 (N_18213,N_17418,N_17791);
xnor U18214 (N_18214,N_17898,N_17632);
and U18215 (N_18215,N_17686,N_17420);
and U18216 (N_18216,N_17687,N_17635);
and U18217 (N_18217,N_17642,N_17688);
nand U18218 (N_18218,N_17482,N_17532);
nor U18219 (N_18219,N_17421,N_17517);
nand U18220 (N_18220,N_17868,N_17851);
and U18221 (N_18221,N_17548,N_17756);
xnor U18222 (N_18222,N_17700,N_17961);
nor U18223 (N_18223,N_17755,N_17696);
nor U18224 (N_18224,N_17810,N_17417);
or U18225 (N_18225,N_17590,N_17969);
xnor U18226 (N_18226,N_17746,N_17510);
and U18227 (N_18227,N_17458,N_17549);
nand U18228 (N_18228,N_17667,N_17571);
and U18229 (N_18229,N_17892,N_17637);
and U18230 (N_18230,N_17464,N_17759);
nand U18231 (N_18231,N_17533,N_17574);
or U18232 (N_18232,N_17819,N_17663);
xnor U18233 (N_18233,N_17846,N_17672);
nor U18234 (N_18234,N_17973,N_17782);
nand U18235 (N_18235,N_17650,N_17515);
and U18236 (N_18236,N_17966,N_17905);
and U18237 (N_18237,N_17772,N_17501);
or U18238 (N_18238,N_17641,N_17620);
nor U18239 (N_18239,N_17914,N_17539);
xnor U18240 (N_18240,N_17479,N_17764);
xnor U18241 (N_18241,N_17459,N_17804);
xor U18242 (N_18242,N_17820,N_17694);
xor U18243 (N_18243,N_17775,N_17584);
nor U18244 (N_18244,N_17596,N_17995);
nand U18245 (N_18245,N_17465,N_17967);
or U18246 (N_18246,N_17585,N_17932);
and U18247 (N_18247,N_17697,N_17499);
and U18248 (N_18248,N_17711,N_17492);
or U18249 (N_18249,N_17831,N_17601);
and U18250 (N_18250,N_17773,N_17930);
xnor U18251 (N_18251,N_17789,N_17793);
and U18252 (N_18252,N_17983,N_17580);
xnor U18253 (N_18253,N_17837,N_17842);
nand U18254 (N_18254,N_17890,N_17827);
or U18255 (N_18255,N_17741,N_17560);
or U18256 (N_18256,N_17668,N_17419);
nor U18257 (N_18257,N_17463,N_17402);
nand U18258 (N_18258,N_17518,N_17910);
nor U18259 (N_18259,N_17947,N_17538);
xor U18260 (N_18260,N_17987,N_17902);
and U18261 (N_18261,N_17695,N_17671);
xnor U18262 (N_18262,N_17602,N_17736);
xor U18263 (N_18263,N_17588,N_17924);
nor U18264 (N_18264,N_17803,N_17643);
and U18265 (N_18265,N_17513,N_17740);
and U18266 (N_18266,N_17885,N_17714);
or U18267 (N_18267,N_17881,N_17496);
or U18268 (N_18268,N_17766,N_17439);
nand U18269 (N_18269,N_17625,N_17485);
and U18270 (N_18270,N_17717,N_17760);
and U18271 (N_18271,N_17860,N_17907);
nor U18272 (N_18272,N_17920,N_17468);
and U18273 (N_18273,N_17487,N_17788);
nor U18274 (N_18274,N_17950,N_17891);
and U18275 (N_18275,N_17974,N_17469);
xor U18276 (N_18276,N_17473,N_17666);
xnor U18277 (N_18277,N_17456,N_17497);
xnor U18278 (N_18278,N_17400,N_17807);
nand U18279 (N_18279,N_17622,N_17676);
nand U18280 (N_18280,N_17996,N_17906);
nor U18281 (N_18281,N_17916,N_17405);
and U18282 (N_18282,N_17785,N_17839);
nor U18283 (N_18283,N_17938,N_17564);
nor U18284 (N_18284,N_17426,N_17466);
xor U18285 (N_18285,N_17735,N_17586);
nand U18286 (N_18286,N_17423,N_17754);
or U18287 (N_18287,N_17491,N_17651);
xor U18288 (N_18288,N_17937,N_17498);
or U18289 (N_18289,N_17732,N_17553);
and U18290 (N_18290,N_17483,N_17971);
and U18291 (N_18291,N_17718,N_17504);
or U18292 (N_18292,N_17923,N_17838);
or U18293 (N_18293,N_17925,N_17530);
or U18294 (N_18294,N_17680,N_17486);
or U18295 (N_18295,N_17883,N_17887);
xnor U18296 (N_18296,N_17815,N_17809);
nand U18297 (N_18297,N_17488,N_17621);
xnor U18298 (N_18298,N_17943,N_17452);
nor U18299 (N_18299,N_17886,N_17822);
xor U18300 (N_18300,N_17893,N_17813);
or U18301 (N_18301,N_17968,N_17853);
xnor U18302 (N_18302,N_17662,N_17626);
or U18303 (N_18303,N_17528,N_17923);
or U18304 (N_18304,N_17962,N_17556);
nor U18305 (N_18305,N_17945,N_17498);
nand U18306 (N_18306,N_17527,N_17813);
nand U18307 (N_18307,N_17834,N_17947);
or U18308 (N_18308,N_17989,N_17404);
xnor U18309 (N_18309,N_17728,N_17521);
nand U18310 (N_18310,N_17744,N_17954);
nand U18311 (N_18311,N_17401,N_17493);
nor U18312 (N_18312,N_17428,N_17949);
nor U18313 (N_18313,N_17461,N_17596);
or U18314 (N_18314,N_17566,N_17984);
and U18315 (N_18315,N_17642,N_17928);
nor U18316 (N_18316,N_17768,N_17754);
and U18317 (N_18317,N_17822,N_17988);
or U18318 (N_18318,N_17543,N_17673);
or U18319 (N_18319,N_17859,N_17459);
xnor U18320 (N_18320,N_17611,N_17499);
nand U18321 (N_18321,N_17628,N_17895);
and U18322 (N_18322,N_17679,N_17839);
nand U18323 (N_18323,N_17944,N_17579);
or U18324 (N_18324,N_17560,N_17480);
and U18325 (N_18325,N_17472,N_17400);
xnor U18326 (N_18326,N_17664,N_17478);
nand U18327 (N_18327,N_17676,N_17824);
or U18328 (N_18328,N_17528,N_17619);
xnor U18329 (N_18329,N_17419,N_17496);
xnor U18330 (N_18330,N_17999,N_17548);
nor U18331 (N_18331,N_17780,N_17650);
xnor U18332 (N_18332,N_17954,N_17679);
or U18333 (N_18333,N_17601,N_17857);
and U18334 (N_18334,N_17762,N_17548);
and U18335 (N_18335,N_17608,N_17723);
and U18336 (N_18336,N_17883,N_17510);
and U18337 (N_18337,N_17636,N_17678);
and U18338 (N_18338,N_17437,N_17849);
nor U18339 (N_18339,N_17409,N_17715);
or U18340 (N_18340,N_17441,N_17693);
nand U18341 (N_18341,N_17561,N_17907);
nand U18342 (N_18342,N_17751,N_17410);
or U18343 (N_18343,N_17954,N_17536);
nand U18344 (N_18344,N_17825,N_17923);
or U18345 (N_18345,N_17675,N_17827);
xnor U18346 (N_18346,N_17644,N_17726);
or U18347 (N_18347,N_17872,N_17730);
or U18348 (N_18348,N_17438,N_17563);
xor U18349 (N_18349,N_17444,N_17695);
xor U18350 (N_18350,N_17585,N_17991);
nand U18351 (N_18351,N_17463,N_17720);
or U18352 (N_18352,N_17611,N_17732);
nand U18353 (N_18353,N_17667,N_17681);
xnor U18354 (N_18354,N_17949,N_17680);
xor U18355 (N_18355,N_17606,N_17461);
nand U18356 (N_18356,N_17594,N_17538);
and U18357 (N_18357,N_17424,N_17726);
xor U18358 (N_18358,N_17717,N_17618);
xor U18359 (N_18359,N_17550,N_17945);
xor U18360 (N_18360,N_17591,N_17733);
or U18361 (N_18361,N_17784,N_17667);
nor U18362 (N_18362,N_17505,N_17501);
and U18363 (N_18363,N_17909,N_17881);
or U18364 (N_18364,N_17694,N_17763);
nor U18365 (N_18365,N_17610,N_17615);
nand U18366 (N_18366,N_17705,N_17942);
nor U18367 (N_18367,N_17841,N_17575);
and U18368 (N_18368,N_17782,N_17459);
and U18369 (N_18369,N_17725,N_17567);
nor U18370 (N_18370,N_17819,N_17588);
or U18371 (N_18371,N_17671,N_17751);
or U18372 (N_18372,N_17576,N_17456);
and U18373 (N_18373,N_17817,N_17949);
or U18374 (N_18374,N_17834,N_17524);
or U18375 (N_18375,N_17644,N_17873);
xnor U18376 (N_18376,N_17993,N_17419);
and U18377 (N_18377,N_17971,N_17723);
nor U18378 (N_18378,N_17843,N_17644);
nor U18379 (N_18379,N_17594,N_17713);
nand U18380 (N_18380,N_17582,N_17477);
or U18381 (N_18381,N_17916,N_17582);
nand U18382 (N_18382,N_17530,N_17797);
nand U18383 (N_18383,N_17856,N_17725);
or U18384 (N_18384,N_17857,N_17725);
nand U18385 (N_18385,N_17465,N_17999);
xnor U18386 (N_18386,N_17758,N_17530);
or U18387 (N_18387,N_17923,N_17964);
xnor U18388 (N_18388,N_17532,N_17989);
and U18389 (N_18389,N_17519,N_17583);
nand U18390 (N_18390,N_17847,N_17532);
nor U18391 (N_18391,N_17609,N_17540);
or U18392 (N_18392,N_17989,N_17668);
and U18393 (N_18393,N_17743,N_17443);
nand U18394 (N_18394,N_17470,N_17803);
and U18395 (N_18395,N_17786,N_17614);
nor U18396 (N_18396,N_17562,N_17421);
nand U18397 (N_18397,N_17412,N_17492);
or U18398 (N_18398,N_17746,N_17452);
and U18399 (N_18399,N_17605,N_17923);
xnor U18400 (N_18400,N_17911,N_17797);
and U18401 (N_18401,N_17852,N_17861);
and U18402 (N_18402,N_17475,N_17972);
or U18403 (N_18403,N_17856,N_17749);
xnor U18404 (N_18404,N_17696,N_17682);
nand U18405 (N_18405,N_17816,N_17832);
and U18406 (N_18406,N_17951,N_17790);
nor U18407 (N_18407,N_17576,N_17978);
or U18408 (N_18408,N_17594,N_17613);
nand U18409 (N_18409,N_17936,N_17511);
nand U18410 (N_18410,N_17856,N_17884);
or U18411 (N_18411,N_17946,N_17897);
xor U18412 (N_18412,N_17443,N_17698);
or U18413 (N_18413,N_17672,N_17488);
xor U18414 (N_18414,N_17542,N_17920);
or U18415 (N_18415,N_17908,N_17713);
nand U18416 (N_18416,N_17851,N_17717);
nor U18417 (N_18417,N_17832,N_17763);
xor U18418 (N_18418,N_17713,N_17941);
xnor U18419 (N_18419,N_17402,N_17533);
and U18420 (N_18420,N_17584,N_17671);
or U18421 (N_18421,N_17405,N_17983);
nor U18422 (N_18422,N_17515,N_17585);
xor U18423 (N_18423,N_17766,N_17789);
or U18424 (N_18424,N_17668,N_17821);
nand U18425 (N_18425,N_17493,N_17761);
and U18426 (N_18426,N_17913,N_17615);
or U18427 (N_18427,N_17887,N_17637);
and U18428 (N_18428,N_17757,N_17771);
xnor U18429 (N_18429,N_17872,N_17793);
nor U18430 (N_18430,N_17494,N_17444);
nor U18431 (N_18431,N_17615,N_17813);
xor U18432 (N_18432,N_17595,N_17585);
nor U18433 (N_18433,N_17771,N_17476);
xnor U18434 (N_18434,N_17909,N_17603);
or U18435 (N_18435,N_17771,N_17745);
or U18436 (N_18436,N_17442,N_17557);
nand U18437 (N_18437,N_17454,N_17452);
xor U18438 (N_18438,N_17923,N_17960);
or U18439 (N_18439,N_17471,N_17608);
nand U18440 (N_18440,N_17922,N_17732);
xnor U18441 (N_18441,N_17410,N_17666);
xnor U18442 (N_18442,N_17673,N_17702);
and U18443 (N_18443,N_17907,N_17969);
nor U18444 (N_18444,N_17651,N_17588);
nand U18445 (N_18445,N_17561,N_17609);
nand U18446 (N_18446,N_17518,N_17951);
or U18447 (N_18447,N_17544,N_17935);
xor U18448 (N_18448,N_17581,N_17639);
xor U18449 (N_18449,N_17954,N_17669);
nor U18450 (N_18450,N_17721,N_17430);
nor U18451 (N_18451,N_17586,N_17606);
nand U18452 (N_18452,N_17429,N_17947);
or U18453 (N_18453,N_17699,N_17456);
nand U18454 (N_18454,N_17845,N_17971);
nor U18455 (N_18455,N_17867,N_17449);
and U18456 (N_18456,N_17892,N_17734);
or U18457 (N_18457,N_17747,N_17546);
nand U18458 (N_18458,N_17421,N_17670);
nor U18459 (N_18459,N_17707,N_17600);
nand U18460 (N_18460,N_17434,N_17707);
or U18461 (N_18461,N_17932,N_17936);
or U18462 (N_18462,N_17642,N_17795);
nor U18463 (N_18463,N_17926,N_17776);
xor U18464 (N_18464,N_17423,N_17903);
nor U18465 (N_18465,N_17605,N_17500);
nand U18466 (N_18466,N_17624,N_17502);
and U18467 (N_18467,N_17549,N_17976);
nor U18468 (N_18468,N_17798,N_17893);
and U18469 (N_18469,N_17724,N_17838);
nor U18470 (N_18470,N_17734,N_17940);
nor U18471 (N_18471,N_17433,N_17815);
or U18472 (N_18472,N_17456,N_17981);
xor U18473 (N_18473,N_17761,N_17821);
nor U18474 (N_18474,N_17783,N_17472);
nand U18475 (N_18475,N_17998,N_17701);
nand U18476 (N_18476,N_17779,N_17899);
nor U18477 (N_18477,N_17436,N_17939);
and U18478 (N_18478,N_17495,N_17812);
nor U18479 (N_18479,N_17707,N_17566);
xnor U18480 (N_18480,N_17898,N_17825);
or U18481 (N_18481,N_17743,N_17505);
nor U18482 (N_18482,N_17508,N_17438);
nor U18483 (N_18483,N_17616,N_17800);
and U18484 (N_18484,N_17765,N_17899);
nor U18485 (N_18485,N_17520,N_17679);
xnor U18486 (N_18486,N_17435,N_17437);
nor U18487 (N_18487,N_17744,N_17875);
or U18488 (N_18488,N_17593,N_17461);
nor U18489 (N_18489,N_17425,N_17620);
and U18490 (N_18490,N_17972,N_17820);
nor U18491 (N_18491,N_17576,N_17696);
nand U18492 (N_18492,N_17709,N_17877);
nor U18493 (N_18493,N_17633,N_17747);
or U18494 (N_18494,N_17482,N_17814);
nand U18495 (N_18495,N_17982,N_17717);
nand U18496 (N_18496,N_17435,N_17916);
and U18497 (N_18497,N_17832,N_17858);
xor U18498 (N_18498,N_17860,N_17680);
nand U18499 (N_18499,N_17486,N_17748);
nand U18500 (N_18500,N_17746,N_17451);
nor U18501 (N_18501,N_17625,N_17586);
and U18502 (N_18502,N_17684,N_17852);
xnor U18503 (N_18503,N_17971,N_17599);
xor U18504 (N_18504,N_17800,N_17906);
or U18505 (N_18505,N_17980,N_17752);
xnor U18506 (N_18506,N_17739,N_17782);
or U18507 (N_18507,N_17644,N_17862);
or U18508 (N_18508,N_17633,N_17446);
xor U18509 (N_18509,N_17678,N_17892);
nor U18510 (N_18510,N_17795,N_17645);
or U18511 (N_18511,N_17899,N_17872);
nor U18512 (N_18512,N_17929,N_17543);
and U18513 (N_18513,N_17649,N_17699);
or U18514 (N_18514,N_17883,N_17590);
nand U18515 (N_18515,N_17445,N_17956);
nor U18516 (N_18516,N_17679,N_17662);
nor U18517 (N_18517,N_17481,N_17484);
xor U18518 (N_18518,N_17673,N_17712);
and U18519 (N_18519,N_17966,N_17723);
nor U18520 (N_18520,N_17518,N_17425);
xnor U18521 (N_18521,N_17469,N_17500);
and U18522 (N_18522,N_17448,N_17702);
nor U18523 (N_18523,N_17676,N_17718);
nand U18524 (N_18524,N_17515,N_17963);
nor U18525 (N_18525,N_17803,N_17558);
xor U18526 (N_18526,N_17569,N_17414);
nand U18527 (N_18527,N_17676,N_17576);
and U18528 (N_18528,N_17515,N_17420);
nand U18529 (N_18529,N_17761,N_17679);
or U18530 (N_18530,N_17946,N_17756);
or U18531 (N_18531,N_17736,N_17729);
xnor U18532 (N_18532,N_17836,N_17915);
nand U18533 (N_18533,N_17730,N_17594);
and U18534 (N_18534,N_17768,N_17954);
and U18535 (N_18535,N_17561,N_17689);
or U18536 (N_18536,N_17742,N_17489);
and U18537 (N_18537,N_17520,N_17618);
and U18538 (N_18538,N_17745,N_17615);
nand U18539 (N_18539,N_17876,N_17620);
nor U18540 (N_18540,N_17710,N_17945);
nand U18541 (N_18541,N_17879,N_17774);
nor U18542 (N_18542,N_17482,N_17563);
nand U18543 (N_18543,N_17480,N_17651);
nor U18544 (N_18544,N_17550,N_17950);
or U18545 (N_18545,N_17957,N_17424);
xor U18546 (N_18546,N_17996,N_17781);
xnor U18547 (N_18547,N_17787,N_17411);
nand U18548 (N_18548,N_17908,N_17483);
nor U18549 (N_18549,N_17994,N_17587);
nor U18550 (N_18550,N_17906,N_17508);
xor U18551 (N_18551,N_17523,N_17428);
xor U18552 (N_18552,N_17831,N_17676);
xnor U18553 (N_18553,N_17499,N_17770);
nor U18554 (N_18554,N_17727,N_17791);
and U18555 (N_18555,N_17671,N_17852);
xnor U18556 (N_18556,N_17598,N_17622);
and U18557 (N_18557,N_17653,N_17734);
xnor U18558 (N_18558,N_17588,N_17943);
and U18559 (N_18559,N_17925,N_17613);
nand U18560 (N_18560,N_17546,N_17642);
or U18561 (N_18561,N_17618,N_17595);
nor U18562 (N_18562,N_17954,N_17970);
nand U18563 (N_18563,N_17787,N_17881);
and U18564 (N_18564,N_17453,N_17527);
nor U18565 (N_18565,N_17751,N_17824);
nand U18566 (N_18566,N_17714,N_17783);
and U18567 (N_18567,N_17886,N_17415);
xor U18568 (N_18568,N_17793,N_17981);
nor U18569 (N_18569,N_17898,N_17922);
nor U18570 (N_18570,N_17648,N_17616);
xor U18571 (N_18571,N_17579,N_17895);
and U18572 (N_18572,N_17992,N_17876);
and U18573 (N_18573,N_17699,N_17752);
nor U18574 (N_18574,N_17832,N_17782);
xnor U18575 (N_18575,N_17924,N_17832);
or U18576 (N_18576,N_17987,N_17503);
and U18577 (N_18577,N_17974,N_17873);
xnor U18578 (N_18578,N_17790,N_17729);
nand U18579 (N_18579,N_17965,N_17571);
and U18580 (N_18580,N_17571,N_17526);
or U18581 (N_18581,N_17982,N_17899);
xnor U18582 (N_18582,N_17937,N_17921);
or U18583 (N_18583,N_17426,N_17626);
or U18584 (N_18584,N_17794,N_17866);
xnor U18585 (N_18585,N_17624,N_17629);
nand U18586 (N_18586,N_17435,N_17403);
nand U18587 (N_18587,N_17431,N_17576);
nor U18588 (N_18588,N_17923,N_17913);
nand U18589 (N_18589,N_17480,N_17511);
and U18590 (N_18590,N_17670,N_17771);
nor U18591 (N_18591,N_17625,N_17596);
nor U18592 (N_18592,N_17543,N_17851);
nand U18593 (N_18593,N_17621,N_17951);
nor U18594 (N_18594,N_17426,N_17547);
and U18595 (N_18595,N_17547,N_17903);
nand U18596 (N_18596,N_17617,N_17699);
or U18597 (N_18597,N_17680,N_17540);
xnor U18598 (N_18598,N_17755,N_17524);
and U18599 (N_18599,N_17525,N_17724);
nor U18600 (N_18600,N_18499,N_18010);
or U18601 (N_18601,N_18572,N_18035);
xor U18602 (N_18602,N_18279,N_18204);
xor U18603 (N_18603,N_18305,N_18262);
and U18604 (N_18604,N_18354,N_18285);
xor U18605 (N_18605,N_18199,N_18238);
or U18606 (N_18606,N_18104,N_18289);
nor U18607 (N_18607,N_18290,N_18312);
and U18608 (N_18608,N_18527,N_18464);
nor U18609 (N_18609,N_18007,N_18114);
nand U18610 (N_18610,N_18457,N_18268);
xor U18611 (N_18611,N_18095,N_18599);
nor U18612 (N_18612,N_18167,N_18232);
xnor U18613 (N_18613,N_18040,N_18200);
xnor U18614 (N_18614,N_18433,N_18297);
or U18615 (N_18615,N_18001,N_18031);
or U18616 (N_18616,N_18447,N_18544);
xor U18617 (N_18617,N_18539,N_18397);
and U18618 (N_18618,N_18392,N_18582);
xor U18619 (N_18619,N_18049,N_18584);
nand U18620 (N_18620,N_18191,N_18381);
and U18621 (N_18621,N_18281,N_18562);
and U18622 (N_18622,N_18355,N_18249);
nand U18623 (N_18623,N_18023,N_18261);
and U18624 (N_18624,N_18195,N_18319);
nand U18625 (N_18625,N_18549,N_18436);
xnor U18626 (N_18626,N_18346,N_18330);
nor U18627 (N_18627,N_18583,N_18428);
or U18628 (N_18628,N_18387,N_18175);
nand U18629 (N_18629,N_18404,N_18231);
nand U18630 (N_18630,N_18022,N_18301);
xor U18631 (N_18631,N_18034,N_18111);
nand U18632 (N_18632,N_18203,N_18337);
and U18633 (N_18633,N_18278,N_18431);
and U18634 (N_18634,N_18252,N_18536);
nor U18635 (N_18635,N_18395,N_18521);
or U18636 (N_18636,N_18359,N_18465);
and U18637 (N_18637,N_18157,N_18540);
nand U18638 (N_18638,N_18481,N_18103);
or U18639 (N_18639,N_18304,N_18089);
xnor U18640 (N_18640,N_18420,N_18245);
or U18641 (N_18641,N_18258,N_18011);
nor U18642 (N_18642,N_18505,N_18283);
nand U18643 (N_18643,N_18240,N_18223);
and U18644 (N_18644,N_18339,N_18019);
xor U18645 (N_18645,N_18077,N_18419);
and U18646 (N_18646,N_18506,N_18026);
nor U18647 (N_18647,N_18538,N_18320);
or U18648 (N_18648,N_18323,N_18058);
or U18649 (N_18649,N_18250,N_18568);
or U18650 (N_18650,N_18020,N_18518);
and U18651 (N_18651,N_18550,N_18291);
or U18652 (N_18652,N_18298,N_18528);
nor U18653 (N_18653,N_18585,N_18327);
nand U18654 (N_18654,N_18311,N_18124);
and U18655 (N_18655,N_18091,N_18567);
xnor U18656 (N_18656,N_18452,N_18213);
nor U18657 (N_18657,N_18147,N_18293);
xnor U18658 (N_18658,N_18561,N_18377);
nand U18659 (N_18659,N_18318,N_18141);
or U18660 (N_18660,N_18149,N_18072);
xor U18661 (N_18661,N_18070,N_18229);
and U18662 (N_18662,N_18079,N_18125);
and U18663 (N_18663,N_18186,N_18430);
nand U18664 (N_18664,N_18492,N_18423);
or U18665 (N_18665,N_18033,N_18140);
or U18666 (N_18666,N_18520,N_18593);
nand U18667 (N_18667,N_18483,N_18029);
xnor U18668 (N_18668,N_18398,N_18371);
xnor U18669 (N_18669,N_18047,N_18315);
or U18670 (N_18670,N_18313,N_18542);
nor U18671 (N_18671,N_18519,N_18565);
nand U18672 (N_18672,N_18106,N_18440);
nand U18673 (N_18673,N_18090,N_18597);
nand U18674 (N_18674,N_18185,N_18437);
xnor U18675 (N_18675,N_18166,N_18324);
nor U18676 (N_18676,N_18037,N_18448);
nand U18677 (N_18677,N_18099,N_18449);
and U18678 (N_18678,N_18131,N_18129);
nor U18679 (N_18679,N_18073,N_18331);
and U18680 (N_18680,N_18165,N_18490);
nor U18681 (N_18681,N_18206,N_18391);
or U18682 (N_18682,N_18112,N_18343);
and U18683 (N_18683,N_18458,N_18406);
nand U18684 (N_18684,N_18155,N_18260);
or U18685 (N_18685,N_18142,N_18135);
xnor U18686 (N_18686,N_18153,N_18389);
nor U18687 (N_18687,N_18393,N_18571);
nor U18688 (N_18688,N_18021,N_18588);
xor U18689 (N_18689,N_18286,N_18531);
xor U18690 (N_18690,N_18533,N_18515);
and U18691 (N_18691,N_18052,N_18192);
xnor U18692 (N_18692,N_18065,N_18445);
nand U18693 (N_18693,N_18592,N_18000);
nor U18694 (N_18694,N_18030,N_18338);
nand U18695 (N_18695,N_18508,N_18004);
or U18696 (N_18696,N_18470,N_18154);
or U18697 (N_18697,N_18352,N_18274);
nand U18698 (N_18698,N_18081,N_18367);
or U18699 (N_18699,N_18182,N_18161);
and U18700 (N_18700,N_18267,N_18045);
nor U18701 (N_18701,N_18292,N_18187);
or U18702 (N_18702,N_18378,N_18317);
and U18703 (N_18703,N_18284,N_18425);
xor U18704 (N_18704,N_18384,N_18068);
nor U18705 (N_18705,N_18064,N_18224);
nor U18706 (N_18706,N_18435,N_18221);
xnor U18707 (N_18707,N_18478,N_18265);
nor U18708 (N_18708,N_18108,N_18422);
nor U18709 (N_18709,N_18294,N_18369);
and U18710 (N_18710,N_18054,N_18085);
and U18711 (N_18711,N_18078,N_18136);
or U18712 (N_18712,N_18014,N_18546);
nor U18713 (N_18713,N_18442,N_18247);
and U18714 (N_18714,N_18362,N_18342);
nor U18715 (N_18715,N_18174,N_18248);
nand U18716 (N_18716,N_18237,N_18418);
nand U18717 (N_18717,N_18375,N_18368);
nand U18718 (N_18718,N_18137,N_18380);
or U18719 (N_18719,N_18590,N_18178);
and U18720 (N_18720,N_18408,N_18488);
or U18721 (N_18721,N_18122,N_18444);
or U18722 (N_18722,N_18183,N_18042);
xor U18723 (N_18723,N_18471,N_18441);
xnor U18724 (N_18724,N_18390,N_18236);
and U18725 (N_18725,N_18512,N_18446);
xor U18726 (N_18726,N_18353,N_18476);
nand U18727 (N_18727,N_18553,N_18427);
nand U18728 (N_18728,N_18219,N_18024);
nand U18729 (N_18729,N_18205,N_18190);
and U18730 (N_18730,N_18098,N_18494);
and U18731 (N_18731,N_18578,N_18316);
or U18732 (N_18732,N_18573,N_18207);
or U18733 (N_18733,N_18295,N_18489);
or U18734 (N_18734,N_18576,N_18027);
or U18735 (N_18735,N_18579,N_18351);
nor U18736 (N_18736,N_18028,N_18556);
xor U18737 (N_18737,N_18156,N_18438);
or U18738 (N_18738,N_18580,N_18560);
nor U18739 (N_18739,N_18211,N_18171);
nand U18740 (N_18740,N_18475,N_18414);
xnor U18741 (N_18741,N_18176,N_18009);
and U18742 (N_18742,N_18517,N_18598);
nor U18743 (N_18743,N_18075,N_18459);
or U18744 (N_18744,N_18242,N_18253);
or U18745 (N_18745,N_18363,N_18409);
and U18746 (N_18746,N_18288,N_18310);
and U18747 (N_18747,N_18039,N_18596);
or U18748 (N_18748,N_18256,N_18116);
or U18749 (N_18749,N_18497,N_18059);
nor U18750 (N_18750,N_18455,N_18480);
or U18751 (N_18751,N_18210,N_18595);
and U18752 (N_18752,N_18227,N_18328);
nor U18753 (N_18753,N_18373,N_18524);
nor U18754 (N_18754,N_18087,N_18074);
nand U18755 (N_18755,N_18463,N_18209);
xor U18756 (N_18756,N_18016,N_18434);
or U18757 (N_18757,N_18566,N_18426);
nand U18758 (N_18758,N_18127,N_18314);
xor U18759 (N_18759,N_18080,N_18255);
nand U18760 (N_18760,N_18547,N_18117);
or U18761 (N_18761,N_18100,N_18530);
xor U18762 (N_18762,N_18118,N_18225);
nand U18763 (N_18763,N_18350,N_18143);
or U18764 (N_18764,N_18300,N_18145);
nor U18765 (N_18765,N_18244,N_18275);
nand U18766 (N_18766,N_18060,N_18150);
nor U18767 (N_18767,N_18370,N_18541);
nor U18768 (N_18768,N_18329,N_18469);
nor U18769 (N_18769,N_18144,N_18102);
or U18770 (N_18770,N_18364,N_18454);
nor U18771 (N_18771,N_18076,N_18243);
xor U18772 (N_18772,N_18554,N_18152);
nand U18773 (N_18773,N_18482,N_18333);
xor U18774 (N_18774,N_18197,N_18461);
nand U18775 (N_18775,N_18516,N_18336);
or U18776 (N_18776,N_18208,N_18133);
xor U18777 (N_18777,N_18510,N_18462);
and U18778 (N_18778,N_18189,N_18372);
nor U18779 (N_18779,N_18509,N_18202);
nor U18780 (N_18780,N_18321,N_18163);
nand U18781 (N_18781,N_18405,N_18069);
and U18782 (N_18782,N_18061,N_18109);
nor U18783 (N_18783,N_18421,N_18067);
xnor U18784 (N_18784,N_18218,N_18594);
nor U18785 (N_18785,N_18050,N_18066);
nand U18786 (N_18786,N_18012,N_18139);
or U18787 (N_18787,N_18097,N_18071);
nand U18788 (N_18788,N_18589,N_18115);
nand U18789 (N_18789,N_18365,N_18162);
nand U18790 (N_18790,N_18005,N_18299);
xnor U18791 (N_18791,N_18486,N_18093);
nor U18792 (N_18792,N_18062,N_18344);
nand U18793 (N_18793,N_18063,N_18335);
xnor U18794 (N_18794,N_18485,N_18374);
and U18795 (N_18795,N_18101,N_18591);
or U18796 (N_18796,N_18326,N_18086);
nand U18797 (N_18797,N_18332,N_18417);
nand U18798 (N_18798,N_18453,N_18041);
and U18799 (N_18799,N_18123,N_18280);
xnor U18800 (N_18800,N_18559,N_18025);
and U18801 (N_18801,N_18113,N_18450);
nor U18802 (N_18802,N_18226,N_18241);
or U18803 (N_18803,N_18151,N_18056);
or U18804 (N_18804,N_18357,N_18082);
nand U18805 (N_18805,N_18504,N_18046);
and U18806 (N_18806,N_18558,N_18230);
nor U18807 (N_18807,N_18500,N_18358);
and U18808 (N_18808,N_18239,N_18128);
or U18809 (N_18809,N_18564,N_18487);
nor U18810 (N_18810,N_18017,N_18407);
and U18811 (N_18811,N_18271,N_18537);
xor U18812 (N_18812,N_18130,N_18277);
or U18813 (N_18813,N_18308,N_18270);
or U18814 (N_18814,N_18502,N_18410);
xnor U18815 (N_18815,N_18439,N_18134);
and U18816 (N_18816,N_18545,N_18188);
nand U18817 (N_18817,N_18503,N_18094);
or U18818 (N_18818,N_18164,N_18169);
or U18819 (N_18819,N_18084,N_18348);
nor U18820 (N_18820,N_18303,N_18003);
nor U18821 (N_18821,N_18511,N_18287);
or U18822 (N_18822,N_18443,N_18382);
xor U18823 (N_18823,N_18148,N_18160);
and U18824 (N_18824,N_18259,N_18105);
nand U18825 (N_18825,N_18386,N_18366);
or U18826 (N_18826,N_18451,N_18460);
nand U18827 (N_18827,N_18473,N_18376);
and U18828 (N_18828,N_18083,N_18467);
nor U18829 (N_18829,N_18472,N_18574);
and U18830 (N_18830,N_18361,N_18273);
nor U18831 (N_18831,N_18254,N_18587);
and U18832 (N_18832,N_18092,N_18356);
nor U18833 (N_18833,N_18322,N_18535);
nor U18834 (N_18834,N_18416,N_18008);
and U18835 (N_18835,N_18557,N_18569);
or U18836 (N_18836,N_18309,N_18477);
xor U18837 (N_18837,N_18586,N_18302);
nor U18838 (N_18838,N_18532,N_18184);
or U18839 (N_18839,N_18513,N_18307);
xnor U18840 (N_18840,N_18048,N_18401);
xnor U18841 (N_18841,N_18170,N_18493);
nor U18842 (N_18842,N_18051,N_18120);
xor U18843 (N_18843,N_18235,N_18194);
nor U18844 (N_18844,N_18212,N_18055);
and U18845 (N_18845,N_18514,N_18570);
or U18846 (N_18846,N_18306,N_18296);
xor U18847 (N_18847,N_18181,N_18216);
and U18848 (N_18848,N_18347,N_18269);
and U18849 (N_18849,N_18038,N_18466);
xnor U18850 (N_18850,N_18126,N_18383);
or U18851 (N_18851,N_18529,N_18507);
xnor U18852 (N_18852,N_18349,N_18096);
nor U18853 (N_18853,N_18214,N_18032);
nor U18854 (N_18854,N_18217,N_18501);
nor U18855 (N_18855,N_18522,N_18415);
nor U18856 (N_18856,N_18534,N_18179);
nand U18857 (N_18857,N_18456,N_18013);
xnor U18858 (N_18858,N_18015,N_18173);
nand U18859 (N_18859,N_18002,N_18484);
nor U18860 (N_18860,N_18399,N_18138);
nand U18861 (N_18861,N_18400,N_18474);
nand U18862 (N_18862,N_18555,N_18379);
nor U18863 (N_18863,N_18334,N_18119);
nand U18864 (N_18864,N_18429,N_18276);
nor U18865 (N_18865,N_18411,N_18575);
or U18866 (N_18866,N_18132,N_18325);
xnor U18867 (N_18867,N_18403,N_18548);
or U18868 (N_18868,N_18394,N_18491);
xnor U18869 (N_18869,N_18581,N_18523);
nand U18870 (N_18870,N_18088,N_18264);
or U18871 (N_18871,N_18180,N_18551);
or U18872 (N_18872,N_18228,N_18222);
or U18873 (N_18873,N_18234,N_18177);
xor U18874 (N_18874,N_18110,N_18121);
xor U18875 (N_18875,N_18360,N_18266);
xor U18876 (N_18876,N_18198,N_18468);
or U18877 (N_18877,N_18257,N_18018);
xnor U18878 (N_18878,N_18282,N_18053);
or U18879 (N_18879,N_18526,N_18263);
xor U18880 (N_18880,N_18495,N_18246);
and U18881 (N_18881,N_18196,N_18107);
or U18882 (N_18882,N_18158,N_18044);
xor U18883 (N_18883,N_18233,N_18412);
nor U18884 (N_18884,N_18168,N_18385);
nand U18885 (N_18885,N_18498,N_18251);
xor U18886 (N_18886,N_18402,N_18525);
nor U18887 (N_18887,N_18172,N_18543);
or U18888 (N_18888,N_18193,N_18146);
nand U18889 (N_18889,N_18340,N_18345);
and U18890 (N_18890,N_18563,N_18577);
nor U18891 (N_18891,N_18432,N_18413);
nand U18892 (N_18892,N_18036,N_18552);
nor U18893 (N_18893,N_18496,N_18057);
nor U18894 (N_18894,N_18220,N_18388);
nand U18895 (N_18895,N_18341,N_18424);
nand U18896 (N_18896,N_18272,N_18043);
nor U18897 (N_18897,N_18159,N_18479);
or U18898 (N_18898,N_18215,N_18396);
nor U18899 (N_18899,N_18201,N_18006);
nor U18900 (N_18900,N_18067,N_18261);
nand U18901 (N_18901,N_18189,N_18532);
and U18902 (N_18902,N_18393,N_18179);
and U18903 (N_18903,N_18107,N_18541);
xor U18904 (N_18904,N_18500,N_18372);
xor U18905 (N_18905,N_18478,N_18557);
xnor U18906 (N_18906,N_18571,N_18465);
nand U18907 (N_18907,N_18595,N_18181);
or U18908 (N_18908,N_18101,N_18433);
and U18909 (N_18909,N_18201,N_18537);
nor U18910 (N_18910,N_18397,N_18310);
or U18911 (N_18911,N_18152,N_18445);
nor U18912 (N_18912,N_18027,N_18270);
and U18913 (N_18913,N_18484,N_18372);
nand U18914 (N_18914,N_18312,N_18207);
and U18915 (N_18915,N_18386,N_18301);
nor U18916 (N_18916,N_18493,N_18158);
xor U18917 (N_18917,N_18334,N_18121);
and U18918 (N_18918,N_18577,N_18310);
nand U18919 (N_18919,N_18490,N_18538);
and U18920 (N_18920,N_18317,N_18189);
and U18921 (N_18921,N_18403,N_18202);
nor U18922 (N_18922,N_18412,N_18240);
or U18923 (N_18923,N_18179,N_18304);
xor U18924 (N_18924,N_18280,N_18286);
nor U18925 (N_18925,N_18561,N_18272);
nand U18926 (N_18926,N_18012,N_18058);
xnor U18927 (N_18927,N_18571,N_18190);
and U18928 (N_18928,N_18081,N_18481);
and U18929 (N_18929,N_18376,N_18036);
nand U18930 (N_18930,N_18398,N_18150);
nor U18931 (N_18931,N_18434,N_18481);
and U18932 (N_18932,N_18138,N_18345);
nor U18933 (N_18933,N_18293,N_18139);
nand U18934 (N_18934,N_18355,N_18363);
nor U18935 (N_18935,N_18245,N_18369);
and U18936 (N_18936,N_18503,N_18189);
nor U18937 (N_18937,N_18132,N_18225);
nor U18938 (N_18938,N_18460,N_18241);
xnor U18939 (N_18939,N_18201,N_18467);
and U18940 (N_18940,N_18557,N_18539);
xnor U18941 (N_18941,N_18587,N_18548);
xor U18942 (N_18942,N_18567,N_18437);
nor U18943 (N_18943,N_18382,N_18143);
nand U18944 (N_18944,N_18495,N_18233);
or U18945 (N_18945,N_18391,N_18034);
nor U18946 (N_18946,N_18578,N_18516);
nand U18947 (N_18947,N_18200,N_18580);
and U18948 (N_18948,N_18541,N_18589);
nand U18949 (N_18949,N_18498,N_18125);
nor U18950 (N_18950,N_18376,N_18359);
or U18951 (N_18951,N_18021,N_18519);
nor U18952 (N_18952,N_18249,N_18173);
or U18953 (N_18953,N_18495,N_18556);
nand U18954 (N_18954,N_18173,N_18557);
nor U18955 (N_18955,N_18300,N_18250);
or U18956 (N_18956,N_18407,N_18567);
or U18957 (N_18957,N_18025,N_18038);
nand U18958 (N_18958,N_18318,N_18010);
xnor U18959 (N_18959,N_18005,N_18096);
nand U18960 (N_18960,N_18421,N_18015);
xor U18961 (N_18961,N_18171,N_18010);
nor U18962 (N_18962,N_18210,N_18199);
or U18963 (N_18963,N_18222,N_18185);
and U18964 (N_18964,N_18019,N_18313);
nand U18965 (N_18965,N_18229,N_18331);
nor U18966 (N_18966,N_18204,N_18573);
and U18967 (N_18967,N_18341,N_18437);
nor U18968 (N_18968,N_18302,N_18054);
or U18969 (N_18969,N_18362,N_18537);
or U18970 (N_18970,N_18408,N_18256);
xor U18971 (N_18971,N_18112,N_18178);
and U18972 (N_18972,N_18322,N_18138);
and U18973 (N_18973,N_18424,N_18497);
nand U18974 (N_18974,N_18047,N_18126);
nand U18975 (N_18975,N_18409,N_18586);
and U18976 (N_18976,N_18078,N_18121);
nor U18977 (N_18977,N_18149,N_18266);
and U18978 (N_18978,N_18303,N_18422);
xor U18979 (N_18979,N_18192,N_18302);
nand U18980 (N_18980,N_18575,N_18481);
nor U18981 (N_18981,N_18581,N_18383);
or U18982 (N_18982,N_18148,N_18270);
nand U18983 (N_18983,N_18198,N_18414);
nand U18984 (N_18984,N_18337,N_18254);
nor U18985 (N_18985,N_18543,N_18173);
nor U18986 (N_18986,N_18059,N_18384);
nand U18987 (N_18987,N_18265,N_18229);
and U18988 (N_18988,N_18147,N_18024);
xor U18989 (N_18989,N_18327,N_18044);
and U18990 (N_18990,N_18504,N_18267);
and U18991 (N_18991,N_18042,N_18267);
xor U18992 (N_18992,N_18538,N_18360);
nor U18993 (N_18993,N_18021,N_18159);
xnor U18994 (N_18994,N_18501,N_18346);
nand U18995 (N_18995,N_18100,N_18152);
nor U18996 (N_18996,N_18274,N_18323);
or U18997 (N_18997,N_18288,N_18491);
nand U18998 (N_18998,N_18003,N_18016);
xnor U18999 (N_18999,N_18108,N_18499);
nand U19000 (N_19000,N_18201,N_18005);
nor U19001 (N_19001,N_18559,N_18021);
and U19002 (N_19002,N_18076,N_18044);
or U19003 (N_19003,N_18212,N_18285);
nand U19004 (N_19004,N_18348,N_18572);
xnor U19005 (N_19005,N_18416,N_18272);
and U19006 (N_19006,N_18341,N_18138);
nand U19007 (N_19007,N_18503,N_18365);
nand U19008 (N_19008,N_18242,N_18215);
nand U19009 (N_19009,N_18399,N_18214);
and U19010 (N_19010,N_18030,N_18390);
nor U19011 (N_19011,N_18191,N_18552);
or U19012 (N_19012,N_18237,N_18040);
nand U19013 (N_19013,N_18439,N_18079);
xor U19014 (N_19014,N_18014,N_18187);
and U19015 (N_19015,N_18191,N_18023);
xor U19016 (N_19016,N_18344,N_18534);
or U19017 (N_19017,N_18121,N_18194);
and U19018 (N_19018,N_18458,N_18135);
or U19019 (N_19019,N_18207,N_18348);
nand U19020 (N_19020,N_18516,N_18070);
xor U19021 (N_19021,N_18300,N_18315);
nand U19022 (N_19022,N_18461,N_18582);
xor U19023 (N_19023,N_18033,N_18535);
and U19024 (N_19024,N_18318,N_18046);
and U19025 (N_19025,N_18573,N_18113);
nor U19026 (N_19026,N_18244,N_18565);
nor U19027 (N_19027,N_18303,N_18374);
nor U19028 (N_19028,N_18006,N_18547);
nor U19029 (N_19029,N_18062,N_18503);
xor U19030 (N_19030,N_18017,N_18210);
and U19031 (N_19031,N_18309,N_18286);
xor U19032 (N_19032,N_18503,N_18467);
nand U19033 (N_19033,N_18170,N_18393);
nor U19034 (N_19034,N_18113,N_18548);
xnor U19035 (N_19035,N_18468,N_18220);
xnor U19036 (N_19036,N_18416,N_18531);
nand U19037 (N_19037,N_18408,N_18132);
nand U19038 (N_19038,N_18216,N_18413);
xor U19039 (N_19039,N_18207,N_18476);
nand U19040 (N_19040,N_18030,N_18128);
and U19041 (N_19041,N_18219,N_18349);
nor U19042 (N_19042,N_18336,N_18533);
and U19043 (N_19043,N_18541,N_18226);
and U19044 (N_19044,N_18252,N_18130);
xnor U19045 (N_19045,N_18400,N_18571);
nor U19046 (N_19046,N_18158,N_18161);
or U19047 (N_19047,N_18375,N_18198);
and U19048 (N_19048,N_18267,N_18058);
nand U19049 (N_19049,N_18487,N_18211);
nand U19050 (N_19050,N_18507,N_18394);
nand U19051 (N_19051,N_18523,N_18440);
nor U19052 (N_19052,N_18105,N_18194);
or U19053 (N_19053,N_18492,N_18418);
nor U19054 (N_19054,N_18264,N_18545);
and U19055 (N_19055,N_18357,N_18526);
and U19056 (N_19056,N_18597,N_18217);
nor U19057 (N_19057,N_18373,N_18412);
and U19058 (N_19058,N_18405,N_18445);
nand U19059 (N_19059,N_18061,N_18358);
nor U19060 (N_19060,N_18390,N_18450);
and U19061 (N_19061,N_18242,N_18333);
nand U19062 (N_19062,N_18157,N_18358);
or U19063 (N_19063,N_18263,N_18453);
and U19064 (N_19064,N_18188,N_18433);
nand U19065 (N_19065,N_18054,N_18198);
nand U19066 (N_19066,N_18297,N_18002);
or U19067 (N_19067,N_18071,N_18538);
and U19068 (N_19068,N_18105,N_18033);
or U19069 (N_19069,N_18055,N_18568);
and U19070 (N_19070,N_18372,N_18001);
nor U19071 (N_19071,N_18363,N_18426);
and U19072 (N_19072,N_18130,N_18587);
xnor U19073 (N_19073,N_18134,N_18493);
xnor U19074 (N_19074,N_18199,N_18437);
or U19075 (N_19075,N_18309,N_18012);
xor U19076 (N_19076,N_18179,N_18540);
xnor U19077 (N_19077,N_18520,N_18216);
nor U19078 (N_19078,N_18194,N_18265);
nand U19079 (N_19079,N_18181,N_18404);
or U19080 (N_19080,N_18562,N_18231);
and U19081 (N_19081,N_18471,N_18537);
nor U19082 (N_19082,N_18194,N_18058);
xor U19083 (N_19083,N_18069,N_18121);
nor U19084 (N_19084,N_18286,N_18041);
xnor U19085 (N_19085,N_18003,N_18158);
or U19086 (N_19086,N_18228,N_18413);
nand U19087 (N_19087,N_18221,N_18560);
nand U19088 (N_19088,N_18084,N_18332);
nor U19089 (N_19089,N_18574,N_18466);
or U19090 (N_19090,N_18565,N_18522);
xor U19091 (N_19091,N_18005,N_18287);
nand U19092 (N_19092,N_18244,N_18198);
nand U19093 (N_19093,N_18184,N_18370);
nand U19094 (N_19094,N_18587,N_18015);
and U19095 (N_19095,N_18439,N_18420);
nand U19096 (N_19096,N_18174,N_18554);
or U19097 (N_19097,N_18427,N_18138);
nand U19098 (N_19098,N_18086,N_18489);
xnor U19099 (N_19099,N_18038,N_18033);
or U19100 (N_19100,N_18234,N_18267);
or U19101 (N_19101,N_18194,N_18035);
xnor U19102 (N_19102,N_18399,N_18425);
nor U19103 (N_19103,N_18388,N_18077);
or U19104 (N_19104,N_18388,N_18367);
nor U19105 (N_19105,N_18427,N_18504);
nor U19106 (N_19106,N_18001,N_18593);
and U19107 (N_19107,N_18280,N_18213);
and U19108 (N_19108,N_18202,N_18140);
nor U19109 (N_19109,N_18506,N_18531);
nor U19110 (N_19110,N_18558,N_18352);
nand U19111 (N_19111,N_18137,N_18205);
nand U19112 (N_19112,N_18419,N_18434);
nor U19113 (N_19113,N_18106,N_18119);
xor U19114 (N_19114,N_18435,N_18284);
nor U19115 (N_19115,N_18212,N_18270);
or U19116 (N_19116,N_18217,N_18322);
nor U19117 (N_19117,N_18455,N_18484);
nand U19118 (N_19118,N_18207,N_18211);
or U19119 (N_19119,N_18221,N_18557);
xnor U19120 (N_19120,N_18444,N_18179);
and U19121 (N_19121,N_18075,N_18505);
or U19122 (N_19122,N_18233,N_18476);
nand U19123 (N_19123,N_18586,N_18344);
xor U19124 (N_19124,N_18509,N_18404);
and U19125 (N_19125,N_18040,N_18542);
and U19126 (N_19126,N_18316,N_18504);
and U19127 (N_19127,N_18413,N_18025);
and U19128 (N_19128,N_18109,N_18080);
or U19129 (N_19129,N_18493,N_18472);
nand U19130 (N_19130,N_18031,N_18008);
and U19131 (N_19131,N_18289,N_18144);
nand U19132 (N_19132,N_18328,N_18468);
or U19133 (N_19133,N_18370,N_18578);
or U19134 (N_19134,N_18009,N_18308);
and U19135 (N_19135,N_18061,N_18576);
nand U19136 (N_19136,N_18403,N_18238);
nand U19137 (N_19137,N_18095,N_18006);
or U19138 (N_19138,N_18369,N_18091);
nand U19139 (N_19139,N_18495,N_18162);
nand U19140 (N_19140,N_18543,N_18224);
nand U19141 (N_19141,N_18100,N_18290);
and U19142 (N_19142,N_18130,N_18506);
xnor U19143 (N_19143,N_18525,N_18240);
nand U19144 (N_19144,N_18599,N_18409);
and U19145 (N_19145,N_18071,N_18090);
nand U19146 (N_19146,N_18125,N_18558);
xor U19147 (N_19147,N_18014,N_18380);
nor U19148 (N_19148,N_18204,N_18219);
nand U19149 (N_19149,N_18512,N_18318);
nand U19150 (N_19150,N_18377,N_18349);
nand U19151 (N_19151,N_18068,N_18591);
or U19152 (N_19152,N_18037,N_18391);
xor U19153 (N_19153,N_18508,N_18371);
xor U19154 (N_19154,N_18365,N_18131);
xor U19155 (N_19155,N_18560,N_18490);
and U19156 (N_19156,N_18349,N_18554);
or U19157 (N_19157,N_18062,N_18461);
nor U19158 (N_19158,N_18486,N_18179);
or U19159 (N_19159,N_18378,N_18435);
nand U19160 (N_19160,N_18347,N_18438);
and U19161 (N_19161,N_18093,N_18103);
or U19162 (N_19162,N_18549,N_18141);
or U19163 (N_19163,N_18424,N_18259);
and U19164 (N_19164,N_18370,N_18258);
or U19165 (N_19165,N_18033,N_18120);
nor U19166 (N_19166,N_18328,N_18150);
and U19167 (N_19167,N_18587,N_18470);
nor U19168 (N_19168,N_18492,N_18080);
nor U19169 (N_19169,N_18365,N_18229);
and U19170 (N_19170,N_18041,N_18214);
nor U19171 (N_19171,N_18108,N_18502);
or U19172 (N_19172,N_18503,N_18136);
and U19173 (N_19173,N_18356,N_18137);
xnor U19174 (N_19174,N_18318,N_18439);
nand U19175 (N_19175,N_18488,N_18049);
nand U19176 (N_19176,N_18181,N_18464);
xor U19177 (N_19177,N_18070,N_18329);
nor U19178 (N_19178,N_18139,N_18222);
nand U19179 (N_19179,N_18197,N_18064);
and U19180 (N_19180,N_18176,N_18149);
xnor U19181 (N_19181,N_18269,N_18437);
xor U19182 (N_19182,N_18575,N_18021);
xnor U19183 (N_19183,N_18083,N_18412);
xor U19184 (N_19184,N_18349,N_18324);
or U19185 (N_19185,N_18019,N_18174);
nor U19186 (N_19186,N_18151,N_18336);
and U19187 (N_19187,N_18132,N_18265);
xnor U19188 (N_19188,N_18345,N_18234);
and U19189 (N_19189,N_18533,N_18442);
xnor U19190 (N_19190,N_18552,N_18483);
nand U19191 (N_19191,N_18523,N_18285);
xnor U19192 (N_19192,N_18544,N_18396);
nand U19193 (N_19193,N_18086,N_18063);
xnor U19194 (N_19194,N_18004,N_18255);
nor U19195 (N_19195,N_18182,N_18551);
and U19196 (N_19196,N_18511,N_18077);
nand U19197 (N_19197,N_18320,N_18334);
nor U19198 (N_19198,N_18146,N_18062);
and U19199 (N_19199,N_18417,N_18596);
and U19200 (N_19200,N_18682,N_19188);
and U19201 (N_19201,N_18894,N_18959);
xnor U19202 (N_19202,N_18849,N_18859);
nor U19203 (N_19203,N_19139,N_19025);
nand U19204 (N_19204,N_18962,N_19110);
xnor U19205 (N_19205,N_18947,N_18882);
nand U19206 (N_19206,N_19128,N_18843);
xor U19207 (N_19207,N_18711,N_19073);
nand U19208 (N_19208,N_18747,N_18616);
nor U19209 (N_19209,N_18762,N_19052);
or U19210 (N_19210,N_18748,N_19172);
or U19211 (N_19211,N_18660,N_19086);
or U19212 (N_19212,N_19053,N_19132);
nand U19213 (N_19213,N_18898,N_19047);
xnor U19214 (N_19214,N_19100,N_18984);
nand U19215 (N_19215,N_18804,N_19013);
nand U19216 (N_19216,N_18760,N_18963);
or U19217 (N_19217,N_19083,N_19037);
nor U19218 (N_19218,N_18968,N_19043);
xnor U19219 (N_19219,N_18789,N_19026);
xnor U19220 (N_19220,N_18887,N_18815);
nor U19221 (N_19221,N_18672,N_19007);
and U19222 (N_19222,N_18647,N_19035);
nor U19223 (N_19223,N_18869,N_18839);
xor U19224 (N_19224,N_18720,N_19167);
xor U19225 (N_19225,N_18946,N_18606);
xor U19226 (N_19226,N_18793,N_19046);
xnor U19227 (N_19227,N_18733,N_19005);
and U19228 (N_19228,N_18796,N_18927);
nand U19229 (N_19229,N_19049,N_19122);
or U19230 (N_19230,N_18812,N_19018);
xnor U19231 (N_19231,N_18677,N_19089);
or U19232 (N_19232,N_19180,N_18925);
nand U19233 (N_19233,N_19150,N_18691);
or U19234 (N_19234,N_19003,N_18888);
and U19235 (N_19235,N_19121,N_18792);
xnor U19236 (N_19236,N_19011,N_18979);
nand U19237 (N_19237,N_19042,N_18614);
xor U19238 (N_19238,N_19071,N_18610);
nor U19239 (N_19239,N_19189,N_19105);
xor U19240 (N_19240,N_18814,N_18922);
xor U19241 (N_19241,N_19140,N_19145);
xor U19242 (N_19242,N_18974,N_19095);
or U19243 (N_19243,N_18870,N_18678);
xnor U19244 (N_19244,N_18794,N_18955);
or U19245 (N_19245,N_18695,N_19117);
or U19246 (N_19246,N_18665,N_18625);
and U19247 (N_19247,N_18611,N_19171);
nor U19248 (N_19248,N_18639,N_19144);
or U19249 (N_19249,N_18653,N_18645);
nor U19250 (N_19250,N_18938,N_18832);
nor U19251 (N_19251,N_19069,N_18817);
nand U19252 (N_19252,N_18634,N_19165);
or U19253 (N_19253,N_18854,N_18713);
nand U19254 (N_19254,N_18821,N_19190);
xnor U19255 (N_19255,N_18829,N_18640);
xor U19256 (N_19256,N_18709,N_19106);
nand U19257 (N_19257,N_19155,N_19153);
xnor U19258 (N_19258,N_19077,N_19068);
nor U19259 (N_19259,N_19184,N_19045);
nor U19260 (N_19260,N_18631,N_19029);
or U19261 (N_19261,N_18750,N_18826);
or U19262 (N_19262,N_18995,N_19084);
nor U19263 (N_19263,N_18694,N_19143);
and U19264 (N_19264,N_19131,N_19157);
or U19265 (N_19265,N_18809,N_18803);
nand U19266 (N_19266,N_18891,N_18836);
and U19267 (N_19267,N_18851,N_19065);
nor U19268 (N_19268,N_18884,N_18676);
xnor U19269 (N_19269,N_18737,N_18648);
or U19270 (N_19270,N_18749,N_18726);
nor U19271 (N_19271,N_19186,N_18976);
nor U19272 (N_19272,N_19075,N_19032);
or U19273 (N_19273,N_18761,N_18702);
and U19274 (N_19274,N_18656,N_18680);
or U19275 (N_19275,N_19174,N_19087);
xor U19276 (N_19276,N_18623,N_18717);
nand U19277 (N_19277,N_18655,N_18861);
nand U19278 (N_19278,N_18918,N_18936);
and U19279 (N_19279,N_19182,N_18802);
or U19280 (N_19280,N_19094,N_18742);
xor U19281 (N_19281,N_18970,N_18950);
or U19282 (N_19282,N_19010,N_19170);
and U19283 (N_19283,N_19156,N_19063);
xor U19284 (N_19284,N_19097,N_19112);
and U19285 (N_19285,N_18977,N_18624);
nand U19286 (N_19286,N_18899,N_18909);
or U19287 (N_19287,N_18806,N_18732);
nand U19288 (N_19288,N_19193,N_19024);
xnor U19289 (N_19289,N_18904,N_18704);
and U19290 (N_19290,N_18828,N_19034);
nand U19291 (N_19291,N_19054,N_19123);
or U19292 (N_19292,N_18845,N_18881);
nand U19293 (N_19293,N_18981,N_18774);
or U19294 (N_19294,N_19183,N_18915);
xor U19295 (N_19295,N_19078,N_19133);
xor U19296 (N_19296,N_18951,N_18790);
nor U19297 (N_19297,N_18605,N_18818);
xor U19298 (N_19298,N_18613,N_18902);
and U19299 (N_19299,N_19137,N_18958);
nand U19300 (N_19300,N_18889,N_19038);
nand U19301 (N_19301,N_19022,N_19126);
nand U19302 (N_19302,N_19019,N_18863);
or U19303 (N_19303,N_19161,N_19093);
xnor U19304 (N_19304,N_18693,N_18940);
or U19305 (N_19305,N_18913,N_18763);
nor U19306 (N_19306,N_18654,N_19058);
nand U19307 (N_19307,N_18673,N_18727);
nand U19308 (N_19308,N_18905,N_18692);
nand U19309 (N_19309,N_18852,N_18866);
nand U19310 (N_19310,N_19080,N_19050);
and U19311 (N_19311,N_18607,N_18716);
nor U19312 (N_19312,N_18808,N_18874);
nand U19313 (N_19313,N_18816,N_19012);
or U19314 (N_19314,N_18679,N_19185);
nand U19315 (N_19315,N_19055,N_18683);
or U19316 (N_19316,N_19159,N_19027);
or U19317 (N_19317,N_18651,N_18671);
xnor U19318 (N_19318,N_18819,N_19127);
or U19319 (N_19319,N_19002,N_18893);
nand U19320 (N_19320,N_19001,N_18919);
nor U19321 (N_19321,N_19099,N_19191);
xor U19322 (N_19322,N_18746,N_18949);
nor U19323 (N_19323,N_19057,N_18797);
nand U19324 (N_19324,N_18764,N_18699);
and U19325 (N_19325,N_19168,N_18901);
nor U19326 (N_19326,N_18779,N_18771);
xnor U19327 (N_19327,N_19044,N_19160);
xnor U19328 (N_19328,N_19000,N_18621);
or U19329 (N_19329,N_18911,N_19192);
or U19330 (N_19330,N_18715,N_18706);
and U19331 (N_19331,N_18662,N_18932);
or U19332 (N_19332,N_18751,N_19173);
xnor U19333 (N_19333,N_18707,N_18945);
xnor U19334 (N_19334,N_18772,N_19102);
nand U19335 (N_19335,N_19120,N_18633);
xnor U19336 (N_19336,N_18877,N_18622);
nand U19337 (N_19337,N_18853,N_18987);
or U19338 (N_19338,N_18862,N_18739);
xnor U19339 (N_19339,N_18840,N_18752);
or U19340 (N_19340,N_19135,N_19028);
xnor U19341 (N_19341,N_19021,N_19004);
and U19342 (N_19342,N_18738,N_18965);
and U19343 (N_19343,N_18994,N_18907);
nor U19344 (N_19344,N_18883,N_18719);
nand U19345 (N_19345,N_18867,N_18784);
xnor U19346 (N_19346,N_19141,N_18873);
xnor U19347 (N_19347,N_18658,N_18753);
and U19348 (N_19348,N_18967,N_18833);
or U19349 (N_19349,N_18910,N_18787);
nand U19350 (N_19350,N_18657,N_18697);
and U19351 (N_19351,N_19076,N_18856);
xor U19352 (N_19352,N_18666,N_18628);
and U19353 (N_19353,N_18933,N_19014);
nor U19354 (N_19354,N_18777,N_18834);
xor U19355 (N_19355,N_18937,N_18928);
xor U19356 (N_19356,N_18600,N_18961);
and U19357 (N_19357,N_18988,N_18780);
and U19358 (N_19358,N_19179,N_19147);
xor U19359 (N_19359,N_19067,N_18886);
nor U19360 (N_19360,N_19138,N_18646);
nand U19361 (N_19361,N_18942,N_18824);
nor U19362 (N_19362,N_18674,N_19166);
and U19363 (N_19363,N_19064,N_19091);
or U19364 (N_19364,N_18973,N_18602);
nand U19365 (N_19365,N_18811,N_19072);
xnor U19366 (N_19366,N_18810,N_18791);
nand U19367 (N_19367,N_18844,N_18885);
xor U19368 (N_19368,N_18953,N_18681);
or U19369 (N_19369,N_18822,N_19195);
xnor U19370 (N_19370,N_18759,N_18795);
nor U19371 (N_19371,N_18754,N_18944);
nand U19372 (N_19372,N_18858,N_19119);
or U19373 (N_19373,N_19092,N_18848);
xnor U19374 (N_19374,N_18982,N_18620);
and U19375 (N_19375,N_18931,N_18825);
or U19376 (N_19376,N_19146,N_18686);
nor U19377 (N_19377,N_18990,N_19151);
and U19378 (N_19378,N_19148,N_19197);
xor U19379 (N_19379,N_18855,N_19124);
nor U19380 (N_19380,N_18871,N_18705);
nor U19381 (N_19381,N_18629,N_18986);
or U19382 (N_19382,N_18743,N_19108);
and U19383 (N_19383,N_18916,N_18917);
nor U19384 (N_19384,N_18842,N_19074);
nand U19385 (N_19385,N_18775,N_19113);
nor U19386 (N_19386,N_18929,N_18661);
xor U19387 (N_19387,N_19006,N_18667);
xnor U19388 (N_19388,N_18670,N_18914);
xnor U19389 (N_19389,N_19107,N_18729);
nor U19390 (N_19390,N_18685,N_19096);
nand U19391 (N_19391,N_19152,N_19114);
nor U19392 (N_19392,N_18926,N_18934);
nand U19393 (N_19393,N_18805,N_19125);
or U19394 (N_19394,N_18807,N_18698);
or U19395 (N_19395,N_18690,N_19062);
nor U19396 (N_19396,N_19030,N_19059);
nand U19397 (N_19397,N_19136,N_18770);
nand U19398 (N_19398,N_18608,N_19082);
or U19399 (N_19399,N_19101,N_19041);
xor U19400 (N_19400,N_19104,N_19176);
xnor U19401 (N_19401,N_18798,N_18714);
or U19402 (N_19402,N_18786,N_18920);
nand U19403 (N_19403,N_18778,N_18703);
xor U19404 (N_19404,N_18688,N_18708);
xnor U19405 (N_19405,N_18989,N_19163);
xor U19406 (N_19406,N_19118,N_19090);
nor U19407 (N_19407,N_18892,N_18735);
nor U19408 (N_19408,N_19115,N_18998);
nand U19409 (N_19409,N_18701,N_19154);
xor U19410 (N_19410,N_19036,N_18785);
nor U19411 (N_19411,N_18609,N_18601);
nand U19412 (N_19412,N_19177,N_18827);
and U19413 (N_19413,N_19178,N_18734);
nand U19414 (N_19414,N_18930,N_18993);
nand U19415 (N_19415,N_18923,N_18723);
xnor U19416 (N_19416,N_18687,N_18758);
nor U19417 (N_19417,N_18971,N_18972);
nand U19418 (N_19418,N_18943,N_18831);
and U19419 (N_19419,N_18684,N_18992);
and U19420 (N_19420,N_18903,N_19061);
or U19421 (N_19421,N_19129,N_18868);
nand U19422 (N_19422,N_18924,N_18700);
nor U19423 (N_19423,N_19088,N_18740);
and U19424 (N_19424,N_18835,N_18636);
nor U19425 (N_19425,N_18736,N_18906);
or U19426 (N_19426,N_18637,N_18980);
nor U19427 (N_19427,N_18801,N_18664);
or U19428 (N_19428,N_18879,N_19085);
and U19429 (N_19429,N_18712,N_18604);
and U19430 (N_19430,N_18964,N_19130);
or U19431 (N_19431,N_18941,N_18895);
or U19432 (N_19432,N_18939,N_18837);
xor U19433 (N_19433,N_18897,N_18782);
xor U19434 (N_19434,N_19009,N_18721);
nor U19435 (N_19435,N_18878,N_18765);
nand U19436 (N_19436,N_19116,N_18652);
nand U19437 (N_19437,N_18756,N_18788);
nor U19438 (N_19438,N_18725,N_18718);
xnor U19439 (N_19439,N_19103,N_19060);
or U19440 (N_19440,N_18956,N_19031);
or U19441 (N_19441,N_18663,N_19066);
nor U19442 (N_19442,N_18997,N_18847);
nand U19443 (N_19443,N_19017,N_18650);
or U19444 (N_19444,N_19111,N_19142);
and U19445 (N_19445,N_18872,N_19056);
xor U19446 (N_19446,N_18948,N_18991);
or U19447 (N_19447,N_18978,N_18776);
nand U19448 (N_19448,N_18800,N_19181);
nor U19449 (N_19449,N_18983,N_18921);
or U19450 (N_19450,N_19070,N_18783);
nand U19451 (N_19451,N_19020,N_19169);
nand U19452 (N_19452,N_18767,N_18612);
nor U19453 (N_19453,N_18630,N_19198);
xor U19454 (N_19454,N_18860,N_18865);
nor U19455 (N_19455,N_19016,N_18952);
nor U19456 (N_19456,N_18799,N_18954);
nand U19457 (N_19457,N_18757,N_19199);
and U19458 (N_19458,N_18985,N_18850);
or U19459 (N_19459,N_19008,N_18966);
nand U19460 (N_19460,N_18668,N_18830);
or U19461 (N_19461,N_19175,N_18643);
nand U19462 (N_19462,N_18669,N_18912);
or U19463 (N_19463,N_18975,N_19040);
nand U19464 (N_19464,N_18823,N_18999);
xor U19465 (N_19465,N_18781,N_18880);
and U19466 (N_19466,N_18766,N_19023);
nand U19467 (N_19467,N_18744,N_18641);
nor U19468 (N_19468,N_19187,N_18846);
nor U19469 (N_19469,N_18813,N_18768);
xnor U19470 (N_19470,N_18755,N_18638);
nand U19471 (N_19471,N_18635,N_18675);
nor U19472 (N_19472,N_19015,N_19149);
nand U19473 (N_19473,N_19134,N_18722);
and U19474 (N_19474,N_18626,N_18960);
or U19475 (N_19475,N_18730,N_19051);
or U19476 (N_19476,N_18728,N_18890);
and U19477 (N_19477,N_19109,N_18908);
xnor U19478 (N_19478,N_19098,N_19048);
and U19479 (N_19479,N_18644,N_18864);
or U19480 (N_19480,N_18820,N_18857);
and U19481 (N_19481,N_18619,N_19194);
or U19482 (N_19482,N_18838,N_18773);
nor U19483 (N_19483,N_18659,N_18617);
or U19484 (N_19484,N_19033,N_18618);
nand U19485 (N_19485,N_18876,N_18615);
nor U19486 (N_19486,N_18769,N_19164);
and U19487 (N_19487,N_18900,N_18841);
xor U19488 (N_19488,N_19079,N_18741);
xnor U19489 (N_19489,N_18745,N_19039);
xor U19490 (N_19490,N_18632,N_19162);
nor U19491 (N_19491,N_18969,N_18896);
or U19492 (N_19492,N_18724,N_18935);
or U19493 (N_19493,N_18642,N_19081);
nor U19494 (N_19494,N_18603,N_18996);
nand U19495 (N_19495,N_18731,N_18696);
nor U19496 (N_19496,N_18957,N_19158);
xor U19497 (N_19497,N_18627,N_18710);
nand U19498 (N_19498,N_18649,N_18875);
nand U19499 (N_19499,N_19196,N_18689);
and U19500 (N_19500,N_19065,N_18660);
xor U19501 (N_19501,N_18758,N_18814);
xnor U19502 (N_19502,N_19179,N_18899);
and U19503 (N_19503,N_18669,N_18627);
or U19504 (N_19504,N_18874,N_19123);
and U19505 (N_19505,N_18821,N_18882);
and U19506 (N_19506,N_18664,N_18802);
or U19507 (N_19507,N_19113,N_19004);
and U19508 (N_19508,N_18709,N_19067);
xor U19509 (N_19509,N_19038,N_19150);
nor U19510 (N_19510,N_18755,N_19099);
and U19511 (N_19511,N_18629,N_18653);
or U19512 (N_19512,N_19009,N_19148);
or U19513 (N_19513,N_19014,N_18680);
and U19514 (N_19514,N_19040,N_19142);
or U19515 (N_19515,N_18749,N_19155);
or U19516 (N_19516,N_19178,N_19046);
and U19517 (N_19517,N_18956,N_19006);
nand U19518 (N_19518,N_19103,N_18831);
nor U19519 (N_19519,N_18914,N_19016);
or U19520 (N_19520,N_19147,N_18911);
and U19521 (N_19521,N_19197,N_18700);
xor U19522 (N_19522,N_19010,N_18721);
and U19523 (N_19523,N_18995,N_19187);
or U19524 (N_19524,N_18776,N_19086);
and U19525 (N_19525,N_18930,N_18956);
nor U19526 (N_19526,N_18981,N_18755);
or U19527 (N_19527,N_19179,N_18944);
or U19528 (N_19528,N_18829,N_18997);
xnor U19529 (N_19529,N_19155,N_19022);
nor U19530 (N_19530,N_18737,N_18890);
nand U19531 (N_19531,N_18959,N_18799);
or U19532 (N_19532,N_18932,N_19086);
or U19533 (N_19533,N_18770,N_19104);
nor U19534 (N_19534,N_18705,N_18899);
nor U19535 (N_19535,N_19040,N_18883);
and U19536 (N_19536,N_18805,N_18711);
nor U19537 (N_19537,N_18944,N_18603);
or U19538 (N_19538,N_18910,N_19180);
xor U19539 (N_19539,N_18908,N_18710);
xnor U19540 (N_19540,N_19045,N_18703);
nor U19541 (N_19541,N_18704,N_18857);
nor U19542 (N_19542,N_19003,N_18912);
or U19543 (N_19543,N_18887,N_18788);
xnor U19544 (N_19544,N_18967,N_18643);
nor U19545 (N_19545,N_18638,N_18632);
and U19546 (N_19546,N_19057,N_19061);
nor U19547 (N_19547,N_18668,N_18692);
or U19548 (N_19548,N_18930,N_19174);
xnor U19549 (N_19549,N_18930,N_18616);
nor U19550 (N_19550,N_18999,N_19049);
and U19551 (N_19551,N_19199,N_18862);
or U19552 (N_19552,N_18824,N_18970);
or U19553 (N_19553,N_18905,N_19015);
xnor U19554 (N_19554,N_18817,N_19062);
xnor U19555 (N_19555,N_18799,N_18974);
or U19556 (N_19556,N_18740,N_18639);
xnor U19557 (N_19557,N_18722,N_19096);
or U19558 (N_19558,N_18643,N_18787);
nor U19559 (N_19559,N_18695,N_19169);
and U19560 (N_19560,N_18903,N_19140);
nor U19561 (N_19561,N_19012,N_18745);
nor U19562 (N_19562,N_19076,N_18732);
xor U19563 (N_19563,N_18668,N_19028);
and U19564 (N_19564,N_18602,N_18821);
nor U19565 (N_19565,N_18829,N_18781);
nand U19566 (N_19566,N_18791,N_18920);
or U19567 (N_19567,N_18822,N_18909);
xnor U19568 (N_19568,N_18600,N_19066);
xnor U19569 (N_19569,N_18857,N_19056);
or U19570 (N_19570,N_18775,N_18742);
nand U19571 (N_19571,N_18782,N_18875);
or U19572 (N_19572,N_18840,N_18918);
xor U19573 (N_19573,N_19108,N_18909);
xnor U19574 (N_19574,N_18872,N_19004);
or U19575 (N_19575,N_19037,N_18701);
or U19576 (N_19576,N_18914,N_19057);
and U19577 (N_19577,N_18702,N_18692);
nor U19578 (N_19578,N_18928,N_19193);
or U19579 (N_19579,N_19143,N_18676);
xnor U19580 (N_19580,N_18802,N_18914);
nand U19581 (N_19581,N_19121,N_18933);
nor U19582 (N_19582,N_18729,N_19092);
xor U19583 (N_19583,N_18741,N_18637);
or U19584 (N_19584,N_18841,N_18656);
nor U19585 (N_19585,N_18967,N_18788);
xnor U19586 (N_19586,N_19039,N_19163);
xnor U19587 (N_19587,N_18951,N_18787);
or U19588 (N_19588,N_18879,N_19138);
or U19589 (N_19589,N_18614,N_19014);
and U19590 (N_19590,N_18661,N_18699);
or U19591 (N_19591,N_18869,N_18940);
or U19592 (N_19592,N_19012,N_18733);
nand U19593 (N_19593,N_19150,N_18969);
xnor U19594 (N_19594,N_19164,N_18829);
or U19595 (N_19595,N_18944,N_18721);
nor U19596 (N_19596,N_19112,N_18711);
or U19597 (N_19597,N_18924,N_19102);
and U19598 (N_19598,N_19127,N_18924);
nand U19599 (N_19599,N_19117,N_18868);
or U19600 (N_19600,N_18964,N_18745);
nand U19601 (N_19601,N_18676,N_18685);
xor U19602 (N_19602,N_19194,N_18841);
nand U19603 (N_19603,N_18864,N_18706);
xnor U19604 (N_19604,N_18679,N_19136);
nor U19605 (N_19605,N_18704,N_18709);
and U19606 (N_19606,N_18757,N_18946);
and U19607 (N_19607,N_18672,N_18874);
nor U19608 (N_19608,N_18656,N_18764);
xor U19609 (N_19609,N_18873,N_18748);
xnor U19610 (N_19610,N_18731,N_19028);
or U19611 (N_19611,N_19165,N_18919);
or U19612 (N_19612,N_18667,N_18986);
xor U19613 (N_19613,N_19012,N_19127);
xnor U19614 (N_19614,N_18672,N_19139);
xnor U19615 (N_19615,N_19050,N_18928);
or U19616 (N_19616,N_18875,N_18667);
xor U19617 (N_19617,N_18756,N_18831);
and U19618 (N_19618,N_18796,N_19001);
nand U19619 (N_19619,N_18978,N_19061);
nand U19620 (N_19620,N_19097,N_18975);
xor U19621 (N_19621,N_18724,N_18857);
or U19622 (N_19622,N_19027,N_18845);
nor U19623 (N_19623,N_18965,N_18606);
and U19624 (N_19624,N_18697,N_19192);
nand U19625 (N_19625,N_18672,N_18723);
xnor U19626 (N_19626,N_18900,N_18993);
nand U19627 (N_19627,N_18827,N_18679);
nand U19628 (N_19628,N_18923,N_18608);
and U19629 (N_19629,N_18659,N_18769);
and U19630 (N_19630,N_19135,N_18718);
nor U19631 (N_19631,N_19155,N_18693);
nor U19632 (N_19632,N_18728,N_18796);
nand U19633 (N_19633,N_18814,N_19115);
xor U19634 (N_19634,N_18896,N_18636);
nand U19635 (N_19635,N_19078,N_19176);
and U19636 (N_19636,N_18837,N_18770);
nor U19637 (N_19637,N_19034,N_18608);
nor U19638 (N_19638,N_18821,N_18696);
and U19639 (N_19639,N_19171,N_19179);
nor U19640 (N_19640,N_18972,N_19187);
nor U19641 (N_19641,N_18728,N_18968);
or U19642 (N_19642,N_19064,N_18816);
and U19643 (N_19643,N_18921,N_18814);
nor U19644 (N_19644,N_18616,N_18711);
nand U19645 (N_19645,N_19119,N_18827);
nand U19646 (N_19646,N_18840,N_19033);
or U19647 (N_19647,N_18748,N_19130);
or U19648 (N_19648,N_18830,N_18601);
nand U19649 (N_19649,N_18645,N_18952);
xnor U19650 (N_19650,N_19068,N_18615);
nor U19651 (N_19651,N_19001,N_19002);
and U19652 (N_19652,N_19176,N_18731);
nor U19653 (N_19653,N_18771,N_18696);
and U19654 (N_19654,N_18940,N_18640);
and U19655 (N_19655,N_19077,N_18976);
xor U19656 (N_19656,N_18719,N_18930);
xnor U19657 (N_19657,N_18720,N_18601);
xor U19658 (N_19658,N_19160,N_18928);
or U19659 (N_19659,N_18936,N_19012);
xnor U19660 (N_19660,N_19117,N_19070);
nor U19661 (N_19661,N_18713,N_19195);
and U19662 (N_19662,N_19063,N_19111);
nor U19663 (N_19663,N_19042,N_18795);
nand U19664 (N_19664,N_18730,N_18994);
nand U19665 (N_19665,N_19103,N_18990);
or U19666 (N_19666,N_19167,N_18927);
and U19667 (N_19667,N_18959,N_19184);
and U19668 (N_19668,N_19009,N_18789);
or U19669 (N_19669,N_19010,N_18810);
and U19670 (N_19670,N_19010,N_18974);
xor U19671 (N_19671,N_18600,N_18802);
or U19672 (N_19672,N_19035,N_19025);
nor U19673 (N_19673,N_18948,N_18761);
or U19674 (N_19674,N_19134,N_18725);
xnor U19675 (N_19675,N_19175,N_19093);
or U19676 (N_19676,N_19079,N_18706);
or U19677 (N_19677,N_19017,N_18680);
and U19678 (N_19678,N_18711,N_19104);
and U19679 (N_19679,N_19190,N_18964);
nor U19680 (N_19680,N_19121,N_18900);
nand U19681 (N_19681,N_19179,N_19050);
nor U19682 (N_19682,N_18851,N_18695);
xor U19683 (N_19683,N_19006,N_18891);
nor U19684 (N_19684,N_18919,N_18937);
nor U19685 (N_19685,N_18610,N_19121);
or U19686 (N_19686,N_19173,N_18807);
xor U19687 (N_19687,N_18784,N_18892);
and U19688 (N_19688,N_18663,N_18915);
xnor U19689 (N_19689,N_19191,N_18712);
xor U19690 (N_19690,N_18676,N_18874);
and U19691 (N_19691,N_18626,N_19162);
xnor U19692 (N_19692,N_19049,N_18991);
xor U19693 (N_19693,N_19006,N_18999);
xor U19694 (N_19694,N_19158,N_19119);
or U19695 (N_19695,N_19039,N_18854);
nor U19696 (N_19696,N_18787,N_18600);
xor U19697 (N_19697,N_18745,N_19187);
or U19698 (N_19698,N_19091,N_18986);
or U19699 (N_19699,N_19123,N_18611);
or U19700 (N_19700,N_18658,N_18808);
and U19701 (N_19701,N_18750,N_18974);
and U19702 (N_19702,N_19103,N_18819);
nand U19703 (N_19703,N_19098,N_19196);
xor U19704 (N_19704,N_18963,N_18852);
nor U19705 (N_19705,N_18762,N_18818);
xnor U19706 (N_19706,N_18971,N_18669);
nor U19707 (N_19707,N_19135,N_19145);
nand U19708 (N_19708,N_18742,N_18862);
nand U19709 (N_19709,N_18738,N_18859);
and U19710 (N_19710,N_19079,N_18747);
nand U19711 (N_19711,N_18874,N_18938);
nor U19712 (N_19712,N_18969,N_19040);
or U19713 (N_19713,N_19085,N_19044);
and U19714 (N_19714,N_19108,N_18804);
and U19715 (N_19715,N_18899,N_18644);
and U19716 (N_19716,N_18861,N_18786);
nor U19717 (N_19717,N_18726,N_18979);
xnor U19718 (N_19718,N_19028,N_19151);
or U19719 (N_19719,N_18810,N_19186);
xnor U19720 (N_19720,N_18961,N_19183);
nand U19721 (N_19721,N_18693,N_18658);
and U19722 (N_19722,N_18644,N_18767);
xnor U19723 (N_19723,N_18970,N_18847);
nor U19724 (N_19724,N_18927,N_18915);
or U19725 (N_19725,N_18993,N_18725);
or U19726 (N_19726,N_19002,N_18943);
or U19727 (N_19727,N_18979,N_19104);
or U19728 (N_19728,N_18787,N_18701);
or U19729 (N_19729,N_18951,N_18885);
xnor U19730 (N_19730,N_18884,N_18970);
nor U19731 (N_19731,N_18633,N_18603);
nor U19732 (N_19732,N_18895,N_18643);
or U19733 (N_19733,N_18724,N_19018);
nor U19734 (N_19734,N_18806,N_19047);
or U19735 (N_19735,N_19061,N_18716);
nor U19736 (N_19736,N_18652,N_18943);
xnor U19737 (N_19737,N_18651,N_18870);
nor U19738 (N_19738,N_18890,N_19002);
nand U19739 (N_19739,N_19127,N_19024);
xnor U19740 (N_19740,N_18867,N_18744);
and U19741 (N_19741,N_19004,N_18993);
nor U19742 (N_19742,N_19096,N_18831);
and U19743 (N_19743,N_19117,N_18716);
nor U19744 (N_19744,N_18604,N_19107);
xor U19745 (N_19745,N_18744,N_18883);
or U19746 (N_19746,N_19079,N_18924);
nand U19747 (N_19747,N_18770,N_18985);
nand U19748 (N_19748,N_19107,N_18692);
and U19749 (N_19749,N_19069,N_19111);
xor U19750 (N_19750,N_19041,N_18887);
nor U19751 (N_19751,N_19118,N_18645);
nand U19752 (N_19752,N_19192,N_18903);
nand U19753 (N_19753,N_18926,N_18993);
nand U19754 (N_19754,N_18754,N_18925);
or U19755 (N_19755,N_18623,N_19174);
or U19756 (N_19756,N_18709,N_18777);
or U19757 (N_19757,N_18791,N_18724);
xor U19758 (N_19758,N_19055,N_19198);
and U19759 (N_19759,N_18777,N_18838);
xor U19760 (N_19760,N_18731,N_19015);
and U19761 (N_19761,N_19116,N_18855);
and U19762 (N_19762,N_18938,N_19007);
and U19763 (N_19763,N_18984,N_19146);
or U19764 (N_19764,N_19033,N_18709);
xor U19765 (N_19765,N_18730,N_18757);
or U19766 (N_19766,N_18714,N_19097);
or U19767 (N_19767,N_18827,N_19175);
nand U19768 (N_19768,N_18695,N_18830);
nor U19769 (N_19769,N_19129,N_18994);
xnor U19770 (N_19770,N_18884,N_19147);
and U19771 (N_19771,N_18969,N_18742);
or U19772 (N_19772,N_18643,N_19016);
nor U19773 (N_19773,N_18883,N_18679);
xor U19774 (N_19774,N_18725,N_19111);
or U19775 (N_19775,N_19143,N_18824);
nor U19776 (N_19776,N_18966,N_18782);
or U19777 (N_19777,N_19153,N_19123);
nand U19778 (N_19778,N_19113,N_19063);
nand U19779 (N_19779,N_18722,N_18608);
xor U19780 (N_19780,N_18818,N_18638);
or U19781 (N_19781,N_19150,N_18648);
xor U19782 (N_19782,N_18769,N_18762);
nand U19783 (N_19783,N_19027,N_18705);
or U19784 (N_19784,N_18705,N_19179);
and U19785 (N_19785,N_18668,N_18936);
nand U19786 (N_19786,N_18760,N_18666);
nand U19787 (N_19787,N_18882,N_19116);
or U19788 (N_19788,N_18787,N_18601);
nor U19789 (N_19789,N_19125,N_19192);
or U19790 (N_19790,N_18903,N_19113);
or U19791 (N_19791,N_18611,N_19003);
xor U19792 (N_19792,N_18699,N_18886);
nand U19793 (N_19793,N_19029,N_19055);
or U19794 (N_19794,N_18779,N_18712);
nand U19795 (N_19795,N_18746,N_18771);
xnor U19796 (N_19796,N_19021,N_19079);
nand U19797 (N_19797,N_19123,N_18995);
or U19798 (N_19798,N_19090,N_19084);
and U19799 (N_19799,N_18914,N_19174);
or U19800 (N_19800,N_19497,N_19561);
nand U19801 (N_19801,N_19568,N_19709);
nor U19802 (N_19802,N_19513,N_19333);
xnor U19803 (N_19803,N_19583,N_19684);
or U19804 (N_19804,N_19677,N_19464);
nand U19805 (N_19805,N_19711,N_19643);
and U19806 (N_19806,N_19300,N_19452);
nor U19807 (N_19807,N_19616,N_19748);
nand U19808 (N_19808,N_19761,N_19437);
nand U19809 (N_19809,N_19678,N_19779);
nand U19810 (N_19810,N_19518,N_19278);
nor U19811 (N_19811,N_19390,N_19345);
nor U19812 (N_19812,N_19537,N_19439);
and U19813 (N_19813,N_19474,N_19758);
or U19814 (N_19814,N_19253,N_19687);
xor U19815 (N_19815,N_19732,N_19455);
nor U19816 (N_19816,N_19394,N_19468);
and U19817 (N_19817,N_19381,N_19329);
nand U19818 (N_19818,N_19630,N_19438);
or U19819 (N_19819,N_19344,N_19231);
or U19820 (N_19820,N_19224,N_19773);
and U19821 (N_19821,N_19782,N_19375);
xor U19822 (N_19822,N_19641,N_19338);
and U19823 (N_19823,N_19774,N_19636);
nand U19824 (N_19824,N_19533,N_19543);
xor U19825 (N_19825,N_19429,N_19729);
xor U19826 (N_19826,N_19760,N_19622);
nand U19827 (N_19827,N_19637,N_19649);
and U19828 (N_19828,N_19451,N_19646);
and U19829 (N_19829,N_19784,N_19236);
nor U19830 (N_19830,N_19431,N_19698);
nor U19831 (N_19831,N_19564,N_19785);
or U19832 (N_19832,N_19306,N_19220);
nand U19833 (N_19833,N_19744,N_19660);
xor U19834 (N_19834,N_19418,N_19434);
nor U19835 (N_19835,N_19415,N_19588);
nand U19836 (N_19836,N_19250,N_19466);
xor U19837 (N_19837,N_19395,N_19465);
and U19838 (N_19838,N_19509,N_19682);
nand U19839 (N_19839,N_19757,N_19221);
nand U19840 (N_19840,N_19204,N_19659);
and U19841 (N_19841,N_19288,N_19461);
and U19842 (N_19842,N_19502,N_19712);
or U19843 (N_19843,N_19282,N_19740);
nor U19844 (N_19844,N_19320,N_19410);
and U19845 (N_19845,N_19789,N_19491);
xnor U19846 (N_19846,N_19627,N_19673);
nand U19847 (N_19847,N_19535,N_19398);
and U19848 (N_19848,N_19402,N_19353);
nor U19849 (N_19849,N_19367,N_19668);
and U19850 (N_19850,N_19790,N_19430);
xor U19851 (N_19851,N_19484,N_19728);
nor U19852 (N_19852,N_19585,N_19610);
nor U19853 (N_19853,N_19263,N_19523);
or U19854 (N_19854,N_19735,N_19490);
xnor U19855 (N_19855,N_19244,N_19623);
nor U19856 (N_19856,N_19373,N_19731);
nand U19857 (N_19857,N_19544,N_19794);
xnor U19858 (N_19858,N_19493,N_19412);
nor U19859 (N_19859,N_19619,N_19498);
xnor U19860 (N_19860,N_19267,N_19615);
nand U19861 (N_19861,N_19446,N_19587);
nor U19862 (N_19862,N_19571,N_19462);
and U19863 (N_19863,N_19207,N_19631);
and U19864 (N_19864,N_19440,N_19213);
and U19865 (N_19865,N_19792,N_19422);
nor U19866 (N_19866,N_19246,N_19256);
nor U19867 (N_19867,N_19396,N_19601);
and U19868 (N_19868,N_19596,N_19399);
and U19869 (N_19869,N_19548,N_19203);
and U19870 (N_19870,N_19304,N_19458);
nor U19871 (N_19871,N_19397,N_19679);
nand U19872 (N_19872,N_19621,N_19211);
nand U19873 (N_19873,N_19352,N_19232);
or U19874 (N_19874,N_19692,N_19209);
nand U19875 (N_19875,N_19614,N_19536);
or U19876 (N_19876,N_19481,N_19460);
xnor U19877 (N_19877,N_19274,N_19756);
nand U19878 (N_19878,N_19666,N_19348);
and U19879 (N_19879,N_19701,N_19473);
and U19880 (N_19880,N_19295,N_19293);
nand U19881 (N_19881,N_19442,N_19405);
and U19882 (N_19882,N_19765,N_19307);
or U19883 (N_19883,N_19443,N_19590);
nor U19884 (N_19884,N_19285,N_19272);
xnor U19885 (N_19885,N_19362,N_19233);
xnor U19886 (N_19886,N_19663,N_19693);
nand U19887 (N_19887,N_19634,N_19382);
or U19888 (N_19888,N_19477,N_19549);
xnor U19889 (N_19889,N_19715,N_19552);
and U19890 (N_19890,N_19741,N_19763);
nor U19891 (N_19891,N_19551,N_19403);
or U19892 (N_19892,N_19457,N_19241);
or U19893 (N_19893,N_19448,N_19234);
xor U19894 (N_19894,N_19360,N_19605);
xor U19895 (N_19895,N_19432,N_19230);
and U19896 (N_19896,N_19525,N_19516);
nand U19897 (N_19897,N_19328,N_19556);
xnor U19898 (N_19898,N_19414,N_19228);
nor U19899 (N_19899,N_19734,N_19714);
xnor U19900 (N_19900,N_19742,N_19512);
nand U19901 (N_19901,N_19769,N_19686);
nor U19902 (N_19902,N_19326,N_19424);
and U19903 (N_19903,N_19771,N_19553);
and U19904 (N_19904,N_19582,N_19308);
or U19905 (N_19905,N_19235,N_19644);
xnor U19906 (N_19906,N_19695,N_19459);
nand U19907 (N_19907,N_19472,N_19495);
and U19908 (N_19908,N_19633,N_19517);
and U19909 (N_19909,N_19317,N_19662);
nand U19910 (N_19910,N_19594,N_19425);
or U19911 (N_19911,N_19661,N_19566);
nand U19912 (N_19912,N_19450,N_19793);
xnor U19913 (N_19913,N_19648,N_19377);
nor U19914 (N_19914,N_19799,N_19355);
nand U19915 (N_19915,N_19505,N_19324);
xor U19916 (N_19916,N_19416,N_19389);
nor U19917 (N_19917,N_19413,N_19261);
nand U19918 (N_19918,N_19563,N_19266);
nor U19919 (N_19919,N_19584,N_19730);
nand U19920 (N_19920,N_19745,N_19264);
xnor U19921 (N_19921,N_19768,N_19762);
nand U19922 (N_19922,N_19541,N_19485);
and U19923 (N_19923,N_19640,N_19565);
nand U19924 (N_19924,N_19401,N_19704);
or U19925 (N_19925,N_19339,N_19656);
nor U19926 (N_19926,N_19453,N_19606);
and U19927 (N_19927,N_19423,N_19651);
xnor U19928 (N_19928,N_19515,N_19208);
or U19929 (N_19929,N_19751,N_19707);
nor U19930 (N_19930,N_19546,N_19327);
and U19931 (N_19931,N_19524,N_19555);
nand U19932 (N_19932,N_19371,N_19618);
nand U19933 (N_19933,N_19528,N_19289);
or U19934 (N_19934,N_19725,N_19444);
and U19935 (N_19935,N_19420,N_19589);
and U19936 (N_19936,N_19297,N_19503);
xor U19937 (N_19937,N_19316,N_19341);
nor U19938 (N_19938,N_19545,N_19212);
xnor U19939 (N_19939,N_19522,N_19222);
or U19940 (N_19940,N_19342,N_19540);
nor U19941 (N_19941,N_19617,N_19268);
nand U19942 (N_19942,N_19237,N_19226);
xnor U19943 (N_19943,N_19454,N_19358);
nand U19944 (N_19944,N_19672,N_19318);
and U19945 (N_19945,N_19499,N_19754);
or U19946 (N_19946,N_19626,N_19319);
and U19947 (N_19947,N_19788,N_19508);
or U19948 (N_19948,N_19593,N_19717);
and U19949 (N_19949,N_19550,N_19296);
nor U19950 (N_19950,N_19277,N_19383);
and U19951 (N_19951,N_19354,N_19721);
nor U19952 (N_19952,N_19343,N_19624);
nor U19953 (N_19953,N_19218,N_19560);
or U19954 (N_19954,N_19538,N_19727);
nor U19955 (N_19955,N_19558,N_19609);
nand U19956 (N_19956,N_19259,N_19325);
or U19957 (N_19957,N_19767,N_19569);
and U19958 (N_19958,N_19305,N_19724);
xor U19959 (N_19959,N_19392,N_19676);
and U19960 (N_19960,N_19510,N_19303);
or U19961 (N_19961,N_19733,N_19675);
or U19962 (N_19962,N_19706,N_19478);
and U19963 (N_19963,N_19612,N_19689);
nand U19964 (N_19964,N_19795,N_19488);
or U19965 (N_19965,N_19719,N_19554);
nor U19966 (N_19966,N_19531,N_19419);
nor U19967 (N_19967,N_19653,N_19273);
nand U19968 (N_19968,N_19321,N_19770);
xnor U19969 (N_19969,N_19703,N_19384);
xnor U19970 (N_19970,N_19281,N_19294);
or U19971 (N_19971,N_19625,N_19200);
or U19972 (N_19972,N_19298,N_19700);
nor U19973 (N_19973,N_19572,N_19716);
or U19974 (N_19974,N_19337,N_19501);
nor U19975 (N_19975,N_19702,N_19409);
xnor U19976 (N_19976,N_19628,N_19750);
nand U19977 (N_19977,N_19369,N_19796);
and U19978 (N_19978,N_19331,N_19657);
and U19979 (N_19979,N_19747,N_19665);
or U19980 (N_19980,N_19559,N_19705);
or U19981 (N_19981,N_19346,N_19311);
xor U19982 (N_19982,N_19275,N_19205);
and U19983 (N_19983,N_19262,N_19694);
and U19984 (N_19984,N_19445,N_19376);
nand U19985 (N_19985,N_19567,N_19364);
xnor U19986 (N_19986,N_19699,N_19500);
nand U19987 (N_19987,N_19313,N_19210);
nand U19988 (N_19988,N_19519,N_19737);
xnor U19989 (N_19989,N_19539,N_19562);
xor U19990 (N_19990,N_19476,N_19607);
nand U19991 (N_19991,N_19467,N_19269);
nor U19992 (N_19992,N_19449,N_19520);
nand U19993 (N_19993,N_19652,N_19547);
xnor U19994 (N_19994,N_19496,N_19279);
xnor U19995 (N_19995,N_19507,N_19766);
or U19996 (N_19996,N_19671,N_19691);
xor U19997 (N_19997,N_19664,N_19577);
nand U19998 (N_19998,N_19489,N_19280);
and U19999 (N_19999,N_19215,N_19494);
and U20000 (N_20000,N_19579,N_19746);
xor U20001 (N_20001,N_19260,N_19683);
nand U20002 (N_20002,N_19271,N_19388);
xnor U20003 (N_20003,N_19290,N_19340);
and U20004 (N_20004,N_19580,N_19781);
nor U20005 (N_20005,N_19214,N_19690);
and U20006 (N_20006,N_19791,N_19408);
xor U20007 (N_20007,N_19265,N_19254);
nand U20008 (N_20008,N_19755,N_19591);
and U20009 (N_20009,N_19310,N_19435);
nand U20010 (N_20010,N_19645,N_19611);
xor U20011 (N_20011,N_19635,N_19238);
and U20012 (N_20012,N_19312,N_19219);
xor U20013 (N_20013,N_19688,N_19713);
and U20014 (N_20014,N_19284,N_19726);
or U20015 (N_20015,N_19526,N_19391);
nand U20016 (N_20016,N_19372,N_19650);
and U20017 (N_20017,N_19753,N_19239);
nor U20018 (N_20018,N_19576,N_19336);
nor U20019 (N_20019,N_19787,N_19456);
nand U20020 (N_20020,N_19595,N_19302);
nor U20021 (N_20021,N_19603,N_19447);
xnor U20022 (N_20022,N_19251,N_19685);
nor U20023 (N_20023,N_19529,N_19385);
xnor U20024 (N_20024,N_19243,N_19411);
xor U20025 (N_20025,N_19578,N_19479);
and U20026 (N_20026,N_19357,N_19374);
or U20027 (N_20027,N_19469,N_19764);
or U20028 (N_20028,N_19287,N_19778);
nand U20029 (N_20029,N_19720,N_19323);
nand U20030 (N_20030,N_19475,N_19597);
xnor U20031 (N_20031,N_19667,N_19710);
xnor U20032 (N_20032,N_19247,N_19242);
xnor U20033 (N_20033,N_19433,N_19776);
xor U20034 (N_20034,N_19613,N_19223);
nor U20035 (N_20035,N_19581,N_19632);
nor U20036 (N_20036,N_19680,N_19249);
xnor U20037 (N_20037,N_19647,N_19570);
and U20038 (N_20038,N_19257,N_19723);
xnor U20039 (N_20039,N_19255,N_19404);
nor U20040 (N_20040,N_19542,N_19286);
xor U20041 (N_20041,N_19608,N_19330);
xnor U20042 (N_20042,N_19428,N_19521);
or U20043 (N_20043,N_19530,N_19506);
xnor U20044 (N_20044,N_19798,N_19736);
nor U20045 (N_20045,N_19332,N_19532);
nand U20046 (N_20046,N_19361,N_19363);
and U20047 (N_20047,N_19598,N_19217);
nor U20048 (N_20048,N_19334,N_19441);
and U20049 (N_20049,N_19270,N_19229);
nand U20050 (N_20050,N_19301,N_19315);
nor U20051 (N_20051,N_19240,N_19696);
or U20052 (N_20052,N_19592,N_19669);
and U20053 (N_20053,N_19514,N_19349);
or U20054 (N_20054,N_19658,N_19436);
nand U20055 (N_20055,N_19480,N_19575);
nand U20056 (N_20056,N_19786,N_19620);
or U20057 (N_20057,N_19604,N_19492);
nor U20058 (N_20058,N_19482,N_19335);
nor U20059 (N_20059,N_19586,N_19674);
and U20060 (N_20060,N_19573,N_19322);
nand U20061 (N_20061,N_19427,N_19670);
nand U20062 (N_20062,N_19504,N_19202);
nand U20063 (N_20063,N_19417,N_19638);
xnor U20064 (N_20064,N_19629,N_19527);
xnor U20065 (N_20065,N_19252,N_19350);
xor U20066 (N_20066,N_19393,N_19718);
and U20067 (N_20067,N_19406,N_19201);
or U20068 (N_20068,N_19642,N_19743);
xor U20069 (N_20069,N_19206,N_19370);
and U20070 (N_20070,N_19681,N_19739);
nor U20071 (N_20071,N_19574,N_19356);
xnor U20072 (N_20072,N_19471,N_19276);
xnor U20073 (N_20073,N_19379,N_19463);
nor U20074 (N_20074,N_19599,N_19749);
nand U20075 (N_20075,N_19557,N_19245);
nor U20076 (N_20076,N_19225,N_19347);
nor U20077 (N_20077,N_19486,N_19722);
xor U20078 (N_20078,N_19291,N_19602);
xnor U20079 (N_20079,N_19600,N_19314);
or U20080 (N_20080,N_19534,N_19759);
nand U20081 (N_20081,N_19421,N_19780);
xor U20082 (N_20082,N_19365,N_19483);
xnor U20083 (N_20083,N_19380,N_19772);
and U20084 (N_20084,N_19407,N_19708);
xor U20085 (N_20085,N_19697,N_19283);
nor U20086 (N_20086,N_19299,N_19248);
xor U20087 (N_20087,N_19400,N_19487);
or U20088 (N_20088,N_19783,N_19797);
nand U20089 (N_20089,N_19738,N_19366);
and U20090 (N_20090,N_19654,N_19777);
nor U20091 (N_20091,N_19386,N_19426);
nand U20092 (N_20092,N_19292,N_19309);
or U20093 (N_20093,N_19227,N_19258);
xnor U20094 (N_20094,N_19387,N_19368);
nand U20095 (N_20095,N_19216,N_19775);
or U20096 (N_20096,N_19359,N_19351);
nor U20097 (N_20097,N_19470,N_19655);
nor U20098 (N_20098,N_19752,N_19639);
and U20099 (N_20099,N_19511,N_19378);
nand U20100 (N_20100,N_19481,N_19603);
xnor U20101 (N_20101,N_19787,N_19780);
nand U20102 (N_20102,N_19539,N_19705);
xor U20103 (N_20103,N_19742,N_19476);
nor U20104 (N_20104,N_19758,N_19755);
or U20105 (N_20105,N_19430,N_19247);
and U20106 (N_20106,N_19442,N_19782);
and U20107 (N_20107,N_19408,N_19698);
and U20108 (N_20108,N_19382,N_19546);
nand U20109 (N_20109,N_19533,N_19469);
nor U20110 (N_20110,N_19249,N_19602);
and U20111 (N_20111,N_19648,N_19296);
nor U20112 (N_20112,N_19781,N_19354);
nor U20113 (N_20113,N_19732,N_19457);
and U20114 (N_20114,N_19641,N_19784);
and U20115 (N_20115,N_19553,N_19556);
and U20116 (N_20116,N_19610,N_19422);
nor U20117 (N_20117,N_19439,N_19536);
nor U20118 (N_20118,N_19621,N_19430);
or U20119 (N_20119,N_19615,N_19731);
nor U20120 (N_20120,N_19436,N_19768);
or U20121 (N_20121,N_19502,N_19379);
and U20122 (N_20122,N_19452,N_19636);
nand U20123 (N_20123,N_19428,N_19560);
nor U20124 (N_20124,N_19628,N_19684);
and U20125 (N_20125,N_19409,N_19591);
or U20126 (N_20126,N_19537,N_19475);
nor U20127 (N_20127,N_19683,N_19310);
xnor U20128 (N_20128,N_19484,N_19771);
nand U20129 (N_20129,N_19651,N_19667);
nand U20130 (N_20130,N_19544,N_19484);
or U20131 (N_20131,N_19792,N_19275);
and U20132 (N_20132,N_19303,N_19253);
nor U20133 (N_20133,N_19677,N_19634);
nand U20134 (N_20134,N_19487,N_19218);
nor U20135 (N_20135,N_19684,N_19600);
and U20136 (N_20136,N_19435,N_19684);
nor U20137 (N_20137,N_19306,N_19345);
xor U20138 (N_20138,N_19329,N_19235);
xnor U20139 (N_20139,N_19545,N_19472);
nor U20140 (N_20140,N_19382,N_19448);
and U20141 (N_20141,N_19259,N_19738);
nor U20142 (N_20142,N_19716,N_19657);
nand U20143 (N_20143,N_19695,N_19315);
and U20144 (N_20144,N_19428,N_19472);
nand U20145 (N_20145,N_19310,N_19781);
xor U20146 (N_20146,N_19252,N_19506);
xnor U20147 (N_20147,N_19300,N_19579);
xnor U20148 (N_20148,N_19570,N_19771);
or U20149 (N_20149,N_19420,N_19415);
nand U20150 (N_20150,N_19297,N_19322);
or U20151 (N_20151,N_19727,N_19258);
and U20152 (N_20152,N_19612,N_19706);
xor U20153 (N_20153,N_19590,N_19726);
and U20154 (N_20154,N_19537,N_19332);
and U20155 (N_20155,N_19349,N_19351);
nand U20156 (N_20156,N_19466,N_19461);
nand U20157 (N_20157,N_19550,N_19457);
nor U20158 (N_20158,N_19459,N_19507);
nand U20159 (N_20159,N_19687,N_19479);
xnor U20160 (N_20160,N_19263,N_19444);
nand U20161 (N_20161,N_19556,N_19782);
nor U20162 (N_20162,N_19669,N_19775);
and U20163 (N_20163,N_19561,N_19786);
and U20164 (N_20164,N_19785,N_19464);
xnor U20165 (N_20165,N_19384,N_19410);
xnor U20166 (N_20166,N_19677,N_19599);
nor U20167 (N_20167,N_19393,N_19751);
or U20168 (N_20168,N_19711,N_19207);
and U20169 (N_20169,N_19475,N_19783);
and U20170 (N_20170,N_19230,N_19686);
nor U20171 (N_20171,N_19781,N_19248);
and U20172 (N_20172,N_19433,N_19237);
nor U20173 (N_20173,N_19782,N_19529);
nor U20174 (N_20174,N_19441,N_19562);
nand U20175 (N_20175,N_19489,N_19573);
nor U20176 (N_20176,N_19748,N_19610);
nand U20177 (N_20177,N_19721,N_19748);
and U20178 (N_20178,N_19457,N_19380);
xor U20179 (N_20179,N_19644,N_19419);
xnor U20180 (N_20180,N_19666,N_19404);
nor U20181 (N_20181,N_19757,N_19772);
nand U20182 (N_20182,N_19452,N_19522);
nor U20183 (N_20183,N_19755,N_19239);
and U20184 (N_20184,N_19712,N_19350);
nand U20185 (N_20185,N_19498,N_19419);
nand U20186 (N_20186,N_19444,N_19266);
nand U20187 (N_20187,N_19775,N_19419);
nand U20188 (N_20188,N_19684,N_19620);
nor U20189 (N_20189,N_19371,N_19345);
and U20190 (N_20190,N_19551,N_19224);
nand U20191 (N_20191,N_19274,N_19412);
nor U20192 (N_20192,N_19540,N_19277);
nand U20193 (N_20193,N_19589,N_19649);
nor U20194 (N_20194,N_19443,N_19463);
nand U20195 (N_20195,N_19596,N_19480);
xnor U20196 (N_20196,N_19721,N_19316);
and U20197 (N_20197,N_19313,N_19471);
nor U20198 (N_20198,N_19305,N_19719);
nor U20199 (N_20199,N_19437,N_19527);
nand U20200 (N_20200,N_19460,N_19545);
xnor U20201 (N_20201,N_19685,N_19253);
or U20202 (N_20202,N_19274,N_19223);
nand U20203 (N_20203,N_19418,N_19583);
nand U20204 (N_20204,N_19420,N_19271);
and U20205 (N_20205,N_19319,N_19717);
nor U20206 (N_20206,N_19223,N_19726);
nor U20207 (N_20207,N_19400,N_19532);
and U20208 (N_20208,N_19325,N_19339);
nor U20209 (N_20209,N_19393,N_19383);
nand U20210 (N_20210,N_19477,N_19679);
and U20211 (N_20211,N_19733,N_19444);
nand U20212 (N_20212,N_19230,N_19594);
nor U20213 (N_20213,N_19719,N_19691);
xnor U20214 (N_20214,N_19784,N_19455);
nand U20215 (N_20215,N_19211,N_19253);
nand U20216 (N_20216,N_19758,N_19539);
nand U20217 (N_20217,N_19598,N_19588);
nand U20218 (N_20218,N_19649,N_19393);
xnor U20219 (N_20219,N_19764,N_19275);
nand U20220 (N_20220,N_19390,N_19355);
and U20221 (N_20221,N_19331,N_19404);
nand U20222 (N_20222,N_19463,N_19531);
nand U20223 (N_20223,N_19684,N_19488);
and U20224 (N_20224,N_19618,N_19352);
and U20225 (N_20225,N_19300,N_19657);
or U20226 (N_20226,N_19666,N_19500);
nor U20227 (N_20227,N_19464,N_19488);
and U20228 (N_20228,N_19795,N_19783);
nand U20229 (N_20229,N_19323,N_19550);
and U20230 (N_20230,N_19390,N_19696);
and U20231 (N_20231,N_19332,N_19245);
and U20232 (N_20232,N_19603,N_19682);
and U20233 (N_20233,N_19541,N_19441);
nor U20234 (N_20234,N_19352,N_19387);
nor U20235 (N_20235,N_19721,N_19602);
nand U20236 (N_20236,N_19266,N_19283);
xor U20237 (N_20237,N_19286,N_19301);
nor U20238 (N_20238,N_19766,N_19285);
or U20239 (N_20239,N_19294,N_19743);
xnor U20240 (N_20240,N_19206,N_19233);
nand U20241 (N_20241,N_19282,N_19770);
and U20242 (N_20242,N_19715,N_19568);
and U20243 (N_20243,N_19734,N_19314);
and U20244 (N_20244,N_19550,N_19494);
or U20245 (N_20245,N_19282,N_19364);
nand U20246 (N_20246,N_19790,N_19709);
nor U20247 (N_20247,N_19501,N_19602);
xor U20248 (N_20248,N_19340,N_19643);
and U20249 (N_20249,N_19579,N_19683);
xnor U20250 (N_20250,N_19500,N_19384);
or U20251 (N_20251,N_19455,N_19556);
or U20252 (N_20252,N_19732,N_19674);
xnor U20253 (N_20253,N_19640,N_19513);
nor U20254 (N_20254,N_19253,N_19769);
xnor U20255 (N_20255,N_19729,N_19222);
nor U20256 (N_20256,N_19597,N_19314);
and U20257 (N_20257,N_19505,N_19513);
or U20258 (N_20258,N_19420,N_19793);
xnor U20259 (N_20259,N_19339,N_19688);
nand U20260 (N_20260,N_19633,N_19523);
or U20261 (N_20261,N_19470,N_19614);
nor U20262 (N_20262,N_19717,N_19251);
or U20263 (N_20263,N_19618,N_19624);
nor U20264 (N_20264,N_19421,N_19372);
nor U20265 (N_20265,N_19614,N_19398);
and U20266 (N_20266,N_19497,N_19725);
nor U20267 (N_20267,N_19585,N_19203);
nor U20268 (N_20268,N_19250,N_19564);
or U20269 (N_20269,N_19217,N_19300);
nand U20270 (N_20270,N_19551,N_19663);
nor U20271 (N_20271,N_19223,N_19293);
xnor U20272 (N_20272,N_19417,N_19768);
nor U20273 (N_20273,N_19292,N_19214);
nand U20274 (N_20274,N_19525,N_19793);
xnor U20275 (N_20275,N_19259,N_19315);
nand U20276 (N_20276,N_19392,N_19433);
xnor U20277 (N_20277,N_19651,N_19600);
or U20278 (N_20278,N_19716,N_19675);
and U20279 (N_20279,N_19715,N_19642);
or U20280 (N_20280,N_19622,N_19769);
and U20281 (N_20281,N_19651,N_19603);
nor U20282 (N_20282,N_19420,N_19210);
or U20283 (N_20283,N_19200,N_19532);
nor U20284 (N_20284,N_19602,N_19209);
and U20285 (N_20285,N_19279,N_19546);
or U20286 (N_20286,N_19660,N_19646);
nand U20287 (N_20287,N_19325,N_19204);
nor U20288 (N_20288,N_19220,N_19205);
and U20289 (N_20289,N_19700,N_19222);
and U20290 (N_20290,N_19545,N_19451);
xor U20291 (N_20291,N_19218,N_19216);
nor U20292 (N_20292,N_19593,N_19689);
nor U20293 (N_20293,N_19490,N_19406);
xnor U20294 (N_20294,N_19682,N_19695);
and U20295 (N_20295,N_19316,N_19408);
xor U20296 (N_20296,N_19723,N_19253);
nor U20297 (N_20297,N_19337,N_19215);
xor U20298 (N_20298,N_19576,N_19418);
xor U20299 (N_20299,N_19762,N_19602);
nand U20300 (N_20300,N_19296,N_19338);
nor U20301 (N_20301,N_19250,N_19350);
nand U20302 (N_20302,N_19512,N_19529);
nor U20303 (N_20303,N_19536,N_19282);
or U20304 (N_20304,N_19260,N_19746);
and U20305 (N_20305,N_19441,N_19252);
or U20306 (N_20306,N_19408,N_19668);
or U20307 (N_20307,N_19767,N_19382);
or U20308 (N_20308,N_19375,N_19257);
and U20309 (N_20309,N_19736,N_19719);
xnor U20310 (N_20310,N_19361,N_19524);
or U20311 (N_20311,N_19484,N_19448);
nor U20312 (N_20312,N_19379,N_19398);
or U20313 (N_20313,N_19657,N_19386);
nor U20314 (N_20314,N_19222,N_19490);
and U20315 (N_20315,N_19369,N_19766);
xnor U20316 (N_20316,N_19370,N_19719);
nand U20317 (N_20317,N_19777,N_19436);
or U20318 (N_20318,N_19202,N_19741);
nand U20319 (N_20319,N_19542,N_19283);
nor U20320 (N_20320,N_19319,N_19320);
xor U20321 (N_20321,N_19262,N_19355);
or U20322 (N_20322,N_19573,N_19311);
and U20323 (N_20323,N_19676,N_19591);
or U20324 (N_20324,N_19429,N_19597);
or U20325 (N_20325,N_19209,N_19413);
nor U20326 (N_20326,N_19382,N_19430);
xor U20327 (N_20327,N_19216,N_19348);
xor U20328 (N_20328,N_19501,N_19280);
or U20329 (N_20329,N_19309,N_19562);
and U20330 (N_20330,N_19601,N_19549);
nand U20331 (N_20331,N_19306,N_19310);
nand U20332 (N_20332,N_19554,N_19387);
and U20333 (N_20333,N_19278,N_19202);
nor U20334 (N_20334,N_19269,N_19304);
nand U20335 (N_20335,N_19464,N_19583);
nand U20336 (N_20336,N_19286,N_19420);
and U20337 (N_20337,N_19325,N_19226);
xnor U20338 (N_20338,N_19306,N_19588);
and U20339 (N_20339,N_19732,N_19330);
nor U20340 (N_20340,N_19767,N_19324);
and U20341 (N_20341,N_19759,N_19452);
or U20342 (N_20342,N_19505,N_19653);
and U20343 (N_20343,N_19408,N_19204);
or U20344 (N_20344,N_19751,N_19660);
and U20345 (N_20345,N_19295,N_19645);
and U20346 (N_20346,N_19792,N_19299);
and U20347 (N_20347,N_19728,N_19570);
nor U20348 (N_20348,N_19334,N_19622);
nand U20349 (N_20349,N_19442,N_19374);
xnor U20350 (N_20350,N_19497,N_19383);
nor U20351 (N_20351,N_19269,N_19546);
nand U20352 (N_20352,N_19482,N_19531);
and U20353 (N_20353,N_19455,N_19413);
xnor U20354 (N_20354,N_19443,N_19425);
and U20355 (N_20355,N_19387,N_19330);
and U20356 (N_20356,N_19223,N_19563);
nand U20357 (N_20357,N_19318,N_19517);
and U20358 (N_20358,N_19680,N_19308);
nand U20359 (N_20359,N_19475,N_19257);
or U20360 (N_20360,N_19789,N_19223);
nand U20361 (N_20361,N_19745,N_19459);
xnor U20362 (N_20362,N_19530,N_19203);
nor U20363 (N_20363,N_19278,N_19607);
or U20364 (N_20364,N_19485,N_19498);
xor U20365 (N_20365,N_19437,N_19263);
and U20366 (N_20366,N_19252,N_19421);
nor U20367 (N_20367,N_19523,N_19517);
or U20368 (N_20368,N_19220,N_19722);
xor U20369 (N_20369,N_19405,N_19302);
and U20370 (N_20370,N_19415,N_19485);
nor U20371 (N_20371,N_19380,N_19408);
nor U20372 (N_20372,N_19311,N_19487);
nand U20373 (N_20373,N_19354,N_19213);
or U20374 (N_20374,N_19367,N_19673);
xor U20375 (N_20375,N_19685,N_19442);
nand U20376 (N_20376,N_19560,N_19491);
or U20377 (N_20377,N_19543,N_19622);
and U20378 (N_20378,N_19538,N_19640);
nand U20379 (N_20379,N_19691,N_19320);
nand U20380 (N_20380,N_19435,N_19754);
or U20381 (N_20381,N_19437,N_19346);
xor U20382 (N_20382,N_19548,N_19740);
or U20383 (N_20383,N_19333,N_19465);
or U20384 (N_20384,N_19679,N_19271);
nand U20385 (N_20385,N_19776,N_19721);
and U20386 (N_20386,N_19491,N_19613);
or U20387 (N_20387,N_19449,N_19524);
xnor U20388 (N_20388,N_19538,N_19251);
nand U20389 (N_20389,N_19709,N_19529);
or U20390 (N_20390,N_19724,N_19528);
xnor U20391 (N_20391,N_19706,N_19777);
xnor U20392 (N_20392,N_19238,N_19217);
xor U20393 (N_20393,N_19742,N_19573);
xor U20394 (N_20394,N_19658,N_19220);
and U20395 (N_20395,N_19630,N_19797);
nand U20396 (N_20396,N_19388,N_19772);
and U20397 (N_20397,N_19296,N_19553);
nand U20398 (N_20398,N_19617,N_19250);
or U20399 (N_20399,N_19611,N_19253);
or U20400 (N_20400,N_20293,N_20084);
nor U20401 (N_20401,N_19955,N_19802);
nor U20402 (N_20402,N_20327,N_20281);
nor U20403 (N_20403,N_20344,N_19899);
xnor U20404 (N_20404,N_20081,N_20011);
nor U20405 (N_20405,N_20039,N_19906);
nor U20406 (N_20406,N_20192,N_20115);
and U20407 (N_20407,N_19979,N_19880);
and U20408 (N_20408,N_19877,N_20332);
nor U20409 (N_20409,N_20162,N_19915);
nor U20410 (N_20410,N_19984,N_20130);
nor U20411 (N_20411,N_19889,N_20204);
or U20412 (N_20412,N_20388,N_20376);
nor U20413 (N_20413,N_19865,N_20278);
or U20414 (N_20414,N_20315,N_20035);
nand U20415 (N_20415,N_20339,N_20156);
nand U20416 (N_20416,N_20172,N_20213);
nand U20417 (N_20417,N_19818,N_20124);
nor U20418 (N_20418,N_19909,N_19943);
nor U20419 (N_20419,N_20238,N_19828);
nand U20420 (N_20420,N_20045,N_19836);
or U20421 (N_20421,N_20225,N_20307);
and U20422 (N_20422,N_20228,N_20069);
nand U20423 (N_20423,N_20348,N_20230);
nand U20424 (N_20424,N_20032,N_19800);
and U20425 (N_20425,N_20209,N_20166);
and U20426 (N_20426,N_20159,N_19824);
or U20427 (N_20427,N_19840,N_19956);
xor U20428 (N_20428,N_20061,N_20294);
nor U20429 (N_20429,N_20272,N_19826);
xor U20430 (N_20430,N_19959,N_20181);
and U20431 (N_20431,N_20093,N_20302);
nand U20432 (N_20432,N_20029,N_19985);
or U20433 (N_20433,N_19991,N_19971);
xnor U20434 (N_20434,N_20211,N_20333);
or U20435 (N_20435,N_20023,N_20067);
or U20436 (N_20436,N_20167,N_20224);
or U20437 (N_20437,N_20105,N_20353);
nand U20438 (N_20438,N_20070,N_20231);
nand U20439 (N_20439,N_19813,N_20351);
nand U20440 (N_20440,N_20373,N_19910);
nand U20441 (N_20441,N_20132,N_20176);
xor U20442 (N_20442,N_19928,N_20384);
or U20443 (N_20443,N_20382,N_20013);
nor U20444 (N_20444,N_20169,N_19805);
xnor U20445 (N_20445,N_19849,N_20256);
nand U20446 (N_20446,N_20305,N_19966);
xor U20447 (N_20447,N_19975,N_20379);
xnor U20448 (N_20448,N_20273,N_19987);
or U20449 (N_20449,N_19812,N_20022);
and U20450 (N_20450,N_19963,N_19852);
or U20451 (N_20451,N_19839,N_20289);
and U20452 (N_20452,N_20180,N_20098);
xor U20453 (N_20453,N_20247,N_19986);
and U20454 (N_20454,N_20075,N_19886);
nor U20455 (N_20455,N_19990,N_20251);
xor U20456 (N_20456,N_20325,N_20129);
nor U20457 (N_20457,N_20354,N_20131);
nor U20458 (N_20458,N_20016,N_19933);
xor U20459 (N_20459,N_20168,N_20076);
xnor U20460 (N_20460,N_19875,N_20367);
or U20461 (N_20461,N_19831,N_20006);
or U20462 (N_20462,N_19902,N_20189);
or U20463 (N_20463,N_19923,N_20027);
nand U20464 (N_20464,N_20377,N_19919);
nor U20465 (N_20465,N_19938,N_19858);
and U20466 (N_20466,N_19892,N_20163);
xnor U20467 (N_20467,N_19816,N_20310);
nand U20468 (N_20468,N_20145,N_20242);
nand U20469 (N_20469,N_20057,N_20047);
nor U20470 (N_20470,N_20317,N_20255);
or U20471 (N_20471,N_20198,N_19854);
and U20472 (N_20472,N_20000,N_20316);
xnor U20473 (N_20473,N_20349,N_20195);
or U20474 (N_20474,N_20074,N_20106);
and U20475 (N_20475,N_20210,N_20308);
and U20476 (N_20476,N_20196,N_20234);
nor U20477 (N_20477,N_20345,N_20218);
xnor U20478 (N_20478,N_20018,N_20356);
xor U20479 (N_20479,N_20083,N_20346);
and U20480 (N_20480,N_19894,N_20220);
nor U20481 (N_20481,N_20341,N_20226);
nand U20482 (N_20482,N_20268,N_19900);
nand U20483 (N_20483,N_20236,N_20001);
or U20484 (N_20484,N_19873,N_20017);
nand U20485 (N_20485,N_20263,N_20393);
nand U20486 (N_20486,N_20313,N_20003);
and U20487 (N_20487,N_20138,N_20221);
or U20488 (N_20488,N_20337,N_20136);
or U20489 (N_20489,N_19890,N_20335);
xor U20490 (N_20490,N_20154,N_19842);
and U20491 (N_20491,N_19939,N_20298);
nand U20492 (N_20492,N_20383,N_20107);
xor U20493 (N_20493,N_20342,N_19860);
and U20494 (N_20494,N_20128,N_19898);
nor U20495 (N_20495,N_20068,N_20064);
nor U20496 (N_20496,N_20311,N_19859);
and U20497 (N_20497,N_20085,N_19926);
and U20498 (N_20498,N_20004,N_20222);
nand U20499 (N_20499,N_19870,N_20177);
nand U20500 (N_20500,N_20285,N_20365);
or U20501 (N_20501,N_19965,N_19825);
xor U20502 (N_20502,N_20215,N_19996);
or U20503 (N_20503,N_19885,N_20260);
nand U20504 (N_20504,N_20364,N_19827);
or U20505 (N_20505,N_19961,N_19801);
xnor U20506 (N_20506,N_20287,N_20157);
nor U20507 (N_20507,N_20126,N_19843);
and U20508 (N_20508,N_19822,N_20276);
xor U20509 (N_20509,N_20122,N_19871);
xnor U20510 (N_20510,N_19920,N_19989);
or U20511 (N_20511,N_20271,N_19935);
nor U20512 (N_20512,N_20030,N_20100);
nand U20513 (N_20513,N_20171,N_20261);
and U20514 (N_20514,N_20241,N_20253);
or U20515 (N_20515,N_20274,N_20229);
or U20516 (N_20516,N_20153,N_20051);
nor U20517 (N_20517,N_20060,N_19867);
xor U20518 (N_20518,N_20203,N_19911);
xor U20519 (N_20519,N_20088,N_19841);
xnor U20520 (N_20520,N_20329,N_19964);
and U20521 (N_20521,N_20270,N_19810);
nor U20522 (N_20522,N_19863,N_20205);
or U20523 (N_20523,N_20330,N_19887);
nand U20524 (N_20524,N_20063,N_19807);
or U20525 (N_20525,N_20217,N_20007);
and U20526 (N_20526,N_20186,N_20368);
or U20527 (N_20527,N_19969,N_20087);
and U20528 (N_20528,N_20043,N_19993);
or U20529 (N_20529,N_20277,N_20326);
and U20530 (N_20530,N_20385,N_19932);
or U20531 (N_20531,N_19878,N_19951);
or U20532 (N_20532,N_20080,N_20135);
nand U20533 (N_20533,N_19850,N_19952);
or U20534 (N_20534,N_19942,N_20362);
and U20535 (N_20535,N_20134,N_20331);
nand U20536 (N_20536,N_19838,N_20227);
nor U20537 (N_20537,N_20340,N_20086);
nor U20538 (N_20538,N_20321,N_19835);
nand U20539 (N_20539,N_20328,N_20071);
xor U20540 (N_20540,N_20359,N_20036);
or U20541 (N_20541,N_20301,N_20194);
nand U20542 (N_20542,N_20054,N_19853);
xor U20543 (N_20543,N_20355,N_20096);
nand U20544 (N_20544,N_20292,N_20279);
and U20545 (N_20545,N_20397,N_19982);
nand U20546 (N_20546,N_19917,N_20252);
nand U20547 (N_20547,N_20389,N_20002);
xor U20548 (N_20548,N_20258,N_19862);
xor U20549 (N_20549,N_20164,N_20319);
nand U20550 (N_20550,N_20077,N_19861);
nand U20551 (N_20551,N_19833,N_20232);
xnor U20552 (N_20552,N_19882,N_20173);
xor U20553 (N_20553,N_20140,N_20089);
nand U20554 (N_20554,N_19834,N_20020);
nor U20555 (N_20555,N_19820,N_20235);
or U20556 (N_20556,N_20121,N_19998);
and U20557 (N_20557,N_20314,N_20360);
and U20558 (N_20558,N_20304,N_19904);
xnor U20559 (N_20559,N_20248,N_20374);
and U20560 (N_20560,N_19874,N_20223);
nand U20561 (N_20561,N_19837,N_19888);
nor U20562 (N_20562,N_20207,N_20264);
xor U20563 (N_20563,N_19945,N_20378);
xor U20564 (N_20564,N_20299,N_20240);
xnor U20565 (N_20565,N_19829,N_20078);
or U20566 (N_20566,N_19972,N_19970);
and U20567 (N_20567,N_20320,N_19857);
nand U20568 (N_20568,N_20034,N_19905);
and U20569 (N_20569,N_19872,N_20296);
or U20570 (N_20570,N_20250,N_20275);
and U20571 (N_20571,N_19946,N_20357);
or U20572 (N_20572,N_20147,N_20245);
xnor U20573 (N_20573,N_20118,N_20111);
xnor U20574 (N_20574,N_19819,N_20033);
nor U20575 (N_20575,N_19927,N_19988);
and U20576 (N_20576,N_19949,N_19983);
and U20577 (N_20577,N_19958,N_20371);
nor U20578 (N_20578,N_19994,N_20101);
xor U20579 (N_20579,N_19846,N_20216);
or U20580 (N_20580,N_19922,N_20392);
nor U20581 (N_20581,N_20249,N_20246);
nand U20582 (N_20582,N_19941,N_19844);
xor U20583 (N_20583,N_20005,N_20175);
nand U20584 (N_20584,N_20363,N_20352);
nor U20585 (N_20585,N_20178,N_20055);
nor U20586 (N_20586,N_20062,N_19893);
and U20587 (N_20587,N_20323,N_20233);
xor U20588 (N_20588,N_19803,N_20148);
nand U20589 (N_20589,N_19821,N_20160);
nand U20590 (N_20590,N_20137,N_20391);
and U20591 (N_20591,N_19924,N_19895);
and U20592 (N_20592,N_20142,N_20318);
and U20593 (N_20593,N_20028,N_20193);
or U20594 (N_20594,N_19947,N_19903);
or U20595 (N_20595,N_20031,N_20095);
and U20596 (N_20596,N_19868,N_20021);
xor U20597 (N_20597,N_20297,N_20306);
and U20598 (N_20598,N_19916,N_20267);
and U20599 (N_20599,N_19879,N_19845);
nand U20600 (N_20600,N_19980,N_20380);
xnor U20601 (N_20601,N_19832,N_20197);
and U20602 (N_20602,N_19876,N_19976);
xor U20603 (N_20603,N_20208,N_19855);
nor U20604 (N_20604,N_19847,N_20091);
nand U20605 (N_20605,N_19891,N_20184);
nand U20606 (N_20606,N_19809,N_20394);
nor U20607 (N_20607,N_19974,N_19957);
nand U20608 (N_20608,N_20324,N_20026);
nand U20609 (N_20609,N_20219,N_20109);
and U20610 (N_20610,N_19954,N_20350);
or U20611 (N_20611,N_20312,N_19856);
and U20612 (N_20612,N_19973,N_19962);
xnor U20613 (N_20613,N_20361,N_19968);
nand U20614 (N_20614,N_20058,N_20014);
and U20615 (N_20615,N_19866,N_20262);
nand U20616 (N_20616,N_20119,N_20123);
nand U20617 (N_20617,N_19937,N_20120);
nand U20618 (N_20618,N_20288,N_20040);
xor U20619 (N_20619,N_19806,N_20052);
nand U20620 (N_20620,N_20049,N_19848);
xnor U20621 (N_20621,N_20127,N_19950);
nand U20622 (N_20622,N_20056,N_19977);
nor U20623 (N_20623,N_20008,N_19997);
or U20624 (N_20624,N_19804,N_19851);
nor U20625 (N_20625,N_19864,N_20165);
xnor U20626 (N_20626,N_20170,N_19934);
nand U20627 (N_20627,N_20200,N_20090);
and U20628 (N_20628,N_20125,N_20396);
or U20629 (N_20629,N_19830,N_20042);
xnor U20630 (N_20630,N_20010,N_20370);
xnor U20631 (N_20631,N_20102,N_20141);
nor U20632 (N_20632,N_20336,N_20239);
nor U20633 (N_20633,N_20265,N_19811);
nor U20634 (N_20634,N_20053,N_19918);
nor U20635 (N_20635,N_20338,N_20322);
nand U20636 (N_20636,N_20185,N_20202);
nor U20637 (N_20637,N_20290,N_20065);
nand U20638 (N_20638,N_19815,N_20369);
xor U20639 (N_20639,N_20399,N_20073);
and U20640 (N_20640,N_19960,N_20347);
xnor U20641 (N_20641,N_20072,N_20110);
nor U20642 (N_20642,N_20191,N_19999);
nor U20643 (N_20643,N_19914,N_19925);
nor U20644 (N_20644,N_19936,N_20206);
nand U20645 (N_20645,N_20190,N_20188);
and U20646 (N_20646,N_20015,N_19929);
nand U20647 (N_20647,N_20151,N_20187);
nor U20648 (N_20648,N_20097,N_20366);
nor U20649 (N_20649,N_19808,N_19948);
nor U20650 (N_20650,N_20254,N_19883);
xor U20651 (N_20651,N_20144,N_19940);
or U20652 (N_20652,N_20284,N_19967);
and U20653 (N_20653,N_20161,N_20183);
nand U20654 (N_20654,N_19913,N_20050);
xnor U20655 (N_20655,N_19931,N_19884);
and U20656 (N_20656,N_20243,N_19930);
and U20657 (N_20657,N_20266,N_20386);
nand U20658 (N_20658,N_20143,N_20291);
xnor U20659 (N_20659,N_20334,N_20113);
xor U20660 (N_20660,N_20112,N_19869);
nand U20661 (N_20661,N_20082,N_20182);
or U20662 (N_20662,N_20038,N_19978);
nand U20663 (N_20663,N_20024,N_20199);
nor U20664 (N_20664,N_20395,N_20092);
xor U20665 (N_20665,N_19901,N_20158);
nor U20666 (N_20666,N_20009,N_20300);
or U20667 (N_20667,N_20116,N_20103);
or U20668 (N_20668,N_20041,N_20398);
and U20669 (N_20669,N_19907,N_19995);
nand U20670 (N_20670,N_19814,N_20257);
xnor U20671 (N_20671,N_20133,N_19896);
xor U20672 (N_20672,N_20375,N_20048);
xor U20673 (N_20673,N_20139,N_20212);
nand U20674 (N_20674,N_19944,N_20286);
nand U20675 (N_20675,N_19817,N_20381);
or U20676 (N_20676,N_20019,N_20044);
and U20677 (N_20677,N_20201,N_20282);
nand U20678 (N_20678,N_19823,N_20104);
xnor U20679 (N_20679,N_20295,N_20390);
or U20680 (N_20680,N_20358,N_20343);
nand U20681 (N_20681,N_20214,N_20114);
xor U20682 (N_20682,N_20046,N_20309);
xnor U20683 (N_20683,N_20179,N_20283);
and U20684 (N_20684,N_20066,N_19953);
nor U20685 (N_20685,N_19908,N_20155);
nor U20686 (N_20686,N_20152,N_20387);
xor U20687 (N_20687,N_20037,N_20150);
nand U20688 (N_20688,N_20303,N_20146);
nor U20689 (N_20689,N_20117,N_19881);
and U20690 (N_20690,N_19897,N_20237);
nand U20691 (N_20691,N_20244,N_20094);
nand U20692 (N_20692,N_20372,N_20149);
or U20693 (N_20693,N_20012,N_20025);
nor U20694 (N_20694,N_20108,N_20099);
xor U20695 (N_20695,N_20079,N_19981);
and U20696 (N_20696,N_20059,N_19992);
nor U20697 (N_20697,N_20269,N_20174);
nand U20698 (N_20698,N_20280,N_19921);
or U20699 (N_20699,N_20259,N_19912);
or U20700 (N_20700,N_20093,N_19955);
or U20701 (N_20701,N_20287,N_20372);
xor U20702 (N_20702,N_19855,N_19842);
or U20703 (N_20703,N_19945,N_20003);
and U20704 (N_20704,N_20087,N_20030);
and U20705 (N_20705,N_20084,N_20244);
nor U20706 (N_20706,N_19934,N_19979);
xor U20707 (N_20707,N_19935,N_19848);
nand U20708 (N_20708,N_20002,N_19944);
or U20709 (N_20709,N_20283,N_19866);
nor U20710 (N_20710,N_20010,N_19976);
or U20711 (N_20711,N_20190,N_20269);
and U20712 (N_20712,N_20002,N_20135);
nand U20713 (N_20713,N_20145,N_20224);
nand U20714 (N_20714,N_19903,N_20157);
or U20715 (N_20715,N_19895,N_19879);
nand U20716 (N_20716,N_20269,N_19825);
nor U20717 (N_20717,N_19844,N_20151);
nor U20718 (N_20718,N_19884,N_20399);
nand U20719 (N_20719,N_19902,N_20171);
nor U20720 (N_20720,N_19846,N_20196);
nor U20721 (N_20721,N_19869,N_20277);
or U20722 (N_20722,N_20190,N_20051);
xor U20723 (N_20723,N_19876,N_20170);
nand U20724 (N_20724,N_20345,N_20222);
and U20725 (N_20725,N_20331,N_20276);
nor U20726 (N_20726,N_20032,N_20185);
xnor U20727 (N_20727,N_20084,N_19903);
and U20728 (N_20728,N_20159,N_20052);
nor U20729 (N_20729,N_20245,N_20210);
xor U20730 (N_20730,N_20228,N_20005);
nor U20731 (N_20731,N_19838,N_19918);
xnor U20732 (N_20732,N_20329,N_20208);
or U20733 (N_20733,N_19873,N_20166);
xor U20734 (N_20734,N_19865,N_19963);
xor U20735 (N_20735,N_20176,N_20031);
and U20736 (N_20736,N_20120,N_20059);
xnor U20737 (N_20737,N_20176,N_20084);
and U20738 (N_20738,N_20025,N_20010);
xor U20739 (N_20739,N_19946,N_20189);
nor U20740 (N_20740,N_20179,N_20012);
or U20741 (N_20741,N_20341,N_19864);
or U20742 (N_20742,N_19940,N_20350);
nand U20743 (N_20743,N_20326,N_20118);
and U20744 (N_20744,N_19935,N_20332);
nor U20745 (N_20745,N_20260,N_19888);
and U20746 (N_20746,N_20235,N_20385);
xor U20747 (N_20747,N_19808,N_19849);
xor U20748 (N_20748,N_19808,N_19912);
and U20749 (N_20749,N_20273,N_20281);
nor U20750 (N_20750,N_20258,N_20197);
xor U20751 (N_20751,N_20074,N_20310);
nor U20752 (N_20752,N_20357,N_20360);
and U20753 (N_20753,N_19885,N_20070);
xnor U20754 (N_20754,N_19933,N_19969);
nand U20755 (N_20755,N_19817,N_20118);
nand U20756 (N_20756,N_20024,N_19944);
xor U20757 (N_20757,N_20151,N_20055);
nor U20758 (N_20758,N_20122,N_20300);
and U20759 (N_20759,N_20134,N_20310);
xor U20760 (N_20760,N_19869,N_19937);
and U20761 (N_20761,N_20266,N_20341);
xnor U20762 (N_20762,N_20290,N_19972);
and U20763 (N_20763,N_20016,N_20200);
nor U20764 (N_20764,N_19870,N_20384);
xor U20765 (N_20765,N_19985,N_19873);
xnor U20766 (N_20766,N_20298,N_20100);
nor U20767 (N_20767,N_20029,N_20153);
or U20768 (N_20768,N_20251,N_20124);
nand U20769 (N_20769,N_20019,N_20064);
nor U20770 (N_20770,N_20165,N_19982);
nand U20771 (N_20771,N_20286,N_19827);
or U20772 (N_20772,N_20113,N_20093);
nand U20773 (N_20773,N_20217,N_19800);
and U20774 (N_20774,N_20026,N_20022);
or U20775 (N_20775,N_20098,N_20181);
and U20776 (N_20776,N_19950,N_20295);
xnor U20777 (N_20777,N_20323,N_19836);
nand U20778 (N_20778,N_20123,N_19911);
nand U20779 (N_20779,N_19895,N_20210);
nand U20780 (N_20780,N_19970,N_20013);
nand U20781 (N_20781,N_20224,N_20057);
nor U20782 (N_20782,N_20310,N_20059);
nand U20783 (N_20783,N_20378,N_20377);
and U20784 (N_20784,N_20068,N_19887);
and U20785 (N_20785,N_20111,N_20208);
xnor U20786 (N_20786,N_20036,N_19883);
xnor U20787 (N_20787,N_20285,N_20260);
or U20788 (N_20788,N_19885,N_20238);
or U20789 (N_20789,N_20167,N_19818);
and U20790 (N_20790,N_20219,N_20113);
xor U20791 (N_20791,N_19831,N_20313);
or U20792 (N_20792,N_19865,N_20043);
nand U20793 (N_20793,N_20199,N_20345);
nand U20794 (N_20794,N_20047,N_20210);
nor U20795 (N_20795,N_19889,N_19990);
and U20796 (N_20796,N_20270,N_20350);
xor U20797 (N_20797,N_19931,N_19928);
xnor U20798 (N_20798,N_20018,N_20291);
or U20799 (N_20799,N_20204,N_19890);
nor U20800 (N_20800,N_20061,N_20373);
or U20801 (N_20801,N_20304,N_20374);
xnor U20802 (N_20802,N_20128,N_19847);
nor U20803 (N_20803,N_19818,N_19847);
xnor U20804 (N_20804,N_20313,N_20195);
or U20805 (N_20805,N_20021,N_19975);
nor U20806 (N_20806,N_20288,N_19899);
nand U20807 (N_20807,N_19839,N_20271);
or U20808 (N_20808,N_19883,N_20320);
nor U20809 (N_20809,N_20101,N_20371);
or U20810 (N_20810,N_20058,N_20362);
and U20811 (N_20811,N_20286,N_20272);
xor U20812 (N_20812,N_19965,N_20083);
or U20813 (N_20813,N_20067,N_20277);
xnor U20814 (N_20814,N_20133,N_19813);
and U20815 (N_20815,N_20366,N_20233);
nor U20816 (N_20816,N_19827,N_20192);
nand U20817 (N_20817,N_19983,N_20256);
xnor U20818 (N_20818,N_20307,N_20383);
nand U20819 (N_20819,N_20168,N_20102);
xor U20820 (N_20820,N_20200,N_20168);
or U20821 (N_20821,N_20083,N_19940);
and U20822 (N_20822,N_20254,N_20223);
nand U20823 (N_20823,N_19813,N_19985);
nor U20824 (N_20824,N_20076,N_20277);
nor U20825 (N_20825,N_19976,N_20137);
and U20826 (N_20826,N_20268,N_20133);
nand U20827 (N_20827,N_20227,N_20345);
xnor U20828 (N_20828,N_20139,N_19839);
or U20829 (N_20829,N_20302,N_20073);
or U20830 (N_20830,N_20347,N_20240);
xnor U20831 (N_20831,N_20364,N_20036);
and U20832 (N_20832,N_20126,N_20019);
and U20833 (N_20833,N_19884,N_19851);
nor U20834 (N_20834,N_19836,N_20080);
nor U20835 (N_20835,N_20329,N_20263);
or U20836 (N_20836,N_20363,N_19823);
or U20837 (N_20837,N_20280,N_20089);
and U20838 (N_20838,N_20154,N_20077);
nand U20839 (N_20839,N_20350,N_20214);
or U20840 (N_20840,N_20174,N_19948);
nor U20841 (N_20841,N_19814,N_19846);
nor U20842 (N_20842,N_20354,N_20165);
xnor U20843 (N_20843,N_20226,N_19831);
or U20844 (N_20844,N_19865,N_20243);
xnor U20845 (N_20845,N_20190,N_20316);
nor U20846 (N_20846,N_19858,N_20254);
xnor U20847 (N_20847,N_20284,N_20213);
and U20848 (N_20848,N_20053,N_20300);
nand U20849 (N_20849,N_20254,N_20337);
and U20850 (N_20850,N_19831,N_19883);
or U20851 (N_20851,N_20094,N_20146);
nor U20852 (N_20852,N_20090,N_20103);
or U20853 (N_20853,N_20211,N_19842);
and U20854 (N_20854,N_20188,N_20185);
nor U20855 (N_20855,N_19818,N_20255);
nor U20856 (N_20856,N_19879,N_20020);
and U20857 (N_20857,N_20288,N_20039);
nand U20858 (N_20858,N_20070,N_20310);
xnor U20859 (N_20859,N_20051,N_20371);
nor U20860 (N_20860,N_19834,N_20158);
and U20861 (N_20861,N_20274,N_20234);
nand U20862 (N_20862,N_20012,N_20325);
and U20863 (N_20863,N_20353,N_19991);
nand U20864 (N_20864,N_20201,N_20288);
or U20865 (N_20865,N_20025,N_20017);
nand U20866 (N_20866,N_19935,N_20273);
xor U20867 (N_20867,N_20105,N_20015);
or U20868 (N_20868,N_20338,N_20091);
and U20869 (N_20869,N_20257,N_20366);
nand U20870 (N_20870,N_20391,N_20109);
and U20871 (N_20871,N_20029,N_20324);
nor U20872 (N_20872,N_20201,N_19944);
nand U20873 (N_20873,N_19899,N_19996);
nor U20874 (N_20874,N_19957,N_20116);
or U20875 (N_20875,N_20206,N_20301);
and U20876 (N_20876,N_20050,N_20191);
nor U20877 (N_20877,N_19999,N_19949);
or U20878 (N_20878,N_19936,N_20289);
nor U20879 (N_20879,N_20101,N_19985);
or U20880 (N_20880,N_19996,N_20337);
or U20881 (N_20881,N_19843,N_20094);
xor U20882 (N_20882,N_20371,N_20313);
nor U20883 (N_20883,N_19981,N_19813);
xnor U20884 (N_20884,N_20379,N_20167);
nor U20885 (N_20885,N_20399,N_20200);
nand U20886 (N_20886,N_19894,N_20025);
nor U20887 (N_20887,N_19949,N_20138);
and U20888 (N_20888,N_19960,N_20085);
xor U20889 (N_20889,N_20061,N_20162);
and U20890 (N_20890,N_20233,N_20185);
or U20891 (N_20891,N_20250,N_19970);
or U20892 (N_20892,N_20319,N_20225);
nor U20893 (N_20893,N_19997,N_20052);
nor U20894 (N_20894,N_20090,N_20089);
nor U20895 (N_20895,N_20220,N_20023);
nor U20896 (N_20896,N_19831,N_19921);
nor U20897 (N_20897,N_19833,N_19992);
or U20898 (N_20898,N_19816,N_19869);
and U20899 (N_20899,N_20136,N_20125);
xor U20900 (N_20900,N_20186,N_20029);
xor U20901 (N_20901,N_19962,N_20194);
nand U20902 (N_20902,N_20271,N_19844);
nor U20903 (N_20903,N_19910,N_20254);
nand U20904 (N_20904,N_19848,N_19866);
nand U20905 (N_20905,N_19809,N_19845);
nor U20906 (N_20906,N_20384,N_20156);
nand U20907 (N_20907,N_20062,N_20077);
and U20908 (N_20908,N_19835,N_20379);
nor U20909 (N_20909,N_20317,N_20103);
nand U20910 (N_20910,N_19858,N_19958);
xor U20911 (N_20911,N_19867,N_19998);
and U20912 (N_20912,N_20164,N_20140);
or U20913 (N_20913,N_20176,N_20392);
xor U20914 (N_20914,N_20371,N_20375);
nor U20915 (N_20915,N_19889,N_20091);
nor U20916 (N_20916,N_20107,N_20196);
nand U20917 (N_20917,N_19945,N_19993);
nand U20918 (N_20918,N_20328,N_20181);
and U20919 (N_20919,N_20373,N_20344);
or U20920 (N_20920,N_19833,N_19977);
xor U20921 (N_20921,N_20250,N_20384);
and U20922 (N_20922,N_19989,N_20340);
nor U20923 (N_20923,N_20350,N_20357);
xor U20924 (N_20924,N_20357,N_20270);
and U20925 (N_20925,N_20275,N_20178);
nand U20926 (N_20926,N_19890,N_19968);
nor U20927 (N_20927,N_20171,N_20243);
and U20928 (N_20928,N_20372,N_19883);
xor U20929 (N_20929,N_19832,N_19906);
xor U20930 (N_20930,N_20331,N_20307);
or U20931 (N_20931,N_20133,N_19978);
or U20932 (N_20932,N_20200,N_20035);
or U20933 (N_20933,N_19859,N_19932);
nor U20934 (N_20934,N_20201,N_20286);
nand U20935 (N_20935,N_20086,N_19975);
xnor U20936 (N_20936,N_20020,N_20075);
nor U20937 (N_20937,N_20332,N_19911);
xnor U20938 (N_20938,N_20389,N_20074);
nor U20939 (N_20939,N_19903,N_20082);
and U20940 (N_20940,N_19919,N_20262);
nand U20941 (N_20941,N_19908,N_20194);
and U20942 (N_20942,N_19970,N_20151);
nand U20943 (N_20943,N_20158,N_19804);
xnor U20944 (N_20944,N_19855,N_20303);
nand U20945 (N_20945,N_20380,N_20322);
xnor U20946 (N_20946,N_20283,N_20175);
nand U20947 (N_20947,N_20129,N_19837);
nand U20948 (N_20948,N_20039,N_20392);
xor U20949 (N_20949,N_20261,N_19976);
nand U20950 (N_20950,N_20232,N_19829);
or U20951 (N_20951,N_20163,N_20103);
nor U20952 (N_20952,N_19871,N_20137);
xor U20953 (N_20953,N_20116,N_19805);
and U20954 (N_20954,N_20368,N_20142);
nand U20955 (N_20955,N_19959,N_20239);
nand U20956 (N_20956,N_20170,N_20141);
nand U20957 (N_20957,N_20382,N_19866);
and U20958 (N_20958,N_20061,N_19825);
nand U20959 (N_20959,N_20226,N_20253);
and U20960 (N_20960,N_20199,N_20157);
or U20961 (N_20961,N_20127,N_20311);
and U20962 (N_20962,N_20148,N_20295);
nand U20963 (N_20963,N_20271,N_20384);
and U20964 (N_20964,N_20392,N_19978);
and U20965 (N_20965,N_19840,N_20105);
nand U20966 (N_20966,N_20167,N_20322);
xor U20967 (N_20967,N_19821,N_19801);
nand U20968 (N_20968,N_20309,N_19947);
xnor U20969 (N_20969,N_20096,N_20032);
xnor U20970 (N_20970,N_19946,N_20061);
or U20971 (N_20971,N_19925,N_20068);
or U20972 (N_20972,N_19829,N_20128);
nand U20973 (N_20973,N_19980,N_20379);
and U20974 (N_20974,N_20116,N_19971);
xnor U20975 (N_20975,N_20303,N_20151);
nor U20976 (N_20976,N_19979,N_20283);
nand U20977 (N_20977,N_20045,N_19890);
or U20978 (N_20978,N_20244,N_20007);
and U20979 (N_20979,N_20217,N_20271);
or U20980 (N_20980,N_20316,N_19818);
nor U20981 (N_20981,N_20120,N_20365);
xor U20982 (N_20982,N_19955,N_20376);
xor U20983 (N_20983,N_20153,N_20183);
xor U20984 (N_20984,N_19918,N_20062);
or U20985 (N_20985,N_19970,N_20070);
nand U20986 (N_20986,N_20147,N_19955);
xor U20987 (N_20987,N_19863,N_19984);
or U20988 (N_20988,N_20390,N_20285);
or U20989 (N_20989,N_20292,N_19953);
or U20990 (N_20990,N_19896,N_20382);
xnor U20991 (N_20991,N_20091,N_20249);
nand U20992 (N_20992,N_20152,N_20312);
and U20993 (N_20993,N_20006,N_19861);
nor U20994 (N_20994,N_19887,N_20120);
xor U20995 (N_20995,N_20388,N_20001);
nor U20996 (N_20996,N_19806,N_20111);
nor U20997 (N_20997,N_20392,N_20045);
nor U20998 (N_20998,N_20065,N_19968);
or U20999 (N_20999,N_19952,N_20131);
or U21000 (N_21000,N_20956,N_20899);
nor U21001 (N_21001,N_20888,N_20403);
nor U21002 (N_21002,N_20459,N_20949);
nand U21003 (N_21003,N_20487,N_20965);
or U21004 (N_21004,N_20767,N_20655);
or U21005 (N_21005,N_20642,N_20488);
xnor U21006 (N_21006,N_20740,N_20651);
nor U21007 (N_21007,N_20737,N_20747);
nor U21008 (N_21008,N_20451,N_20827);
xnor U21009 (N_21009,N_20952,N_20530);
nor U21010 (N_21010,N_20969,N_20863);
nand U21011 (N_21011,N_20817,N_20497);
nand U21012 (N_21012,N_20919,N_20445);
and U21013 (N_21013,N_20885,N_20839);
nand U21014 (N_21014,N_20677,N_20558);
nand U21015 (N_21015,N_20668,N_20473);
nand U21016 (N_21016,N_20407,N_20995);
or U21017 (N_21017,N_20743,N_20753);
nor U21018 (N_21018,N_20752,N_20734);
and U21019 (N_21019,N_20596,N_20970);
or U21020 (N_21020,N_20908,N_20667);
or U21021 (N_21021,N_20463,N_20462);
nand U21022 (N_21022,N_20957,N_20939);
and U21023 (N_21023,N_20953,N_20542);
nor U21024 (N_21024,N_20825,N_20793);
nand U21025 (N_21025,N_20537,N_20441);
xor U21026 (N_21026,N_20599,N_20664);
xnor U21027 (N_21027,N_20910,N_20516);
xor U21028 (N_21028,N_20418,N_20581);
xnor U21029 (N_21029,N_20590,N_20884);
nand U21030 (N_21030,N_20773,N_20517);
or U21031 (N_21031,N_20658,N_20615);
nor U21032 (N_21032,N_20679,N_20778);
nor U21033 (N_21033,N_20649,N_20751);
nand U21034 (N_21034,N_20733,N_20788);
or U21035 (N_21035,N_20727,N_20657);
nor U21036 (N_21036,N_20566,N_20836);
nand U21037 (N_21037,N_20573,N_20510);
nand U21038 (N_21038,N_20475,N_20474);
or U21039 (N_21039,N_20849,N_20898);
xnor U21040 (N_21040,N_20998,N_20992);
nand U21041 (N_21041,N_20728,N_20822);
or U21042 (N_21042,N_20812,N_20993);
and U21043 (N_21043,N_20963,N_20729);
nand U21044 (N_21044,N_20997,N_20500);
xnor U21045 (N_21045,N_20948,N_20868);
and U21046 (N_21046,N_20567,N_20521);
nor U21047 (N_21047,N_20821,N_20968);
nor U21048 (N_21048,N_20659,N_20961);
xor U21049 (N_21049,N_20433,N_20635);
nand U21050 (N_21050,N_20913,N_20643);
or U21051 (N_21051,N_20576,N_20860);
xnor U21052 (N_21052,N_20835,N_20414);
nor U21053 (N_21053,N_20833,N_20660);
and U21054 (N_21054,N_20632,N_20801);
or U21055 (N_21055,N_20617,N_20518);
xor U21056 (N_21056,N_20994,N_20757);
nand U21057 (N_21057,N_20719,N_20675);
and U21058 (N_21058,N_20597,N_20772);
or U21059 (N_21059,N_20620,N_20449);
and U21060 (N_21060,N_20569,N_20564);
nand U21061 (N_21061,N_20781,N_20831);
nand U21062 (N_21062,N_20670,N_20843);
xor U21063 (N_21063,N_20647,N_20689);
nor U21064 (N_21064,N_20830,N_20716);
nand U21065 (N_21065,N_20798,N_20935);
nand U21066 (N_21066,N_20857,N_20591);
or U21067 (N_21067,N_20535,N_20622);
xnor U21068 (N_21068,N_20905,N_20624);
xor U21069 (N_21069,N_20958,N_20946);
nor U21070 (N_21070,N_20945,N_20442);
nor U21071 (N_21071,N_20524,N_20749);
nor U21072 (N_21072,N_20425,N_20483);
and U21073 (N_21073,N_20858,N_20761);
and U21074 (N_21074,N_20400,N_20731);
or U21075 (N_21075,N_20654,N_20413);
and U21076 (N_21076,N_20648,N_20875);
xnor U21077 (N_21077,N_20979,N_20936);
nand U21078 (N_21078,N_20794,N_20560);
nand U21079 (N_21079,N_20437,N_20807);
and U21080 (N_21080,N_20603,N_20686);
nor U21081 (N_21081,N_20426,N_20577);
nor U21082 (N_21082,N_20411,N_20882);
or U21083 (N_21083,N_20528,N_20493);
and U21084 (N_21084,N_20850,N_20423);
or U21085 (N_21085,N_20894,N_20621);
xor U21086 (N_21086,N_20549,N_20937);
xnor U21087 (N_21087,N_20881,N_20691);
nand U21088 (N_21088,N_20420,N_20851);
nand U21089 (N_21089,N_20429,N_20787);
xnor U21090 (N_21090,N_20797,N_20763);
xor U21091 (N_21091,N_20819,N_20903);
or U21092 (N_21092,N_20906,N_20457);
or U21093 (N_21093,N_20924,N_20687);
nand U21094 (N_21094,N_20578,N_20934);
or U21095 (N_21095,N_20674,N_20570);
nand U21096 (N_21096,N_20783,N_20694);
xnor U21097 (N_21097,N_20893,N_20818);
nand U21098 (N_21098,N_20738,N_20550);
nor U21099 (N_21099,N_20450,N_20713);
or U21100 (N_21100,N_20813,N_20460);
nand U21101 (N_21101,N_20628,N_20703);
nor U21102 (N_21102,N_20816,N_20974);
xnor U21103 (N_21103,N_20792,N_20623);
xor U21104 (N_21104,N_20575,N_20726);
and U21105 (N_21105,N_20472,N_20593);
nor U21106 (N_21106,N_20556,N_20975);
xor U21107 (N_21107,N_20631,N_20741);
or U21108 (N_21108,N_20840,N_20532);
nor U21109 (N_21109,N_20874,N_20630);
nand U21110 (N_21110,N_20444,N_20774);
xnor U21111 (N_21111,N_20877,N_20718);
nor U21112 (N_21112,N_20533,N_20987);
nand U21113 (N_21113,N_20810,N_20984);
nor U21114 (N_21114,N_20522,N_20452);
nand U21115 (N_21115,N_20436,N_20955);
nor U21116 (N_21116,N_20847,N_20465);
xnor U21117 (N_21117,N_20904,N_20525);
or U21118 (N_21118,N_20534,N_20769);
nand U21119 (N_21119,N_20896,N_20795);
nor U21120 (N_21120,N_20468,N_20653);
xnor U21121 (N_21121,N_20768,N_20775);
nand U21122 (N_21122,N_20824,N_20770);
and U21123 (N_21123,N_20732,N_20431);
xor U21124 (N_21124,N_20496,N_20940);
nand U21125 (N_21125,N_20714,N_20607);
and U21126 (N_21126,N_20477,N_20614);
nor U21127 (N_21127,N_20717,N_20501);
and U21128 (N_21128,N_20688,N_20705);
xnor U21129 (N_21129,N_20921,N_20920);
and U21130 (N_21130,N_20941,N_20582);
nor U21131 (N_21131,N_20478,N_20618);
nand U21132 (N_21132,N_20455,N_20848);
nand U21133 (N_21133,N_20644,N_20683);
nor U21134 (N_21134,N_20744,N_20990);
or U21135 (N_21135,N_20922,N_20739);
xor U21136 (N_21136,N_20480,N_20595);
nand U21137 (N_21137,N_20439,N_20467);
xnor U21138 (N_21138,N_20484,N_20799);
and U21139 (N_21139,N_20514,N_20708);
and U21140 (N_21140,N_20639,N_20986);
nor U21141 (N_21141,N_20855,N_20861);
nand U21142 (N_21142,N_20856,N_20704);
xor U21143 (N_21143,N_20585,N_20806);
and U21144 (N_21144,N_20665,N_20443);
or U21145 (N_21145,N_20434,N_20417);
nor U21146 (N_21146,N_20765,N_20976);
nand U21147 (N_21147,N_20927,N_20545);
nor U21148 (N_21148,N_20890,N_20762);
nand U21149 (N_21149,N_20959,N_20917);
nor U21150 (N_21150,N_20492,N_20912);
or U21151 (N_21151,N_20634,N_20693);
nor U21152 (N_21152,N_20479,N_20470);
xnor U21153 (N_21153,N_20780,N_20918);
xor U21154 (N_21154,N_20766,N_20458);
nor U21155 (N_21155,N_20754,N_20938);
nor U21156 (N_21156,N_20489,N_20523);
xnor U21157 (N_21157,N_20610,N_20779);
or U21158 (N_21158,N_20402,N_20950);
nand U21159 (N_21159,N_20989,N_20901);
or U21160 (N_21160,N_20823,N_20419);
nor U21161 (N_21161,N_20561,N_20867);
xnor U21162 (N_21162,N_20844,N_20645);
or U21163 (N_21163,N_20876,N_20422);
or U21164 (N_21164,N_20435,N_20711);
or U21165 (N_21165,N_20800,N_20404);
and U21166 (N_21166,N_20791,N_20415);
or U21167 (N_21167,N_20854,N_20692);
nand U21168 (N_21168,N_20656,N_20509);
or U21169 (N_21169,N_20699,N_20897);
and U21170 (N_21170,N_20942,N_20671);
or U21171 (N_21171,N_20784,N_20482);
or U21172 (N_21172,N_20672,N_20895);
and U21173 (N_21173,N_20865,N_20789);
or U21174 (N_21174,N_20606,N_20702);
nand U21175 (N_21175,N_20495,N_20902);
nand U21176 (N_21176,N_20446,N_20641);
xnor U21177 (N_21177,N_20598,N_20837);
nor U21178 (N_21178,N_20814,N_20464);
or U21179 (N_21179,N_20829,N_20580);
nor U21180 (N_21180,N_20915,N_20796);
or U21181 (N_21181,N_20828,N_20662);
xnor U21182 (N_21182,N_20682,N_20512);
nand U21183 (N_21183,N_20834,N_20421);
and U21184 (N_21184,N_20612,N_20503);
xnor U21185 (N_21185,N_20553,N_20730);
xnor U21186 (N_21186,N_20526,N_20491);
or U21187 (N_21187,N_20494,N_20572);
xnor U21188 (N_21188,N_20954,N_20646);
xnor U21189 (N_21189,N_20709,N_20605);
nand U21190 (N_21190,N_20430,N_20967);
or U21191 (N_21191,N_20758,N_20878);
and U21192 (N_21192,N_20625,N_20506);
or U21193 (N_21193,N_20760,N_20406);
nor U21194 (N_21194,N_20519,N_20755);
nor U21195 (N_21195,N_20771,N_20454);
and U21196 (N_21196,N_20539,N_20568);
xor U21197 (N_21197,N_20685,N_20600);
xor U21198 (N_21198,N_20589,N_20914);
and U21199 (N_21199,N_20759,N_20476);
nand U21200 (N_21200,N_20579,N_20978);
xnor U21201 (N_21201,N_20527,N_20808);
nor U21202 (N_21202,N_20438,N_20410);
nor U21203 (N_21203,N_20681,N_20706);
xor U21204 (N_21204,N_20619,N_20669);
xor U21205 (N_21205,N_20985,N_20932);
xor U21206 (N_21206,N_20424,N_20627);
nor U21207 (N_21207,N_20661,N_20983);
xnor U21208 (N_21208,N_20973,N_20574);
or U21209 (N_21209,N_20637,N_20636);
xor U21210 (N_21210,N_20826,N_20991);
xnor U21211 (N_21211,N_20611,N_20412);
or U21212 (N_21212,N_20745,N_20925);
or U21213 (N_21213,N_20832,N_20604);
nand U21214 (N_21214,N_20852,N_20548);
nand U21215 (N_21215,N_20933,N_20736);
xor U21216 (N_21216,N_20988,N_20531);
xnor U21217 (N_21217,N_20947,N_20887);
nor U21218 (N_21218,N_20584,N_20962);
nor U21219 (N_21219,N_20432,N_20698);
xor U21220 (N_21220,N_20841,N_20690);
or U21221 (N_21221,N_20499,N_20427);
xor U21222 (N_21222,N_20866,N_20859);
xor U21223 (N_21223,N_20507,N_20715);
xor U21224 (N_21224,N_20815,N_20790);
nand U21225 (N_21225,N_20802,N_20809);
nor U21226 (N_21226,N_20536,N_20724);
and U21227 (N_21227,N_20701,N_20498);
xnor U21228 (N_21228,N_20972,N_20873);
or U21229 (N_21229,N_20552,N_20466);
nand U21230 (N_21230,N_20696,N_20633);
nand U21231 (N_21231,N_20588,N_20416);
xnor U21232 (N_21232,N_20871,N_20471);
or U21233 (N_21233,N_20504,N_20999);
xnor U21234 (N_21234,N_20544,N_20695);
or U21235 (N_21235,N_20864,N_20508);
xor U21236 (N_21236,N_20891,N_20944);
xor U21237 (N_21237,N_20721,N_20461);
nor U21238 (N_21238,N_20486,N_20511);
nand U21239 (N_21239,N_20966,N_20629);
nor U21240 (N_21240,N_20401,N_20543);
nor U21241 (N_21241,N_20723,N_20602);
and U21242 (N_21242,N_20481,N_20587);
nand U21243 (N_21243,N_20928,N_20909);
nand U21244 (N_21244,N_20777,N_20640);
nor U21245 (N_21245,N_20879,N_20663);
nor U21246 (N_21246,N_20929,N_20538);
nand U21247 (N_21247,N_20870,N_20931);
nand U21248 (N_21248,N_20448,N_20756);
or U21249 (N_21249,N_20892,N_20559);
nand U21250 (N_21250,N_20977,N_20613);
xnor U21251 (N_21251,N_20546,N_20529);
or U21252 (N_21252,N_20785,N_20565);
nor U21253 (N_21253,N_20786,N_20750);
nand U21254 (N_21254,N_20811,N_20409);
xnor U21255 (N_21255,N_20926,N_20886);
xnor U21256 (N_21256,N_20916,N_20742);
nor U21257 (N_21257,N_20846,N_20697);
nand U21258 (N_21258,N_20626,N_20900);
nand U21259 (N_21259,N_20700,N_20601);
nor U21260 (N_21260,N_20554,N_20453);
xor U21261 (N_21261,N_20562,N_20680);
nor U21262 (N_21262,N_20880,N_20485);
xor U21263 (N_21263,N_20666,N_20515);
xnor U21264 (N_21264,N_20776,N_20505);
nor U21265 (N_21265,N_20638,N_20720);
and U21266 (N_21266,N_20712,N_20735);
nand U21267 (N_21267,N_20583,N_20490);
nand U21268 (N_21268,N_20803,N_20405);
or U21269 (N_21269,N_20609,N_20447);
or U21270 (N_21270,N_20862,N_20456);
nor U21271 (N_21271,N_20555,N_20502);
and U21272 (N_21272,N_20673,N_20520);
xnor U21273 (N_21273,N_20980,N_20845);
xnor U21274 (N_21274,N_20676,N_20746);
and U21275 (N_21275,N_20592,N_20748);
nor U21276 (N_21276,N_20764,N_20820);
nand U21277 (N_21277,N_20594,N_20838);
nor U21278 (N_21278,N_20571,N_20541);
nor U21279 (N_21279,N_20557,N_20684);
nor U21280 (N_21280,N_20869,N_20616);
nor U21281 (N_21281,N_20678,N_20540);
and U21282 (N_21282,N_20586,N_20911);
or U21283 (N_21283,N_20960,N_20513);
nor U21284 (N_21284,N_20971,N_20996);
or U21285 (N_21285,N_20440,N_20842);
and U21286 (N_21286,N_20652,N_20408);
or U21287 (N_21287,N_20982,N_20853);
nand U21288 (N_21288,N_20951,N_20428);
or U21289 (N_21289,N_20889,N_20883);
nor U21290 (N_21290,N_20722,N_20608);
or U21291 (N_21291,N_20710,N_20872);
xnor U21292 (N_21292,N_20547,N_20907);
or U21293 (N_21293,N_20650,N_20725);
nand U21294 (N_21294,N_20805,N_20943);
nor U21295 (N_21295,N_20930,N_20923);
and U21296 (N_21296,N_20981,N_20469);
nor U21297 (N_21297,N_20804,N_20707);
nand U21298 (N_21298,N_20563,N_20551);
or U21299 (N_21299,N_20964,N_20782);
and U21300 (N_21300,N_20551,N_20666);
xnor U21301 (N_21301,N_20770,N_20817);
and U21302 (N_21302,N_20401,N_20818);
nor U21303 (N_21303,N_20899,N_20428);
xor U21304 (N_21304,N_20708,N_20959);
xnor U21305 (N_21305,N_20630,N_20963);
and U21306 (N_21306,N_20898,N_20894);
nand U21307 (N_21307,N_20690,N_20788);
or U21308 (N_21308,N_20874,N_20606);
xor U21309 (N_21309,N_20770,N_20726);
and U21310 (N_21310,N_20543,N_20882);
nor U21311 (N_21311,N_20571,N_20404);
nand U21312 (N_21312,N_20689,N_20535);
or U21313 (N_21313,N_20813,N_20455);
nand U21314 (N_21314,N_20436,N_20570);
nor U21315 (N_21315,N_20774,N_20668);
and U21316 (N_21316,N_20876,N_20628);
nand U21317 (N_21317,N_20747,N_20676);
or U21318 (N_21318,N_20735,N_20552);
nor U21319 (N_21319,N_20510,N_20890);
or U21320 (N_21320,N_20771,N_20706);
xor U21321 (N_21321,N_20621,N_20599);
and U21322 (N_21322,N_20666,N_20462);
nand U21323 (N_21323,N_20455,N_20899);
nand U21324 (N_21324,N_20671,N_20453);
or U21325 (N_21325,N_20506,N_20667);
nand U21326 (N_21326,N_20418,N_20728);
or U21327 (N_21327,N_20430,N_20571);
xor U21328 (N_21328,N_20856,N_20760);
and U21329 (N_21329,N_20717,N_20693);
or U21330 (N_21330,N_20800,N_20732);
or U21331 (N_21331,N_20964,N_20520);
and U21332 (N_21332,N_20477,N_20858);
or U21333 (N_21333,N_20991,N_20773);
and U21334 (N_21334,N_20893,N_20618);
or U21335 (N_21335,N_20584,N_20424);
nor U21336 (N_21336,N_20949,N_20425);
xnor U21337 (N_21337,N_20839,N_20756);
and U21338 (N_21338,N_20437,N_20900);
or U21339 (N_21339,N_20851,N_20414);
xnor U21340 (N_21340,N_20404,N_20708);
nand U21341 (N_21341,N_20573,N_20713);
nand U21342 (N_21342,N_20974,N_20860);
nand U21343 (N_21343,N_20584,N_20963);
nand U21344 (N_21344,N_20926,N_20928);
and U21345 (N_21345,N_20550,N_20749);
nor U21346 (N_21346,N_20706,N_20945);
or U21347 (N_21347,N_20700,N_20977);
xor U21348 (N_21348,N_20905,N_20629);
nor U21349 (N_21349,N_20805,N_20537);
nor U21350 (N_21350,N_20863,N_20935);
nand U21351 (N_21351,N_20969,N_20834);
or U21352 (N_21352,N_20946,N_20631);
nand U21353 (N_21353,N_20891,N_20458);
nor U21354 (N_21354,N_20456,N_20813);
and U21355 (N_21355,N_20888,N_20529);
nor U21356 (N_21356,N_20750,N_20723);
and U21357 (N_21357,N_20500,N_20743);
nor U21358 (N_21358,N_20672,N_20453);
or U21359 (N_21359,N_20598,N_20933);
nand U21360 (N_21360,N_20964,N_20928);
xor U21361 (N_21361,N_20712,N_20625);
nand U21362 (N_21362,N_20519,N_20535);
xnor U21363 (N_21363,N_20582,N_20932);
nor U21364 (N_21364,N_20440,N_20672);
xor U21365 (N_21365,N_20873,N_20556);
nand U21366 (N_21366,N_20819,N_20859);
or U21367 (N_21367,N_20719,N_20756);
nand U21368 (N_21368,N_20712,N_20788);
xnor U21369 (N_21369,N_20423,N_20511);
or U21370 (N_21370,N_20667,N_20689);
nor U21371 (N_21371,N_20980,N_20569);
nand U21372 (N_21372,N_20492,N_20482);
nand U21373 (N_21373,N_20417,N_20549);
and U21374 (N_21374,N_20425,N_20662);
nor U21375 (N_21375,N_20967,N_20688);
nand U21376 (N_21376,N_20665,N_20942);
nor U21377 (N_21377,N_20944,N_20767);
nand U21378 (N_21378,N_20765,N_20653);
or U21379 (N_21379,N_20620,N_20790);
or U21380 (N_21380,N_20687,N_20917);
or U21381 (N_21381,N_20985,N_20937);
xnor U21382 (N_21382,N_20690,N_20974);
nand U21383 (N_21383,N_20413,N_20700);
or U21384 (N_21384,N_20475,N_20916);
and U21385 (N_21385,N_20606,N_20832);
or U21386 (N_21386,N_20462,N_20750);
and U21387 (N_21387,N_20585,N_20917);
and U21388 (N_21388,N_20688,N_20975);
and U21389 (N_21389,N_20847,N_20437);
nand U21390 (N_21390,N_20857,N_20872);
or U21391 (N_21391,N_20583,N_20411);
xnor U21392 (N_21392,N_20728,N_20722);
xor U21393 (N_21393,N_20478,N_20583);
nor U21394 (N_21394,N_20761,N_20588);
nand U21395 (N_21395,N_20423,N_20862);
nor U21396 (N_21396,N_20855,N_20991);
xnor U21397 (N_21397,N_20700,N_20948);
xor U21398 (N_21398,N_20568,N_20791);
xor U21399 (N_21399,N_20505,N_20939);
and U21400 (N_21400,N_20854,N_20988);
nand U21401 (N_21401,N_20798,N_20714);
nand U21402 (N_21402,N_20590,N_20403);
or U21403 (N_21403,N_20684,N_20871);
and U21404 (N_21404,N_20696,N_20993);
nor U21405 (N_21405,N_20471,N_20413);
nand U21406 (N_21406,N_20962,N_20447);
nor U21407 (N_21407,N_20813,N_20899);
nand U21408 (N_21408,N_20618,N_20939);
or U21409 (N_21409,N_20499,N_20697);
nor U21410 (N_21410,N_20475,N_20785);
nand U21411 (N_21411,N_20615,N_20574);
nor U21412 (N_21412,N_20744,N_20752);
nand U21413 (N_21413,N_20485,N_20939);
nor U21414 (N_21414,N_20773,N_20514);
xor U21415 (N_21415,N_20679,N_20713);
and U21416 (N_21416,N_20563,N_20950);
or U21417 (N_21417,N_20682,N_20755);
and U21418 (N_21418,N_20850,N_20616);
nor U21419 (N_21419,N_20623,N_20833);
and U21420 (N_21420,N_20771,N_20893);
xnor U21421 (N_21421,N_20708,N_20557);
or U21422 (N_21422,N_20444,N_20710);
nor U21423 (N_21423,N_20914,N_20856);
and U21424 (N_21424,N_20661,N_20868);
xor U21425 (N_21425,N_20978,N_20703);
or U21426 (N_21426,N_20920,N_20643);
xnor U21427 (N_21427,N_20990,N_20768);
or U21428 (N_21428,N_20732,N_20763);
or U21429 (N_21429,N_20653,N_20831);
and U21430 (N_21430,N_20543,N_20503);
nor U21431 (N_21431,N_20917,N_20895);
and U21432 (N_21432,N_20625,N_20692);
nand U21433 (N_21433,N_20813,N_20596);
and U21434 (N_21434,N_20874,N_20998);
xnor U21435 (N_21435,N_20848,N_20866);
xor U21436 (N_21436,N_20997,N_20617);
nand U21437 (N_21437,N_20734,N_20851);
nand U21438 (N_21438,N_20788,N_20725);
xor U21439 (N_21439,N_20568,N_20979);
nand U21440 (N_21440,N_20401,N_20757);
nand U21441 (N_21441,N_20820,N_20969);
xnor U21442 (N_21442,N_20635,N_20920);
or U21443 (N_21443,N_20604,N_20652);
nor U21444 (N_21444,N_20911,N_20977);
xnor U21445 (N_21445,N_20509,N_20694);
or U21446 (N_21446,N_20562,N_20849);
nor U21447 (N_21447,N_20689,N_20448);
xnor U21448 (N_21448,N_20793,N_20950);
or U21449 (N_21449,N_20438,N_20450);
or U21450 (N_21450,N_20753,N_20983);
and U21451 (N_21451,N_20470,N_20790);
and U21452 (N_21452,N_20538,N_20923);
nand U21453 (N_21453,N_20673,N_20463);
xor U21454 (N_21454,N_20841,N_20563);
nand U21455 (N_21455,N_20555,N_20593);
xor U21456 (N_21456,N_20460,N_20829);
xnor U21457 (N_21457,N_20927,N_20914);
nor U21458 (N_21458,N_20986,N_20697);
nand U21459 (N_21459,N_20556,N_20439);
and U21460 (N_21460,N_20814,N_20901);
nand U21461 (N_21461,N_20877,N_20762);
xnor U21462 (N_21462,N_20714,N_20864);
nor U21463 (N_21463,N_20897,N_20974);
and U21464 (N_21464,N_20621,N_20463);
xor U21465 (N_21465,N_20535,N_20668);
and U21466 (N_21466,N_20506,N_20430);
xor U21467 (N_21467,N_20678,N_20994);
and U21468 (N_21468,N_20546,N_20953);
and U21469 (N_21469,N_20996,N_20521);
nand U21470 (N_21470,N_20513,N_20492);
or U21471 (N_21471,N_20914,N_20562);
or U21472 (N_21472,N_20780,N_20460);
nand U21473 (N_21473,N_20939,N_20436);
nand U21474 (N_21474,N_20939,N_20938);
and U21475 (N_21475,N_20918,N_20478);
or U21476 (N_21476,N_20400,N_20704);
and U21477 (N_21477,N_20608,N_20486);
and U21478 (N_21478,N_20518,N_20555);
xor U21479 (N_21479,N_20474,N_20703);
xor U21480 (N_21480,N_20956,N_20693);
or U21481 (N_21481,N_20716,N_20923);
nor U21482 (N_21482,N_20779,N_20776);
and U21483 (N_21483,N_20795,N_20882);
or U21484 (N_21484,N_20833,N_20647);
and U21485 (N_21485,N_20937,N_20593);
or U21486 (N_21486,N_20857,N_20475);
xor U21487 (N_21487,N_20401,N_20876);
and U21488 (N_21488,N_20840,N_20721);
xor U21489 (N_21489,N_20940,N_20624);
or U21490 (N_21490,N_20850,N_20915);
or U21491 (N_21491,N_20898,N_20491);
xnor U21492 (N_21492,N_20737,N_20575);
nor U21493 (N_21493,N_20782,N_20722);
or U21494 (N_21494,N_20541,N_20674);
xnor U21495 (N_21495,N_20453,N_20597);
nor U21496 (N_21496,N_20449,N_20430);
nor U21497 (N_21497,N_20456,N_20466);
nor U21498 (N_21498,N_20897,N_20879);
nor U21499 (N_21499,N_20541,N_20700);
and U21500 (N_21500,N_20643,N_20591);
and U21501 (N_21501,N_20498,N_20995);
xor U21502 (N_21502,N_20646,N_20999);
or U21503 (N_21503,N_20499,N_20669);
nor U21504 (N_21504,N_20419,N_20940);
nand U21505 (N_21505,N_20645,N_20793);
nor U21506 (N_21506,N_20444,N_20775);
xor U21507 (N_21507,N_20704,N_20697);
nand U21508 (N_21508,N_20907,N_20731);
or U21509 (N_21509,N_20649,N_20834);
nor U21510 (N_21510,N_20858,N_20989);
xnor U21511 (N_21511,N_20603,N_20951);
nand U21512 (N_21512,N_20960,N_20853);
nor U21513 (N_21513,N_20500,N_20557);
xor U21514 (N_21514,N_20668,N_20708);
and U21515 (N_21515,N_20474,N_20674);
xnor U21516 (N_21516,N_20957,N_20434);
or U21517 (N_21517,N_20789,N_20602);
or U21518 (N_21518,N_20499,N_20522);
and U21519 (N_21519,N_20471,N_20462);
xor U21520 (N_21520,N_20602,N_20641);
nor U21521 (N_21521,N_20747,N_20799);
and U21522 (N_21522,N_20966,N_20797);
and U21523 (N_21523,N_20954,N_20707);
and U21524 (N_21524,N_20747,N_20970);
nand U21525 (N_21525,N_20629,N_20615);
or U21526 (N_21526,N_20454,N_20497);
nand U21527 (N_21527,N_20503,N_20836);
nand U21528 (N_21528,N_20968,N_20629);
nand U21529 (N_21529,N_20500,N_20463);
and U21530 (N_21530,N_20463,N_20654);
nor U21531 (N_21531,N_20444,N_20670);
or U21532 (N_21532,N_20919,N_20972);
and U21533 (N_21533,N_20671,N_20592);
xnor U21534 (N_21534,N_20611,N_20919);
and U21535 (N_21535,N_20424,N_20637);
xnor U21536 (N_21536,N_20505,N_20855);
xor U21537 (N_21537,N_20411,N_20409);
nand U21538 (N_21538,N_20609,N_20855);
and U21539 (N_21539,N_20432,N_20575);
and U21540 (N_21540,N_20993,N_20871);
nor U21541 (N_21541,N_20761,N_20692);
and U21542 (N_21542,N_20423,N_20771);
xor U21543 (N_21543,N_20694,N_20865);
nor U21544 (N_21544,N_20628,N_20967);
nand U21545 (N_21545,N_20950,N_20592);
or U21546 (N_21546,N_20523,N_20788);
xnor U21547 (N_21547,N_20690,N_20860);
xnor U21548 (N_21548,N_20657,N_20827);
or U21549 (N_21549,N_20962,N_20903);
and U21550 (N_21550,N_20865,N_20506);
and U21551 (N_21551,N_20791,N_20498);
or U21552 (N_21552,N_20431,N_20836);
xor U21553 (N_21553,N_20936,N_20582);
xor U21554 (N_21554,N_20805,N_20627);
nand U21555 (N_21555,N_20670,N_20600);
nor U21556 (N_21556,N_20837,N_20799);
xor U21557 (N_21557,N_20985,N_20859);
and U21558 (N_21558,N_20933,N_20588);
xor U21559 (N_21559,N_20598,N_20722);
nor U21560 (N_21560,N_20599,N_20979);
xnor U21561 (N_21561,N_20868,N_20784);
nor U21562 (N_21562,N_20672,N_20595);
and U21563 (N_21563,N_20754,N_20663);
nor U21564 (N_21564,N_20709,N_20940);
xnor U21565 (N_21565,N_20973,N_20480);
nand U21566 (N_21566,N_20652,N_20574);
and U21567 (N_21567,N_20512,N_20953);
or U21568 (N_21568,N_20767,N_20968);
nand U21569 (N_21569,N_20567,N_20944);
nand U21570 (N_21570,N_20717,N_20910);
and U21571 (N_21571,N_20947,N_20464);
nand U21572 (N_21572,N_20408,N_20546);
nor U21573 (N_21573,N_20767,N_20741);
nand U21574 (N_21574,N_20593,N_20539);
and U21575 (N_21575,N_20549,N_20828);
or U21576 (N_21576,N_20705,N_20626);
xor U21577 (N_21577,N_20436,N_20789);
nor U21578 (N_21578,N_20680,N_20724);
nor U21579 (N_21579,N_20876,N_20666);
xor U21580 (N_21580,N_20680,N_20648);
nor U21581 (N_21581,N_20879,N_20480);
and U21582 (N_21582,N_20729,N_20921);
or U21583 (N_21583,N_20879,N_20998);
xor U21584 (N_21584,N_20466,N_20823);
xnor U21585 (N_21585,N_20821,N_20541);
and U21586 (N_21586,N_20492,N_20917);
and U21587 (N_21587,N_20754,N_20706);
or U21588 (N_21588,N_20542,N_20921);
nor U21589 (N_21589,N_20998,N_20970);
or U21590 (N_21590,N_20989,N_20885);
and U21591 (N_21591,N_20555,N_20918);
nor U21592 (N_21592,N_20864,N_20608);
nand U21593 (N_21593,N_20600,N_20544);
xnor U21594 (N_21594,N_20793,N_20756);
nor U21595 (N_21595,N_20576,N_20438);
nand U21596 (N_21596,N_20684,N_20862);
nand U21597 (N_21597,N_20937,N_20524);
or U21598 (N_21598,N_20484,N_20929);
nor U21599 (N_21599,N_20804,N_20783);
and U21600 (N_21600,N_21167,N_21047);
xor U21601 (N_21601,N_21505,N_21147);
or U21602 (N_21602,N_21054,N_21477);
or U21603 (N_21603,N_21071,N_21248);
nor U21604 (N_21604,N_21299,N_21205);
or U21605 (N_21605,N_21144,N_21373);
nand U21606 (N_21606,N_21235,N_21595);
nand U21607 (N_21607,N_21128,N_21319);
nand U21608 (N_21608,N_21192,N_21202);
or U21609 (N_21609,N_21050,N_21525);
nor U21610 (N_21610,N_21499,N_21177);
xnor U21611 (N_21611,N_21511,N_21256);
nor U21612 (N_21612,N_21093,N_21358);
xnor U21613 (N_21613,N_21101,N_21046);
and U21614 (N_21614,N_21360,N_21385);
and U21615 (N_21615,N_21535,N_21020);
xor U21616 (N_21616,N_21179,N_21011);
or U21617 (N_21617,N_21269,N_21145);
xnor U21618 (N_21618,N_21409,N_21129);
nand U21619 (N_21619,N_21201,N_21270);
and U21620 (N_21620,N_21545,N_21188);
nand U21621 (N_21621,N_21591,N_21295);
or U21622 (N_21622,N_21033,N_21582);
xnor U21623 (N_21623,N_21118,N_21051);
xor U21624 (N_21624,N_21002,N_21095);
nor U21625 (N_21625,N_21277,N_21075);
and U21626 (N_21626,N_21066,N_21371);
and U21627 (N_21627,N_21586,N_21484);
nor U21628 (N_21628,N_21379,N_21340);
nand U21629 (N_21629,N_21022,N_21289);
and U21630 (N_21630,N_21544,N_21569);
and U21631 (N_21631,N_21434,N_21162);
nor U21632 (N_21632,N_21483,N_21313);
xnor U21633 (N_21633,N_21194,N_21567);
nor U21634 (N_21634,N_21330,N_21042);
nor U21635 (N_21635,N_21412,N_21305);
xnor U21636 (N_21636,N_21234,N_21007);
nand U21637 (N_21637,N_21443,N_21088);
nand U21638 (N_21638,N_21522,N_21326);
and U21639 (N_21639,N_21456,N_21082);
or U21640 (N_21640,N_21331,N_21476);
nand U21641 (N_21641,N_21490,N_21405);
nand U21642 (N_21642,N_21260,N_21424);
and U21643 (N_21643,N_21265,N_21450);
or U21644 (N_21644,N_21414,N_21131);
or U21645 (N_21645,N_21159,N_21148);
nor U21646 (N_21646,N_21553,N_21052);
or U21647 (N_21647,N_21200,N_21403);
nor U21648 (N_21648,N_21296,N_21485);
or U21649 (N_21649,N_21151,N_21049);
or U21650 (N_21650,N_21551,N_21139);
xor U21651 (N_21651,N_21130,N_21398);
xnor U21652 (N_21652,N_21143,N_21221);
nor U21653 (N_21653,N_21074,N_21195);
nand U21654 (N_21654,N_21264,N_21348);
xor U21655 (N_21655,N_21516,N_21367);
or U21656 (N_21656,N_21261,N_21132);
nand U21657 (N_21657,N_21232,N_21362);
nand U21658 (N_21658,N_21353,N_21172);
and U21659 (N_21659,N_21464,N_21383);
nor U21660 (N_21660,N_21255,N_21573);
or U21661 (N_21661,N_21557,N_21470);
nor U21662 (N_21662,N_21543,N_21336);
xor U21663 (N_21663,N_21279,N_21380);
nand U21664 (N_21664,N_21041,N_21428);
xor U21665 (N_21665,N_21574,N_21210);
or U21666 (N_21666,N_21491,N_21559);
xnor U21667 (N_21667,N_21363,N_21252);
nor U21668 (N_21668,N_21273,N_21396);
and U21669 (N_21669,N_21445,N_21486);
and U21670 (N_21670,N_21572,N_21266);
xor U21671 (N_21671,N_21571,N_21587);
or U21672 (N_21672,N_21400,N_21199);
or U21673 (N_21673,N_21060,N_21004);
nor U21674 (N_21674,N_21006,N_21423);
or U21675 (N_21675,N_21012,N_21211);
and U21676 (N_21676,N_21286,N_21564);
or U21677 (N_21677,N_21016,N_21366);
xor U21678 (N_21678,N_21113,N_21302);
nand U21679 (N_21679,N_21268,N_21480);
xnor U21680 (N_21680,N_21588,N_21080);
or U21681 (N_21681,N_21005,N_21365);
xor U21682 (N_21682,N_21287,N_21184);
nor U21683 (N_21683,N_21078,N_21213);
xor U21684 (N_21684,N_21070,N_21029);
nand U21685 (N_21685,N_21059,N_21244);
nor U21686 (N_21686,N_21243,N_21419);
or U21687 (N_21687,N_21431,N_21369);
and U21688 (N_21688,N_21533,N_21173);
or U21689 (N_21689,N_21351,N_21422);
nor U21690 (N_21690,N_21108,N_21001);
and U21691 (N_21691,N_21164,N_21182);
or U21692 (N_21692,N_21149,N_21315);
xor U21693 (N_21693,N_21537,N_21216);
or U21694 (N_21694,N_21469,N_21432);
nand U21695 (N_21695,N_21121,N_21361);
xnor U21696 (N_21696,N_21250,N_21272);
nor U21697 (N_21697,N_21061,N_21152);
and U21698 (N_21698,N_21514,N_21158);
or U21699 (N_21699,N_21318,N_21554);
xor U21700 (N_21700,N_21301,N_21442);
or U21701 (N_21701,N_21109,N_21104);
xor U21702 (N_21702,N_21136,N_21417);
xor U21703 (N_21703,N_21407,N_21370);
nor U21704 (N_21704,N_21241,N_21566);
or U21705 (N_21705,N_21325,N_21359);
nor U21706 (N_21706,N_21251,N_21242);
or U21707 (N_21707,N_21257,N_21411);
or U21708 (N_21708,N_21284,N_21263);
and U21709 (N_21709,N_21048,N_21576);
nand U21710 (N_21710,N_21427,N_21057);
xor U21711 (N_21711,N_21585,N_21030);
and U21712 (N_21712,N_21141,N_21085);
and U21713 (N_21713,N_21096,N_21013);
nor U21714 (N_21714,N_21119,N_21040);
xnor U21715 (N_21715,N_21283,N_21519);
or U21716 (N_21716,N_21226,N_21032);
xnor U21717 (N_21717,N_21408,N_21364);
or U21718 (N_21718,N_21198,N_21397);
nor U21719 (N_21719,N_21222,N_21328);
and U21720 (N_21720,N_21352,N_21563);
or U21721 (N_21721,N_21441,N_21570);
xor U21722 (N_21722,N_21237,N_21482);
nor U21723 (N_21723,N_21027,N_21290);
nor U21724 (N_21724,N_21240,N_21133);
xor U21725 (N_21725,N_21189,N_21540);
xnor U21726 (N_21726,N_21247,N_21117);
nand U21727 (N_21727,N_21446,N_21138);
nor U21728 (N_21728,N_21274,N_21126);
xnor U21729 (N_21729,N_21308,N_21034);
or U21730 (N_21730,N_21298,N_21097);
xnor U21731 (N_21731,N_21528,N_21455);
xnor U21732 (N_21732,N_21094,N_21510);
and U21733 (N_21733,N_21125,N_21347);
or U21734 (N_21734,N_21062,N_21171);
or U21735 (N_21735,N_21521,N_21539);
nor U21736 (N_21736,N_21390,N_21324);
nor U21737 (N_21737,N_21561,N_21463);
or U21738 (N_21738,N_21281,N_21438);
or U21739 (N_21739,N_21120,N_21067);
and U21740 (N_21740,N_21418,N_21479);
nand U21741 (N_21741,N_21003,N_21212);
or U21742 (N_21742,N_21026,N_21376);
nand U21743 (N_21743,N_21249,N_21481);
and U21744 (N_21744,N_21112,N_21219);
and U21745 (N_21745,N_21339,N_21000);
nand U21746 (N_21746,N_21223,N_21087);
or U21747 (N_21747,N_21449,N_21401);
xor U21748 (N_21748,N_21160,N_21531);
nand U21749 (N_21749,N_21236,N_21494);
and U21750 (N_21750,N_21106,N_21036);
or U21751 (N_21751,N_21154,N_21452);
nor U21752 (N_21752,N_21024,N_21025);
nor U21753 (N_21753,N_21107,N_21337);
nand U21754 (N_21754,N_21447,N_21526);
and U21755 (N_21755,N_21204,N_21415);
or U21756 (N_21756,N_21218,N_21388);
nor U21757 (N_21757,N_21292,N_21191);
nand U21758 (N_21758,N_21342,N_21069);
and U21759 (N_21759,N_21598,N_21303);
xor U21760 (N_21760,N_21150,N_21406);
nand U21761 (N_21761,N_21596,N_21534);
xnor U21762 (N_21762,N_21555,N_21239);
or U21763 (N_21763,N_21161,N_21382);
or U21764 (N_21764,N_21377,N_21375);
and U21765 (N_21765,N_21384,N_21542);
xnor U21766 (N_21766,N_21053,N_21115);
nor U21767 (N_21767,N_21580,N_21043);
xor U21768 (N_21768,N_21142,N_21157);
and U21769 (N_21769,N_21503,N_21170);
or U21770 (N_21770,N_21124,N_21044);
xor U21771 (N_21771,N_21317,N_21497);
nand U21772 (N_21772,N_21552,N_21562);
nor U21773 (N_21773,N_21393,N_21500);
nand U21774 (N_21774,N_21246,N_21245);
nand U21775 (N_21775,N_21114,N_21076);
and U21776 (N_21776,N_21293,N_21338);
xor U21777 (N_21777,N_21448,N_21183);
and U21778 (N_21778,N_21495,N_21310);
and U21779 (N_21779,N_21530,N_21518);
or U21780 (N_21780,N_21517,N_21341);
or U21781 (N_21781,N_21037,N_21506);
or U21782 (N_21782,N_21233,N_21072);
or U21783 (N_21783,N_21304,N_21178);
and U21784 (N_21784,N_21015,N_21238);
nand U21785 (N_21785,N_21321,N_21579);
nand U21786 (N_21786,N_21231,N_21541);
nand U21787 (N_21787,N_21254,N_21073);
or U21788 (N_21788,N_21225,N_21402);
xor U21789 (N_21789,N_21590,N_21462);
or U21790 (N_21790,N_21322,N_21593);
xnor U21791 (N_21791,N_21465,N_21058);
or U21792 (N_21792,N_21467,N_21578);
and U21793 (N_21793,N_21134,N_21089);
nor U21794 (N_21794,N_21155,N_21473);
and U21795 (N_21795,N_21391,N_21181);
or U21796 (N_21796,N_21056,N_21451);
or U21797 (N_21797,N_21459,N_21187);
nand U21798 (N_21798,N_21291,N_21214);
nand U21799 (N_21799,N_21014,N_21258);
or U21800 (N_21800,N_21532,N_21513);
nor U21801 (N_21801,N_21426,N_21594);
xor U21802 (N_21802,N_21496,N_21116);
or U21803 (N_21803,N_21174,N_21294);
nand U21804 (N_21804,N_21548,N_21259);
xor U21805 (N_21805,N_21207,N_21357);
xnor U21806 (N_21806,N_21461,N_21453);
nand U21807 (N_21807,N_21153,N_21487);
xnor U21808 (N_21808,N_21507,N_21413);
nand U21809 (N_21809,N_21086,N_21589);
and U21810 (N_21810,N_21489,N_21560);
nand U21811 (N_21811,N_21436,N_21420);
nand U21812 (N_21812,N_21230,N_21343);
nand U21813 (N_21813,N_21017,N_21297);
xnor U21814 (N_21814,N_21081,N_21504);
nor U21815 (N_21815,N_21556,N_21288);
nand U21816 (N_21816,N_21520,N_21100);
and U21817 (N_21817,N_21549,N_21253);
or U21818 (N_21818,N_21193,N_21156);
or U21819 (N_21819,N_21039,N_21092);
xor U21820 (N_21820,N_21140,N_21471);
or U21821 (N_21821,N_21175,N_21217);
nor U21822 (N_21822,N_21227,N_21098);
xnor U21823 (N_21823,N_21565,N_21444);
and U21824 (N_21824,N_21440,N_21224);
xnor U21825 (N_21825,N_21394,N_21008);
nor U21826 (N_21826,N_21329,N_21038);
xnor U21827 (N_21827,N_21165,N_21278);
nor U21828 (N_21828,N_21169,N_21334);
nand U21829 (N_21829,N_21502,N_21421);
and U21830 (N_21830,N_21135,N_21498);
xnor U21831 (N_21831,N_21435,N_21009);
nand U21832 (N_21832,N_21285,N_21267);
xnor U21833 (N_21833,N_21311,N_21512);
and U21834 (N_21834,N_21316,N_21454);
nor U21835 (N_21835,N_21381,N_21378);
xor U21836 (N_21836,N_21508,N_21524);
nor U21837 (N_21837,N_21546,N_21327);
and U21838 (N_21838,N_21583,N_21399);
nor U21839 (N_21839,N_21433,N_21084);
or U21840 (N_21840,N_21387,N_21314);
or U21841 (N_21841,N_21475,N_21190);
nand U21842 (N_21842,N_21460,N_21090);
nand U21843 (N_21843,N_21068,N_21350);
and U21844 (N_21844,N_21309,N_21478);
nor U21845 (N_21845,N_21439,N_21262);
nand U21846 (N_21846,N_21091,N_21110);
nor U21847 (N_21847,N_21079,N_21035);
and U21848 (N_21848,N_21346,N_21332);
nor U21849 (N_21849,N_21077,N_21206);
or U21850 (N_21850,N_21166,N_21344);
and U21851 (N_21851,N_21523,N_21501);
or U21852 (N_21852,N_21215,N_21122);
and U21853 (N_21853,N_21599,N_21457);
or U21854 (N_21854,N_21186,N_21306);
nand U21855 (N_21855,N_21584,N_21354);
nand U21856 (N_21856,N_21123,N_21064);
or U21857 (N_21857,N_21168,N_21282);
nor U21858 (N_21858,N_21509,N_21276);
and U21859 (N_21859,N_21312,N_21031);
or U21860 (N_21860,N_21105,N_21389);
and U21861 (N_21861,N_21127,N_21597);
or U21862 (N_21862,N_21180,N_21063);
nand U21863 (N_21863,N_21345,N_21271);
nor U21864 (N_21864,N_21458,N_21220);
xnor U21865 (N_21865,N_21300,N_21536);
or U21866 (N_21866,N_21568,N_21395);
nor U21867 (N_21867,N_21515,N_21045);
nor U21868 (N_21868,N_21472,N_21021);
and U21869 (N_21869,N_21437,N_21176);
nor U21870 (N_21870,N_21203,N_21335);
nand U21871 (N_21871,N_21083,N_21197);
nor U21872 (N_21872,N_21275,N_21538);
and U21873 (N_21873,N_21185,N_21229);
xor U21874 (N_21874,N_21349,N_21163);
and U21875 (N_21875,N_21529,N_21374);
xnor U21876 (N_21876,N_21055,N_21333);
or U21877 (N_21877,N_21019,N_21323);
or U21878 (N_21878,N_21493,N_21209);
xor U21879 (N_21879,N_21137,N_21429);
nor U21880 (N_21880,N_21102,N_21492);
nor U21881 (N_21881,N_21018,N_21425);
nor U21882 (N_21882,N_21355,N_21320);
or U21883 (N_21883,N_21575,N_21410);
and U21884 (N_21884,N_21558,N_21550);
nand U21885 (N_21885,N_21592,N_21372);
and U21886 (N_21886,N_21468,N_21547);
nor U21887 (N_21887,N_21099,N_21466);
or U21888 (N_21888,N_21474,N_21146);
or U21889 (N_21889,N_21392,N_21577);
nand U21890 (N_21890,N_21010,N_21307);
or U21891 (N_21891,N_21368,N_21028);
and U21892 (N_21892,N_21208,N_21228);
and U21893 (N_21893,N_21404,N_21416);
nor U21894 (N_21894,N_21581,N_21196);
nand U21895 (N_21895,N_21280,N_21430);
xor U21896 (N_21896,N_21488,N_21023);
xnor U21897 (N_21897,N_21527,N_21386);
and U21898 (N_21898,N_21065,N_21356);
nand U21899 (N_21899,N_21111,N_21103);
xor U21900 (N_21900,N_21158,N_21110);
or U21901 (N_21901,N_21502,N_21486);
and U21902 (N_21902,N_21405,N_21345);
nor U21903 (N_21903,N_21366,N_21090);
and U21904 (N_21904,N_21109,N_21091);
or U21905 (N_21905,N_21369,N_21051);
and U21906 (N_21906,N_21379,N_21004);
nor U21907 (N_21907,N_21276,N_21254);
nor U21908 (N_21908,N_21482,N_21328);
xnor U21909 (N_21909,N_21360,N_21066);
nand U21910 (N_21910,N_21282,N_21289);
or U21911 (N_21911,N_21301,N_21074);
nor U21912 (N_21912,N_21075,N_21081);
and U21913 (N_21913,N_21076,N_21331);
xnor U21914 (N_21914,N_21594,N_21040);
or U21915 (N_21915,N_21128,N_21382);
and U21916 (N_21916,N_21083,N_21006);
nand U21917 (N_21917,N_21032,N_21438);
xnor U21918 (N_21918,N_21408,N_21106);
or U21919 (N_21919,N_21559,N_21359);
nand U21920 (N_21920,N_21108,N_21166);
xor U21921 (N_21921,N_21112,N_21513);
or U21922 (N_21922,N_21047,N_21267);
nor U21923 (N_21923,N_21542,N_21375);
or U21924 (N_21924,N_21187,N_21543);
and U21925 (N_21925,N_21021,N_21490);
or U21926 (N_21926,N_21410,N_21084);
nand U21927 (N_21927,N_21220,N_21596);
and U21928 (N_21928,N_21432,N_21241);
nor U21929 (N_21929,N_21228,N_21220);
nand U21930 (N_21930,N_21412,N_21423);
nor U21931 (N_21931,N_21392,N_21238);
nor U21932 (N_21932,N_21552,N_21247);
or U21933 (N_21933,N_21018,N_21150);
or U21934 (N_21934,N_21358,N_21321);
nor U21935 (N_21935,N_21208,N_21350);
and U21936 (N_21936,N_21429,N_21253);
xnor U21937 (N_21937,N_21573,N_21519);
nor U21938 (N_21938,N_21422,N_21430);
and U21939 (N_21939,N_21413,N_21586);
xnor U21940 (N_21940,N_21448,N_21084);
nor U21941 (N_21941,N_21468,N_21163);
and U21942 (N_21942,N_21082,N_21517);
or U21943 (N_21943,N_21291,N_21031);
xnor U21944 (N_21944,N_21472,N_21499);
or U21945 (N_21945,N_21304,N_21581);
nor U21946 (N_21946,N_21115,N_21463);
nor U21947 (N_21947,N_21306,N_21110);
or U21948 (N_21948,N_21571,N_21275);
or U21949 (N_21949,N_21308,N_21119);
xnor U21950 (N_21950,N_21251,N_21588);
or U21951 (N_21951,N_21092,N_21584);
nand U21952 (N_21952,N_21313,N_21004);
nor U21953 (N_21953,N_21482,N_21230);
and U21954 (N_21954,N_21135,N_21081);
xnor U21955 (N_21955,N_21454,N_21411);
nor U21956 (N_21956,N_21356,N_21327);
and U21957 (N_21957,N_21329,N_21132);
xnor U21958 (N_21958,N_21106,N_21476);
or U21959 (N_21959,N_21132,N_21573);
and U21960 (N_21960,N_21550,N_21392);
xor U21961 (N_21961,N_21368,N_21291);
nand U21962 (N_21962,N_21079,N_21443);
nor U21963 (N_21963,N_21180,N_21471);
nand U21964 (N_21964,N_21598,N_21507);
or U21965 (N_21965,N_21341,N_21593);
and U21966 (N_21966,N_21469,N_21036);
or U21967 (N_21967,N_21593,N_21520);
nand U21968 (N_21968,N_21013,N_21317);
nor U21969 (N_21969,N_21555,N_21285);
nor U21970 (N_21970,N_21185,N_21242);
nand U21971 (N_21971,N_21542,N_21430);
and U21972 (N_21972,N_21590,N_21580);
or U21973 (N_21973,N_21406,N_21541);
and U21974 (N_21974,N_21073,N_21423);
or U21975 (N_21975,N_21142,N_21235);
and U21976 (N_21976,N_21284,N_21007);
nor U21977 (N_21977,N_21577,N_21407);
nor U21978 (N_21978,N_21018,N_21499);
and U21979 (N_21979,N_21161,N_21422);
or U21980 (N_21980,N_21306,N_21118);
or U21981 (N_21981,N_21561,N_21291);
xor U21982 (N_21982,N_21261,N_21471);
nand U21983 (N_21983,N_21302,N_21126);
and U21984 (N_21984,N_21024,N_21522);
nand U21985 (N_21985,N_21358,N_21572);
or U21986 (N_21986,N_21404,N_21344);
nor U21987 (N_21987,N_21310,N_21573);
or U21988 (N_21988,N_21404,N_21069);
nor U21989 (N_21989,N_21121,N_21409);
nand U21990 (N_21990,N_21033,N_21167);
or U21991 (N_21991,N_21200,N_21456);
nor U21992 (N_21992,N_21137,N_21274);
and U21993 (N_21993,N_21166,N_21486);
xor U21994 (N_21994,N_21472,N_21391);
or U21995 (N_21995,N_21401,N_21422);
or U21996 (N_21996,N_21115,N_21214);
xnor U21997 (N_21997,N_21024,N_21177);
xnor U21998 (N_21998,N_21370,N_21333);
nor U21999 (N_21999,N_21414,N_21323);
or U22000 (N_22000,N_21596,N_21544);
or U22001 (N_22001,N_21508,N_21236);
nand U22002 (N_22002,N_21426,N_21206);
xnor U22003 (N_22003,N_21525,N_21189);
or U22004 (N_22004,N_21128,N_21290);
and U22005 (N_22005,N_21215,N_21027);
xnor U22006 (N_22006,N_21434,N_21005);
and U22007 (N_22007,N_21165,N_21214);
nor U22008 (N_22008,N_21114,N_21520);
xnor U22009 (N_22009,N_21123,N_21402);
nand U22010 (N_22010,N_21463,N_21265);
and U22011 (N_22011,N_21437,N_21348);
nand U22012 (N_22012,N_21257,N_21016);
or U22013 (N_22013,N_21284,N_21505);
nand U22014 (N_22014,N_21156,N_21598);
and U22015 (N_22015,N_21355,N_21114);
and U22016 (N_22016,N_21507,N_21266);
nand U22017 (N_22017,N_21561,N_21259);
and U22018 (N_22018,N_21032,N_21503);
nand U22019 (N_22019,N_21150,N_21316);
nor U22020 (N_22020,N_21505,N_21126);
nand U22021 (N_22021,N_21568,N_21534);
and U22022 (N_22022,N_21519,N_21334);
nor U22023 (N_22023,N_21277,N_21086);
nor U22024 (N_22024,N_21549,N_21072);
and U22025 (N_22025,N_21198,N_21046);
nor U22026 (N_22026,N_21056,N_21194);
and U22027 (N_22027,N_21452,N_21528);
or U22028 (N_22028,N_21072,N_21228);
nand U22029 (N_22029,N_21168,N_21093);
nor U22030 (N_22030,N_21518,N_21556);
nor U22031 (N_22031,N_21125,N_21438);
nand U22032 (N_22032,N_21058,N_21098);
nand U22033 (N_22033,N_21506,N_21085);
xnor U22034 (N_22034,N_21566,N_21531);
or U22035 (N_22035,N_21168,N_21035);
xor U22036 (N_22036,N_21036,N_21515);
xor U22037 (N_22037,N_21205,N_21336);
nand U22038 (N_22038,N_21359,N_21360);
or U22039 (N_22039,N_21438,N_21158);
xnor U22040 (N_22040,N_21589,N_21567);
or U22041 (N_22041,N_21114,N_21006);
nor U22042 (N_22042,N_21560,N_21166);
nor U22043 (N_22043,N_21036,N_21099);
nand U22044 (N_22044,N_21440,N_21507);
and U22045 (N_22045,N_21000,N_21244);
nand U22046 (N_22046,N_21022,N_21112);
or U22047 (N_22047,N_21013,N_21534);
and U22048 (N_22048,N_21197,N_21323);
and U22049 (N_22049,N_21381,N_21383);
xor U22050 (N_22050,N_21404,N_21304);
and U22051 (N_22051,N_21390,N_21400);
nor U22052 (N_22052,N_21089,N_21511);
nor U22053 (N_22053,N_21059,N_21476);
or U22054 (N_22054,N_21325,N_21207);
xnor U22055 (N_22055,N_21276,N_21124);
xor U22056 (N_22056,N_21435,N_21343);
nor U22057 (N_22057,N_21598,N_21167);
xnor U22058 (N_22058,N_21207,N_21053);
nor U22059 (N_22059,N_21252,N_21021);
and U22060 (N_22060,N_21392,N_21279);
nor U22061 (N_22061,N_21462,N_21082);
and U22062 (N_22062,N_21426,N_21539);
xor U22063 (N_22063,N_21428,N_21329);
and U22064 (N_22064,N_21414,N_21321);
or U22065 (N_22065,N_21441,N_21443);
nand U22066 (N_22066,N_21215,N_21351);
or U22067 (N_22067,N_21258,N_21368);
xnor U22068 (N_22068,N_21523,N_21261);
xnor U22069 (N_22069,N_21561,N_21311);
or U22070 (N_22070,N_21310,N_21106);
nor U22071 (N_22071,N_21023,N_21092);
or U22072 (N_22072,N_21204,N_21141);
or U22073 (N_22073,N_21426,N_21081);
xor U22074 (N_22074,N_21413,N_21215);
xor U22075 (N_22075,N_21411,N_21040);
xnor U22076 (N_22076,N_21455,N_21008);
nor U22077 (N_22077,N_21545,N_21321);
xnor U22078 (N_22078,N_21320,N_21445);
nor U22079 (N_22079,N_21064,N_21435);
xor U22080 (N_22080,N_21349,N_21105);
nand U22081 (N_22081,N_21599,N_21519);
nand U22082 (N_22082,N_21205,N_21303);
and U22083 (N_22083,N_21119,N_21276);
or U22084 (N_22084,N_21127,N_21595);
nand U22085 (N_22085,N_21170,N_21237);
nor U22086 (N_22086,N_21154,N_21079);
and U22087 (N_22087,N_21230,N_21056);
nor U22088 (N_22088,N_21339,N_21045);
and U22089 (N_22089,N_21313,N_21540);
nor U22090 (N_22090,N_21509,N_21109);
or U22091 (N_22091,N_21174,N_21348);
or U22092 (N_22092,N_21025,N_21486);
or U22093 (N_22093,N_21435,N_21294);
xnor U22094 (N_22094,N_21554,N_21071);
nor U22095 (N_22095,N_21366,N_21396);
and U22096 (N_22096,N_21595,N_21578);
and U22097 (N_22097,N_21004,N_21328);
or U22098 (N_22098,N_21062,N_21480);
and U22099 (N_22099,N_21248,N_21178);
nor U22100 (N_22100,N_21401,N_21536);
nor U22101 (N_22101,N_21567,N_21442);
xor U22102 (N_22102,N_21581,N_21384);
nor U22103 (N_22103,N_21279,N_21073);
and U22104 (N_22104,N_21045,N_21083);
and U22105 (N_22105,N_21286,N_21155);
and U22106 (N_22106,N_21050,N_21008);
nor U22107 (N_22107,N_21524,N_21274);
nand U22108 (N_22108,N_21003,N_21581);
nor U22109 (N_22109,N_21491,N_21172);
or U22110 (N_22110,N_21589,N_21132);
and U22111 (N_22111,N_21162,N_21241);
xor U22112 (N_22112,N_21374,N_21339);
nand U22113 (N_22113,N_21581,N_21292);
nand U22114 (N_22114,N_21375,N_21093);
nand U22115 (N_22115,N_21546,N_21208);
xnor U22116 (N_22116,N_21417,N_21392);
xor U22117 (N_22117,N_21125,N_21571);
nor U22118 (N_22118,N_21081,N_21020);
xor U22119 (N_22119,N_21343,N_21015);
and U22120 (N_22120,N_21566,N_21302);
nor U22121 (N_22121,N_21494,N_21130);
or U22122 (N_22122,N_21453,N_21093);
nor U22123 (N_22123,N_21180,N_21124);
or U22124 (N_22124,N_21571,N_21335);
and U22125 (N_22125,N_21496,N_21130);
nand U22126 (N_22126,N_21178,N_21016);
xor U22127 (N_22127,N_21351,N_21167);
nand U22128 (N_22128,N_21150,N_21482);
nand U22129 (N_22129,N_21116,N_21308);
nor U22130 (N_22130,N_21064,N_21108);
xor U22131 (N_22131,N_21484,N_21543);
nor U22132 (N_22132,N_21101,N_21021);
xor U22133 (N_22133,N_21066,N_21337);
nor U22134 (N_22134,N_21497,N_21433);
and U22135 (N_22135,N_21458,N_21215);
and U22136 (N_22136,N_21346,N_21255);
nor U22137 (N_22137,N_21179,N_21025);
or U22138 (N_22138,N_21102,N_21173);
nor U22139 (N_22139,N_21519,N_21087);
nand U22140 (N_22140,N_21232,N_21199);
nor U22141 (N_22141,N_21388,N_21238);
nor U22142 (N_22142,N_21362,N_21435);
xor U22143 (N_22143,N_21294,N_21409);
or U22144 (N_22144,N_21014,N_21130);
and U22145 (N_22145,N_21305,N_21386);
xnor U22146 (N_22146,N_21465,N_21522);
and U22147 (N_22147,N_21289,N_21462);
or U22148 (N_22148,N_21466,N_21440);
and U22149 (N_22149,N_21091,N_21595);
or U22150 (N_22150,N_21325,N_21347);
or U22151 (N_22151,N_21070,N_21053);
nor U22152 (N_22152,N_21469,N_21445);
nand U22153 (N_22153,N_21499,N_21236);
nor U22154 (N_22154,N_21529,N_21206);
xor U22155 (N_22155,N_21275,N_21572);
nand U22156 (N_22156,N_21473,N_21239);
nand U22157 (N_22157,N_21481,N_21236);
or U22158 (N_22158,N_21510,N_21099);
xor U22159 (N_22159,N_21252,N_21518);
nand U22160 (N_22160,N_21133,N_21326);
nor U22161 (N_22161,N_21018,N_21214);
or U22162 (N_22162,N_21588,N_21332);
nor U22163 (N_22163,N_21578,N_21316);
and U22164 (N_22164,N_21076,N_21214);
xnor U22165 (N_22165,N_21057,N_21256);
nor U22166 (N_22166,N_21079,N_21102);
nand U22167 (N_22167,N_21235,N_21426);
and U22168 (N_22168,N_21127,N_21467);
and U22169 (N_22169,N_21172,N_21030);
nand U22170 (N_22170,N_21031,N_21160);
nor U22171 (N_22171,N_21429,N_21117);
and U22172 (N_22172,N_21365,N_21271);
and U22173 (N_22173,N_21282,N_21055);
nand U22174 (N_22174,N_21517,N_21216);
and U22175 (N_22175,N_21046,N_21570);
nor U22176 (N_22176,N_21535,N_21368);
nand U22177 (N_22177,N_21412,N_21435);
or U22178 (N_22178,N_21554,N_21485);
nor U22179 (N_22179,N_21257,N_21485);
xor U22180 (N_22180,N_21225,N_21163);
xor U22181 (N_22181,N_21573,N_21473);
nand U22182 (N_22182,N_21055,N_21173);
or U22183 (N_22183,N_21172,N_21442);
nand U22184 (N_22184,N_21152,N_21147);
xor U22185 (N_22185,N_21586,N_21293);
and U22186 (N_22186,N_21288,N_21084);
xor U22187 (N_22187,N_21002,N_21548);
nand U22188 (N_22188,N_21522,N_21300);
and U22189 (N_22189,N_21224,N_21185);
xor U22190 (N_22190,N_21083,N_21005);
and U22191 (N_22191,N_21233,N_21143);
nor U22192 (N_22192,N_21284,N_21559);
and U22193 (N_22193,N_21338,N_21157);
xor U22194 (N_22194,N_21532,N_21144);
and U22195 (N_22195,N_21060,N_21300);
nand U22196 (N_22196,N_21169,N_21421);
nor U22197 (N_22197,N_21078,N_21180);
xor U22198 (N_22198,N_21335,N_21373);
xnor U22199 (N_22199,N_21581,N_21096);
or U22200 (N_22200,N_22173,N_22111);
xnor U22201 (N_22201,N_21980,N_21858);
xnor U22202 (N_22202,N_21816,N_21946);
xnor U22203 (N_22203,N_21734,N_22056);
nor U22204 (N_22204,N_21633,N_21803);
and U22205 (N_22205,N_21975,N_21753);
nor U22206 (N_22206,N_22027,N_22162);
nand U22207 (N_22207,N_22151,N_21733);
xor U22208 (N_22208,N_22185,N_22070);
or U22209 (N_22209,N_21658,N_21773);
nor U22210 (N_22210,N_21872,N_21792);
nor U22211 (N_22211,N_22004,N_21786);
and U22212 (N_22212,N_21842,N_22082);
nor U22213 (N_22213,N_21862,N_21993);
xor U22214 (N_22214,N_21759,N_21983);
or U22215 (N_22215,N_21672,N_21802);
or U22216 (N_22216,N_22050,N_22023);
or U22217 (N_22217,N_21697,N_21906);
nor U22218 (N_22218,N_22181,N_21984);
or U22219 (N_22219,N_21891,N_22064);
nor U22220 (N_22220,N_21806,N_21965);
nor U22221 (N_22221,N_22096,N_21882);
xnor U22222 (N_22222,N_21784,N_21772);
nor U22223 (N_22223,N_21605,N_22199);
or U22224 (N_22224,N_21704,N_22104);
nor U22225 (N_22225,N_21995,N_21673);
nand U22226 (N_22226,N_21699,N_22179);
and U22227 (N_22227,N_21927,N_21774);
and U22228 (N_22228,N_22143,N_21838);
xor U22229 (N_22229,N_21837,N_21741);
nand U22230 (N_22230,N_21840,N_22063);
xor U22231 (N_22231,N_21903,N_21620);
nor U22232 (N_22232,N_21726,N_21933);
nand U22233 (N_22233,N_21963,N_21950);
or U22234 (N_22234,N_21740,N_21607);
nand U22235 (N_22235,N_21700,N_21931);
nor U22236 (N_22236,N_22045,N_21650);
xnor U22237 (N_22237,N_21789,N_21920);
or U22238 (N_22238,N_21897,N_21643);
xor U22239 (N_22239,N_21818,N_22041);
nor U22240 (N_22240,N_21628,N_21994);
and U22241 (N_22241,N_22134,N_21738);
nor U22242 (N_22242,N_22095,N_21793);
nand U22243 (N_22243,N_21695,N_22080);
and U22244 (N_22244,N_21747,N_21796);
or U22245 (N_22245,N_21798,N_22046);
xnor U22246 (N_22246,N_21725,N_21641);
xnor U22247 (N_22247,N_22019,N_22093);
nor U22248 (N_22248,N_22036,N_21601);
xor U22249 (N_22249,N_21832,N_21604);
or U22250 (N_22250,N_22117,N_21805);
nor U22251 (N_22251,N_22069,N_21890);
nand U22252 (N_22252,N_22032,N_22140);
or U22253 (N_22253,N_22057,N_21855);
or U22254 (N_22254,N_21622,N_21947);
or U22255 (N_22255,N_21696,N_21752);
or U22256 (N_22256,N_21720,N_21916);
and U22257 (N_22257,N_21790,N_22109);
nor U22258 (N_22258,N_22024,N_21757);
xnor U22259 (N_22259,N_22010,N_21710);
and U22260 (N_22260,N_21936,N_21848);
nor U22261 (N_22261,N_22110,N_21886);
xor U22262 (N_22262,N_22137,N_21690);
nand U22263 (N_22263,N_21618,N_21626);
nor U22264 (N_22264,N_21959,N_21724);
nand U22265 (N_22265,N_21657,N_22141);
xor U22266 (N_22266,N_21887,N_22139);
nor U22267 (N_22267,N_21787,N_21996);
and U22268 (N_22268,N_21717,N_22171);
xnor U22269 (N_22269,N_22077,N_21804);
nor U22270 (N_22270,N_21870,N_21934);
nand U22271 (N_22271,N_21736,N_22175);
or U22272 (N_22272,N_21871,N_22194);
and U22273 (N_22273,N_21971,N_21619);
or U22274 (N_22274,N_21844,N_22145);
xor U22275 (N_22275,N_21865,N_22060);
nand U22276 (N_22276,N_21925,N_21714);
nand U22277 (N_22277,N_21692,N_22102);
or U22278 (N_22278,N_21705,N_22103);
and U22279 (N_22279,N_21991,N_21610);
or U22280 (N_22280,N_21797,N_21681);
and U22281 (N_22281,N_21986,N_21914);
nor U22282 (N_22282,N_21666,N_22062);
nand U22283 (N_22283,N_22028,N_21908);
xnor U22284 (N_22284,N_21809,N_21867);
and U22285 (N_22285,N_22066,N_21721);
or U22286 (N_22286,N_21990,N_21910);
xor U22287 (N_22287,N_21782,N_21881);
nor U22288 (N_22288,N_21964,N_21821);
and U22289 (N_22289,N_21754,N_21636);
nand U22290 (N_22290,N_22116,N_22067);
nor U22291 (N_22291,N_21667,N_21864);
xor U22292 (N_22292,N_22124,N_22106);
nor U22293 (N_22293,N_21877,N_22051);
or U22294 (N_22294,N_22005,N_21621);
nand U22295 (N_22295,N_21829,N_22108);
nor U22296 (N_22296,N_22125,N_21999);
xnor U22297 (N_22297,N_21716,N_22091);
nand U22298 (N_22298,N_21711,N_21679);
and U22299 (N_22299,N_21830,N_21654);
and U22300 (N_22300,N_21823,N_21889);
or U22301 (N_22301,N_21630,N_22118);
or U22302 (N_22302,N_21969,N_21879);
nor U22303 (N_22303,N_21686,N_21954);
nand U22304 (N_22304,N_22012,N_22039);
xor U22305 (N_22305,N_21857,N_21613);
or U22306 (N_22306,N_22163,N_22044);
or U22307 (N_22307,N_21730,N_21776);
xor U22308 (N_22308,N_22138,N_21694);
nand U22309 (N_22309,N_22015,N_22161);
nor U22310 (N_22310,N_21744,N_21913);
nor U22311 (N_22311,N_22088,N_21850);
or U22312 (N_22312,N_21751,N_22089);
or U22313 (N_22313,N_22136,N_22198);
nor U22314 (N_22314,N_22182,N_22186);
or U22315 (N_22315,N_21836,N_21684);
nand U22316 (N_22316,N_21712,N_21888);
and U22317 (N_22317,N_22094,N_22043);
nand U22318 (N_22318,N_22018,N_21884);
nor U22319 (N_22319,N_22029,N_21631);
or U22320 (N_22320,N_21616,N_22196);
and U22321 (N_22321,N_21670,N_21860);
xor U22322 (N_22322,N_21928,N_21939);
and U22323 (N_22323,N_22142,N_21849);
and U22324 (N_22324,N_22065,N_21750);
nand U22325 (N_22325,N_21737,N_21861);
nand U22326 (N_22326,N_22052,N_21761);
or U22327 (N_22327,N_21831,N_21943);
nand U22328 (N_22328,N_21693,N_22086);
and U22329 (N_22329,N_21788,N_22147);
nand U22330 (N_22330,N_21834,N_21680);
or U22331 (N_22331,N_22033,N_21957);
nand U22332 (N_22332,N_21899,N_21968);
nand U22333 (N_22333,N_22030,N_22164);
or U22334 (N_22334,N_21634,N_22007);
or U22335 (N_22335,N_21687,N_22105);
xnor U22336 (N_22336,N_21824,N_22100);
and U22337 (N_22337,N_22191,N_21929);
nor U22338 (N_22338,N_21677,N_21958);
or U22339 (N_22339,N_21742,N_21791);
or U22340 (N_22340,N_21602,N_21952);
and U22341 (N_22341,N_21880,N_22107);
or U22342 (N_22342,N_22017,N_21825);
and U22343 (N_22343,N_22058,N_21612);
nor U22344 (N_22344,N_21876,N_21770);
or U22345 (N_22345,N_21907,N_21745);
xnor U22346 (N_22346,N_21852,N_21767);
nor U22347 (N_22347,N_22155,N_22148);
nand U22348 (N_22348,N_22183,N_22002);
nand U22349 (N_22349,N_21854,N_22011);
nor U22350 (N_22350,N_21718,N_22079);
or U22351 (N_22351,N_21807,N_22092);
xor U22352 (N_22352,N_21894,N_22189);
nor U22353 (N_22353,N_21649,N_22072);
and U22354 (N_22354,N_21841,N_21760);
or U22355 (N_22355,N_22031,N_21924);
nand U22356 (N_22356,N_21977,N_21935);
and U22357 (N_22357,N_22022,N_21902);
nor U22358 (N_22358,N_21780,N_22193);
nand U22359 (N_22359,N_22123,N_21951);
and U22360 (N_22360,N_21685,N_21659);
or U22361 (N_22361,N_21937,N_21708);
xnor U22362 (N_22362,N_21938,N_22037);
nor U22363 (N_22363,N_22025,N_22034);
and U22364 (N_22364,N_21988,N_21702);
nand U22365 (N_22365,N_21691,N_21748);
nor U22366 (N_22366,N_21715,N_22153);
nor U22367 (N_22367,N_22048,N_21828);
and U22368 (N_22368,N_21810,N_21648);
and U22369 (N_22369,N_21663,N_21981);
or U22370 (N_22370,N_21635,N_21956);
and U22371 (N_22371,N_22087,N_21811);
and U22372 (N_22372,N_22190,N_21678);
or U22373 (N_22373,N_22167,N_21723);
and U22374 (N_22374,N_21851,N_22075);
and U22375 (N_22375,N_21632,N_22135);
nand U22376 (N_22376,N_22192,N_22038);
nor U22377 (N_22377,N_21982,N_22131);
nor U22378 (N_22378,N_22068,N_21698);
or U22379 (N_22379,N_21972,N_22009);
nand U22380 (N_22380,N_21728,N_21664);
or U22381 (N_22381,N_21683,N_22008);
and U22382 (N_22382,N_22099,N_21966);
nand U22383 (N_22383,N_21978,N_22047);
and U22384 (N_22384,N_21921,N_21671);
nor U22385 (N_22385,N_21662,N_22166);
and U22386 (N_22386,N_21703,N_21668);
xnor U22387 (N_22387,N_21960,N_22059);
xnor U22388 (N_22388,N_21945,N_22078);
and U22389 (N_22389,N_21606,N_21615);
nor U22390 (N_22390,N_22083,N_21701);
nor U22391 (N_22391,N_21617,N_22021);
xor U22392 (N_22392,N_21746,N_21755);
or U22393 (N_22393,N_22128,N_22150);
nand U22394 (N_22394,N_21846,N_21608);
nand U22395 (N_22395,N_21813,N_21713);
xor U22396 (N_22396,N_21727,N_21898);
and U22397 (N_22397,N_21765,N_21729);
nand U22398 (N_22398,N_21799,N_21785);
nor U22399 (N_22399,N_22156,N_22154);
nor U22400 (N_22400,N_22177,N_21896);
xor U22401 (N_22401,N_21669,N_22000);
nor U22402 (N_22402,N_21859,N_21992);
xnor U22403 (N_22403,N_21874,N_22149);
nand U22404 (N_22404,N_21800,N_21778);
nor U22405 (N_22405,N_22114,N_21652);
nor U22406 (N_22406,N_21904,N_21900);
nand U22407 (N_22407,N_22126,N_22188);
nand U22408 (N_22408,N_22054,N_22049);
xnor U22409 (N_22409,N_21783,N_22014);
nand U22410 (N_22410,N_21614,N_22129);
xor U22411 (N_22411,N_21843,N_21771);
xnor U22412 (N_22412,N_21624,N_21893);
or U22413 (N_22413,N_21707,N_21922);
or U22414 (N_22414,N_22195,N_21651);
and U22415 (N_22415,N_21820,N_22146);
nand U22416 (N_22416,N_22152,N_22003);
nor U22417 (N_22417,N_21719,N_21709);
nand U22418 (N_22418,N_21839,N_21973);
nor U22419 (N_22419,N_22112,N_22026);
xor U22420 (N_22420,N_21682,N_21918);
or U22421 (N_22421,N_22130,N_21629);
nor U22422 (N_22422,N_22170,N_21762);
and U22423 (N_22423,N_22165,N_22178);
and U22424 (N_22424,N_21827,N_22157);
xnor U22425 (N_22425,N_22174,N_21892);
nand U22426 (N_22426,N_22073,N_22035);
and U22427 (N_22427,N_21637,N_22119);
xnor U22428 (N_22428,N_22081,N_21656);
xor U22429 (N_22429,N_21625,N_22121);
nor U22430 (N_22430,N_21756,N_22144);
nor U22431 (N_22431,N_21835,N_21781);
nor U22432 (N_22432,N_21941,N_21847);
xnor U22433 (N_22433,N_21795,N_22169);
xnor U22434 (N_22434,N_22120,N_21801);
or U22435 (N_22435,N_21905,N_22172);
or U22436 (N_22436,N_21812,N_22001);
xor U22437 (N_22437,N_21642,N_21688);
nor U22438 (N_22438,N_21763,N_22076);
xnor U22439 (N_22439,N_22016,N_21653);
nor U22440 (N_22440,N_21808,N_21955);
or U22441 (N_22441,N_21998,N_21749);
xnor U22442 (N_22442,N_21940,N_21675);
nor U22443 (N_22443,N_21609,N_22040);
nor U22444 (N_22444,N_22115,N_21627);
and U22445 (N_22445,N_22122,N_22042);
or U22446 (N_22446,N_21962,N_22176);
or U22447 (N_22447,N_22053,N_22006);
nor U22448 (N_22448,N_21961,N_21895);
nor U22449 (N_22449,N_21731,N_21623);
nand U22450 (N_22450,N_21647,N_21911);
nor U22451 (N_22451,N_21953,N_21970);
nor U22452 (N_22452,N_22074,N_21901);
or U22453 (N_22453,N_22127,N_21976);
nand U22454 (N_22454,N_21853,N_21644);
xor U22455 (N_22455,N_22020,N_21868);
or U22456 (N_22456,N_22113,N_21640);
or U22457 (N_22457,N_22133,N_21646);
xnor U22458 (N_22458,N_21775,N_21815);
xor U22459 (N_22459,N_21676,N_22085);
nor U22460 (N_22460,N_21639,N_21794);
nand U22461 (N_22461,N_22098,N_21777);
nand U22462 (N_22462,N_22197,N_21766);
or U22463 (N_22463,N_21979,N_21764);
and U22464 (N_22464,N_21826,N_22061);
xor U22465 (N_22465,N_21743,N_21768);
nand U22466 (N_22466,N_21735,N_21689);
or U22467 (N_22467,N_21674,N_22084);
and U22468 (N_22468,N_21817,N_22180);
or U22469 (N_22469,N_22184,N_21967);
or U22470 (N_22470,N_21987,N_21989);
nand U22471 (N_22471,N_21638,N_21665);
or U22472 (N_22472,N_21779,N_21878);
xor U22473 (N_22473,N_21923,N_21739);
nand U22474 (N_22474,N_21603,N_21926);
and U22475 (N_22475,N_22101,N_21814);
nand U22476 (N_22476,N_21944,N_22187);
nand U22477 (N_22477,N_21997,N_21706);
or U22478 (N_22478,N_22013,N_22090);
and U22479 (N_22479,N_21869,N_21915);
and U22480 (N_22480,N_21949,N_21985);
nand U22481 (N_22481,N_21660,N_21883);
or U22482 (N_22482,N_22168,N_22055);
or U22483 (N_22483,N_21661,N_22159);
and U22484 (N_22484,N_21600,N_21833);
or U22485 (N_22485,N_21769,N_21645);
or U22486 (N_22486,N_21732,N_21866);
and U22487 (N_22487,N_21611,N_21919);
nand U22488 (N_22488,N_21942,N_21655);
or U22489 (N_22489,N_21819,N_21885);
nor U22490 (N_22490,N_21822,N_21758);
nand U22491 (N_22491,N_22097,N_21932);
xnor U22492 (N_22492,N_21722,N_21930);
or U22493 (N_22493,N_21863,N_21856);
nor U22494 (N_22494,N_22158,N_21845);
xnor U22495 (N_22495,N_21948,N_22071);
xnor U22496 (N_22496,N_21912,N_21917);
and U22497 (N_22497,N_21873,N_21875);
and U22498 (N_22498,N_21909,N_21974);
and U22499 (N_22499,N_22160,N_22132);
xnor U22500 (N_22500,N_21687,N_21738);
or U22501 (N_22501,N_22085,N_21911);
xor U22502 (N_22502,N_21882,N_22130);
nand U22503 (N_22503,N_21891,N_21655);
and U22504 (N_22504,N_22029,N_21923);
xor U22505 (N_22505,N_21719,N_21663);
and U22506 (N_22506,N_21767,N_21978);
or U22507 (N_22507,N_21963,N_21616);
nand U22508 (N_22508,N_21871,N_21678);
and U22509 (N_22509,N_21669,N_21899);
nor U22510 (N_22510,N_21717,N_21872);
and U22511 (N_22511,N_22084,N_22094);
and U22512 (N_22512,N_21615,N_21858);
and U22513 (N_22513,N_21812,N_22007);
nand U22514 (N_22514,N_21782,N_22041);
nor U22515 (N_22515,N_22139,N_21722);
or U22516 (N_22516,N_21735,N_22141);
nand U22517 (N_22517,N_22039,N_21878);
xnor U22518 (N_22518,N_22096,N_21657);
or U22519 (N_22519,N_21743,N_21956);
xor U22520 (N_22520,N_21810,N_22173);
and U22521 (N_22521,N_22096,N_21917);
nand U22522 (N_22522,N_22078,N_22042);
nand U22523 (N_22523,N_21704,N_21649);
and U22524 (N_22524,N_22155,N_21777);
or U22525 (N_22525,N_21907,N_22020);
nand U22526 (N_22526,N_21783,N_21611);
or U22527 (N_22527,N_21720,N_22099);
nor U22528 (N_22528,N_22185,N_21718);
nand U22529 (N_22529,N_21967,N_22118);
xnor U22530 (N_22530,N_21859,N_21827);
xor U22531 (N_22531,N_21601,N_21628);
nand U22532 (N_22532,N_21709,N_21624);
nand U22533 (N_22533,N_21951,N_21928);
or U22534 (N_22534,N_21978,N_21981);
nand U22535 (N_22535,N_21980,N_22045);
or U22536 (N_22536,N_22189,N_21768);
and U22537 (N_22537,N_22071,N_21742);
or U22538 (N_22538,N_22020,N_22178);
and U22539 (N_22539,N_21621,N_21677);
nor U22540 (N_22540,N_21749,N_21919);
and U22541 (N_22541,N_22194,N_21935);
nor U22542 (N_22542,N_21753,N_22022);
nor U22543 (N_22543,N_21804,N_21859);
nor U22544 (N_22544,N_21820,N_21995);
nor U22545 (N_22545,N_21907,N_22059);
nand U22546 (N_22546,N_21963,N_21758);
nor U22547 (N_22547,N_21907,N_21997);
xor U22548 (N_22548,N_21621,N_21717);
and U22549 (N_22549,N_21681,N_21868);
or U22550 (N_22550,N_21969,N_22015);
and U22551 (N_22551,N_21626,N_21982);
and U22552 (N_22552,N_21730,N_21857);
and U22553 (N_22553,N_22156,N_21673);
nand U22554 (N_22554,N_22191,N_22037);
or U22555 (N_22555,N_22026,N_22042);
or U22556 (N_22556,N_21658,N_22070);
nand U22557 (N_22557,N_22122,N_22028);
nand U22558 (N_22558,N_21685,N_21798);
or U22559 (N_22559,N_22140,N_22182);
and U22560 (N_22560,N_21618,N_21921);
and U22561 (N_22561,N_22173,N_21862);
nor U22562 (N_22562,N_22029,N_21951);
nor U22563 (N_22563,N_21789,N_21999);
nor U22564 (N_22564,N_21681,N_21731);
xor U22565 (N_22565,N_21891,N_21805);
nand U22566 (N_22566,N_21661,N_22081);
xor U22567 (N_22567,N_21617,N_22012);
nand U22568 (N_22568,N_22063,N_21973);
nor U22569 (N_22569,N_21871,N_21791);
nor U22570 (N_22570,N_21757,N_22032);
and U22571 (N_22571,N_22006,N_21780);
or U22572 (N_22572,N_21686,N_22148);
nand U22573 (N_22573,N_22039,N_21805);
or U22574 (N_22574,N_21672,N_22109);
and U22575 (N_22575,N_21657,N_21724);
and U22576 (N_22576,N_21865,N_21805);
xnor U22577 (N_22577,N_22159,N_21627);
nor U22578 (N_22578,N_22059,N_21983);
nor U22579 (N_22579,N_21732,N_21657);
nor U22580 (N_22580,N_21775,N_21759);
nor U22581 (N_22581,N_21886,N_21837);
nor U22582 (N_22582,N_21955,N_21753);
nor U22583 (N_22583,N_22179,N_21964);
nand U22584 (N_22584,N_22020,N_21724);
nor U22585 (N_22585,N_21916,N_21923);
and U22586 (N_22586,N_22123,N_21603);
or U22587 (N_22587,N_22188,N_21955);
xnor U22588 (N_22588,N_22069,N_22145);
and U22589 (N_22589,N_22097,N_21758);
nor U22590 (N_22590,N_21712,N_21613);
or U22591 (N_22591,N_21737,N_22192);
nor U22592 (N_22592,N_21926,N_22041);
nor U22593 (N_22593,N_21822,N_21870);
and U22594 (N_22594,N_21663,N_21772);
nand U22595 (N_22595,N_21656,N_21882);
or U22596 (N_22596,N_22155,N_21762);
or U22597 (N_22597,N_21860,N_21817);
nand U22598 (N_22598,N_21896,N_21627);
or U22599 (N_22599,N_21940,N_21963);
xnor U22600 (N_22600,N_22173,N_22123);
xnor U22601 (N_22601,N_22087,N_21867);
nor U22602 (N_22602,N_21742,N_22157);
or U22603 (N_22603,N_21849,N_21696);
nor U22604 (N_22604,N_21707,N_22101);
xor U22605 (N_22605,N_21651,N_22055);
nor U22606 (N_22606,N_21884,N_22185);
xor U22607 (N_22607,N_21939,N_22015);
nand U22608 (N_22608,N_21971,N_21924);
nor U22609 (N_22609,N_22100,N_21960);
nor U22610 (N_22610,N_21835,N_22052);
or U22611 (N_22611,N_22046,N_21946);
or U22612 (N_22612,N_21973,N_22091);
xor U22613 (N_22613,N_22145,N_21772);
and U22614 (N_22614,N_21901,N_22062);
and U22615 (N_22615,N_21856,N_21922);
nor U22616 (N_22616,N_21995,N_21649);
xor U22617 (N_22617,N_21806,N_21769);
and U22618 (N_22618,N_21776,N_21631);
nor U22619 (N_22619,N_21972,N_21793);
xnor U22620 (N_22620,N_21948,N_21797);
nor U22621 (N_22621,N_21674,N_21881);
nor U22622 (N_22622,N_21809,N_21701);
or U22623 (N_22623,N_22154,N_21641);
nand U22624 (N_22624,N_22198,N_21714);
xor U22625 (N_22625,N_21653,N_22170);
or U22626 (N_22626,N_21686,N_22024);
nor U22627 (N_22627,N_21797,N_21782);
or U22628 (N_22628,N_22162,N_21747);
and U22629 (N_22629,N_22048,N_21948);
and U22630 (N_22630,N_21969,N_21666);
xor U22631 (N_22631,N_21868,N_22056);
nand U22632 (N_22632,N_22106,N_21692);
and U22633 (N_22633,N_21634,N_21734);
xnor U22634 (N_22634,N_22094,N_22110);
xor U22635 (N_22635,N_22061,N_22026);
xnor U22636 (N_22636,N_22065,N_21989);
and U22637 (N_22637,N_21794,N_21846);
nor U22638 (N_22638,N_22053,N_21844);
and U22639 (N_22639,N_21833,N_22009);
nor U22640 (N_22640,N_21626,N_21711);
or U22641 (N_22641,N_21750,N_21797);
or U22642 (N_22642,N_22037,N_22125);
nor U22643 (N_22643,N_22077,N_21703);
and U22644 (N_22644,N_21834,N_21715);
and U22645 (N_22645,N_22115,N_21899);
or U22646 (N_22646,N_21729,N_22128);
xnor U22647 (N_22647,N_21943,N_22092);
or U22648 (N_22648,N_21730,N_22137);
nand U22649 (N_22649,N_22095,N_21895);
xnor U22650 (N_22650,N_22140,N_21839);
xnor U22651 (N_22651,N_22053,N_21753);
or U22652 (N_22652,N_21643,N_22038);
nand U22653 (N_22653,N_21610,N_21998);
or U22654 (N_22654,N_21798,N_22142);
xor U22655 (N_22655,N_22118,N_22186);
and U22656 (N_22656,N_22089,N_21916);
xnor U22657 (N_22657,N_21893,N_21835);
xor U22658 (N_22658,N_21709,N_21906);
nand U22659 (N_22659,N_22131,N_22030);
and U22660 (N_22660,N_22048,N_22049);
nand U22661 (N_22661,N_22043,N_22004);
nand U22662 (N_22662,N_22146,N_21917);
nor U22663 (N_22663,N_21701,N_21859);
xnor U22664 (N_22664,N_22076,N_21818);
nor U22665 (N_22665,N_21717,N_21701);
and U22666 (N_22666,N_21690,N_21778);
or U22667 (N_22667,N_21969,N_22193);
nor U22668 (N_22668,N_21719,N_21881);
or U22669 (N_22669,N_21704,N_21939);
xor U22670 (N_22670,N_21756,N_22060);
or U22671 (N_22671,N_21604,N_21633);
or U22672 (N_22672,N_22088,N_21663);
and U22673 (N_22673,N_21716,N_21680);
xor U22674 (N_22674,N_21751,N_21955);
nand U22675 (N_22675,N_21975,N_21934);
xnor U22676 (N_22676,N_21858,N_22099);
xnor U22677 (N_22677,N_22148,N_21720);
or U22678 (N_22678,N_21967,N_22033);
or U22679 (N_22679,N_21610,N_21840);
nor U22680 (N_22680,N_22150,N_21698);
or U22681 (N_22681,N_21763,N_21938);
nand U22682 (N_22682,N_21976,N_21620);
nand U22683 (N_22683,N_21942,N_22099);
nand U22684 (N_22684,N_22064,N_21885);
and U22685 (N_22685,N_21905,N_21609);
xor U22686 (N_22686,N_22075,N_21686);
or U22687 (N_22687,N_22030,N_22011);
and U22688 (N_22688,N_21917,N_22121);
nand U22689 (N_22689,N_21987,N_21846);
or U22690 (N_22690,N_21917,N_21601);
xnor U22691 (N_22691,N_22023,N_21685);
nand U22692 (N_22692,N_21738,N_21996);
xnor U22693 (N_22693,N_22079,N_22077);
nor U22694 (N_22694,N_21893,N_22052);
and U22695 (N_22695,N_21693,N_22103);
nand U22696 (N_22696,N_21833,N_22004);
or U22697 (N_22697,N_21904,N_21789);
nand U22698 (N_22698,N_21973,N_22066);
and U22699 (N_22699,N_21728,N_21973);
and U22700 (N_22700,N_21600,N_21617);
or U22701 (N_22701,N_21790,N_21629);
nor U22702 (N_22702,N_22055,N_21754);
nand U22703 (N_22703,N_21710,N_22073);
nor U22704 (N_22704,N_22165,N_22065);
nor U22705 (N_22705,N_21967,N_21914);
nand U22706 (N_22706,N_21672,N_21715);
nand U22707 (N_22707,N_21803,N_21654);
nand U22708 (N_22708,N_21958,N_22191);
and U22709 (N_22709,N_21985,N_22026);
xnor U22710 (N_22710,N_22001,N_21929);
or U22711 (N_22711,N_21961,N_21606);
and U22712 (N_22712,N_21751,N_21849);
nor U22713 (N_22713,N_22126,N_21688);
or U22714 (N_22714,N_21730,N_22085);
xor U22715 (N_22715,N_21978,N_21620);
xnor U22716 (N_22716,N_22003,N_22186);
or U22717 (N_22717,N_21728,N_21692);
and U22718 (N_22718,N_21968,N_21817);
or U22719 (N_22719,N_22033,N_21737);
nor U22720 (N_22720,N_22142,N_22154);
nand U22721 (N_22721,N_21983,N_21806);
and U22722 (N_22722,N_22071,N_22068);
nor U22723 (N_22723,N_22155,N_22111);
and U22724 (N_22724,N_21931,N_22007);
nand U22725 (N_22725,N_21897,N_21707);
or U22726 (N_22726,N_21725,N_21845);
nor U22727 (N_22727,N_21915,N_22034);
nand U22728 (N_22728,N_21806,N_21978);
xor U22729 (N_22729,N_21642,N_22156);
and U22730 (N_22730,N_21844,N_21995);
or U22731 (N_22731,N_22118,N_21739);
nand U22732 (N_22732,N_22178,N_22026);
xor U22733 (N_22733,N_21986,N_22083);
xnor U22734 (N_22734,N_21947,N_22140);
xnor U22735 (N_22735,N_22111,N_22110);
or U22736 (N_22736,N_21866,N_21843);
or U22737 (N_22737,N_22170,N_21634);
nand U22738 (N_22738,N_21829,N_22088);
or U22739 (N_22739,N_21647,N_22129);
and U22740 (N_22740,N_21743,N_21747);
nand U22741 (N_22741,N_22074,N_21705);
xnor U22742 (N_22742,N_21782,N_21743);
and U22743 (N_22743,N_21929,N_21922);
nor U22744 (N_22744,N_22122,N_21649);
nor U22745 (N_22745,N_21871,N_21929);
nor U22746 (N_22746,N_21614,N_22054);
nand U22747 (N_22747,N_22076,N_22139);
and U22748 (N_22748,N_22155,N_21952);
and U22749 (N_22749,N_22195,N_21951);
and U22750 (N_22750,N_21642,N_21783);
nor U22751 (N_22751,N_21765,N_21758);
nor U22752 (N_22752,N_21724,N_21839);
nand U22753 (N_22753,N_21939,N_22198);
nand U22754 (N_22754,N_21667,N_21694);
nand U22755 (N_22755,N_22154,N_21896);
xor U22756 (N_22756,N_21835,N_21916);
or U22757 (N_22757,N_21717,N_21996);
and U22758 (N_22758,N_21641,N_21639);
nand U22759 (N_22759,N_21749,N_22141);
and U22760 (N_22760,N_21773,N_21825);
or U22761 (N_22761,N_21888,N_21688);
nand U22762 (N_22762,N_21843,N_21877);
nand U22763 (N_22763,N_21919,N_21657);
nand U22764 (N_22764,N_22111,N_21636);
and U22765 (N_22765,N_21652,N_22108);
nor U22766 (N_22766,N_21863,N_21785);
nand U22767 (N_22767,N_21608,N_21748);
nand U22768 (N_22768,N_22172,N_22189);
nor U22769 (N_22769,N_22191,N_22082);
or U22770 (N_22770,N_21773,N_21850);
and U22771 (N_22771,N_22131,N_22153);
or U22772 (N_22772,N_21672,N_21740);
nor U22773 (N_22773,N_21740,N_21679);
or U22774 (N_22774,N_22125,N_21764);
nor U22775 (N_22775,N_21701,N_22189);
nor U22776 (N_22776,N_21680,N_22165);
xnor U22777 (N_22777,N_21700,N_22083);
nand U22778 (N_22778,N_21889,N_21930);
nor U22779 (N_22779,N_22193,N_22009);
and U22780 (N_22780,N_22058,N_22107);
and U22781 (N_22781,N_22142,N_21776);
and U22782 (N_22782,N_22097,N_21768);
nand U22783 (N_22783,N_21930,N_21777);
and U22784 (N_22784,N_21998,N_21854);
nor U22785 (N_22785,N_21751,N_21987);
nand U22786 (N_22786,N_21685,N_21932);
xnor U22787 (N_22787,N_21629,N_22040);
or U22788 (N_22788,N_21657,N_21812);
nor U22789 (N_22789,N_21979,N_22044);
or U22790 (N_22790,N_22085,N_21704);
and U22791 (N_22791,N_21953,N_22096);
or U22792 (N_22792,N_21939,N_21803);
or U22793 (N_22793,N_21733,N_21660);
and U22794 (N_22794,N_21885,N_22174);
or U22795 (N_22795,N_21812,N_21625);
nor U22796 (N_22796,N_21961,N_22016);
or U22797 (N_22797,N_21740,N_22115);
and U22798 (N_22798,N_21750,N_21833);
or U22799 (N_22799,N_21818,N_21756);
nand U22800 (N_22800,N_22585,N_22512);
xnor U22801 (N_22801,N_22457,N_22525);
nor U22802 (N_22802,N_22355,N_22578);
nand U22803 (N_22803,N_22269,N_22752);
xor U22804 (N_22804,N_22539,N_22491);
and U22805 (N_22805,N_22440,N_22348);
and U22806 (N_22806,N_22568,N_22679);
or U22807 (N_22807,N_22455,N_22729);
xor U22808 (N_22808,N_22330,N_22765);
xnor U22809 (N_22809,N_22774,N_22763);
xnor U22810 (N_22810,N_22597,N_22283);
nor U22811 (N_22811,N_22481,N_22308);
nand U22812 (N_22812,N_22604,N_22490);
or U22813 (N_22813,N_22452,N_22533);
nand U22814 (N_22814,N_22767,N_22785);
or U22815 (N_22815,N_22246,N_22621);
and U22816 (N_22816,N_22319,N_22587);
and U22817 (N_22817,N_22248,N_22221);
nor U22818 (N_22818,N_22636,N_22385);
nand U22819 (N_22819,N_22418,N_22462);
or U22820 (N_22820,N_22227,N_22312);
and U22821 (N_22821,N_22356,N_22697);
nand U22822 (N_22822,N_22438,N_22640);
and U22823 (N_22823,N_22701,N_22476);
nor U22824 (N_22824,N_22734,N_22324);
xnor U22825 (N_22825,N_22793,N_22625);
nand U22826 (N_22826,N_22673,N_22505);
and U22827 (N_22827,N_22523,N_22226);
and U22828 (N_22828,N_22725,N_22721);
and U22829 (N_22829,N_22419,N_22633);
xor U22830 (N_22830,N_22428,N_22754);
and U22831 (N_22831,N_22635,N_22304);
nor U22832 (N_22832,N_22574,N_22486);
nand U22833 (N_22833,N_22396,N_22557);
xnor U22834 (N_22834,N_22708,N_22589);
nor U22835 (N_22835,N_22688,N_22572);
and U22836 (N_22836,N_22658,N_22655);
and U22837 (N_22837,N_22427,N_22397);
nand U22838 (N_22838,N_22576,N_22593);
and U22839 (N_22839,N_22219,N_22443);
nand U22840 (N_22840,N_22249,N_22584);
nor U22841 (N_22841,N_22493,N_22750);
or U22842 (N_22842,N_22445,N_22607);
and U22843 (N_22843,N_22497,N_22757);
nor U22844 (N_22844,N_22361,N_22535);
or U22845 (N_22845,N_22739,N_22732);
xnor U22846 (N_22846,N_22284,N_22528);
xnor U22847 (N_22847,N_22360,N_22748);
and U22848 (N_22848,N_22511,N_22614);
and U22849 (N_22849,N_22606,N_22233);
nor U22850 (N_22850,N_22513,N_22494);
nor U22851 (N_22851,N_22292,N_22524);
or U22852 (N_22852,N_22676,N_22345);
nand U22853 (N_22853,N_22693,N_22617);
or U22854 (N_22854,N_22579,N_22403);
xor U22855 (N_22855,N_22600,N_22482);
nand U22856 (N_22856,N_22619,N_22791);
and U22857 (N_22857,N_22276,N_22260);
nor U22858 (N_22858,N_22517,N_22254);
or U22859 (N_22859,N_22660,N_22464);
nor U22860 (N_22860,N_22352,N_22797);
xnor U22861 (N_22861,N_22700,N_22434);
and U22862 (N_22862,N_22646,N_22545);
nor U22863 (N_22863,N_22777,N_22424);
nand U22864 (N_22864,N_22288,N_22372);
xnor U22865 (N_22865,N_22258,N_22740);
nor U22866 (N_22866,N_22310,N_22690);
or U22867 (N_22867,N_22442,N_22240);
and U22868 (N_22868,N_22277,N_22451);
xnor U22869 (N_22869,N_22780,N_22703);
nor U22870 (N_22870,N_22205,N_22376);
and U22871 (N_22871,N_22390,N_22668);
and U22872 (N_22872,N_22799,N_22723);
nor U22873 (N_22873,N_22544,N_22571);
xor U22874 (N_22874,N_22437,N_22650);
xor U22875 (N_22875,N_22425,N_22598);
nand U22876 (N_22876,N_22622,N_22549);
nand U22877 (N_22877,N_22569,N_22346);
or U22878 (N_22878,N_22521,N_22235);
nand U22879 (N_22879,N_22328,N_22641);
xor U22880 (N_22880,N_22720,N_22753);
and U22881 (N_22881,N_22272,N_22689);
xnor U22882 (N_22882,N_22247,N_22466);
and U22883 (N_22883,N_22303,N_22685);
and U22884 (N_22884,N_22210,N_22514);
nand U22885 (N_22885,N_22558,N_22731);
nor U22886 (N_22886,N_22506,N_22415);
nor U22887 (N_22887,N_22699,N_22762);
nor U22888 (N_22888,N_22648,N_22379);
and U22889 (N_22889,N_22702,N_22215);
nand U22890 (N_22890,N_22592,N_22499);
and U22891 (N_22891,N_22392,N_22294);
or U22892 (N_22892,N_22522,N_22423);
or U22893 (N_22893,N_22488,N_22567);
xor U22894 (N_22894,N_22792,N_22552);
xor U22895 (N_22895,N_22575,N_22296);
xnor U22896 (N_22896,N_22719,N_22639);
nor U22897 (N_22897,N_22331,N_22766);
nand U22898 (N_22898,N_22461,N_22550);
nor U22899 (N_22899,N_22231,N_22588);
xor U22900 (N_22900,N_22469,N_22208);
nor U22901 (N_22901,N_22484,N_22630);
xor U22902 (N_22902,N_22787,N_22237);
xor U22903 (N_22903,N_22228,N_22479);
and U22904 (N_22904,N_22322,N_22282);
nand U22905 (N_22905,N_22480,N_22412);
and U22906 (N_22906,N_22323,N_22760);
and U22907 (N_22907,N_22782,N_22239);
nor U22908 (N_22908,N_22402,N_22562);
nor U22909 (N_22909,N_22783,N_22665);
or U22910 (N_22910,N_22381,N_22671);
xor U22911 (N_22911,N_22460,N_22678);
and U22912 (N_22912,N_22620,N_22370);
nor U22913 (N_22913,N_22315,N_22200);
nor U22914 (N_22914,N_22580,N_22244);
or U22915 (N_22915,N_22431,N_22386);
nor U22916 (N_22916,N_22382,N_22662);
and U22917 (N_22917,N_22744,N_22314);
and U22918 (N_22918,N_22264,N_22623);
xor U22919 (N_22919,N_22353,N_22771);
and U22920 (N_22920,N_22610,N_22224);
nor U22921 (N_22921,N_22709,N_22770);
nand U22922 (N_22922,N_22682,N_22285);
nor U22923 (N_22923,N_22629,N_22691);
or U22924 (N_22924,N_22798,N_22408);
or U22925 (N_22925,N_22642,N_22238);
xor U22926 (N_22926,N_22243,N_22516);
nand U22927 (N_22927,N_22686,N_22616);
nand U22928 (N_22928,N_22295,N_22540);
nand U22929 (N_22929,N_22764,N_22400);
or U22930 (N_22930,N_22632,N_22391);
nand U22931 (N_22931,N_22320,N_22422);
or U22932 (N_22932,N_22393,N_22223);
and U22933 (N_22933,N_22795,N_22500);
nand U22934 (N_22934,N_22374,N_22465);
nor U22935 (N_22935,N_22775,N_22738);
or U22936 (N_22936,N_22339,N_22316);
nand U22937 (N_22937,N_22297,N_22559);
nor U22938 (N_22938,N_22326,N_22548);
nor U22939 (N_22939,N_22344,N_22496);
nor U22940 (N_22940,N_22667,N_22745);
xor U22941 (N_22941,N_22664,N_22649);
xor U22942 (N_22942,N_22212,N_22713);
xor U22943 (N_22943,N_22281,N_22541);
or U22944 (N_22944,N_22242,N_22204);
nor U22945 (N_22945,N_22551,N_22519);
nand U22946 (N_22946,N_22354,N_22430);
nand U22947 (N_22947,N_22608,N_22270);
nand U22948 (N_22948,N_22234,N_22410);
or U22949 (N_22949,N_22309,N_22463);
xnor U22950 (N_22950,N_22776,N_22426);
nor U22951 (N_22951,N_22784,N_22216);
nor U22952 (N_22952,N_22201,N_22542);
xnor U22953 (N_22953,N_22680,N_22417);
and U22954 (N_22954,N_22411,N_22279);
and U22955 (N_22955,N_22388,N_22458);
and U22956 (N_22956,N_22229,N_22778);
xor U22957 (N_22957,N_22577,N_22526);
or U22958 (N_22958,N_22436,N_22715);
or U22959 (N_22959,N_22265,N_22409);
xnor U22960 (N_22960,N_22478,N_22251);
nor U22961 (N_22961,N_22489,N_22538);
nand U22962 (N_22962,N_22380,N_22341);
and U22963 (N_22963,N_22357,N_22599);
or U22964 (N_22964,N_22786,N_22718);
nand U22965 (N_22965,N_22217,N_22332);
and U22966 (N_22966,N_22651,N_22756);
or U22967 (N_22967,N_22564,N_22278);
or U22968 (N_22968,N_22759,N_22573);
nor U22969 (N_22969,N_22647,N_22214);
xor U22970 (N_22970,N_22300,N_22373);
nor U22971 (N_22971,N_22218,N_22325);
or U22972 (N_22972,N_22448,N_22675);
or U22973 (N_22973,N_22362,N_22444);
nand U22974 (N_22974,N_22327,N_22358);
nand U22975 (N_22975,N_22439,N_22267);
nor U22976 (N_22976,N_22547,N_22416);
nand U22977 (N_22977,N_22624,N_22586);
nor U22978 (N_22978,N_22730,N_22203);
xnor U22979 (N_22979,N_22518,N_22405);
or U22980 (N_22980,N_22634,N_22727);
xor U22981 (N_22981,N_22274,N_22726);
and U22982 (N_22982,N_22298,N_22611);
nor U22983 (N_22983,N_22746,N_22613);
nand U22984 (N_22984,N_22363,N_22565);
xor U22985 (N_22985,N_22681,N_22749);
and U22986 (N_22986,N_22241,N_22475);
xnor U22987 (N_22987,N_22710,N_22663);
nor U22988 (N_22988,N_22566,N_22626);
nand U22989 (N_22989,N_22507,N_22275);
or U22990 (N_22990,N_22378,N_22515);
and U22991 (N_22991,N_22334,N_22601);
nand U22992 (N_22992,N_22206,N_22395);
nor U22993 (N_22993,N_22307,N_22446);
xor U22994 (N_22994,N_22696,N_22609);
and U22995 (N_22995,N_22377,N_22329);
nand U22996 (N_22996,N_22311,N_22259);
nand U22997 (N_22997,N_22692,N_22333);
xnor U22998 (N_22998,N_22594,N_22368);
or U22999 (N_22999,N_22383,N_22672);
and U23000 (N_23000,N_22706,N_22483);
or U23001 (N_23001,N_22794,N_22302);
nor U23002 (N_23002,N_22659,N_22485);
or U23003 (N_23003,N_22364,N_22456);
nor U23004 (N_23004,N_22349,N_22318);
or U23005 (N_23005,N_22751,N_22470);
or U23006 (N_23006,N_22728,N_22340);
and U23007 (N_23007,N_22705,N_22435);
and U23008 (N_23008,N_22406,N_22652);
and U23009 (N_23009,N_22398,N_22342);
and U23010 (N_23010,N_22714,N_22273);
and U23011 (N_23011,N_22543,N_22306);
nand U23012 (N_23012,N_22474,N_22503);
nor U23013 (N_23013,N_22637,N_22367);
nor U23014 (N_23014,N_22769,N_22789);
and U23015 (N_23015,N_22472,N_22560);
nand U23016 (N_23016,N_22250,N_22399);
xor U23017 (N_23017,N_22755,N_22501);
xnor U23018 (N_23018,N_22387,N_22694);
nor U23019 (N_23019,N_22401,N_22220);
nor U23020 (N_23020,N_22553,N_22321);
and U23021 (N_23021,N_22656,N_22527);
and U23022 (N_23022,N_22413,N_22643);
xnor U23023 (N_23023,N_22450,N_22737);
nand U23024 (N_23024,N_22618,N_22781);
nor U23025 (N_23025,N_22202,N_22266);
xnor U23026 (N_23026,N_22293,N_22317);
nand U23027 (N_23027,N_22603,N_22209);
nand U23028 (N_23028,N_22790,N_22628);
nor U23029 (N_23029,N_22590,N_22773);
and U23030 (N_23030,N_22271,N_22747);
or U23031 (N_23031,N_22669,N_22495);
nor U23032 (N_23032,N_22245,N_22530);
nand U23033 (N_23033,N_22256,N_22529);
nor U23034 (N_23034,N_22447,N_22627);
nor U23035 (N_23035,N_22291,N_22359);
xnor U23036 (N_23036,N_22467,N_22432);
or U23037 (N_23037,N_22449,N_22638);
nand U23038 (N_23038,N_22563,N_22779);
and U23039 (N_23039,N_22742,N_22645);
or U23040 (N_23040,N_22369,N_22561);
nor U23041 (N_23041,N_22225,N_22429);
nor U23042 (N_23042,N_22612,N_22741);
xnor U23043 (N_23043,N_22421,N_22704);
and U23044 (N_23044,N_22657,N_22581);
nor U23045 (N_23045,N_22520,N_22365);
and U23046 (N_23046,N_22335,N_22602);
nor U23047 (N_23047,N_22257,N_22743);
or U23048 (N_23048,N_22487,N_22509);
or U23049 (N_23049,N_22596,N_22687);
and U23050 (N_23050,N_22252,N_22532);
nand U23051 (N_23051,N_22375,N_22394);
nor U23052 (N_23052,N_22498,N_22631);
and U23053 (N_23053,N_22684,N_22351);
nand U23054 (N_23054,N_22280,N_22471);
and U23055 (N_23055,N_22289,N_22644);
xnor U23056 (N_23056,N_22453,N_22707);
or U23057 (N_23057,N_22414,N_22468);
nand U23058 (N_23058,N_22459,N_22232);
nand U23059 (N_23059,N_22290,N_22261);
xor U23060 (N_23060,N_22313,N_22554);
and U23061 (N_23061,N_22695,N_22716);
or U23062 (N_23062,N_22537,N_22768);
xnor U23063 (N_23063,N_22717,N_22531);
and U23064 (N_23064,N_22211,N_22712);
or U23065 (N_23065,N_22736,N_22473);
nand U23066 (N_23066,N_22796,N_22722);
and U23067 (N_23067,N_22222,N_22477);
or U23068 (N_23068,N_22677,N_22761);
or U23069 (N_23069,N_22591,N_22724);
and U23070 (N_23070,N_22299,N_22733);
or U23071 (N_23071,N_22653,N_22711);
and U23072 (N_23072,N_22268,N_22263);
and U23073 (N_23073,N_22583,N_22389);
nand U23074 (N_23074,N_22758,N_22262);
nand U23075 (N_23075,N_22337,N_22556);
nand U23076 (N_23076,N_22347,N_22433);
and U23077 (N_23077,N_22255,N_22454);
and U23078 (N_23078,N_22504,N_22683);
nor U23079 (N_23079,N_22366,N_22287);
nand U23080 (N_23080,N_22336,N_22305);
and U23081 (N_23081,N_22615,N_22508);
nor U23082 (N_23082,N_22788,N_22772);
nor U23083 (N_23083,N_22536,N_22605);
nor U23084 (N_23084,N_22407,N_22546);
and U23085 (N_23085,N_22213,N_22502);
and U23086 (N_23086,N_22236,N_22404);
or U23087 (N_23087,N_22674,N_22301);
nor U23088 (N_23088,N_22350,N_22661);
nor U23089 (N_23089,N_22286,N_22666);
nor U23090 (N_23090,N_22371,N_22253);
nand U23091 (N_23091,N_22492,N_22420);
nor U23092 (N_23092,N_22343,N_22735);
nand U23093 (N_23093,N_22698,N_22441);
xor U23094 (N_23094,N_22670,N_22595);
and U23095 (N_23095,N_22582,N_22570);
and U23096 (N_23096,N_22534,N_22654);
and U23097 (N_23097,N_22555,N_22230);
nand U23098 (N_23098,N_22207,N_22338);
or U23099 (N_23099,N_22510,N_22384);
and U23100 (N_23100,N_22386,N_22490);
and U23101 (N_23101,N_22497,N_22786);
nor U23102 (N_23102,N_22735,N_22476);
and U23103 (N_23103,N_22246,N_22450);
nand U23104 (N_23104,N_22451,N_22666);
and U23105 (N_23105,N_22511,N_22461);
or U23106 (N_23106,N_22510,N_22702);
and U23107 (N_23107,N_22461,N_22702);
nand U23108 (N_23108,N_22413,N_22745);
nor U23109 (N_23109,N_22538,N_22498);
and U23110 (N_23110,N_22283,N_22393);
and U23111 (N_23111,N_22561,N_22341);
and U23112 (N_23112,N_22297,N_22639);
xnor U23113 (N_23113,N_22369,N_22675);
nand U23114 (N_23114,N_22252,N_22741);
xnor U23115 (N_23115,N_22712,N_22204);
or U23116 (N_23116,N_22215,N_22480);
xor U23117 (N_23117,N_22489,N_22696);
xnor U23118 (N_23118,N_22310,N_22348);
xnor U23119 (N_23119,N_22740,N_22436);
nor U23120 (N_23120,N_22616,N_22693);
nor U23121 (N_23121,N_22384,N_22798);
nor U23122 (N_23122,N_22517,N_22337);
nand U23123 (N_23123,N_22234,N_22467);
and U23124 (N_23124,N_22713,N_22729);
nand U23125 (N_23125,N_22647,N_22558);
xnor U23126 (N_23126,N_22410,N_22388);
or U23127 (N_23127,N_22323,N_22324);
nor U23128 (N_23128,N_22377,N_22441);
xnor U23129 (N_23129,N_22280,N_22360);
or U23130 (N_23130,N_22240,N_22746);
nor U23131 (N_23131,N_22443,N_22391);
nor U23132 (N_23132,N_22425,N_22466);
or U23133 (N_23133,N_22467,N_22243);
and U23134 (N_23134,N_22384,N_22514);
nor U23135 (N_23135,N_22344,N_22575);
nand U23136 (N_23136,N_22247,N_22373);
and U23137 (N_23137,N_22378,N_22236);
or U23138 (N_23138,N_22749,N_22798);
and U23139 (N_23139,N_22213,N_22324);
xor U23140 (N_23140,N_22513,N_22320);
nand U23141 (N_23141,N_22489,N_22343);
or U23142 (N_23142,N_22330,N_22486);
and U23143 (N_23143,N_22388,N_22763);
nor U23144 (N_23144,N_22662,N_22650);
and U23145 (N_23145,N_22370,N_22705);
nor U23146 (N_23146,N_22781,N_22281);
nor U23147 (N_23147,N_22669,N_22493);
or U23148 (N_23148,N_22439,N_22208);
and U23149 (N_23149,N_22574,N_22491);
nor U23150 (N_23150,N_22746,N_22325);
nor U23151 (N_23151,N_22249,N_22471);
nor U23152 (N_23152,N_22306,N_22485);
nand U23153 (N_23153,N_22207,N_22563);
xnor U23154 (N_23154,N_22684,N_22572);
and U23155 (N_23155,N_22639,N_22444);
and U23156 (N_23156,N_22618,N_22220);
xnor U23157 (N_23157,N_22386,N_22225);
xor U23158 (N_23158,N_22714,N_22286);
xnor U23159 (N_23159,N_22584,N_22655);
xor U23160 (N_23160,N_22601,N_22626);
and U23161 (N_23161,N_22367,N_22532);
nor U23162 (N_23162,N_22429,N_22674);
and U23163 (N_23163,N_22698,N_22539);
xnor U23164 (N_23164,N_22363,N_22207);
and U23165 (N_23165,N_22409,N_22351);
or U23166 (N_23166,N_22235,N_22643);
nand U23167 (N_23167,N_22647,N_22523);
and U23168 (N_23168,N_22332,N_22788);
nor U23169 (N_23169,N_22289,N_22720);
or U23170 (N_23170,N_22561,N_22647);
or U23171 (N_23171,N_22763,N_22771);
nor U23172 (N_23172,N_22215,N_22498);
or U23173 (N_23173,N_22731,N_22488);
and U23174 (N_23174,N_22343,N_22330);
xnor U23175 (N_23175,N_22654,N_22589);
nand U23176 (N_23176,N_22450,N_22423);
nor U23177 (N_23177,N_22387,N_22487);
xnor U23178 (N_23178,N_22278,N_22352);
xor U23179 (N_23179,N_22436,N_22384);
or U23180 (N_23180,N_22358,N_22243);
nand U23181 (N_23181,N_22366,N_22530);
or U23182 (N_23182,N_22255,N_22380);
or U23183 (N_23183,N_22458,N_22754);
nand U23184 (N_23184,N_22762,N_22558);
nand U23185 (N_23185,N_22534,N_22652);
xnor U23186 (N_23186,N_22343,N_22645);
nor U23187 (N_23187,N_22207,N_22629);
nand U23188 (N_23188,N_22669,N_22581);
and U23189 (N_23189,N_22765,N_22551);
nand U23190 (N_23190,N_22589,N_22788);
and U23191 (N_23191,N_22591,N_22208);
or U23192 (N_23192,N_22494,N_22590);
and U23193 (N_23193,N_22675,N_22429);
nand U23194 (N_23194,N_22407,N_22442);
and U23195 (N_23195,N_22640,N_22684);
xnor U23196 (N_23196,N_22251,N_22318);
nand U23197 (N_23197,N_22765,N_22414);
nor U23198 (N_23198,N_22729,N_22261);
or U23199 (N_23199,N_22752,N_22605);
nor U23200 (N_23200,N_22464,N_22282);
or U23201 (N_23201,N_22472,N_22442);
nor U23202 (N_23202,N_22566,N_22657);
or U23203 (N_23203,N_22454,N_22766);
nand U23204 (N_23204,N_22479,N_22642);
and U23205 (N_23205,N_22239,N_22514);
nor U23206 (N_23206,N_22519,N_22355);
or U23207 (N_23207,N_22616,N_22403);
nor U23208 (N_23208,N_22494,N_22645);
or U23209 (N_23209,N_22486,N_22320);
or U23210 (N_23210,N_22357,N_22588);
nand U23211 (N_23211,N_22585,N_22479);
xor U23212 (N_23212,N_22781,N_22271);
nor U23213 (N_23213,N_22396,N_22798);
xor U23214 (N_23214,N_22398,N_22668);
or U23215 (N_23215,N_22327,N_22452);
xor U23216 (N_23216,N_22222,N_22791);
nand U23217 (N_23217,N_22713,N_22374);
and U23218 (N_23218,N_22614,N_22204);
or U23219 (N_23219,N_22417,N_22573);
or U23220 (N_23220,N_22744,N_22382);
or U23221 (N_23221,N_22594,N_22259);
and U23222 (N_23222,N_22401,N_22480);
and U23223 (N_23223,N_22354,N_22351);
xnor U23224 (N_23224,N_22774,N_22268);
and U23225 (N_23225,N_22734,N_22334);
or U23226 (N_23226,N_22278,N_22284);
or U23227 (N_23227,N_22533,N_22755);
nor U23228 (N_23228,N_22434,N_22464);
nand U23229 (N_23229,N_22349,N_22428);
and U23230 (N_23230,N_22217,N_22765);
nor U23231 (N_23231,N_22769,N_22526);
or U23232 (N_23232,N_22446,N_22296);
nand U23233 (N_23233,N_22572,N_22583);
nor U23234 (N_23234,N_22735,N_22310);
xnor U23235 (N_23235,N_22467,N_22569);
or U23236 (N_23236,N_22432,N_22726);
nor U23237 (N_23237,N_22573,N_22274);
nand U23238 (N_23238,N_22475,N_22448);
nor U23239 (N_23239,N_22576,N_22363);
or U23240 (N_23240,N_22651,N_22740);
xor U23241 (N_23241,N_22676,N_22576);
nor U23242 (N_23242,N_22538,N_22670);
and U23243 (N_23243,N_22329,N_22689);
or U23244 (N_23244,N_22598,N_22378);
xor U23245 (N_23245,N_22766,N_22597);
nand U23246 (N_23246,N_22738,N_22487);
xnor U23247 (N_23247,N_22564,N_22637);
nand U23248 (N_23248,N_22767,N_22526);
and U23249 (N_23249,N_22328,N_22231);
or U23250 (N_23250,N_22357,N_22351);
xor U23251 (N_23251,N_22332,N_22484);
and U23252 (N_23252,N_22751,N_22646);
nor U23253 (N_23253,N_22684,N_22489);
nand U23254 (N_23254,N_22467,N_22341);
nand U23255 (N_23255,N_22493,N_22430);
and U23256 (N_23256,N_22527,N_22487);
xor U23257 (N_23257,N_22360,N_22630);
and U23258 (N_23258,N_22547,N_22446);
nor U23259 (N_23259,N_22368,N_22330);
nand U23260 (N_23260,N_22286,N_22233);
nor U23261 (N_23261,N_22252,N_22419);
nor U23262 (N_23262,N_22590,N_22701);
and U23263 (N_23263,N_22586,N_22583);
or U23264 (N_23264,N_22288,N_22363);
or U23265 (N_23265,N_22694,N_22365);
nor U23266 (N_23266,N_22758,N_22416);
xor U23267 (N_23267,N_22574,N_22356);
nor U23268 (N_23268,N_22283,N_22482);
or U23269 (N_23269,N_22500,N_22796);
nor U23270 (N_23270,N_22315,N_22605);
and U23271 (N_23271,N_22231,N_22356);
and U23272 (N_23272,N_22617,N_22700);
nor U23273 (N_23273,N_22488,N_22281);
and U23274 (N_23274,N_22743,N_22500);
nor U23275 (N_23275,N_22720,N_22568);
nand U23276 (N_23276,N_22625,N_22575);
nor U23277 (N_23277,N_22752,N_22313);
or U23278 (N_23278,N_22724,N_22314);
nor U23279 (N_23279,N_22627,N_22244);
xnor U23280 (N_23280,N_22697,N_22369);
and U23281 (N_23281,N_22316,N_22781);
xnor U23282 (N_23282,N_22557,N_22382);
or U23283 (N_23283,N_22654,N_22785);
or U23284 (N_23284,N_22772,N_22596);
and U23285 (N_23285,N_22778,N_22429);
nand U23286 (N_23286,N_22421,N_22652);
or U23287 (N_23287,N_22287,N_22421);
xnor U23288 (N_23288,N_22622,N_22730);
nor U23289 (N_23289,N_22596,N_22373);
and U23290 (N_23290,N_22698,N_22374);
nand U23291 (N_23291,N_22332,N_22705);
and U23292 (N_23292,N_22690,N_22594);
nor U23293 (N_23293,N_22351,N_22517);
and U23294 (N_23294,N_22444,N_22689);
nor U23295 (N_23295,N_22266,N_22624);
or U23296 (N_23296,N_22375,N_22477);
nand U23297 (N_23297,N_22483,N_22414);
nand U23298 (N_23298,N_22566,N_22736);
nor U23299 (N_23299,N_22322,N_22769);
nor U23300 (N_23300,N_22356,N_22511);
xnor U23301 (N_23301,N_22350,N_22675);
or U23302 (N_23302,N_22301,N_22682);
and U23303 (N_23303,N_22412,N_22765);
nor U23304 (N_23304,N_22431,N_22571);
nor U23305 (N_23305,N_22627,N_22718);
nand U23306 (N_23306,N_22662,N_22575);
and U23307 (N_23307,N_22338,N_22440);
xor U23308 (N_23308,N_22664,N_22282);
nor U23309 (N_23309,N_22281,N_22269);
xor U23310 (N_23310,N_22244,N_22734);
nand U23311 (N_23311,N_22747,N_22405);
and U23312 (N_23312,N_22446,N_22336);
or U23313 (N_23313,N_22335,N_22542);
xnor U23314 (N_23314,N_22637,N_22467);
and U23315 (N_23315,N_22783,N_22539);
xor U23316 (N_23316,N_22644,N_22616);
and U23317 (N_23317,N_22330,N_22515);
nor U23318 (N_23318,N_22757,N_22482);
xor U23319 (N_23319,N_22698,N_22618);
nor U23320 (N_23320,N_22429,N_22431);
or U23321 (N_23321,N_22719,N_22395);
or U23322 (N_23322,N_22388,N_22725);
or U23323 (N_23323,N_22512,N_22760);
nor U23324 (N_23324,N_22763,N_22389);
nand U23325 (N_23325,N_22470,N_22431);
nor U23326 (N_23326,N_22440,N_22663);
and U23327 (N_23327,N_22320,N_22730);
xnor U23328 (N_23328,N_22633,N_22606);
xor U23329 (N_23329,N_22687,N_22532);
nand U23330 (N_23330,N_22691,N_22569);
nand U23331 (N_23331,N_22229,N_22298);
nand U23332 (N_23332,N_22616,N_22243);
and U23333 (N_23333,N_22525,N_22337);
nand U23334 (N_23334,N_22599,N_22447);
and U23335 (N_23335,N_22509,N_22443);
xor U23336 (N_23336,N_22226,N_22442);
nor U23337 (N_23337,N_22746,N_22493);
nand U23338 (N_23338,N_22581,N_22450);
xnor U23339 (N_23339,N_22652,N_22665);
nand U23340 (N_23340,N_22211,N_22318);
or U23341 (N_23341,N_22539,N_22718);
or U23342 (N_23342,N_22310,N_22751);
and U23343 (N_23343,N_22255,N_22461);
and U23344 (N_23344,N_22240,N_22744);
and U23345 (N_23345,N_22785,N_22622);
or U23346 (N_23346,N_22241,N_22238);
xor U23347 (N_23347,N_22280,N_22270);
nand U23348 (N_23348,N_22786,N_22735);
xor U23349 (N_23349,N_22229,N_22476);
and U23350 (N_23350,N_22506,N_22380);
or U23351 (N_23351,N_22303,N_22244);
or U23352 (N_23352,N_22228,N_22509);
nor U23353 (N_23353,N_22553,N_22322);
and U23354 (N_23354,N_22449,N_22522);
and U23355 (N_23355,N_22581,N_22410);
or U23356 (N_23356,N_22624,N_22476);
nor U23357 (N_23357,N_22223,N_22508);
xor U23358 (N_23358,N_22244,N_22769);
xnor U23359 (N_23359,N_22676,N_22427);
nor U23360 (N_23360,N_22724,N_22331);
xnor U23361 (N_23361,N_22793,N_22449);
and U23362 (N_23362,N_22311,N_22471);
nand U23363 (N_23363,N_22794,N_22473);
nand U23364 (N_23364,N_22212,N_22221);
xor U23365 (N_23365,N_22453,N_22663);
nand U23366 (N_23366,N_22693,N_22697);
nand U23367 (N_23367,N_22233,N_22417);
nand U23368 (N_23368,N_22793,N_22582);
nor U23369 (N_23369,N_22441,N_22240);
nor U23370 (N_23370,N_22675,N_22214);
nand U23371 (N_23371,N_22565,N_22500);
and U23372 (N_23372,N_22345,N_22763);
and U23373 (N_23373,N_22784,N_22473);
nand U23374 (N_23374,N_22777,N_22248);
nand U23375 (N_23375,N_22586,N_22701);
xnor U23376 (N_23376,N_22538,N_22229);
nand U23377 (N_23377,N_22433,N_22715);
and U23378 (N_23378,N_22619,N_22747);
nor U23379 (N_23379,N_22598,N_22326);
and U23380 (N_23380,N_22772,N_22219);
nor U23381 (N_23381,N_22692,N_22276);
nor U23382 (N_23382,N_22510,N_22552);
nand U23383 (N_23383,N_22788,N_22609);
and U23384 (N_23384,N_22506,N_22250);
xnor U23385 (N_23385,N_22322,N_22672);
nand U23386 (N_23386,N_22416,N_22230);
xor U23387 (N_23387,N_22402,N_22627);
and U23388 (N_23388,N_22754,N_22249);
xnor U23389 (N_23389,N_22391,N_22357);
nor U23390 (N_23390,N_22527,N_22218);
or U23391 (N_23391,N_22341,N_22662);
nand U23392 (N_23392,N_22445,N_22491);
and U23393 (N_23393,N_22440,N_22785);
xor U23394 (N_23394,N_22359,N_22280);
and U23395 (N_23395,N_22786,N_22532);
nor U23396 (N_23396,N_22720,N_22572);
or U23397 (N_23397,N_22401,N_22554);
or U23398 (N_23398,N_22265,N_22773);
and U23399 (N_23399,N_22373,N_22534);
xor U23400 (N_23400,N_23139,N_23083);
nor U23401 (N_23401,N_23085,N_23326);
or U23402 (N_23402,N_22926,N_22800);
and U23403 (N_23403,N_23192,N_23340);
xnor U23404 (N_23404,N_22807,N_22973);
or U23405 (N_23405,N_23271,N_23319);
or U23406 (N_23406,N_23124,N_22806);
and U23407 (N_23407,N_23067,N_23213);
nand U23408 (N_23408,N_22801,N_22820);
and U23409 (N_23409,N_23351,N_22898);
xnor U23410 (N_23410,N_23395,N_23365);
and U23411 (N_23411,N_23148,N_22963);
and U23412 (N_23412,N_23211,N_23047);
nor U23413 (N_23413,N_23380,N_23277);
xnor U23414 (N_23414,N_23250,N_22860);
xnor U23415 (N_23415,N_23002,N_23115);
and U23416 (N_23416,N_23074,N_23038);
xor U23417 (N_23417,N_23332,N_23204);
xor U23418 (N_23418,N_23007,N_22941);
or U23419 (N_23419,N_22974,N_22985);
or U23420 (N_23420,N_23011,N_23033);
nor U23421 (N_23421,N_22938,N_22904);
nor U23422 (N_23422,N_22982,N_23249);
nor U23423 (N_23423,N_23082,N_23255);
and U23424 (N_23424,N_23162,N_22864);
xor U23425 (N_23425,N_22816,N_23164);
xnor U23426 (N_23426,N_22840,N_22825);
nor U23427 (N_23427,N_23168,N_23086);
and U23428 (N_23428,N_22879,N_22895);
and U23429 (N_23429,N_23137,N_23110);
or U23430 (N_23430,N_23344,N_23101);
or U23431 (N_23431,N_23312,N_23034);
xor U23432 (N_23432,N_23366,N_22949);
and U23433 (N_23433,N_22869,N_22900);
nor U23434 (N_23434,N_23203,N_23237);
xor U23435 (N_23435,N_23309,N_23088);
and U23436 (N_23436,N_23031,N_23313);
nor U23437 (N_23437,N_22843,N_23129);
xnor U23438 (N_23438,N_23235,N_23079);
or U23439 (N_23439,N_23132,N_22835);
nor U23440 (N_23440,N_23108,N_23364);
or U23441 (N_23441,N_23353,N_22964);
nor U23442 (N_23442,N_23144,N_23356);
and U23443 (N_23443,N_22855,N_22833);
and U23444 (N_23444,N_23315,N_22813);
nor U23445 (N_23445,N_23143,N_23343);
or U23446 (N_23446,N_23260,N_23274);
nor U23447 (N_23447,N_23111,N_23342);
or U23448 (N_23448,N_22922,N_23258);
or U23449 (N_23449,N_23102,N_23278);
nor U23450 (N_23450,N_22810,N_23140);
or U23451 (N_23451,N_23024,N_23217);
nand U23452 (N_23452,N_23321,N_23292);
and U23453 (N_23453,N_22814,N_23003);
nor U23454 (N_23454,N_23265,N_23163);
or U23455 (N_23455,N_23236,N_23021);
or U23456 (N_23456,N_23176,N_22874);
nand U23457 (N_23457,N_23092,N_23390);
nor U23458 (N_23458,N_23361,N_23050);
xnor U23459 (N_23459,N_23290,N_23109);
xnor U23460 (N_23460,N_23195,N_22978);
and U23461 (N_23461,N_23360,N_22858);
nand U23462 (N_23462,N_23284,N_23262);
and U23463 (N_23463,N_23149,N_23010);
and U23464 (N_23464,N_23205,N_23389);
or U23465 (N_23465,N_23374,N_23130);
or U23466 (N_23466,N_22880,N_23091);
xor U23467 (N_23467,N_23046,N_22892);
and U23468 (N_23468,N_23026,N_23141);
nand U23469 (N_23469,N_23378,N_22865);
and U23470 (N_23470,N_23329,N_23166);
xnor U23471 (N_23471,N_22862,N_22920);
or U23472 (N_23472,N_23081,N_23297);
nor U23473 (N_23473,N_22824,N_22931);
nor U23474 (N_23474,N_22822,N_22987);
nor U23475 (N_23475,N_23302,N_22834);
or U23476 (N_23476,N_22991,N_23397);
nand U23477 (N_23477,N_22805,N_22866);
nor U23478 (N_23478,N_23314,N_23293);
or U23479 (N_23479,N_22945,N_23275);
and U23480 (N_23480,N_23363,N_22950);
and U23481 (N_23481,N_22886,N_23349);
nand U23482 (N_23482,N_23207,N_22859);
nand U23483 (N_23483,N_22959,N_23198);
nand U23484 (N_23484,N_23125,N_22966);
nand U23485 (N_23485,N_23151,N_23379);
xor U23486 (N_23486,N_23068,N_23122);
nor U23487 (N_23487,N_23177,N_22925);
or U23488 (N_23488,N_22956,N_23385);
nor U23489 (N_23489,N_23269,N_22861);
or U23490 (N_23490,N_23208,N_23288);
xor U23491 (N_23491,N_22995,N_23063);
nand U23492 (N_23492,N_22986,N_22934);
nor U23493 (N_23493,N_23370,N_22850);
xor U23494 (N_23494,N_23223,N_22940);
xor U23495 (N_23495,N_23027,N_23280);
xnor U23496 (N_23496,N_22914,N_22854);
nor U23497 (N_23497,N_23387,N_23224);
nand U23498 (N_23498,N_23113,N_23099);
and U23499 (N_23499,N_22918,N_23214);
and U23500 (N_23500,N_23120,N_22811);
xor U23501 (N_23501,N_22836,N_23320);
nor U23502 (N_23502,N_22980,N_22911);
or U23503 (N_23503,N_23317,N_23335);
or U23504 (N_23504,N_22808,N_22952);
nand U23505 (N_23505,N_22916,N_23076);
and U23506 (N_23506,N_23042,N_23017);
or U23507 (N_23507,N_23308,N_22970);
or U23508 (N_23508,N_23221,N_23248);
nor U23509 (N_23509,N_23234,N_23306);
xor U23510 (N_23510,N_22829,N_23041);
xor U23511 (N_23511,N_23165,N_22888);
nand U23512 (N_23512,N_23327,N_22975);
or U23513 (N_23513,N_23362,N_22832);
and U23514 (N_23514,N_22981,N_22972);
or U23515 (N_23515,N_22983,N_23194);
nand U23516 (N_23516,N_23167,N_23106);
xnor U23517 (N_23517,N_23078,N_23368);
nand U23518 (N_23518,N_23283,N_23045);
nor U23519 (N_23519,N_22996,N_22872);
xnor U23520 (N_23520,N_22851,N_23231);
nand U23521 (N_23521,N_23253,N_23090);
or U23522 (N_23522,N_23218,N_23098);
nand U23523 (N_23523,N_23294,N_23105);
nor U23524 (N_23524,N_22933,N_22809);
and U23525 (N_23525,N_22988,N_22868);
nor U23526 (N_23526,N_22893,N_23393);
nand U23527 (N_23527,N_23094,N_23112);
nor U23528 (N_23528,N_22821,N_22883);
and U23529 (N_23529,N_23123,N_23240);
nor U23530 (N_23530,N_22881,N_23004);
xor U23531 (N_23531,N_23199,N_23065);
xor U23532 (N_23532,N_23295,N_23259);
nand U23533 (N_23533,N_22917,N_23187);
and U23534 (N_23534,N_23013,N_23341);
nor U23535 (N_23535,N_22944,N_23219);
or U23536 (N_23536,N_23398,N_22812);
and U23537 (N_23537,N_22932,N_23273);
nand U23538 (N_23538,N_23061,N_23044);
and U23539 (N_23539,N_22910,N_23336);
nor U23540 (N_23540,N_23348,N_23396);
nand U23541 (N_23541,N_23119,N_22803);
xnor U23542 (N_23542,N_23062,N_23300);
nor U23543 (N_23543,N_23037,N_23305);
and U23544 (N_23544,N_22876,N_23048);
and U23545 (N_23545,N_23324,N_23104);
nor U23546 (N_23546,N_23242,N_23333);
or U23547 (N_23547,N_23202,N_22894);
xnor U23548 (N_23548,N_23058,N_23241);
nor U23549 (N_23549,N_23000,N_22977);
xor U23550 (N_23550,N_23228,N_23225);
nand U23551 (N_23551,N_23029,N_22935);
and U23552 (N_23552,N_23247,N_23382);
and U23553 (N_23553,N_22849,N_22896);
nor U23554 (N_23554,N_23345,N_22817);
and U23555 (N_23555,N_23220,N_22908);
nand U23556 (N_23556,N_23136,N_22905);
and U23557 (N_23557,N_22847,N_23070);
nand U23558 (N_23558,N_23032,N_22942);
or U23559 (N_23559,N_22962,N_23286);
nor U23560 (N_23560,N_22857,N_23392);
xnor U23561 (N_23561,N_22903,N_23386);
and U23562 (N_23562,N_23006,N_23264);
and U23563 (N_23563,N_22936,N_23311);
and U23564 (N_23564,N_22841,N_23189);
nor U23565 (N_23565,N_23197,N_22902);
nor U23566 (N_23566,N_23135,N_23056);
or U23567 (N_23567,N_22971,N_23193);
and U23568 (N_23568,N_22984,N_22828);
or U23569 (N_23569,N_22939,N_23118);
nand U23570 (N_23570,N_22830,N_23150);
and U23571 (N_23571,N_23072,N_23084);
and U23572 (N_23572,N_22837,N_23337);
nor U23573 (N_23573,N_23210,N_23131);
xnor U23574 (N_23574,N_22955,N_23188);
nor U23575 (N_23575,N_23376,N_23054);
nand U23576 (N_23576,N_23191,N_23399);
nor U23577 (N_23577,N_23178,N_23229);
nor U23578 (N_23578,N_23239,N_22819);
nand U23579 (N_23579,N_22839,N_22853);
nand U23580 (N_23580,N_23388,N_23127);
nand U23581 (N_23581,N_23276,N_23075);
or U23582 (N_23582,N_22919,N_23161);
nand U23583 (N_23583,N_23051,N_22951);
nand U23584 (N_23584,N_23303,N_22946);
xnor U23585 (N_23585,N_23238,N_22915);
nand U23586 (N_23586,N_23121,N_23077);
xnor U23587 (N_23587,N_22943,N_23206);
nand U23588 (N_23588,N_23299,N_23049);
or U23589 (N_23589,N_23359,N_23172);
or U23590 (N_23590,N_22889,N_23226);
nor U23591 (N_23591,N_22826,N_22842);
xnor U23592 (N_23592,N_23158,N_23243);
nor U23593 (N_23593,N_23296,N_23355);
xnor U23594 (N_23594,N_23174,N_23212);
nand U23595 (N_23595,N_22969,N_23316);
or U23596 (N_23596,N_23175,N_23138);
and U23597 (N_23597,N_23023,N_23185);
or U23598 (N_23598,N_22961,N_23173);
xnor U23599 (N_23599,N_23028,N_22887);
and U23600 (N_23600,N_23018,N_23040);
xor U23601 (N_23601,N_22844,N_23330);
nor U23602 (N_23602,N_22815,N_22958);
nand U23603 (N_23603,N_22997,N_23272);
nand U23604 (N_23604,N_23036,N_23394);
nor U23605 (N_23605,N_23257,N_23096);
or U23606 (N_23606,N_23279,N_23145);
nor U23607 (N_23607,N_23268,N_23134);
nand U23608 (N_23608,N_23383,N_23254);
nor U23609 (N_23609,N_22965,N_23080);
or U23610 (N_23610,N_23093,N_22930);
xnor U23611 (N_23611,N_23153,N_23244);
or U23612 (N_23612,N_23357,N_23222);
and U23613 (N_23613,N_23001,N_23020);
or U23614 (N_23614,N_22827,N_23052);
and U23615 (N_23615,N_22968,N_22831);
and U23616 (N_23616,N_23128,N_22878);
or U23617 (N_23617,N_23155,N_23323);
and U23618 (N_23618,N_23022,N_23246);
and U23619 (N_23619,N_23200,N_23069);
and U23620 (N_23620,N_23377,N_23301);
xor U23621 (N_23621,N_23256,N_23180);
nand U23622 (N_23622,N_22882,N_23270);
nand U23623 (N_23623,N_23012,N_23350);
nand U23624 (N_23624,N_23227,N_23035);
nor U23625 (N_23625,N_23201,N_22989);
and U23626 (N_23626,N_22891,N_22990);
and U23627 (N_23627,N_23182,N_22998);
xnor U23628 (N_23628,N_23057,N_23373);
nand U23629 (N_23629,N_23066,N_23015);
and U23630 (N_23630,N_23116,N_22804);
nor U23631 (N_23631,N_23157,N_23089);
xor U23632 (N_23632,N_23285,N_23183);
and U23633 (N_23633,N_23181,N_23325);
nor U23634 (N_23634,N_23160,N_22848);
nor U23635 (N_23635,N_22870,N_23107);
and U23636 (N_23636,N_22867,N_23338);
or U23637 (N_23637,N_23170,N_22929);
xnor U23638 (N_23638,N_22999,N_23005);
xor U23639 (N_23639,N_22899,N_22913);
nor U23640 (N_23640,N_23146,N_22823);
and U23641 (N_23641,N_23196,N_23322);
and U23642 (N_23642,N_22912,N_23060);
xnor U23643 (N_23643,N_23347,N_23331);
nor U23644 (N_23644,N_23053,N_23358);
xor U23645 (N_23645,N_23087,N_22890);
nor U23646 (N_23646,N_23100,N_22863);
nand U23647 (N_23647,N_23391,N_22921);
xnor U23648 (N_23648,N_23008,N_22838);
and U23649 (N_23649,N_23291,N_23354);
or U23650 (N_23650,N_23014,N_22802);
and U23651 (N_23651,N_22907,N_23339);
nor U23652 (N_23652,N_23266,N_22885);
and U23653 (N_23653,N_22897,N_23169);
nand U23654 (N_23654,N_22960,N_23281);
and U23655 (N_23655,N_23133,N_23097);
and U23656 (N_23656,N_23073,N_23064);
and U23657 (N_23657,N_22856,N_23289);
nor U23658 (N_23658,N_23307,N_23043);
nand U23659 (N_23659,N_23209,N_23367);
or U23660 (N_23660,N_23304,N_23152);
and U23661 (N_23661,N_22953,N_22884);
nand U23662 (N_23662,N_23287,N_22871);
nand U23663 (N_23663,N_22845,N_23179);
and U23664 (N_23664,N_23159,N_23030);
nand U23665 (N_23665,N_23184,N_23346);
xnor U23666 (N_23666,N_22927,N_23055);
nor U23667 (N_23667,N_23318,N_22909);
xor U23668 (N_23668,N_22954,N_23381);
nand U23669 (N_23669,N_23369,N_22957);
nor U23670 (N_23670,N_23009,N_23263);
or U23671 (N_23671,N_22976,N_22901);
xnor U23672 (N_23672,N_23372,N_23186);
or U23673 (N_23673,N_23117,N_23114);
nand U23674 (N_23674,N_23142,N_22852);
or U23675 (N_23675,N_22873,N_23384);
xor U23676 (N_23676,N_23310,N_22979);
nor U23677 (N_23677,N_22928,N_23334);
xnor U23678 (N_23678,N_23252,N_23059);
xor U23679 (N_23679,N_23171,N_22924);
nor U23680 (N_23680,N_23352,N_23328);
and U23681 (N_23681,N_23245,N_22994);
nand U23682 (N_23682,N_23371,N_23233);
nand U23683 (N_23683,N_23016,N_22846);
nor U23684 (N_23684,N_23156,N_23375);
nor U23685 (N_23685,N_22906,N_23095);
xnor U23686 (N_23686,N_22947,N_22875);
xnor U23687 (N_23687,N_22993,N_23126);
or U23688 (N_23688,N_23216,N_22923);
and U23689 (N_23689,N_23215,N_22948);
and U23690 (N_23690,N_23190,N_22877);
or U23691 (N_23691,N_23103,N_23267);
xor U23692 (N_23692,N_23071,N_23261);
and U23693 (N_23693,N_22967,N_23232);
or U23694 (N_23694,N_23039,N_22937);
and U23695 (N_23695,N_23025,N_22992);
xor U23696 (N_23696,N_23298,N_23147);
xor U23697 (N_23697,N_23251,N_23230);
nor U23698 (N_23698,N_23019,N_23154);
and U23699 (N_23699,N_22818,N_23282);
nand U23700 (N_23700,N_22918,N_22851);
nor U23701 (N_23701,N_23143,N_23382);
or U23702 (N_23702,N_23263,N_23290);
nor U23703 (N_23703,N_22898,N_23245);
nand U23704 (N_23704,N_22909,N_22902);
nand U23705 (N_23705,N_23232,N_23171);
and U23706 (N_23706,N_23031,N_23322);
nor U23707 (N_23707,N_22969,N_23157);
and U23708 (N_23708,N_23222,N_23110);
and U23709 (N_23709,N_22873,N_23052);
xor U23710 (N_23710,N_22977,N_22991);
nand U23711 (N_23711,N_23312,N_22980);
xor U23712 (N_23712,N_22938,N_23310);
nand U23713 (N_23713,N_22829,N_23260);
xor U23714 (N_23714,N_22910,N_23387);
and U23715 (N_23715,N_23304,N_22902);
nand U23716 (N_23716,N_23285,N_23343);
and U23717 (N_23717,N_23083,N_23005);
xnor U23718 (N_23718,N_22958,N_22835);
xnor U23719 (N_23719,N_23183,N_23260);
and U23720 (N_23720,N_23286,N_22802);
and U23721 (N_23721,N_22836,N_23012);
or U23722 (N_23722,N_23182,N_23162);
xnor U23723 (N_23723,N_22906,N_22978);
nand U23724 (N_23724,N_23316,N_23024);
nor U23725 (N_23725,N_23281,N_23293);
nor U23726 (N_23726,N_23266,N_23135);
nand U23727 (N_23727,N_23389,N_22907);
nand U23728 (N_23728,N_22903,N_22865);
or U23729 (N_23729,N_23356,N_23193);
and U23730 (N_23730,N_23373,N_23387);
or U23731 (N_23731,N_23014,N_23017);
xnor U23732 (N_23732,N_23389,N_22974);
nor U23733 (N_23733,N_22838,N_22905);
and U23734 (N_23734,N_22904,N_22903);
xnor U23735 (N_23735,N_22998,N_23127);
and U23736 (N_23736,N_23112,N_22820);
or U23737 (N_23737,N_22984,N_23058);
or U23738 (N_23738,N_23268,N_23156);
or U23739 (N_23739,N_23033,N_23118);
nor U23740 (N_23740,N_23111,N_23159);
xor U23741 (N_23741,N_23034,N_22927);
xnor U23742 (N_23742,N_22851,N_22861);
nand U23743 (N_23743,N_23132,N_23094);
nand U23744 (N_23744,N_22929,N_22989);
or U23745 (N_23745,N_23019,N_23213);
nor U23746 (N_23746,N_23326,N_23310);
nor U23747 (N_23747,N_22950,N_22885);
or U23748 (N_23748,N_22891,N_23235);
nand U23749 (N_23749,N_23052,N_22977);
xor U23750 (N_23750,N_22878,N_23353);
and U23751 (N_23751,N_23000,N_23138);
xnor U23752 (N_23752,N_23214,N_23200);
nor U23753 (N_23753,N_22898,N_22960);
nand U23754 (N_23754,N_23029,N_22821);
and U23755 (N_23755,N_23048,N_22866);
nor U23756 (N_23756,N_22967,N_23183);
xnor U23757 (N_23757,N_23369,N_22937);
or U23758 (N_23758,N_23089,N_23097);
xnor U23759 (N_23759,N_23039,N_23207);
nor U23760 (N_23760,N_22802,N_23087);
and U23761 (N_23761,N_23101,N_23297);
or U23762 (N_23762,N_23352,N_23032);
xnor U23763 (N_23763,N_22916,N_23293);
and U23764 (N_23764,N_22818,N_22871);
xor U23765 (N_23765,N_23375,N_23089);
xor U23766 (N_23766,N_23221,N_23082);
nor U23767 (N_23767,N_23324,N_23373);
or U23768 (N_23768,N_23202,N_22863);
xor U23769 (N_23769,N_22844,N_23306);
xor U23770 (N_23770,N_22805,N_22922);
nand U23771 (N_23771,N_23332,N_23218);
nand U23772 (N_23772,N_23317,N_23000);
xor U23773 (N_23773,N_23175,N_23190);
xnor U23774 (N_23774,N_23039,N_23138);
xnor U23775 (N_23775,N_23131,N_23326);
or U23776 (N_23776,N_23020,N_23357);
nand U23777 (N_23777,N_22888,N_23083);
nor U23778 (N_23778,N_23221,N_23292);
xor U23779 (N_23779,N_23227,N_22975);
or U23780 (N_23780,N_22918,N_23222);
xnor U23781 (N_23781,N_22991,N_22961);
xor U23782 (N_23782,N_23135,N_22909);
or U23783 (N_23783,N_22868,N_22866);
or U23784 (N_23784,N_23379,N_22985);
or U23785 (N_23785,N_23108,N_22956);
or U23786 (N_23786,N_23151,N_23215);
nor U23787 (N_23787,N_22842,N_23103);
and U23788 (N_23788,N_23323,N_22953);
nor U23789 (N_23789,N_23090,N_22931);
or U23790 (N_23790,N_23090,N_23303);
nor U23791 (N_23791,N_22947,N_22982);
and U23792 (N_23792,N_23165,N_23151);
and U23793 (N_23793,N_23282,N_22969);
xor U23794 (N_23794,N_23353,N_22898);
nor U23795 (N_23795,N_23188,N_23276);
nand U23796 (N_23796,N_23216,N_22867);
or U23797 (N_23797,N_22902,N_22824);
and U23798 (N_23798,N_22902,N_23085);
or U23799 (N_23799,N_23204,N_23038);
nand U23800 (N_23800,N_23021,N_23084);
nor U23801 (N_23801,N_23118,N_23240);
nand U23802 (N_23802,N_23143,N_23319);
xor U23803 (N_23803,N_23076,N_23259);
nand U23804 (N_23804,N_23024,N_22951);
nand U23805 (N_23805,N_23229,N_22813);
xnor U23806 (N_23806,N_22946,N_23191);
nor U23807 (N_23807,N_23267,N_23344);
and U23808 (N_23808,N_23009,N_23010);
or U23809 (N_23809,N_22941,N_23371);
xor U23810 (N_23810,N_23203,N_23213);
or U23811 (N_23811,N_22888,N_22875);
and U23812 (N_23812,N_23273,N_23379);
nand U23813 (N_23813,N_23252,N_22825);
nand U23814 (N_23814,N_23098,N_23361);
or U23815 (N_23815,N_23301,N_22933);
or U23816 (N_23816,N_22842,N_23390);
nand U23817 (N_23817,N_22859,N_23004);
or U23818 (N_23818,N_22932,N_22817);
nor U23819 (N_23819,N_23080,N_23186);
and U23820 (N_23820,N_23117,N_23154);
nand U23821 (N_23821,N_22966,N_22819);
nand U23822 (N_23822,N_22942,N_23329);
nor U23823 (N_23823,N_23388,N_22961);
nand U23824 (N_23824,N_23295,N_22950);
xnor U23825 (N_23825,N_23041,N_23350);
and U23826 (N_23826,N_22965,N_23235);
and U23827 (N_23827,N_23177,N_23206);
and U23828 (N_23828,N_23041,N_22804);
nand U23829 (N_23829,N_22942,N_23282);
nand U23830 (N_23830,N_23107,N_23348);
nor U23831 (N_23831,N_23316,N_22888);
nand U23832 (N_23832,N_22880,N_23012);
and U23833 (N_23833,N_22980,N_23168);
and U23834 (N_23834,N_23061,N_23072);
nand U23835 (N_23835,N_23058,N_22958);
or U23836 (N_23836,N_22814,N_22923);
nor U23837 (N_23837,N_23044,N_23220);
xor U23838 (N_23838,N_23169,N_23002);
and U23839 (N_23839,N_23140,N_23291);
or U23840 (N_23840,N_23319,N_23294);
and U23841 (N_23841,N_23070,N_23300);
xor U23842 (N_23842,N_23379,N_23238);
or U23843 (N_23843,N_22975,N_22887);
and U23844 (N_23844,N_23287,N_23317);
xnor U23845 (N_23845,N_22917,N_22914);
nor U23846 (N_23846,N_23057,N_23062);
nor U23847 (N_23847,N_23315,N_22982);
and U23848 (N_23848,N_23297,N_23174);
and U23849 (N_23849,N_23031,N_22823);
nor U23850 (N_23850,N_22813,N_23347);
or U23851 (N_23851,N_22842,N_23066);
nand U23852 (N_23852,N_23263,N_23045);
or U23853 (N_23853,N_23202,N_23030);
or U23854 (N_23854,N_22926,N_22898);
nor U23855 (N_23855,N_23068,N_23016);
nor U23856 (N_23856,N_22836,N_22890);
xnor U23857 (N_23857,N_22916,N_22860);
nand U23858 (N_23858,N_23169,N_22802);
nor U23859 (N_23859,N_22934,N_23129);
xnor U23860 (N_23860,N_23137,N_23399);
nand U23861 (N_23861,N_22933,N_23092);
nor U23862 (N_23862,N_22894,N_23329);
and U23863 (N_23863,N_22879,N_22971);
nand U23864 (N_23864,N_22994,N_23323);
nand U23865 (N_23865,N_23026,N_23288);
nand U23866 (N_23866,N_23228,N_22879);
or U23867 (N_23867,N_22947,N_22820);
nor U23868 (N_23868,N_23242,N_23288);
xor U23869 (N_23869,N_23368,N_22996);
xnor U23870 (N_23870,N_23121,N_23212);
nand U23871 (N_23871,N_23069,N_23213);
nand U23872 (N_23872,N_23050,N_22830);
xor U23873 (N_23873,N_23350,N_22913);
or U23874 (N_23874,N_23372,N_22936);
xor U23875 (N_23875,N_22966,N_23396);
nor U23876 (N_23876,N_22862,N_23360);
nand U23877 (N_23877,N_23086,N_23119);
nand U23878 (N_23878,N_22943,N_23183);
or U23879 (N_23879,N_22852,N_22868);
or U23880 (N_23880,N_22948,N_23265);
nor U23881 (N_23881,N_23321,N_22975);
nand U23882 (N_23882,N_22995,N_23175);
or U23883 (N_23883,N_23321,N_23285);
and U23884 (N_23884,N_23375,N_22937);
nor U23885 (N_23885,N_22954,N_23046);
nor U23886 (N_23886,N_23393,N_23347);
nand U23887 (N_23887,N_23112,N_23367);
xor U23888 (N_23888,N_23221,N_22978);
and U23889 (N_23889,N_22980,N_22803);
xor U23890 (N_23890,N_23132,N_22986);
nor U23891 (N_23891,N_23139,N_23360);
nor U23892 (N_23892,N_23230,N_23339);
nor U23893 (N_23893,N_22915,N_23075);
xor U23894 (N_23894,N_23371,N_22851);
or U23895 (N_23895,N_23314,N_22807);
nand U23896 (N_23896,N_23248,N_23266);
nand U23897 (N_23897,N_23129,N_23240);
or U23898 (N_23898,N_23153,N_22852);
or U23899 (N_23899,N_22952,N_22916);
or U23900 (N_23900,N_23066,N_23396);
nand U23901 (N_23901,N_23120,N_23008);
and U23902 (N_23902,N_23023,N_23135);
nor U23903 (N_23903,N_23295,N_22896);
and U23904 (N_23904,N_23281,N_23149);
and U23905 (N_23905,N_23287,N_23124);
xor U23906 (N_23906,N_23165,N_23087);
nor U23907 (N_23907,N_22875,N_23240);
and U23908 (N_23908,N_23281,N_22872);
nand U23909 (N_23909,N_23202,N_23259);
and U23910 (N_23910,N_23197,N_22828);
nor U23911 (N_23911,N_23216,N_23015);
xnor U23912 (N_23912,N_23095,N_23392);
and U23913 (N_23913,N_23002,N_23292);
and U23914 (N_23914,N_22902,N_22907);
xor U23915 (N_23915,N_23312,N_23288);
or U23916 (N_23916,N_23165,N_23360);
or U23917 (N_23917,N_23365,N_22824);
nand U23918 (N_23918,N_23244,N_23344);
nand U23919 (N_23919,N_23275,N_23004);
or U23920 (N_23920,N_22931,N_22933);
or U23921 (N_23921,N_23392,N_23100);
and U23922 (N_23922,N_22894,N_22991);
nand U23923 (N_23923,N_23108,N_23337);
and U23924 (N_23924,N_23222,N_22928);
nand U23925 (N_23925,N_22906,N_23237);
or U23926 (N_23926,N_22930,N_22884);
and U23927 (N_23927,N_23119,N_23313);
nand U23928 (N_23928,N_23072,N_23017);
or U23929 (N_23929,N_23262,N_23203);
nor U23930 (N_23930,N_22816,N_23030);
nor U23931 (N_23931,N_23130,N_23176);
or U23932 (N_23932,N_23395,N_23192);
nor U23933 (N_23933,N_23270,N_23285);
nand U23934 (N_23934,N_23094,N_23236);
xnor U23935 (N_23935,N_22950,N_23362);
and U23936 (N_23936,N_23104,N_22837);
xnor U23937 (N_23937,N_23034,N_23096);
nor U23938 (N_23938,N_22941,N_23216);
nor U23939 (N_23939,N_23037,N_23374);
and U23940 (N_23940,N_23353,N_23012);
xor U23941 (N_23941,N_23064,N_23135);
nand U23942 (N_23942,N_23076,N_22978);
or U23943 (N_23943,N_22954,N_23277);
or U23944 (N_23944,N_23316,N_22925);
nand U23945 (N_23945,N_23152,N_23079);
xnor U23946 (N_23946,N_23335,N_23203);
and U23947 (N_23947,N_23355,N_23200);
nor U23948 (N_23948,N_23077,N_23130);
nand U23949 (N_23949,N_22899,N_23354);
or U23950 (N_23950,N_23297,N_23226);
and U23951 (N_23951,N_22984,N_23272);
and U23952 (N_23952,N_23088,N_23252);
xor U23953 (N_23953,N_23387,N_22859);
xor U23954 (N_23954,N_23253,N_22876);
and U23955 (N_23955,N_23094,N_23388);
xor U23956 (N_23956,N_23260,N_23042);
nand U23957 (N_23957,N_23189,N_22814);
and U23958 (N_23958,N_22950,N_22869);
nor U23959 (N_23959,N_22950,N_22891);
nand U23960 (N_23960,N_23339,N_23344);
and U23961 (N_23961,N_23019,N_23294);
nor U23962 (N_23962,N_23309,N_22807);
xnor U23963 (N_23963,N_22807,N_23144);
and U23964 (N_23964,N_23008,N_22968);
nand U23965 (N_23965,N_23234,N_23270);
xnor U23966 (N_23966,N_23121,N_23021);
and U23967 (N_23967,N_23029,N_23132);
xnor U23968 (N_23968,N_22813,N_23160);
or U23969 (N_23969,N_22986,N_23196);
xnor U23970 (N_23970,N_23250,N_23171);
nand U23971 (N_23971,N_23069,N_23236);
or U23972 (N_23972,N_23369,N_23184);
xnor U23973 (N_23973,N_22820,N_23064);
and U23974 (N_23974,N_22938,N_22805);
nor U23975 (N_23975,N_23367,N_23062);
xor U23976 (N_23976,N_23207,N_22910);
xor U23977 (N_23977,N_23044,N_23034);
nand U23978 (N_23978,N_22958,N_23330);
nand U23979 (N_23979,N_23130,N_23062);
and U23980 (N_23980,N_23043,N_23119);
or U23981 (N_23981,N_23316,N_22910);
nor U23982 (N_23982,N_23017,N_22896);
xnor U23983 (N_23983,N_23049,N_22961);
nand U23984 (N_23984,N_23330,N_23042);
nor U23985 (N_23985,N_22819,N_23144);
or U23986 (N_23986,N_22820,N_23253);
or U23987 (N_23987,N_23350,N_23204);
and U23988 (N_23988,N_22831,N_23301);
xnor U23989 (N_23989,N_23129,N_23171);
and U23990 (N_23990,N_22936,N_22887);
xnor U23991 (N_23991,N_23396,N_22919);
and U23992 (N_23992,N_23365,N_23311);
and U23993 (N_23993,N_23244,N_23256);
or U23994 (N_23994,N_22905,N_22996);
nand U23995 (N_23995,N_23076,N_22899);
nand U23996 (N_23996,N_22940,N_22828);
and U23997 (N_23997,N_22813,N_22823);
and U23998 (N_23998,N_22854,N_22982);
xnor U23999 (N_23999,N_22949,N_22872);
and U24000 (N_24000,N_23538,N_23441);
and U24001 (N_24001,N_23509,N_23950);
and U24002 (N_24002,N_23819,N_23725);
and U24003 (N_24003,N_23772,N_23626);
and U24004 (N_24004,N_23412,N_23569);
nand U24005 (N_24005,N_23526,N_23546);
and U24006 (N_24006,N_23891,N_23826);
nor U24007 (N_24007,N_23991,N_23755);
or U24008 (N_24008,N_23847,N_23622);
nor U24009 (N_24009,N_23705,N_23972);
or U24010 (N_24010,N_23932,N_23408);
or U24011 (N_24011,N_23924,N_23874);
and U24012 (N_24012,N_23607,N_23999);
xor U24013 (N_24013,N_23736,N_23775);
and U24014 (N_24014,N_23856,N_23915);
nor U24015 (N_24015,N_23816,N_23811);
xor U24016 (N_24016,N_23898,N_23522);
and U24017 (N_24017,N_23824,N_23849);
or U24018 (N_24018,N_23692,N_23964);
and U24019 (N_24019,N_23696,N_23630);
nand U24020 (N_24020,N_23473,N_23794);
nand U24021 (N_24021,N_23894,N_23873);
xnor U24022 (N_24022,N_23529,N_23415);
or U24023 (N_24023,N_23957,N_23475);
or U24024 (N_24024,N_23591,N_23628);
and U24025 (N_24025,N_23491,N_23449);
or U24026 (N_24026,N_23733,N_23767);
xnor U24027 (N_24027,N_23930,N_23836);
nand U24028 (N_24028,N_23629,N_23676);
nand U24029 (N_24029,N_23618,N_23784);
nand U24030 (N_24030,N_23872,N_23625);
or U24031 (N_24031,N_23425,N_23603);
nand U24032 (N_24032,N_23890,N_23610);
xor U24033 (N_24033,N_23837,N_23627);
nand U24034 (N_24034,N_23430,N_23765);
nand U24035 (N_24035,N_23520,N_23481);
nor U24036 (N_24036,N_23620,N_23853);
xnor U24037 (N_24037,N_23446,N_23785);
nand U24038 (N_24038,N_23869,N_23909);
nand U24039 (N_24039,N_23472,N_23967);
nand U24040 (N_24040,N_23442,N_23694);
nor U24041 (N_24041,N_23619,N_23443);
and U24042 (N_24042,N_23731,N_23668);
xor U24043 (N_24043,N_23411,N_23745);
and U24044 (N_24044,N_23969,N_23877);
and U24045 (N_24045,N_23571,N_23848);
nor U24046 (N_24046,N_23584,N_23482);
xor U24047 (N_24047,N_23783,N_23455);
xnor U24048 (N_24048,N_23746,N_23899);
nor U24049 (N_24049,N_23786,N_23928);
nand U24050 (N_24050,N_23406,N_23465);
xor U24051 (N_24051,N_23519,N_23421);
and U24052 (N_24052,N_23748,N_23822);
nand U24053 (N_24053,N_23807,N_23750);
or U24054 (N_24054,N_23914,N_23801);
and U24055 (N_24055,N_23921,N_23881);
xor U24056 (N_24056,N_23402,N_23580);
xnor U24057 (N_24057,N_23466,N_23712);
nor U24058 (N_24058,N_23492,N_23693);
nand U24059 (N_24059,N_23825,N_23617);
xor U24060 (N_24060,N_23865,N_23568);
nor U24061 (N_24061,N_23863,N_23660);
nor U24062 (N_24062,N_23714,N_23722);
nor U24063 (N_24063,N_23771,N_23742);
nor U24064 (N_24064,N_23700,N_23933);
nor U24065 (N_24065,N_23685,N_23457);
xnor U24066 (N_24066,N_23684,N_23959);
nand U24067 (N_24067,N_23669,N_23403);
and U24068 (N_24068,N_23615,N_23806);
and U24069 (N_24069,N_23754,N_23947);
xnor U24070 (N_24070,N_23536,N_23943);
or U24071 (N_24071,N_23946,N_23850);
nand U24072 (N_24072,N_23737,N_23562);
or U24073 (N_24073,N_23878,N_23587);
nor U24074 (N_24074,N_23920,N_23506);
nor U24075 (N_24075,N_23908,N_23780);
nor U24076 (N_24076,N_23897,N_23458);
or U24077 (N_24077,N_23813,N_23554);
nand U24078 (N_24078,N_23505,N_23977);
nor U24079 (N_24079,N_23489,N_23936);
nor U24080 (N_24080,N_23595,N_23799);
nor U24081 (N_24081,N_23711,N_23675);
and U24082 (N_24082,N_23414,N_23471);
or U24083 (N_24083,N_23662,N_23533);
and U24084 (N_24084,N_23564,N_23624);
xor U24085 (N_24085,N_23931,N_23576);
and U24086 (N_24086,N_23949,N_23980);
and U24087 (N_24087,N_23439,N_23462);
xnor U24088 (N_24088,N_23616,N_23996);
nor U24089 (N_24089,N_23800,N_23792);
nor U24090 (N_24090,N_23905,N_23706);
or U24091 (N_24091,N_23703,N_23641);
nor U24092 (N_24092,N_23487,N_23718);
xor U24093 (N_24093,N_23695,N_23507);
or U24094 (N_24094,N_23958,N_23868);
nand U24095 (N_24095,N_23761,N_23757);
nor U24096 (N_24096,N_23532,N_23893);
xnor U24097 (N_24097,N_23404,N_23829);
or U24098 (N_24098,N_23774,N_23919);
nand U24099 (N_24099,N_23479,N_23553);
or U24100 (N_24100,N_23555,N_23859);
or U24101 (N_24101,N_23987,N_23524);
nand U24102 (N_24102,N_23420,N_23447);
nor U24103 (N_24103,N_23955,N_23778);
nor U24104 (N_24104,N_23787,N_23812);
and U24105 (N_24105,N_23835,N_23779);
or U24106 (N_24106,N_23497,N_23839);
nor U24107 (N_24107,N_23469,N_23486);
or U24108 (N_24108,N_23478,N_23585);
or U24109 (N_24109,N_23503,N_23752);
nor U24110 (N_24110,N_23770,N_23876);
nor U24111 (N_24111,N_23727,N_23940);
nand U24112 (N_24112,N_23852,N_23510);
nand U24113 (N_24113,N_23884,N_23612);
and U24114 (N_24114,N_23918,N_23713);
nor U24115 (N_24115,N_23961,N_23611);
nand U24116 (N_24116,N_23781,N_23913);
and U24117 (N_24117,N_23652,N_23866);
nor U24118 (N_24118,N_23638,N_23658);
nor U24119 (N_24119,N_23593,N_23719);
xnor U24120 (N_24120,N_23756,N_23892);
and U24121 (N_24121,N_23704,N_23753);
nor U24122 (N_24122,N_23547,N_23710);
nand U24123 (N_24123,N_23508,N_23802);
nor U24124 (N_24124,N_23600,N_23896);
xnor U24125 (N_24125,N_23689,N_23614);
xnor U24126 (N_24126,N_23838,N_23743);
xor U24127 (N_24127,N_23724,N_23515);
and U24128 (N_24128,N_23682,N_23966);
and U24129 (N_24129,N_23567,N_23906);
and U24130 (N_24130,N_23574,N_23424);
xnor U24131 (N_24131,N_23855,N_23831);
nor U24132 (N_24132,N_23860,N_23644);
and U24133 (N_24133,N_23605,N_23598);
nor U24134 (N_24134,N_23531,N_23577);
and U24135 (N_24135,N_23688,N_23938);
xnor U24136 (N_24136,N_23416,N_23606);
nand U24137 (N_24137,N_23960,N_23922);
nor U24138 (N_24138,N_23432,N_23895);
nor U24139 (N_24139,N_23460,N_23461);
xnor U24140 (N_24140,N_23766,N_23609);
or U24141 (N_24141,N_23400,N_23521);
nor U24142 (N_24142,N_23976,N_23740);
and U24143 (N_24143,N_23631,N_23534);
xnor U24144 (N_24144,N_23832,N_23545);
or U24145 (N_24145,N_23602,N_23764);
or U24146 (N_24146,N_23582,N_23604);
xor U24147 (N_24147,N_23565,N_23566);
or U24148 (N_24148,N_23975,N_23667);
nand U24149 (N_24149,N_23648,N_23516);
and U24150 (N_24150,N_23483,N_23539);
nor U24151 (N_24151,N_23923,N_23708);
or U24152 (N_24152,N_23671,N_23841);
and U24153 (N_24153,N_23594,N_23809);
nand U24154 (N_24154,N_23759,N_23716);
and U24155 (N_24155,N_23499,N_23805);
or U24156 (N_24156,N_23744,N_23962);
nor U24157 (N_24157,N_23552,N_23985);
nor U24158 (N_24158,N_23470,N_23444);
or U24159 (N_24159,N_23570,N_23879);
nor U24160 (N_24160,N_23581,N_23840);
nor U24161 (N_24161,N_23844,N_23769);
or U24162 (N_24162,N_23608,N_23513);
and U24163 (N_24163,N_23548,N_23715);
and U24164 (N_24164,N_23464,N_23561);
nor U24165 (N_24165,N_23965,N_23454);
xor U24166 (N_24166,N_23834,N_23563);
nand U24167 (N_24167,N_23749,N_23514);
xnor U24168 (N_24168,N_23815,N_23670);
xor U24169 (N_24169,N_23490,N_23912);
and U24170 (N_24170,N_23687,N_23496);
or U24171 (N_24171,N_23929,N_23954);
or U24172 (N_24172,N_23867,N_23798);
xnor U24173 (N_24173,N_23992,N_23973);
nand U24174 (N_24174,N_23735,N_23937);
xnor U24175 (N_24175,N_23953,N_23663);
and U24176 (N_24176,N_23951,N_23431);
or U24177 (N_24177,N_23640,N_23636);
nand U24178 (N_24178,N_23418,N_23945);
or U24179 (N_24179,N_23575,N_23527);
nor U24180 (N_24180,N_23817,N_23583);
nor U24181 (N_24181,N_23741,N_23528);
and U24182 (N_24182,N_23407,N_23782);
xnor U24183 (N_24183,N_23907,N_23998);
xnor U24184 (N_24184,N_23948,N_23665);
and U24185 (N_24185,N_23440,N_23790);
xor U24186 (N_24186,N_23886,N_23474);
or U24187 (N_24187,N_23875,N_23550);
and U24188 (N_24188,N_23702,N_23437);
and U24189 (N_24189,N_23511,N_23572);
or U24190 (N_24190,N_23677,N_23535);
xnor U24191 (N_24191,N_23730,N_23788);
nand U24192 (N_24192,N_23558,N_23468);
and U24193 (N_24193,N_23666,N_23726);
or U24194 (N_24194,N_23984,N_23690);
xnor U24195 (N_24195,N_23747,N_23986);
and U24196 (N_24196,N_23678,N_23401);
nor U24197 (N_24197,N_23463,N_23941);
nor U24198 (N_24198,N_23871,N_23653);
nor U24199 (N_24199,N_23453,N_23997);
xnor U24200 (N_24200,N_23927,N_23827);
and U24201 (N_24201,N_23588,N_23413);
xor U24202 (N_24202,N_23760,N_23803);
or U24203 (N_24203,N_23823,N_23632);
nor U24204 (N_24204,N_23709,N_23902);
or U24205 (N_24205,N_23974,N_23501);
nor U24206 (N_24206,N_23493,N_23592);
nor U24207 (N_24207,N_23544,N_23728);
nor U24208 (N_24208,N_23707,N_23883);
xor U24209 (N_24209,N_23979,N_23720);
xnor U24210 (N_24210,N_23995,N_23858);
and U24211 (N_24211,N_23732,N_23729);
and U24212 (N_24212,N_23990,N_23993);
or U24213 (N_24213,N_23651,N_23542);
nor U24214 (N_24214,N_23983,N_23523);
xor U24215 (N_24215,N_23763,N_23797);
nor U24216 (N_24216,N_23517,N_23559);
nand U24217 (N_24217,N_23525,N_23916);
xor U24218 (N_24218,N_23818,N_23723);
or U24219 (N_24219,N_23655,N_23643);
xor U24220 (N_24220,N_23541,N_23939);
and U24221 (N_24221,N_23795,N_23427);
nand U24222 (N_24222,N_23910,N_23861);
xnor U24223 (N_24223,N_23656,N_23904);
and U24224 (N_24224,N_23549,N_23699);
nand U24225 (N_24225,N_23500,N_23701);
nand U24226 (N_24226,N_23808,N_23498);
nand U24227 (N_24227,N_23804,N_23925);
xnor U24228 (N_24228,N_23661,N_23433);
or U24229 (N_24229,N_23777,N_23672);
xor U24230 (N_24230,N_23485,N_23504);
and U24231 (N_24231,N_23683,N_23762);
and U24232 (N_24232,N_23935,N_23845);
or U24233 (N_24233,N_23480,N_23968);
or U24234 (N_24234,N_23579,N_23880);
and U24235 (N_24235,N_23679,N_23642);
and U24236 (N_24236,N_23476,N_23851);
nor U24237 (N_24237,N_23599,N_23673);
nand U24238 (N_24238,N_23842,N_23882);
and U24239 (N_24239,N_23970,N_23978);
nand U24240 (N_24240,N_23654,N_23657);
nand U24241 (N_24241,N_23551,N_23900);
or U24242 (N_24242,N_23451,N_23560);
xor U24243 (N_24243,N_23426,N_23681);
nand U24244 (N_24244,N_23452,N_23870);
nand U24245 (N_24245,N_23601,N_23739);
nor U24246 (N_24246,N_23751,N_23589);
xor U24247 (N_24247,N_23495,N_23814);
xnor U24248 (N_24248,N_23846,N_23647);
or U24249 (N_24249,N_23512,N_23646);
and U24250 (N_24250,N_23857,N_23926);
xor U24251 (N_24251,N_23956,N_23410);
nor U24252 (N_24252,N_23537,N_23911);
and U24253 (N_24253,N_23793,N_23674);
and U24254 (N_24254,N_23810,N_23428);
nor U24255 (N_24255,N_23650,N_23423);
and U24256 (N_24256,N_23738,N_23789);
xnor U24257 (N_24257,N_23456,N_23821);
nand U24258 (N_24258,N_23944,N_23623);
and U24259 (N_24259,N_23734,N_23540);
nor U24260 (N_24260,N_23830,N_23971);
or U24261 (N_24261,N_23409,N_23989);
or U24262 (N_24262,N_23637,N_23435);
nand U24263 (N_24263,N_23721,N_23691);
and U24264 (N_24264,N_23438,N_23635);
nor U24265 (N_24265,N_23448,N_23952);
xnor U24266 (N_24266,N_23864,N_23459);
and U24267 (N_24267,N_23988,N_23776);
nand U24268 (N_24268,N_23982,N_23934);
and U24269 (N_24269,N_23697,N_23596);
xnor U24270 (N_24270,N_23590,N_23917);
and U24271 (N_24271,N_23994,N_23791);
and U24272 (N_24272,N_23901,N_23820);
nor U24273 (N_24273,N_23477,N_23634);
and U24274 (N_24274,N_23717,N_23686);
and U24275 (N_24275,N_23494,N_23885);
and U24276 (N_24276,N_23405,N_23664);
nand U24277 (N_24277,N_23862,N_23543);
nand U24278 (N_24278,N_23586,N_23981);
nand U24279 (N_24279,N_23578,N_23484);
nor U24280 (N_24280,N_23613,N_23573);
nand U24281 (N_24281,N_23419,N_23621);
and U24282 (N_24282,N_23502,N_23758);
or U24283 (N_24283,N_23773,N_23942);
xnor U24284 (N_24284,N_23796,N_23597);
xnor U24285 (N_24285,N_23649,N_23445);
xnor U24286 (N_24286,N_23888,N_23556);
nor U24287 (N_24287,N_23833,N_23467);
or U24288 (N_24288,N_23422,N_23903);
nor U24289 (N_24289,N_23530,N_23639);
and U24290 (N_24290,N_23828,N_23633);
xor U24291 (N_24291,N_23659,N_23450);
or U24292 (N_24292,N_23417,N_23645);
or U24293 (N_24293,N_23843,N_23429);
or U24294 (N_24294,N_23963,N_23434);
or U24295 (N_24295,N_23436,N_23557);
xnor U24296 (N_24296,N_23518,N_23698);
and U24297 (N_24297,N_23680,N_23854);
nor U24298 (N_24298,N_23889,N_23887);
xnor U24299 (N_24299,N_23488,N_23768);
xnor U24300 (N_24300,N_23804,N_23789);
nand U24301 (N_24301,N_23489,N_23971);
and U24302 (N_24302,N_23434,N_23820);
nand U24303 (N_24303,N_23885,N_23608);
xor U24304 (N_24304,N_23601,N_23786);
xor U24305 (N_24305,N_23718,N_23565);
or U24306 (N_24306,N_23704,N_23974);
xor U24307 (N_24307,N_23536,N_23620);
xor U24308 (N_24308,N_23479,N_23513);
or U24309 (N_24309,N_23570,N_23744);
xor U24310 (N_24310,N_23570,N_23855);
nand U24311 (N_24311,N_23460,N_23645);
xnor U24312 (N_24312,N_23611,N_23719);
and U24313 (N_24313,N_23716,N_23532);
or U24314 (N_24314,N_23680,N_23523);
xnor U24315 (N_24315,N_23414,N_23599);
and U24316 (N_24316,N_23939,N_23512);
and U24317 (N_24317,N_23735,N_23899);
nand U24318 (N_24318,N_23791,N_23663);
xnor U24319 (N_24319,N_23996,N_23754);
and U24320 (N_24320,N_23968,N_23880);
and U24321 (N_24321,N_23631,N_23593);
and U24322 (N_24322,N_23714,N_23465);
nor U24323 (N_24323,N_23614,N_23908);
or U24324 (N_24324,N_23873,N_23671);
xor U24325 (N_24325,N_23643,N_23709);
and U24326 (N_24326,N_23771,N_23975);
nor U24327 (N_24327,N_23509,N_23758);
or U24328 (N_24328,N_23401,N_23717);
and U24329 (N_24329,N_23483,N_23749);
nand U24330 (N_24330,N_23666,N_23988);
xor U24331 (N_24331,N_23922,N_23565);
and U24332 (N_24332,N_23415,N_23723);
nor U24333 (N_24333,N_23635,N_23835);
xnor U24334 (N_24334,N_23858,N_23480);
xnor U24335 (N_24335,N_23784,N_23541);
and U24336 (N_24336,N_23814,N_23662);
nand U24337 (N_24337,N_23586,N_23917);
or U24338 (N_24338,N_23913,N_23547);
or U24339 (N_24339,N_23650,N_23572);
nand U24340 (N_24340,N_23864,N_23844);
and U24341 (N_24341,N_23948,N_23520);
xor U24342 (N_24342,N_23511,N_23752);
nor U24343 (N_24343,N_23773,N_23416);
nor U24344 (N_24344,N_23727,N_23598);
xnor U24345 (N_24345,N_23753,N_23927);
nand U24346 (N_24346,N_23648,N_23922);
nor U24347 (N_24347,N_23425,N_23611);
xnor U24348 (N_24348,N_23761,N_23494);
and U24349 (N_24349,N_23499,N_23965);
xor U24350 (N_24350,N_23746,N_23566);
and U24351 (N_24351,N_23982,N_23955);
nand U24352 (N_24352,N_23953,N_23523);
and U24353 (N_24353,N_23933,N_23874);
and U24354 (N_24354,N_23823,N_23752);
nor U24355 (N_24355,N_23849,N_23835);
and U24356 (N_24356,N_23865,N_23683);
xor U24357 (N_24357,N_23607,N_23652);
xor U24358 (N_24358,N_23705,N_23600);
nand U24359 (N_24359,N_23701,N_23851);
nand U24360 (N_24360,N_23913,N_23650);
xnor U24361 (N_24361,N_23407,N_23966);
or U24362 (N_24362,N_23925,N_23813);
nand U24363 (N_24363,N_23554,N_23564);
nand U24364 (N_24364,N_23953,N_23529);
or U24365 (N_24365,N_23861,N_23841);
nand U24366 (N_24366,N_23902,N_23521);
nor U24367 (N_24367,N_23555,N_23561);
nand U24368 (N_24368,N_23700,N_23781);
nor U24369 (N_24369,N_23620,N_23616);
xor U24370 (N_24370,N_23914,N_23789);
nand U24371 (N_24371,N_23923,N_23487);
nor U24372 (N_24372,N_23826,N_23854);
nor U24373 (N_24373,N_23527,N_23413);
and U24374 (N_24374,N_23422,N_23827);
and U24375 (N_24375,N_23827,N_23610);
and U24376 (N_24376,N_23758,N_23775);
or U24377 (N_24377,N_23890,N_23721);
xor U24378 (N_24378,N_23841,N_23594);
nand U24379 (N_24379,N_23972,N_23658);
nor U24380 (N_24380,N_23701,N_23867);
nand U24381 (N_24381,N_23697,N_23956);
or U24382 (N_24382,N_23769,N_23735);
nor U24383 (N_24383,N_23558,N_23499);
nand U24384 (N_24384,N_23860,N_23588);
xnor U24385 (N_24385,N_23402,N_23649);
nor U24386 (N_24386,N_23624,N_23915);
or U24387 (N_24387,N_23939,N_23436);
nor U24388 (N_24388,N_23842,N_23916);
xnor U24389 (N_24389,N_23652,N_23515);
nor U24390 (N_24390,N_23741,N_23467);
nor U24391 (N_24391,N_23798,N_23727);
and U24392 (N_24392,N_23681,N_23569);
xnor U24393 (N_24393,N_23584,N_23921);
or U24394 (N_24394,N_23526,N_23817);
nor U24395 (N_24395,N_23435,N_23495);
or U24396 (N_24396,N_23643,N_23637);
and U24397 (N_24397,N_23402,N_23557);
xnor U24398 (N_24398,N_23414,N_23424);
nor U24399 (N_24399,N_23867,N_23452);
or U24400 (N_24400,N_23779,N_23857);
xor U24401 (N_24401,N_23759,N_23526);
or U24402 (N_24402,N_23999,N_23931);
nor U24403 (N_24403,N_23717,N_23492);
xor U24404 (N_24404,N_23587,N_23988);
nor U24405 (N_24405,N_23947,N_23690);
nand U24406 (N_24406,N_23746,N_23858);
or U24407 (N_24407,N_23898,N_23435);
xnor U24408 (N_24408,N_23674,N_23513);
and U24409 (N_24409,N_23512,N_23830);
nand U24410 (N_24410,N_23993,N_23744);
or U24411 (N_24411,N_23951,N_23502);
and U24412 (N_24412,N_23658,N_23957);
nand U24413 (N_24413,N_23736,N_23642);
and U24414 (N_24414,N_23505,N_23871);
xnor U24415 (N_24415,N_23979,N_23718);
nand U24416 (N_24416,N_23818,N_23473);
nor U24417 (N_24417,N_23710,N_23410);
nor U24418 (N_24418,N_23939,N_23460);
xor U24419 (N_24419,N_23681,N_23977);
or U24420 (N_24420,N_23843,N_23554);
or U24421 (N_24421,N_23898,N_23948);
nor U24422 (N_24422,N_23891,N_23511);
nand U24423 (N_24423,N_23548,N_23681);
and U24424 (N_24424,N_23902,N_23772);
nand U24425 (N_24425,N_23811,N_23940);
xor U24426 (N_24426,N_23890,N_23718);
xor U24427 (N_24427,N_23754,N_23495);
nor U24428 (N_24428,N_23706,N_23988);
nand U24429 (N_24429,N_23747,N_23578);
xnor U24430 (N_24430,N_23420,N_23482);
nor U24431 (N_24431,N_23725,N_23446);
and U24432 (N_24432,N_23407,N_23759);
xnor U24433 (N_24433,N_23570,N_23918);
nor U24434 (N_24434,N_23487,N_23736);
nor U24435 (N_24435,N_23545,N_23814);
or U24436 (N_24436,N_23453,N_23983);
nand U24437 (N_24437,N_23860,N_23501);
xnor U24438 (N_24438,N_23876,N_23912);
nor U24439 (N_24439,N_23444,N_23703);
nor U24440 (N_24440,N_23582,N_23430);
nand U24441 (N_24441,N_23540,N_23417);
and U24442 (N_24442,N_23993,N_23816);
nand U24443 (N_24443,N_23735,N_23815);
xnor U24444 (N_24444,N_23988,N_23450);
xnor U24445 (N_24445,N_23521,N_23774);
and U24446 (N_24446,N_23902,N_23849);
nor U24447 (N_24447,N_23687,N_23408);
or U24448 (N_24448,N_23800,N_23818);
and U24449 (N_24449,N_23692,N_23630);
nor U24450 (N_24450,N_23952,N_23553);
nand U24451 (N_24451,N_23564,N_23995);
xnor U24452 (N_24452,N_23988,N_23546);
nor U24453 (N_24453,N_23492,N_23818);
nor U24454 (N_24454,N_23879,N_23851);
and U24455 (N_24455,N_23965,N_23676);
xnor U24456 (N_24456,N_23679,N_23899);
and U24457 (N_24457,N_23705,N_23527);
or U24458 (N_24458,N_23739,N_23869);
nor U24459 (N_24459,N_23966,N_23951);
nor U24460 (N_24460,N_23913,N_23767);
or U24461 (N_24461,N_23868,N_23411);
nor U24462 (N_24462,N_23504,N_23845);
and U24463 (N_24463,N_23798,N_23440);
or U24464 (N_24464,N_23822,N_23896);
or U24465 (N_24465,N_23557,N_23554);
nor U24466 (N_24466,N_23466,N_23510);
and U24467 (N_24467,N_23898,N_23803);
and U24468 (N_24468,N_23934,N_23559);
or U24469 (N_24469,N_23580,N_23891);
xor U24470 (N_24470,N_23791,N_23866);
nor U24471 (N_24471,N_23617,N_23482);
and U24472 (N_24472,N_23750,N_23529);
xnor U24473 (N_24473,N_23704,N_23637);
xnor U24474 (N_24474,N_23882,N_23706);
nand U24475 (N_24475,N_23917,N_23536);
nor U24476 (N_24476,N_23675,N_23505);
nand U24477 (N_24477,N_23943,N_23459);
nand U24478 (N_24478,N_23614,N_23968);
xnor U24479 (N_24479,N_23477,N_23774);
nand U24480 (N_24480,N_23862,N_23539);
nor U24481 (N_24481,N_23459,N_23575);
nor U24482 (N_24482,N_23773,N_23619);
xor U24483 (N_24483,N_23538,N_23792);
xnor U24484 (N_24484,N_23824,N_23791);
nand U24485 (N_24485,N_23722,N_23540);
xor U24486 (N_24486,N_23710,N_23809);
xor U24487 (N_24487,N_23491,N_23770);
and U24488 (N_24488,N_23594,N_23567);
xnor U24489 (N_24489,N_23531,N_23415);
and U24490 (N_24490,N_23516,N_23418);
xnor U24491 (N_24491,N_23968,N_23414);
nand U24492 (N_24492,N_23868,N_23567);
nand U24493 (N_24493,N_23648,N_23585);
nor U24494 (N_24494,N_23465,N_23835);
or U24495 (N_24495,N_23965,N_23715);
nand U24496 (N_24496,N_23466,N_23814);
or U24497 (N_24497,N_23999,N_23520);
xor U24498 (N_24498,N_23868,N_23786);
or U24499 (N_24499,N_23631,N_23967);
or U24500 (N_24500,N_23776,N_23556);
or U24501 (N_24501,N_23571,N_23920);
nand U24502 (N_24502,N_23643,N_23958);
xor U24503 (N_24503,N_23417,N_23745);
xor U24504 (N_24504,N_23824,N_23583);
and U24505 (N_24505,N_23557,N_23437);
and U24506 (N_24506,N_23702,N_23844);
xor U24507 (N_24507,N_23878,N_23733);
xnor U24508 (N_24508,N_23706,N_23992);
or U24509 (N_24509,N_23767,N_23625);
or U24510 (N_24510,N_23627,N_23684);
xor U24511 (N_24511,N_23650,N_23765);
and U24512 (N_24512,N_23963,N_23427);
and U24513 (N_24513,N_23410,N_23583);
and U24514 (N_24514,N_23646,N_23963);
nor U24515 (N_24515,N_23781,N_23588);
and U24516 (N_24516,N_23895,N_23731);
and U24517 (N_24517,N_23899,N_23776);
or U24518 (N_24518,N_23930,N_23558);
or U24519 (N_24519,N_23779,N_23828);
or U24520 (N_24520,N_23945,N_23420);
or U24521 (N_24521,N_23723,N_23945);
or U24522 (N_24522,N_23453,N_23523);
xor U24523 (N_24523,N_23724,N_23877);
nand U24524 (N_24524,N_23593,N_23886);
and U24525 (N_24525,N_23638,N_23405);
or U24526 (N_24526,N_23452,N_23895);
nor U24527 (N_24527,N_23460,N_23635);
nor U24528 (N_24528,N_23702,N_23695);
and U24529 (N_24529,N_23724,N_23748);
xnor U24530 (N_24530,N_23858,N_23930);
nor U24531 (N_24531,N_23735,N_23791);
or U24532 (N_24532,N_23641,N_23489);
xor U24533 (N_24533,N_23596,N_23615);
nor U24534 (N_24534,N_23768,N_23755);
xor U24535 (N_24535,N_23747,N_23992);
or U24536 (N_24536,N_23794,N_23409);
nor U24537 (N_24537,N_23760,N_23707);
nand U24538 (N_24538,N_23607,N_23810);
and U24539 (N_24539,N_23735,N_23629);
and U24540 (N_24540,N_23550,N_23863);
xnor U24541 (N_24541,N_23479,N_23840);
nand U24542 (N_24542,N_23588,N_23505);
and U24543 (N_24543,N_23637,N_23512);
xnor U24544 (N_24544,N_23546,N_23560);
nand U24545 (N_24545,N_23773,N_23857);
xor U24546 (N_24546,N_23888,N_23568);
xnor U24547 (N_24547,N_23820,N_23421);
nand U24548 (N_24548,N_23406,N_23496);
nand U24549 (N_24549,N_23996,N_23740);
xor U24550 (N_24550,N_23792,N_23455);
xor U24551 (N_24551,N_23792,N_23760);
nand U24552 (N_24552,N_23676,N_23711);
or U24553 (N_24553,N_23915,N_23945);
or U24554 (N_24554,N_23998,N_23933);
and U24555 (N_24555,N_23974,N_23710);
nor U24556 (N_24556,N_23751,N_23983);
or U24557 (N_24557,N_23623,N_23573);
nand U24558 (N_24558,N_23603,N_23939);
nand U24559 (N_24559,N_23679,N_23437);
and U24560 (N_24560,N_23791,N_23882);
nor U24561 (N_24561,N_23493,N_23917);
and U24562 (N_24562,N_23602,N_23960);
xor U24563 (N_24563,N_23483,N_23422);
nand U24564 (N_24564,N_23430,N_23827);
or U24565 (N_24565,N_23815,N_23865);
nand U24566 (N_24566,N_23402,N_23774);
and U24567 (N_24567,N_23470,N_23747);
xnor U24568 (N_24568,N_23445,N_23730);
or U24569 (N_24569,N_23572,N_23707);
nor U24570 (N_24570,N_23833,N_23989);
or U24571 (N_24571,N_23793,N_23707);
and U24572 (N_24572,N_23610,N_23648);
nor U24573 (N_24573,N_23976,N_23426);
xor U24574 (N_24574,N_23531,N_23651);
nand U24575 (N_24575,N_23893,N_23861);
xor U24576 (N_24576,N_23796,N_23945);
nor U24577 (N_24577,N_23594,N_23775);
nand U24578 (N_24578,N_23730,N_23987);
or U24579 (N_24579,N_23577,N_23501);
and U24580 (N_24580,N_23915,N_23491);
nand U24581 (N_24581,N_23428,N_23668);
or U24582 (N_24582,N_23718,N_23421);
nor U24583 (N_24583,N_23403,N_23952);
or U24584 (N_24584,N_23794,N_23470);
xor U24585 (N_24585,N_23745,N_23898);
or U24586 (N_24586,N_23880,N_23697);
xor U24587 (N_24587,N_23611,N_23519);
and U24588 (N_24588,N_23700,N_23636);
xnor U24589 (N_24589,N_23656,N_23931);
or U24590 (N_24590,N_23421,N_23433);
and U24591 (N_24591,N_23686,N_23723);
or U24592 (N_24592,N_23953,N_23719);
or U24593 (N_24593,N_23673,N_23465);
and U24594 (N_24594,N_23807,N_23646);
nor U24595 (N_24595,N_23471,N_23826);
nor U24596 (N_24596,N_23675,N_23848);
xnor U24597 (N_24597,N_23471,N_23828);
nand U24598 (N_24598,N_23897,N_23702);
nand U24599 (N_24599,N_23584,N_23626);
nand U24600 (N_24600,N_24049,N_24042);
nand U24601 (N_24601,N_24181,N_24356);
nor U24602 (N_24602,N_24502,N_24322);
xnor U24603 (N_24603,N_24384,N_24589);
nor U24604 (N_24604,N_24586,N_24430);
and U24605 (N_24605,N_24422,N_24063);
nor U24606 (N_24606,N_24341,N_24228);
and U24607 (N_24607,N_24131,N_24568);
and U24608 (N_24608,N_24510,N_24167);
nand U24609 (N_24609,N_24015,N_24230);
nor U24610 (N_24610,N_24386,N_24345);
or U24611 (N_24611,N_24296,N_24151);
or U24612 (N_24612,N_24118,N_24154);
and U24613 (N_24613,N_24056,N_24252);
xor U24614 (N_24614,N_24213,N_24378);
nor U24615 (N_24615,N_24104,N_24125);
or U24616 (N_24616,N_24145,N_24244);
or U24617 (N_24617,N_24306,N_24451);
xor U24618 (N_24618,N_24459,N_24518);
or U24619 (N_24619,N_24307,N_24256);
xor U24620 (N_24620,N_24381,N_24025);
nand U24621 (N_24621,N_24082,N_24168);
xor U24622 (N_24622,N_24446,N_24544);
xnor U24623 (N_24623,N_24418,N_24203);
or U24624 (N_24624,N_24376,N_24475);
or U24625 (N_24625,N_24423,N_24062);
and U24626 (N_24626,N_24262,N_24204);
nand U24627 (N_24627,N_24408,N_24585);
and U24628 (N_24628,N_24476,N_24570);
nor U24629 (N_24629,N_24165,N_24157);
nand U24630 (N_24630,N_24404,N_24300);
or U24631 (N_24631,N_24482,N_24431);
or U24632 (N_24632,N_24147,N_24597);
xnor U24633 (N_24633,N_24057,N_24517);
xnor U24634 (N_24634,N_24286,N_24089);
nand U24635 (N_24635,N_24508,N_24578);
or U24636 (N_24636,N_24511,N_24486);
xor U24637 (N_24637,N_24311,N_24263);
and U24638 (N_24638,N_24011,N_24447);
xor U24639 (N_24639,N_24008,N_24474);
xnor U24640 (N_24640,N_24559,N_24044);
nor U24641 (N_24641,N_24093,N_24555);
xnor U24642 (N_24642,N_24548,N_24318);
nor U24643 (N_24643,N_24182,N_24357);
and U24644 (N_24644,N_24484,N_24584);
or U24645 (N_24645,N_24205,N_24143);
nor U24646 (N_24646,N_24196,N_24366);
nand U24647 (N_24647,N_24481,N_24138);
and U24648 (N_24648,N_24110,N_24516);
nor U24649 (N_24649,N_24074,N_24297);
and U24650 (N_24650,N_24149,N_24190);
xnor U24651 (N_24651,N_24577,N_24206);
nand U24652 (N_24652,N_24173,N_24081);
xnor U24653 (N_24653,N_24347,N_24348);
nor U24654 (N_24654,N_24417,N_24462);
xor U24655 (N_24655,N_24009,N_24227);
nor U24656 (N_24656,N_24551,N_24420);
nor U24657 (N_24657,N_24222,N_24461);
xor U24658 (N_24658,N_24403,N_24097);
or U24659 (N_24659,N_24241,N_24253);
nand U24660 (N_24660,N_24188,N_24092);
and U24661 (N_24661,N_24028,N_24268);
xor U24662 (N_24662,N_24444,N_24237);
and U24663 (N_24663,N_24083,N_24365);
xor U24664 (N_24664,N_24591,N_24288);
xnor U24665 (N_24665,N_24330,N_24274);
and U24666 (N_24666,N_24471,N_24080);
and U24667 (N_24667,N_24593,N_24562);
or U24668 (N_24668,N_24304,N_24533);
and U24669 (N_24669,N_24560,N_24160);
nor U24670 (N_24670,N_24034,N_24052);
or U24671 (N_24671,N_24248,N_24477);
or U24672 (N_24672,N_24424,N_24442);
xnor U24673 (N_24673,N_24309,N_24497);
nor U24674 (N_24674,N_24116,N_24023);
nand U24675 (N_24675,N_24117,N_24195);
xnor U24676 (N_24676,N_24111,N_24538);
xor U24677 (N_24677,N_24321,N_24436);
nor U24678 (N_24678,N_24529,N_24488);
xor U24679 (N_24679,N_24349,N_24421);
or U24680 (N_24680,N_24358,N_24257);
xnor U24681 (N_24681,N_24519,N_24212);
nand U24682 (N_24682,N_24105,N_24460);
nand U24683 (N_24683,N_24338,N_24229);
or U24684 (N_24684,N_24491,N_24284);
nor U24685 (N_24685,N_24298,N_24554);
nor U24686 (N_24686,N_24547,N_24148);
nand U24687 (N_24687,N_24184,N_24087);
or U24688 (N_24688,N_24490,N_24264);
nor U24689 (N_24689,N_24084,N_24079);
and U24690 (N_24690,N_24058,N_24536);
or U24691 (N_24691,N_24383,N_24394);
nor U24692 (N_24692,N_24124,N_24070);
or U24693 (N_24693,N_24438,N_24113);
and U24694 (N_24694,N_24251,N_24277);
nand U24695 (N_24695,N_24275,N_24326);
nor U24696 (N_24696,N_24520,N_24119);
nand U24697 (N_24697,N_24019,N_24329);
nor U24698 (N_24698,N_24594,N_24246);
nor U24699 (N_24699,N_24361,N_24328);
nand U24700 (N_24700,N_24158,N_24353);
or U24701 (N_24701,N_24595,N_24342);
nand U24702 (N_24702,N_24514,N_24416);
nand U24703 (N_24703,N_24433,N_24231);
or U24704 (N_24704,N_24027,N_24579);
xnor U24705 (N_24705,N_24458,N_24265);
or U24706 (N_24706,N_24278,N_24054);
and U24707 (N_24707,N_24535,N_24463);
nor U24708 (N_24708,N_24343,N_24272);
xnor U24709 (N_24709,N_24498,N_24374);
nand U24710 (N_24710,N_24260,N_24130);
or U24711 (N_24711,N_24128,N_24106);
nor U24712 (N_24712,N_24572,N_24359);
or U24713 (N_24713,N_24325,N_24472);
or U24714 (N_24714,N_24245,N_24144);
xnor U24715 (N_24715,N_24367,N_24454);
or U24716 (N_24716,N_24164,N_24410);
nand U24717 (N_24717,N_24197,N_24234);
and U24718 (N_24718,N_24363,N_24409);
nand U24719 (N_24719,N_24426,N_24558);
or U24720 (N_24720,N_24189,N_24177);
or U24721 (N_24721,N_24140,N_24292);
and U24722 (N_24722,N_24440,N_24061);
nand U24723 (N_24723,N_24012,N_24240);
xnor U24724 (N_24724,N_24503,N_24532);
and U24725 (N_24725,N_24443,N_24333);
nand U24726 (N_24726,N_24317,N_24220);
xnor U24727 (N_24727,N_24521,N_24073);
or U24728 (N_24728,N_24495,N_24392);
and U24729 (N_24729,N_24527,N_24100);
or U24730 (N_24730,N_24166,N_24280);
nor U24731 (N_24731,N_24171,N_24088);
or U24732 (N_24732,N_24053,N_24159);
or U24733 (N_24733,N_24439,N_24437);
nand U24734 (N_24734,N_24095,N_24501);
and U24735 (N_24735,N_24468,N_24287);
or U24736 (N_24736,N_24223,N_24219);
nor U24737 (N_24737,N_24552,N_24340);
and U24738 (N_24738,N_24448,N_24543);
nand U24739 (N_24739,N_24592,N_24085);
nand U24740 (N_24740,N_24065,N_24169);
xor U24741 (N_24741,N_24121,N_24530);
nand U24742 (N_24742,N_24068,N_24139);
and U24743 (N_24743,N_24003,N_24269);
or U24744 (N_24744,N_24243,N_24441);
or U24745 (N_24745,N_24395,N_24494);
and U24746 (N_24746,N_24055,N_24232);
and U24747 (N_24747,N_24249,N_24183);
xnor U24748 (N_24748,N_24320,N_24567);
nand U24749 (N_24749,N_24487,N_24563);
or U24750 (N_24750,N_24550,N_24001);
xor U24751 (N_24751,N_24045,N_24035);
and U24752 (N_24752,N_24282,N_24492);
or U24753 (N_24753,N_24489,N_24150);
nand U24754 (N_24754,N_24236,N_24090);
nor U24755 (N_24755,N_24467,N_24308);
nand U24756 (N_24756,N_24526,N_24324);
and U24757 (N_24757,N_24515,N_24323);
and U24758 (N_24758,N_24014,N_24261);
nand U24759 (N_24759,N_24344,N_24200);
or U24760 (N_24760,N_24037,N_24499);
nor U24761 (N_24761,N_24017,N_24071);
nor U24762 (N_24762,N_24496,N_24135);
xnor U24763 (N_24763,N_24029,N_24315);
and U24764 (N_24764,N_24201,N_24466);
xor U24765 (N_24765,N_24290,N_24575);
nand U24766 (N_24766,N_24332,N_24120);
or U24767 (N_24767,N_24242,N_24411);
nand U24768 (N_24768,N_24346,N_24393);
and U24769 (N_24769,N_24388,N_24507);
nand U24770 (N_24770,N_24406,N_24129);
nand U24771 (N_24771,N_24313,N_24557);
nand U24772 (N_24772,N_24218,N_24078);
or U24773 (N_24773,N_24141,N_24096);
nand U24774 (N_24774,N_24194,N_24271);
or U24775 (N_24775,N_24258,N_24414);
nand U24776 (N_24776,N_24186,N_24362);
nand U24777 (N_24777,N_24146,N_24123);
or U24778 (N_24778,N_24390,N_24077);
nor U24779 (N_24779,N_24170,N_24137);
xnor U24780 (N_24780,N_24480,N_24209);
or U24781 (N_24781,N_24449,N_24576);
nand U24782 (N_24782,N_24339,N_24109);
nor U24783 (N_24783,N_24556,N_24504);
and U24784 (N_24784,N_24156,N_24180);
and U24785 (N_24785,N_24596,N_24191);
or U24786 (N_24786,N_24214,N_24522);
and U24787 (N_24787,N_24115,N_24226);
nor U24788 (N_24788,N_24402,N_24452);
and U24789 (N_24789,N_24401,N_24295);
or U24790 (N_24790,N_24018,N_24046);
nor U24791 (N_24791,N_24122,N_24179);
and U24792 (N_24792,N_24005,N_24587);
nor U24793 (N_24793,N_24569,N_24133);
xor U24794 (N_24794,N_24161,N_24373);
or U24795 (N_24795,N_24375,N_24493);
or U24796 (N_24796,N_24250,N_24112);
nand U24797 (N_24797,N_24217,N_24285);
or U24798 (N_24798,N_24002,N_24478);
and U24799 (N_24799,N_24281,N_24291);
xnor U24800 (N_24800,N_24331,N_24380);
xnor U24801 (N_24801,N_24108,N_24407);
nor U24802 (N_24802,N_24294,N_24043);
nand U24803 (N_24803,N_24176,N_24368);
nor U24804 (N_24804,N_24127,N_24233);
or U24805 (N_24805,N_24583,N_24152);
xnor U24806 (N_24806,N_24465,N_24064);
xnor U24807 (N_24807,N_24412,N_24050);
nand U24808 (N_24808,N_24435,N_24500);
nor U24809 (N_24809,N_24473,N_24523);
nand U24810 (N_24810,N_24126,N_24387);
nand U24811 (N_24811,N_24210,N_24091);
and U24812 (N_24812,N_24136,N_24199);
xor U24813 (N_24813,N_24069,N_24549);
or U24814 (N_24814,N_24221,N_24153);
nor U24815 (N_24815,N_24479,N_24561);
nor U24816 (N_24816,N_24364,N_24048);
xor U24817 (N_24817,N_24372,N_24247);
nand U24818 (N_24818,N_24539,N_24428);
and U24819 (N_24819,N_24445,N_24581);
nand U24820 (N_24820,N_24314,N_24267);
xor U24821 (N_24821,N_24155,N_24270);
and U24822 (N_24822,N_24036,N_24542);
nor U24823 (N_24823,N_24060,N_24013);
nor U24824 (N_24824,N_24382,N_24582);
xnor U24825 (N_24825,N_24016,N_24198);
nor U24826 (N_24826,N_24351,N_24007);
nor U24827 (N_24827,N_24033,N_24216);
or U24828 (N_24828,N_24310,N_24178);
xnor U24829 (N_24829,N_24512,N_24098);
xor U24830 (N_24830,N_24470,N_24385);
and U24831 (N_24831,N_24534,N_24531);
nor U24832 (N_24832,N_24103,N_24072);
nand U24833 (N_24833,N_24429,N_24293);
xnor U24834 (N_24834,N_24360,N_24238);
xor U24835 (N_24835,N_24255,N_24312);
and U24836 (N_24836,N_24506,N_24415);
xor U24837 (N_24837,N_24546,N_24588);
or U24838 (N_24838,N_24305,N_24303);
nand U24839 (N_24839,N_24211,N_24094);
nand U24840 (N_24840,N_24020,N_24371);
and U24841 (N_24841,N_24134,N_24509);
or U24842 (N_24842,N_24599,N_24354);
and U24843 (N_24843,N_24334,N_24525);
nor U24844 (N_24844,N_24336,N_24059);
nand U24845 (N_24845,N_24202,N_24102);
nand U24846 (N_24846,N_24469,N_24051);
nand U24847 (N_24847,N_24397,N_24208);
xor U24848 (N_24848,N_24319,N_24299);
and U24849 (N_24849,N_24022,N_24337);
and U24850 (N_24850,N_24142,N_24379);
nor U24851 (N_24851,N_24540,N_24193);
nor U24852 (N_24852,N_24224,N_24235);
nor U24853 (N_24853,N_24541,N_24391);
nor U24854 (N_24854,N_24276,N_24039);
and U24855 (N_24855,N_24398,N_24419);
nor U24856 (N_24856,N_24352,N_24427);
nor U24857 (N_24857,N_24505,N_24041);
nor U24858 (N_24858,N_24483,N_24101);
nand U24859 (N_24859,N_24040,N_24566);
and U24860 (N_24860,N_24289,N_24350);
nor U24861 (N_24861,N_24545,N_24425);
xor U24862 (N_24862,N_24032,N_24075);
nor U24863 (N_24863,N_24175,N_24400);
and U24864 (N_24864,N_24031,N_24564);
and U24865 (N_24865,N_24396,N_24377);
nor U24866 (N_24866,N_24010,N_24574);
and U24867 (N_24867,N_24405,N_24000);
xor U24868 (N_24868,N_24185,N_24162);
nand U24869 (N_24869,N_24192,N_24455);
xor U24870 (N_24870,N_24432,N_24279);
and U24871 (N_24871,N_24370,N_24413);
nand U24872 (N_24872,N_24524,N_24590);
nor U24873 (N_24873,N_24187,N_24225);
and U24874 (N_24874,N_24021,N_24215);
nand U24875 (N_24875,N_24066,N_24389);
or U24876 (N_24876,N_24456,N_24565);
xnor U24877 (N_24877,N_24369,N_24024);
or U24878 (N_24878,N_24099,N_24172);
nand U24879 (N_24879,N_24026,N_24571);
or U24880 (N_24880,N_24006,N_24254);
and U24881 (N_24881,N_24283,N_24132);
xnor U24882 (N_24882,N_24485,N_24086);
nor U24883 (N_24883,N_24163,N_24259);
or U24884 (N_24884,N_24513,N_24273);
and U24885 (N_24885,N_24528,N_24174);
or U24886 (N_24886,N_24038,N_24399);
nand U24887 (N_24887,N_24537,N_24457);
nand U24888 (N_24888,N_24107,N_24047);
or U24889 (N_24889,N_24076,N_24004);
xor U24890 (N_24890,N_24553,N_24067);
xnor U24891 (N_24891,N_24030,N_24580);
nand U24892 (N_24892,N_24355,N_24598);
nand U24893 (N_24893,N_24573,N_24301);
and U24894 (N_24894,N_24453,N_24450);
nand U24895 (N_24895,N_24239,N_24316);
nand U24896 (N_24896,N_24302,N_24207);
and U24897 (N_24897,N_24114,N_24266);
nor U24898 (N_24898,N_24335,N_24464);
nor U24899 (N_24899,N_24434,N_24327);
and U24900 (N_24900,N_24414,N_24185);
or U24901 (N_24901,N_24153,N_24556);
and U24902 (N_24902,N_24348,N_24501);
or U24903 (N_24903,N_24119,N_24364);
xnor U24904 (N_24904,N_24084,N_24529);
and U24905 (N_24905,N_24083,N_24585);
and U24906 (N_24906,N_24192,N_24420);
nand U24907 (N_24907,N_24597,N_24231);
nand U24908 (N_24908,N_24409,N_24012);
and U24909 (N_24909,N_24388,N_24535);
and U24910 (N_24910,N_24272,N_24374);
nand U24911 (N_24911,N_24557,N_24581);
xnor U24912 (N_24912,N_24378,N_24201);
nand U24913 (N_24913,N_24310,N_24165);
nand U24914 (N_24914,N_24079,N_24247);
and U24915 (N_24915,N_24358,N_24108);
or U24916 (N_24916,N_24597,N_24526);
xnor U24917 (N_24917,N_24098,N_24387);
nor U24918 (N_24918,N_24095,N_24020);
or U24919 (N_24919,N_24014,N_24093);
nand U24920 (N_24920,N_24163,N_24286);
nor U24921 (N_24921,N_24058,N_24090);
nor U24922 (N_24922,N_24261,N_24249);
nand U24923 (N_24923,N_24336,N_24516);
nand U24924 (N_24924,N_24041,N_24417);
xor U24925 (N_24925,N_24003,N_24372);
or U24926 (N_24926,N_24579,N_24509);
nand U24927 (N_24927,N_24470,N_24300);
nand U24928 (N_24928,N_24194,N_24327);
nand U24929 (N_24929,N_24372,N_24298);
nor U24930 (N_24930,N_24297,N_24271);
and U24931 (N_24931,N_24590,N_24582);
nand U24932 (N_24932,N_24478,N_24435);
nand U24933 (N_24933,N_24322,N_24276);
or U24934 (N_24934,N_24367,N_24042);
and U24935 (N_24935,N_24200,N_24021);
or U24936 (N_24936,N_24108,N_24174);
or U24937 (N_24937,N_24455,N_24217);
nand U24938 (N_24938,N_24011,N_24362);
nand U24939 (N_24939,N_24269,N_24483);
or U24940 (N_24940,N_24012,N_24543);
xnor U24941 (N_24941,N_24039,N_24433);
nand U24942 (N_24942,N_24011,N_24047);
and U24943 (N_24943,N_24088,N_24548);
and U24944 (N_24944,N_24082,N_24561);
xnor U24945 (N_24945,N_24252,N_24310);
xnor U24946 (N_24946,N_24420,N_24359);
and U24947 (N_24947,N_24455,N_24257);
xnor U24948 (N_24948,N_24155,N_24589);
and U24949 (N_24949,N_24489,N_24426);
or U24950 (N_24950,N_24313,N_24365);
nand U24951 (N_24951,N_24005,N_24053);
and U24952 (N_24952,N_24411,N_24000);
nor U24953 (N_24953,N_24229,N_24465);
nand U24954 (N_24954,N_24510,N_24152);
nor U24955 (N_24955,N_24405,N_24126);
and U24956 (N_24956,N_24043,N_24540);
nand U24957 (N_24957,N_24026,N_24474);
nor U24958 (N_24958,N_24197,N_24380);
xnor U24959 (N_24959,N_24020,N_24534);
and U24960 (N_24960,N_24587,N_24277);
and U24961 (N_24961,N_24175,N_24112);
and U24962 (N_24962,N_24597,N_24474);
or U24963 (N_24963,N_24418,N_24516);
xnor U24964 (N_24964,N_24421,N_24283);
and U24965 (N_24965,N_24438,N_24576);
nor U24966 (N_24966,N_24156,N_24483);
nor U24967 (N_24967,N_24088,N_24282);
or U24968 (N_24968,N_24179,N_24047);
nor U24969 (N_24969,N_24140,N_24586);
nor U24970 (N_24970,N_24562,N_24423);
or U24971 (N_24971,N_24041,N_24020);
nand U24972 (N_24972,N_24152,N_24433);
nor U24973 (N_24973,N_24251,N_24404);
and U24974 (N_24974,N_24085,N_24186);
nor U24975 (N_24975,N_24405,N_24312);
nor U24976 (N_24976,N_24246,N_24165);
and U24977 (N_24977,N_24059,N_24120);
and U24978 (N_24978,N_24390,N_24389);
or U24979 (N_24979,N_24548,N_24428);
nand U24980 (N_24980,N_24405,N_24338);
and U24981 (N_24981,N_24077,N_24013);
nor U24982 (N_24982,N_24220,N_24182);
and U24983 (N_24983,N_24448,N_24425);
xnor U24984 (N_24984,N_24194,N_24445);
or U24985 (N_24985,N_24524,N_24067);
and U24986 (N_24986,N_24041,N_24490);
or U24987 (N_24987,N_24537,N_24531);
nor U24988 (N_24988,N_24507,N_24170);
nand U24989 (N_24989,N_24049,N_24097);
or U24990 (N_24990,N_24000,N_24076);
nand U24991 (N_24991,N_24205,N_24542);
xnor U24992 (N_24992,N_24229,N_24150);
nand U24993 (N_24993,N_24517,N_24060);
nand U24994 (N_24994,N_24012,N_24102);
and U24995 (N_24995,N_24473,N_24338);
or U24996 (N_24996,N_24192,N_24525);
nor U24997 (N_24997,N_24262,N_24177);
nand U24998 (N_24998,N_24315,N_24186);
xnor U24999 (N_24999,N_24276,N_24504);
xor U25000 (N_25000,N_24443,N_24372);
and U25001 (N_25001,N_24206,N_24155);
xor U25002 (N_25002,N_24256,N_24156);
nor U25003 (N_25003,N_24009,N_24013);
and U25004 (N_25004,N_24265,N_24362);
and U25005 (N_25005,N_24326,N_24596);
nand U25006 (N_25006,N_24421,N_24439);
and U25007 (N_25007,N_24369,N_24402);
nor U25008 (N_25008,N_24414,N_24014);
xnor U25009 (N_25009,N_24095,N_24399);
or U25010 (N_25010,N_24589,N_24323);
and U25011 (N_25011,N_24540,N_24303);
or U25012 (N_25012,N_24564,N_24502);
or U25013 (N_25013,N_24160,N_24313);
xnor U25014 (N_25014,N_24438,N_24515);
xor U25015 (N_25015,N_24194,N_24238);
or U25016 (N_25016,N_24125,N_24342);
or U25017 (N_25017,N_24273,N_24327);
nor U25018 (N_25018,N_24225,N_24385);
nand U25019 (N_25019,N_24578,N_24047);
nand U25020 (N_25020,N_24194,N_24064);
xor U25021 (N_25021,N_24578,N_24477);
and U25022 (N_25022,N_24166,N_24169);
or U25023 (N_25023,N_24260,N_24063);
nand U25024 (N_25024,N_24528,N_24082);
xor U25025 (N_25025,N_24530,N_24249);
nand U25026 (N_25026,N_24465,N_24554);
or U25027 (N_25027,N_24406,N_24507);
nand U25028 (N_25028,N_24275,N_24465);
xnor U25029 (N_25029,N_24472,N_24199);
nand U25030 (N_25030,N_24106,N_24006);
and U25031 (N_25031,N_24295,N_24064);
and U25032 (N_25032,N_24481,N_24139);
nor U25033 (N_25033,N_24085,N_24107);
nand U25034 (N_25034,N_24540,N_24041);
or U25035 (N_25035,N_24487,N_24253);
xor U25036 (N_25036,N_24120,N_24363);
and U25037 (N_25037,N_24083,N_24526);
nor U25038 (N_25038,N_24464,N_24443);
and U25039 (N_25039,N_24121,N_24304);
and U25040 (N_25040,N_24244,N_24113);
nor U25041 (N_25041,N_24483,N_24435);
xnor U25042 (N_25042,N_24231,N_24458);
nand U25043 (N_25043,N_24161,N_24465);
xnor U25044 (N_25044,N_24283,N_24570);
nand U25045 (N_25045,N_24517,N_24216);
or U25046 (N_25046,N_24099,N_24429);
and U25047 (N_25047,N_24524,N_24113);
nand U25048 (N_25048,N_24553,N_24252);
nand U25049 (N_25049,N_24159,N_24063);
nor U25050 (N_25050,N_24086,N_24348);
nand U25051 (N_25051,N_24547,N_24055);
xnor U25052 (N_25052,N_24219,N_24096);
nand U25053 (N_25053,N_24549,N_24349);
and U25054 (N_25054,N_24368,N_24316);
and U25055 (N_25055,N_24231,N_24123);
nor U25056 (N_25056,N_24419,N_24011);
nand U25057 (N_25057,N_24286,N_24029);
xnor U25058 (N_25058,N_24576,N_24346);
and U25059 (N_25059,N_24232,N_24287);
nor U25060 (N_25060,N_24124,N_24472);
xnor U25061 (N_25061,N_24515,N_24542);
xnor U25062 (N_25062,N_24396,N_24063);
and U25063 (N_25063,N_24431,N_24144);
nor U25064 (N_25064,N_24465,N_24558);
and U25065 (N_25065,N_24515,N_24436);
xor U25066 (N_25066,N_24131,N_24455);
nand U25067 (N_25067,N_24167,N_24029);
and U25068 (N_25068,N_24262,N_24559);
and U25069 (N_25069,N_24053,N_24214);
nand U25070 (N_25070,N_24489,N_24497);
or U25071 (N_25071,N_24159,N_24196);
nor U25072 (N_25072,N_24202,N_24408);
nor U25073 (N_25073,N_24437,N_24447);
and U25074 (N_25074,N_24172,N_24217);
xor U25075 (N_25075,N_24244,N_24127);
nand U25076 (N_25076,N_24029,N_24195);
nand U25077 (N_25077,N_24332,N_24588);
nand U25078 (N_25078,N_24062,N_24246);
nand U25079 (N_25079,N_24366,N_24411);
nor U25080 (N_25080,N_24279,N_24401);
nor U25081 (N_25081,N_24151,N_24376);
nand U25082 (N_25082,N_24055,N_24132);
nor U25083 (N_25083,N_24138,N_24270);
nor U25084 (N_25084,N_24423,N_24234);
nor U25085 (N_25085,N_24537,N_24120);
and U25086 (N_25086,N_24442,N_24326);
nor U25087 (N_25087,N_24308,N_24092);
or U25088 (N_25088,N_24278,N_24125);
and U25089 (N_25089,N_24327,N_24091);
xnor U25090 (N_25090,N_24385,N_24520);
nand U25091 (N_25091,N_24045,N_24092);
xnor U25092 (N_25092,N_24375,N_24510);
nand U25093 (N_25093,N_24571,N_24599);
nand U25094 (N_25094,N_24190,N_24211);
xor U25095 (N_25095,N_24034,N_24113);
nor U25096 (N_25096,N_24089,N_24243);
and U25097 (N_25097,N_24157,N_24425);
xnor U25098 (N_25098,N_24484,N_24595);
or U25099 (N_25099,N_24271,N_24554);
nor U25100 (N_25100,N_24325,N_24090);
nor U25101 (N_25101,N_24110,N_24311);
xor U25102 (N_25102,N_24383,N_24041);
and U25103 (N_25103,N_24069,N_24159);
nand U25104 (N_25104,N_24378,N_24101);
or U25105 (N_25105,N_24574,N_24327);
nor U25106 (N_25106,N_24287,N_24044);
or U25107 (N_25107,N_24154,N_24009);
xnor U25108 (N_25108,N_24142,N_24450);
xnor U25109 (N_25109,N_24584,N_24244);
and U25110 (N_25110,N_24072,N_24056);
or U25111 (N_25111,N_24004,N_24385);
and U25112 (N_25112,N_24348,N_24246);
nand U25113 (N_25113,N_24499,N_24237);
and U25114 (N_25114,N_24514,N_24063);
and U25115 (N_25115,N_24278,N_24076);
and U25116 (N_25116,N_24314,N_24152);
nor U25117 (N_25117,N_24410,N_24258);
and U25118 (N_25118,N_24086,N_24441);
xor U25119 (N_25119,N_24231,N_24167);
nor U25120 (N_25120,N_24142,N_24330);
xnor U25121 (N_25121,N_24450,N_24129);
xor U25122 (N_25122,N_24180,N_24187);
nand U25123 (N_25123,N_24256,N_24561);
nor U25124 (N_25124,N_24569,N_24570);
nand U25125 (N_25125,N_24494,N_24037);
and U25126 (N_25126,N_24532,N_24205);
nor U25127 (N_25127,N_24460,N_24173);
or U25128 (N_25128,N_24036,N_24038);
or U25129 (N_25129,N_24290,N_24138);
or U25130 (N_25130,N_24294,N_24274);
xor U25131 (N_25131,N_24158,N_24007);
nand U25132 (N_25132,N_24390,N_24140);
nand U25133 (N_25133,N_24396,N_24562);
and U25134 (N_25134,N_24523,N_24221);
nor U25135 (N_25135,N_24079,N_24296);
and U25136 (N_25136,N_24232,N_24336);
nor U25137 (N_25137,N_24477,N_24414);
nor U25138 (N_25138,N_24386,N_24531);
nor U25139 (N_25139,N_24406,N_24425);
and U25140 (N_25140,N_24367,N_24538);
nor U25141 (N_25141,N_24028,N_24481);
nand U25142 (N_25142,N_24369,N_24131);
nand U25143 (N_25143,N_24542,N_24006);
nor U25144 (N_25144,N_24005,N_24526);
xor U25145 (N_25145,N_24025,N_24093);
nor U25146 (N_25146,N_24055,N_24533);
nor U25147 (N_25147,N_24023,N_24438);
nand U25148 (N_25148,N_24488,N_24266);
nand U25149 (N_25149,N_24096,N_24254);
or U25150 (N_25150,N_24292,N_24137);
nand U25151 (N_25151,N_24361,N_24542);
and U25152 (N_25152,N_24188,N_24426);
and U25153 (N_25153,N_24087,N_24182);
xor U25154 (N_25154,N_24439,N_24183);
or U25155 (N_25155,N_24471,N_24187);
or U25156 (N_25156,N_24092,N_24305);
and U25157 (N_25157,N_24334,N_24371);
nand U25158 (N_25158,N_24365,N_24465);
xnor U25159 (N_25159,N_24357,N_24218);
nand U25160 (N_25160,N_24244,N_24274);
xor U25161 (N_25161,N_24037,N_24549);
xor U25162 (N_25162,N_24535,N_24543);
xor U25163 (N_25163,N_24343,N_24427);
or U25164 (N_25164,N_24549,N_24011);
nor U25165 (N_25165,N_24444,N_24343);
and U25166 (N_25166,N_24488,N_24235);
xnor U25167 (N_25167,N_24201,N_24527);
or U25168 (N_25168,N_24529,N_24509);
or U25169 (N_25169,N_24373,N_24186);
and U25170 (N_25170,N_24200,N_24418);
nand U25171 (N_25171,N_24549,N_24251);
and U25172 (N_25172,N_24437,N_24388);
or U25173 (N_25173,N_24246,N_24256);
nor U25174 (N_25174,N_24369,N_24125);
nor U25175 (N_25175,N_24447,N_24308);
and U25176 (N_25176,N_24277,N_24334);
nor U25177 (N_25177,N_24594,N_24479);
nand U25178 (N_25178,N_24103,N_24104);
and U25179 (N_25179,N_24098,N_24329);
nor U25180 (N_25180,N_24434,N_24279);
nand U25181 (N_25181,N_24188,N_24323);
or U25182 (N_25182,N_24081,N_24231);
and U25183 (N_25183,N_24214,N_24452);
nand U25184 (N_25184,N_24254,N_24074);
or U25185 (N_25185,N_24126,N_24190);
or U25186 (N_25186,N_24577,N_24284);
and U25187 (N_25187,N_24270,N_24509);
and U25188 (N_25188,N_24172,N_24491);
and U25189 (N_25189,N_24481,N_24564);
nor U25190 (N_25190,N_24211,N_24198);
nand U25191 (N_25191,N_24385,N_24348);
nand U25192 (N_25192,N_24528,N_24497);
nand U25193 (N_25193,N_24483,N_24539);
or U25194 (N_25194,N_24571,N_24317);
nor U25195 (N_25195,N_24373,N_24033);
and U25196 (N_25196,N_24453,N_24220);
xor U25197 (N_25197,N_24405,N_24188);
or U25198 (N_25198,N_24515,N_24181);
nor U25199 (N_25199,N_24024,N_24306);
xnor U25200 (N_25200,N_25127,N_24655);
nand U25201 (N_25201,N_24610,N_24744);
and U25202 (N_25202,N_24693,N_24681);
or U25203 (N_25203,N_24638,N_24921);
or U25204 (N_25204,N_25153,N_24828);
nor U25205 (N_25205,N_24682,N_24779);
and U25206 (N_25206,N_24657,N_24847);
nor U25207 (N_25207,N_25154,N_24618);
and U25208 (N_25208,N_25059,N_24943);
and U25209 (N_25209,N_24628,N_25175);
nor U25210 (N_25210,N_24683,N_24709);
xnor U25211 (N_25211,N_25198,N_24733);
nor U25212 (N_25212,N_25194,N_24864);
xor U25213 (N_25213,N_24947,N_25079);
and U25214 (N_25214,N_25117,N_24926);
or U25215 (N_25215,N_25073,N_25080);
or U25216 (N_25216,N_24901,N_24957);
nand U25217 (N_25217,N_24692,N_24656);
and U25218 (N_25218,N_24713,N_24839);
or U25219 (N_25219,N_24939,N_24814);
nor U25220 (N_25220,N_24953,N_24803);
nor U25221 (N_25221,N_24626,N_24894);
nand U25222 (N_25222,N_24609,N_24930);
nand U25223 (N_25223,N_24867,N_24677);
or U25224 (N_25224,N_25142,N_24885);
xor U25225 (N_25225,N_24750,N_24646);
or U25226 (N_25226,N_25022,N_25109);
nand U25227 (N_25227,N_24938,N_25169);
nand U25228 (N_25228,N_24747,N_25129);
xnor U25229 (N_25229,N_24667,N_24798);
nand U25230 (N_25230,N_24740,N_24652);
or U25231 (N_25231,N_25160,N_24844);
and U25232 (N_25232,N_24927,N_25078);
and U25233 (N_25233,N_24691,N_25102);
xor U25234 (N_25234,N_24600,N_24820);
nand U25235 (N_25235,N_24634,N_24823);
nand U25236 (N_25236,N_24649,N_25062);
nor U25237 (N_25237,N_25068,N_24995);
nor U25238 (N_25238,N_25170,N_24605);
and U25239 (N_25239,N_25005,N_25106);
xor U25240 (N_25240,N_25029,N_24854);
xor U25241 (N_25241,N_25074,N_24853);
nor U25242 (N_25242,N_24857,N_24822);
nor U25243 (N_25243,N_24819,N_24883);
nand U25244 (N_25244,N_25152,N_25027);
nand U25245 (N_25245,N_24678,N_24862);
nand U25246 (N_25246,N_24909,N_24759);
or U25247 (N_25247,N_25049,N_24698);
and U25248 (N_25248,N_25051,N_24662);
and U25249 (N_25249,N_24623,N_25008);
nor U25250 (N_25250,N_24858,N_25077);
and U25251 (N_25251,N_25112,N_25017);
or U25252 (N_25252,N_24635,N_24888);
or U25253 (N_25253,N_24933,N_24992);
and U25254 (N_25254,N_24919,N_24711);
and U25255 (N_25255,N_25039,N_24818);
nand U25256 (N_25256,N_24726,N_25067);
or U25257 (N_25257,N_25124,N_25081);
or U25258 (N_25258,N_24615,N_24967);
nand U25259 (N_25259,N_25173,N_25013);
and U25260 (N_25260,N_24602,N_24668);
nor U25261 (N_25261,N_24684,N_24651);
nor U25262 (N_25262,N_24703,N_24714);
xor U25263 (N_25263,N_24948,N_25133);
nand U25264 (N_25264,N_24757,N_25063);
and U25265 (N_25265,N_24986,N_25018);
and U25266 (N_25266,N_24619,N_25024);
nor U25267 (N_25267,N_25099,N_24984);
and U25268 (N_25268,N_24834,N_25189);
or U25269 (N_25269,N_24617,N_24647);
nor U25270 (N_25270,N_24731,N_24643);
or U25271 (N_25271,N_25108,N_24782);
and U25272 (N_25272,N_24763,N_24800);
and U25273 (N_25273,N_24846,N_25033);
and U25274 (N_25274,N_25015,N_24879);
and U25275 (N_25275,N_24966,N_25178);
xnor U25276 (N_25276,N_24767,N_24704);
or U25277 (N_25277,N_24607,N_25149);
and U25278 (N_25278,N_25076,N_25028);
and U25279 (N_25279,N_24810,N_25016);
or U25280 (N_25280,N_24781,N_24971);
nor U25281 (N_25281,N_24701,N_24985);
nand U25282 (N_25282,N_25192,N_24778);
and U25283 (N_25283,N_24771,N_25146);
nor U25284 (N_25284,N_25058,N_24848);
or U25285 (N_25285,N_25164,N_24842);
or U25286 (N_25286,N_25085,N_24755);
or U25287 (N_25287,N_24809,N_24812);
nand U25288 (N_25288,N_24764,N_25140);
nand U25289 (N_25289,N_24807,N_25054);
and U25290 (N_25290,N_25092,N_25158);
and U25291 (N_25291,N_24849,N_24949);
nor U25292 (N_25292,N_25037,N_25019);
and U25293 (N_25293,N_24608,N_24772);
or U25294 (N_25294,N_24773,N_24811);
nand U25295 (N_25295,N_24843,N_25100);
and U25296 (N_25296,N_25126,N_25188);
xnor U25297 (N_25297,N_24737,N_24994);
or U25298 (N_25298,N_24951,N_24792);
xor U25299 (N_25299,N_24793,N_24787);
or U25300 (N_25300,N_25143,N_25093);
xor U25301 (N_25301,N_24753,N_24616);
or U25302 (N_25302,N_24614,N_24936);
nor U25303 (N_25303,N_24650,N_24718);
and U25304 (N_25304,N_24940,N_25199);
nand U25305 (N_25305,N_24962,N_24913);
nor U25306 (N_25306,N_24873,N_24897);
xnor U25307 (N_25307,N_25057,N_24836);
or U25308 (N_25308,N_24606,N_25046);
and U25309 (N_25309,N_24659,N_24769);
or U25310 (N_25310,N_25113,N_25052);
or U25311 (N_25311,N_25044,N_24878);
and U25312 (N_25312,N_25034,N_25196);
xnor U25313 (N_25313,N_25134,N_25191);
xor U25314 (N_25314,N_25061,N_24892);
nand U25315 (N_25315,N_24841,N_24983);
and U25316 (N_25316,N_24804,N_24770);
nor U25317 (N_25317,N_25171,N_24723);
and U25318 (N_25318,N_24738,N_24776);
and U25319 (N_25319,N_25165,N_24758);
nor U25320 (N_25320,N_24861,N_25050);
nand U25321 (N_25321,N_25090,N_25060);
nor U25322 (N_25322,N_24956,N_24993);
and U25323 (N_25323,N_24838,N_24870);
or U25324 (N_25324,N_24761,N_24627);
or U25325 (N_25325,N_25003,N_24826);
and U25326 (N_25326,N_24961,N_24912);
xor U25327 (N_25327,N_25066,N_24699);
and U25328 (N_25328,N_24790,N_24968);
nor U25329 (N_25329,N_25184,N_24998);
nand U25330 (N_25330,N_24697,N_24902);
nor U25331 (N_25331,N_24831,N_24664);
xor U25332 (N_25332,N_24722,N_25098);
or U25333 (N_25333,N_24815,N_25159);
or U25334 (N_25334,N_24702,N_24910);
or U25335 (N_25335,N_24881,N_25130);
nor U25336 (N_25336,N_24629,N_24865);
or U25337 (N_25337,N_25135,N_24869);
and U25338 (N_25338,N_24695,N_25040);
xnor U25339 (N_25339,N_24945,N_24988);
nor U25340 (N_25340,N_24884,N_24837);
or U25341 (N_25341,N_24777,N_24908);
nor U25342 (N_25342,N_24954,N_25045);
and U25343 (N_25343,N_24641,N_25089);
and U25344 (N_25344,N_24795,N_25055);
nor U25345 (N_25345,N_24707,N_24970);
xor U25346 (N_25346,N_25035,N_24708);
nor U25347 (N_25347,N_25101,N_24710);
xnor U25348 (N_25348,N_24705,N_25123);
and U25349 (N_25349,N_24904,N_24712);
or U25350 (N_25350,N_24833,N_24775);
nand U25351 (N_25351,N_25043,N_25048);
and U25352 (N_25352,N_25095,N_24687);
xnor U25353 (N_25353,N_25163,N_24829);
or U25354 (N_25354,N_24794,N_24788);
or U25355 (N_25355,N_24631,N_24832);
xnor U25356 (N_25356,N_24673,N_25084);
and U25357 (N_25357,N_25125,N_25172);
and U25358 (N_25358,N_24745,N_24715);
nor U25359 (N_25359,N_24907,N_24625);
or U25360 (N_25360,N_24851,N_24721);
nand U25361 (N_25361,N_24696,N_24982);
and U25362 (N_25362,N_24613,N_24825);
xor U25363 (N_25363,N_24932,N_24784);
nand U25364 (N_25364,N_25021,N_24654);
or U25365 (N_25365,N_24855,N_24665);
xnor U25366 (N_25366,N_24931,N_25150);
nor U25367 (N_25367,N_25010,N_25197);
nor U25368 (N_25368,N_24866,N_25011);
and U25369 (N_25369,N_25156,N_24887);
nor U25370 (N_25370,N_24955,N_24974);
nor U25371 (N_25371,N_25183,N_24666);
xnor U25372 (N_25372,N_24964,N_25138);
nor U25373 (N_25373,N_24690,N_25069);
and U25374 (N_25374,N_25176,N_24632);
xnor U25375 (N_25375,N_24719,N_24989);
nand U25376 (N_25376,N_24746,N_24880);
nand U25377 (N_25377,N_24679,N_24969);
and U25378 (N_25378,N_24856,N_24742);
nor U25379 (N_25379,N_25025,N_24749);
or U25380 (N_25380,N_24729,N_24941);
or U25381 (N_25381,N_24845,N_24893);
and U25382 (N_25382,N_25121,N_24735);
nor U25383 (N_25383,N_24706,N_25185);
xor U25384 (N_25384,N_24813,N_25056);
nor U25385 (N_25385,N_24914,N_25071);
xnor U25386 (N_25386,N_25120,N_24876);
and U25387 (N_25387,N_24694,N_24996);
nand U25388 (N_25388,N_24975,N_25190);
xnor U25389 (N_25389,N_25026,N_24896);
xor U25390 (N_25390,N_24630,N_24816);
nor U25391 (N_25391,N_24760,N_24732);
xnor U25392 (N_25392,N_24890,N_24979);
nor U25393 (N_25393,N_25115,N_24612);
nor U25394 (N_25394,N_24863,N_24724);
nor U25395 (N_25395,N_24959,N_25122);
or U25396 (N_25396,N_24801,N_24817);
xnor U25397 (N_25397,N_24925,N_24754);
and U25398 (N_25398,N_24874,N_24802);
xor U25399 (N_25399,N_25104,N_24648);
or U25400 (N_25400,N_25137,N_24923);
nor U25401 (N_25401,N_24725,N_25179);
and U25402 (N_25402,N_24620,N_24700);
or U25403 (N_25403,N_25180,N_24786);
xor U25404 (N_25404,N_25001,N_24736);
nor U25405 (N_25405,N_24601,N_25082);
xor U25406 (N_25406,N_24688,N_24999);
nand U25407 (N_25407,N_24644,N_24860);
xnor U25408 (N_25408,N_24899,N_25144);
nor U25409 (N_25409,N_25166,N_25128);
nand U25410 (N_25410,N_25031,N_25155);
and U25411 (N_25411,N_24937,N_25131);
and U25412 (N_25412,N_25009,N_25187);
xor U25413 (N_25413,N_25147,N_24877);
and U25414 (N_25414,N_25020,N_24972);
xnor U25415 (N_25415,N_24977,N_24751);
nand U25416 (N_25416,N_24689,N_24903);
nor U25417 (N_25417,N_25107,N_24991);
nor U25418 (N_25418,N_25119,N_24642);
xor U25419 (N_25419,N_24676,N_24835);
and U25420 (N_25420,N_25000,N_24720);
nor U25421 (N_25421,N_24680,N_24730);
or U25422 (N_25422,N_24850,N_25105);
and U25423 (N_25423,N_25086,N_25139);
nand U25424 (N_25424,N_24789,N_24739);
nor U25425 (N_25425,N_24889,N_25116);
nand U25426 (N_25426,N_24743,N_25036);
nand U25427 (N_25427,N_24797,N_25168);
and U25428 (N_25428,N_25014,N_24780);
and U25429 (N_25429,N_24960,N_24895);
and U25430 (N_25430,N_24728,N_25002);
nand U25431 (N_25431,N_25174,N_24980);
and U25432 (N_25432,N_24952,N_24603);
or U25433 (N_25433,N_24633,N_24727);
nand U25434 (N_25434,N_25177,N_24990);
and U25435 (N_25435,N_24882,N_24906);
or U25436 (N_25436,N_25157,N_25151);
nand U25437 (N_25437,N_25110,N_25181);
nand U25438 (N_25438,N_25096,N_25004);
and U25439 (N_25439,N_25097,N_24924);
and U25440 (N_25440,N_25023,N_24840);
nand U25441 (N_25441,N_24935,N_24766);
nor U25442 (N_25442,N_25103,N_24660);
or U25443 (N_25443,N_24734,N_24671);
and U25444 (N_25444,N_25012,N_24827);
or U25445 (N_25445,N_24808,N_24796);
nand U25446 (N_25446,N_24859,N_24920);
nor U25447 (N_25447,N_24950,N_24783);
and U25448 (N_25448,N_25042,N_25053);
nor U25449 (N_25449,N_25145,N_25141);
and U25450 (N_25450,N_24674,N_24963);
nor U25451 (N_25451,N_24922,N_24806);
xnor U25452 (N_25452,N_25193,N_25148);
or U25453 (N_25453,N_24765,N_24645);
or U25454 (N_25454,N_25006,N_24748);
and U25455 (N_25455,N_25094,N_24622);
and U25456 (N_25456,N_24762,N_25041);
nand U25457 (N_25457,N_25162,N_25065);
nor U25458 (N_25458,N_24672,N_24653);
and U25459 (N_25459,N_24987,N_25182);
nand U25460 (N_25460,N_25064,N_24958);
and U25461 (N_25461,N_24685,N_24621);
xor U25462 (N_25462,N_24717,N_24934);
nor U25463 (N_25463,N_24791,N_25195);
or U25464 (N_25464,N_25186,N_25075);
nand U25465 (N_25465,N_25161,N_24670);
or U25466 (N_25466,N_24973,N_24978);
and U25467 (N_25467,N_24821,N_24875);
nand U25468 (N_25468,N_24965,N_25030);
and U25469 (N_25469,N_24752,N_24799);
xor U25470 (N_25470,N_25118,N_25087);
nand U25471 (N_25471,N_24872,N_25032);
nand U25472 (N_25472,N_25083,N_24917);
or U25473 (N_25473,N_25114,N_24916);
or U25474 (N_25474,N_24658,N_24774);
or U25475 (N_25475,N_25111,N_24944);
nand U25476 (N_25476,N_24981,N_24604);
nand U25477 (N_25477,N_24686,N_24886);
nor U25478 (N_25478,N_24905,N_24942);
nand U25479 (N_25479,N_25132,N_25088);
and U25480 (N_25480,N_24898,N_25047);
or U25481 (N_25481,N_25091,N_24915);
xnor U25482 (N_25482,N_25072,N_24637);
and U25483 (N_25483,N_24624,N_24928);
nor U25484 (N_25484,N_25070,N_25167);
nand U25485 (N_25485,N_24716,N_24830);
nor U25486 (N_25486,N_24824,N_24663);
or U25487 (N_25487,N_25038,N_24871);
nor U25488 (N_25488,N_24768,N_24611);
or U25489 (N_25489,N_24741,N_25007);
and U25490 (N_25490,N_24900,N_24675);
or U25491 (N_25491,N_24946,N_25136);
xnor U25492 (N_25492,N_24661,N_24756);
and U25493 (N_25493,N_24639,N_24868);
xnor U25494 (N_25494,N_24976,N_24852);
nor U25495 (N_25495,N_24805,N_24640);
nor U25496 (N_25496,N_24891,N_24636);
xnor U25497 (N_25497,N_24997,N_24918);
nor U25498 (N_25498,N_24929,N_24911);
nand U25499 (N_25499,N_24785,N_24669);
xnor U25500 (N_25500,N_24608,N_24884);
nor U25501 (N_25501,N_25065,N_24695);
or U25502 (N_25502,N_24655,N_24955);
nor U25503 (N_25503,N_25124,N_24626);
nor U25504 (N_25504,N_24745,N_25180);
nor U25505 (N_25505,N_25193,N_24974);
nor U25506 (N_25506,N_24921,N_24842);
xor U25507 (N_25507,N_24762,N_24791);
xnor U25508 (N_25508,N_24905,N_24780);
xor U25509 (N_25509,N_25042,N_24922);
nand U25510 (N_25510,N_24862,N_25191);
xor U25511 (N_25511,N_24654,N_24835);
or U25512 (N_25512,N_24600,N_24818);
or U25513 (N_25513,N_25145,N_25153);
and U25514 (N_25514,N_24798,N_24899);
nand U25515 (N_25515,N_24915,N_24982);
nand U25516 (N_25516,N_24968,N_24650);
and U25517 (N_25517,N_24704,N_24999);
nand U25518 (N_25518,N_25131,N_24927);
or U25519 (N_25519,N_24733,N_25006);
xnor U25520 (N_25520,N_24665,N_24743);
xnor U25521 (N_25521,N_24940,N_24972);
or U25522 (N_25522,N_24883,N_24814);
or U25523 (N_25523,N_25007,N_24678);
and U25524 (N_25524,N_24868,N_25045);
nand U25525 (N_25525,N_25125,N_24817);
xnor U25526 (N_25526,N_24786,N_24995);
or U25527 (N_25527,N_24736,N_25068);
nand U25528 (N_25528,N_25154,N_24687);
and U25529 (N_25529,N_24686,N_24773);
or U25530 (N_25530,N_25199,N_25049);
nor U25531 (N_25531,N_24654,N_24875);
nand U25532 (N_25532,N_24991,N_24861);
and U25533 (N_25533,N_24680,N_24810);
nor U25534 (N_25534,N_24969,N_25146);
nand U25535 (N_25535,N_24718,N_24659);
xnor U25536 (N_25536,N_24758,N_24784);
and U25537 (N_25537,N_24741,N_24925);
nor U25538 (N_25538,N_24636,N_25183);
or U25539 (N_25539,N_24683,N_24680);
nand U25540 (N_25540,N_24702,N_24646);
and U25541 (N_25541,N_25143,N_24611);
xor U25542 (N_25542,N_24720,N_25003);
or U25543 (N_25543,N_24984,N_25006);
or U25544 (N_25544,N_24785,N_24682);
and U25545 (N_25545,N_25034,N_24652);
and U25546 (N_25546,N_24829,N_24616);
nor U25547 (N_25547,N_25064,N_24867);
nor U25548 (N_25548,N_24901,N_25064);
xnor U25549 (N_25549,N_24880,N_25070);
nor U25550 (N_25550,N_24930,N_24858);
and U25551 (N_25551,N_24906,N_25187);
or U25552 (N_25552,N_24951,N_24955);
and U25553 (N_25553,N_24759,N_24978);
xnor U25554 (N_25554,N_25047,N_24753);
and U25555 (N_25555,N_25016,N_24794);
nor U25556 (N_25556,N_24644,N_24669);
and U25557 (N_25557,N_24978,N_24896);
xnor U25558 (N_25558,N_25035,N_25164);
xor U25559 (N_25559,N_24908,N_24763);
nand U25560 (N_25560,N_24710,N_25165);
or U25561 (N_25561,N_24854,N_24820);
or U25562 (N_25562,N_25031,N_25164);
or U25563 (N_25563,N_25106,N_24868);
nand U25564 (N_25564,N_24714,N_25180);
xor U25565 (N_25565,N_24980,N_24935);
nor U25566 (N_25566,N_24896,N_24805);
nand U25567 (N_25567,N_24880,N_25150);
and U25568 (N_25568,N_24794,N_25034);
nor U25569 (N_25569,N_25149,N_24618);
and U25570 (N_25570,N_24871,N_24912);
nand U25571 (N_25571,N_25083,N_24680);
xnor U25572 (N_25572,N_24631,N_25152);
and U25573 (N_25573,N_25152,N_24944);
nor U25574 (N_25574,N_24930,N_24920);
nor U25575 (N_25575,N_25170,N_24845);
nor U25576 (N_25576,N_25039,N_24757);
nand U25577 (N_25577,N_24831,N_24878);
nor U25578 (N_25578,N_24618,N_24838);
nor U25579 (N_25579,N_24663,N_24784);
xnor U25580 (N_25580,N_24843,N_25142);
nor U25581 (N_25581,N_24657,N_24959);
xor U25582 (N_25582,N_24965,N_24636);
nor U25583 (N_25583,N_24742,N_24778);
and U25584 (N_25584,N_24852,N_25032);
xor U25585 (N_25585,N_25032,N_24961);
nand U25586 (N_25586,N_24979,N_25021);
or U25587 (N_25587,N_24648,N_25010);
and U25588 (N_25588,N_25026,N_24792);
nor U25589 (N_25589,N_25107,N_25074);
nor U25590 (N_25590,N_24977,N_25038);
nor U25591 (N_25591,N_24865,N_24639);
or U25592 (N_25592,N_24951,N_24717);
and U25593 (N_25593,N_24618,N_25041);
xor U25594 (N_25594,N_24904,N_24971);
nand U25595 (N_25595,N_24706,N_25181);
nor U25596 (N_25596,N_25179,N_25102);
or U25597 (N_25597,N_24733,N_24695);
nor U25598 (N_25598,N_25188,N_24673);
xnor U25599 (N_25599,N_24820,N_24617);
nand U25600 (N_25600,N_24631,N_24702);
nor U25601 (N_25601,N_24989,N_24882);
nand U25602 (N_25602,N_24889,N_24865);
and U25603 (N_25603,N_24677,N_24976);
nor U25604 (N_25604,N_25060,N_25150);
or U25605 (N_25605,N_24946,N_24744);
nor U25606 (N_25606,N_25121,N_24751);
nand U25607 (N_25607,N_25092,N_24862);
or U25608 (N_25608,N_25100,N_25059);
or U25609 (N_25609,N_24960,N_24643);
and U25610 (N_25610,N_24907,N_25064);
or U25611 (N_25611,N_24676,N_25184);
nor U25612 (N_25612,N_24898,N_24600);
nand U25613 (N_25613,N_24991,N_24792);
nor U25614 (N_25614,N_25186,N_24726);
nor U25615 (N_25615,N_25080,N_24709);
nor U25616 (N_25616,N_25002,N_24873);
xnor U25617 (N_25617,N_25052,N_24668);
xnor U25618 (N_25618,N_25034,N_24765);
xor U25619 (N_25619,N_25095,N_24882);
xnor U25620 (N_25620,N_24771,N_24765);
and U25621 (N_25621,N_24837,N_24908);
or U25622 (N_25622,N_25039,N_25173);
xor U25623 (N_25623,N_24744,N_25096);
and U25624 (N_25624,N_25009,N_24748);
nor U25625 (N_25625,N_24948,N_24750);
xor U25626 (N_25626,N_25021,N_24996);
nand U25627 (N_25627,N_24750,N_25091);
nand U25628 (N_25628,N_25154,N_24647);
nor U25629 (N_25629,N_25030,N_24795);
and U25630 (N_25630,N_25057,N_24863);
or U25631 (N_25631,N_25036,N_24734);
or U25632 (N_25632,N_24633,N_24995);
xor U25633 (N_25633,N_25145,N_24943);
nand U25634 (N_25634,N_24648,N_24848);
nand U25635 (N_25635,N_24745,N_24699);
nand U25636 (N_25636,N_24623,N_25002);
nand U25637 (N_25637,N_25024,N_24831);
nand U25638 (N_25638,N_24785,N_24614);
nor U25639 (N_25639,N_25103,N_25030);
nor U25640 (N_25640,N_24963,N_25147);
nand U25641 (N_25641,N_25043,N_24783);
nor U25642 (N_25642,N_24880,N_25176);
nand U25643 (N_25643,N_24672,N_24725);
xor U25644 (N_25644,N_25120,N_25091);
xor U25645 (N_25645,N_25149,N_24723);
or U25646 (N_25646,N_24804,N_24808);
nand U25647 (N_25647,N_24893,N_24710);
nor U25648 (N_25648,N_24693,N_25166);
nor U25649 (N_25649,N_25072,N_24654);
nand U25650 (N_25650,N_25085,N_24766);
nor U25651 (N_25651,N_24722,N_25001);
or U25652 (N_25652,N_24982,N_24816);
and U25653 (N_25653,N_24837,N_24612);
nand U25654 (N_25654,N_24960,N_25185);
or U25655 (N_25655,N_24865,N_24840);
nand U25656 (N_25656,N_25113,N_24953);
nand U25657 (N_25657,N_24944,N_24870);
xnor U25658 (N_25658,N_25042,N_24695);
xnor U25659 (N_25659,N_25072,N_24628);
nor U25660 (N_25660,N_25176,N_24950);
and U25661 (N_25661,N_25093,N_25062);
nor U25662 (N_25662,N_24862,N_24982);
nand U25663 (N_25663,N_24960,N_24890);
nor U25664 (N_25664,N_24668,N_24633);
xor U25665 (N_25665,N_25172,N_25126);
xor U25666 (N_25666,N_25116,N_24984);
nand U25667 (N_25667,N_24815,N_25037);
nor U25668 (N_25668,N_24935,N_25101);
and U25669 (N_25669,N_24858,N_24696);
nand U25670 (N_25670,N_24837,N_25040);
nand U25671 (N_25671,N_24979,N_24724);
nor U25672 (N_25672,N_25046,N_25168);
xnor U25673 (N_25673,N_25138,N_24639);
nor U25674 (N_25674,N_25115,N_25112);
or U25675 (N_25675,N_24899,N_24690);
nor U25676 (N_25676,N_24748,N_24621);
and U25677 (N_25677,N_25055,N_24611);
or U25678 (N_25678,N_24701,N_25160);
and U25679 (N_25679,N_25159,N_24861);
and U25680 (N_25680,N_24874,N_25177);
xor U25681 (N_25681,N_24619,N_24613);
nor U25682 (N_25682,N_24957,N_25173);
and U25683 (N_25683,N_24832,N_24791);
or U25684 (N_25684,N_24938,N_24871);
nor U25685 (N_25685,N_25105,N_24879);
nor U25686 (N_25686,N_24792,N_24770);
and U25687 (N_25687,N_24681,N_25185);
or U25688 (N_25688,N_24695,N_25142);
xor U25689 (N_25689,N_24836,N_24735);
and U25690 (N_25690,N_24922,N_24909);
nor U25691 (N_25691,N_24780,N_24936);
or U25692 (N_25692,N_24899,N_24734);
xnor U25693 (N_25693,N_24917,N_24678);
nor U25694 (N_25694,N_24862,N_25159);
xnor U25695 (N_25695,N_25170,N_24839);
and U25696 (N_25696,N_25094,N_24816);
nor U25697 (N_25697,N_24846,N_25140);
or U25698 (N_25698,N_24963,N_24999);
xor U25699 (N_25699,N_24920,N_24735);
nor U25700 (N_25700,N_24938,N_25018);
nand U25701 (N_25701,N_24611,N_25174);
and U25702 (N_25702,N_25009,N_24986);
xnor U25703 (N_25703,N_25160,N_25168);
xor U25704 (N_25704,N_24662,N_24659);
or U25705 (N_25705,N_24975,N_25116);
xor U25706 (N_25706,N_25081,N_24871);
nor U25707 (N_25707,N_25123,N_25076);
or U25708 (N_25708,N_25039,N_24960);
nand U25709 (N_25709,N_24887,N_24831);
nand U25710 (N_25710,N_25168,N_25107);
nand U25711 (N_25711,N_25078,N_24730);
and U25712 (N_25712,N_25004,N_24763);
xnor U25713 (N_25713,N_25155,N_25059);
or U25714 (N_25714,N_24702,N_24744);
nand U25715 (N_25715,N_24946,N_24950);
nor U25716 (N_25716,N_24815,N_24980);
and U25717 (N_25717,N_24828,N_25087);
nor U25718 (N_25718,N_24781,N_24807);
nor U25719 (N_25719,N_24805,N_24648);
and U25720 (N_25720,N_25160,N_25186);
nand U25721 (N_25721,N_24788,N_24944);
nand U25722 (N_25722,N_24859,N_25166);
and U25723 (N_25723,N_24848,N_24898);
nor U25724 (N_25724,N_24798,N_25133);
or U25725 (N_25725,N_25104,N_24983);
nand U25726 (N_25726,N_24606,N_24770);
nand U25727 (N_25727,N_24757,N_24707);
xnor U25728 (N_25728,N_24672,N_25061);
or U25729 (N_25729,N_24775,N_24828);
or U25730 (N_25730,N_24711,N_24888);
nor U25731 (N_25731,N_25002,N_25107);
xor U25732 (N_25732,N_25024,N_24840);
and U25733 (N_25733,N_24634,N_25125);
or U25734 (N_25734,N_24913,N_25039);
nor U25735 (N_25735,N_24620,N_24994);
nand U25736 (N_25736,N_24866,N_24613);
xor U25737 (N_25737,N_24613,N_25039);
xnor U25738 (N_25738,N_24815,N_24632);
nand U25739 (N_25739,N_24648,N_24975);
nand U25740 (N_25740,N_25161,N_24990);
nor U25741 (N_25741,N_24987,N_24838);
xnor U25742 (N_25742,N_25144,N_25181);
or U25743 (N_25743,N_25002,N_25141);
nor U25744 (N_25744,N_25129,N_25127);
and U25745 (N_25745,N_24750,N_24762);
nor U25746 (N_25746,N_24795,N_25079);
nor U25747 (N_25747,N_24989,N_24951);
or U25748 (N_25748,N_25045,N_24670);
nor U25749 (N_25749,N_24635,N_24611);
and U25750 (N_25750,N_24965,N_24664);
xnor U25751 (N_25751,N_24755,N_24825);
and U25752 (N_25752,N_24657,N_25002);
or U25753 (N_25753,N_24694,N_25156);
xor U25754 (N_25754,N_24722,N_25151);
or U25755 (N_25755,N_24970,N_25038);
nand U25756 (N_25756,N_24714,N_24791);
xnor U25757 (N_25757,N_24751,N_24884);
or U25758 (N_25758,N_25102,N_24787);
xor U25759 (N_25759,N_24787,N_25168);
xor U25760 (N_25760,N_24689,N_25164);
or U25761 (N_25761,N_25146,N_24788);
or U25762 (N_25762,N_24684,N_25109);
and U25763 (N_25763,N_25146,N_25042);
nor U25764 (N_25764,N_24631,N_25157);
or U25765 (N_25765,N_24724,N_25145);
nand U25766 (N_25766,N_24965,N_25050);
nor U25767 (N_25767,N_24830,N_24713);
xnor U25768 (N_25768,N_24790,N_25059);
xnor U25769 (N_25769,N_24971,N_24988);
and U25770 (N_25770,N_24879,N_25147);
or U25771 (N_25771,N_24891,N_24853);
nand U25772 (N_25772,N_24770,N_24796);
nor U25773 (N_25773,N_24894,N_25173);
and U25774 (N_25774,N_24991,N_24934);
nor U25775 (N_25775,N_25128,N_24847);
or U25776 (N_25776,N_24934,N_25026);
xor U25777 (N_25777,N_24755,N_24946);
or U25778 (N_25778,N_24840,N_24890);
or U25779 (N_25779,N_24751,N_24827);
nand U25780 (N_25780,N_24956,N_24633);
or U25781 (N_25781,N_24808,N_24647);
xnor U25782 (N_25782,N_25189,N_24916);
xor U25783 (N_25783,N_25147,N_24842);
nand U25784 (N_25784,N_24610,N_24917);
and U25785 (N_25785,N_24661,N_24950);
xnor U25786 (N_25786,N_25003,N_24824);
or U25787 (N_25787,N_24949,N_24762);
nand U25788 (N_25788,N_24698,N_24953);
and U25789 (N_25789,N_25086,N_24909);
xnor U25790 (N_25790,N_24711,N_24724);
and U25791 (N_25791,N_24616,N_24609);
or U25792 (N_25792,N_24807,N_24916);
nand U25793 (N_25793,N_24931,N_24648);
and U25794 (N_25794,N_24769,N_25019);
nor U25795 (N_25795,N_24780,N_24887);
xnor U25796 (N_25796,N_25012,N_25198);
and U25797 (N_25797,N_24624,N_25170);
or U25798 (N_25798,N_24715,N_24750);
or U25799 (N_25799,N_24987,N_25145);
nand U25800 (N_25800,N_25408,N_25401);
nor U25801 (N_25801,N_25773,N_25209);
or U25802 (N_25802,N_25200,N_25521);
xor U25803 (N_25803,N_25469,N_25792);
nand U25804 (N_25804,N_25686,N_25749);
and U25805 (N_25805,N_25238,N_25623);
nor U25806 (N_25806,N_25246,N_25205);
xor U25807 (N_25807,N_25433,N_25418);
or U25808 (N_25808,N_25705,N_25780);
nand U25809 (N_25809,N_25625,N_25414);
xnor U25810 (N_25810,N_25606,N_25510);
nor U25811 (N_25811,N_25384,N_25497);
nand U25812 (N_25812,N_25612,N_25277);
and U25813 (N_25813,N_25797,N_25397);
nor U25814 (N_25814,N_25770,N_25366);
or U25815 (N_25815,N_25380,N_25585);
and U25816 (N_25816,N_25581,N_25647);
and U25817 (N_25817,N_25755,N_25421);
or U25818 (N_25818,N_25786,N_25640);
nor U25819 (N_25819,N_25642,N_25412);
and U25820 (N_25820,N_25717,N_25697);
and U25821 (N_25821,N_25610,N_25300);
xor U25822 (N_25822,N_25374,N_25458);
xnor U25823 (N_25823,N_25325,N_25646);
nor U25824 (N_25824,N_25701,N_25628);
and U25825 (N_25825,N_25688,N_25724);
and U25826 (N_25826,N_25662,N_25315);
or U25827 (N_25827,N_25594,N_25314);
xor U25828 (N_25828,N_25626,N_25472);
xor U25829 (N_25829,N_25290,N_25482);
and U25830 (N_25830,N_25243,N_25535);
nand U25831 (N_25831,N_25547,N_25536);
nand U25832 (N_25832,N_25379,N_25709);
nand U25833 (N_25833,N_25228,N_25293);
nand U25834 (N_25834,N_25789,N_25618);
nor U25835 (N_25835,N_25227,N_25583);
nor U25836 (N_25836,N_25526,N_25236);
nand U25837 (N_25837,N_25367,N_25377);
xor U25838 (N_25838,N_25253,N_25653);
xor U25839 (N_25839,N_25465,N_25604);
nor U25840 (N_25840,N_25648,N_25307);
and U25841 (N_25841,N_25217,N_25423);
nor U25842 (N_25842,N_25250,N_25344);
xor U25843 (N_25843,N_25760,N_25339);
xor U25844 (N_25844,N_25321,N_25263);
or U25845 (N_25845,N_25406,N_25534);
nor U25846 (N_25846,N_25475,N_25434);
nor U25847 (N_25847,N_25793,N_25566);
and U25848 (N_25848,N_25447,N_25663);
or U25849 (N_25849,N_25771,N_25448);
and U25850 (N_25850,N_25638,N_25726);
nor U25851 (N_25851,N_25256,N_25511);
and U25852 (N_25852,N_25621,N_25545);
nand U25853 (N_25853,N_25260,N_25282);
or U25854 (N_25854,N_25525,N_25455);
and U25855 (N_25855,N_25540,N_25287);
xor U25856 (N_25856,N_25629,N_25453);
xnor U25857 (N_25857,N_25788,N_25441);
and U25858 (N_25858,N_25439,N_25716);
and U25859 (N_25859,N_25201,N_25775);
nand U25860 (N_25860,N_25303,N_25267);
and U25861 (N_25861,N_25301,N_25283);
and U25862 (N_25862,N_25722,N_25495);
xor U25863 (N_25863,N_25393,N_25635);
nand U25864 (N_25864,N_25590,N_25402);
and U25865 (N_25865,N_25241,N_25302);
nor U25866 (N_25866,N_25332,N_25729);
nor U25867 (N_25867,N_25313,N_25644);
xor U25868 (N_25868,N_25661,N_25557);
and U25869 (N_25869,N_25349,N_25262);
xnor U25870 (N_25870,N_25387,N_25669);
nand U25871 (N_25871,N_25711,N_25440);
and U25872 (N_25872,N_25504,N_25291);
nor U25873 (N_25873,N_25474,N_25312);
nand U25874 (N_25874,N_25296,N_25257);
xor U25875 (N_25875,N_25350,N_25231);
nor U25876 (N_25876,N_25477,N_25326);
and U25877 (N_25877,N_25405,N_25533);
nor U25878 (N_25878,N_25672,N_25278);
xnor U25879 (N_25879,N_25654,N_25490);
nand U25880 (N_25880,N_25316,N_25764);
nand U25881 (N_25881,N_25436,N_25643);
nand U25882 (N_25882,N_25608,N_25299);
and U25883 (N_25883,N_25216,N_25233);
or U25884 (N_25884,N_25487,N_25754);
nand U25885 (N_25885,N_25211,N_25356);
and U25886 (N_25886,N_25322,N_25294);
nand U25887 (N_25887,N_25410,N_25342);
xnor U25888 (N_25888,N_25273,N_25558);
nand U25889 (N_25889,N_25288,N_25551);
nor U25890 (N_25890,N_25703,N_25503);
xnor U25891 (N_25891,N_25693,N_25435);
nand U25892 (N_25892,N_25687,N_25328);
nor U25893 (N_25893,N_25550,N_25685);
xor U25894 (N_25894,N_25343,N_25753);
nand U25895 (N_25895,N_25578,N_25645);
or U25896 (N_25896,N_25799,N_25275);
nand U25897 (N_25897,N_25665,N_25268);
nor U25898 (N_25898,N_25620,N_25427);
or U25899 (N_25899,N_25784,N_25376);
xnor U25900 (N_25900,N_25781,N_25471);
nor U25901 (N_25901,N_25403,N_25779);
and U25902 (N_25902,N_25420,N_25619);
xnor U25903 (N_25903,N_25554,N_25763);
xnor U25904 (N_25904,N_25428,N_25776);
or U25905 (N_25905,N_25708,N_25532);
nor U25906 (N_25906,N_25598,N_25787);
and U25907 (N_25907,N_25244,N_25668);
nand U25908 (N_25908,N_25508,N_25212);
and U25909 (N_25909,N_25602,N_25768);
xnor U25910 (N_25910,N_25655,N_25354);
nand U25911 (N_25911,N_25580,N_25348);
nor U25912 (N_25912,N_25422,N_25255);
nand U25913 (N_25913,N_25750,N_25398);
nand U25914 (N_25914,N_25746,N_25235);
and U25915 (N_25915,N_25530,N_25695);
or U25916 (N_25916,N_25735,N_25264);
and U25917 (N_25917,N_25527,N_25446);
and U25918 (N_25918,N_25591,N_25476);
nor U25919 (N_25919,N_25457,N_25549);
nand U25920 (N_25920,N_25215,N_25395);
nor U25921 (N_25921,N_25631,N_25794);
nand U25922 (N_25922,N_25528,N_25486);
nor U25923 (N_25923,N_25737,N_25564);
or U25924 (N_25924,N_25700,N_25470);
xnor U25925 (N_25925,N_25556,N_25637);
nor U25926 (N_25926,N_25353,N_25603);
and U25927 (N_25927,N_25432,N_25286);
or U25928 (N_25928,N_25514,N_25285);
nand U25929 (N_25929,N_25727,N_25203);
nor U25930 (N_25930,N_25666,N_25281);
nand U25931 (N_25931,N_25759,N_25577);
and U25932 (N_25932,N_25237,N_25515);
and U25933 (N_25933,N_25505,N_25372);
and U25934 (N_25934,N_25736,N_25468);
or U25935 (N_25935,N_25289,N_25667);
nor U25936 (N_25936,N_25502,N_25245);
or U25937 (N_25937,N_25396,N_25559);
nand U25938 (N_25938,N_25553,N_25785);
xor U25939 (N_25939,N_25740,N_25338);
and U25940 (N_25940,N_25388,N_25451);
and U25941 (N_25941,N_25459,N_25499);
xnor U25942 (N_25942,N_25323,N_25224);
and U25943 (N_25943,N_25587,N_25728);
or U25944 (N_25944,N_25333,N_25251);
and U25945 (N_25945,N_25383,N_25284);
nand U25946 (N_25946,N_25649,N_25745);
nand U25947 (N_25947,N_25225,N_25513);
or U25948 (N_25948,N_25493,N_25713);
xnor U25949 (N_25949,N_25769,N_25498);
xor U25950 (N_25950,N_25444,N_25632);
nor U25951 (N_25951,N_25607,N_25630);
xor U25952 (N_25952,N_25543,N_25531);
xnor U25953 (N_25953,N_25699,N_25778);
nor U25954 (N_25954,N_25341,N_25673);
nand U25955 (N_25955,N_25491,N_25450);
xnor U25956 (N_25956,N_25568,N_25596);
xnor U25957 (N_25957,N_25707,N_25651);
nand U25958 (N_25958,N_25617,N_25572);
xnor U25959 (N_25959,N_25270,N_25674);
and U25960 (N_25960,N_25798,N_25473);
and U25961 (N_25961,N_25202,N_25742);
or U25962 (N_25962,N_25624,N_25570);
xnor U25963 (N_25963,N_25324,N_25478);
or U25964 (N_25964,N_25239,N_25252);
xnor U25965 (N_25965,N_25795,N_25274);
nand U25966 (N_25966,N_25271,N_25466);
nor U25967 (N_25967,N_25467,N_25219);
nand U25968 (N_25968,N_25691,N_25417);
nand U25969 (N_25969,N_25519,N_25364);
and U25970 (N_25970,N_25494,N_25351);
xor U25971 (N_25971,N_25518,N_25306);
nor U25972 (N_25972,N_25352,N_25744);
nand U25973 (N_25973,N_25445,N_25452);
or U25974 (N_25974,N_25357,N_25415);
nor U25975 (N_25975,N_25331,N_25681);
or U25976 (N_25976,N_25438,N_25579);
or U25977 (N_25977,N_25600,N_25454);
or U25978 (N_25978,N_25391,N_25548);
nand U25979 (N_25979,N_25652,N_25346);
nor U25980 (N_25980,N_25777,N_25774);
xor U25981 (N_25981,N_25258,N_25766);
nor U25982 (N_25982,N_25360,N_25517);
and U25983 (N_25983,N_25539,N_25714);
nand U25984 (N_25984,N_25622,N_25659);
xor U25985 (N_25985,N_25247,N_25751);
or U25986 (N_25986,N_25743,N_25463);
nor U25987 (N_25987,N_25680,N_25409);
or U25988 (N_25988,N_25425,N_25242);
nor U25989 (N_25989,N_25639,N_25501);
nor U25990 (N_25990,N_25689,N_25589);
xor U25991 (N_25991,N_25230,N_25298);
and U25992 (N_25992,N_25456,N_25611);
nor U25993 (N_25993,N_25259,N_25741);
or U25994 (N_25994,N_25232,N_25492);
or U25995 (N_25995,N_25758,N_25330);
or U25996 (N_25996,N_25650,N_25748);
nand U25997 (N_25997,N_25392,N_25292);
or U25998 (N_25998,N_25615,N_25730);
nor U25999 (N_25999,N_25368,N_25222);
or U26000 (N_26000,N_25783,N_25756);
or U26001 (N_26001,N_25679,N_25555);
xor U26002 (N_26002,N_25279,N_25381);
xor U26003 (N_26003,N_25683,N_25449);
xor U26004 (N_26004,N_25520,N_25221);
or U26005 (N_26005,N_25407,N_25682);
and U26006 (N_26006,N_25584,N_25461);
and U26007 (N_26007,N_25204,N_25529);
or U26008 (N_26008,N_25399,N_25522);
nand U26009 (N_26009,N_25223,N_25336);
nand U26010 (N_26010,N_25375,N_25226);
or U26011 (N_26011,N_25280,N_25507);
xor U26012 (N_26012,N_25369,N_25370);
nand U26013 (N_26013,N_25214,N_25569);
or U26014 (N_26014,N_25460,N_25721);
nand U26015 (N_26015,N_25462,N_25419);
nand U26016 (N_26016,N_25340,N_25389);
nor U26017 (N_26017,N_25442,N_25582);
and U26018 (N_26018,N_25254,N_25706);
xor U26019 (N_26019,N_25481,N_25576);
nand U26020 (N_26020,N_25480,N_25248);
xnor U26021 (N_26021,N_25429,N_25677);
and U26022 (N_26022,N_25361,N_25309);
nand U26023 (N_26023,N_25329,N_25712);
and U26024 (N_26024,N_25304,N_25586);
or U26025 (N_26025,N_25404,N_25641);
xnor U26026 (N_26026,N_25249,N_25319);
or U26027 (N_26027,N_25765,N_25544);
or U26028 (N_26028,N_25295,N_25413);
nor U26029 (N_26029,N_25240,N_25390);
xor U26030 (N_26030,N_25269,N_25208);
nand U26031 (N_26031,N_25593,N_25430);
xor U26032 (N_26032,N_25464,N_25739);
nand U26033 (N_26033,N_25762,N_25334);
or U26034 (N_26034,N_25738,N_25400);
nor U26035 (N_26035,N_25373,N_25297);
and U26036 (N_26036,N_25546,N_25443);
nand U26037 (N_26037,N_25561,N_25335);
and U26038 (N_26038,N_25565,N_25605);
nor U26039 (N_26039,N_25715,N_25720);
nor U26040 (N_26040,N_25347,N_25318);
xor U26041 (N_26041,N_25772,N_25571);
and U26042 (N_26042,N_25305,N_25371);
nand U26043 (N_26043,N_25218,N_25506);
and U26044 (N_26044,N_25675,N_25266);
or U26045 (N_26045,N_25563,N_25660);
and U26046 (N_26046,N_25614,N_25485);
and U26047 (N_26047,N_25320,N_25310);
and U26048 (N_26048,N_25698,N_25424);
nor U26049 (N_26049,N_25378,N_25311);
or U26050 (N_26050,N_25437,N_25734);
xnor U26051 (N_26051,N_25358,N_25394);
nor U26052 (N_26052,N_25489,N_25692);
and U26053 (N_26053,N_25541,N_25678);
or U26054 (N_26054,N_25592,N_25595);
nor U26055 (N_26055,N_25575,N_25732);
nor U26056 (N_26056,N_25702,N_25609);
nor U26057 (N_26057,N_25516,N_25671);
or U26058 (N_26058,N_25796,N_25704);
or U26059 (N_26059,N_25213,N_25791);
xnor U26060 (N_26060,N_25597,N_25317);
nand U26061 (N_26061,N_25723,N_25483);
nor U26062 (N_26062,N_25601,N_25337);
and U26063 (N_26063,N_25757,N_25731);
nor U26064 (N_26064,N_25411,N_25588);
nand U26065 (N_26065,N_25613,N_25627);
nor U26066 (N_26066,N_25365,N_25509);
xnor U26067 (N_26067,N_25599,N_25426);
or U26068 (N_26068,N_25633,N_25496);
and U26069 (N_26069,N_25500,N_25386);
nand U26070 (N_26070,N_25676,N_25210);
nand U26071 (N_26071,N_25719,N_25694);
nor U26072 (N_26072,N_25790,N_25634);
and U26073 (N_26073,N_25363,N_25567);
xor U26074 (N_26074,N_25234,N_25573);
nor U26075 (N_26075,N_25560,N_25479);
or U26076 (N_26076,N_25537,N_25276);
and U26077 (N_26077,N_25690,N_25636);
xnor U26078 (N_26078,N_25265,N_25562);
nand U26079 (N_26079,N_25761,N_25752);
or U26080 (N_26080,N_25207,N_25220);
nor U26081 (N_26081,N_25261,N_25523);
xor U26082 (N_26082,N_25385,N_25538);
xor U26083 (N_26083,N_25710,N_25552);
or U26084 (N_26084,N_25345,N_25229);
xnor U26085 (N_26085,N_25658,N_25382);
xor U26086 (N_26086,N_25488,N_25670);
nor U26087 (N_26087,N_25327,N_25574);
or U26088 (N_26088,N_25747,N_25512);
or U26089 (N_26089,N_25362,N_25416);
nor U26090 (N_26090,N_25206,N_25733);
and U26091 (N_26091,N_25782,N_25542);
or U26092 (N_26092,N_25272,N_25684);
and U26093 (N_26093,N_25725,N_25524);
and U26094 (N_26094,N_25656,N_25355);
xnor U26095 (N_26095,N_25718,N_25308);
nand U26096 (N_26096,N_25696,N_25359);
xor U26097 (N_26097,N_25767,N_25616);
xor U26098 (N_26098,N_25664,N_25657);
nor U26099 (N_26099,N_25431,N_25484);
and U26100 (N_26100,N_25291,N_25217);
xnor U26101 (N_26101,N_25705,N_25202);
xnor U26102 (N_26102,N_25293,N_25586);
nand U26103 (N_26103,N_25751,N_25249);
or U26104 (N_26104,N_25449,N_25572);
or U26105 (N_26105,N_25268,N_25569);
nand U26106 (N_26106,N_25526,N_25237);
xor U26107 (N_26107,N_25727,N_25376);
nand U26108 (N_26108,N_25550,N_25610);
nand U26109 (N_26109,N_25732,N_25632);
xnor U26110 (N_26110,N_25673,N_25664);
xor U26111 (N_26111,N_25681,N_25292);
and U26112 (N_26112,N_25404,N_25352);
and U26113 (N_26113,N_25248,N_25518);
nor U26114 (N_26114,N_25628,N_25394);
nand U26115 (N_26115,N_25230,N_25563);
or U26116 (N_26116,N_25270,N_25699);
or U26117 (N_26117,N_25705,N_25769);
or U26118 (N_26118,N_25316,N_25660);
nand U26119 (N_26119,N_25716,N_25357);
or U26120 (N_26120,N_25322,N_25670);
and U26121 (N_26121,N_25591,N_25601);
xor U26122 (N_26122,N_25729,N_25611);
xor U26123 (N_26123,N_25505,N_25405);
xor U26124 (N_26124,N_25789,N_25274);
xor U26125 (N_26125,N_25699,N_25456);
and U26126 (N_26126,N_25766,N_25266);
nor U26127 (N_26127,N_25444,N_25501);
or U26128 (N_26128,N_25473,N_25531);
and U26129 (N_26129,N_25236,N_25506);
xor U26130 (N_26130,N_25686,N_25415);
and U26131 (N_26131,N_25700,N_25517);
or U26132 (N_26132,N_25269,N_25550);
nand U26133 (N_26133,N_25357,N_25313);
and U26134 (N_26134,N_25544,N_25240);
or U26135 (N_26135,N_25646,N_25213);
xnor U26136 (N_26136,N_25740,N_25425);
or U26137 (N_26137,N_25464,N_25339);
nand U26138 (N_26138,N_25488,N_25433);
xor U26139 (N_26139,N_25574,N_25325);
nand U26140 (N_26140,N_25204,N_25657);
xor U26141 (N_26141,N_25484,N_25289);
nand U26142 (N_26142,N_25269,N_25280);
and U26143 (N_26143,N_25361,N_25494);
nor U26144 (N_26144,N_25279,N_25697);
or U26145 (N_26145,N_25709,N_25468);
nand U26146 (N_26146,N_25565,N_25625);
xnor U26147 (N_26147,N_25567,N_25552);
or U26148 (N_26148,N_25277,N_25311);
xnor U26149 (N_26149,N_25742,N_25297);
or U26150 (N_26150,N_25763,N_25624);
and U26151 (N_26151,N_25434,N_25441);
and U26152 (N_26152,N_25623,N_25316);
and U26153 (N_26153,N_25563,N_25527);
xor U26154 (N_26154,N_25234,N_25777);
and U26155 (N_26155,N_25464,N_25462);
nor U26156 (N_26156,N_25619,N_25692);
or U26157 (N_26157,N_25740,N_25205);
nand U26158 (N_26158,N_25309,N_25285);
and U26159 (N_26159,N_25300,N_25771);
and U26160 (N_26160,N_25759,N_25565);
xnor U26161 (N_26161,N_25420,N_25371);
xnor U26162 (N_26162,N_25587,N_25378);
and U26163 (N_26163,N_25260,N_25479);
nor U26164 (N_26164,N_25434,N_25523);
and U26165 (N_26165,N_25474,N_25621);
or U26166 (N_26166,N_25453,N_25201);
or U26167 (N_26167,N_25678,N_25606);
nor U26168 (N_26168,N_25690,N_25477);
nor U26169 (N_26169,N_25783,N_25342);
nand U26170 (N_26170,N_25551,N_25594);
nand U26171 (N_26171,N_25703,N_25607);
nor U26172 (N_26172,N_25744,N_25639);
nand U26173 (N_26173,N_25437,N_25273);
nand U26174 (N_26174,N_25450,N_25486);
nand U26175 (N_26175,N_25358,N_25312);
nor U26176 (N_26176,N_25609,N_25215);
nand U26177 (N_26177,N_25435,N_25702);
nand U26178 (N_26178,N_25239,N_25455);
nor U26179 (N_26179,N_25556,N_25737);
or U26180 (N_26180,N_25782,N_25363);
or U26181 (N_26181,N_25512,N_25261);
and U26182 (N_26182,N_25574,N_25577);
xor U26183 (N_26183,N_25264,N_25668);
nor U26184 (N_26184,N_25714,N_25296);
nor U26185 (N_26185,N_25697,N_25404);
xor U26186 (N_26186,N_25749,N_25668);
and U26187 (N_26187,N_25239,N_25550);
nand U26188 (N_26188,N_25338,N_25295);
or U26189 (N_26189,N_25421,N_25515);
or U26190 (N_26190,N_25779,N_25342);
or U26191 (N_26191,N_25389,N_25479);
and U26192 (N_26192,N_25577,N_25479);
xor U26193 (N_26193,N_25323,N_25423);
or U26194 (N_26194,N_25568,N_25215);
xnor U26195 (N_26195,N_25772,N_25298);
nor U26196 (N_26196,N_25217,N_25288);
or U26197 (N_26197,N_25412,N_25531);
nand U26198 (N_26198,N_25215,N_25295);
or U26199 (N_26199,N_25752,N_25348);
nor U26200 (N_26200,N_25766,N_25704);
nor U26201 (N_26201,N_25562,N_25788);
or U26202 (N_26202,N_25715,N_25605);
xnor U26203 (N_26203,N_25769,N_25720);
nand U26204 (N_26204,N_25774,N_25636);
nor U26205 (N_26205,N_25683,N_25325);
nand U26206 (N_26206,N_25781,N_25544);
nand U26207 (N_26207,N_25506,N_25728);
nor U26208 (N_26208,N_25644,N_25275);
and U26209 (N_26209,N_25671,N_25378);
nand U26210 (N_26210,N_25564,N_25219);
nor U26211 (N_26211,N_25744,N_25606);
nand U26212 (N_26212,N_25224,N_25509);
xor U26213 (N_26213,N_25695,N_25703);
xnor U26214 (N_26214,N_25251,N_25499);
nand U26215 (N_26215,N_25609,N_25370);
or U26216 (N_26216,N_25352,N_25359);
xnor U26217 (N_26217,N_25466,N_25702);
or U26218 (N_26218,N_25784,N_25706);
and U26219 (N_26219,N_25572,N_25342);
or U26220 (N_26220,N_25406,N_25670);
nor U26221 (N_26221,N_25750,N_25586);
nor U26222 (N_26222,N_25530,N_25429);
and U26223 (N_26223,N_25278,N_25640);
and U26224 (N_26224,N_25632,N_25404);
xnor U26225 (N_26225,N_25300,N_25590);
nand U26226 (N_26226,N_25267,N_25296);
and U26227 (N_26227,N_25710,N_25770);
and U26228 (N_26228,N_25596,N_25669);
or U26229 (N_26229,N_25387,N_25295);
xor U26230 (N_26230,N_25284,N_25573);
nor U26231 (N_26231,N_25474,N_25412);
nand U26232 (N_26232,N_25710,N_25413);
nand U26233 (N_26233,N_25433,N_25537);
xnor U26234 (N_26234,N_25295,N_25283);
nand U26235 (N_26235,N_25735,N_25562);
or U26236 (N_26236,N_25790,N_25410);
nor U26237 (N_26237,N_25212,N_25469);
or U26238 (N_26238,N_25360,N_25724);
and U26239 (N_26239,N_25738,N_25511);
nor U26240 (N_26240,N_25431,N_25608);
nor U26241 (N_26241,N_25799,N_25334);
nor U26242 (N_26242,N_25541,N_25398);
xor U26243 (N_26243,N_25254,N_25597);
nor U26244 (N_26244,N_25616,N_25746);
nand U26245 (N_26245,N_25585,N_25560);
and U26246 (N_26246,N_25289,N_25308);
xor U26247 (N_26247,N_25728,N_25579);
xnor U26248 (N_26248,N_25648,N_25689);
nor U26249 (N_26249,N_25568,N_25534);
xor U26250 (N_26250,N_25291,N_25299);
xnor U26251 (N_26251,N_25488,N_25340);
and U26252 (N_26252,N_25368,N_25434);
and U26253 (N_26253,N_25768,N_25609);
or U26254 (N_26254,N_25475,N_25561);
or U26255 (N_26255,N_25277,N_25675);
or U26256 (N_26256,N_25554,N_25585);
xor U26257 (N_26257,N_25709,N_25457);
nor U26258 (N_26258,N_25356,N_25387);
and U26259 (N_26259,N_25509,N_25729);
xnor U26260 (N_26260,N_25261,N_25458);
and U26261 (N_26261,N_25523,N_25654);
nor U26262 (N_26262,N_25602,N_25434);
or U26263 (N_26263,N_25365,N_25785);
nor U26264 (N_26264,N_25289,N_25314);
nor U26265 (N_26265,N_25745,N_25382);
nor U26266 (N_26266,N_25767,N_25415);
nor U26267 (N_26267,N_25650,N_25370);
nand U26268 (N_26268,N_25399,N_25202);
nand U26269 (N_26269,N_25452,N_25412);
and U26270 (N_26270,N_25253,N_25602);
nand U26271 (N_26271,N_25593,N_25738);
nand U26272 (N_26272,N_25259,N_25626);
nand U26273 (N_26273,N_25264,N_25675);
nor U26274 (N_26274,N_25408,N_25344);
or U26275 (N_26275,N_25786,N_25494);
xnor U26276 (N_26276,N_25475,N_25750);
nor U26277 (N_26277,N_25509,N_25626);
nor U26278 (N_26278,N_25354,N_25624);
and U26279 (N_26279,N_25273,N_25637);
nor U26280 (N_26280,N_25661,N_25384);
and U26281 (N_26281,N_25383,N_25766);
or U26282 (N_26282,N_25209,N_25455);
nor U26283 (N_26283,N_25524,N_25340);
xor U26284 (N_26284,N_25338,N_25780);
nor U26285 (N_26285,N_25247,N_25286);
nand U26286 (N_26286,N_25273,N_25485);
and U26287 (N_26287,N_25250,N_25634);
nor U26288 (N_26288,N_25285,N_25699);
nand U26289 (N_26289,N_25516,N_25296);
and U26290 (N_26290,N_25725,N_25734);
or U26291 (N_26291,N_25760,N_25464);
and U26292 (N_26292,N_25661,N_25649);
nand U26293 (N_26293,N_25746,N_25482);
nor U26294 (N_26294,N_25560,N_25733);
nor U26295 (N_26295,N_25747,N_25714);
nor U26296 (N_26296,N_25347,N_25647);
nor U26297 (N_26297,N_25269,N_25425);
nor U26298 (N_26298,N_25241,N_25476);
nand U26299 (N_26299,N_25680,N_25720);
nor U26300 (N_26300,N_25397,N_25252);
and U26301 (N_26301,N_25208,N_25261);
xnor U26302 (N_26302,N_25393,N_25520);
or U26303 (N_26303,N_25551,N_25470);
nor U26304 (N_26304,N_25793,N_25482);
nor U26305 (N_26305,N_25747,N_25347);
and U26306 (N_26306,N_25539,N_25675);
nor U26307 (N_26307,N_25650,N_25351);
xor U26308 (N_26308,N_25388,N_25352);
xnor U26309 (N_26309,N_25444,N_25344);
and U26310 (N_26310,N_25585,N_25455);
nand U26311 (N_26311,N_25741,N_25456);
and U26312 (N_26312,N_25740,N_25718);
xnor U26313 (N_26313,N_25723,N_25276);
or U26314 (N_26314,N_25654,N_25220);
xor U26315 (N_26315,N_25691,N_25589);
nand U26316 (N_26316,N_25273,N_25405);
xnor U26317 (N_26317,N_25697,N_25260);
xnor U26318 (N_26318,N_25726,N_25598);
or U26319 (N_26319,N_25240,N_25686);
or U26320 (N_26320,N_25355,N_25445);
and U26321 (N_26321,N_25752,N_25454);
nand U26322 (N_26322,N_25723,N_25411);
and U26323 (N_26323,N_25527,N_25247);
nand U26324 (N_26324,N_25402,N_25372);
xor U26325 (N_26325,N_25568,N_25527);
xnor U26326 (N_26326,N_25718,N_25219);
and U26327 (N_26327,N_25698,N_25211);
nand U26328 (N_26328,N_25341,N_25215);
xor U26329 (N_26329,N_25214,N_25387);
xnor U26330 (N_26330,N_25552,N_25682);
nor U26331 (N_26331,N_25536,N_25535);
nand U26332 (N_26332,N_25222,N_25674);
or U26333 (N_26333,N_25407,N_25517);
xnor U26334 (N_26334,N_25509,N_25363);
or U26335 (N_26335,N_25480,N_25675);
nand U26336 (N_26336,N_25740,N_25287);
nor U26337 (N_26337,N_25620,N_25378);
nand U26338 (N_26338,N_25500,N_25225);
nand U26339 (N_26339,N_25211,N_25324);
nand U26340 (N_26340,N_25243,N_25209);
nand U26341 (N_26341,N_25386,N_25433);
xor U26342 (N_26342,N_25747,N_25383);
or U26343 (N_26343,N_25629,N_25279);
nor U26344 (N_26344,N_25262,N_25641);
and U26345 (N_26345,N_25221,N_25380);
nor U26346 (N_26346,N_25285,N_25432);
or U26347 (N_26347,N_25360,N_25798);
or U26348 (N_26348,N_25740,N_25507);
or U26349 (N_26349,N_25335,N_25306);
or U26350 (N_26350,N_25423,N_25428);
and U26351 (N_26351,N_25390,N_25565);
nand U26352 (N_26352,N_25568,N_25210);
xnor U26353 (N_26353,N_25578,N_25276);
nand U26354 (N_26354,N_25426,N_25640);
nand U26355 (N_26355,N_25430,N_25713);
nor U26356 (N_26356,N_25765,N_25622);
and U26357 (N_26357,N_25686,N_25345);
nand U26358 (N_26358,N_25782,N_25511);
or U26359 (N_26359,N_25290,N_25210);
or U26360 (N_26360,N_25210,N_25272);
or U26361 (N_26361,N_25341,N_25407);
or U26362 (N_26362,N_25767,N_25677);
and U26363 (N_26363,N_25404,N_25766);
or U26364 (N_26364,N_25211,N_25426);
nand U26365 (N_26365,N_25333,N_25430);
or U26366 (N_26366,N_25396,N_25357);
nor U26367 (N_26367,N_25499,N_25655);
xor U26368 (N_26368,N_25342,N_25543);
nor U26369 (N_26369,N_25612,N_25532);
nand U26370 (N_26370,N_25771,N_25390);
and U26371 (N_26371,N_25567,N_25519);
xnor U26372 (N_26372,N_25640,N_25740);
nor U26373 (N_26373,N_25337,N_25380);
and U26374 (N_26374,N_25463,N_25738);
and U26375 (N_26375,N_25277,N_25358);
nand U26376 (N_26376,N_25749,N_25209);
or U26377 (N_26377,N_25699,N_25208);
xor U26378 (N_26378,N_25395,N_25414);
xnor U26379 (N_26379,N_25223,N_25447);
or U26380 (N_26380,N_25726,N_25279);
and U26381 (N_26381,N_25477,N_25342);
nand U26382 (N_26382,N_25747,N_25581);
nor U26383 (N_26383,N_25534,N_25764);
and U26384 (N_26384,N_25585,N_25495);
nand U26385 (N_26385,N_25328,N_25718);
nand U26386 (N_26386,N_25773,N_25633);
nor U26387 (N_26387,N_25200,N_25585);
and U26388 (N_26388,N_25724,N_25244);
and U26389 (N_26389,N_25508,N_25740);
or U26390 (N_26390,N_25290,N_25419);
and U26391 (N_26391,N_25669,N_25314);
or U26392 (N_26392,N_25416,N_25305);
xnor U26393 (N_26393,N_25791,N_25743);
xor U26394 (N_26394,N_25565,N_25521);
nand U26395 (N_26395,N_25570,N_25673);
nand U26396 (N_26396,N_25756,N_25647);
xnor U26397 (N_26397,N_25692,N_25675);
or U26398 (N_26398,N_25474,N_25520);
xnor U26399 (N_26399,N_25205,N_25290);
xnor U26400 (N_26400,N_26356,N_25855);
xnor U26401 (N_26401,N_26288,N_26018);
xor U26402 (N_26402,N_26274,N_26367);
nand U26403 (N_26403,N_26043,N_26286);
xnor U26404 (N_26404,N_26306,N_25982);
nor U26405 (N_26405,N_26250,N_26296);
nor U26406 (N_26406,N_26217,N_26010);
nor U26407 (N_26407,N_25834,N_26205);
xnor U26408 (N_26408,N_26111,N_26366);
and U26409 (N_26409,N_26307,N_25963);
xnor U26410 (N_26410,N_26284,N_26207);
or U26411 (N_26411,N_26131,N_25840);
nor U26412 (N_26412,N_26123,N_25891);
nand U26413 (N_26413,N_26329,N_25958);
xnor U26414 (N_26414,N_25972,N_26373);
and U26415 (N_26415,N_25992,N_26012);
nand U26416 (N_26416,N_25980,N_26099);
nor U26417 (N_26417,N_25813,N_25959);
and U26418 (N_26418,N_26232,N_26140);
nor U26419 (N_26419,N_26095,N_26362);
xor U26420 (N_26420,N_25938,N_25951);
nor U26421 (N_26421,N_26086,N_26093);
or U26422 (N_26422,N_26110,N_26187);
nor U26423 (N_26423,N_26080,N_25805);
xor U26424 (N_26424,N_26006,N_26069);
nand U26425 (N_26425,N_25875,N_26067);
and U26426 (N_26426,N_26100,N_26292);
nand U26427 (N_26427,N_26029,N_26231);
and U26428 (N_26428,N_25912,N_26312);
and U26429 (N_26429,N_26026,N_26386);
nand U26430 (N_26430,N_26127,N_26293);
nor U26431 (N_26431,N_26090,N_26215);
or U26432 (N_26432,N_26188,N_26039);
nand U26433 (N_26433,N_26098,N_26190);
or U26434 (N_26434,N_25970,N_25864);
or U26435 (N_26435,N_26271,N_26020);
xor U26436 (N_26436,N_26024,N_26339);
nor U26437 (N_26437,N_26199,N_26049);
xnor U26438 (N_26438,N_25858,N_26017);
or U26439 (N_26439,N_25818,N_25978);
nor U26440 (N_26440,N_26255,N_26332);
and U26441 (N_26441,N_26028,N_26163);
and U26442 (N_26442,N_25983,N_25872);
nor U26443 (N_26443,N_26139,N_26397);
xnor U26444 (N_26444,N_25894,N_26112);
xor U26445 (N_26445,N_26166,N_26096);
and U26446 (N_26446,N_26125,N_26240);
nand U26447 (N_26447,N_26372,N_26181);
nor U26448 (N_26448,N_25852,N_26005);
xor U26449 (N_26449,N_26036,N_25874);
or U26450 (N_26450,N_26137,N_26082);
and U26451 (N_26451,N_25800,N_26044);
and U26452 (N_26452,N_26243,N_26088);
or U26453 (N_26453,N_26394,N_25839);
or U26454 (N_26454,N_26389,N_26183);
nand U26455 (N_26455,N_26279,N_26229);
nor U26456 (N_26456,N_25842,N_26105);
xor U26457 (N_26457,N_26239,N_26132);
xnor U26458 (N_26458,N_26195,N_26073);
and U26459 (N_26459,N_26299,N_25907);
nand U26460 (N_26460,N_25808,N_25802);
and U26461 (N_26461,N_25847,N_26167);
nor U26462 (N_26462,N_25900,N_26056);
or U26463 (N_26463,N_26155,N_26013);
nor U26464 (N_26464,N_26103,N_26282);
or U26465 (N_26465,N_26050,N_25942);
nor U26466 (N_26466,N_26055,N_26101);
nor U26467 (N_26467,N_26025,N_25917);
nor U26468 (N_26468,N_26378,N_25865);
nand U26469 (N_26469,N_26331,N_26186);
and U26470 (N_26470,N_25944,N_26377);
xnor U26471 (N_26471,N_25923,N_26237);
or U26472 (N_26472,N_25962,N_26084);
xor U26473 (N_26473,N_26130,N_26149);
xnor U26474 (N_26474,N_26047,N_26064);
nor U26475 (N_26475,N_25868,N_26180);
and U26476 (N_26476,N_26168,N_26008);
and U26477 (N_26477,N_25835,N_26364);
xnor U26478 (N_26478,N_26325,N_26011);
or U26479 (N_26479,N_26152,N_26189);
xor U26480 (N_26480,N_26285,N_25908);
nor U26481 (N_26481,N_26330,N_25928);
xnor U26482 (N_26482,N_26388,N_26015);
xnor U26483 (N_26483,N_25999,N_25981);
nor U26484 (N_26484,N_26057,N_25904);
and U26485 (N_26485,N_26358,N_26294);
nand U26486 (N_26486,N_26194,N_26256);
and U26487 (N_26487,N_26048,N_26261);
xnor U26488 (N_26488,N_26041,N_25889);
and U26489 (N_26489,N_26122,N_26276);
and U26490 (N_26490,N_25987,N_26160);
nor U26491 (N_26491,N_26387,N_26248);
and U26492 (N_26492,N_25946,N_25961);
nor U26493 (N_26493,N_25861,N_26072);
and U26494 (N_26494,N_25906,N_26233);
xnor U26495 (N_26495,N_26398,N_25979);
or U26496 (N_26496,N_26310,N_26283);
or U26497 (N_26497,N_26003,N_25853);
nor U26498 (N_26498,N_25823,N_25899);
or U26499 (N_26499,N_26118,N_26263);
xor U26500 (N_26500,N_25817,N_26081);
nand U26501 (N_26501,N_25939,N_26382);
xor U26502 (N_26502,N_26230,N_26342);
nor U26503 (N_26503,N_25950,N_26319);
nand U26504 (N_26504,N_26291,N_26119);
or U26505 (N_26505,N_26000,N_26390);
nand U26506 (N_26506,N_26318,N_25914);
xor U26507 (N_26507,N_26254,N_25824);
or U26508 (N_26508,N_26363,N_26175);
or U26509 (N_26509,N_26204,N_26259);
or U26510 (N_26510,N_26009,N_25831);
nor U26511 (N_26511,N_26311,N_25867);
nor U26512 (N_26512,N_26275,N_25838);
nand U26513 (N_26513,N_25888,N_26385);
nor U26514 (N_26514,N_26128,N_25940);
or U26515 (N_26515,N_26162,N_26345);
and U26516 (N_26516,N_25827,N_26223);
xor U26517 (N_26517,N_26260,N_25971);
or U26518 (N_26518,N_26120,N_26225);
xnor U26519 (N_26519,N_26198,N_26265);
or U26520 (N_26520,N_26066,N_25816);
or U26521 (N_26521,N_25932,N_25828);
and U26522 (N_26522,N_25916,N_25991);
nor U26523 (N_26523,N_25869,N_26138);
nor U26524 (N_26524,N_26316,N_25954);
xor U26525 (N_26525,N_25856,N_25814);
xnor U26526 (N_26526,N_25969,N_26300);
and U26527 (N_26527,N_26034,N_25993);
and U26528 (N_26528,N_26091,N_26344);
and U26529 (N_26529,N_25929,N_25819);
xor U26530 (N_26530,N_25880,N_25968);
xnor U26531 (N_26531,N_26109,N_25952);
xnor U26532 (N_26532,N_25822,N_25803);
xor U26533 (N_26533,N_25809,N_25903);
nand U26534 (N_26534,N_25885,N_26359);
nor U26535 (N_26535,N_26063,N_25851);
nor U26536 (N_26536,N_26249,N_26102);
nand U26537 (N_26537,N_26145,N_26371);
and U26538 (N_26538,N_26161,N_26170);
and U26539 (N_26539,N_25873,N_26245);
or U26540 (N_26540,N_26246,N_26115);
and U26541 (N_26541,N_25989,N_25930);
nand U26542 (N_26542,N_26206,N_26121);
or U26543 (N_26543,N_26171,N_26032);
nand U26544 (N_26544,N_26257,N_26060);
or U26545 (N_26545,N_26165,N_26236);
xor U26546 (N_26546,N_26308,N_26244);
nor U26547 (N_26547,N_26164,N_26320);
nand U26548 (N_26548,N_26361,N_25833);
nor U26549 (N_26549,N_26226,N_26335);
or U26550 (N_26550,N_25804,N_25882);
nor U26551 (N_26551,N_26376,N_26391);
nand U26552 (N_26552,N_25941,N_25883);
xnor U26553 (N_26553,N_25896,N_26169);
xor U26554 (N_26554,N_25815,N_25964);
nand U26555 (N_26555,N_26304,N_26079);
nor U26556 (N_26556,N_26228,N_26357);
or U26557 (N_26557,N_26322,N_26258);
or U26558 (N_26558,N_25812,N_26077);
and U26559 (N_26559,N_26174,N_26191);
or U26560 (N_26560,N_26143,N_26369);
xor U26561 (N_26561,N_26117,N_26089);
and U26562 (N_26562,N_26305,N_26301);
xor U26563 (N_26563,N_25863,N_25931);
and U26564 (N_26564,N_26173,N_26042);
nand U26565 (N_26565,N_26220,N_26019);
nor U26566 (N_26566,N_26347,N_25850);
xnor U26567 (N_26567,N_26251,N_26197);
nand U26568 (N_26568,N_26134,N_25965);
and U26569 (N_26569,N_26272,N_25871);
and U26570 (N_26570,N_26178,N_26092);
nand U26571 (N_26571,N_26336,N_25984);
xnor U26572 (N_26572,N_26287,N_26070);
or U26573 (N_26573,N_26062,N_26201);
nor U26574 (N_26574,N_26177,N_26348);
nor U26575 (N_26575,N_26213,N_26150);
and U26576 (N_26576,N_25830,N_26303);
nor U26577 (N_26577,N_25947,N_26295);
and U26578 (N_26578,N_26212,N_26326);
and U26579 (N_26579,N_25943,N_25821);
or U26580 (N_26580,N_26315,N_25876);
xnor U26581 (N_26581,N_26002,N_26352);
or U26582 (N_26582,N_26076,N_26214);
xnor U26583 (N_26583,N_26065,N_26346);
or U26584 (N_26584,N_26269,N_26341);
nand U26585 (N_26585,N_26040,N_26083);
nor U26586 (N_26586,N_26061,N_26297);
nand U26587 (N_26587,N_25998,N_25966);
or U26588 (N_26588,N_26349,N_26046);
nor U26589 (N_26589,N_26350,N_26222);
nand U26590 (N_26590,N_26298,N_26266);
or U26591 (N_26591,N_26146,N_26124);
nor U26592 (N_26592,N_26192,N_26333);
xnor U26593 (N_26593,N_26153,N_25977);
or U26594 (N_26594,N_26075,N_25886);
nor U26595 (N_26595,N_26219,N_25953);
nand U26596 (N_26596,N_26211,N_25948);
nand U26597 (N_26597,N_26196,N_25811);
nor U26598 (N_26598,N_25897,N_25973);
xor U26599 (N_26599,N_25937,N_26370);
nand U26600 (N_26600,N_26375,N_25994);
nand U26601 (N_26601,N_26224,N_26338);
xnor U26602 (N_26602,N_26097,N_25846);
xor U26603 (N_26603,N_26221,N_26277);
xnor U26604 (N_26604,N_26054,N_26104);
and U26605 (N_26605,N_26156,N_25920);
nand U26606 (N_26606,N_25806,N_26053);
and U26607 (N_26607,N_26147,N_25935);
nand U26608 (N_26608,N_26085,N_25967);
nor U26609 (N_26609,N_26379,N_26045);
xor U26610 (N_26610,N_26135,N_26384);
and U26611 (N_26611,N_26136,N_26126);
nor U26612 (N_26612,N_26396,N_25960);
nand U26613 (N_26613,N_26252,N_26354);
xor U26614 (N_26614,N_26216,N_26253);
and U26615 (N_26615,N_26157,N_26203);
nand U26616 (N_26616,N_25974,N_26328);
and U26617 (N_26617,N_26151,N_26129);
nand U26618 (N_26618,N_25915,N_26133);
nor U26619 (N_26619,N_25841,N_25919);
or U26620 (N_26620,N_25878,N_25843);
and U26621 (N_26621,N_25866,N_25859);
nand U26622 (N_26622,N_25837,N_26392);
nor U26623 (N_26623,N_26242,N_25902);
nand U26624 (N_26624,N_26068,N_25810);
nor U26625 (N_26625,N_26321,N_26324);
and U26626 (N_26626,N_25934,N_26159);
nor U26627 (N_26627,N_25832,N_26353);
xor U26628 (N_26628,N_26393,N_26148);
xor U26629 (N_26629,N_25975,N_26154);
and U26630 (N_26630,N_26038,N_25825);
or U26631 (N_26631,N_26193,N_26247);
and U26632 (N_26632,N_26383,N_26340);
nor U26633 (N_26633,N_26327,N_25895);
nand U26634 (N_26634,N_26051,N_25957);
and U26635 (N_26635,N_26023,N_26030);
or U26636 (N_26636,N_26141,N_25955);
or U26637 (N_26637,N_25918,N_26202);
nand U26638 (N_26638,N_26262,N_26314);
or U26639 (N_26639,N_26343,N_26027);
nand U26640 (N_26640,N_26035,N_25936);
nand U26641 (N_26641,N_26158,N_25924);
xnor U26642 (N_26642,N_25986,N_25890);
or U26643 (N_26643,N_25926,N_25949);
nand U26644 (N_26644,N_26142,N_26380);
and U26645 (N_26645,N_26113,N_26280);
and U26646 (N_26646,N_25901,N_26176);
xnor U26647 (N_26647,N_25945,N_25881);
nand U26648 (N_26648,N_26087,N_25892);
nand U26649 (N_26649,N_25893,N_26399);
and U26650 (N_26650,N_26270,N_26031);
or U26651 (N_26651,N_25836,N_25925);
or U26652 (N_26652,N_25887,N_25913);
xor U26653 (N_26653,N_26241,N_26273);
or U26654 (N_26654,N_26278,N_26052);
and U26655 (N_26655,N_25857,N_26374);
nand U26656 (N_26656,N_26094,N_25933);
xor U26657 (N_26657,N_26014,N_25801);
or U26658 (N_26658,N_26116,N_25898);
nand U26659 (N_26659,N_25879,N_26337);
nor U26660 (N_26660,N_26078,N_26037);
nor U26661 (N_26661,N_25862,N_26264);
or U26662 (N_26662,N_25985,N_26395);
xnor U26663 (N_26663,N_26004,N_25956);
and U26664 (N_26664,N_26033,N_25848);
xor U26665 (N_26665,N_26281,N_26114);
and U26666 (N_26666,N_26218,N_26209);
xnor U26667 (N_26667,N_25854,N_25990);
or U26668 (N_26668,N_25829,N_26355);
nor U26669 (N_26669,N_26200,N_26227);
nand U26670 (N_26670,N_26360,N_25844);
nor U26671 (N_26671,N_26365,N_25988);
xor U26672 (N_26672,N_26058,N_26144);
nand U26673 (N_26673,N_26022,N_26179);
or U26674 (N_26674,N_26172,N_26238);
and U26675 (N_26675,N_26368,N_26106);
nor U26676 (N_26676,N_25976,N_25870);
xnor U26677 (N_26677,N_26071,N_25884);
or U26678 (N_26678,N_25997,N_26381);
nor U26679 (N_26679,N_26059,N_25996);
xor U26680 (N_26680,N_25849,N_25820);
and U26681 (N_26681,N_26267,N_26351);
nand U26682 (N_26682,N_25995,N_25910);
nand U26683 (N_26683,N_25807,N_26313);
nand U26684 (N_26684,N_26185,N_26210);
xor U26685 (N_26685,N_26184,N_26074);
and U26686 (N_26686,N_25905,N_25826);
xor U26687 (N_26687,N_26016,N_26108);
and U26688 (N_26688,N_26268,N_25927);
and U26689 (N_26689,N_26208,N_26235);
or U26690 (N_26690,N_25845,N_26334);
xor U26691 (N_26691,N_26234,N_26021);
or U26692 (N_26692,N_25877,N_25922);
nand U26693 (N_26693,N_25911,N_26302);
or U26694 (N_26694,N_26290,N_26182);
xor U26695 (N_26695,N_25860,N_25909);
nand U26696 (N_26696,N_26107,N_25921);
and U26697 (N_26697,N_26317,N_26007);
nand U26698 (N_26698,N_26323,N_26001);
nand U26699 (N_26699,N_26309,N_26289);
nor U26700 (N_26700,N_26062,N_26254);
xnor U26701 (N_26701,N_26364,N_25910);
and U26702 (N_26702,N_26030,N_26350);
or U26703 (N_26703,N_26296,N_25980);
nand U26704 (N_26704,N_25805,N_25949);
or U26705 (N_26705,N_26113,N_26028);
and U26706 (N_26706,N_25980,N_25872);
and U26707 (N_26707,N_26351,N_26150);
nand U26708 (N_26708,N_25918,N_25990);
nand U26709 (N_26709,N_25886,N_26052);
and U26710 (N_26710,N_26099,N_25974);
and U26711 (N_26711,N_25826,N_26218);
nor U26712 (N_26712,N_25949,N_26241);
nor U26713 (N_26713,N_25886,N_26167);
nand U26714 (N_26714,N_26041,N_26371);
nor U26715 (N_26715,N_25987,N_26222);
or U26716 (N_26716,N_26189,N_25973);
xnor U26717 (N_26717,N_25890,N_25899);
or U26718 (N_26718,N_26213,N_25938);
nand U26719 (N_26719,N_25903,N_26393);
or U26720 (N_26720,N_26294,N_26169);
or U26721 (N_26721,N_26383,N_26054);
xnor U26722 (N_26722,N_26129,N_26371);
nor U26723 (N_26723,N_26308,N_25878);
nor U26724 (N_26724,N_26024,N_26052);
xnor U26725 (N_26725,N_26050,N_25957);
xnor U26726 (N_26726,N_26233,N_25976);
nor U26727 (N_26727,N_26339,N_26049);
or U26728 (N_26728,N_26068,N_25828);
xor U26729 (N_26729,N_25874,N_26003);
xnor U26730 (N_26730,N_26356,N_25972);
nand U26731 (N_26731,N_26250,N_26273);
xor U26732 (N_26732,N_25867,N_26364);
xor U26733 (N_26733,N_26257,N_26019);
or U26734 (N_26734,N_25802,N_25926);
nand U26735 (N_26735,N_26356,N_26257);
nand U26736 (N_26736,N_26170,N_26200);
and U26737 (N_26737,N_26341,N_26358);
and U26738 (N_26738,N_26251,N_25856);
nor U26739 (N_26739,N_25836,N_26368);
and U26740 (N_26740,N_26124,N_26232);
xor U26741 (N_26741,N_26134,N_26075);
nand U26742 (N_26742,N_25892,N_26038);
and U26743 (N_26743,N_26236,N_25979);
nand U26744 (N_26744,N_25991,N_26056);
nand U26745 (N_26745,N_25856,N_25865);
nand U26746 (N_26746,N_26208,N_25819);
nor U26747 (N_26747,N_25928,N_25999);
nand U26748 (N_26748,N_26036,N_25960);
nor U26749 (N_26749,N_25964,N_26153);
and U26750 (N_26750,N_25857,N_26019);
nand U26751 (N_26751,N_26037,N_26280);
nand U26752 (N_26752,N_25921,N_26126);
and U26753 (N_26753,N_25870,N_26258);
nand U26754 (N_26754,N_25930,N_26326);
or U26755 (N_26755,N_26265,N_26289);
and U26756 (N_26756,N_25940,N_26259);
and U26757 (N_26757,N_26269,N_25909);
xor U26758 (N_26758,N_26193,N_26342);
xor U26759 (N_26759,N_25935,N_25911);
nor U26760 (N_26760,N_26164,N_26130);
nand U26761 (N_26761,N_26216,N_26023);
and U26762 (N_26762,N_26239,N_25866);
nand U26763 (N_26763,N_26378,N_26264);
nand U26764 (N_26764,N_25916,N_26213);
nor U26765 (N_26765,N_26246,N_26373);
nand U26766 (N_26766,N_26130,N_26294);
nor U26767 (N_26767,N_25948,N_26263);
nor U26768 (N_26768,N_26316,N_26348);
and U26769 (N_26769,N_25974,N_25950);
xnor U26770 (N_26770,N_26391,N_25921);
nor U26771 (N_26771,N_26369,N_26316);
nand U26772 (N_26772,N_26318,N_26331);
or U26773 (N_26773,N_25819,N_25941);
nand U26774 (N_26774,N_25830,N_25890);
and U26775 (N_26775,N_25883,N_26089);
xor U26776 (N_26776,N_25946,N_26376);
xnor U26777 (N_26777,N_26034,N_25862);
and U26778 (N_26778,N_25843,N_26011);
nor U26779 (N_26779,N_26169,N_26044);
or U26780 (N_26780,N_25952,N_26040);
or U26781 (N_26781,N_26270,N_26392);
and U26782 (N_26782,N_26250,N_25807);
nor U26783 (N_26783,N_26075,N_25949);
nor U26784 (N_26784,N_26357,N_26223);
or U26785 (N_26785,N_26256,N_26323);
nor U26786 (N_26786,N_26152,N_25920);
or U26787 (N_26787,N_25944,N_25890);
or U26788 (N_26788,N_26140,N_26188);
xor U26789 (N_26789,N_25986,N_25805);
nand U26790 (N_26790,N_26388,N_25841);
and U26791 (N_26791,N_25952,N_26395);
and U26792 (N_26792,N_26164,N_26220);
xnor U26793 (N_26793,N_25888,N_25904);
nor U26794 (N_26794,N_26027,N_25988);
nor U26795 (N_26795,N_26029,N_25865);
and U26796 (N_26796,N_25855,N_26080);
nor U26797 (N_26797,N_25960,N_25986);
nor U26798 (N_26798,N_25924,N_25826);
xor U26799 (N_26799,N_26267,N_25853);
xor U26800 (N_26800,N_25983,N_25915);
or U26801 (N_26801,N_25848,N_26182);
or U26802 (N_26802,N_26345,N_25871);
xnor U26803 (N_26803,N_26077,N_26088);
nand U26804 (N_26804,N_26112,N_26233);
or U26805 (N_26805,N_25957,N_26307);
and U26806 (N_26806,N_25862,N_25876);
and U26807 (N_26807,N_26178,N_25919);
or U26808 (N_26808,N_25813,N_26303);
or U26809 (N_26809,N_26369,N_26241);
nand U26810 (N_26810,N_25911,N_25964);
xnor U26811 (N_26811,N_25900,N_26271);
nor U26812 (N_26812,N_25873,N_25965);
and U26813 (N_26813,N_25912,N_26228);
or U26814 (N_26814,N_25967,N_25904);
or U26815 (N_26815,N_26190,N_26208);
nor U26816 (N_26816,N_25996,N_26184);
or U26817 (N_26817,N_25901,N_25868);
or U26818 (N_26818,N_25929,N_25828);
nand U26819 (N_26819,N_26109,N_26054);
xor U26820 (N_26820,N_25820,N_26345);
and U26821 (N_26821,N_25902,N_26315);
nand U26822 (N_26822,N_25916,N_25903);
nand U26823 (N_26823,N_26389,N_26057);
and U26824 (N_26824,N_26079,N_25851);
and U26825 (N_26825,N_26134,N_25901);
xor U26826 (N_26826,N_26045,N_25927);
xnor U26827 (N_26827,N_26133,N_25851);
nor U26828 (N_26828,N_25861,N_26174);
xor U26829 (N_26829,N_26313,N_26048);
xnor U26830 (N_26830,N_26298,N_25935);
or U26831 (N_26831,N_26287,N_26363);
nand U26832 (N_26832,N_25930,N_25987);
nor U26833 (N_26833,N_25946,N_26220);
xor U26834 (N_26834,N_26309,N_26077);
nor U26835 (N_26835,N_25833,N_26118);
and U26836 (N_26836,N_26030,N_26200);
nand U26837 (N_26837,N_25955,N_26189);
xnor U26838 (N_26838,N_26215,N_26213);
or U26839 (N_26839,N_26384,N_26312);
xor U26840 (N_26840,N_26132,N_26301);
and U26841 (N_26841,N_25869,N_26393);
nand U26842 (N_26842,N_26177,N_26172);
nand U26843 (N_26843,N_26238,N_26326);
and U26844 (N_26844,N_26172,N_26039);
nor U26845 (N_26845,N_26306,N_25942);
and U26846 (N_26846,N_26233,N_26201);
nor U26847 (N_26847,N_26147,N_25838);
nand U26848 (N_26848,N_25887,N_25890);
and U26849 (N_26849,N_26255,N_26134);
nand U26850 (N_26850,N_25825,N_26152);
xor U26851 (N_26851,N_25820,N_25933);
xor U26852 (N_26852,N_26235,N_26261);
or U26853 (N_26853,N_25808,N_25888);
xor U26854 (N_26854,N_26100,N_26394);
and U26855 (N_26855,N_25993,N_26311);
and U26856 (N_26856,N_26092,N_26205);
xnor U26857 (N_26857,N_26258,N_25808);
xnor U26858 (N_26858,N_26116,N_26165);
nor U26859 (N_26859,N_26215,N_25816);
or U26860 (N_26860,N_26358,N_26217);
and U26861 (N_26861,N_26004,N_26368);
nor U26862 (N_26862,N_26272,N_25806);
nor U26863 (N_26863,N_26245,N_26021);
nand U26864 (N_26864,N_26127,N_26095);
xor U26865 (N_26865,N_26131,N_26326);
or U26866 (N_26866,N_26246,N_26185);
xor U26867 (N_26867,N_26201,N_26351);
nand U26868 (N_26868,N_26246,N_26392);
and U26869 (N_26869,N_26263,N_25859);
nand U26870 (N_26870,N_25900,N_25805);
xor U26871 (N_26871,N_26246,N_26243);
or U26872 (N_26872,N_26058,N_26273);
nor U26873 (N_26873,N_26388,N_26201);
and U26874 (N_26874,N_26357,N_26099);
nand U26875 (N_26875,N_25991,N_26044);
and U26876 (N_26876,N_26356,N_26398);
nand U26877 (N_26877,N_25823,N_26179);
nand U26878 (N_26878,N_25923,N_25974);
or U26879 (N_26879,N_26236,N_26117);
xnor U26880 (N_26880,N_25884,N_26177);
xor U26881 (N_26881,N_26015,N_26164);
nor U26882 (N_26882,N_25860,N_25897);
and U26883 (N_26883,N_26201,N_26009);
nor U26884 (N_26884,N_25818,N_26315);
nor U26885 (N_26885,N_26378,N_26381);
nand U26886 (N_26886,N_25906,N_26108);
xor U26887 (N_26887,N_25819,N_25916);
or U26888 (N_26888,N_25979,N_26254);
nand U26889 (N_26889,N_26164,N_25891);
or U26890 (N_26890,N_26114,N_26355);
nand U26891 (N_26891,N_26315,N_26024);
nor U26892 (N_26892,N_25926,N_25947);
or U26893 (N_26893,N_26370,N_26262);
or U26894 (N_26894,N_26311,N_26321);
and U26895 (N_26895,N_26060,N_26128);
xnor U26896 (N_26896,N_26219,N_25864);
nor U26897 (N_26897,N_26112,N_26027);
xor U26898 (N_26898,N_25982,N_25822);
nand U26899 (N_26899,N_25818,N_25932);
nand U26900 (N_26900,N_26046,N_25885);
or U26901 (N_26901,N_26325,N_26381);
and U26902 (N_26902,N_25899,N_26345);
and U26903 (N_26903,N_26168,N_26379);
nor U26904 (N_26904,N_26327,N_26141);
or U26905 (N_26905,N_25817,N_26144);
xor U26906 (N_26906,N_26202,N_25952);
and U26907 (N_26907,N_26119,N_25920);
xnor U26908 (N_26908,N_26144,N_26281);
and U26909 (N_26909,N_26180,N_25900);
and U26910 (N_26910,N_26281,N_25938);
or U26911 (N_26911,N_26008,N_26033);
nand U26912 (N_26912,N_26243,N_26065);
nor U26913 (N_26913,N_26102,N_25973);
and U26914 (N_26914,N_26135,N_25956);
xor U26915 (N_26915,N_26126,N_26383);
xnor U26916 (N_26916,N_26349,N_26072);
xor U26917 (N_26917,N_26016,N_26345);
nor U26918 (N_26918,N_26321,N_26351);
nor U26919 (N_26919,N_26299,N_26291);
and U26920 (N_26920,N_26178,N_26321);
and U26921 (N_26921,N_26042,N_25992);
and U26922 (N_26922,N_26289,N_26144);
nor U26923 (N_26923,N_26053,N_26155);
or U26924 (N_26924,N_26286,N_26169);
and U26925 (N_26925,N_26344,N_26130);
and U26926 (N_26926,N_25997,N_26119);
nor U26927 (N_26927,N_26370,N_26357);
and U26928 (N_26928,N_25942,N_26072);
and U26929 (N_26929,N_25802,N_25918);
xnor U26930 (N_26930,N_25883,N_26245);
nand U26931 (N_26931,N_26189,N_26289);
nor U26932 (N_26932,N_26295,N_25874);
xor U26933 (N_26933,N_26041,N_26059);
or U26934 (N_26934,N_26063,N_25982);
xor U26935 (N_26935,N_25961,N_25964);
nor U26936 (N_26936,N_26013,N_25978);
and U26937 (N_26937,N_26016,N_26158);
and U26938 (N_26938,N_26222,N_26273);
nand U26939 (N_26939,N_26024,N_26195);
xor U26940 (N_26940,N_25949,N_26029);
or U26941 (N_26941,N_26397,N_25892);
or U26942 (N_26942,N_26077,N_25894);
nand U26943 (N_26943,N_26237,N_25901);
or U26944 (N_26944,N_26010,N_26239);
and U26945 (N_26945,N_26034,N_26233);
xor U26946 (N_26946,N_25999,N_26066);
xnor U26947 (N_26947,N_26090,N_25852);
xor U26948 (N_26948,N_25968,N_26292);
or U26949 (N_26949,N_25911,N_25946);
xnor U26950 (N_26950,N_26390,N_25849);
and U26951 (N_26951,N_26394,N_25870);
or U26952 (N_26952,N_26310,N_25926);
nand U26953 (N_26953,N_26040,N_26049);
and U26954 (N_26954,N_25923,N_26224);
xor U26955 (N_26955,N_26178,N_26144);
or U26956 (N_26956,N_25949,N_25884);
xnor U26957 (N_26957,N_25816,N_26166);
xor U26958 (N_26958,N_26208,N_26091);
xor U26959 (N_26959,N_26270,N_26339);
nor U26960 (N_26960,N_25906,N_25983);
nor U26961 (N_26961,N_26004,N_25875);
and U26962 (N_26962,N_26340,N_26398);
and U26963 (N_26963,N_25809,N_26287);
and U26964 (N_26964,N_26370,N_25998);
or U26965 (N_26965,N_25884,N_25844);
nand U26966 (N_26966,N_25893,N_25859);
or U26967 (N_26967,N_26384,N_26372);
or U26968 (N_26968,N_25948,N_25820);
xor U26969 (N_26969,N_26194,N_26202);
and U26970 (N_26970,N_26201,N_26165);
nand U26971 (N_26971,N_26044,N_26099);
nand U26972 (N_26972,N_25893,N_25949);
xor U26973 (N_26973,N_26028,N_25872);
xnor U26974 (N_26974,N_26369,N_26255);
nand U26975 (N_26975,N_26315,N_26012);
or U26976 (N_26976,N_25900,N_25940);
nand U26977 (N_26977,N_26203,N_26343);
or U26978 (N_26978,N_26222,N_26220);
xor U26979 (N_26979,N_26232,N_26085);
nor U26980 (N_26980,N_26371,N_25916);
xnor U26981 (N_26981,N_26144,N_25973);
nand U26982 (N_26982,N_26234,N_26033);
and U26983 (N_26983,N_26055,N_26258);
or U26984 (N_26984,N_26386,N_25995);
or U26985 (N_26985,N_26127,N_26280);
nor U26986 (N_26986,N_25995,N_26125);
and U26987 (N_26987,N_26346,N_26047);
and U26988 (N_26988,N_26199,N_26390);
nand U26989 (N_26989,N_26288,N_26307);
or U26990 (N_26990,N_25940,N_26119);
and U26991 (N_26991,N_26020,N_25873);
nand U26992 (N_26992,N_26193,N_25903);
or U26993 (N_26993,N_25816,N_26050);
nand U26994 (N_26994,N_26100,N_26053);
and U26995 (N_26995,N_26113,N_25848);
nand U26996 (N_26996,N_26035,N_26249);
xor U26997 (N_26997,N_26379,N_26108);
xnor U26998 (N_26998,N_26008,N_25969);
xnor U26999 (N_26999,N_25940,N_26319);
xor U27000 (N_27000,N_26534,N_26511);
nand U27001 (N_27001,N_26430,N_26881);
xor U27002 (N_27002,N_26497,N_26965);
nand U27003 (N_27003,N_26767,N_26475);
nor U27004 (N_27004,N_26436,N_26720);
or U27005 (N_27005,N_26569,N_26692);
xnor U27006 (N_27006,N_26760,N_26893);
and U27007 (N_27007,N_26581,N_26558);
nand U27008 (N_27008,N_26509,N_26606);
nand U27009 (N_27009,N_26525,N_26707);
xnor U27010 (N_27010,N_26660,N_26638);
and U27011 (N_27011,N_26764,N_26761);
xnor U27012 (N_27012,N_26409,N_26712);
or U27013 (N_27013,N_26535,N_26536);
or U27014 (N_27014,N_26822,N_26626);
nor U27015 (N_27015,N_26728,N_26461);
or U27016 (N_27016,N_26680,N_26715);
xnor U27017 (N_27017,N_26691,N_26485);
nand U27018 (N_27018,N_26916,N_26957);
or U27019 (N_27019,N_26665,N_26912);
nor U27020 (N_27020,N_26890,N_26421);
xnor U27021 (N_27021,N_26827,N_26533);
nand U27022 (N_27022,N_26964,N_26997);
xnor U27023 (N_27023,N_26849,N_26984);
and U27024 (N_27024,N_26620,N_26555);
and U27025 (N_27025,N_26447,N_26587);
nor U27026 (N_27026,N_26867,N_26631);
nor U27027 (N_27027,N_26412,N_26943);
nor U27028 (N_27028,N_26426,N_26995);
and U27029 (N_27029,N_26757,N_26592);
xnor U27030 (N_27030,N_26899,N_26448);
and U27031 (N_27031,N_26579,N_26801);
nor U27032 (N_27032,N_26891,N_26422);
nand U27033 (N_27033,N_26806,N_26809);
nor U27034 (N_27034,N_26419,N_26736);
and U27035 (N_27035,N_26664,N_26451);
nor U27036 (N_27036,N_26578,N_26753);
xnor U27037 (N_27037,N_26634,N_26953);
or U27038 (N_27038,N_26661,N_26940);
xnor U27039 (N_27039,N_26700,N_26679);
or U27040 (N_27040,N_26817,N_26971);
xor U27041 (N_27041,N_26591,N_26919);
and U27042 (N_27042,N_26793,N_26945);
xor U27043 (N_27043,N_26988,N_26411);
nand U27044 (N_27044,N_26444,N_26505);
nor U27045 (N_27045,N_26462,N_26671);
xor U27046 (N_27046,N_26568,N_26788);
or U27047 (N_27047,N_26762,N_26994);
or U27048 (N_27048,N_26790,N_26433);
or U27049 (N_27049,N_26922,N_26752);
xnor U27050 (N_27050,N_26657,N_26585);
nor U27051 (N_27051,N_26494,N_26835);
and U27052 (N_27052,N_26754,N_26812);
xnor U27053 (N_27053,N_26561,N_26501);
xnor U27054 (N_27054,N_26763,N_26539);
nand U27055 (N_27055,N_26550,N_26863);
xor U27056 (N_27056,N_26903,N_26844);
nand U27057 (N_27057,N_26693,N_26482);
and U27058 (N_27058,N_26552,N_26711);
or U27059 (N_27059,N_26888,N_26948);
nand U27060 (N_27060,N_26427,N_26658);
nand U27061 (N_27061,N_26437,N_26493);
xnor U27062 (N_27062,N_26589,N_26554);
or U27063 (N_27063,N_26416,N_26443);
and U27064 (N_27064,N_26960,N_26842);
xor U27065 (N_27065,N_26926,N_26405);
and U27066 (N_27066,N_26771,N_26567);
and U27067 (N_27067,N_26489,N_26998);
or U27068 (N_27068,N_26406,N_26531);
and U27069 (N_27069,N_26713,N_26845);
nor U27070 (N_27070,N_26871,N_26769);
and U27071 (N_27071,N_26513,N_26917);
or U27072 (N_27072,N_26966,N_26928);
or U27073 (N_27073,N_26467,N_26478);
and U27074 (N_27074,N_26963,N_26481);
or U27075 (N_27075,N_26751,N_26559);
or U27076 (N_27076,N_26446,N_26802);
and U27077 (N_27077,N_26933,N_26521);
nor U27078 (N_27078,N_26843,N_26516);
or U27079 (N_27079,N_26607,N_26429);
xnor U27080 (N_27080,N_26770,N_26600);
nor U27081 (N_27081,N_26732,N_26435);
xor U27082 (N_27082,N_26886,N_26854);
xnor U27083 (N_27083,N_26979,N_26833);
or U27084 (N_27084,N_26684,N_26519);
nand U27085 (N_27085,N_26683,N_26413);
and U27086 (N_27086,N_26955,N_26847);
or U27087 (N_27087,N_26924,N_26479);
nand U27088 (N_27088,N_26520,N_26417);
nand U27089 (N_27089,N_26706,N_26738);
nor U27090 (N_27090,N_26789,N_26915);
nand U27091 (N_27091,N_26611,N_26441);
or U27092 (N_27092,N_26425,N_26852);
or U27093 (N_27093,N_26887,N_26911);
or U27094 (N_27094,N_26604,N_26747);
nor U27095 (N_27095,N_26947,N_26541);
nand U27096 (N_27096,N_26820,N_26543);
nand U27097 (N_27097,N_26609,N_26708);
nor U27098 (N_27098,N_26458,N_26583);
nand U27099 (N_27099,N_26480,N_26510);
xor U27100 (N_27100,N_26838,N_26618);
and U27101 (N_27101,N_26885,N_26623);
and U27102 (N_27102,N_26724,N_26526);
and U27103 (N_27103,N_26449,N_26640);
and U27104 (N_27104,N_26949,N_26872);
nor U27105 (N_27105,N_26938,N_26841);
and U27106 (N_27106,N_26798,N_26597);
or U27107 (N_27107,N_26402,N_26704);
nor U27108 (N_27108,N_26766,N_26666);
nand U27109 (N_27109,N_26682,N_26669);
and U27110 (N_27110,N_26678,N_26564);
nand U27111 (N_27111,N_26676,N_26641);
nand U27112 (N_27112,N_26726,N_26976);
nand U27113 (N_27113,N_26821,N_26637);
or U27114 (N_27114,N_26931,N_26951);
xnor U27115 (N_27115,N_26659,N_26644);
and U27116 (N_27116,N_26791,N_26783);
nand U27117 (N_27117,N_26981,N_26935);
nor U27118 (N_27118,N_26892,N_26739);
nor U27119 (N_27119,N_26962,N_26452);
nand U27120 (N_27120,N_26703,N_26839);
and U27121 (N_27121,N_26990,N_26826);
xnor U27122 (N_27122,N_26909,N_26616);
xor U27123 (N_27123,N_26746,N_26484);
nand U27124 (N_27124,N_26818,N_26792);
xor U27125 (N_27125,N_26829,N_26648);
or U27126 (N_27126,N_26614,N_26908);
xor U27127 (N_27127,N_26491,N_26824);
nand U27128 (N_27128,N_26407,N_26512);
or U27129 (N_27129,N_26400,N_26575);
and U27130 (N_27130,N_26741,N_26950);
nand U27131 (N_27131,N_26701,N_26477);
xor U27132 (N_27132,N_26819,N_26864);
nand U27133 (N_27133,N_26492,N_26488);
and U27134 (N_27134,N_26621,N_26813);
nand U27135 (N_27135,N_26923,N_26808);
nand U27136 (N_27136,N_26929,N_26972);
or U27137 (N_27137,N_26530,N_26508);
nor U27138 (N_27138,N_26978,N_26776);
xnor U27139 (N_27139,N_26410,N_26557);
or U27140 (N_27140,N_26667,N_26731);
and U27141 (N_27141,N_26651,N_26906);
or U27142 (N_27142,N_26765,N_26471);
and U27143 (N_27143,N_26628,N_26782);
nand U27144 (N_27144,N_26549,N_26642);
or U27145 (N_27145,N_26855,N_26743);
nand U27146 (N_27146,N_26727,N_26499);
or U27147 (N_27147,N_26875,N_26565);
or U27148 (N_27148,N_26897,N_26846);
or U27149 (N_27149,N_26681,N_26830);
and U27150 (N_27150,N_26880,N_26959);
or U27151 (N_27151,N_26689,N_26463);
or U27152 (N_27152,N_26930,N_26517);
and U27153 (N_27153,N_26570,N_26528);
xor U27154 (N_27154,N_26551,N_26453);
and U27155 (N_27155,N_26869,N_26744);
and U27156 (N_27156,N_26646,N_26457);
xor U27157 (N_27157,N_26672,N_26889);
and U27158 (N_27158,N_26828,N_26944);
xor U27159 (N_27159,N_26755,N_26850);
nor U27160 (N_27160,N_26615,N_26851);
nand U27161 (N_27161,N_26625,N_26487);
nand U27162 (N_27162,N_26901,N_26857);
xor U27163 (N_27163,N_26454,N_26633);
nand U27164 (N_27164,N_26627,N_26469);
or U27165 (N_27165,N_26431,N_26905);
or U27166 (N_27166,N_26445,N_26939);
and U27167 (N_27167,N_26593,N_26868);
or U27168 (N_27168,N_26612,N_26836);
or U27169 (N_27169,N_26927,N_26450);
xor U27170 (N_27170,N_26473,N_26687);
xnor U27171 (N_27171,N_26987,N_26690);
xnor U27172 (N_27172,N_26415,N_26538);
xor U27173 (N_27173,N_26999,N_26879);
nand U27174 (N_27174,N_26582,N_26418);
xor U27175 (N_27175,N_26737,N_26702);
and U27176 (N_27176,N_26942,N_26518);
nand U27177 (N_27177,N_26540,N_26653);
nor U27178 (N_27178,N_26932,N_26602);
or U27179 (N_27179,N_26865,N_26874);
and U27180 (N_27180,N_26476,N_26803);
and U27181 (N_27181,N_26870,N_26758);
and U27182 (N_27182,N_26723,N_26810);
or U27183 (N_27183,N_26749,N_26975);
xor U27184 (N_27184,N_26668,N_26502);
nand U27185 (N_27185,N_26853,N_26785);
and U27186 (N_27186,N_26688,N_26556);
xnor U27187 (N_27187,N_26455,N_26725);
nand U27188 (N_27188,N_26778,N_26873);
xnor U27189 (N_27189,N_26925,N_26710);
nand U27190 (N_27190,N_26652,N_26663);
nand U27191 (N_27191,N_26805,N_26670);
xor U27192 (N_27192,N_26442,N_26647);
nand U27193 (N_27193,N_26734,N_26622);
nand U27194 (N_27194,N_26472,N_26866);
or U27195 (N_27195,N_26639,N_26542);
or U27196 (N_27196,N_26617,N_26861);
nor U27197 (N_27197,N_26548,N_26636);
and U27198 (N_27198,N_26498,N_26496);
xnor U27199 (N_27199,N_26795,N_26807);
nor U27200 (N_27200,N_26895,N_26596);
nor U27201 (N_27201,N_26748,N_26759);
nor U27202 (N_27202,N_26774,N_26576);
xnor U27203 (N_27203,N_26650,N_26896);
nand U27204 (N_27204,N_26654,N_26946);
nand U27205 (N_27205,N_26577,N_26465);
and U27206 (N_27206,N_26649,N_26506);
xor U27207 (N_27207,N_26860,N_26694);
and U27208 (N_27208,N_26717,N_26401);
or U27209 (N_27209,N_26490,N_26794);
or U27210 (N_27210,N_26674,N_26958);
nand U27211 (N_27211,N_26503,N_26982);
or U27212 (N_27212,N_26884,N_26574);
xor U27213 (N_27213,N_26424,N_26719);
and U27214 (N_27214,N_26718,N_26466);
nand U27215 (N_27215,N_26594,N_26643);
nand U27216 (N_27216,N_26936,N_26941);
nor U27217 (N_27217,N_26848,N_26775);
nor U27218 (N_27218,N_26745,N_26740);
or U27219 (N_27219,N_26883,N_26722);
xnor U27220 (N_27220,N_26544,N_26991);
or U27221 (N_27221,N_26705,N_26952);
nand U27222 (N_27222,N_26730,N_26980);
xor U27223 (N_27223,N_26629,N_26632);
xnor U27224 (N_27224,N_26527,N_26546);
nor U27225 (N_27225,N_26697,N_26537);
or U27226 (N_27226,N_26474,N_26913);
nor U27227 (N_27227,N_26877,N_26856);
or U27228 (N_27228,N_26656,N_26709);
xor U27229 (N_27229,N_26598,N_26900);
nand U27230 (N_27230,N_26750,N_26514);
nor U27231 (N_27231,N_26560,N_26986);
nor U27232 (N_27232,N_26993,N_26500);
nand U27233 (N_27233,N_26563,N_26428);
xnor U27234 (N_27234,N_26523,N_26655);
and U27235 (N_27235,N_26721,N_26772);
nor U27236 (N_27236,N_26504,N_26876);
nand U27237 (N_27237,N_26483,N_26777);
xor U27238 (N_27238,N_26831,N_26414);
and U27239 (N_27239,N_26675,N_26786);
xnor U27240 (N_27240,N_26662,N_26586);
or U27241 (N_27241,N_26645,N_26434);
nand U27242 (N_27242,N_26815,N_26545);
nor U27243 (N_27243,N_26677,N_26588);
or U27244 (N_27244,N_26460,N_26459);
and U27245 (N_27245,N_26572,N_26862);
nand U27246 (N_27246,N_26486,N_26956);
nand U27247 (N_27247,N_26686,N_26403);
xnor U27248 (N_27248,N_26605,N_26440);
xor U27249 (N_27249,N_26773,N_26907);
xnor U27250 (N_27250,N_26804,N_26635);
nand U27251 (N_27251,N_26756,N_26522);
nand U27252 (N_27252,N_26524,N_26529);
nor U27253 (N_27253,N_26832,N_26977);
or U27254 (N_27254,N_26799,N_26989);
xor U27255 (N_27255,N_26624,N_26470);
nand U27256 (N_27256,N_26811,N_26797);
or U27257 (N_27257,N_26408,N_26495);
nor U27258 (N_27258,N_26404,N_26601);
nand U27259 (N_27259,N_26571,N_26698);
nand U27260 (N_27260,N_26902,N_26468);
and U27261 (N_27261,N_26456,N_26599);
or U27262 (N_27262,N_26898,N_26729);
nor U27263 (N_27263,N_26800,N_26547);
xnor U27264 (N_27264,N_26937,N_26553);
nor U27265 (N_27265,N_26630,N_26882);
xor U27266 (N_27266,N_26904,N_26595);
nand U27267 (N_27267,N_26969,N_26858);
nor U27268 (N_27268,N_26673,N_26910);
or U27269 (N_27269,N_26432,N_26970);
nor U27270 (N_27270,N_26584,N_26921);
nor U27271 (N_27271,N_26696,N_26716);
xor U27272 (N_27272,N_26996,N_26781);
xor U27273 (N_27273,N_26784,N_26573);
or U27274 (N_27274,N_26608,N_26973);
nor U27275 (N_27275,N_26934,N_26735);
or U27276 (N_27276,N_26439,N_26920);
nand U27277 (N_27277,N_26992,N_26796);
nand U27278 (N_27278,N_26566,N_26837);
xnor U27279 (N_27279,N_26714,N_26918);
nor U27280 (N_27280,N_26834,N_26814);
and U27281 (N_27281,N_26878,N_26768);
xnor U27282 (N_27282,N_26954,N_26685);
nand U27283 (N_27283,N_26859,N_26695);
nand U27284 (N_27284,N_26983,N_26742);
nor U27285 (N_27285,N_26423,N_26507);
nand U27286 (N_27286,N_26603,N_26464);
or U27287 (N_27287,N_26816,N_26619);
xor U27288 (N_27288,N_26825,N_26967);
nand U27289 (N_27289,N_26590,N_26515);
and U27290 (N_27290,N_26610,N_26733);
or U27291 (N_27291,N_26438,N_26699);
or U27292 (N_27292,N_26613,N_26787);
nand U27293 (N_27293,N_26894,N_26840);
or U27294 (N_27294,N_26914,N_26968);
nor U27295 (N_27295,N_26532,N_26420);
or U27296 (N_27296,N_26580,N_26780);
or U27297 (N_27297,N_26961,N_26985);
nor U27298 (N_27298,N_26779,N_26974);
or U27299 (N_27299,N_26823,N_26562);
or U27300 (N_27300,N_26685,N_26910);
nor U27301 (N_27301,N_26603,N_26840);
xnor U27302 (N_27302,N_26486,N_26531);
or U27303 (N_27303,N_26592,N_26693);
or U27304 (N_27304,N_26713,N_26417);
xor U27305 (N_27305,N_26918,N_26897);
nor U27306 (N_27306,N_26759,N_26680);
nor U27307 (N_27307,N_26838,N_26538);
xor U27308 (N_27308,N_26853,N_26463);
or U27309 (N_27309,N_26877,N_26638);
nor U27310 (N_27310,N_26493,N_26512);
or U27311 (N_27311,N_26768,N_26503);
xor U27312 (N_27312,N_26635,N_26509);
or U27313 (N_27313,N_26643,N_26923);
nand U27314 (N_27314,N_26628,N_26679);
xor U27315 (N_27315,N_26997,N_26871);
or U27316 (N_27316,N_26630,N_26784);
xnor U27317 (N_27317,N_26853,N_26953);
xor U27318 (N_27318,N_26907,N_26723);
nor U27319 (N_27319,N_26538,N_26463);
xnor U27320 (N_27320,N_26943,N_26579);
xor U27321 (N_27321,N_26430,N_26909);
xor U27322 (N_27322,N_26524,N_26873);
or U27323 (N_27323,N_26429,N_26867);
or U27324 (N_27324,N_26634,N_26780);
nand U27325 (N_27325,N_26541,N_26932);
and U27326 (N_27326,N_26598,N_26476);
and U27327 (N_27327,N_26464,N_26949);
nand U27328 (N_27328,N_26438,N_26416);
xnor U27329 (N_27329,N_26832,N_26439);
nand U27330 (N_27330,N_26896,N_26634);
xnor U27331 (N_27331,N_26770,N_26502);
and U27332 (N_27332,N_26432,N_26992);
nand U27333 (N_27333,N_26758,N_26940);
or U27334 (N_27334,N_26604,N_26545);
nor U27335 (N_27335,N_26846,N_26949);
xnor U27336 (N_27336,N_26894,N_26479);
and U27337 (N_27337,N_26776,N_26948);
nor U27338 (N_27338,N_26704,N_26869);
nand U27339 (N_27339,N_26850,N_26721);
and U27340 (N_27340,N_26919,N_26976);
or U27341 (N_27341,N_26877,N_26640);
or U27342 (N_27342,N_26579,N_26881);
xor U27343 (N_27343,N_26572,N_26567);
or U27344 (N_27344,N_26457,N_26528);
xor U27345 (N_27345,N_26492,N_26922);
xor U27346 (N_27346,N_26622,N_26773);
and U27347 (N_27347,N_26620,N_26632);
or U27348 (N_27348,N_26822,N_26924);
nor U27349 (N_27349,N_26706,N_26407);
nor U27350 (N_27350,N_26949,N_26867);
and U27351 (N_27351,N_26457,N_26894);
nor U27352 (N_27352,N_26950,N_26915);
xor U27353 (N_27353,N_26545,N_26500);
or U27354 (N_27354,N_26427,N_26778);
nor U27355 (N_27355,N_26823,N_26470);
nand U27356 (N_27356,N_26413,N_26857);
and U27357 (N_27357,N_26470,N_26999);
xor U27358 (N_27358,N_26463,N_26740);
and U27359 (N_27359,N_26705,N_26822);
nor U27360 (N_27360,N_26958,N_26480);
nand U27361 (N_27361,N_26897,N_26428);
and U27362 (N_27362,N_26648,N_26544);
or U27363 (N_27363,N_26752,N_26569);
xnor U27364 (N_27364,N_26405,N_26874);
xnor U27365 (N_27365,N_26511,N_26835);
and U27366 (N_27366,N_26586,N_26749);
nor U27367 (N_27367,N_26526,N_26643);
xor U27368 (N_27368,N_26453,N_26918);
or U27369 (N_27369,N_26551,N_26466);
nor U27370 (N_27370,N_26760,N_26474);
xor U27371 (N_27371,N_26565,N_26569);
and U27372 (N_27372,N_26546,N_26483);
and U27373 (N_27373,N_26692,N_26420);
or U27374 (N_27374,N_26554,N_26559);
nand U27375 (N_27375,N_26791,N_26531);
or U27376 (N_27376,N_26954,N_26955);
nand U27377 (N_27377,N_26883,N_26643);
and U27378 (N_27378,N_26436,N_26667);
and U27379 (N_27379,N_26705,N_26662);
or U27380 (N_27380,N_26978,N_26484);
nor U27381 (N_27381,N_26580,N_26932);
and U27382 (N_27382,N_26748,N_26657);
nand U27383 (N_27383,N_26743,N_26568);
nor U27384 (N_27384,N_26428,N_26430);
nor U27385 (N_27385,N_26433,N_26692);
nor U27386 (N_27386,N_26688,N_26673);
and U27387 (N_27387,N_26628,N_26479);
nand U27388 (N_27388,N_26937,N_26472);
nor U27389 (N_27389,N_26464,N_26978);
nor U27390 (N_27390,N_26406,N_26756);
nor U27391 (N_27391,N_26800,N_26467);
and U27392 (N_27392,N_26442,N_26698);
xnor U27393 (N_27393,N_26498,N_26583);
nand U27394 (N_27394,N_26956,N_26869);
nor U27395 (N_27395,N_26681,N_26629);
xor U27396 (N_27396,N_26908,N_26720);
and U27397 (N_27397,N_26942,N_26888);
and U27398 (N_27398,N_26524,N_26890);
xor U27399 (N_27399,N_26855,N_26963);
xnor U27400 (N_27400,N_26696,N_26782);
nor U27401 (N_27401,N_26919,N_26565);
nor U27402 (N_27402,N_26943,N_26960);
nand U27403 (N_27403,N_26427,N_26520);
or U27404 (N_27404,N_26998,N_26928);
nor U27405 (N_27405,N_26662,N_26804);
and U27406 (N_27406,N_26455,N_26402);
or U27407 (N_27407,N_26540,N_26677);
nor U27408 (N_27408,N_26945,N_26607);
nor U27409 (N_27409,N_26793,N_26805);
or U27410 (N_27410,N_26702,N_26424);
or U27411 (N_27411,N_26457,N_26701);
nand U27412 (N_27412,N_26777,N_26752);
or U27413 (N_27413,N_26866,N_26452);
or U27414 (N_27414,N_26548,N_26563);
and U27415 (N_27415,N_26497,N_26619);
nand U27416 (N_27416,N_26877,N_26522);
nor U27417 (N_27417,N_26551,N_26701);
xor U27418 (N_27418,N_26989,N_26742);
nand U27419 (N_27419,N_26455,N_26912);
xnor U27420 (N_27420,N_26665,N_26916);
nand U27421 (N_27421,N_26962,N_26706);
xnor U27422 (N_27422,N_26860,N_26479);
nand U27423 (N_27423,N_26860,N_26601);
and U27424 (N_27424,N_26697,N_26674);
xor U27425 (N_27425,N_26544,N_26416);
or U27426 (N_27426,N_26896,N_26994);
or U27427 (N_27427,N_26912,N_26608);
and U27428 (N_27428,N_26534,N_26562);
or U27429 (N_27429,N_26842,N_26715);
or U27430 (N_27430,N_26852,N_26696);
xnor U27431 (N_27431,N_26623,N_26753);
nor U27432 (N_27432,N_26611,N_26705);
nor U27433 (N_27433,N_26875,N_26786);
xor U27434 (N_27434,N_26471,N_26633);
and U27435 (N_27435,N_26849,N_26965);
and U27436 (N_27436,N_26992,N_26553);
nor U27437 (N_27437,N_26532,N_26499);
nor U27438 (N_27438,N_26975,N_26639);
and U27439 (N_27439,N_26502,N_26976);
and U27440 (N_27440,N_26537,N_26789);
nand U27441 (N_27441,N_26783,N_26851);
nand U27442 (N_27442,N_26979,N_26822);
and U27443 (N_27443,N_26489,N_26767);
xnor U27444 (N_27444,N_26730,N_26764);
nand U27445 (N_27445,N_26671,N_26925);
xor U27446 (N_27446,N_26980,N_26940);
nand U27447 (N_27447,N_26943,N_26583);
or U27448 (N_27448,N_26648,N_26911);
nor U27449 (N_27449,N_26922,N_26993);
or U27450 (N_27450,N_26482,N_26602);
nor U27451 (N_27451,N_26665,N_26739);
nand U27452 (N_27452,N_26515,N_26849);
nor U27453 (N_27453,N_26441,N_26610);
nor U27454 (N_27454,N_26478,N_26944);
nor U27455 (N_27455,N_26456,N_26704);
or U27456 (N_27456,N_26420,N_26845);
nand U27457 (N_27457,N_26678,N_26505);
nor U27458 (N_27458,N_26563,N_26701);
or U27459 (N_27459,N_26448,N_26624);
or U27460 (N_27460,N_26876,N_26411);
and U27461 (N_27461,N_26965,N_26991);
nand U27462 (N_27462,N_26706,N_26690);
or U27463 (N_27463,N_26944,N_26740);
nand U27464 (N_27464,N_26881,N_26643);
nand U27465 (N_27465,N_26633,N_26840);
nand U27466 (N_27466,N_26820,N_26586);
nor U27467 (N_27467,N_26673,N_26654);
nand U27468 (N_27468,N_26455,N_26910);
nand U27469 (N_27469,N_26849,N_26845);
nand U27470 (N_27470,N_26606,N_26857);
nor U27471 (N_27471,N_26550,N_26695);
or U27472 (N_27472,N_26982,N_26677);
xor U27473 (N_27473,N_26961,N_26808);
xnor U27474 (N_27474,N_26670,N_26830);
or U27475 (N_27475,N_26694,N_26731);
and U27476 (N_27476,N_26964,N_26479);
xor U27477 (N_27477,N_26843,N_26732);
or U27478 (N_27478,N_26872,N_26491);
xnor U27479 (N_27479,N_26592,N_26975);
nand U27480 (N_27480,N_26441,N_26685);
xor U27481 (N_27481,N_26596,N_26580);
nor U27482 (N_27482,N_26438,N_26478);
or U27483 (N_27483,N_26877,N_26973);
or U27484 (N_27484,N_26776,N_26686);
or U27485 (N_27485,N_26905,N_26588);
or U27486 (N_27486,N_26902,N_26910);
nand U27487 (N_27487,N_26695,N_26493);
and U27488 (N_27488,N_26972,N_26928);
nand U27489 (N_27489,N_26921,N_26922);
xor U27490 (N_27490,N_26676,N_26767);
or U27491 (N_27491,N_26606,N_26576);
nand U27492 (N_27492,N_26745,N_26845);
or U27493 (N_27493,N_26472,N_26731);
nor U27494 (N_27494,N_26953,N_26607);
or U27495 (N_27495,N_26721,N_26963);
and U27496 (N_27496,N_26543,N_26496);
nand U27497 (N_27497,N_26854,N_26936);
and U27498 (N_27498,N_26408,N_26671);
nand U27499 (N_27499,N_26637,N_26782);
nor U27500 (N_27500,N_26884,N_26810);
and U27501 (N_27501,N_26692,N_26982);
and U27502 (N_27502,N_26836,N_26781);
nand U27503 (N_27503,N_26853,N_26563);
nor U27504 (N_27504,N_26979,N_26897);
and U27505 (N_27505,N_26596,N_26481);
and U27506 (N_27506,N_26807,N_26460);
nor U27507 (N_27507,N_26646,N_26541);
xor U27508 (N_27508,N_26614,N_26667);
or U27509 (N_27509,N_26809,N_26733);
nor U27510 (N_27510,N_26739,N_26988);
xor U27511 (N_27511,N_26457,N_26478);
and U27512 (N_27512,N_26669,N_26574);
nor U27513 (N_27513,N_26528,N_26549);
nand U27514 (N_27514,N_26938,N_26652);
nor U27515 (N_27515,N_26755,N_26449);
xnor U27516 (N_27516,N_26402,N_26978);
xor U27517 (N_27517,N_26633,N_26765);
and U27518 (N_27518,N_26470,N_26538);
nor U27519 (N_27519,N_26869,N_26459);
nor U27520 (N_27520,N_26866,N_26789);
xor U27521 (N_27521,N_26498,N_26997);
nor U27522 (N_27522,N_26604,N_26811);
nand U27523 (N_27523,N_26801,N_26714);
xor U27524 (N_27524,N_26753,N_26553);
nor U27525 (N_27525,N_26921,N_26413);
nand U27526 (N_27526,N_26945,N_26491);
xnor U27527 (N_27527,N_26921,N_26581);
nor U27528 (N_27528,N_26510,N_26736);
and U27529 (N_27529,N_26921,N_26443);
xnor U27530 (N_27530,N_26587,N_26702);
and U27531 (N_27531,N_26813,N_26971);
or U27532 (N_27532,N_26818,N_26491);
or U27533 (N_27533,N_26701,N_26892);
xnor U27534 (N_27534,N_26618,N_26937);
nor U27535 (N_27535,N_26541,N_26470);
nand U27536 (N_27536,N_26605,N_26830);
and U27537 (N_27537,N_26898,N_26668);
or U27538 (N_27538,N_26627,N_26688);
and U27539 (N_27539,N_26688,N_26928);
or U27540 (N_27540,N_26437,N_26634);
nor U27541 (N_27541,N_26724,N_26958);
xnor U27542 (N_27542,N_26854,N_26619);
xor U27543 (N_27543,N_26698,N_26965);
and U27544 (N_27544,N_26442,N_26403);
nand U27545 (N_27545,N_26659,N_26906);
and U27546 (N_27546,N_26521,N_26504);
nor U27547 (N_27547,N_26475,N_26516);
xnor U27548 (N_27548,N_26604,N_26999);
and U27549 (N_27549,N_26667,N_26771);
or U27550 (N_27550,N_26475,N_26910);
nor U27551 (N_27551,N_26550,N_26504);
nand U27552 (N_27552,N_26489,N_26966);
nand U27553 (N_27553,N_26644,N_26639);
xnor U27554 (N_27554,N_26461,N_26524);
and U27555 (N_27555,N_26404,N_26506);
nor U27556 (N_27556,N_26748,N_26848);
nand U27557 (N_27557,N_26883,N_26929);
xor U27558 (N_27558,N_26771,N_26902);
nand U27559 (N_27559,N_26954,N_26501);
or U27560 (N_27560,N_26549,N_26739);
nand U27561 (N_27561,N_26696,N_26829);
and U27562 (N_27562,N_26637,N_26618);
xor U27563 (N_27563,N_26511,N_26867);
nand U27564 (N_27564,N_26642,N_26400);
or U27565 (N_27565,N_26701,N_26858);
nor U27566 (N_27566,N_26797,N_26837);
nand U27567 (N_27567,N_26506,N_26916);
nand U27568 (N_27568,N_26473,N_26753);
and U27569 (N_27569,N_26693,N_26935);
nor U27570 (N_27570,N_26897,N_26429);
xor U27571 (N_27571,N_26416,N_26976);
xor U27572 (N_27572,N_26463,N_26728);
and U27573 (N_27573,N_26555,N_26609);
or U27574 (N_27574,N_26608,N_26851);
xor U27575 (N_27575,N_26444,N_26503);
and U27576 (N_27576,N_26464,N_26675);
nor U27577 (N_27577,N_26727,N_26870);
nand U27578 (N_27578,N_26992,N_26873);
and U27579 (N_27579,N_26426,N_26975);
nor U27580 (N_27580,N_26458,N_26664);
xnor U27581 (N_27581,N_26506,N_26419);
xor U27582 (N_27582,N_26910,N_26706);
nor U27583 (N_27583,N_26494,N_26414);
nor U27584 (N_27584,N_26589,N_26498);
or U27585 (N_27585,N_26608,N_26765);
and U27586 (N_27586,N_26940,N_26989);
nand U27587 (N_27587,N_26599,N_26872);
or U27588 (N_27588,N_26724,N_26462);
or U27589 (N_27589,N_26436,N_26857);
and U27590 (N_27590,N_26919,N_26548);
nand U27591 (N_27591,N_26769,N_26592);
nand U27592 (N_27592,N_26803,N_26506);
xor U27593 (N_27593,N_26627,N_26508);
and U27594 (N_27594,N_26795,N_26560);
xnor U27595 (N_27595,N_26611,N_26502);
and U27596 (N_27596,N_26721,N_26813);
nor U27597 (N_27597,N_26724,N_26651);
xnor U27598 (N_27598,N_26946,N_26971);
nand U27599 (N_27599,N_26588,N_26839);
and U27600 (N_27600,N_27267,N_27196);
or U27601 (N_27601,N_27249,N_27154);
or U27602 (N_27602,N_27318,N_27399);
xor U27603 (N_27603,N_27537,N_27026);
and U27604 (N_27604,N_27572,N_27522);
nor U27605 (N_27605,N_27342,N_27588);
nor U27606 (N_27606,N_27083,N_27103);
nor U27607 (N_27607,N_27218,N_27570);
nand U27608 (N_27608,N_27238,N_27430);
or U27609 (N_27609,N_27304,N_27346);
xor U27610 (N_27610,N_27118,N_27356);
and U27611 (N_27611,N_27289,N_27428);
nand U27612 (N_27612,N_27112,N_27021);
and U27613 (N_27613,N_27188,N_27373);
or U27614 (N_27614,N_27000,N_27398);
and U27615 (N_27615,N_27234,N_27444);
nor U27616 (N_27616,N_27183,N_27578);
or U27617 (N_27617,N_27278,N_27003);
nand U27618 (N_27618,N_27546,N_27458);
and U27619 (N_27619,N_27394,N_27055);
xor U27620 (N_27620,N_27284,N_27493);
or U27621 (N_27621,N_27053,N_27349);
nand U27622 (N_27622,N_27038,N_27464);
and U27623 (N_27623,N_27479,N_27224);
xor U27624 (N_27624,N_27301,N_27380);
nor U27625 (N_27625,N_27169,N_27475);
xnor U27626 (N_27626,N_27147,N_27175);
and U27627 (N_27627,N_27040,N_27060);
xnor U27628 (N_27628,N_27483,N_27311);
nor U27629 (N_27629,N_27240,N_27269);
xor U27630 (N_27630,N_27592,N_27363);
nand U27631 (N_27631,N_27273,N_27037);
or U27632 (N_27632,N_27200,N_27160);
and U27633 (N_27633,N_27272,N_27085);
xor U27634 (N_27634,N_27137,N_27396);
and U27635 (N_27635,N_27437,N_27534);
or U27636 (N_27636,N_27128,N_27164);
xnor U27637 (N_27637,N_27533,N_27443);
or U27638 (N_27638,N_27386,N_27331);
nor U27639 (N_27639,N_27321,N_27024);
xor U27640 (N_27640,N_27333,N_27462);
or U27641 (N_27641,N_27012,N_27456);
and U27642 (N_27642,N_27410,N_27292);
and U27643 (N_27643,N_27302,N_27006);
nor U27644 (N_27644,N_27193,N_27189);
nor U27645 (N_27645,N_27376,N_27436);
and U27646 (N_27646,N_27484,N_27498);
nand U27647 (N_27647,N_27497,N_27069);
xnor U27648 (N_27648,N_27126,N_27113);
xor U27649 (N_27649,N_27288,N_27583);
nor U27650 (N_27650,N_27477,N_27567);
and U27651 (N_27651,N_27461,N_27305);
or U27652 (N_27652,N_27553,N_27448);
xor U27653 (N_27653,N_27178,N_27098);
and U27654 (N_27654,N_27313,N_27229);
xor U27655 (N_27655,N_27097,N_27576);
and U27656 (N_27656,N_27020,N_27170);
or U27657 (N_27657,N_27237,N_27157);
xor U27658 (N_27658,N_27133,N_27540);
or U27659 (N_27659,N_27018,N_27110);
xnor U27660 (N_27660,N_27243,N_27381);
and U27661 (N_27661,N_27545,N_27127);
nor U27662 (N_27662,N_27139,N_27491);
and U27663 (N_27663,N_27210,N_27090);
or U27664 (N_27664,N_27595,N_27582);
and U27665 (N_27665,N_27262,N_27556);
nor U27666 (N_27666,N_27338,N_27208);
and U27667 (N_27667,N_27418,N_27174);
nand U27668 (N_27668,N_27259,N_27368);
nor U27669 (N_27669,N_27403,N_27030);
nand U27670 (N_27670,N_27153,N_27408);
nor U27671 (N_27671,N_27124,N_27334);
xor U27672 (N_27672,N_27426,N_27283);
nand U27673 (N_27673,N_27370,N_27463);
xnor U27674 (N_27674,N_27106,N_27514);
nand U27675 (N_27675,N_27511,N_27599);
or U27676 (N_27676,N_27114,N_27045);
xnor U27677 (N_27677,N_27389,N_27447);
nand U27678 (N_27678,N_27395,N_27379);
xnor U27679 (N_27679,N_27494,N_27587);
nand U27680 (N_27680,N_27427,N_27422);
xnor U27681 (N_27681,N_27235,N_27270);
or U27682 (N_27682,N_27049,N_27315);
and U27683 (N_27683,N_27508,N_27415);
or U27684 (N_27684,N_27168,N_27074);
nand U27685 (N_27685,N_27316,N_27505);
xnor U27686 (N_27686,N_27266,N_27451);
xnor U27687 (N_27687,N_27034,N_27227);
xnor U27688 (N_27688,N_27594,N_27228);
nand U27689 (N_27689,N_27192,N_27405);
nand U27690 (N_27690,N_27590,N_27521);
or U27691 (N_27691,N_27271,N_27579);
nor U27692 (N_27692,N_27375,N_27165);
and U27693 (N_27693,N_27423,N_27470);
nor U27694 (N_27694,N_27080,N_27219);
or U27695 (N_27695,N_27166,N_27059);
and U27696 (N_27696,N_27377,N_27032);
or U27697 (N_27697,N_27144,N_27258);
and U27698 (N_27698,N_27041,N_27028);
and U27699 (N_27699,N_27509,N_27528);
nor U27700 (N_27700,N_27312,N_27467);
nand U27701 (N_27701,N_27217,N_27432);
nand U27702 (N_27702,N_27440,N_27205);
or U27703 (N_27703,N_27094,N_27061);
nand U27704 (N_27704,N_27009,N_27323);
nand U27705 (N_27705,N_27145,N_27541);
xor U27706 (N_27706,N_27075,N_27568);
nand U27707 (N_27707,N_27487,N_27010);
and U27708 (N_27708,N_27455,N_27435);
and U27709 (N_27709,N_27029,N_27067);
and U27710 (N_27710,N_27337,N_27476);
or U27711 (N_27711,N_27092,N_27383);
nor U27712 (N_27712,N_27387,N_27099);
xnor U27713 (N_27713,N_27581,N_27317);
nand U27714 (N_27714,N_27152,N_27295);
xor U27715 (N_27715,N_27364,N_27185);
and U27716 (N_27716,N_27148,N_27176);
nor U27717 (N_27717,N_27136,N_27179);
nand U27718 (N_27718,N_27204,N_27241);
nor U27719 (N_27719,N_27485,N_27253);
nor U27720 (N_27720,N_27186,N_27566);
xnor U27721 (N_27721,N_27504,N_27257);
xnor U27722 (N_27722,N_27560,N_27182);
nor U27723 (N_27723,N_27369,N_27431);
and U27724 (N_27724,N_27231,N_27008);
xnor U27725 (N_27725,N_27328,N_27254);
and U27726 (N_27726,N_27402,N_27524);
nand U27727 (N_27727,N_27255,N_27523);
nor U27728 (N_27728,N_27209,N_27197);
or U27729 (N_27729,N_27088,N_27223);
nor U27730 (N_27730,N_27282,N_27500);
nor U27731 (N_27731,N_27093,N_27057);
xor U27732 (N_27732,N_27052,N_27158);
xnor U27733 (N_27733,N_27551,N_27274);
or U27734 (N_27734,N_27544,N_27480);
and U27735 (N_27735,N_27181,N_27575);
or U27736 (N_27736,N_27388,N_27344);
or U27737 (N_27737,N_27471,N_27486);
nor U27738 (N_27738,N_27416,N_27236);
or U27739 (N_27739,N_27107,N_27539);
or U27740 (N_27740,N_27125,N_27033);
and U27741 (N_27741,N_27299,N_27354);
nand U27742 (N_27742,N_27076,N_27340);
and U27743 (N_27743,N_27216,N_27367);
nor U27744 (N_27744,N_27362,N_27132);
nor U27745 (N_27745,N_27314,N_27279);
and U27746 (N_27746,N_27105,N_27332);
nor U27747 (N_27747,N_27047,N_27489);
xor U27748 (N_27748,N_27120,N_27413);
xnor U27749 (N_27749,N_27225,N_27457);
xor U27750 (N_27750,N_27100,N_27374);
xnor U27751 (N_27751,N_27438,N_27382);
nor U27752 (N_27752,N_27345,N_27251);
and U27753 (N_27753,N_27087,N_27122);
and U27754 (N_27754,N_27096,N_27529);
nand U27755 (N_27755,N_27220,N_27056);
nor U27756 (N_27756,N_27535,N_27180);
or U27757 (N_27757,N_27355,N_27372);
nand U27758 (N_27758,N_27163,N_27330);
and U27759 (N_27759,N_27177,N_27239);
nor U27760 (N_27760,N_27559,N_27135);
xor U27761 (N_27761,N_27261,N_27488);
nor U27762 (N_27762,N_27101,N_27482);
nor U27763 (N_27763,N_27411,N_27525);
or U27764 (N_27764,N_27063,N_27361);
and U27765 (N_27765,N_27326,N_27002);
xor U27766 (N_27766,N_27420,N_27242);
and U27767 (N_27767,N_27391,N_27536);
nand U27768 (N_27768,N_27138,N_27111);
xor U27769 (N_27769,N_27256,N_27001);
xor U27770 (N_27770,N_27213,N_27401);
xnor U27771 (N_27771,N_27348,N_27459);
xnor U27772 (N_27772,N_27442,N_27407);
or U27773 (N_27773,N_27425,N_27390);
xnor U27774 (N_27774,N_27571,N_27460);
xnor U27775 (N_27775,N_27450,N_27468);
nand U27776 (N_27776,N_27065,N_27184);
and U27777 (N_27777,N_27079,N_27286);
and U27778 (N_27778,N_27466,N_27247);
nand U27779 (N_27779,N_27134,N_27336);
nand U27780 (N_27780,N_27226,N_27058);
xnor U27781 (N_27781,N_27327,N_27140);
xor U27782 (N_27782,N_27531,N_27538);
nor U27783 (N_27783,N_27445,N_27048);
nand U27784 (N_27784,N_27473,N_27378);
nand U27785 (N_27785,N_27573,N_27025);
nand U27786 (N_27786,N_27171,N_27516);
or U27787 (N_27787,N_27146,N_27296);
and U27788 (N_27788,N_27042,N_27062);
nor U27789 (N_27789,N_27404,N_27195);
nor U27790 (N_27790,N_27517,N_27050);
or U27791 (N_27791,N_27357,N_27406);
and U27792 (N_27792,N_27064,N_27142);
nor U27793 (N_27793,N_27151,N_27206);
xor U27794 (N_27794,N_27481,N_27584);
or U27795 (N_27795,N_27141,N_27117);
xor U27796 (N_27796,N_27591,N_27202);
and U27797 (N_27797,N_27597,N_27596);
or U27798 (N_27798,N_27071,N_27417);
nand U27799 (N_27799,N_27512,N_27248);
and U27800 (N_27800,N_27108,N_27194);
xor U27801 (N_27801,N_27414,N_27421);
xor U27802 (N_27802,N_27066,N_27172);
nor U27803 (N_27803,N_27232,N_27469);
nor U27804 (N_27804,N_27550,N_27082);
or U27805 (N_27805,N_27474,N_27358);
nor U27806 (N_27806,N_27054,N_27123);
xor U27807 (N_27807,N_27077,N_27078);
nor U27808 (N_27808,N_27293,N_27518);
or U27809 (N_27809,N_27084,N_27412);
nor U27810 (N_27810,N_27023,N_27173);
nand U27811 (N_27811,N_27320,N_27046);
or U27812 (N_27812,N_27548,N_27569);
nor U27813 (N_27813,N_27397,N_27385);
nand U27814 (N_27814,N_27441,N_27297);
and U27815 (N_27815,N_27563,N_27351);
and U27816 (N_27816,N_27530,N_27547);
nand U27817 (N_27817,N_27562,N_27353);
nand U27818 (N_27818,N_27501,N_27439);
and U27819 (N_27819,N_27306,N_27260);
nor U27820 (N_27820,N_27091,N_27005);
xnor U27821 (N_27821,N_27446,N_27580);
nor U27822 (N_27822,N_27419,N_27324);
nand U27823 (N_27823,N_27507,N_27513);
or U27824 (N_27824,N_27285,N_27086);
nand U27825 (N_27825,N_27519,N_27325);
xnor U27826 (N_27826,N_27424,N_27263);
xor U27827 (N_27827,N_27492,N_27233);
and U27828 (N_27828,N_27156,N_27070);
xnor U27829 (N_27829,N_27207,N_27198);
or U27830 (N_27830,N_27212,N_27250);
or U27831 (N_27831,N_27400,N_27268);
or U27832 (N_27832,N_27554,N_27309);
xor U27833 (N_27833,N_27072,N_27557);
nor U27834 (N_27834,N_27287,N_27359);
or U27835 (N_27835,N_27503,N_27201);
nand U27836 (N_27836,N_27121,N_27453);
nor U27837 (N_27837,N_27454,N_27520);
and U27838 (N_27838,N_27161,N_27019);
nor U27839 (N_27839,N_27490,N_27496);
and U27840 (N_27840,N_27167,N_27561);
nor U27841 (N_27841,N_27130,N_27280);
or U27842 (N_27842,N_27300,N_27015);
or U27843 (N_27843,N_27319,N_27119);
xor U27844 (N_27844,N_27499,N_27203);
nand U27845 (N_27845,N_27007,N_27199);
xor U27846 (N_27846,N_27221,N_27598);
nand U27847 (N_27847,N_27162,N_27542);
nand U27848 (N_27848,N_27478,N_27068);
xor U27849 (N_27849,N_27035,N_27392);
and U27850 (N_27850,N_27366,N_27095);
xor U27851 (N_27851,N_27244,N_27290);
nor U27852 (N_27852,N_27409,N_27190);
nand U27853 (N_27853,N_27036,N_27433);
and U27854 (N_27854,N_27039,N_27043);
nor U27855 (N_27855,N_27429,N_27465);
and U27856 (N_27856,N_27215,N_27527);
xor U27857 (N_27857,N_27564,N_27434);
nand U27858 (N_27858,N_27129,N_27371);
xor U27859 (N_27859,N_27187,N_27495);
and U27860 (N_27860,N_27281,N_27150);
nor U27861 (N_27861,N_27452,N_27502);
and U27862 (N_27862,N_27384,N_27155);
nand U27863 (N_27863,N_27360,N_27565);
and U27864 (N_27864,N_27276,N_27222);
nor U27865 (N_27865,N_27277,N_27245);
nor U27866 (N_27866,N_27149,N_27308);
nor U27867 (N_27867,N_27109,N_27044);
or U27868 (N_27868,N_27365,N_27011);
and U27869 (N_27869,N_27073,N_27089);
or U27870 (N_27870,N_27586,N_27294);
and U27871 (N_27871,N_27343,N_27027);
xor U27872 (N_27872,N_27593,N_27552);
nor U27873 (N_27873,N_27051,N_27214);
xnor U27874 (N_27874,N_27555,N_27303);
and U27875 (N_27875,N_27472,N_27131);
or U27876 (N_27876,N_27307,N_27014);
or U27877 (N_27877,N_27246,N_27339);
xor U27878 (N_27878,N_27574,N_27115);
or U27879 (N_27879,N_27104,N_27510);
nor U27880 (N_27880,N_27449,N_27393);
and U27881 (N_27881,N_27532,N_27275);
or U27882 (N_27882,N_27143,N_27017);
and U27883 (N_27883,N_27031,N_27322);
nor U27884 (N_27884,N_27310,N_27102);
nor U27885 (N_27885,N_27335,N_27081);
nor U27886 (N_27886,N_27291,N_27230);
nor U27887 (N_27887,N_27589,N_27577);
nand U27888 (N_27888,N_27264,N_27543);
nor U27889 (N_27889,N_27252,N_27329);
and U27890 (N_27890,N_27016,N_27022);
or U27891 (N_27891,N_27585,N_27526);
and U27892 (N_27892,N_27298,N_27347);
nor U27893 (N_27893,N_27013,N_27350);
nand U27894 (N_27894,N_27558,N_27352);
and U27895 (N_27895,N_27506,N_27549);
and U27896 (N_27896,N_27116,N_27341);
xnor U27897 (N_27897,N_27265,N_27211);
nor U27898 (N_27898,N_27159,N_27191);
or U27899 (N_27899,N_27515,N_27004);
nand U27900 (N_27900,N_27478,N_27351);
or U27901 (N_27901,N_27319,N_27236);
or U27902 (N_27902,N_27188,N_27286);
xnor U27903 (N_27903,N_27435,N_27443);
or U27904 (N_27904,N_27342,N_27596);
xor U27905 (N_27905,N_27251,N_27273);
xnor U27906 (N_27906,N_27038,N_27398);
and U27907 (N_27907,N_27242,N_27098);
nand U27908 (N_27908,N_27082,N_27468);
nor U27909 (N_27909,N_27469,N_27445);
nand U27910 (N_27910,N_27488,N_27021);
xnor U27911 (N_27911,N_27183,N_27316);
nor U27912 (N_27912,N_27427,N_27226);
xor U27913 (N_27913,N_27592,N_27101);
or U27914 (N_27914,N_27105,N_27563);
nand U27915 (N_27915,N_27497,N_27522);
nor U27916 (N_27916,N_27584,N_27466);
nor U27917 (N_27917,N_27335,N_27494);
or U27918 (N_27918,N_27404,N_27572);
xor U27919 (N_27919,N_27114,N_27398);
nor U27920 (N_27920,N_27118,N_27162);
nand U27921 (N_27921,N_27153,N_27588);
nor U27922 (N_27922,N_27420,N_27570);
and U27923 (N_27923,N_27057,N_27070);
nand U27924 (N_27924,N_27579,N_27367);
nor U27925 (N_27925,N_27574,N_27571);
nand U27926 (N_27926,N_27368,N_27187);
or U27927 (N_27927,N_27278,N_27466);
or U27928 (N_27928,N_27417,N_27064);
nor U27929 (N_27929,N_27049,N_27334);
xnor U27930 (N_27930,N_27165,N_27029);
nor U27931 (N_27931,N_27159,N_27411);
nor U27932 (N_27932,N_27568,N_27291);
nand U27933 (N_27933,N_27205,N_27052);
nor U27934 (N_27934,N_27586,N_27025);
nor U27935 (N_27935,N_27137,N_27010);
xor U27936 (N_27936,N_27555,N_27424);
nand U27937 (N_27937,N_27526,N_27302);
nor U27938 (N_27938,N_27302,N_27247);
nand U27939 (N_27939,N_27102,N_27144);
xor U27940 (N_27940,N_27185,N_27515);
nor U27941 (N_27941,N_27533,N_27550);
nor U27942 (N_27942,N_27063,N_27416);
or U27943 (N_27943,N_27294,N_27098);
xor U27944 (N_27944,N_27049,N_27559);
or U27945 (N_27945,N_27507,N_27054);
and U27946 (N_27946,N_27306,N_27572);
or U27947 (N_27947,N_27361,N_27255);
and U27948 (N_27948,N_27478,N_27146);
or U27949 (N_27949,N_27515,N_27272);
nor U27950 (N_27950,N_27109,N_27140);
and U27951 (N_27951,N_27097,N_27358);
or U27952 (N_27952,N_27232,N_27502);
nor U27953 (N_27953,N_27385,N_27010);
and U27954 (N_27954,N_27361,N_27536);
nor U27955 (N_27955,N_27379,N_27492);
or U27956 (N_27956,N_27365,N_27524);
xor U27957 (N_27957,N_27125,N_27244);
nand U27958 (N_27958,N_27180,N_27431);
nor U27959 (N_27959,N_27504,N_27003);
or U27960 (N_27960,N_27186,N_27431);
and U27961 (N_27961,N_27481,N_27084);
and U27962 (N_27962,N_27311,N_27376);
nand U27963 (N_27963,N_27407,N_27473);
xor U27964 (N_27964,N_27158,N_27212);
xnor U27965 (N_27965,N_27454,N_27392);
nand U27966 (N_27966,N_27441,N_27581);
nor U27967 (N_27967,N_27535,N_27402);
and U27968 (N_27968,N_27049,N_27311);
nor U27969 (N_27969,N_27529,N_27108);
nor U27970 (N_27970,N_27559,N_27349);
nand U27971 (N_27971,N_27145,N_27095);
xor U27972 (N_27972,N_27459,N_27556);
nand U27973 (N_27973,N_27565,N_27473);
xor U27974 (N_27974,N_27312,N_27229);
nor U27975 (N_27975,N_27445,N_27120);
nand U27976 (N_27976,N_27469,N_27453);
and U27977 (N_27977,N_27120,N_27208);
xnor U27978 (N_27978,N_27131,N_27005);
and U27979 (N_27979,N_27105,N_27539);
nor U27980 (N_27980,N_27377,N_27169);
nor U27981 (N_27981,N_27219,N_27058);
nand U27982 (N_27982,N_27147,N_27558);
or U27983 (N_27983,N_27530,N_27464);
or U27984 (N_27984,N_27011,N_27344);
and U27985 (N_27985,N_27197,N_27336);
nor U27986 (N_27986,N_27562,N_27524);
and U27987 (N_27987,N_27267,N_27597);
xor U27988 (N_27988,N_27256,N_27581);
and U27989 (N_27989,N_27579,N_27034);
xnor U27990 (N_27990,N_27266,N_27444);
and U27991 (N_27991,N_27532,N_27337);
nand U27992 (N_27992,N_27444,N_27470);
or U27993 (N_27993,N_27268,N_27336);
or U27994 (N_27994,N_27103,N_27429);
and U27995 (N_27995,N_27210,N_27254);
or U27996 (N_27996,N_27418,N_27127);
nand U27997 (N_27997,N_27303,N_27517);
nand U27998 (N_27998,N_27067,N_27311);
or U27999 (N_27999,N_27179,N_27326);
nor U28000 (N_28000,N_27189,N_27085);
or U28001 (N_28001,N_27383,N_27592);
nand U28002 (N_28002,N_27013,N_27309);
and U28003 (N_28003,N_27457,N_27448);
nand U28004 (N_28004,N_27238,N_27384);
and U28005 (N_28005,N_27082,N_27544);
xor U28006 (N_28006,N_27062,N_27287);
nand U28007 (N_28007,N_27270,N_27404);
and U28008 (N_28008,N_27297,N_27541);
or U28009 (N_28009,N_27137,N_27015);
nand U28010 (N_28010,N_27307,N_27300);
xnor U28011 (N_28011,N_27041,N_27472);
and U28012 (N_28012,N_27572,N_27135);
xor U28013 (N_28013,N_27308,N_27145);
and U28014 (N_28014,N_27154,N_27518);
nand U28015 (N_28015,N_27138,N_27385);
and U28016 (N_28016,N_27044,N_27179);
nand U28017 (N_28017,N_27390,N_27165);
nand U28018 (N_28018,N_27305,N_27467);
nor U28019 (N_28019,N_27437,N_27268);
and U28020 (N_28020,N_27209,N_27248);
nor U28021 (N_28021,N_27067,N_27428);
or U28022 (N_28022,N_27126,N_27383);
xor U28023 (N_28023,N_27074,N_27446);
nor U28024 (N_28024,N_27017,N_27286);
nor U28025 (N_28025,N_27493,N_27300);
or U28026 (N_28026,N_27460,N_27023);
nand U28027 (N_28027,N_27168,N_27142);
nor U28028 (N_28028,N_27546,N_27281);
nand U28029 (N_28029,N_27209,N_27283);
and U28030 (N_28030,N_27071,N_27266);
nor U28031 (N_28031,N_27246,N_27070);
and U28032 (N_28032,N_27579,N_27583);
or U28033 (N_28033,N_27387,N_27552);
and U28034 (N_28034,N_27238,N_27447);
nand U28035 (N_28035,N_27036,N_27124);
nor U28036 (N_28036,N_27079,N_27024);
xnor U28037 (N_28037,N_27468,N_27493);
and U28038 (N_28038,N_27327,N_27188);
and U28039 (N_28039,N_27330,N_27104);
xor U28040 (N_28040,N_27209,N_27194);
nor U28041 (N_28041,N_27572,N_27548);
nand U28042 (N_28042,N_27234,N_27163);
nand U28043 (N_28043,N_27394,N_27517);
xor U28044 (N_28044,N_27312,N_27149);
nand U28045 (N_28045,N_27034,N_27166);
nor U28046 (N_28046,N_27384,N_27404);
xnor U28047 (N_28047,N_27181,N_27144);
nor U28048 (N_28048,N_27452,N_27565);
xor U28049 (N_28049,N_27589,N_27543);
and U28050 (N_28050,N_27039,N_27156);
and U28051 (N_28051,N_27541,N_27030);
xnor U28052 (N_28052,N_27034,N_27143);
nand U28053 (N_28053,N_27291,N_27338);
and U28054 (N_28054,N_27509,N_27151);
xnor U28055 (N_28055,N_27331,N_27306);
and U28056 (N_28056,N_27340,N_27557);
nand U28057 (N_28057,N_27495,N_27109);
nor U28058 (N_28058,N_27024,N_27542);
nor U28059 (N_28059,N_27415,N_27296);
or U28060 (N_28060,N_27092,N_27531);
or U28061 (N_28061,N_27174,N_27443);
nand U28062 (N_28062,N_27188,N_27208);
nor U28063 (N_28063,N_27151,N_27134);
and U28064 (N_28064,N_27425,N_27294);
or U28065 (N_28065,N_27579,N_27521);
xor U28066 (N_28066,N_27151,N_27414);
xor U28067 (N_28067,N_27345,N_27123);
xnor U28068 (N_28068,N_27529,N_27509);
or U28069 (N_28069,N_27336,N_27327);
nor U28070 (N_28070,N_27065,N_27330);
or U28071 (N_28071,N_27572,N_27067);
or U28072 (N_28072,N_27563,N_27056);
nor U28073 (N_28073,N_27268,N_27000);
nor U28074 (N_28074,N_27580,N_27196);
and U28075 (N_28075,N_27499,N_27056);
nand U28076 (N_28076,N_27445,N_27525);
xor U28077 (N_28077,N_27188,N_27246);
nand U28078 (N_28078,N_27294,N_27500);
nor U28079 (N_28079,N_27070,N_27305);
nor U28080 (N_28080,N_27443,N_27149);
or U28081 (N_28081,N_27069,N_27009);
nand U28082 (N_28082,N_27379,N_27479);
and U28083 (N_28083,N_27342,N_27195);
and U28084 (N_28084,N_27392,N_27512);
or U28085 (N_28085,N_27244,N_27527);
xnor U28086 (N_28086,N_27545,N_27476);
or U28087 (N_28087,N_27565,N_27460);
and U28088 (N_28088,N_27079,N_27360);
nor U28089 (N_28089,N_27208,N_27427);
or U28090 (N_28090,N_27076,N_27440);
and U28091 (N_28091,N_27353,N_27032);
nor U28092 (N_28092,N_27325,N_27341);
and U28093 (N_28093,N_27300,N_27020);
xnor U28094 (N_28094,N_27196,N_27519);
xnor U28095 (N_28095,N_27009,N_27282);
or U28096 (N_28096,N_27475,N_27405);
and U28097 (N_28097,N_27091,N_27186);
nand U28098 (N_28098,N_27095,N_27311);
nor U28099 (N_28099,N_27454,N_27564);
and U28100 (N_28100,N_27545,N_27566);
nand U28101 (N_28101,N_27117,N_27171);
or U28102 (N_28102,N_27540,N_27351);
or U28103 (N_28103,N_27485,N_27023);
nand U28104 (N_28104,N_27303,N_27533);
nor U28105 (N_28105,N_27372,N_27197);
nand U28106 (N_28106,N_27399,N_27231);
nor U28107 (N_28107,N_27296,N_27158);
or U28108 (N_28108,N_27131,N_27572);
nor U28109 (N_28109,N_27300,N_27321);
nor U28110 (N_28110,N_27019,N_27581);
nand U28111 (N_28111,N_27214,N_27556);
nand U28112 (N_28112,N_27533,N_27574);
or U28113 (N_28113,N_27125,N_27461);
xor U28114 (N_28114,N_27445,N_27240);
nor U28115 (N_28115,N_27238,N_27183);
nor U28116 (N_28116,N_27131,N_27464);
and U28117 (N_28117,N_27278,N_27162);
and U28118 (N_28118,N_27363,N_27000);
nor U28119 (N_28119,N_27057,N_27360);
nor U28120 (N_28120,N_27389,N_27346);
and U28121 (N_28121,N_27061,N_27077);
xnor U28122 (N_28122,N_27347,N_27531);
nand U28123 (N_28123,N_27487,N_27434);
nor U28124 (N_28124,N_27284,N_27040);
nor U28125 (N_28125,N_27584,N_27382);
or U28126 (N_28126,N_27007,N_27419);
nand U28127 (N_28127,N_27430,N_27594);
or U28128 (N_28128,N_27479,N_27292);
nand U28129 (N_28129,N_27599,N_27519);
and U28130 (N_28130,N_27351,N_27437);
xor U28131 (N_28131,N_27041,N_27067);
nor U28132 (N_28132,N_27103,N_27295);
or U28133 (N_28133,N_27238,N_27165);
nand U28134 (N_28134,N_27150,N_27539);
xor U28135 (N_28135,N_27040,N_27310);
xor U28136 (N_28136,N_27121,N_27265);
nand U28137 (N_28137,N_27239,N_27077);
nand U28138 (N_28138,N_27417,N_27460);
or U28139 (N_28139,N_27211,N_27587);
nand U28140 (N_28140,N_27559,N_27122);
or U28141 (N_28141,N_27342,N_27205);
and U28142 (N_28142,N_27285,N_27174);
and U28143 (N_28143,N_27094,N_27173);
xnor U28144 (N_28144,N_27191,N_27060);
xnor U28145 (N_28145,N_27587,N_27113);
nand U28146 (N_28146,N_27383,N_27168);
xor U28147 (N_28147,N_27067,N_27318);
nor U28148 (N_28148,N_27274,N_27374);
nand U28149 (N_28149,N_27517,N_27437);
xor U28150 (N_28150,N_27489,N_27265);
or U28151 (N_28151,N_27528,N_27570);
nor U28152 (N_28152,N_27232,N_27020);
nand U28153 (N_28153,N_27276,N_27058);
nand U28154 (N_28154,N_27469,N_27260);
or U28155 (N_28155,N_27303,N_27409);
xnor U28156 (N_28156,N_27086,N_27278);
or U28157 (N_28157,N_27490,N_27282);
nand U28158 (N_28158,N_27056,N_27458);
or U28159 (N_28159,N_27145,N_27391);
xnor U28160 (N_28160,N_27046,N_27014);
and U28161 (N_28161,N_27453,N_27573);
xor U28162 (N_28162,N_27426,N_27530);
nand U28163 (N_28163,N_27174,N_27224);
nand U28164 (N_28164,N_27049,N_27326);
nor U28165 (N_28165,N_27130,N_27546);
nor U28166 (N_28166,N_27449,N_27358);
and U28167 (N_28167,N_27298,N_27369);
and U28168 (N_28168,N_27190,N_27198);
xnor U28169 (N_28169,N_27379,N_27423);
or U28170 (N_28170,N_27015,N_27133);
or U28171 (N_28171,N_27168,N_27494);
or U28172 (N_28172,N_27290,N_27323);
nand U28173 (N_28173,N_27180,N_27176);
and U28174 (N_28174,N_27251,N_27393);
or U28175 (N_28175,N_27064,N_27531);
xor U28176 (N_28176,N_27540,N_27303);
nor U28177 (N_28177,N_27034,N_27585);
or U28178 (N_28178,N_27519,N_27542);
and U28179 (N_28179,N_27216,N_27048);
nor U28180 (N_28180,N_27318,N_27076);
xnor U28181 (N_28181,N_27071,N_27306);
xnor U28182 (N_28182,N_27018,N_27254);
nor U28183 (N_28183,N_27013,N_27394);
nor U28184 (N_28184,N_27566,N_27005);
and U28185 (N_28185,N_27426,N_27388);
nor U28186 (N_28186,N_27321,N_27357);
and U28187 (N_28187,N_27466,N_27229);
and U28188 (N_28188,N_27252,N_27223);
nor U28189 (N_28189,N_27415,N_27216);
nor U28190 (N_28190,N_27480,N_27580);
or U28191 (N_28191,N_27477,N_27188);
or U28192 (N_28192,N_27176,N_27080);
nand U28193 (N_28193,N_27239,N_27407);
and U28194 (N_28194,N_27528,N_27220);
xor U28195 (N_28195,N_27571,N_27324);
or U28196 (N_28196,N_27253,N_27114);
and U28197 (N_28197,N_27426,N_27126);
or U28198 (N_28198,N_27389,N_27233);
nand U28199 (N_28199,N_27139,N_27441);
or U28200 (N_28200,N_28096,N_28121);
xor U28201 (N_28201,N_27792,N_27918);
and U28202 (N_28202,N_28042,N_28095);
nand U28203 (N_28203,N_27606,N_27762);
nand U28204 (N_28204,N_27706,N_27707);
nand U28205 (N_28205,N_27842,N_27702);
or U28206 (N_28206,N_27978,N_28059);
nor U28207 (N_28207,N_28089,N_27872);
nand U28208 (N_28208,N_27867,N_27733);
nand U28209 (N_28209,N_27881,N_27808);
nor U28210 (N_28210,N_27697,N_28085);
nor U28211 (N_28211,N_28160,N_28175);
nand U28212 (N_28212,N_27664,N_27700);
or U28213 (N_28213,N_27941,N_27734);
nand U28214 (N_28214,N_27802,N_27995);
and U28215 (N_28215,N_28140,N_27758);
nor U28216 (N_28216,N_28035,N_27783);
and U28217 (N_28217,N_27648,N_27622);
nand U28218 (N_28218,N_28046,N_27753);
xor U28219 (N_28219,N_28161,N_27711);
nand U28220 (N_28220,N_27732,N_28019);
nand U28221 (N_28221,N_27938,N_28006);
xor U28222 (N_28222,N_27774,N_28052);
nand U28223 (N_28223,N_27832,N_28015);
xor U28224 (N_28224,N_27831,N_27666);
or U28225 (N_28225,N_27903,N_28166);
and U28226 (N_28226,N_28113,N_27725);
nand U28227 (N_28227,N_28021,N_27931);
xor U28228 (N_28228,N_27628,N_27954);
nor U28229 (N_28229,N_27912,N_27811);
xor U28230 (N_28230,N_27804,N_27916);
nand U28231 (N_28231,N_27806,N_28002);
nor U28232 (N_28232,N_28011,N_28056);
xor U28233 (N_28233,N_28040,N_27679);
nand U28234 (N_28234,N_27636,N_27671);
or U28235 (N_28235,N_27830,N_27997);
nor U28236 (N_28236,N_27647,N_28125);
xnor U28237 (N_28237,N_27866,N_27801);
and U28238 (N_28238,N_28107,N_27935);
or U28239 (N_28239,N_28139,N_28181);
xnor U28240 (N_28240,N_28116,N_27724);
or U28241 (N_28241,N_28092,N_27676);
and U28242 (N_28242,N_27678,N_27601);
and U28243 (N_28243,N_28047,N_27630);
xor U28244 (N_28244,N_28167,N_27996);
or U28245 (N_28245,N_27654,N_27943);
nand U28246 (N_28246,N_28106,N_27855);
nand U28247 (N_28247,N_28098,N_28124);
nor U28248 (N_28248,N_27876,N_27992);
and U28249 (N_28249,N_27719,N_27788);
or U28250 (N_28250,N_28178,N_28193);
or U28251 (N_28251,N_27930,N_28008);
and U28252 (N_28252,N_28126,N_27746);
and U28253 (N_28253,N_28182,N_28164);
nand U28254 (N_28254,N_27991,N_27735);
and U28255 (N_28255,N_27993,N_27875);
nor U28256 (N_28256,N_27626,N_27764);
nand U28257 (N_28257,N_28142,N_28173);
xnor U28258 (N_28258,N_27785,N_28060);
nor U28259 (N_28259,N_27977,N_27698);
nor U28260 (N_28260,N_28038,N_28159);
xnor U28261 (N_28261,N_28058,N_28109);
and U28262 (N_28262,N_27983,N_28063);
nand U28263 (N_28263,N_27965,N_27895);
or U28264 (N_28264,N_28103,N_27945);
nand U28265 (N_28265,N_27906,N_27981);
nand U28266 (N_28266,N_27794,N_28131);
or U28267 (N_28267,N_27932,N_27685);
or U28268 (N_28268,N_27959,N_28027);
nor U28269 (N_28269,N_27760,N_28065);
nand U28270 (N_28270,N_27948,N_27791);
nand U28271 (N_28271,N_27772,N_27882);
or U28272 (N_28272,N_28143,N_28184);
nor U28273 (N_28273,N_28022,N_27793);
and U28274 (N_28274,N_27990,N_28099);
nand U28275 (N_28275,N_27957,N_28194);
and U28276 (N_28276,N_28196,N_27950);
xnor U28277 (N_28277,N_28188,N_27694);
or U28278 (N_28278,N_27728,N_27869);
or U28279 (N_28279,N_27665,N_28189);
and U28280 (N_28280,N_27845,N_27909);
nor U28281 (N_28281,N_27956,N_27844);
and U28282 (N_28282,N_27754,N_27898);
or U28283 (N_28283,N_27780,N_27994);
or U28284 (N_28284,N_27973,N_27718);
nor U28285 (N_28285,N_28162,N_27674);
and U28286 (N_28286,N_27657,N_27638);
and U28287 (N_28287,N_28150,N_28153);
xnor U28288 (N_28288,N_28149,N_28134);
xnor U28289 (N_28289,N_27825,N_27737);
xor U28290 (N_28290,N_27656,N_27926);
nor U28291 (N_28291,N_27857,N_28148);
xnor U28292 (N_28292,N_27921,N_27602);
xnor U28293 (N_28293,N_28000,N_28062);
and U28294 (N_28294,N_28133,N_27815);
or U28295 (N_28295,N_27980,N_28064);
xnor U28296 (N_28296,N_27797,N_28014);
or U28297 (N_28297,N_27765,N_28190);
xnor U28298 (N_28298,N_28013,N_27796);
nand U28299 (N_28299,N_27879,N_27951);
xor U28300 (N_28300,N_27800,N_28079);
xor U28301 (N_28301,N_27984,N_27917);
xor U28302 (N_28302,N_28165,N_27803);
or U28303 (N_28303,N_28177,N_28078);
nand U28304 (N_28304,N_27610,N_27720);
and U28305 (N_28305,N_27805,N_27986);
nor U28306 (N_28306,N_28016,N_27982);
nand U28307 (N_28307,N_27861,N_27816);
and U28308 (N_28308,N_27618,N_27858);
and U28309 (N_28309,N_27692,N_27829);
nand U28310 (N_28310,N_27949,N_27639);
nand U28311 (N_28311,N_27778,N_27766);
nor U28312 (N_28312,N_27634,N_27669);
nand U28313 (N_28313,N_27809,N_27722);
nand U28314 (N_28314,N_28043,N_27874);
xnor U28315 (N_28315,N_28151,N_27848);
or U28316 (N_28316,N_28075,N_28132);
or U28317 (N_28317,N_28025,N_28071);
or U28318 (N_28318,N_27668,N_28045);
nand U28319 (N_28319,N_27911,N_27904);
nand U28320 (N_28320,N_27742,N_27641);
nand U28321 (N_28321,N_27854,N_27726);
xnor U28322 (N_28322,N_27976,N_27643);
nand U28323 (N_28323,N_28057,N_28101);
xnor U28324 (N_28324,N_27755,N_27924);
or U28325 (N_28325,N_28074,N_28127);
nor U28326 (N_28326,N_27709,N_27773);
nand U28327 (N_28327,N_27814,N_28195);
xnor U28328 (N_28328,N_28136,N_27684);
xor U28329 (N_28329,N_28135,N_28156);
nand U28330 (N_28330,N_27953,N_28172);
nand U28331 (N_28331,N_27786,N_27936);
nand U28332 (N_28332,N_28028,N_28141);
xnor U28333 (N_28333,N_27900,N_28197);
or U28334 (N_28334,N_28061,N_27836);
nand U28335 (N_28335,N_27812,N_27840);
xor U28336 (N_28336,N_27987,N_28048);
xor U28337 (N_28337,N_28128,N_28050);
nand U28338 (N_28338,N_27972,N_27969);
xor U28339 (N_28339,N_27907,N_27777);
nor U28340 (N_28340,N_27891,N_28171);
and U28341 (N_28341,N_27860,N_27738);
xor U28342 (N_28342,N_28137,N_27751);
nor U28343 (N_28343,N_27768,N_27999);
and U28344 (N_28344,N_28102,N_28155);
xor U28345 (N_28345,N_28012,N_27672);
nand U28346 (N_28346,N_27940,N_27998);
nor U28347 (N_28347,N_27871,N_27631);
or U28348 (N_28348,N_27819,N_27759);
nand U28349 (N_28349,N_27682,N_27644);
or U28350 (N_28350,N_27795,N_27856);
or U28351 (N_28351,N_28157,N_27810);
and U28352 (N_28352,N_27704,N_28199);
nor U28353 (N_28353,N_27888,N_27710);
xor U28354 (N_28354,N_27962,N_27868);
nand U28355 (N_28355,N_27649,N_28018);
nor U28356 (N_28356,N_27627,N_27988);
xnor U28357 (N_28357,N_27789,N_27933);
xnor U28358 (N_28358,N_27667,N_27713);
or U28359 (N_28359,N_28054,N_28147);
or U28360 (N_28360,N_27749,N_28007);
nand U28361 (N_28361,N_27885,N_27934);
nor U28362 (N_28362,N_27889,N_28146);
xor U28363 (N_28363,N_28129,N_28097);
nand U28364 (N_28364,N_27779,N_28034);
or U28365 (N_28365,N_27901,N_27970);
and U28366 (N_28366,N_27769,N_28031);
and U28367 (N_28367,N_28017,N_28003);
nor U28368 (N_28368,N_27745,N_27877);
and U28369 (N_28369,N_28083,N_27699);
or U28370 (N_28370,N_28029,N_28115);
nor U28371 (N_28371,N_27971,N_27818);
nor U28372 (N_28372,N_27723,N_27946);
nand U28373 (N_28373,N_27756,N_27646);
xor U28374 (N_28374,N_28049,N_27850);
nor U28375 (N_28375,N_27928,N_27937);
nor U28376 (N_28376,N_27712,N_28158);
xor U28377 (N_28377,N_27897,N_28069);
nor U28378 (N_28378,N_27989,N_28004);
nand U28379 (N_28379,N_27731,N_27975);
nand U28380 (N_28380,N_27873,N_27767);
nand U28381 (N_28381,N_27899,N_27862);
nand U28382 (N_28382,N_27663,N_27919);
xnor U28383 (N_28383,N_27955,N_28020);
nand U28384 (N_28384,N_28070,N_27683);
nand U28385 (N_28385,N_27750,N_27614);
and U28386 (N_28386,N_27880,N_27629);
xnor U28387 (N_28387,N_27859,N_28192);
or U28388 (N_28388,N_27616,N_27966);
nand U28389 (N_28389,N_27799,N_28010);
nand U28390 (N_28390,N_27890,N_27691);
nand U28391 (N_28391,N_27823,N_27822);
or U28392 (N_28392,N_27675,N_27905);
xnor U28393 (N_28393,N_28093,N_27673);
and U28394 (N_28394,N_27696,N_27894);
nor U28395 (N_28395,N_27979,N_27782);
xor U28396 (N_28396,N_28105,N_28174);
xor U28397 (N_28397,N_27608,N_27775);
nor U28398 (N_28398,N_27841,N_27770);
and U28399 (N_28399,N_27621,N_27607);
and U28400 (N_28400,N_27910,N_27705);
xor U28401 (N_28401,N_27961,N_27717);
and U28402 (N_28402,N_28039,N_28067);
nand U28403 (N_28403,N_27680,N_27662);
nand U28404 (N_28404,N_27923,N_27837);
and U28405 (N_28405,N_28198,N_27915);
and U28406 (N_28406,N_27776,N_27687);
or U28407 (N_28407,N_27701,N_28044);
nor U28408 (N_28408,N_27703,N_27820);
xnor U28409 (N_28409,N_27693,N_27849);
or U28410 (N_28410,N_27615,N_27736);
nand U28411 (N_28411,N_27964,N_27851);
or U28412 (N_28412,N_27893,N_28082);
and U28413 (N_28413,N_28053,N_27878);
nor U28414 (N_28414,N_27958,N_27833);
nand U28415 (N_28415,N_27744,N_28001);
and U28416 (N_28416,N_27920,N_27613);
nand U28417 (N_28417,N_28114,N_27828);
nor U28418 (N_28418,N_28111,N_27847);
nor U28419 (N_28419,N_27985,N_27838);
xor U28420 (N_28420,N_27908,N_27690);
xnor U28421 (N_28421,N_28051,N_27681);
and U28422 (N_28422,N_27743,N_27807);
xnor U28423 (N_28423,N_27974,N_27784);
or U28424 (N_28424,N_28138,N_27887);
nand U28425 (N_28425,N_28072,N_28120);
or U28426 (N_28426,N_27952,N_27863);
and U28427 (N_28427,N_27865,N_27927);
xor U28428 (N_28428,N_28119,N_27939);
or U28429 (N_28429,N_27813,N_27624);
and U28430 (N_28430,N_27650,N_27611);
xnor U28431 (N_28431,N_27896,N_27914);
xnor U28432 (N_28432,N_28076,N_28055);
nor U28433 (N_28433,N_28100,N_27884);
nand U28434 (N_28434,N_28168,N_27716);
nand U28435 (N_28435,N_27947,N_28169);
or U28436 (N_28436,N_27642,N_28077);
or U28437 (N_28437,N_28084,N_27612);
nor U28438 (N_28438,N_27821,N_27660);
xnor U28439 (N_28439,N_28112,N_27967);
xnor U28440 (N_28440,N_28026,N_27913);
xnor U28441 (N_28441,N_27963,N_27827);
or U28442 (N_28442,N_28036,N_27787);
xor U28443 (N_28443,N_27730,N_27883);
or U28444 (N_28444,N_27790,N_27925);
nor U28445 (N_28445,N_27886,N_27741);
xor U28446 (N_28446,N_27619,N_27620);
nand U28447 (N_28447,N_28037,N_28066);
or U28448 (N_28448,N_27968,N_28191);
xnor U28449 (N_28449,N_27686,N_27670);
or U28450 (N_28450,N_27853,N_28086);
nor U28451 (N_28451,N_27689,N_27623);
nand U28452 (N_28452,N_27846,N_28123);
xor U28453 (N_28453,N_28110,N_28180);
and U28454 (N_28454,N_28183,N_27651);
or U28455 (N_28455,N_27729,N_27870);
nor U28456 (N_28456,N_27695,N_27739);
or U28457 (N_28457,N_28041,N_27824);
and U28458 (N_28458,N_27817,N_28144);
nand U28459 (N_28459,N_27645,N_28090);
and U28460 (N_28460,N_27834,N_28033);
and U28461 (N_28461,N_27892,N_27747);
and U28462 (N_28462,N_28009,N_27798);
or U28463 (N_28463,N_28024,N_27632);
and U28464 (N_28464,N_27839,N_27600);
xor U28465 (N_28465,N_28081,N_28068);
xnor U28466 (N_28466,N_28154,N_27625);
nor U28467 (N_28467,N_28186,N_27761);
or U28468 (N_28468,N_27721,N_28179);
and U28469 (N_28469,N_27752,N_27944);
and U28470 (N_28470,N_27640,N_27843);
or U28471 (N_28471,N_28145,N_28170);
xor U28472 (N_28472,N_27864,N_28104);
nand U28473 (N_28473,N_27835,N_28030);
nand U28474 (N_28474,N_27633,N_27655);
nor U28475 (N_28475,N_28080,N_28163);
and U28476 (N_28476,N_27637,N_28152);
and U28477 (N_28477,N_27661,N_27715);
or U28478 (N_28478,N_27603,N_27771);
xnor U28479 (N_28479,N_27727,N_27652);
and U28480 (N_28480,N_27781,N_28073);
xor U28481 (N_28481,N_28094,N_27677);
and U28482 (N_28482,N_27658,N_27617);
xor U28483 (N_28483,N_28005,N_27929);
xor U28484 (N_28484,N_27763,N_28130);
xnor U28485 (N_28485,N_27635,N_27653);
nand U28486 (N_28486,N_28108,N_27902);
and U28487 (N_28487,N_28032,N_27942);
xor U28488 (N_28488,N_27708,N_27688);
xor U28489 (N_28489,N_27922,N_28087);
nand U28490 (N_28490,N_27748,N_28117);
and U28491 (N_28491,N_28118,N_28122);
or U28492 (N_28492,N_28176,N_28185);
nor U28493 (N_28493,N_27852,N_27960);
xnor U28494 (N_28494,N_27714,N_28023);
or U28495 (N_28495,N_27740,N_27659);
or U28496 (N_28496,N_27604,N_28088);
or U28497 (N_28497,N_28091,N_28187);
nor U28498 (N_28498,N_27609,N_27757);
and U28499 (N_28499,N_27605,N_27826);
xnor U28500 (N_28500,N_27769,N_27918);
xnor U28501 (N_28501,N_27715,N_27722);
nor U28502 (N_28502,N_28145,N_27741);
nand U28503 (N_28503,N_28095,N_27902);
nor U28504 (N_28504,N_27862,N_28033);
nor U28505 (N_28505,N_27740,N_28043);
nor U28506 (N_28506,N_27805,N_27771);
nor U28507 (N_28507,N_27618,N_27658);
and U28508 (N_28508,N_27688,N_27669);
xor U28509 (N_28509,N_27949,N_27842);
nand U28510 (N_28510,N_28148,N_28041);
and U28511 (N_28511,N_27897,N_27784);
or U28512 (N_28512,N_27992,N_27784);
nor U28513 (N_28513,N_27775,N_27613);
nor U28514 (N_28514,N_27817,N_27916);
or U28515 (N_28515,N_27748,N_28169);
or U28516 (N_28516,N_27699,N_27842);
or U28517 (N_28517,N_27678,N_28125);
and U28518 (N_28518,N_28190,N_28186);
and U28519 (N_28519,N_27769,N_27896);
or U28520 (N_28520,N_27916,N_27936);
nor U28521 (N_28521,N_27722,N_28007);
and U28522 (N_28522,N_28109,N_28099);
nand U28523 (N_28523,N_27646,N_28163);
nand U28524 (N_28524,N_27966,N_28017);
and U28525 (N_28525,N_27957,N_27695);
nor U28526 (N_28526,N_27666,N_28085);
or U28527 (N_28527,N_27688,N_27888);
nor U28528 (N_28528,N_27750,N_27755);
or U28529 (N_28529,N_28096,N_27694);
and U28530 (N_28530,N_27995,N_27840);
nor U28531 (N_28531,N_27850,N_27805);
and U28532 (N_28532,N_28103,N_27636);
xor U28533 (N_28533,N_28034,N_27661);
xnor U28534 (N_28534,N_27915,N_27634);
or U28535 (N_28535,N_27832,N_28162);
or U28536 (N_28536,N_28171,N_27825);
nand U28537 (N_28537,N_27857,N_27868);
or U28538 (N_28538,N_27737,N_27788);
or U28539 (N_28539,N_27982,N_28182);
xnor U28540 (N_28540,N_27669,N_28180);
and U28541 (N_28541,N_27798,N_27662);
and U28542 (N_28542,N_27676,N_27808);
xor U28543 (N_28543,N_27666,N_27856);
nor U28544 (N_28544,N_27712,N_27867);
nand U28545 (N_28545,N_27722,N_27967);
and U28546 (N_28546,N_27760,N_28024);
nand U28547 (N_28547,N_27838,N_27763);
nor U28548 (N_28548,N_27995,N_27633);
xnor U28549 (N_28549,N_27721,N_27712);
and U28550 (N_28550,N_27909,N_27943);
xnor U28551 (N_28551,N_28199,N_28051);
or U28552 (N_28552,N_28177,N_27616);
nor U28553 (N_28553,N_27758,N_28132);
nor U28554 (N_28554,N_27920,N_27642);
and U28555 (N_28555,N_27640,N_27929);
and U28556 (N_28556,N_27827,N_28031);
nand U28557 (N_28557,N_28133,N_28149);
nand U28558 (N_28558,N_27816,N_28089);
xnor U28559 (N_28559,N_28197,N_27919);
nand U28560 (N_28560,N_27949,N_27655);
nand U28561 (N_28561,N_27969,N_27743);
nand U28562 (N_28562,N_28036,N_28002);
or U28563 (N_28563,N_27980,N_27604);
nand U28564 (N_28564,N_27606,N_27693);
or U28565 (N_28565,N_28132,N_27679);
or U28566 (N_28566,N_28147,N_27681);
xor U28567 (N_28567,N_28129,N_27660);
nor U28568 (N_28568,N_27733,N_27782);
nor U28569 (N_28569,N_27658,N_28183);
or U28570 (N_28570,N_27972,N_28098);
xor U28571 (N_28571,N_28075,N_27936);
nor U28572 (N_28572,N_27888,N_28007);
nor U28573 (N_28573,N_27714,N_28167);
nand U28574 (N_28574,N_27926,N_27814);
nor U28575 (N_28575,N_27781,N_28028);
nand U28576 (N_28576,N_27830,N_28004);
nand U28577 (N_28577,N_27949,N_27829);
nand U28578 (N_28578,N_28135,N_28113);
nand U28579 (N_28579,N_27682,N_27734);
xnor U28580 (N_28580,N_27846,N_27627);
and U28581 (N_28581,N_28184,N_27691);
nor U28582 (N_28582,N_28082,N_27917);
or U28583 (N_28583,N_27853,N_28003);
and U28584 (N_28584,N_27775,N_28020);
nor U28585 (N_28585,N_27810,N_27819);
nand U28586 (N_28586,N_27773,N_27870);
xor U28587 (N_28587,N_27868,N_27678);
and U28588 (N_28588,N_28056,N_28098);
xnor U28589 (N_28589,N_27661,N_27666);
nand U28590 (N_28590,N_27875,N_27710);
and U28591 (N_28591,N_27635,N_28189);
or U28592 (N_28592,N_27693,N_27702);
nand U28593 (N_28593,N_27942,N_28125);
xnor U28594 (N_28594,N_28176,N_28065);
nand U28595 (N_28595,N_28145,N_27978);
and U28596 (N_28596,N_27975,N_27944);
xnor U28597 (N_28597,N_28172,N_27867);
nor U28598 (N_28598,N_28008,N_28147);
and U28599 (N_28599,N_28116,N_27827);
and U28600 (N_28600,N_28132,N_27728);
and U28601 (N_28601,N_28137,N_28133);
or U28602 (N_28602,N_27657,N_27624);
nand U28603 (N_28603,N_28197,N_28071);
xnor U28604 (N_28604,N_27969,N_27725);
nand U28605 (N_28605,N_27734,N_27875);
and U28606 (N_28606,N_28028,N_27891);
or U28607 (N_28607,N_28087,N_27998);
nand U28608 (N_28608,N_28113,N_28040);
nand U28609 (N_28609,N_27699,N_27866);
or U28610 (N_28610,N_27871,N_28085);
and U28611 (N_28611,N_27601,N_28086);
and U28612 (N_28612,N_27750,N_27851);
xnor U28613 (N_28613,N_27679,N_27699);
or U28614 (N_28614,N_27670,N_27832);
and U28615 (N_28615,N_27617,N_27744);
or U28616 (N_28616,N_27643,N_27677);
nor U28617 (N_28617,N_28184,N_27783);
or U28618 (N_28618,N_27696,N_27998);
and U28619 (N_28619,N_28101,N_28097);
nor U28620 (N_28620,N_27615,N_27756);
nor U28621 (N_28621,N_27716,N_27739);
or U28622 (N_28622,N_28081,N_28015);
nand U28623 (N_28623,N_28117,N_27927);
xor U28624 (N_28624,N_28131,N_27838);
and U28625 (N_28625,N_27953,N_27629);
or U28626 (N_28626,N_27903,N_28018);
nor U28627 (N_28627,N_28072,N_28141);
xnor U28628 (N_28628,N_27733,N_27897);
nor U28629 (N_28629,N_27753,N_27848);
or U28630 (N_28630,N_27756,N_27723);
and U28631 (N_28631,N_28023,N_27939);
nand U28632 (N_28632,N_28018,N_27652);
and U28633 (N_28633,N_27971,N_28196);
or U28634 (N_28634,N_27862,N_27996);
xor U28635 (N_28635,N_27966,N_27768);
xor U28636 (N_28636,N_28172,N_27648);
or U28637 (N_28637,N_27864,N_27782);
nand U28638 (N_28638,N_28170,N_27952);
or U28639 (N_28639,N_27916,N_27843);
or U28640 (N_28640,N_27682,N_28187);
and U28641 (N_28641,N_27951,N_27991);
nand U28642 (N_28642,N_28188,N_27668);
nor U28643 (N_28643,N_28063,N_27889);
nand U28644 (N_28644,N_27759,N_28133);
and U28645 (N_28645,N_27657,N_27755);
and U28646 (N_28646,N_27904,N_27616);
or U28647 (N_28647,N_28012,N_28001);
or U28648 (N_28648,N_27962,N_27796);
and U28649 (N_28649,N_27989,N_27689);
or U28650 (N_28650,N_27994,N_28144);
xor U28651 (N_28651,N_28078,N_28136);
or U28652 (N_28652,N_28017,N_28043);
nand U28653 (N_28653,N_27929,N_27723);
nor U28654 (N_28654,N_27908,N_27724);
or U28655 (N_28655,N_27631,N_27705);
nand U28656 (N_28656,N_28046,N_27832);
nor U28657 (N_28657,N_27897,N_27861);
nand U28658 (N_28658,N_27694,N_28064);
and U28659 (N_28659,N_28024,N_27863);
nor U28660 (N_28660,N_27692,N_28176);
xor U28661 (N_28661,N_27998,N_28009);
nor U28662 (N_28662,N_28179,N_27969);
nor U28663 (N_28663,N_27902,N_27607);
nand U28664 (N_28664,N_28094,N_27844);
xnor U28665 (N_28665,N_27981,N_28077);
xnor U28666 (N_28666,N_28173,N_27976);
nand U28667 (N_28667,N_27821,N_27781);
nand U28668 (N_28668,N_27910,N_27904);
xor U28669 (N_28669,N_28049,N_28103);
nor U28670 (N_28670,N_28195,N_27704);
xor U28671 (N_28671,N_27858,N_27884);
xnor U28672 (N_28672,N_28024,N_27995);
nor U28673 (N_28673,N_28100,N_28066);
nand U28674 (N_28674,N_27960,N_27928);
nor U28675 (N_28675,N_28012,N_27608);
xor U28676 (N_28676,N_27705,N_27785);
xnor U28677 (N_28677,N_27933,N_27831);
xor U28678 (N_28678,N_27780,N_27658);
nand U28679 (N_28679,N_27919,N_27720);
nor U28680 (N_28680,N_28048,N_28120);
or U28681 (N_28681,N_27772,N_27971);
or U28682 (N_28682,N_27608,N_27904);
nand U28683 (N_28683,N_28137,N_27645);
or U28684 (N_28684,N_28004,N_27785);
and U28685 (N_28685,N_27969,N_27791);
nor U28686 (N_28686,N_27941,N_27645);
nor U28687 (N_28687,N_27794,N_28134);
nand U28688 (N_28688,N_27833,N_27689);
nand U28689 (N_28689,N_27875,N_27947);
or U28690 (N_28690,N_28090,N_27756);
or U28691 (N_28691,N_27870,N_28197);
nor U28692 (N_28692,N_28101,N_27766);
or U28693 (N_28693,N_27680,N_27641);
nand U28694 (N_28694,N_27965,N_27876);
xnor U28695 (N_28695,N_27627,N_27628);
xor U28696 (N_28696,N_27970,N_27986);
nand U28697 (N_28697,N_27976,N_28127);
nor U28698 (N_28698,N_27949,N_27613);
or U28699 (N_28699,N_28095,N_27960);
nor U28700 (N_28700,N_28051,N_28151);
xor U28701 (N_28701,N_27843,N_27697);
and U28702 (N_28702,N_28003,N_27774);
and U28703 (N_28703,N_27992,N_27601);
or U28704 (N_28704,N_27773,N_28030);
and U28705 (N_28705,N_28126,N_27955);
or U28706 (N_28706,N_27827,N_27623);
nor U28707 (N_28707,N_28151,N_27650);
xnor U28708 (N_28708,N_27803,N_28064);
nand U28709 (N_28709,N_27861,N_27981);
nand U28710 (N_28710,N_27773,N_27913);
xnor U28711 (N_28711,N_28039,N_27939);
nor U28712 (N_28712,N_27776,N_27608);
or U28713 (N_28713,N_27629,N_28162);
nor U28714 (N_28714,N_28053,N_27826);
nor U28715 (N_28715,N_27787,N_27886);
xor U28716 (N_28716,N_28097,N_27722);
and U28717 (N_28717,N_27996,N_27816);
nor U28718 (N_28718,N_27779,N_27630);
or U28719 (N_28719,N_27951,N_27625);
xnor U28720 (N_28720,N_27765,N_27945);
or U28721 (N_28721,N_27729,N_28121);
and U28722 (N_28722,N_27809,N_28169);
xor U28723 (N_28723,N_27966,N_28032);
xor U28724 (N_28724,N_27882,N_28016);
and U28725 (N_28725,N_27762,N_27702);
nor U28726 (N_28726,N_27608,N_27761);
nor U28727 (N_28727,N_28134,N_27649);
and U28728 (N_28728,N_27794,N_27699);
nor U28729 (N_28729,N_27712,N_28011);
nor U28730 (N_28730,N_27934,N_27891);
nand U28731 (N_28731,N_27866,N_28125);
or U28732 (N_28732,N_28111,N_27920);
nor U28733 (N_28733,N_28188,N_28046);
or U28734 (N_28734,N_27868,N_28102);
xor U28735 (N_28735,N_28184,N_27927);
nand U28736 (N_28736,N_28161,N_28101);
or U28737 (N_28737,N_27879,N_27976);
nor U28738 (N_28738,N_27845,N_27856);
and U28739 (N_28739,N_27685,N_27933);
xnor U28740 (N_28740,N_27882,N_27913);
nand U28741 (N_28741,N_28157,N_27988);
nor U28742 (N_28742,N_28069,N_27630);
or U28743 (N_28743,N_28097,N_27655);
and U28744 (N_28744,N_27761,N_27687);
nand U28745 (N_28745,N_28108,N_27806);
xor U28746 (N_28746,N_28173,N_27947);
or U28747 (N_28747,N_28128,N_27939);
nand U28748 (N_28748,N_27789,N_28081);
nor U28749 (N_28749,N_27906,N_28176);
xnor U28750 (N_28750,N_27999,N_28163);
and U28751 (N_28751,N_27782,N_27982);
and U28752 (N_28752,N_28196,N_27856);
or U28753 (N_28753,N_27625,N_27822);
or U28754 (N_28754,N_27922,N_28034);
xor U28755 (N_28755,N_27692,N_28146);
nor U28756 (N_28756,N_28114,N_27971);
nor U28757 (N_28757,N_28189,N_28120);
and U28758 (N_28758,N_27737,N_27689);
nand U28759 (N_28759,N_28021,N_27677);
nand U28760 (N_28760,N_27961,N_28130);
or U28761 (N_28761,N_27685,N_27775);
or U28762 (N_28762,N_27683,N_27879);
xor U28763 (N_28763,N_28077,N_28187);
nor U28764 (N_28764,N_27859,N_27850);
xor U28765 (N_28765,N_28085,N_28133);
nand U28766 (N_28766,N_28129,N_28173);
and U28767 (N_28767,N_28184,N_27640);
nor U28768 (N_28768,N_27985,N_27703);
nor U28769 (N_28769,N_28106,N_27782);
and U28770 (N_28770,N_27798,N_27850);
nor U28771 (N_28771,N_28177,N_27823);
nand U28772 (N_28772,N_27794,N_27760);
or U28773 (N_28773,N_27836,N_27621);
nand U28774 (N_28774,N_27930,N_28102);
nand U28775 (N_28775,N_27778,N_28128);
nor U28776 (N_28776,N_28108,N_27949);
xor U28777 (N_28777,N_27869,N_27836);
or U28778 (N_28778,N_28184,N_28016);
and U28779 (N_28779,N_27788,N_27840);
nor U28780 (N_28780,N_28196,N_27682);
and U28781 (N_28781,N_27946,N_28124);
and U28782 (N_28782,N_28087,N_27962);
xnor U28783 (N_28783,N_27920,N_28188);
or U28784 (N_28784,N_27631,N_28008);
nand U28785 (N_28785,N_27967,N_28126);
or U28786 (N_28786,N_27965,N_28085);
nand U28787 (N_28787,N_27724,N_28103);
nor U28788 (N_28788,N_27659,N_27640);
nand U28789 (N_28789,N_27908,N_28098);
nor U28790 (N_28790,N_27714,N_27759);
xor U28791 (N_28791,N_27916,N_28174);
nand U28792 (N_28792,N_28183,N_28015);
or U28793 (N_28793,N_28016,N_27645);
and U28794 (N_28794,N_28038,N_27661);
nor U28795 (N_28795,N_27897,N_28076);
xor U28796 (N_28796,N_27620,N_28153);
nor U28797 (N_28797,N_27729,N_27689);
nor U28798 (N_28798,N_27734,N_28075);
nand U28799 (N_28799,N_27719,N_27681);
xnor U28800 (N_28800,N_28733,N_28620);
and U28801 (N_28801,N_28637,N_28482);
xnor U28802 (N_28802,N_28508,N_28486);
or U28803 (N_28803,N_28567,N_28248);
xnor U28804 (N_28804,N_28371,N_28354);
xnor U28805 (N_28805,N_28468,N_28747);
nand U28806 (N_28806,N_28613,N_28296);
nand U28807 (N_28807,N_28343,N_28385);
xnor U28808 (N_28808,N_28284,N_28741);
nand U28809 (N_28809,N_28616,N_28539);
or U28810 (N_28810,N_28570,N_28303);
xnor U28811 (N_28811,N_28345,N_28222);
nand U28812 (N_28812,N_28648,N_28207);
nand U28813 (N_28813,N_28753,N_28210);
and U28814 (N_28814,N_28458,N_28464);
xnor U28815 (N_28815,N_28367,N_28203);
or U28816 (N_28816,N_28557,N_28555);
and U28817 (N_28817,N_28756,N_28399);
nand U28818 (N_28818,N_28790,N_28693);
and U28819 (N_28819,N_28642,N_28766);
or U28820 (N_28820,N_28260,N_28734);
or U28821 (N_28821,N_28626,N_28772);
nand U28822 (N_28822,N_28730,N_28579);
or U28823 (N_28823,N_28434,N_28307);
nor U28824 (N_28824,N_28699,N_28256);
nand U28825 (N_28825,N_28624,N_28668);
nor U28826 (N_28826,N_28749,N_28584);
nor U28827 (N_28827,N_28606,N_28475);
xnor U28828 (N_28828,N_28576,N_28587);
xnor U28829 (N_28829,N_28568,N_28241);
and U28830 (N_28830,N_28578,N_28332);
xnor U28831 (N_28831,N_28411,N_28706);
nor U28832 (N_28832,N_28751,N_28655);
or U28833 (N_28833,N_28436,N_28299);
nand U28834 (N_28834,N_28205,N_28270);
and U28835 (N_28835,N_28533,N_28612);
or U28836 (N_28836,N_28268,N_28489);
or U28837 (N_28837,N_28378,N_28546);
nor U28838 (N_28838,N_28431,N_28283);
and U28839 (N_28839,N_28532,N_28602);
or U28840 (N_28840,N_28603,N_28477);
xnor U28841 (N_28841,N_28252,N_28690);
nor U28842 (N_28842,N_28561,N_28691);
or U28843 (N_28843,N_28535,N_28405);
xnor U28844 (N_28844,N_28279,N_28287);
nor U28845 (N_28845,N_28365,N_28630);
nand U28846 (N_28846,N_28590,N_28660);
or U28847 (N_28847,N_28285,N_28649);
and U28848 (N_28848,N_28764,N_28597);
and U28849 (N_28849,N_28615,N_28676);
xnor U28850 (N_28850,N_28293,N_28582);
and U28851 (N_28851,N_28692,N_28379);
and U28852 (N_28852,N_28485,N_28502);
xor U28853 (N_28853,N_28202,N_28524);
nand U28854 (N_28854,N_28674,N_28384);
nand U28855 (N_28855,N_28495,N_28233);
nor U28856 (N_28856,N_28552,N_28726);
xor U28857 (N_28857,N_28718,N_28407);
nor U28858 (N_28858,N_28586,N_28314);
or U28859 (N_28859,N_28439,N_28460);
nor U28860 (N_28860,N_28374,N_28491);
xnor U28861 (N_28861,N_28481,N_28452);
nor U28862 (N_28862,N_28498,N_28294);
nand U28863 (N_28863,N_28330,N_28640);
nand U28864 (N_28864,N_28271,N_28373);
or U28865 (N_28865,N_28480,N_28647);
nand U28866 (N_28866,N_28440,N_28797);
xnor U28867 (N_28867,N_28522,N_28664);
nor U28868 (N_28868,N_28243,N_28743);
xnor U28869 (N_28869,N_28698,N_28438);
and U28870 (N_28870,N_28705,N_28636);
nor U28871 (N_28871,N_28351,N_28449);
or U28872 (N_28872,N_28686,N_28467);
and U28873 (N_28873,N_28781,N_28657);
nor U28874 (N_28874,N_28462,N_28617);
or U28875 (N_28875,N_28221,N_28350);
and U28876 (N_28876,N_28391,N_28762);
xor U28877 (N_28877,N_28583,N_28518);
or U28878 (N_28878,N_28277,N_28656);
xnor U28879 (N_28879,N_28380,N_28638);
or U28880 (N_28880,N_28473,N_28707);
or U28881 (N_28881,N_28218,N_28445);
nand U28882 (N_28882,N_28635,N_28739);
and U28883 (N_28883,N_28750,N_28731);
or U28884 (N_28884,N_28684,N_28711);
nand U28885 (N_28885,N_28398,N_28775);
or U28886 (N_28886,N_28700,N_28703);
xnor U28887 (N_28887,N_28608,N_28776);
nand U28888 (N_28888,N_28499,N_28618);
nand U28889 (N_28889,N_28421,N_28665);
or U28890 (N_28890,N_28738,N_28249);
or U28891 (N_28891,N_28712,N_28235);
xnor U28892 (N_28892,N_28784,N_28304);
or U28893 (N_28893,N_28538,N_28329);
xor U28894 (N_28894,N_28396,N_28672);
and U28895 (N_28895,N_28461,N_28729);
nor U28896 (N_28896,N_28589,N_28250);
nand U28897 (N_28897,N_28497,N_28782);
or U28898 (N_28898,N_28791,N_28503);
nor U28899 (N_28899,N_28265,N_28798);
nor U28900 (N_28900,N_28383,N_28397);
nand U28901 (N_28901,N_28417,N_28326);
and U28902 (N_28902,N_28695,N_28621);
nor U28903 (N_28903,N_28785,N_28269);
nand U28904 (N_28904,N_28275,N_28607);
nand U28905 (N_28905,N_28795,N_28220);
or U28906 (N_28906,N_28216,N_28722);
nor U28907 (N_28907,N_28257,N_28771);
xnor U28908 (N_28908,N_28504,N_28321);
nor U28909 (N_28909,N_28496,N_28591);
and U28910 (N_28910,N_28356,N_28404);
nand U28911 (N_28911,N_28346,N_28459);
and U28912 (N_28912,N_28448,N_28789);
or U28913 (N_28913,N_28540,N_28702);
xnor U28914 (N_28914,N_28236,N_28646);
nor U28915 (N_28915,N_28315,N_28742);
and U28916 (N_28916,N_28454,N_28574);
xor U28917 (N_28917,N_28773,N_28752);
and U28918 (N_28918,N_28788,N_28357);
xor U28919 (N_28919,N_28687,N_28286);
or U28920 (N_28920,N_28768,N_28573);
xnor U28921 (N_28921,N_28488,N_28760);
nor U28922 (N_28922,N_28312,N_28728);
and U28923 (N_28923,N_28395,N_28639);
and U28924 (N_28924,N_28588,N_28231);
nor U28925 (N_28925,N_28331,N_28359);
or U28926 (N_28926,N_28644,N_28320);
and U28927 (N_28927,N_28564,N_28451);
nor U28928 (N_28928,N_28759,N_28337);
nand U28929 (N_28929,N_28453,N_28667);
nor U28930 (N_28930,N_28215,N_28387);
nand U28931 (N_28931,N_28364,N_28765);
xnor U28932 (N_28932,N_28470,N_28289);
nor U28933 (N_28933,N_28554,N_28677);
nor U28934 (N_28934,N_28758,N_28678);
nor U28935 (N_28935,N_28562,N_28406);
nand U28936 (N_28936,N_28336,N_28510);
and U28937 (N_28937,N_28605,N_28600);
nand U28938 (N_28938,N_28372,N_28507);
and U28939 (N_28939,N_28599,N_28575);
nand U28940 (N_28940,N_28394,N_28509);
or U28941 (N_28941,N_28292,N_28368);
nor U28942 (N_28942,N_28778,N_28519);
or U28943 (N_28943,N_28469,N_28247);
nor U28944 (N_28944,N_28536,N_28670);
nand U28945 (N_28945,N_28401,N_28541);
nand U28946 (N_28946,N_28594,N_28349);
nand U28947 (N_28947,N_28754,N_28446);
and U28948 (N_28948,N_28344,N_28457);
nor U28949 (N_28949,N_28263,N_28709);
and U28950 (N_28950,N_28413,N_28466);
xnor U28951 (N_28951,N_28681,N_28422);
nand U28952 (N_28952,N_28770,N_28757);
or U28953 (N_28953,N_28455,N_28200);
xor U28954 (N_28954,N_28529,N_28386);
or U28955 (N_28955,N_28290,N_28416);
or U28956 (N_28956,N_28226,N_28340);
nor U28957 (N_28957,N_28366,N_28558);
or U28958 (N_28958,N_28737,N_28382);
and U28959 (N_28959,N_28242,N_28774);
nor U28960 (N_28960,N_28763,N_28680);
or U28961 (N_28961,N_28651,N_28361);
nor U28962 (N_28962,N_28724,N_28305);
xnor U28963 (N_28963,N_28537,N_28297);
nor U28964 (N_28964,N_28259,N_28325);
and U28965 (N_28965,N_28273,N_28426);
xor U28966 (N_28966,N_28338,N_28542);
or U28967 (N_28967,N_28643,N_28238);
and U28968 (N_28968,N_28484,N_28794);
nand U28969 (N_28969,N_28355,N_28360);
or U28970 (N_28970,N_28623,N_28441);
and U28971 (N_28971,N_28217,N_28736);
and U28972 (N_28972,N_28531,N_28585);
nand U28973 (N_28973,N_28258,N_28209);
xor U28974 (N_28974,N_28412,N_28375);
nor U28975 (N_28975,N_28609,N_28362);
and U28976 (N_28976,N_28553,N_28409);
or U28977 (N_28977,N_28725,N_28628);
xnor U28978 (N_28978,N_28232,N_28427);
xor U28979 (N_28979,N_28746,N_28339);
or U28980 (N_28980,N_28548,N_28596);
nor U28981 (N_28981,N_28633,N_28214);
nand U28982 (N_28982,N_28632,N_28272);
or U28983 (N_28983,N_28428,N_28240);
xor U28984 (N_28984,N_28424,N_28223);
and U28985 (N_28985,N_28526,N_28423);
xnor U28986 (N_28986,N_28713,N_28653);
xnor U28987 (N_28987,N_28525,N_28493);
nand U28988 (N_28988,N_28652,N_28201);
nor U28989 (N_28989,N_28245,N_28334);
or U28990 (N_28990,N_28517,N_28661);
xor U28991 (N_28991,N_28761,N_28310);
nor U28992 (N_28992,N_28219,N_28571);
nor U28993 (N_28993,N_28363,N_28474);
nor U28994 (N_28994,N_28534,N_28316);
xor U28995 (N_28995,N_28313,N_28261);
or U28996 (N_28996,N_28550,N_28402);
and U28997 (N_28997,N_28543,N_28559);
nand U28998 (N_28998,N_28521,N_28476);
nor U28999 (N_28999,N_28530,N_28370);
nor U29000 (N_29000,N_28601,N_28282);
xnor U29001 (N_29001,N_28487,N_28388);
and U29002 (N_29002,N_28246,N_28450);
xor U29003 (N_29003,N_28704,N_28429);
or U29004 (N_29004,N_28443,N_28228);
nand U29005 (N_29005,N_28719,N_28442);
xor U29006 (N_29006,N_28377,N_28244);
and U29007 (N_29007,N_28627,N_28437);
nand U29008 (N_29008,N_28547,N_28463);
xnor U29009 (N_29009,N_28572,N_28727);
xnor U29010 (N_29010,N_28280,N_28319);
nor U29011 (N_29011,N_28237,N_28211);
xnor U29012 (N_29012,N_28322,N_28318);
or U29013 (N_29013,N_28456,N_28779);
and U29014 (N_29014,N_28565,N_28631);
and U29015 (N_29015,N_28777,N_28212);
xnor U29016 (N_29016,N_28716,N_28513);
nor U29017 (N_29017,N_28328,N_28381);
and U29018 (N_29018,N_28471,N_28604);
or U29019 (N_29019,N_28444,N_28786);
and U29020 (N_29020,N_28295,N_28641);
nand U29021 (N_29021,N_28433,N_28291);
nand U29022 (N_29022,N_28714,N_28253);
xor U29023 (N_29023,N_28796,N_28683);
or U29024 (N_29024,N_28347,N_28494);
xor U29025 (N_29025,N_28267,N_28302);
and U29026 (N_29026,N_28682,N_28420);
nor U29027 (N_29027,N_28717,N_28430);
xor U29028 (N_29028,N_28685,N_28419);
nor U29029 (N_29029,N_28662,N_28309);
nor U29030 (N_29030,N_28593,N_28392);
and U29031 (N_29031,N_28204,N_28629);
xor U29032 (N_29032,N_28276,N_28697);
nor U29033 (N_29033,N_28274,N_28769);
and U29034 (N_29034,N_28720,N_28208);
nor U29035 (N_29035,N_28516,N_28645);
nor U29036 (N_29036,N_28675,N_28306);
nor U29037 (N_29037,N_28688,N_28352);
nand U29038 (N_29038,N_28254,N_28580);
nand U29039 (N_29039,N_28732,N_28425);
and U29040 (N_29040,N_28472,N_28255);
nor U29041 (N_29041,N_28663,N_28595);
nor U29042 (N_29042,N_28658,N_28740);
nor U29043 (N_29043,N_28671,N_28654);
xnor U29044 (N_29044,N_28432,N_28225);
and U29045 (N_29045,N_28610,N_28483);
or U29046 (N_29046,N_28342,N_28435);
xor U29047 (N_29047,N_28414,N_28324);
nor U29048 (N_29048,N_28611,N_28376);
nand U29049 (N_29049,N_28544,N_28234);
nand U29050 (N_29050,N_28696,N_28666);
xor U29051 (N_29051,N_28634,N_28560);
xor U29052 (N_29052,N_28679,N_28229);
nor U29053 (N_29053,N_28792,N_28300);
nand U29054 (N_29054,N_28569,N_28505);
or U29055 (N_29055,N_28669,N_28353);
xnor U29056 (N_29056,N_28598,N_28708);
nor U29057 (N_29057,N_28369,N_28659);
or U29058 (N_29058,N_28551,N_28614);
nand U29059 (N_29059,N_28327,N_28619);
or U29060 (N_29060,N_28787,N_28710);
nand U29061 (N_29061,N_28767,N_28563);
or U29062 (N_29062,N_28748,N_28520);
xor U29063 (N_29063,N_28556,N_28514);
and U29064 (N_29064,N_28224,N_28506);
and U29065 (N_29065,N_28577,N_28418);
nand U29066 (N_29066,N_28527,N_28755);
xnor U29067 (N_29067,N_28266,N_28317);
and U29068 (N_29068,N_28492,N_28239);
nand U29069 (N_29069,N_28780,N_28622);
nor U29070 (N_29070,N_28393,N_28298);
nor U29071 (N_29071,N_28447,N_28206);
nand U29072 (N_29072,N_28358,N_28715);
nor U29073 (N_29073,N_28288,N_28478);
and U29074 (N_29074,N_28251,N_28262);
and U29075 (N_29075,N_28479,N_28515);
xor U29076 (N_29076,N_28301,N_28511);
or U29077 (N_29077,N_28227,N_28694);
or U29078 (N_29078,N_28723,N_28793);
nor U29079 (N_29079,N_28333,N_28528);
nor U29080 (N_29080,N_28783,N_28490);
and U29081 (N_29081,N_28410,N_28390);
or U29082 (N_29082,N_28389,N_28341);
and U29083 (N_29083,N_28213,N_28400);
xnor U29084 (N_29084,N_28549,N_28592);
or U29085 (N_29085,N_28744,N_28308);
and U29086 (N_29086,N_28673,N_28281);
nand U29087 (N_29087,N_28465,N_28323);
and U29088 (N_29088,N_28415,N_28721);
nor U29089 (N_29089,N_28650,N_28799);
nand U29090 (N_29090,N_28408,N_28348);
or U29091 (N_29091,N_28403,N_28545);
nand U29092 (N_29092,N_28701,N_28566);
and U29093 (N_29093,N_28625,N_28311);
xor U29094 (N_29094,N_28501,N_28278);
xnor U29095 (N_29095,N_28735,N_28500);
or U29096 (N_29096,N_28581,N_28512);
xor U29097 (N_29097,N_28523,N_28745);
or U29098 (N_29098,N_28264,N_28230);
nor U29099 (N_29099,N_28689,N_28335);
nor U29100 (N_29100,N_28317,N_28308);
nor U29101 (N_29101,N_28774,N_28333);
xnor U29102 (N_29102,N_28545,N_28450);
nand U29103 (N_29103,N_28230,N_28698);
and U29104 (N_29104,N_28254,N_28439);
and U29105 (N_29105,N_28525,N_28689);
xor U29106 (N_29106,N_28721,N_28723);
nand U29107 (N_29107,N_28391,N_28395);
nor U29108 (N_29108,N_28726,N_28571);
or U29109 (N_29109,N_28608,N_28372);
or U29110 (N_29110,N_28788,N_28425);
and U29111 (N_29111,N_28231,N_28323);
and U29112 (N_29112,N_28442,N_28651);
and U29113 (N_29113,N_28511,N_28652);
nand U29114 (N_29114,N_28593,N_28369);
nand U29115 (N_29115,N_28350,N_28514);
nand U29116 (N_29116,N_28705,N_28565);
or U29117 (N_29117,N_28645,N_28569);
xnor U29118 (N_29118,N_28471,N_28784);
nor U29119 (N_29119,N_28683,N_28686);
or U29120 (N_29120,N_28674,N_28531);
nor U29121 (N_29121,N_28673,N_28455);
nand U29122 (N_29122,N_28677,N_28382);
nor U29123 (N_29123,N_28243,N_28685);
nor U29124 (N_29124,N_28426,N_28211);
or U29125 (N_29125,N_28442,N_28685);
nor U29126 (N_29126,N_28249,N_28489);
nand U29127 (N_29127,N_28536,N_28266);
nand U29128 (N_29128,N_28726,N_28258);
xnor U29129 (N_29129,N_28201,N_28358);
xor U29130 (N_29130,N_28743,N_28429);
nor U29131 (N_29131,N_28527,N_28714);
xnor U29132 (N_29132,N_28419,N_28752);
nand U29133 (N_29133,N_28347,N_28256);
or U29134 (N_29134,N_28590,N_28498);
xnor U29135 (N_29135,N_28294,N_28411);
nand U29136 (N_29136,N_28577,N_28483);
nor U29137 (N_29137,N_28566,N_28787);
nor U29138 (N_29138,N_28208,N_28600);
nand U29139 (N_29139,N_28692,N_28485);
nor U29140 (N_29140,N_28733,N_28540);
nand U29141 (N_29141,N_28345,N_28615);
nor U29142 (N_29142,N_28245,N_28675);
or U29143 (N_29143,N_28434,N_28421);
xnor U29144 (N_29144,N_28447,N_28443);
and U29145 (N_29145,N_28367,N_28772);
or U29146 (N_29146,N_28398,N_28346);
or U29147 (N_29147,N_28294,N_28588);
and U29148 (N_29148,N_28676,N_28497);
nor U29149 (N_29149,N_28365,N_28419);
nand U29150 (N_29150,N_28785,N_28277);
and U29151 (N_29151,N_28685,N_28370);
or U29152 (N_29152,N_28248,N_28441);
nand U29153 (N_29153,N_28337,N_28649);
nand U29154 (N_29154,N_28505,N_28774);
xor U29155 (N_29155,N_28693,N_28733);
nor U29156 (N_29156,N_28271,N_28426);
xnor U29157 (N_29157,N_28536,N_28488);
nand U29158 (N_29158,N_28365,N_28383);
nand U29159 (N_29159,N_28430,N_28262);
and U29160 (N_29160,N_28696,N_28794);
and U29161 (N_29161,N_28549,N_28345);
and U29162 (N_29162,N_28618,N_28788);
nor U29163 (N_29163,N_28264,N_28773);
nand U29164 (N_29164,N_28492,N_28426);
nor U29165 (N_29165,N_28537,N_28512);
or U29166 (N_29166,N_28344,N_28301);
and U29167 (N_29167,N_28362,N_28603);
nor U29168 (N_29168,N_28757,N_28783);
nor U29169 (N_29169,N_28651,N_28301);
or U29170 (N_29170,N_28485,N_28286);
nand U29171 (N_29171,N_28689,N_28477);
nand U29172 (N_29172,N_28344,N_28342);
xnor U29173 (N_29173,N_28512,N_28307);
nor U29174 (N_29174,N_28748,N_28253);
or U29175 (N_29175,N_28601,N_28577);
xnor U29176 (N_29176,N_28270,N_28343);
xor U29177 (N_29177,N_28507,N_28259);
xor U29178 (N_29178,N_28380,N_28668);
nor U29179 (N_29179,N_28722,N_28593);
or U29180 (N_29180,N_28505,N_28272);
xnor U29181 (N_29181,N_28771,N_28759);
or U29182 (N_29182,N_28636,N_28728);
or U29183 (N_29183,N_28626,N_28633);
nor U29184 (N_29184,N_28334,N_28323);
and U29185 (N_29185,N_28575,N_28230);
nand U29186 (N_29186,N_28630,N_28211);
xnor U29187 (N_29187,N_28794,N_28343);
nand U29188 (N_29188,N_28396,N_28579);
or U29189 (N_29189,N_28371,N_28201);
nand U29190 (N_29190,N_28367,N_28256);
nand U29191 (N_29191,N_28471,N_28333);
nor U29192 (N_29192,N_28411,N_28422);
and U29193 (N_29193,N_28609,N_28654);
xnor U29194 (N_29194,N_28428,N_28334);
and U29195 (N_29195,N_28252,N_28516);
nand U29196 (N_29196,N_28239,N_28466);
nor U29197 (N_29197,N_28570,N_28496);
or U29198 (N_29198,N_28650,N_28239);
nor U29199 (N_29199,N_28666,N_28537);
nor U29200 (N_29200,N_28741,N_28365);
or U29201 (N_29201,N_28775,N_28605);
nor U29202 (N_29202,N_28330,N_28539);
and U29203 (N_29203,N_28256,N_28376);
xnor U29204 (N_29204,N_28775,N_28596);
nand U29205 (N_29205,N_28420,N_28264);
and U29206 (N_29206,N_28616,N_28779);
or U29207 (N_29207,N_28729,N_28387);
nor U29208 (N_29208,N_28383,N_28449);
nor U29209 (N_29209,N_28382,N_28582);
nand U29210 (N_29210,N_28252,N_28737);
or U29211 (N_29211,N_28232,N_28261);
and U29212 (N_29212,N_28668,N_28386);
nor U29213 (N_29213,N_28521,N_28298);
nor U29214 (N_29214,N_28205,N_28545);
xor U29215 (N_29215,N_28233,N_28611);
xor U29216 (N_29216,N_28688,N_28496);
nand U29217 (N_29217,N_28450,N_28451);
xnor U29218 (N_29218,N_28267,N_28576);
nand U29219 (N_29219,N_28637,N_28583);
and U29220 (N_29220,N_28385,N_28428);
nor U29221 (N_29221,N_28556,N_28380);
and U29222 (N_29222,N_28767,N_28342);
and U29223 (N_29223,N_28515,N_28529);
and U29224 (N_29224,N_28419,N_28769);
nor U29225 (N_29225,N_28576,N_28648);
nand U29226 (N_29226,N_28743,N_28552);
nand U29227 (N_29227,N_28773,N_28756);
xor U29228 (N_29228,N_28697,N_28609);
and U29229 (N_29229,N_28551,N_28615);
and U29230 (N_29230,N_28636,N_28577);
nand U29231 (N_29231,N_28301,N_28383);
and U29232 (N_29232,N_28568,N_28408);
and U29233 (N_29233,N_28304,N_28788);
and U29234 (N_29234,N_28488,N_28697);
or U29235 (N_29235,N_28357,N_28518);
or U29236 (N_29236,N_28663,N_28696);
xnor U29237 (N_29237,N_28668,N_28754);
and U29238 (N_29238,N_28496,N_28384);
xor U29239 (N_29239,N_28688,N_28300);
or U29240 (N_29240,N_28795,N_28656);
and U29241 (N_29241,N_28382,N_28579);
and U29242 (N_29242,N_28286,N_28258);
and U29243 (N_29243,N_28567,N_28299);
nor U29244 (N_29244,N_28303,N_28498);
or U29245 (N_29245,N_28679,N_28470);
xor U29246 (N_29246,N_28477,N_28759);
or U29247 (N_29247,N_28487,N_28390);
or U29248 (N_29248,N_28795,N_28522);
and U29249 (N_29249,N_28617,N_28638);
nor U29250 (N_29250,N_28636,N_28268);
nand U29251 (N_29251,N_28683,N_28366);
nand U29252 (N_29252,N_28428,N_28716);
or U29253 (N_29253,N_28424,N_28509);
nor U29254 (N_29254,N_28530,N_28559);
nor U29255 (N_29255,N_28437,N_28457);
nand U29256 (N_29256,N_28567,N_28456);
nand U29257 (N_29257,N_28535,N_28351);
and U29258 (N_29258,N_28565,N_28287);
nor U29259 (N_29259,N_28783,N_28631);
and U29260 (N_29260,N_28340,N_28291);
nand U29261 (N_29261,N_28706,N_28604);
or U29262 (N_29262,N_28653,N_28719);
nand U29263 (N_29263,N_28631,N_28508);
xor U29264 (N_29264,N_28625,N_28251);
nor U29265 (N_29265,N_28569,N_28766);
nand U29266 (N_29266,N_28706,N_28449);
nand U29267 (N_29267,N_28768,N_28600);
and U29268 (N_29268,N_28430,N_28504);
xnor U29269 (N_29269,N_28759,N_28627);
and U29270 (N_29270,N_28500,N_28324);
or U29271 (N_29271,N_28757,N_28588);
nand U29272 (N_29272,N_28772,N_28240);
xor U29273 (N_29273,N_28454,N_28673);
nand U29274 (N_29274,N_28775,N_28434);
nand U29275 (N_29275,N_28612,N_28279);
nand U29276 (N_29276,N_28394,N_28316);
or U29277 (N_29277,N_28206,N_28499);
nand U29278 (N_29278,N_28435,N_28442);
nor U29279 (N_29279,N_28627,N_28724);
or U29280 (N_29280,N_28488,N_28437);
xor U29281 (N_29281,N_28531,N_28611);
nor U29282 (N_29282,N_28554,N_28463);
nand U29283 (N_29283,N_28403,N_28227);
xnor U29284 (N_29284,N_28673,N_28731);
or U29285 (N_29285,N_28668,N_28708);
or U29286 (N_29286,N_28680,N_28262);
or U29287 (N_29287,N_28500,N_28298);
xor U29288 (N_29288,N_28471,N_28627);
or U29289 (N_29289,N_28635,N_28494);
or U29290 (N_29290,N_28793,N_28233);
nand U29291 (N_29291,N_28250,N_28764);
nor U29292 (N_29292,N_28790,N_28642);
nand U29293 (N_29293,N_28447,N_28344);
xnor U29294 (N_29294,N_28784,N_28478);
or U29295 (N_29295,N_28629,N_28609);
and U29296 (N_29296,N_28384,N_28285);
nand U29297 (N_29297,N_28220,N_28503);
xor U29298 (N_29298,N_28684,N_28284);
and U29299 (N_29299,N_28470,N_28745);
and U29300 (N_29300,N_28211,N_28557);
and U29301 (N_29301,N_28596,N_28714);
xor U29302 (N_29302,N_28583,N_28790);
or U29303 (N_29303,N_28252,N_28695);
xor U29304 (N_29304,N_28309,N_28473);
xnor U29305 (N_29305,N_28578,N_28639);
or U29306 (N_29306,N_28378,N_28575);
nand U29307 (N_29307,N_28764,N_28342);
nand U29308 (N_29308,N_28781,N_28737);
or U29309 (N_29309,N_28369,N_28653);
xor U29310 (N_29310,N_28323,N_28661);
nand U29311 (N_29311,N_28459,N_28737);
or U29312 (N_29312,N_28739,N_28525);
or U29313 (N_29313,N_28248,N_28297);
and U29314 (N_29314,N_28695,N_28426);
or U29315 (N_29315,N_28680,N_28759);
xor U29316 (N_29316,N_28345,N_28752);
nor U29317 (N_29317,N_28690,N_28578);
nor U29318 (N_29318,N_28231,N_28643);
or U29319 (N_29319,N_28351,N_28329);
xor U29320 (N_29320,N_28510,N_28305);
nor U29321 (N_29321,N_28307,N_28681);
and U29322 (N_29322,N_28250,N_28651);
or U29323 (N_29323,N_28612,N_28608);
nand U29324 (N_29324,N_28724,N_28295);
xor U29325 (N_29325,N_28304,N_28611);
nor U29326 (N_29326,N_28741,N_28254);
and U29327 (N_29327,N_28644,N_28358);
or U29328 (N_29328,N_28704,N_28342);
and U29329 (N_29329,N_28779,N_28680);
or U29330 (N_29330,N_28664,N_28525);
or U29331 (N_29331,N_28604,N_28507);
nand U29332 (N_29332,N_28548,N_28250);
nand U29333 (N_29333,N_28734,N_28492);
xor U29334 (N_29334,N_28797,N_28420);
xor U29335 (N_29335,N_28769,N_28391);
nor U29336 (N_29336,N_28648,N_28428);
nand U29337 (N_29337,N_28359,N_28246);
nor U29338 (N_29338,N_28675,N_28579);
nor U29339 (N_29339,N_28513,N_28741);
nor U29340 (N_29340,N_28229,N_28370);
nor U29341 (N_29341,N_28577,N_28614);
nand U29342 (N_29342,N_28727,N_28655);
nand U29343 (N_29343,N_28539,N_28576);
xor U29344 (N_29344,N_28573,N_28326);
nor U29345 (N_29345,N_28209,N_28797);
nor U29346 (N_29346,N_28407,N_28485);
nand U29347 (N_29347,N_28649,N_28712);
nor U29348 (N_29348,N_28548,N_28723);
nor U29349 (N_29349,N_28281,N_28729);
xor U29350 (N_29350,N_28631,N_28228);
nor U29351 (N_29351,N_28370,N_28761);
and U29352 (N_29352,N_28709,N_28712);
nand U29353 (N_29353,N_28538,N_28442);
or U29354 (N_29354,N_28687,N_28363);
and U29355 (N_29355,N_28357,N_28418);
nand U29356 (N_29356,N_28777,N_28508);
and U29357 (N_29357,N_28783,N_28798);
or U29358 (N_29358,N_28334,N_28468);
nor U29359 (N_29359,N_28224,N_28478);
and U29360 (N_29360,N_28655,N_28671);
nand U29361 (N_29361,N_28277,N_28754);
xnor U29362 (N_29362,N_28400,N_28537);
nor U29363 (N_29363,N_28455,N_28567);
and U29364 (N_29364,N_28748,N_28564);
and U29365 (N_29365,N_28303,N_28791);
or U29366 (N_29366,N_28419,N_28773);
and U29367 (N_29367,N_28536,N_28675);
nand U29368 (N_29368,N_28344,N_28260);
and U29369 (N_29369,N_28430,N_28479);
and U29370 (N_29370,N_28252,N_28754);
xnor U29371 (N_29371,N_28553,N_28647);
nand U29372 (N_29372,N_28212,N_28338);
nor U29373 (N_29373,N_28774,N_28571);
or U29374 (N_29374,N_28650,N_28360);
nor U29375 (N_29375,N_28701,N_28433);
nand U29376 (N_29376,N_28509,N_28724);
xor U29377 (N_29377,N_28327,N_28490);
xnor U29378 (N_29378,N_28247,N_28480);
xor U29379 (N_29379,N_28756,N_28658);
xnor U29380 (N_29380,N_28483,N_28740);
nor U29381 (N_29381,N_28633,N_28285);
or U29382 (N_29382,N_28636,N_28489);
or U29383 (N_29383,N_28518,N_28484);
nor U29384 (N_29384,N_28686,N_28327);
and U29385 (N_29385,N_28796,N_28733);
nand U29386 (N_29386,N_28284,N_28730);
or U29387 (N_29387,N_28474,N_28670);
nand U29388 (N_29388,N_28476,N_28395);
and U29389 (N_29389,N_28240,N_28720);
or U29390 (N_29390,N_28310,N_28450);
and U29391 (N_29391,N_28464,N_28685);
nand U29392 (N_29392,N_28787,N_28738);
xnor U29393 (N_29393,N_28764,N_28262);
or U29394 (N_29394,N_28439,N_28288);
or U29395 (N_29395,N_28671,N_28756);
xor U29396 (N_29396,N_28487,N_28508);
or U29397 (N_29397,N_28569,N_28529);
nand U29398 (N_29398,N_28692,N_28404);
xor U29399 (N_29399,N_28272,N_28598);
or U29400 (N_29400,N_29035,N_28803);
nor U29401 (N_29401,N_28943,N_29355);
or U29402 (N_29402,N_28997,N_29166);
or U29403 (N_29403,N_28884,N_29347);
or U29404 (N_29404,N_29230,N_28951);
xnor U29405 (N_29405,N_29184,N_28806);
xnor U29406 (N_29406,N_29128,N_28933);
xnor U29407 (N_29407,N_29129,N_29140);
xnor U29408 (N_29408,N_29221,N_29173);
xnor U29409 (N_29409,N_29278,N_28985);
nor U29410 (N_29410,N_28839,N_28905);
and U29411 (N_29411,N_29238,N_29310);
or U29412 (N_29412,N_28804,N_28996);
or U29413 (N_29413,N_29254,N_29303);
and U29414 (N_29414,N_28813,N_29387);
xor U29415 (N_29415,N_29364,N_29397);
xor U29416 (N_29416,N_28827,N_29218);
nand U29417 (N_29417,N_28849,N_29257);
nand U29418 (N_29418,N_29039,N_28970);
xor U29419 (N_29419,N_28936,N_29135);
or U29420 (N_29420,N_28980,N_28807);
xnor U29421 (N_29421,N_28969,N_29088);
nand U29422 (N_29422,N_29319,N_29082);
nand U29423 (N_29423,N_29064,N_28895);
nand U29424 (N_29424,N_29148,N_29106);
nand U29425 (N_29425,N_29248,N_29292);
or U29426 (N_29426,N_28994,N_29205);
or U29427 (N_29427,N_29015,N_29350);
nand U29428 (N_29428,N_28928,N_29127);
or U29429 (N_29429,N_28954,N_29107);
or U29430 (N_29430,N_29019,N_29044);
nand U29431 (N_29431,N_29200,N_28914);
nand U29432 (N_29432,N_29378,N_29045);
nand U29433 (N_29433,N_29123,N_29268);
xor U29434 (N_29434,N_28901,N_29256);
or U29435 (N_29435,N_28992,N_29309);
nor U29436 (N_29436,N_28902,N_29056);
nand U29437 (N_29437,N_29264,N_29185);
nand U29438 (N_29438,N_28857,N_28979);
and U29439 (N_29439,N_28946,N_29004);
or U29440 (N_29440,N_29014,N_28856);
nand U29441 (N_29441,N_28853,N_29274);
nand U29442 (N_29442,N_29149,N_28879);
nor U29443 (N_29443,N_28848,N_29276);
and U29444 (N_29444,N_29340,N_29258);
nand U29445 (N_29445,N_29333,N_28931);
or U29446 (N_29446,N_29161,N_29052);
xor U29447 (N_29447,N_29339,N_29178);
and U29448 (N_29448,N_29365,N_29066);
xor U29449 (N_29449,N_29022,N_28859);
xor U29450 (N_29450,N_29147,N_29210);
nand U29451 (N_29451,N_28843,N_29059);
or U29452 (N_29452,N_28805,N_29020);
nand U29453 (N_29453,N_28810,N_28872);
nand U29454 (N_29454,N_29115,N_29001);
or U29455 (N_29455,N_29202,N_29065);
and U29456 (N_29456,N_29380,N_29083);
nand U29457 (N_29457,N_28941,N_28820);
nand U29458 (N_29458,N_28833,N_29219);
nand U29459 (N_29459,N_28904,N_28973);
and U29460 (N_29460,N_29377,N_29227);
or U29461 (N_29461,N_28938,N_29138);
nand U29462 (N_29462,N_29116,N_29030);
nor U29463 (N_29463,N_29335,N_28865);
xor U29464 (N_29464,N_28814,N_29026);
or U29465 (N_29465,N_29118,N_28966);
and U29466 (N_29466,N_29099,N_28975);
xor U29467 (N_29467,N_28912,N_29192);
xnor U29468 (N_29468,N_29325,N_29301);
and U29469 (N_29469,N_29376,N_29057);
xnor U29470 (N_29470,N_29117,N_28957);
nor U29471 (N_29471,N_28836,N_29121);
or U29472 (N_29472,N_28845,N_29240);
xnor U29473 (N_29473,N_29042,N_29299);
nand U29474 (N_29474,N_29196,N_29320);
nor U29475 (N_29475,N_28982,N_29308);
nor U29476 (N_29476,N_29157,N_29295);
or U29477 (N_29477,N_28801,N_29002);
or U29478 (N_29478,N_29273,N_29012);
xnor U29479 (N_29479,N_29220,N_29396);
nand U29480 (N_29480,N_28963,N_28952);
nand U29481 (N_29481,N_29047,N_29233);
nand U29482 (N_29482,N_29162,N_28923);
and U29483 (N_29483,N_28984,N_29009);
or U29484 (N_29484,N_28882,N_29055);
and U29485 (N_29485,N_29126,N_28911);
and U29486 (N_29486,N_29150,N_29244);
nor U29487 (N_29487,N_29291,N_29062);
or U29488 (N_29488,N_28830,N_29086);
and U29489 (N_29489,N_29224,N_28886);
or U29490 (N_29490,N_29029,N_29368);
nand U29491 (N_29491,N_29006,N_29269);
xnor U29492 (N_29492,N_29089,N_29249);
or U29493 (N_29493,N_28986,N_29179);
or U29494 (N_29494,N_29362,N_28942);
nor U29495 (N_29495,N_29261,N_29262);
or U29496 (N_29496,N_28892,N_29112);
nor U29497 (N_29497,N_28959,N_28903);
nand U29498 (N_29498,N_29027,N_29061);
nor U29499 (N_29499,N_29145,N_29213);
nand U29500 (N_29500,N_29208,N_29399);
and U29501 (N_29501,N_29383,N_29316);
or U29502 (N_29502,N_28965,N_29144);
and U29503 (N_29503,N_29051,N_29102);
and U29504 (N_29504,N_29090,N_28821);
xnor U29505 (N_29505,N_28919,N_29236);
nor U29506 (N_29506,N_29255,N_28876);
xnor U29507 (N_29507,N_28922,N_29391);
xor U29508 (N_29508,N_28899,N_29021);
nand U29509 (N_29509,N_28907,N_29193);
xnor U29510 (N_29510,N_29197,N_29188);
nor U29511 (N_29511,N_28971,N_29160);
nor U29512 (N_29512,N_28953,N_29237);
nand U29513 (N_29513,N_29330,N_29252);
xnor U29514 (N_29514,N_29091,N_28840);
and U29515 (N_29515,N_28877,N_28940);
nor U29516 (N_29516,N_28925,N_29098);
nand U29517 (N_29517,N_29040,N_29060);
xnor U29518 (N_29518,N_29114,N_29007);
or U29519 (N_29519,N_28816,N_28878);
nand U29520 (N_29520,N_29398,N_29351);
or U29521 (N_29521,N_29189,N_29395);
nor U29522 (N_29522,N_28823,N_28866);
or U29523 (N_29523,N_28841,N_29013);
xnor U29524 (N_29524,N_29074,N_28811);
xor U29525 (N_29525,N_28898,N_29263);
nor U29526 (N_29526,N_29000,N_29212);
nor U29527 (N_29527,N_29369,N_28929);
or U29528 (N_29528,N_29180,N_29172);
and U29529 (N_29529,N_29113,N_29169);
and U29530 (N_29530,N_29282,N_28875);
xor U29531 (N_29531,N_29209,N_29287);
nor U29532 (N_29532,N_28838,N_29294);
xor U29533 (N_29533,N_28835,N_28860);
or U29534 (N_29534,N_29228,N_29232);
or U29535 (N_29535,N_28855,N_29008);
and U29536 (N_29536,N_28908,N_29302);
and U29537 (N_29537,N_29037,N_28939);
and U29538 (N_29538,N_29036,N_29242);
or U29539 (N_29539,N_29379,N_29307);
nor U29540 (N_29540,N_29375,N_29080);
xor U29541 (N_29541,N_28837,N_29337);
xor U29542 (N_29542,N_29229,N_29361);
nand U29543 (N_29543,N_28958,N_28854);
nand U29544 (N_29544,N_29217,N_28968);
nor U29545 (N_29545,N_29275,N_29370);
nand U29546 (N_29546,N_29298,N_28888);
nand U29547 (N_29547,N_29181,N_29100);
nand U29548 (N_29548,N_28909,N_28873);
and U29549 (N_29549,N_29314,N_28846);
nand U29550 (N_29550,N_29158,N_29031);
xnor U29551 (N_29551,N_29215,N_29342);
and U29552 (N_29552,N_29131,N_29300);
nand U29553 (N_29553,N_29211,N_29348);
and U29554 (N_29554,N_28978,N_29078);
xor U29555 (N_29555,N_29389,N_29321);
and U29556 (N_29556,N_28847,N_29054);
nor U29557 (N_29557,N_28812,N_29283);
and U29558 (N_29558,N_29304,N_29293);
nand U29559 (N_29559,N_29329,N_29203);
nand U29560 (N_29560,N_29214,N_29267);
xnor U29561 (N_29561,N_29344,N_29124);
nor U29562 (N_29562,N_28864,N_29095);
and U29563 (N_29563,N_28981,N_29394);
or U29564 (N_29564,N_29324,N_28871);
xnor U29565 (N_29565,N_28937,N_29120);
and U29566 (N_29566,N_29289,N_29352);
or U29567 (N_29567,N_28834,N_28817);
nor U29568 (N_29568,N_29048,N_28967);
and U29569 (N_29569,N_29250,N_29315);
and U29570 (N_29570,N_29167,N_29195);
nand U29571 (N_29571,N_29201,N_29143);
and U29572 (N_29572,N_28891,N_29260);
and U29573 (N_29573,N_29306,N_28956);
and U29574 (N_29574,N_29392,N_28927);
nand U29575 (N_29575,N_29171,N_29170);
and U29576 (N_29576,N_29356,N_28990);
xnor U29577 (N_29577,N_29371,N_29103);
nor U29578 (N_29578,N_28945,N_29005);
xnor U29579 (N_29579,N_28831,N_28883);
xnor U29580 (N_29580,N_28993,N_29345);
or U29581 (N_29581,N_29104,N_28972);
and U29582 (N_29582,N_29341,N_29385);
or U29583 (N_29583,N_29288,N_28822);
xor U29584 (N_29584,N_29312,N_28852);
xnor U29585 (N_29585,N_29092,N_28976);
xor U29586 (N_29586,N_29024,N_29041);
or U29587 (N_29587,N_28832,N_28960);
nand U29588 (N_29588,N_28964,N_28863);
nor U29589 (N_29589,N_29108,N_29334);
xnor U29590 (N_29590,N_29245,N_29087);
nand U29591 (N_29591,N_29084,N_28800);
or U29592 (N_29592,N_29073,N_28924);
nor U29593 (N_29593,N_28988,N_29382);
nand U29594 (N_29594,N_29194,N_29243);
and U29595 (N_29595,N_29049,N_29141);
and U29596 (N_29596,N_29216,N_29381);
nor U29597 (N_29597,N_29374,N_29327);
and U29598 (N_29598,N_28913,N_29190);
or U29599 (N_29599,N_28896,N_28881);
nand U29600 (N_29600,N_29253,N_28915);
nand U29601 (N_29601,N_29155,N_29096);
nor U29602 (N_29602,N_29270,N_29038);
and U29603 (N_29603,N_28935,N_28867);
nor U29604 (N_29604,N_29175,N_29182);
or U29605 (N_29605,N_28802,N_29093);
or U29606 (N_29606,N_29367,N_29165);
nor U29607 (N_29607,N_29280,N_29046);
nor U29608 (N_29608,N_29234,N_28987);
and U29609 (N_29609,N_29226,N_29109);
and U29610 (N_29610,N_29317,N_29272);
xor U29611 (N_29611,N_28916,N_29183);
and U29612 (N_29612,N_29266,N_28851);
nor U29613 (N_29613,N_28889,N_29017);
and U29614 (N_29614,N_29011,N_28819);
or U29615 (N_29615,N_28815,N_29346);
and U29616 (N_29616,N_29336,N_28930);
and U29617 (N_29617,N_29393,N_29139);
and U29618 (N_29618,N_29032,N_29153);
nand U29619 (N_29619,N_29366,N_28885);
xor U29620 (N_29620,N_28917,N_28858);
xnor U29621 (N_29621,N_29111,N_29204);
nor U29622 (N_29622,N_28842,N_29286);
nand U29623 (N_29623,N_29070,N_28950);
xnor U29624 (N_29624,N_29318,N_29296);
nand U29625 (N_29625,N_29277,N_29094);
and U29626 (N_29626,N_28989,N_28890);
xor U29627 (N_29627,N_29069,N_28894);
and U29628 (N_29628,N_29177,N_29132);
xnor U29629 (N_29629,N_29353,N_29284);
and U29630 (N_29630,N_29133,N_28995);
nand U29631 (N_29631,N_29290,N_29360);
and U29632 (N_29632,N_29168,N_29328);
or U29633 (N_29633,N_28809,N_29372);
nand U29634 (N_29634,N_28991,N_29297);
and U29635 (N_29635,N_29174,N_28844);
nor U29636 (N_29636,N_28961,N_29034);
and U29637 (N_29637,N_28897,N_29358);
nand U29638 (N_29638,N_29225,N_28880);
xor U29639 (N_29639,N_29222,N_29010);
or U29640 (N_29640,N_29063,N_29068);
or U29641 (N_29641,N_29305,N_29357);
or U29642 (N_29642,N_29259,N_29338);
and U29643 (N_29643,N_29223,N_29313);
or U29644 (N_29644,N_29119,N_28932);
nand U29645 (N_29645,N_29373,N_29206);
or U29646 (N_29646,N_29271,N_28918);
nand U29647 (N_29647,N_29207,N_28921);
or U29648 (N_29648,N_29105,N_29281);
nor U29649 (N_29649,N_29146,N_28862);
or U29650 (N_29650,N_29359,N_29101);
nand U29651 (N_29651,N_29097,N_29187);
or U29652 (N_29652,N_29043,N_29363);
nand U29653 (N_29653,N_28934,N_29331);
xor U29654 (N_29654,N_29050,N_29349);
xnor U29655 (N_29655,N_29279,N_29390);
nand U29656 (N_29656,N_29154,N_28977);
nand U29657 (N_29657,N_29134,N_28983);
nand U29658 (N_29658,N_29075,N_29122);
nor U29659 (N_29659,N_28910,N_29053);
nand U29660 (N_29660,N_29186,N_29354);
and U29661 (N_29661,N_28944,N_29311);
and U29662 (N_29662,N_29231,N_28870);
nor U29663 (N_29663,N_28949,N_28893);
xor U29664 (N_29664,N_29142,N_28926);
or U29665 (N_29665,N_29198,N_28829);
nand U29666 (N_29666,N_29191,N_29003);
nor U29667 (N_29667,N_29343,N_29025);
nor U29668 (N_29668,N_29071,N_29023);
or U29669 (N_29669,N_29159,N_29058);
or U29670 (N_29670,N_29388,N_28826);
xnor U29671 (N_29671,N_28824,N_29136);
nand U29672 (N_29672,N_29076,N_28869);
nor U29673 (N_29673,N_29033,N_28948);
or U29674 (N_29674,N_29018,N_29332);
or U29675 (N_29675,N_28828,N_29285);
xnor U29676 (N_29676,N_29199,N_29164);
xnor U29677 (N_29677,N_28962,N_28861);
nor U29678 (N_29678,N_28998,N_28808);
nor U29679 (N_29679,N_29163,N_28999);
nor U29680 (N_29680,N_29067,N_29085);
xor U29681 (N_29681,N_28947,N_28900);
and U29682 (N_29682,N_28874,N_29077);
and U29683 (N_29683,N_29176,N_29028);
xor U29684 (N_29684,N_29156,N_29079);
nor U29685 (N_29685,N_29110,N_28818);
or U29686 (N_29686,N_28825,N_28850);
or U29687 (N_29687,N_28974,N_29326);
and U29688 (N_29688,N_28920,N_28955);
nor U29689 (N_29689,N_29137,N_29081);
nor U29690 (N_29690,N_29323,N_29130);
xnor U29691 (N_29691,N_29239,N_29151);
xnor U29692 (N_29692,N_28868,N_29386);
nand U29693 (N_29693,N_28887,N_29247);
and U29694 (N_29694,N_29125,N_29152);
xnor U29695 (N_29695,N_29384,N_29072);
and U29696 (N_29696,N_29265,N_28906);
nor U29697 (N_29697,N_29241,N_29246);
and U29698 (N_29698,N_29016,N_29235);
nand U29699 (N_29699,N_29251,N_29322);
xor U29700 (N_29700,N_28937,N_29303);
nor U29701 (N_29701,N_29155,N_28913);
and U29702 (N_29702,N_29120,N_28828);
xor U29703 (N_29703,N_29373,N_29335);
xnor U29704 (N_29704,N_29305,N_29191);
nor U29705 (N_29705,N_28998,N_29060);
and U29706 (N_29706,N_29199,N_28988);
xnor U29707 (N_29707,N_28926,N_29287);
xnor U29708 (N_29708,N_29341,N_29271);
nand U29709 (N_29709,N_29170,N_29254);
and U29710 (N_29710,N_29379,N_29354);
xor U29711 (N_29711,N_29185,N_28975);
nor U29712 (N_29712,N_29230,N_29332);
or U29713 (N_29713,N_29383,N_29110);
and U29714 (N_29714,N_29293,N_28952);
xor U29715 (N_29715,N_29248,N_28959);
or U29716 (N_29716,N_29084,N_29159);
nor U29717 (N_29717,N_28993,N_29311);
and U29718 (N_29718,N_29291,N_29253);
or U29719 (N_29719,N_28941,N_29375);
xor U29720 (N_29720,N_29249,N_29050);
or U29721 (N_29721,N_29277,N_29323);
nand U29722 (N_29722,N_28859,N_28977);
nand U29723 (N_29723,N_28955,N_28861);
nor U29724 (N_29724,N_28907,N_29367);
nand U29725 (N_29725,N_28833,N_29255);
and U29726 (N_29726,N_28902,N_29382);
nor U29727 (N_29727,N_28984,N_29287);
xnor U29728 (N_29728,N_29185,N_28888);
or U29729 (N_29729,N_29079,N_28908);
or U29730 (N_29730,N_29368,N_29297);
and U29731 (N_29731,N_29021,N_28967);
or U29732 (N_29732,N_29258,N_29098);
nor U29733 (N_29733,N_28891,N_28893);
nand U29734 (N_29734,N_29015,N_28939);
and U29735 (N_29735,N_29285,N_29091);
and U29736 (N_29736,N_28941,N_28882);
xnor U29737 (N_29737,N_29036,N_29051);
and U29738 (N_29738,N_29217,N_29054);
nor U29739 (N_29739,N_29020,N_28988);
nand U29740 (N_29740,N_29089,N_28913);
or U29741 (N_29741,N_29057,N_29378);
nand U29742 (N_29742,N_28850,N_29232);
nor U29743 (N_29743,N_29003,N_29061);
or U29744 (N_29744,N_29364,N_29209);
nand U29745 (N_29745,N_29254,N_28964);
and U29746 (N_29746,N_29296,N_28913);
and U29747 (N_29747,N_29212,N_29075);
or U29748 (N_29748,N_29140,N_28817);
nor U29749 (N_29749,N_28932,N_28856);
nor U29750 (N_29750,N_29193,N_28800);
nor U29751 (N_29751,N_29017,N_29029);
and U29752 (N_29752,N_29201,N_28864);
or U29753 (N_29753,N_29260,N_28897);
xnor U29754 (N_29754,N_29123,N_29391);
xor U29755 (N_29755,N_29214,N_28977);
nor U29756 (N_29756,N_29258,N_29281);
nor U29757 (N_29757,N_28953,N_29120);
or U29758 (N_29758,N_28930,N_29297);
or U29759 (N_29759,N_28871,N_29137);
or U29760 (N_29760,N_29023,N_29139);
nor U29761 (N_29761,N_28819,N_29204);
nand U29762 (N_29762,N_29314,N_28877);
and U29763 (N_29763,N_28989,N_28883);
nor U29764 (N_29764,N_29147,N_29039);
xor U29765 (N_29765,N_29299,N_28992);
nand U29766 (N_29766,N_28951,N_29166);
xor U29767 (N_29767,N_29145,N_29016);
or U29768 (N_29768,N_29167,N_29328);
nor U29769 (N_29769,N_29333,N_29198);
nand U29770 (N_29770,N_29299,N_29149);
and U29771 (N_29771,N_28845,N_29064);
and U29772 (N_29772,N_28912,N_29246);
or U29773 (N_29773,N_29269,N_29146);
xnor U29774 (N_29774,N_28802,N_28917);
nand U29775 (N_29775,N_29359,N_28838);
nand U29776 (N_29776,N_29029,N_29271);
and U29777 (N_29777,N_29019,N_28835);
xor U29778 (N_29778,N_29047,N_28923);
xor U29779 (N_29779,N_29378,N_28807);
nor U29780 (N_29780,N_29254,N_29164);
and U29781 (N_29781,N_29342,N_29177);
or U29782 (N_29782,N_29269,N_29124);
nor U29783 (N_29783,N_28808,N_29034);
and U29784 (N_29784,N_28860,N_29101);
xnor U29785 (N_29785,N_29095,N_28942);
xnor U29786 (N_29786,N_29171,N_29031);
nor U29787 (N_29787,N_28824,N_29078);
and U29788 (N_29788,N_29228,N_29040);
nand U29789 (N_29789,N_29134,N_29082);
and U29790 (N_29790,N_28877,N_29296);
or U29791 (N_29791,N_28877,N_28985);
nand U29792 (N_29792,N_28831,N_29152);
xnor U29793 (N_29793,N_29230,N_29228);
nand U29794 (N_29794,N_29133,N_29267);
nor U29795 (N_29795,N_28906,N_28919);
nand U29796 (N_29796,N_28877,N_29001);
nand U29797 (N_29797,N_29281,N_28975);
nor U29798 (N_29798,N_29134,N_29200);
nor U29799 (N_29799,N_29328,N_28889);
nand U29800 (N_29800,N_28894,N_29211);
or U29801 (N_29801,N_29112,N_28937);
or U29802 (N_29802,N_29099,N_28834);
and U29803 (N_29803,N_29381,N_28804);
or U29804 (N_29804,N_29111,N_29374);
xor U29805 (N_29805,N_29374,N_28893);
nor U29806 (N_29806,N_28841,N_29340);
nand U29807 (N_29807,N_28878,N_29094);
and U29808 (N_29808,N_28940,N_28897);
xor U29809 (N_29809,N_29094,N_28897);
or U29810 (N_29810,N_29362,N_28819);
nand U29811 (N_29811,N_29393,N_29277);
xor U29812 (N_29812,N_29072,N_28902);
nand U29813 (N_29813,N_28837,N_28964);
and U29814 (N_29814,N_29119,N_28997);
xnor U29815 (N_29815,N_28880,N_28972);
nand U29816 (N_29816,N_28863,N_28883);
or U29817 (N_29817,N_29045,N_28878);
or U29818 (N_29818,N_28935,N_29339);
and U29819 (N_29819,N_29135,N_28907);
or U29820 (N_29820,N_29111,N_28913);
and U29821 (N_29821,N_29079,N_28981);
xnor U29822 (N_29822,N_29258,N_28852);
xnor U29823 (N_29823,N_29187,N_29162);
nor U29824 (N_29824,N_29235,N_29057);
xnor U29825 (N_29825,N_29237,N_29227);
and U29826 (N_29826,N_29249,N_29188);
or U29827 (N_29827,N_28862,N_29125);
nand U29828 (N_29828,N_29309,N_29322);
and U29829 (N_29829,N_29315,N_29084);
or U29830 (N_29830,N_29084,N_28808);
or U29831 (N_29831,N_29296,N_29025);
or U29832 (N_29832,N_29108,N_29085);
or U29833 (N_29833,N_29103,N_29039);
or U29834 (N_29834,N_29236,N_28842);
xor U29835 (N_29835,N_28846,N_29193);
nor U29836 (N_29836,N_28989,N_28939);
or U29837 (N_29837,N_29046,N_29244);
nor U29838 (N_29838,N_29382,N_29332);
and U29839 (N_29839,N_28992,N_29313);
nand U29840 (N_29840,N_29279,N_28954);
xor U29841 (N_29841,N_28865,N_29171);
or U29842 (N_29842,N_28949,N_28947);
xnor U29843 (N_29843,N_28975,N_29315);
nor U29844 (N_29844,N_28950,N_29206);
and U29845 (N_29845,N_28967,N_29011);
and U29846 (N_29846,N_29314,N_29024);
and U29847 (N_29847,N_29335,N_29217);
nor U29848 (N_29848,N_29015,N_29190);
or U29849 (N_29849,N_28834,N_29008);
nand U29850 (N_29850,N_29234,N_29002);
and U29851 (N_29851,N_29208,N_28809);
or U29852 (N_29852,N_29379,N_28999);
or U29853 (N_29853,N_29190,N_29048);
nand U29854 (N_29854,N_29195,N_28826);
xor U29855 (N_29855,N_29140,N_29121);
nor U29856 (N_29856,N_29389,N_29018);
nor U29857 (N_29857,N_28995,N_28824);
nand U29858 (N_29858,N_29272,N_29006);
nor U29859 (N_29859,N_28804,N_29073);
or U29860 (N_29860,N_28890,N_29374);
and U29861 (N_29861,N_28992,N_28916);
nand U29862 (N_29862,N_29075,N_29366);
xor U29863 (N_29863,N_29074,N_29183);
nor U29864 (N_29864,N_28806,N_28880);
nor U29865 (N_29865,N_29139,N_29225);
nand U29866 (N_29866,N_29299,N_28815);
nor U29867 (N_29867,N_29229,N_29115);
xnor U29868 (N_29868,N_29052,N_28859);
and U29869 (N_29869,N_29250,N_29187);
and U29870 (N_29870,N_29076,N_28949);
or U29871 (N_29871,N_28830,N_29264);
or U29872 (N_29872,N_28898,N_29281);
nand U29873 (N_29873,N_29344,N_28978);
nand U29874 (N_29874,N_29338,N_29133);
nand U29875 (N_29875,N_29028,N_29090);
and U29876 (N_29876,N_29258,N_28812);
nor U29877 (N_29877,N_29136,N_29130);
or U29878 (N_29878,N_29045,N_28978);
nor U29879 (N_29879,N_29319,N_29031);
and U29880 (N_29880,N_29004,N_28889);
xor U29881 (N_29881,N_29214,N_28999);
and U29882 (N_29882,N_28901,N_29040);
xor U29883 (N_29883,N_29071,N_29389);
or U29884 (N_29884,N_29000,N_29328);
nand U29885 (N_29885,N_29153,N_28826);
xor U29886 (N_29886,N_28958,N_28913);
nor U29887 (N_29887,N_28842,N_28923);
xnor U29888 (N_29888,N_29034,N_29355);
xnor U29889 (N_29889,N_29181,N_29061);
xor U29890 (N_29890,N_28992,N_29389);
nand U29891 (N_29891,N_29052,N_29056);
and U29892 (N_29892,N_28968,N_29140);
xor U29893 (N_29893,N_28958,N_28815);
xor U29894 (N_29894,N_28891,N_29185);
and U29895 (N_29895,N_29192,N_29071);
nor U29896 (N_29896,N_29197,N_29155);
nand U29897 (N_29897,N_29384,N_29329);
nand U29898 (N_29898,N_29076,N_29275);
xor U29899 (N_29899,N_29166,N_28851);
and U29900 (N_29900,N_28829,N_29086);
nand U29901 (N_29901,N_29152,N_29102);
nor U29902 (N_29902,N_28801,N_29179);
nor U29903 (N_29903,N_28916,N_29086);
or U29904 (N_29904,N_29050,N_29266);
nor U29905 (N_29905,N_28891,N_29066);
and U29906 (N_29906,N_28815,N_29115);
nand U29907 (N_29907,N_29059,N_29348);
nor U29908 (N_29908,N_29058,N_29349);
nand U29909 (N_29909,N_28901,N_29305);
xor U29910 (N_29910,N_29231,N_29176);
nor U29911 (N_29911,N_28965,N_28931);
and U29912 (N_29912,N_28892,N_29359);
nor U29913 (N_29913,N_29238,N_28880);
nor U29914 (N_29914,N_29009,N_29346);
nand U29915 (N_29915,N_28908,N_29036);
or U29916 (N_29916,N_29005,N_29290);
xor U29917 (N_29917,N_29065,N_28911);
nor U29918 (N_29918,N_29333,N_29169);
nor U29919 (N_29919,N_29110,N_29217);
and U29920 (N_29920,N_29361,N_29291);
nand U29921 (N_29921,N_29034,N_28928);
xor U29922 (N_29922,N_29319,N_29336);
and U29923 (N_29923,N_28833,N_29049);
xor U29924 (N_29924,N_29039,N_28862);
xnor U29925 (N_29925,N_29271,N_28965);
nand U29926 (N_29926,N_29163,N_29157);
nand U29927 (N_29927,N_28921,N_28914);
nand U29928 (N_29928,N_28983,N_29358);
nand U29929 (N_29929,N_29008,N_29366);
nor U29930 (N_29930,N_29076,N_28866);
and U29931 (N_29931,N_29239,N_28946);
and U29932 (N_29932,N_29337,N_28818);
nand U29933 (N_29933,N_29128,N_29087);
and U29934 (N_29934,N_29052,N_29005);
xor U29935 (N_29935,N_29350,N_28838);
nand U29936 (N_29936,N_28916,N_29323);
nand U29937 (N_29937,N_29390,N_28860);
or U29938 (N_29938,N_29256,N_28931);
nor U29939 (N_29939,N_28937,N_29316);
or U29940 (N_29940,N_28908,N_29357);
and U29941 (N_29941,N_29279,N_28886);
or U29942 (N_29942,N_29094,N_28851);
xor U29943 (N_29943,N_28949,N_29299);
nor U29944 (N_29944,N_29146,N_29199);
nand U29945 (N_29945,N_29296,N_29170);
and U29946 (N_29946,N_28843,N_28820);
or U29947 (N_29947,N_29120,N_29237);
nor U29948 (N_29948,N_29290,N_28936);
nor U29949 (N_29949,N_29173,N_29178);
xor U29950 (N_29950,N_28995,N_28885);
nor U29951 (N_29951,N_28837,N_29088);
and U29952 (N_29952,N_29341,N_29021);
nand U29953 (N_29953,N_28932,N_29055);
nor U29954 (N_29954,N_28843,N_29014);
nand U29955 (N_29955,N_29302,N_29279);
nand U29956 (N_29956,N_29346,N_29136);
xor U29957 (N_29957,N_29380,N_29234);
nand U29958 (N_29958,N_29318,N_28908);
xnor U29959 (N_29959,N_29328,N_28826);
nand U29960 (N_29960,N_29017,N_29351);
nand U29961 (N_29961,N_29315,N_29366);
nand U29962 (N_29962,N_29150,N_29232);
xor U29963 (N_29963,N_28832,N_28826);
and U29964 (N_29964,N_28851,N_28822);
nor U29965 (N_29965,N_29337,N_29060);
xor U29966 (N_29966,N_29129,N_29398);
nor U29967 (N_29967,N_28908,N_29323);
xor U29968 (N_29968,N_29072,N_29335);
nor U29969 (N_29969,N_28950,N_28881);
and U29970 (N_29970,N_29383,N_28905);
or U29971 (N_29971,N_28857,N_29309);
or U29972 (N_29972,N_29328,N_29122);
xnor U29973 (N_29973,N_28886,N_29294);
nor U29974 (N_29974,N_29325,N_28833);
and U29975 (N_29975,N_29281,N_29334);
or U29976 (N_29976,N_28810,N_29160);
and U29977 (N_29977,N_28844,N_28834);
or U29978 (N_29978,N_29079,N_29118);
nand U29979 (N_29979,N_29384,N_28950);
nand U29980 (N_29980,N_29369,N_29288);
nor U29981 (N_29981,N_28988,N_29215);
or U29982 (N_29982,N_28875,N_29085);
or U29983 (N_29983,N_29150,N_29097);
nand U29984 (N_29984,N_28809,N_29039);
nor U29985 (N_29985,N_29280,N_29383);
nor U29986 (N_29986,N_29024,N_29296);
and U29987 (N_29987,N_29093,N_29143);
and U29988 (N_29988,N_29260,N_29111);
and U29989 (N_29989,N_29019,N_28873);
nand U29990 (N_29990,N_29095,N_28950);
xor U29991 (N_29991,N_28980,N_29343);
and U29992 (N_29992,N_29331,N_29203);
nor U29993 (N_29993,N_29342,N_28962);
xor U29994 (N_29994,N_28826,N_29222);
or U29995 (N_29995,N_28970,N_29153);
nor U29996 (N_29996,N_29371,N_28806);
xnor U29997 (N_29997,N_29398,N_28907);
or U29998 (N_29998,N_28892,N_28823);
nand U29999 (N_29999,N_29395,N_28870);
or UO_0 (O_0,N_29824,N_29642);
nor UO_1 (O_1,N_29817,N_29970);
or UO_2 (O_2,N_29644,N_29945);
xnor UO_3 (O_3,N_29784,N_29818);
or UO_4 (O_4,N_29622,N_29599);
and UO_5 (O_5,N_29861,N_29688);
and UO_6 (O_6,N_29887,N_29496);
nor UO_7 (O_7,N_29550,N_29542);
and UO_8 (O_8,N_29657,N_29422);
nor UO_9 (O_9,N_29503,N_29801);
xor UO_10 (O_10,N_29694,N_29528);
or UO_11 (O_11,N_29572,N_29778);
xor UO_12 (O_12,N_29493,N_29950);
xnor UO_13 (O_13,N_29934,N_29708);
or UO_14 (O_14,N_29839,N_29783);
and UO_15 (O_15,N_29544,N_29524);
nand UO_16 (O_16,N_29797,N_29799);
or UO_17 (O_17,N_29747,N_29739);
or UO_18 (O_18,N_29712,N_29968);
or UO_19 (O_19,N_29715,N_29508);
nor UO_20 (O_20,N_29854,N_29653);
nor UO_21 (O_21,N_29609,N_29751);
or UO_22 (O_22,N_29757,N_29913);
xor UO_23 (O_23,N_29886,N_29965);
nor UO_24 (O_24,N_29690,N_29648);
nor UO_25 (O_25,N_29734,N_29849);
nor UO_26 (O_26,N_29758,N_29506);
xor UO_27 (O_27,N_29431,N_29717);
xnor UO_28 (O_28,N_29410,N_29462);
and UO_29 (O_29,N_29893,N_29752);
nor UO_30 (O_30,N_29826,N_29838);
and UO_31 (O_31,N_29564,N_29665);
and UO_32 (O_32,N_29967,N_29530);
and UO_33 (O_33,N_29697,N_29980);
nand UO_34 (O_34,N_29600,N_29859);
and UO_35 (O_35,N_29998,N_29951);
or UO_36 (O_36,N_29791,N_29488);
and UO_37 (O_37,N_29847,N_29796);
nor UO_38 (O_38,N_29436,N_29495);
nor UO_39 (O_39,N_29613,N_29721);
nor UO_40 (O_40,N_29914,N_29891);
nor UO_41 (O_41,N_29938,N_29972);
nand UO_42 (O_42,N_29479,N_29946);
and UO_43 (O_43,N_29434,N_29737);
nor UO_44 (O_44,N_29437,N_29701);
nand UO_45 (O_45,N_29947,N_29673);
xor UO_46 (O_46,N_29656,N_29776);
xnor UO_47 (O_47,N_29798,N_29457);
xor UO_48 (O_48,N_29825,N_29441);
or UO_49 (O_49,N_29860,N_29454);
nand UO_50 (O_50,N_29526,N_29408);
xnor UO_51 (O_51,N_29439,N_29513);
or UO_52 (O_52,N_29837,N_29413);
nor UO_53 (O_53,N_29470,N_29821);
nand UO_54 (O_54,N_29900,N_29409);
or UO_55 (O_55,N_29584,N_29522);
nand UO_56 (O_56,N_29562,N_29979);
xor UO_57 (O_57,N_29716,N_29892);
and UO_58 (O_58,N_29786,N_29420);
nand UO_59 (O_59,N_29639,N_29905);
xor UO_60 (O_60,N_29561,N_29875);
and UO_61 (O_61,N_29977,N_29558);
xor UO_62 (O_62,N_29908,N_29925);
nor UO_63 (O_63,N_29632,N_29615);
or UO_64 (O_64,N_29674,N_29517);
nor UO_65 (O_65,N_29961,N_29761);
and UO_66 (O_66,N_29498,N_29624);
nand UO_67 (O_67,N_29813,N_29582);
xor UO_68 (O_68,N_29952,N_29451);
nor UO_69 (O_69,N_29917,N_29702);
and UO_70 (O_70,N_29749,N_29919);
xor UO_71 (O_71,N_29617,N_29733);
or UO_72 (O_72,N_29545,N_29993);
or UO_73 (O_73,N_29475,N_29842);
nand UO_74 (O_74,N_29438,N_29635);
and UO_75 (O_75,N_29548,N_29452);
and UO_76 (O_76,N_29810,N_29966);
xor UO_77 (O_77,N_29627,N_29910);
xor UO_78 (O_78,N_29537,N_29732);
nor UO_79 (O_79,N_29652,N_29792);
nand UO_80 (O_80,N_29446,N_29646);
nor UO_81 (O_81,N_29929,N_29450);
nor UO_82 (O_82,N_29692,N_29724);
nand UO_83 (O_83,N_29480,N_29589);
xor UO_84 (O_84,N_29577,N_29597);
or UO_85 (O_85,N_29501,N_29466);
nand UO_86 (O_86,N_29667,N_29845);
or UO_87 (O_87,N_29411,N_29988);
or UO_88 (O_88,N_29963,N_29707);
xor UO_89 (O_89,N_29868,N_29720);
or UO_90 (O_90,N_29658,N_29606);
and UO_91 (O_91,N_29889,N_29858);
xor UO_92 (O_92,N_29736,N_29766);
and UO_93 (O_93,N_29552,N_29429);
nor UO_94 (O_94,N_29874,N_29704);
and UO_95 (O_95,N_29848,N_29992);
and UO_96 (O_96,N_29478,N_29865);
nor UO_97 (O_97,N_29557,N_29578);
and UO_98 (O_98,N_29922,N_29897);
nor UO_99 (O_99,N_29953,N_29873);
nor UO_100 (O_100,N_29541,N_29996);
nor UO_101 (O_101,N_29430,N_29805);
xnor UO_102 (O_102,N_29985,N_29533);
nor UO_103 (O_103,N_29764,N_29811);
nand UO_104 (O_104,N_29753,N_29406);
xor UO_105 (O_105,N_29756,N_29928);
nor UO_106 (O_106,N_29964,N_29962);
and UO_107 (O_107,N_29465,N_29402);
xnor UO_108 (O_108,N_29554,N_29689);
xor UO_109 (O_109,N_29591,N_29602);
nand UO_110 (O_110,N_29727,N_29955);
nor UO_111 (O_111,N_29435,N_29876);
nor UO_112 (O_112,N_29871,N_29754);
xor UO_113 (O_113,N_29836,N_29691);
xor UO_114 (O_114,N_29417,N_29772);
nor UO_115 (O_115,N_29536,N_29990);
or UO_116 (O_116,N_29573,N_29668);
nand UO_117 (O_117,N_29447,N_29566);
and UO_118 (O_118,N_29949,N_29956);
nand UO_119 (O_119,N_29592,N_29618);
xor UO_120 (O_120,N_29790,N_29612);
and UO_121 (O_121,N_29781,N_29676);
xor UO_122 (O_122,N_29850,N_29647);
nand UO_123 (O_123,N_29696,N_29999);
or UO_124 (O_124,N_29984,N_29585);
nor UO_125 (O_125,N_29802,N_29607);
and UO_126 (O_126,N_29631,N_29546);
nor UO_127 (O_127,N_29835,N_29924);
and UO_128 (O_128,N_29569,N_29782);
xor UO_129 (O_129,N_29789,N_29504);
nor UO_130 (O_130,N_29649,N_29971);
and UO_131 (O_131,N_29487,N_29630);
or UO_132 (O_132,N_29890,N_29492);
and UO_133 (O_133,N_29532,N_29902);
and UO_134 (O_134,N_29746,N_29540);
nor UO_135 (O_135,N_29510,N_29939);
and UO_136 (O_136,N_29471,N_29832);
xor UO_137 (O_137,N_29567,N_29975);
nor UO_138 (O_138,N_29844,N_29903);
and UO_139 (O_139,N_29440,N_29907);
or UO_140 (O_140,N_29943,N_29455);
xnor UO_141 (O_141,N_29449,N_29974);
nor UO_142 (O_142,N_29531,N_29534);
nor UO_143 (O_143,N_29755,N_29490);
nand UO_144 (O_144,N_29678,N_29515);
xnor UO_145 (O_145,N_29426,N_29700);
or UO_146 (O_146,N_29401,N_29834);
or UO_147 (O_147,N_29978,N_29959);
or UO_148 (O_148,N_29500,N_29863);
and UO_149 (O_149,N_29958,N_29738);
nand UO_150 (O_150,N_29941,N_29525);
nand UO_151 (O_151,N_29853,N_29888);
nor UO_152 (O_152,N_29725,N_29477);
and UO_153 (O_153,N_29706,N_29693);
and UO_154 (O_154,N_29827,N_29444);
nand UO_155 (O_155,N_29773,N_29620);
nor UO_156 (O_156,N_29870,N_29458);
or UO_157 (O_157,N_29636,N_29882);
and UO_158 (O_158,N_29872,N_29726);
nand UO_159 (O_159,N_29759,N_29456);
or UO_160 (O_160,N_29740,N_29468);
and UO_161 (O_161,N_29867,N_29601);
nand UO_162 (O_162,N_29660,N_29414);
or UO_163 (O_163,N_29857,N_29877);
nor UO_164 (O_164,N_29745,N_29634);
or UO_165 (O_165,N_29830,N_29671);
or UO_166 (O_166,N_29523,N_29407);
or UO_167 (O_167,N_29586,N_29555);
or UO_168 (O_168,N_29944,N_29485);
and UO_169 (O_169,N_29574,N_29625);
nor UO_170 (O_170,N_29547,N_29695);
xor UO_171 (O_171,N_29957,N_29828);
xnor UO_172 (O_172,N_29991,N_29419);
or UO_173 (O_173,N_29841,N_29682);
nor UO_174 (O_174,N_29484,N_29663);
or UO_175 (O_175,N_29785,N_29427);
nand UO_176 (O_176,N_29741,N_29464);
xor UO_177 (O_177,N_29556,N_29423);
nand UO_178 (O_178,N_29769,N_29800);
nor UO_179 (O_179,N_29594,N_29655);
nand UO_180 (O_180,N_29529,N_29819);
or UO_181 (O_181,N_29509,N_29670);
nand UO_182 (O_182,N_29405,N_29666);
nand UO_183 (O_183,N_29499,N_29816);
and UO_184 (O_184,N_29428,N_29611);
and UO_185 (O_185,N_29549,N_29774);
nand UO_186 (O_186,N_29714,N_29920);
xnor UO_187 (O_187,N_29633,N_29997);
or UO_188 (O_188,N_29491,N_29878);
nand UO_189 (O_189,N_29516,N_29614);
nor UO_190 (O_190,N_29421,N_29425);
xor UO_191 (O_191,N_29559,N_29502);
or UO_192 (O_192,N_29852,N_29942);
nand UO_193 (O_193,N_29935,N_29608);
nor UO_194 (O_194,N_29553,N_29918);
nor UO_195 (O_195,N_29823,N_29629);
nand UO_196 (O_196,N_29855,N_29527);
nand UO_197 (O_197,N_29762,N_29822);
or UO_198 (O_198,N_29467,N_29543);
nor UO_199 (O_199,N_29723,N_29448);
nand UO_200 (O_200,N_29960,N_29519);
nand UO_201 (O_201,N_29815,N_29936);
and UO_202 (O_202,N_29787,N_29424);
nor UO_203 (O_203,N_29469,N_29794);
nand UO_204 (O_204,N_29539,N_29807);
or UO_205 (O_205,N_29596,N_29846);
or UO_206 (O_206,N_29669,N_29560);
nor UO_207 (O_207,N_29699,N_29775);
or UO_208 (O_208,N_29901,N_29587);
xor UO_209 (O_209,N_29954,N_29932);
and UO_210 (O_210,N_29626,N_29461);
xnor UO_211 (O_211,N_29705,N_29583);
or UO_212 (O_212,N_29679,N_29915);
nand UO_213 (O_213,N_29731,N_29687);
xor UO_214 (O_214,N_29684,N_29497);
nand UO_215 (O_215,N_29433,N_29898);
and UO_216 (O_216,N_29686,N_29442);
and UO_217 (O_217,N_29623,N_29538);
xor UO_218 (O_218,N_29703,N_29661);
xnor UO_219 (O_219,N_29463,N_29896);
nor UO_220 (O_220,N_29881,N_29760);
nor UO_221 (O_221,N_29514,N_29982);
xor UO_222 (O_222,N_29474,N_29829);
and UO_223 (O_223,N_29482,N_29416);
xnor UO_224 (O_224,N_29415,N_29808);
or UO_225 (O_225,N_29637,N_29568);
or UO_226 (O_226,N_29742,N_29472);
nand UO_227 (O_227,N_29987,N_29899);
nand UO_228 (O_228,N_29793,N_29595);
and UO_229 (O_229,N_29521,N_29765);
xnor UO_230 (O_230,N_29418,N_29535);
and UO_231 (O_231,N_29486,N_29880);
or UO_232 (O_232,N_29659,N_29843);
nand UO_233 (O_233,N_29443,N_29770);
nor UO_234 (O_234,N_29912,N_29662);
or UO_235 (O_235,N_29598,N_29983);
xnor UO_236 (O_236,N_29869,N_29883);
and UO_237 (O_237,N_29453,N_29820);
and UO_238 (O_238,N_29489,N_29518);
nor UO_239 (O_239,N_29672,N_29812);
and UO_240 (O_240,N_29563,N_29735);
nand UO_241 (O_241,N_29763,N_29603);
and UO_242 (O_242,N_29719,N_29483);
nand UO_243 (O_243,N_29507,N_29809);
nor UO_244 (O_244,N_29989,N_29904);
nand UO_245 (O_245,N_29744,N_29570);
nand UO_246 (O_246,N_29650,N_29604);
xnor UO_247 (O_247,N_29511,N_29654);
or UO_248 (O_248,N_29851,N_29579);
or UO_249 (O_249,N_29885,N_29750);
nand UO_250 (O_250,N_29494,N_29640);
xnor UO_251 (O_251,N_29937,N_29923);
xnor UO_252 (O_252,N_29748,N_29412);
nand UO_253 (O_253,N_29404,N_29767);
or UO_254 (O_254,N_29476,N_29806);
nor UO_255 (O_255,N_29856,N_29581);
nand UO_256 (O_256,N_29638,N_29804);
and UO_257 (O_257,N_29722,N_29565);
and UO_258 (O_258,N_29718,N_29680);
and UO_259 (O_259,N_29862,N_29473);
nand UO_260 (O_260,N_29916,N_29709);
and UO_261 (O_261,N_29571,N_29895);
and UO_262 (O_262,N_29619,N_29520);
and UO_263 (O_263,N_29400,N_29711);
nor UO_264 (O_264,N_29909,N_29933);
nand UO_265 (O_265,N_29879,N_29921);
nor UO_266 (O_266,N_29610,N_29986);
nand UO_267 (O_267,N_29593,N_29729);
or UO_268 (O_268,N_29930,N_29432);
xnor UO_269 (O_269,N_29675,N_29864);
xor UO_270 (O_270,N_29459,N_29803);
nand UO_271 (O_271,N_29777,N_29683);
nor UO_272 (O_272,N_29771,N_29866);
and UO_273 (O_273,N_29681,N_29621);
nand UO_274 (O_274,N_29445,N_29481);
and UO_275 (O_275,N_29995,N_29768);
nor UO_276 (O_276,N_29616,N_29580);
nor UO_277 (O_277,N_29906,N_29884);
nand UO_278 (O_278,N_29831,N_29927);
xnor UO_279 (O_279,N_29840,N_29795);
nor UO_280 (O_280,N_29940,N_29664);
xor UO_281 (O_281,N_29628,N_29976);
nor UO_282 (O_282,N_29948,N_29926);
nand UO_283 (O_283,N_29814,N_29643);
nor UO_284 (O_284,N_29641,N_29713);
xnor UO_285 (O_285,N_29590,N_29730);
xor UO_286 (O_286,N_29710,N_29677);
xor UO_287 (O_287,N_29780,N_29994);
xnor UO_288 (O_288,N_29931,N_29894);
nor UO_289 (O_289,N_29743,N_29588);
nor UO_290 (O_290,N_29833,N_29403);
nor UO_291 (O_291,N_29512,N_29779);
or UO_292 (O_292,N_29911,N_29969);
xor UO_293 (O_293,N_29460,N_29728);
nand UO_294 (O_294,N_29973,N_29651);
nand UO_295 (O_295,N_29576,N_29575);
and UO_296 (O_296,N_29685,N_29698);
nand UO_297 (O_297,N_29505,N_29645);
xor UO_298 (O_298,N_29788,N_29551);
or UO_299 (O_299,N_29605,N_29981);
and UO_300 (O_300,N_29437,N_29904);
xor UO_301 (O_301,N_29639,N_29462);
or UO_302 (O_302,N_29911,N_29602);
nand UO_303 (O_303,N_29491,N_29954);
xnor UO_304 (O_304,N_29817,N_29987);
and UO_305 (O_305,N_29752,N_29750);
and UO_306 (O_306,N_29911,N_29565);
nor UO_307 (O_307,N_29918,N_29606);
nor UO_308 (O_308,N_29409,N_29803);
or UO_309 (O_309,N_29659,N_29967);
nor UO_310 (O_310,N_29833,N_29531);
nand UO_311 (O_311,N_29406,N_29998);
xor UO_312 (O_312,N_29708,N_29571);
xor UO_313 (O_313,N_29762,N_29434);
xnor UO_314 (O_314,N_29540,N_29724);
xnor UO_315 (O_315,N_29527,N_29504);
nor UO_316 (O_316,N_29789,N_29577);
or UO_317 (O_317,N_29639,N_29640);
and UO_318 (O_318,N_29896,N_29558);
or UO_319 (O_319,N_29559,N_29596);
xor UO_320 (O_320,N_29677,N_29665);
and UO_321 (O_321,N_29564,N_29421);
nand UO_322 (O_322,N_29446,N_29400);
and UO_323 (O_323,N_29975,N_29610);
xnor UO_324 (O_324,N_29512,N_29430);
nor UO_325 (O_325,N_29772,N_29735);
or UO_326 (O_326,N_29895,N_29440);
or UO_327 (O_327,N_29764,N_29415);
nor UO_328 (O_328,N_29657,N_29895);
and UO_329 (O_329,N_29658,N_29429);
or UO_330 (O_330,N_29586,N_29403);
nor UO_331 (O_331,N_29647,N_29519);
xnor UO_332 (O_332,N_29916,N_29789);
nand UO_333 (O_333,N_29531,N_29841);
nand UO_334 (O_334,N_29546,N_29872);
nor UO_335 (O_335,N_29477,N_29625);
nand UO_336 (O_336,N_29584,N_29487);
nand UO_337 (O_337,N_29529,N_29453);
xnor UO_338 (O_338,N_29876,N_29492);
xnor UO_339 (O_339,N_29899,N_29521);
or UO_340 (O_340,N_29720,N_29494);
nor UO_341 (O_341,N_29445,N_29468);
nor UO_342 (O_342,N_29553,N_29472);
nand UO_343 (O_343,N_29813,N_29783);
or UO_344 (O_344,N_29523,N_29843);
nand UO_345 (O_345,N_29641,N_29510);
xnor UO_346 (O_346,N_29743,N_29801);
and UO_347 (O_347,N_29745,N_29515);
and UO_348 (O_348,N_29952,N_29574);
xnor UO_349 (O_349,N_29712,N_29773);
xor UO_350 (O_350,N_29608,N_29788);
or UO_351 (O_351,N_29996,N_29597);
or UO_352 (O_352,N_29445,N_29458);
and UO_353 (O_353,N_29639,N_29768);
nor UO_354 (O_354,N_29950,N_29687);
xor UO_355 (O_355,N_29617,N_29574);
nand UO_356 (O_356,N_29986,N_29646);
xor UO_357 (O_357,N_29816,N_29711);
and UO_358 (O_358,N_29843,N_29468);
and UO_359 (O_359,N_29646,N_29771);
xor UO_360 (O_360,N_29936,N_29425);
nor UO_361 (O_361,N_29875,N_29723);
or UO_362 (O_362,N_29541,N_29506);
nor UO_363 (O_363,N_29530,N_29439);
xnor UO_364 (O_364,N_29413,N_29602);
or UO_365 (O_365,N_29729,N_29878);
nand UO_366 (O_366,N_29974,N_29492);
and UO_367 (O_367,N_29484,N_29963);
xnor UO_368 (O_368,N_29483,N_29891);
xor UO_369 (O_369,N_29913,N_29427);
nor UO_370 (O_370,N_29884,N_29730);
and UO_371 (O_371,N_29915,N_29467);
and UO_372 (O_372,N_29672,N_29741);
nor UO_373 (O_373,N_29584,N_29533);
nor UO_374 (O_374,N_29701,N_29624);
and UO_375 (O_375,N_29465,N_29882);
and UO_376 (O_376,N_29465,N_29441);
nor UO_377 (O_377,N_29867,N_29480);
xor UO_378 (O_378,N_29664,N_29937);
or UO_379 (O_379,N_29959,N_29708);
xor UO_380 (O_380,N_29470,N_29563);
nand UO_381 (O_381,N_29976,N_29433);
xnor UO_382 (O_382,N_29978,N_29802);
nor UO_383 (O_383,N_29842,N_29457);
and UO_384 (O_384,N_29718,N_29940);
and UO_385 (O_385,N_29680,N_29825);
nand UO_386 (O_386,N_29704,N_29473);
nor UO_387 (O_387,N_29495,N_29716);
nand UO_388 (O_388,N_29767,N_29879);
nand UO_389 (O_389,N_29649,N_29431);
nand UO_390 (O_390,N_29847,N_29949);
xnor UO_391 (O_391,N_29647,N_29521);
xor UO_392 (O_392,N_29717,N_29423);
nor UO_393 (O_393,N_29651,N_29700);
or UO_394 (O_394,N_29786,N_29858);
and UO_395 (O_395,N_29416,N_29804);
or UO_396 (O_396,N_29627,N_29552);
or UO_397 (O_397,N_29617,N_29720);
or UO_398 (O_398,N_29492,N_29649);
or UO_399 (O_399,N_29533,N_29862);
nor UO_400 (O_400,N_29849,N_29945);
nor UO_401 (O_401,N_29658,N_29760);
or UO_402 (O_402,N_29435,N_29505);
and UO_403 (O_403,N_29903,N_29636);
nor UO_404 (O_404,N_29707,N_29438);
nor UO_405 (O_405,N_29485,N_29599);
nor UO_406 (O_406,N_29514,N_29666);
xnor UO_407 (O_407,N_29461,N_29654);
and UO_408 (O_408,N_29440,N_29629);
xnor UO_409 (O_409,N_29717,N_29883);
or UO_410 (O_410,N_29989,N_29931);
xor UO_411 (O_411,N_29988,N_29538);
xor UO_412 (O_412,N_29795,N_29704);
xor UO_413 (O_413,N_29946,N_29605);
and UO_414 (O_414,N_29675,N_29549);
xor UO_415 (O_415,N_29741,N_29632);
xnor UO_416 (O_416,N_29700,N_29593);
nand UO_417 (O_417,N_29921,N_29564);
nand UO_418 (O_418,N_29738,N_29583);
nand UO_419 (O_419,N_29727,N_29880);
nand UO_420 (O_420,N_29768,N_29428);
nand UO_421 (O_421,N_29420,N_29976);
and UO_422 (O_422,N_29659,N_29724);
nor UO_423 (O_423,N_29669,N_29466);
nand UO_424 (O_424,N_29400,N_29747);
nand UO_425 (O_425,N_29592,N_29848);
nor UO_426 (O_426,N_29448,N_29470);
and UO_427 (O_427,N_29473,N_29493);
xnor UO_428 (O_428,N_29692,N_29454);
xor UO_429 (O_429,N_29921,N_29527);
or UO_430 (O_430,N_29481,N_29497);
nand UO_431 (O_431,N_29665,N_29545);
xor UO_432 (O_432,N_29548,N_29584);
xor UO_433 (O_433,N_29507,N_29676);
and UO_434 (O_434,N_29541,N_29932);
xnor UO_435 (O_435,N_29620,N_29829);
nor UO_436 (O_436,N_29747,N_29402);
and UO_437 (O_437,N_29430,N_29899);
or UO_438 (O_438,N_29970,N_29989);
xnor UO_439 (O_439,N_29614,N_29473);
or UO_440 (O_440,N_29510,N_29970);
or UO_441 (O_441,N_29419,N_29898);
or UO_442 (O_442,N_29984,N_29616);
or UO_443 (O_443,N_29743,N_29607);
and UO_444 (O_444,N_29581,N_29956);
or UO_445 (O_445,N_29761,N_29964);
nor UO_446 (O_446,N_29877,N_29880);
nor UO_447 (O_447,N_29605,N_29501);
and UO_448 (O_448,N_29987,N_29723);
xor UO_449 (O_449,N_29808,N_29549);
nand UO_450 (O_450,N_29500,N_29966);
xor UO_451 (O_451,N_29756,N_29868);
nor UO_452 (O_452,N_29974,N_29415);
or UO_453 (O_453,N_29471,N_29770);
or UO_454 (O_454,N_29824,N_29755);
nand UO_455 (O_455,N_29413,N_29659);
and UO_456 (O_456,N_29524,N_29676);
nor UO_457 (O_457,N_29668,N_29998);
nand UO_458 (O_458,N_29612,N_29530);
and UO_459 (O_459,N_29891,N_29624);
xnor UO_460 (O_460,N_29690,N_29990);
and UO_461 (O_461,N_29850,N_29659);
nor UO_462 (O_462,N_29683,N_29631);
nand UO_463 (O_463,N_29676,N_29494);
or UO_464 (O_464,N_29500,N_29693);
or UO_465 (O_465,N_29858,N_29807);
nor UO_466 (O_466,N_29494,N_29760);
nand UO_467 (O_467,N_29464,N_29989);
xor UO_468 (O_468,N_29559,N_29532);
and UO_469 (O_469,N_29884,N_29969);
xnor UO_470 (O_470,N_29795,N_29782);
nand UO_471 (O_471,N_29431,N_29682);
or UO_472 (O_472,N_29853,N_29679);
nor UO_473 (O_473,N_29451,N_29957);
xor UO_474 (O_474,N_29860,N_29872);
nand UO_475 (O_475,N_29930,N_29866);
nor UO_476 (O_476,N_29592,N_29803);
xor UO_477 (O_477,N_29621,N_29550);
nor UO_478 (O_478,N_29712,N_29861);
xor UO_479 (O_479,N_29731,N_29946);
xnor UO_480 (O_480,N_29561,N_29884);
or UO_481 (O_481,N_29832,N_29785);
nor UO_482 (O_482,N_29660,N_29521);
and UO_483 (O_483,N_29658,N_29739);
nand UO_484 (O_484,N_29699,N_29835);
nor UO_485 (O_485,N_29481,N_29521);
xnor UO_486 (O_486,N_29812,N_29444);
and UO_487 (O_487,N_29761,N_29735);
xnor UO_488 (O_488,N_29627,N_29701);
xor UO_489 (O_489,N_29662,N_29728);
and UO_490 (O_490,N_29873,N_29621);
nand UO_491 (O_491,N_29945,N_29769);
or UO_492 (O_492,N_29734,N_29542);
nor UO_493 (O_493,N_29474,N_29740);
nand UO_494 (O_494,N_29624,N_29993);
or UO_495 (O_495,N_29676,N_29951);
or UO_496 (O_496,N_29428,N_29690);
nor UO_497 (O_497,N_29973,N_29708);
nor UO_498 (O_498,N_29771,N_29527);
nand UO_499 (O_499,N_29877,N_29813);
xnor UO_500 (O_500,N_29586,N_29762);
and UO_501 (O_501,N_29421,N_29615);
or UO_502 (O_502,N_29919,N_29802);
and UO_503 (O_503,N_29876,N_29659);
nand UO_504 (O_504,N_29777,N_29953);
and UO_505 (O_505,N_29482,N_29892);
and UO_506 (O_506,N_29635,N_29744);
and UO_507 (O_507,N_29749,N_29665);
nor UO_508 (O_508,N_29620,N_29862);
nand UO_509 (O_509,N_29531,N_29887);
or UO_510 (O_510,N_29461,N_29458);
or UO_511 (O_511,N_29712,N_29572);
xor UO_512 (O_512,N_29523,N_29926);
nand UO_513 (O_513,N_29549,N_29932);
and UO_514 (O_514,N_29438,N_29583);
xnor UO_515 (O_515,N_29588,N_29786);
nor UO_516 (O_516,N_29896,N_29856);
nor UO_517 (O_517,N_29828,N_29843);
and UO_518 (O_518,N_29425,N_29676);
nor UO_519 (O_519,N_29600,N_29459);
xnor UO_520 (O_520,N_29935,N_29789);
and UO_521 (O_521,N_29456,N_29846);
nand UO_522 (O_522,N_29468,N_29934);
nor UO_523 (O_523,N_29875,N_29953);
nor UO_524 (O_524,N_29926,N_29853);
nand UO_525 (O_525,N_29504,N_29744);
xnor UO_526 (O_526,N_29564,N_29892);
nand UO_527 (O_527,N_29904,N_29724);
and UO_528 (O_528,N_29469,N_29428);
or UO_529 (O_529,N_29651,N_29809);
or UO_530 (O_530,N_29541,N_29632);
and UO_531 (O_531,N_29719,N_29584);
xor UO_532 (O_532,N_29680,N_29421);
or UO_533 (O_533,N_29521,N_29419);
and UO_534 (O_534,N_29774,N_29824);
nand UO_535 (O_535,N_29471,N_29677);
or UO_536 (O_536,N_29812,N_29665);
xor UO_537 (O_537,N_29917,N_29772);
xnor UO_538 (O_538,N_29461,N_29723);
nand UO_539 (O_539,N_29630,N_29628);
xor UO_540 (O_540,N_29508,N_29520);
nand UO_541 (O_541,N_29880,N_29573);
xnor UO_542 (O_542,N_29655,N_29490);
and UO_543 (O_543,N_29440,N_29692);
or UO_544 (O_544,N_29855,N_29970);
or UO_545 (O_545,N_29991,N_29454);
nor UO_546 (O_546,N_29933,N_29808);
or UO_547 (O_547,N_29602,N_29800);
and UO_548 (O_548,N_29537,N_29776);
and UO_549 (O_549,N_29607,N_29440);
nor UO_550 (O_550,N_29601,N_29855);
or UO_551 (O_551,N_29477,N_29865);
nand UO_552 (O_552,N_29564,N_29605);
or UO_553 (O_553,N_29738,N_29585);
nor UO_554 (O_554,N_29449,N_29577);
nand UO_555 (O_555,N_29926,N_29433);
xnor UO_556 (O_556,N_29718,N_29485);
or UO_557 (O_557,N_29845,N_29506);
and UO_558 (O_558,N_29508,N_29996);
and UO_559 (O_559,N_29933,N_29727);
and UO_560 (O_560,N_29833,N_29675);
nand UO_561 (O_561,N_29535,N_29547);
nand UO_562 (O_562,N_29415,N_29428);
or UO_563 (O_563,N_29850,N_29544);
and UO_564 (O_564,N_29457,N_29830);
nor UO_565 (O_565,N_29659,N_29679);
xor UO_566 (O_566,N_29675,N_29679);
and UO_567 (O_567,N_29908,N_29475);
xnor UO_568 (O_568,N_29561,N_29809);
or UO_569 (O_569,N_29544,N_29939);
nor UO_570 (O_570,N_29729,N_29862);
and UO_571 (O_571,N_29421,N_29520);
and UO_572 (O_572,N_29904,N_29498);
xor UO_573 (O_573,N_29843,N_29707);
and UO_574 (O_574,N_29733,N_29867);
xnor UO_575 (O_575,N_29708,N_29437);
or UO_576 (O_576,N_29603,N_29486);
xnor UO_577 (O_577,N_29668,N_29751);
nor UO_578 (O_578,N_29503,N_29925);
and UO_579 (O_579,N_29846,N_29992);
nand UO_580 (O_580,N_29991,N_29705);
and UO_581 (O_581,N_29939,N_29403);
nor UO_582 (O_582,N_29711,N_29485);
nand UO_583 (O_583,N_29569,N_29799);
xor UO_584 (O_584,N_29468,N_29511);
or UO_585 (O_585,N_29763,N_29672);
nand UO_586 (O_586,N_29450,N_29441);
or UO_587 (O_587,N_29528,N_29662);
nor UO_588 (O_588,N_29919,N_29456);
or UO_589 (O_589,N_29758,N_29803);
nand UO_590 (O_590,N_29984,N_29400);
or UO_591 (O_591,N_29942,N_29712);
and UO_592 (O_592,N_29897,N_29747);
or UO_593 (O_593,N_29446,N_29637);
nor UO_594 (O_594,N_29605,N_29884);
or UO_595 (O_595,N_29946,N_29424);
nand UO_596 (O_596,N_29873,N_29473);
or UO_597 (O_597,N_29455,N_29873);
or UO_598 (O_598,N_29412,N_29954);
nor UO_599 (O_599,N_29599,N_29724);
or UO_600 (O_600,N_29683,N_29904);
nor UO_601 (O_601,N_29932,N_29590);
xnor UO_602 (O_602,N_29779,N_29548);
nor UO_603 (O_603,N_29750,N_29532);
or UO_604 (O_604,N_29823,N_29884);
xor UO_605 (O_605,N_29544,N_29818);
xnor UO_606 (O_606,N_29866,N_29415);
nand UO_607 (O_607,N_29634,N_29961);
xnor UO_608 (O_608,N_29583,N_29482);
or UO_609 (O_609,N_29481,N_29413);
or UO_610 (O_610,N_29923,N_29568);
and UO_611 (O_611,N_29811,N_29903);
xnor UO_612 (O_612,N_29722,N_29977);
or UO_613 (O_613,N_29654,N_29666);
xor UO_614 (O_614,N_29616,N_29600);
nor UO_615 (O_615,N_29909,N_29954);
nand UO_616 (O_616,N_29872,N_29908);
xor UO_617 (O_617,N_29811,N_29562);
and UO_618 (O_618,N_29490,N_29920);
xor UO_619 (O_619,N_29847,N_29751);
xor UO_620 (O_620,N_29816,N_29726);
or UO_621 (O_621,N_29978,N_29717);
xor UO_622 (O_622,N_29643,N_29712);
nor UO_623 (O_623,N_29545,N_29927);
nand UO_624 (O_624,N_29784,N_29660);
nand UO_625 (O_625,N_29645,N_29655);
nor UO_626 (O_626,N_29455,N_29888);
xnor UO_627 (O_627,N_29508,N_29918);
xnor UO_628 (O_628,N_29413,N_29782);
nand UO_629 (O_629,N_29938,N_29487);
and UO_630 (O_630,N_29848,N_29724);
or UO_631 (O_631,N_29557,N_29442);
nor UO_632 (O_632,N_29492,N_29528);
nor UO_633 (O_633,N_29852,N_29780);
xnor UO_634 (O_634,N_29751,N_29840);
or UO_635 (O_635,N_29817,N_29634);
xnor UO_636 (O_636,N_29990,N_29915);
nand UO_637 (O_637,N_29813,N_29663);
nor UO_638 (O_638,N_29851,N_29595);
and UO_639 (O_639,N_29644,N_29501);
and UO_640 (O_640,N_29609,N_29607);
and UO_641 (O_641,N_29671,N_29587);
nand UO_642 (O_642,N_29937,N_29656);
xor UO_643 (O_643,N_29628,N_29448);
and UO_644 (O_644,N_29759,N_29889);
or UO_645 (O_645,N_29657,N_29514);
nand UO_646 (O_646,N_29915,N_29852);
or UO_647 (O_647,N_29760,N_29485);
xnor UO_648 (O_648,N_29831,N_29825);
xnor UO_649 (O_649,N_29857,N_29902);
and UO_650 (O_650,N_29407,N_29817);
nand UO_651 (O_651,N_29661,N_29925);
nand UO_652 (O_652,N_29464,N_29938);
nor UO_653 (O_653,N_29987,N_29461);
or UO_654 (O_654,N_29535,N_29768);
xnor UO_655 (O_655,N_29843,N_29801);
or UO_656 (O_656,N_29545,N_29797);
nor UO_657 (O_657,N_29916,N_29403);
or UO_658 (O_658,N_29943,N_29672);
nor UO_659 (O_659,N_29517,N_29721);
nor UO_660 (O_660,N_29438,N_29936);
nor UO_661 (O_661,N_29726,N_29746);
xor UO_662 (O_662,N_29603,N_29443);
xnor UO_663 (O_663,N_29494,N_29604);
and UO_664 (O_664,N_29595,N_29554);
and UO_665 (O_665,N_29588,N_29485);
and UO_666 (O_666,N_29445,N_29400);
nor UO_667 (O_667,N_29955,N_29496);
or UO_668 (O_668,N_29889,N_29755);
xnor UO_669 (O_669,N_29651,N_29951);
or UO_670 (O_670,N_29401,N_29550);
or UO_671 (O_671,N_29948,N_29402);
or UO_672 (O_672,N_29668,N_29515);
or UO_673 (O_673,N_29671,N_29701);
nor UO_674 (O_674,N_29985,N_29683);
xor UO_675 (O_675,N_29827,N_29784);
nand UO_676 (O_676,N_29446,N_29403);
xor UO_677 (O_677,N_29413,N_29681);
or UO_678 (O_678,N_29673,N_29631);
xnor UO_679 (O_679,N_29786,N_29874);
nor UO_680 (O_680,N_29996,N_29653);
nor UO_681 (O_681,N_29516,N_29436);
xnor UO_682 (O_682,N_29774,N_29485);
nand UO_683 (O_683,N_29746,N_29411);
xor UO_684 (O_684,N_29817,N_29471);
nand UO_685 (O_685,N_29413,N_29550);
xor UO_686 (O_686,N_29769,N_29496);
or UO_687 (O_687,N_29929,N_29607);
and UO_688 (O_688,N_29859,N_29997);
and UO_689 (O_689,N_29859,N_29979);
and UO_690 (O_690,N_29627,N_29959);
nand UO_691 (O_691,N_29684,N_29851);
or UO_692 (O_692,N_29648,N_29874);
xor UO_693 (O_693,N_29926,N_29439);
nor UO_694 (O_694,N_29709,N_29908);
and UO_695 (O_695,N_29904,N_29715);
and UO_696 (O_696,N_29924,N_29971);
and UO_697 (O_697,N_29412,N_29633);
xor UO_698 (O_698,N_29925,N_29775);
and UO_699 (O_699,N_29401,N_29645);
and UO_700 (O_700,N_29401,N_29455);
xor UO_701 (O_701,N_29609,N_29473);
and UO_702 (O_702,N_29456,N_29469);
nor UO_703 (O_703,N_29546,N_29968);
and UO_704 (O_704,N_29736,N_29818);
nand UO_705 (O_705,N_29471,N_29933);
xnor UO_706 (O_706,N_29423,N_29680);
and UO_707 (O_707,N_29990,N_29940);
nor UO_708 (O_708,N_29519,N_29716);
and UO_709 (O_709,N_29842,N_29681);
xnor UO_710 (O_710,N_29509,N_29908);
xnor UO_711 (O_711,N_29893,N_29414);
or UO_712 (O_712,N_29464,N_29848);
nor UO_713 (O_713,N_29608,N_29454);
or UO_714 (O_714,N_29481,N_29564);
and UO_715 (O_715,N_29723,N_29762);
xnor UO_716 (O_716,N_29551,N_29408);
or UO_717 (O_717,N_29766,N_29610);
nor UO_718 (O_718,N_29627,N_29535);
nor UO_719 (O_719,N_29415,N_29712);
and UO_720 (O_720,N_29547,N_29775);
and UO_721 (O_721,N_29979,N_29469);
nand UO_722 (O_722,N_29739,N_29504);
and UO_723 (O_723,N_29759,N_29949);
xnor UO_724 (O_724,N_29869,N_29763);
xnor UO_725 (O_725,N_29464,N_29431);
or UO_726 (O_726,N_29921,N_29415);
or UO_727 (O_727,N_29670,N_29640);
nor UO_728 (O_728,N_29601,N_29995);
nand UO_729 (O_729,N_29864,N_29947);
xnor UO_730 (O_730,N_29611,N_29995);
xnor UO_731 (O_731,N_29438,N_29996);
nor UO_732 (O_732,N_29708,N_29562);
xnor UO_733 (O_733,N_29567,N_29889);
or UO_734 (O_734,N_29404,N_29492);
or UO_735 (O_735,N_29795,N_29564);
and UO_736 (O_736,N_29411,N_29744);
or UO_737 (O_737,N_29529,N_29950);
and UO_738 (O_738,N_29788,N_29811);
xnor UO_739 (O_739,N_29466,N_29629);
xnor UO_740 (O_740,N_29810,N_29714);
nand UO_741 (O_741,N_29787,N_29724);
xnor UO_742 (O_742,N_29950,N_29552);
xnor UO_743 (O_743,N_29492,N_29813);
xor UO_744 (O_744,N_29988,N_29799);
or UO_745 (O_745,N_29544,N_29518);
xor UO_746 (O_746,N_29858,N_29557);
nor UO_747 (O_747,N_29466,N_29610);
or UO_748 (O_748,N_29966,N_29532);
xor UO_749 (O_749,N_29625,N_29600);
or UO_750 (O_750,N_29608,N_29857);
xor UO_751 (O_751,N_29706,N_29814);
or UO_752 (O_752,N_29506,N_29448);
or UO_753 (O_753,N_29450,N_29795);
xnor UO_754 (O_754,N_29928,N_29490);
nand UO_755 (O_755,N_29853,N_29692);
nand UO_756 (O_756,N_29477,N_29914);
or UO_757 (O_757,N_29851,N_29925);
and UO_758 (O_758,N_29514,N_29677);
xor UO_759 (O_759,N_29908,N_29584);
xor UO_760 (O_760,N_29573,N_29578);
nor UO_761 (O_761,N_29974,N_29911);
nand UO_762 (O_762,N_29648,N_29997);
xnor UO_763 (O_763,N_29755,N_29964);
and UO_764 (O_764,N_29617,N_29455);
nor UO_765 (O_765,N_29754,N_29670);
nor UO_766 (O_766,N_29962,N_29845);
nand UO_767 (O_767,N_29620,N_29602);
nor UO_768 (O_768,N_29552,N_29639);
nand UO_769 (O_769,N_29860,N_29809);
or UO_770 (O_770,N_29732,N_29982);
nor UO_771 (O_771,N_29931,N_29452);
nor UO_772 (O_772,N_29649,N_29532);
xor UO_773 (O_773,N_29692,N_29433);
or UO_774 (O_774,N_29588,N_29521);
nand UO_775 (O_775,N_29631,N_29661);
xor UO_776 (O_776,N_29636,N_29877);
nand UO_777 (O_777,N_29579,N_29462);
and UO_778 (O_778,N_29425,N_29942);
nand UO_779 (O_779,N_29796,N_29707);
or UO_780 (O_780,N_29576,N_29651);
nor UO_781 (O_781,N_29752,N_29403);
and UO_782 (O_782,N_29683,N_29564);
nand UO_783 (O_783,N_29722,N_29608);
xor UO_784 (O_784,N_29549,N_29911);
nand UO_785 (O_785,N_29739,N_29862);
xnor UO_786 (O_786,N_29917,N_29599);
nand UO_787 (O_787,N_29785,N_29609);
nand UO_788 (O_788,N_29692,N_29735);
nand UO_789 (O_789,N_29889,N_29831);
nor UO_790 (O_790,N_29552,N_29881);
nor UO_791 (O_791,N_29727,N_29912);
xor UO_792 (O_792,N_29603,N_29407);
nand UO_793 (O_793,N_29961,N_29880);
nand UO_794 (O_794,N_29776,N_29706);
xnor UO_795 (O_795,N_29438,N_29956);
and UO_796 (O_796,N_29807,N_29792);
or UO_797 (O_797,N_29447,N_29870);
or UO_798 (O_798,N_29404,N_29481);
nor UO_799 (O_799,N_29968,N_29540);
xor UO_800 (O_800,N_29797,N_29596);
nand UO_801 (O_801,N_29768,N_29982);
or UO_802 (O_802,N_29592,N_29696);
xor UO_803 (O_803,N_29506,N_29842);
and UO_804 (O_804,N_29409,N_29411);
nand UO_805 (O_805,N_29669,N_29659);
nand UO_806 (O_806,N_29438,N_29458);
xnor UO_807 (O_807,N_29887,N_29753);
nand UO_808 (O_808,N_29751,N_29688);
xnor UO_809 (O_809,N_29528,N_29774);
and UO_810 (O_810,N_29711,N_29867);
nor UO_811 (O_811,N_29837,N_29851);
and UO_812 (O_812,N_29875,N_29664);
nor UO_813 (O_813,N_29447,N_29889);
xnor UO_814 (O_814,N_29731,N_29916);
or UO_815 (O_815,N_29415,N_29935);
nand UO_816 (O_816,N_29619,N_29964);
and UO_817 (O_817,N_29929,N_29977);
nand UO_818 (O_818,N_29812,N_29864);
and UO_819 (O_819,N_29811,N_29682);
nand UO_820 (O_820,N_29424,N_29613);
xnor UO_821 (O_821,N_29742,N_29540);
nand UO_822 (O_822,N_29445,N_29659);
xor UO_823 (O_823,N_29594,N_29883);
nor UO_824 (O_824,N_29525,N_29847);
and UO_825 (O_825,N_29443,N_29881);
or UO_826 (O_826,N_29757,N_29494);
nor UO_827 (O_827,N_29786,N_29738);
nor UO_828 (O_828,N_29465,N_29831);
xnor UO_829 (O_829,N_29617,N_29748);
nand UO_830 (O_830,N_29521,N_29593);
and UO_831 (O_831,N_29782,N_29615);
xor UO_832 (O_832,N_29821,N_29932);
nand UO_833 (O_833,N_29545,N_29968);
nand UO_834 (O_834,N_29859,N_29467);
nor UO_835 (O_835,N_29727,N_29562);
nor UO_836 (O_836,N_29609,N_29791);
or UO_837 (O_837,N_29615,N_29593);
nor UO_838 (O_838,N_29808,N_29806);
xor UO_839 (O_839,N_29527,N_29739);
or UO_840 (O_840,N_29502,N_29438);
xor UO_841 (O_841,N_29675,N_29496);
nand UO_842 (O_842,N_29504,N_29603);
and UO_843 (O_843,N_29984,N_29722);
xnor UO_844 (O_844,N_29803,N_29433);
nor UO_845 (O_845,N_29829,N_29564);
nor UO_846 (O_846,N_29824,N_29527);
or UO_847 (O_847,N_29532,N_29941);
nor UO_848 (O_848,N_29658,N_29473);
nor UO_849 (O_849,N_29484,N_29733);
nand UO_850 (O_850,N_29686,N_29509);
nor UO_851 (O_851,N_29939,N_29421);
nand UO_852 (O_852,N_29647,N_29644);
nand UO_853 (O_853,N_29729,N_29621);
or UO_854 (O_854,N_29782,N_29513);
nand UO_855 (O_855,N_29639,N_29786);
and UO_856 (O_856,N_29717,N_29407);
xnor UO_857 (O_857,N_29999,N_29862);
and UO_858 (O_858,N_29612,N_29414);
nand UO_859 (O_859,N_29831,N_29586);
or UO_860 (O_860,N_29857,N_29878);
xor UO_861 (O_861,N_29452,N_29543);
or UO_862 (O_862,N_29873,N_29409);
xor UO_863 (O_863,N_29400,N_29923);
nand UO_864 (O_864,N_29625,N_29617);
nor UO_865 (O_865,N_29821,N_29717);
and UO_866 (O_866,N_29632,N_29452);
and UO_867 (O_867,N_29782,N_29876);
nand UO_868 (O_868,N_29508,N_29461);
nor UO_869 (O_869,N_29674,N_29883);
nor UO_870 (O_870,N_29896,N_29508);
or UO_871 (O_871,N_29682,N_29976);
and UO_872 (O_872,N_29803,N_29745);
and UO_873 (O_873,N_29818,N_29953);
xor UO_874 (O_874,N_29906,N_29689);
and UO_875 (O_875,N_29586,N_29569);
nor UO_876 (O_876,N_29403,N_29952);
nand UO_877 (O_877,N_29480,N_29686);
nor UO_878 (O_878,N_29763,N_29585);
and UO_879 (O_879,N_29834,N_29646);
and UO_880 (O_880,N_29764,N_29827);
nand UO_881 (O_881,N_29476,N_29440);
xnor UO_882 (O_882,N_29785,N_29848);
nand UO_883 (O_883,N_29861,N_29460);
xor UO_884 (O_884,N_29946,N_29410);
and UO_885 (O_885,N_29966,N_29670);
xor UO_886 (O_886,N_29446,N_29482);
nor UO_887 (O_887,N_29592,N_29596);
and UO_888 (O_888,N_29945,N_29881);
nand UO_889 (O_889,N_29601,N_29872);
and UO_890 (O_890,N_29535,N_29417);
nor UO_891 (O_891,N_29641,N_29927);
and UO_892 (O_892,N_29917,N_29899);
nor UO_893 (O_893,N_29673,N_29982);
nand UO_894 (O_894,N_29757,N_29475);
nor UO_895 (O_895,N_29762,N_29596);
or UO_896 (O_896,N_29799,N_29582);
and UO_897 (O_897,N_29685,N_29958);
xnor UO_898 (O_898,N_29951,N_29600);
xnor UO_899 (O_899,N_29401,N_29976);
xor UO_900 (O_900,N_29949,N_29980);
nand UO_901 (O_901,N_29881,N_29883);
and UO_902 (O_902,N_29789,N_29888);
or UO_903 (O_903,N_29847,N_29634);
nor UO_904 (O_904,N_29814,N_29560);
or UO_905 (O_905,N_29847,N_29833);
nor UO_906 (O_906,N_29749,N_29592);
nor UO_907 (O_907,N_29952,N_29790);
xor UO_908 (O_908,N_29634,N_29741);
nand UO_909 (O_909,N_29738,N_29829);
or UO_910 (O_910,N_29482,N_29807);
nand UO_911 (O_911,N_29937,N_29864);
or UO_912 (O_912,N_29541,N_29564);
nor UO_913 (O_913,N_29457,N_29969);
or UO_914 (O_914,N_29853,N_29729);
nor UO_915 (O_915,N_29456,N_29569);
and UO_916 (O_916,N_29625,N_29652);
nor UO_917 (O_917,N_29721,N_29535);
nand UO_918 (O_918,N_29615,N_29751);
nand UO_919 (O_919,N_29923,N_29790);
xor UO_920 (O_920,N_29882,N_29588);
xor UO_921 (O_921,N_29488,N_29834);
or UO_922 (O_922,N_29804,N_29593);
nor UO_923 (O_923,N_29755,N_29879);
nor UO_924 (O_924,N_29569,N_29867);
and UO_925 (O_925,N_29509,N_29528);
and UO_926 (O_926,N_29877,N_29585);
nand UO_927 (O_927,N_29596,N_29699);
and UO_928 (O_928,N_29509,N_29642);
nor UO_929 (O_929,N_29654,N_29500);
and UO_930 (O_930,N_29816,N_29690);
xor UO_931 (O_931,N_29782,N_29613);
and UO_932 (O_932,N_29561,N_29629);
nor UO_933 (O_933,N_29477,N_29938);
nor UO_934 (O_934,N_29598,N_29521);
xnor UO_935 (O_935,N_29507,N_29854);
nor UO_936 (O_936,N_29473,N_29480);
or UO_937 (O_937,N_29625,N_29591);
nand UO_938 (O_938,N_29469,N_29925);
nor UO_939 (O_939,N_29835,N_29756);
xor UO_940 (O_940,N_29696,N_29554);
and UO_941 (O_941,N_29434,N_29479);
nor UO_942 (O_942,N_29759,N_29765);
nor UO_943 (O_943,N_29716,N_29735);
xor UO_944 (O_944,N_29424,N_29829);
xnor UO_945 (O_945,N_29978,N_29982);
xnor UO_946 (O_946,N_29408,N_29940);
nor UO_947 (O_947,N_29576,N_29538);
nand UO_948 (O_948,N_29763,N_29916);
xnor UO_949 (O_949,N_29830,N_29931);
xor UO_950 (O_950,N_29926,N_29962);
and UO_951 (O_951,N_29817,N_29590);
nor UO_952 (O_952,N_29813,N_29418);
and UO_953 (O_953,N_29427,N_29875);
nor UO_954 (O_954,N_29954,N_29507);
nor UO_955 (O_955,N_29772,N_29873);
nor UO_956 (O_956,N_29425,N_29428);
xor UO_957 (O_957,N_29515,N_29974);
and UO_958 (O_958,N_29833,N_29683);
nor UO_959 (O_959,N_29699,N_29568);
nand UO_960 (O_960,N_29913,N_29473);
or UO_961 (O_961,N_29681,N_29951);
or UO_962 (O_962,N_29866,N_29800);
nand UO_963 (O_963,N_29737,N_29899);
xor UO_964 (O_964,N_29667,N_29961);
xnor UO_965 (O_965,N_29497,N_29748);
xnor UO_966 (O_966,N_29808,N_29559);
xnor UO_967 (O_967,N_29506,N_29733);
xor UO_968 (O_968,N_29928,N_29650);
and UO_969 (O_969,N_29925,N_29973);
or UO_970 (O_970,N_29929,N_29813);
xnor UO_971 (O_971,N_29900,N_29590);
or UO_972 (O_972,N_29468,N_29692);
and UO_973 (O_973,N_29515,N_29983);
xor UO_974 (O_974,N_29929,N_29892);
and UO_975 (O_975,N_29768,N_29670);
nand UO_976 (O_976,N_29964,N_29688);
xor UO_977 (O_977,N_29557,N_29655);
or UO_978 (O_978,N_29496,N_29605);
nor UO_979 (O_979,N_29956,N_29606);
nor UO_980 (O_980,N_29802,N_29912);
nand UO_981 (O_981,N_29548,N_29505);
nor UO_982 (O_982,N_29929,N_29536);
nand UO_983 (O_983,N_29683,N_29717);
nor UO_984 (O_984,N_29492,N_29808);
or UO_985 (O_985,N_29746,N_29636);
nand UO_986 (O_986,N_29521,N_29733);
nand UO_987 (O_987,N_29581,N_29685);
and UO_988 (O_988,N_29852,N_29633);
nor UO_989 (O_989,N_29403,N_29520);
or UO_990 (O_990,N_29552,N_29922);
xnor UO_991 (O_991,N_29789,N_29737);
and UO_992 (O_992,N_29808,N_29491);
xor UO_993 (O_993,N_29839,N_29848);
and UO_994 (O_994,N_29441,N_29464);
xor UO_995 (O_995,N_29966,N_29442);
xor UO_996 (O_996,N_29581,N_29944);
nand UO_997 (O_997,N_29616,N_29621);
and UO_998 (O_998,N_29897,N_29766);
xnor UO_999 (O_999,N_29488,N_29993);
nand UO_1000 (O_1000,N_29413,N_29549);
nand UO_1001 (O_1001,N_29477,N_29780);
nor UO_1002 (O_1002,N_29723,N_29623);
or UO_1003 (O_1003,N_29915,N_29826);
xnor UO_1004 (O_1004,N_29660,N_29483);
or UO_1005 (O_1005,N_29505,N_29638);
and UO_1006 (O_1006,N_29634,N_29611);
nand UO_1007 (O_1007,N_29950,N_29553);
xor UO_1008 (O_1008,N_29562,N_29840);
nand UO_1009 (O_1009,N_29710,N_29659);
xor UO_1010 (O_1010,N_29697,N_29491);
nor UO_1011 (O_1011,N_29952,N_29425);
and UO_1012 (O_1012,N_29516,N_29557);
xnor UO_1013 (O_1013,N_29424,N_29465);
or UO_1014 (O_1014,N_29977,N_29897);
xor UO_1015 (O_1015,N_29647,N_29442);
nor UO_1016 (O_1016,N_29946,N_29437);
or UO_1017 (O_1017,N_29929,N_29704);
xnor UO_1018 (O_1018,N_29641,N_29829);
and UO_1019 (O_1019,N_29953,N_29998);
xor UO_1020 (O_1020,N_29691,N_29702);
nor UO_1021 (O_1021,N_29899,N_29657);
xnor UO_1022 (O_1022,N_29462,N_29724);
and UO_1023 (O_1023,N_29403,N_29663);
nand UO_1024 (O_1024,N_29403,N_29613);
or UO_1025 (O_1025,N_29605,N_29914);
xor UO_1026 (O_1026,N_29759,N_29890);
nand UO_1027 (O_1027,N_29587,N_29425);
or UO_1028 (O_1028,N_29679,N_29885);
nand UO_1029 (O_1029,N_29720,N_29996);
nor UO_1030 (O_1030,N_29560,N_29405);
nand UO_1031 (O_1031,N_29864,N_29918);
nand UO_1032 (O_1032,N_29453,N_29932);
xor UO_1033 (O_1033,N_29631,N_29934);
nand UO_1034 (O_1034,N_29493,N_29788);
xnor UO_1035 (O_1035,N_29906,N_29536);
nor UO_1036 (O_1036,N_29928,N_29729);
xnor UO_1037 (O_1037,N_29568,N_29428);
nor UO_1038 (O_1038,N_29975,N_29564);
or UO_1039 (O_1039,N_29742,N_29831);
and UO_1040 (O_1040,N_29471,N_29999);
and UO_1041 (O_1041,N_29902,N_29761);
nand UO_1042 (O_1042,N_29976,N_29430);
or UO_1043 (O_1043,N_29652,N_29630);
nor UO_1044 (O_1044,N_29418,N_29679);
xor UO_1045 (O_1045,N_29544,N_29993);
nand UO_1046 (O_1046,N_29627,N_29669);
nor UO_1047 (O_1047,N_29965,N_29737);
and UO_1048 (O_1048,N_29613,N_29596);
or UO_1049 (O_1049,N_29641,N_29719);
nand UO_1050 (O_1050,N_29811,N_29835);
nor UO_1051 (O_1051,N_29677,N_29879);
and UO_1052 (O_1052,N_29439,N_29869);
and UO_1053 (O_1053,N_29579,N_29721);
and UO_1054 (O_1054,N_29540,N_29723);
or UO_1055 (O_1055,N_29611,N_29890);
or UO_1056 (O_1056,N_29670,N_29963);
nand UO_1057 (O_1057,N_29967,N_29534);
xnor UO_1058 (O_1058,N_29726,N_29490);
nand UO_1059 (O_1059,N_29859,N_29410);
or UO_1060 (O_1060,N_29418,N_29886);
and UO_1061 (O_1061,N_29617,N_29979);
nor UO_1062 (O_1062,N_29849,N_29507);
nand UO_1063 (O_1063,N_29700,N_29802);
xor UO_1064 (O_1064,N_29977,N_29618);
nand UO_1065 (O_1065,N_29866,N_29563);
and UO_1066 (O_1066,N_29703,N_29798);
nor UO_1067 (O_1067,N_29473,N_29639);
xor UO_1068 (O_1068,N_29817,N_29442);
or UO_1069 (O_1069,N_29843,N_29606);
nand UO_1070 (O_1070,N_29881,N_29655);
and UO_1071 (O_1071,N_29681,N_29894);
xor UO_1072 (O_1072,N_29872,N_29406);
and UO_1073 (O_1073,N_29626,N_29712);
nor UO_1074 (O_1074,N_29781,N_29830);
nor UO_1075 (O_1075,N_29737,N_29401);
and UO_1076 (O_1076,N_29991,N_29471);
or UO_1077 (O_1077,N_29415,N_29525);
or UO_1078 (O_1078,N_29778,N_29574);
nor UO_1079 (O_1079,N_29773,N_29839);
xor UO_1080 (O_1080,N_29786,N_29406);
xor UO_1081 (O_1081,N_29820,N_29723);
nor UO_1082 (O_1082,N_29793,N_29557);
or UO_1083 (O_1083,N_29860,N_29952);
nand UO_1084 (O_1084,N_29770,N_29769);
nor UO_1085 (O_1085,N_29805,N_29453);
nor UO_1086 (O_1086,N_29723,N_29492);
nor UO_1087 (O_1087,N_29633,N_29909);
and UO_1088 (O_1088,N_29740,N_29802);
nor UO_1089 (O_1089,N_29466,N_29983);
nand UO_1090 (O_1090,N_29552,N_29421);
xor UO_1091 (O_1091,N_29901,N_29875);
and UO_1092 (O_1092,N_29724,N_29655);
nor UO_1093 (O_1093,N_29838,N_29720);
and UO_1094 (O_1094,N_29884,N_29886);
or UO_1095 (O_1095,N_29917,N_29762);
nor UO_1096 (O_1096,N_29569,N_29606);
nand UO_1097 (O_1097,N_29658,N_29801);
and UO_1098 (O_1098,N_29435,N_29462);
nor UO_1099 (O_1099,N_29519,N_29585);
nand UO_1100 (O_1100,N_29496,N_29543);
and UO_1101 (O_1101,N_29968,N_29927);
and UO_1102 (O_1102,N_29483,N_29990);
xor UO_1103 (O_1103,N_29686,N_29595);
xor UO_1104 (O_1104,N_29472,N_29732);
and UO_1105 (O_1105,N_29699,N_29575);
and UO_1106 (O_1106,N_29854,N_29737);
and UO_1107 (O_1107,N_29773,N_29554);
and UO_1108 (O_1108,N_29766,N_29749);
xor UO_1109 (O_1109,N_29747,N_29764);
nand UO_1110 (O_1110,N_29553,N_29674);
and UO_1111 (O_1111,N_29769,N_29483);
nand UO_1112 (O_1112,N_29523,N_29632);
xnor UO_1113 (O_1113,N_29803,N_29925);
or UO_1114 (O_1114,N_29771,N_29645);
or UO_1115 (O_1115,N_29770,N_29688);
or UO_1116 (O_1116,N_29525,N_29455);
nand UO_1117 (O_1117,N_29474,N_29783);
and UO_1118 (O_1118,N_29411,N_29619);
or UO_1119 (O_1119,N_29488,N_29496);
and UO_1120 (O_1120,N_29525,N_29774);
and UO_1121 (O_1121,N_29428,N_29685);
and UO_1122 (O_1122,N_29965,N_29772);
or UO_1123 (O_1123,N_29735,N_29595);
nand UO_1124 (O_1124,N_29875,N_29841);
nand UO_1125 (O_1125,N_29924,N_29854);
or UO_1126 (O_1126,N_29590,N_29693);
nand UO_1127 (O_1127,N_29595,N_29831);
and UO_1128 (O_1128,N_29518,N_29680);
nand UO_1129 (O_1129,N_29529,N_29945);
nor UO_1130 (O_1130,N_29912,N_29574);
nand UO_1131 (O_1131,N_29535,N_29884);
nand UO_1132 (O_1132,N_29689,N_29463);
and UO_1133 (O_1133,N_29864,N_29668);
or UO_1134 (O_1134,N_29862,N_29795);
and UO_1135 (O_1135,N_29519,N_29538);
or UO_1136 (O_1136,N_29797,N_29668);
or UO_1137 (O_1137,N_29960,N_29585);
nor UO_1138 (O_1138,N_29619,N_29716);
nand UO_1139 (O_1139,N_29927,N_29570);
xnor UO_1140 (O_1140,N_29495,N_29405);
and UO_1141 (O_1141,N_29551,N_29857);
or UO_1142 (O_1142,N_29535,N_29687);
xor UO_1143 (O_1143,N_29780,N_29769);
nor UO_1144 (O_1144,N_29930,N_29736);
nand UO_1145 (O_1145,N_29630,N_29529);
or UO_1146 (O_1146,N_29935,N_29914);
and UO_1147 (O_1147,N_29613,N_29646);
nor UO_1148 (O_1148,N_29531,N_29548);
nor UO_1149 (O_1149,N_29642,N_29488);
nand UO_1150 (O_1150,N_29469,N_29672);
and UO_1151 (O_1151,N_29479,N_29501);
xnor UO_1152 (O_1152,N_29411,N_29840);
nor UO_1153 (O_1153,N_29521,N_29403);
nand UO_1154 (O_1154,N_29541,N_29796);
and UO_1155 (O_1155,N_29462,N_29781);
nor UO_1156 (O_1156,N_29558,N_29501);
nand UO_1157 (O_1157,N_29737,N_29716);
nor UO_1158 (O_1158,N_29632,N_29982);
and UO_1159 (O_1159,N_29430,N_29555);
or UO_1160 (O_1160,N_29965,N_29739);
and UO_1161 (O_1161,N_29714,N_29843);
nand UO_1162 (O_1162,N_29484,N_29901);
nor UO_1163 (O_1163,N_29471,N_29911);
nor UO_1164 (O_1164,N_29740,N_29603);
and UO_1165 (O_1165,N_29449,N_29536);
and UO_1166 (O_1166,N_29820,N_29591);
or UO_1167 (O_1167,N_29918,N_29767);
or UO_1168 (O_1168,N_29591,N_29407);
nor UO_1169 (O_1169,N_29681,N_29640);
and UO_1170 (O_1170,N_29800,N_29857);
xor UO_1171 (O_1171,N_29704,N_29705);
nand UO_1172 (O_1172,N_29754,N_29509);
or UO_1173 (O_1173,N_29677,N_29451);
nor UO_1174 (O_1174,N_29712,N_29802);
and UO_1175 (O_1175,N_29842,N_29401);
and UO_1176 (O_1176,N_29562,N_29577);
nand UO_1177 (O_1177,N_29698,N_29942);
or UO_1178 (O_1178,N_29878,N_29923);
nand UO_1179 (O_1179,N_29621,N_29624);
nor UO_1180 (O_1180,N_29685,N_29716);
nor UO_1181 (O_1181,N_29983,N_29479);
nor UO_1182 (O_1182,N_29823,N_29989);
and UO_1183 (O_1183,N_29733,N_29539);
or UO_1184 (O_1184,N_29520,N_29417);
and UO_1185 (O_1185,N_29836,N_29838);
or UO_1186 (O_1186,N_29568,N_29731);
xnor UO_1187 (O_1187,N_29936,N_29721);
and UO_1188 (O_1188,N_29645,N_29433);
nand UO_1189 (O_1189,N_29911,N_29620);
nor UO_1190 (O_1190,N_29511,N_29431);
nand UO_1191 (O_1191,N_29560,N_29577);
and UO_1192 (O_1192,N_29921,N_29826);
and UO_1193 (O_1193,N_29589,N_29854);
xor UO_1194 (O_1194,N_29505,N_29859);
xor UO_1195 (O_1195,N_29820,N_29943);
xor UO_1196 (O_1196,N_29402,N_29851);
and UO_1197 (O_1197,N_29910,N_29756);
nand UO_1198 (O_1198,N_29975,N_29692);
and UO_1199 (O_1199,N_29888,N_29930);
or UO_1200 (O_1200,N_29561,N_29709);
xnor UO_1201 (O_1201,N_29403,N_29850);
or UO_1202 (O_1202,N_29755,N_29486);
nand UO_1203 (O_1203,N_29837,N_29542);
nor UO_1204 (O_1204,N_29417,N_29867);
nand UO_1205 (O_1205,N_29725,N_29804);
or UO_1206 (O_1206,N_29665,N_29508);
xnor UO_1207 (O_1207,N_29716,N_29905);
nor UO_1208 (O_1208,N_29994,N_29853);
and UO_1209 (O_1209,N_29897,N_29872);
or UO_1210 (O_1210,N_29539,N_29747);
nor UO_1211 (O_1211,N_29853,N_29857);
nand UO_1212 (O_1212,N_29972,N_29700);
nand UO_1213 (O_1213,N_29550,N_29996);
and UO_1214 (O_1214,N_29516,N_29584);
xor UO_1215 (O_1215,N_29470,N_29720);
and UO_1216 (O_1216,N_29658,N_29956);
nand UO_1217 (O_1217,N_29793,N_29989);
nor UO_1218 (O_1218,N_29782,N_29937);
nand UO_1219 (O_1219,N_29598,N_29613);
nor UO_1220 (O_1220,N_29543,N_29670);
and UO_1221 (O_1221,N_29770,N_29668);
xnor UO_1222 (O_1222,N_29645,N_29472);
nor UO_1223 (O_1223,N_29906,N_29941);
nand UO_1224 (O_1224,N_29931,N_29597);
and UO_1225 (O_1225,N_29896,N_29617);
nor UO_1226 (O_1226,N_29420,N_29503);
nand UO_1227 (O_1227,N_29842,N_29922);
nor UO_1228 (O_1228,N_29649,N_29579);
xor UO_1229 (O_1229,N_29830,N_29858);
or UO_1230 (O_1230,N_29736,N_29632);
nand UO_1231 (O_1231,N_29422,N_29925);
or UO_1232 (O_1232,N_29568,N_29940);
xnor UO_1233 (O_1233,N_29403,N_29658);
xnor UO_1234 (O_1234,N_29401,N_29593);
and UO_1235 (O_1235,N_29921,N_29444);
xor UO_1236 (O_1236,N_29812,N_29863);
or UO_1237 (O_1237,N_29906,N_29635);
and UO_1238 (O_1238,N_29646,N_29501);
nand UO_1239 (O_1239,N_29545,N_29785);
or UO_1240 (O_1240,N_29698,N_29859);
and UO_1241 (O_1241,N_29864,N_29530);
or UO_1242 (O_1242,N_29443,N_29521);
or UO_1243 (O_1243,N_29527,N_29432);
nand UO_1244 (O_1244,N_29676,N_29792);
and UO_1245 (O_1245,N_29839,N_29907);
xnor UO_1246 (O_1246,N_29896,N_29947);
or UO_1247 (O_1247,N_29856,N_29449);
or UO_1248 (O_1248,N_29920,N_29533);
or UO_1249 (O_1249,N_29554,N_29850);
and UO_1250 (O_1250,N_29617,N_29735);
nor UO_1251 (O_1251,N_29822,N_29977);
nor UO_1252 (O_1252,N_29882,N_29541);
and UO_1253 (O_1253,N_29447,N_29480);
and UO_1254 (O_1254,N_29677,N_29975);
and UO_1255 (O_1255,N_29623,N_29816);
and UO_1256 (O_1256,N_29870,N_29695);
or UO_1257 (O_1257,N_29661,N_29875);
xor UO_1258 (O_1258,N_29927,N_29939);
or UO_1259 (O_1259,N_29997,N_29854);
and UO_1260 (O_1260,N_29927,N_29522);
nor UO_1261 (O_1261,N_29506,N_29997);
nand UO_1262 (O_1262,N_29625,N_29567);
or UO_1263 (O_1263,N_29448,N_29649);
or UO_1264 (O_1264,N_29485,N_29438);
xor UO_1265 (O_1265,N_29566,N_29933);
or UO_1266 (O_1266,N_29484,N_29496);
or UO_1267 (O_1267,N_29949,N_29824);
xnor UO_1268 (O_1268,N_29679,N_29513);
or UO_1269 (O_1269,N_29660,N_29894);
or UO_1270 (O_1270,N_29793,N_29797);
nand UO_1271 (O_1271,N_29608,N_29429);
nor UO_1272 (O_1272,N_29480,N_29868);
and UO_1273 (O_1273,N_29476,N_29904);
and UO_1274 (O_1274,N_29427,N_29805);
nor UO_1275 (O_1275,N_29447,N_29966);
nand UO_1276 (O_1276,N_29425,N_29899);
or UO_1277 (O_1277,N_29971,N_29637);
nor UO_1278 (O_1278,N_29862,N_29798);
nand UO_1279 (O_1279,N_29765,N_29642);
nand UO_1280 (O_1280,N_29823,N_29434);
or UO_1281 (O_1281,N_29433,N_29854);
xor UO_1282 (O_1282,N_29856,N_29670);
or UO_1283 (O_1283,N_29635,N_29679);
or UO_1284 (O_1284,N_29851,N_29576);
nor UO_1285 (O_1285,N_29935,N_29930);
xor UO_1286 (O_1286,N_29727,N_29584);
nand UO_1287 (O_1287,N_29529,N_29952);
or UO_1288 (O_1288,N_29655,N_29839);
and UO_1289 (O_1289,N_29721,N_29986);
xnor UO_1290 (O_1290,N_29489,N_29414);
or UO_1291 (O_1291,N_29733,N_29645);
nand UO_1292 (O_1292,N_29506,N_29536);
or UO_1293 (O_1293,N_29532,N_29791);
nor UO_1294 (O_1294,N_29564,N_29508);
or UO_1295 (O_1295,N_29443,N_29423);
or UO_1296 (O_1296,N_29974,N_29424);
xor UO_1297 (O_1297,N_29715,N_29563);
or UO_1298 (O_1298,N_29448,N_29513);
or UO_1299 (O_1299,N_29408,N_29457);
or UO_1300 (O_1300,N_29405,N_29824);
and UO_1301 (O_1301,N_29696,N_29737);
nor UO_1302 (O_1302,N_29699,N_29985);
or UO_1303 (O_1303,N_29915,N_29763);
xor UO_1304 (O_1304,N_29672,N_29891);
xor UO_1305 (O_1305,N_29816,N_29548);
xor UO_1306 (O_1306,N_29527,N_29943);
or UO_1307 (O_1307,N_29479,N_29690);
xnor UO_1308 (O_1308,N_29404,N_29821);
nor UO_1309 (O_1309,N_29807,N_29910);
nor UO_1310 (O_1310,N_29988,N_29544);
nand UO_1311 (O_1311,N_29406,N_29413);
or UO_1312 (O_1312,N_29653,N_29552);
and UO_1313 (O_1313,N_29673,N_29780);
nor UO_1314 (O_1314,N_29938,N_29984);
nand UO_1315 (O_1315,N_29567,N_29649);
nor UO_1316 (O_1316,N_29533,N_29669);
nor UO_1317 (O_1317,N_29503,N_29828);
nand UO_1318 (O_1318,N_29983,N_29842);
nor UO_1319 (O_1319,N_29800,N_29940);
xnor UO_1320 (O_1320,N_29881,N_29841);
and UO_1321 (O_1321,N_29817,N_29850);
and UO_1322 (O_1322,N_29772,N_29472);
xnor UO_1323 (O_1323,N_29825,N_29440);
and UO_1324 (O_1324,N_29540,N_29613);
nor UO_1325 (O_1325,N_29638,N_29769);
xor UO_1326 (O_1326,N_29862,N_29941);
and UO_1327 (O_1327,N_29890,N_29429);
nor UO_1328 (O_1328,N_29432,N_29521);
and UO_1329 (O_1329,N_29411,N_29905);
xnor UO_1330 (O_1330,N_29947,N_29511);
nand UO_1331 (O_1331,N_29900,N_29674);
and UO_1332 (O_1332,N_29596,N_29944);
nor UO_1333 (O_1333,N_29562,N_29926);
nand UO_1334 (O_1334,N_29928,N_29655);
and UO_1335 (O_1335,N_29785,N_29647);
nand UO_1336 (O_1336,N_29953,N_29504);
or UO_1337 (O_1337,N_29615,N_29736);
xnor UO_1338 (O_1338,N_29406,N_29807);
nor UO_1339 (O_1339,N_29900,N_29721);
and UO_1340 (O_1340,N_29475,N_29906);
nand UO_1341 (O_1341,N_29903,N_29813);
and UO_1342 (O_1342,N_29767,N_29932);
and UO_1343 (O_1343,N_29750,N_29852);
nand UO_1344 (O_1344,N_29733,N_29816);
nor UO_1345 (O_1345,N_29759,N_29470);
or UO_1346 (O_1346,N_29799,N_29886);
xor UO_1347 (O_1347,N_29620,N_29498);
nand UO_1348 (O_1348,N_29506,N_29598);
nor UO_1349 (O_1349,N_29742,N_29480);
nand UO_1350 (O_1350,N_29954,N_29437);
xnor UO_1351 (O_1351,N_29448,N_29888);
and UO_1352 (O_1352,N_29507,N_29417);
nand UO_1353 (O_1353,N_29500,N_29538);
nand UO_1354 (O_1354,N_29540,N_29864);
nand UO_1355 (O_1355,N_29761,N_29744);
and UO_1356 (O_1356,N_29894,N_29509);
and UO_1357 (O_1357,N_29703,N_29628);
or UO_1358 (O_1358,N_29679,N_29694);
and UO_1359 (O_1359,N_29843,N_29979);
nand UO_1360 (O_1360,N_29420,N_29819);
and UO_1361 (O_1361,N_29425,N_29778);
nor UO_1362 (O_1362,N_29837,N_29740);
or UO_1363 (O_1363,N_29822,N_29952);
nand UO_1364 (O_1364,N_29993,N_29669);
nor UO_1365 (O_1365,N_29858,N_29942);
xor UO_1366 (O_1366,N_29400,N_29579);
nor UO_1367 (O_1367,N_29427,N_29810);
nor UO_1368 (O_1368,N_29513,N_29426);
nand UO_1369 (O_1369,N_29698,N_29816);
nand UO_1370 (O_1370,N_29577,N_29556);
nand UO_1371 (O_1371,N_29425,N_29532);
nor UO_1372 (O_1372,N_29576,N_29504);
nor UO_1373 (O_1373,N_29536,N_29927);
nand UO_1374 (O_1374,N_29734,N_29937);
or UO_1375 (O_1375,N_29864,N_29952);
xor UO_1376 (O_1376,N_29615,N_29548);
nor UO_1377 (O_1377,N_29410,N_29888);
and UO_1378 (O_1378,N_29496,N_29759);
and UO_1379 (O_1379,N_29519,N_29652);
and UO_1380 (O_1380,N_29900,N_29759);
and UO_1381 (O_1381,N_29604,N_29735);
and UO_1382 (O_1382,N_29538,N_29718);
or UO_1383 (O_1383,N_29760,N_29948);
and UO_1384 (O_1384,N_29895,N_29499);
nand UO_1385 (O_1385,N_29641,N_29618);
xor UO_1386 (O_1386,N_29431,N_29680);
nand UO_1387 (O_1387,N_29559,N_29589);
xnor UO_1388 (O_1388,N_29644,N_29616);
xor UO_1389 (O_1389,N_29773,N_29624);
nor UO_1390 (O_1390,N_29868,N_29534);
and UO_1391 (O_1391,N_29648,N_29652);
nand UO_1392 (O_1392,N_29795,N_29937);
nor UO_1393 (O_1393,N_29474,N_29431);
or UO_1394 (O_1394,N_29666,N_29452);
nand UO_1395 (O_1395,N_29886,N_29839);
xnor UO_1396 (O_1396,N_29553,N_29952);
xor UO_1397 (O_1397,N_29980,N_29662);
xnor UO_1398 (O_1398,N_29667,N_29588);
or UO_1399 (O_1399,N_29841,N_29678);
nor UO_1400 (O_1400,N_29582,N_29913);
or UO_1401 (O_1401,N_29439,N_29517);
xnor UO_1402 (O_1402,N_29623,N_29508);
or UO_1403 (O_1403,N_29401,N_29908);
nor UO_1404 (O_1404,N_29647,N_29894);
xnor UO_1405 (O_1405,N_29542,N_29626);
nor UO_1406 (O_1406,N_29520,N_29925);
nor UO_1407 (O_1407,N_29597,N_29510);
nor UO_1408 (O_1408,N_29539,N_29709);
and UO_1409 (O_1409,N_29925,N_29895);
or UO_1410 (O_1410,N_29454,N_29908);
and UO_1411 (O_1411,N_29533,N_29977);
and UO_1412 (O_1412,N_29503,N_29896);
nor UO_1413 (O_1413,N_29671,N_29559);
and UO_1414 (O_1414,N_29742,N_29488);
and UO_1415 (O_1415,N_29688,N_29785);
or UO_1416 (O_1416,N_29608,N_29480);
or UO_1417 (O_1417,N_29634,N_29797);
and UO_1418 (O_1418,N_29512,N_29564);
and UO_1419 (O_1419,N_29495,N_29498);
nor UO_1420 (O_1420,N_29822,N_29914);
nor UO_1421 (O_1421,N_29678,N_29928);
and UO_1422 (O_1422,N_29931,N_29624);
nand UO_1423 (O_1423,N_29490,N_29585);
and UO_1424 (O_1424,N_29746,N_29995);
xnor UO_1425 (O_1425,N_29732,N_29753);
and UO_1426 (O_1426,N_29837,N_29472);
or UO_1427 (O_1427,N_29944,N_29623);
and UO_1428 (O_1428,N_29873,N_29519);
xnor UO_1429 (O_1429,N_29781,N_29542);
or UO_1430 (O_1430,N_29627,N_29423);
xnor UO_1431 (O_1431,N_29545,N_29514);
xor UO_1432 (O_1432,N_29970,N_29462);
nand UO_1433 (O_1433,N_29663,N_29913);
xor UO_1434 (O_1434,N_29904,N_29541);
xor UO_1435 (O_1435,N_29419,N_29947);
and UO_1436 (O_1436,N_29583,N_29806);
xnor UO_1437 (O_1437,N_29917,N_29404);
and UO_1438 (O_1438,N_29755,N_29588);
or UO_1439 (O_1439,N_29422,N_29881);
and UO_1440 (O_1440,N_29675,N_29941);
or UO_1441 (O_1441,N_29915,N_29911);
nand UO_1442 (O_1442,N_29875,N_29405);
nand UO_1443 (O_1443,N_29716,N_29414);
or UO_1444 (O_1444,N_29650,N_29421);
or UO_1445 (O_1445,N_29982,N_29799);
nand UO_1446 (O_1446,N_29629,N_29824);
nor UO_1447 (O_1447,N_29453,N_29585);
nor UO_1448 (O_1448,N_29502,N_29597);
nor UO_1449 (O_1449,N_29903,N_29740);
xnor UO_1450 (O_1450,N_29723,N_29927);
nand UO_1451 (O_1451,N_29741,N_29959);
xnor UO_1452 (O_1452,N_29987,N_29444);
and UO_1453 (O_1453,N_29818,N_29680);
nor UO_1454 (O_1454,N_29540,N_29501);
nor UO_1455 (O_1455,N_29942,N_29800);
and UO_1456 (O_1456,N_29913,N_29559);
nor UO_1457 (O_1457,N_29509,N_29812);
xor UO_1458 (O_1458,N_29648,N_29501);
or UO_1459 (O_1459,N_29695,N_29826);
and UO_1460 (O_1460,N_29718,N_29872);
and UO_1461 (O_1461,N_29539,N_29705);
nand UO_1462 (O_1462,N_29431,N_29490);
and UO_1463 (O_1463,N_29517,N_29705);
nand UO_1464 (O_1464,N_29585,N_29836);
nand UO_1465 (O_1465,N_29896,N_29555);
nor UO_1466 (O_1466,N_29569,N_29587);
nor UO_1467 (O_1467,N_29781,N_29443);
nor UO_1468 (O_1468,N_29457,N_29512);
and UO_1469 (O_1469,N_29891,N_29613);
nor UO_1470 (O_1470,N_29997,N_29639);
or UO_1471 (O_1471,N_29562,N_29435);
nand UO_1472 (O_1472,N_29928,N_29660);
xnor UO_1473 (O_1473,N_29489,N_29942);
or UO_1474 (O_1474,N_29455,N_29625);
nor UO_1475 (O_1475,N_29554,N_29477);
or UO_1476 (O_1476,N_29881,N_29948);
or UO_1477 (O_1477,N_29660,N_29548);
and UO_1478 (O_1478,N_29412,N_29758);
nor UO_1479 (O_1479,N_29587,N_29484);
or UO_1480 (O_1480,N_29559,N_29926);
and UO_1481 (O_1481,N_29828,N_29563);
nor UO_1482 (O_1482,N_29938,N_29810);
and UO_1483 (O_1483,N_29709,N_29471);
xor UO_1484 (O_1484,N_29445,N_29430);
nand UO_1485 (O_1485,N_29498,N_29985);
or UO_1486 (O_1486,N_29450,N_29885);
nand UO_1487 (O_1487,N_29560,N_29614);
xor UO_1488 (O_1488,N_29642,N_29761);
xnor UO_1489 (O_1489,N_29596,N_29510);
and UO_1490 (O_1490,N_29426,N_29554);
nand UO_1491 (O_1491,N_29838,N_29992);
or UO_1492 (O_1492,N_29645,N_29615);
and UO_1493 (O_1493,N_29663,N_29886);
nand UO_1494 (O_1494,N_29946,N_29602);
nand UO_1495 (O_1495,N_29934,N_29633);
or UO_1496 (O_1496,N_29503,N_29712);
nor UO_1497 (O_1497,N_29570,N_29783);
xnor UO_1498 (O_1498,N_29475,N_29931);
nand UO_1499 (O_1499,N_29506,N_29508);
nor UO_1500 (O_1500,N_29921,N_29594);
nand UO_1501 (O_1501,N_29726,N_29592);
and UO_1502 (O_1502,N_29706,N_29886);
and UO_1503 (O_1503,N_29503,N_29402);
and UO_1504 (O_1504,N_29966,N_29774);
nor UO_1505 (O_1505,N_29734,N_29610);
or UO_1506 (O_1506,N_29854,N_29631);
xor UO_1507 (O_1507,N_29510,N_29640);
xor UO_1508 (O_1508,N_29905,N_29748);
nand UO_1509 (O_1509,N_29792,N_29667);
xor UO_1510 (O_1510,N_29477,N_29466);
xnor UO_1511 (O_1511,N_29611,N_29708);
and UO_1512 (O_1512,N_29638,N_29456);
nand UO_1513 (O_1513,N_29776,N_29524);
xnor UO_1514 (O_1514,N_29423,N_29774);
nor UO_1515 (O_1515,N_29479,N_29569);
and UO_1516 (O_1516,N_29482,N_29837);
and UO_1517 (O_1517,N_29640,N_29474);
or UO_1518 (O_1518,N_29941,N_29968);
or UO_1519 (O_1519,N_29888,N_29938);
or UO_1520 (O_1520,N_29871,N_29765);
and UO_1521 (O_1521,N_29863,N_29875);
xnor UO_1522 (O_1522,N_29736,N_29924);
nand UO_1523 (O_1523,N_29513,N_29431);
and UO_1524 (O_1524,N_29816,N_29527);
nand UO_1525 (O_1525,N_29768,N_29413);
and UO_1526 (O_1526,N_29910,N_29993);
or UO_1527 (O_1527,N_29546,N_29434);
and UO_1528 (O_1528,N_29465,N_29985);
and UO_1529 (O_1529,N_29858,N_29665);
and UO_1530 (O_1530,N_29844,N_29463);
and UO_1531 (O_1531,N_29647,N_29789);
xnor UO_1532 (O_1532,N_29637,N_29561);
nor UO_1533 (O_1533,N_29676,N_29613);
nand UO_1534 (O_1534,N_29713,N_29725);
nand UO_1535 (O_1535,N_29444,N_29811);
nand UO_1536 (O_1536,N_29842,N_29691);
nand UO_1537 (O_1537,N_29608,N_29472);
xnor UO_1538 (O_1538,N_29443,N_29637);
or UO_1539 (O_1539,N_29475,N_29726);
and UO_1540 (O_1540,N_29798,N_29934);
nor UO_1541 (O_1541,N_29938,N_29533);
and UO_1542 (O_1542,N_29430,N_29746);
or UO_1543 (O_1543,N_29812,N_29732);
or UO_1544 (O_1544,N_29583,N_29402);
or UO_1545 (O_1545,N_29739,N_29788);
nand UO_1546 (O_1546,N_29450,N_29519);
xnor UO_1547 (O_1547,N_29470,N_29755);
or UO_1548 (O_1548,N_29470,N_29919);
nand UO_1549 (O_1549,N_29863,N_29910);
and UO_1550 (O_1550,N_29654,N_29749);
xnor UO_1551 (O_1551,N_29998,N_29732);
nand UO_1552 (O_1552,N_29920,N_29580);
or UO_1553 (O_1553,N_29451,N_29792);
and UO_1554 (O_1554,N_29428,N_29500);
xor UO_1555 (O_1555,N_29729,N_29660);
and UO_1556 (O_1556,N_29570,N_29434);
and UO_1557 (O_1557,N_29656,N_29565);
xnor UO_1558 (O_1558,N_29571,N_29840);
xor UO_1559 (O_1559,N_29753,N_29678);
xnor UO_1560 (O_1560,N_29920,N_29882);
nand UO_1561 (O_1561,N_29723,N_29781);
xnor UO_1562 (O_1562,N_29878,N_29516);
or UO_1563 (O_1563,N_29760,N_29853);
nand UO_1564 (O_1564,N_29690,N_29573);
nand UO_1565 (O_1565,N_29897,N_29710);
nand UO_1566 (O_1566,N_29993,N_29878);
or UO_1567 (O_1567,N_29479,N_29813);
xnor UO_1568 (O_1568,N_29944,N_29543);
nor UO_1569 (O_1569,N_29631,N_29422);
nor UO_1570 (O_1570,N_29603,N_29575);
nand UO_1571 (O_1571,N_29502,N_29911);
nor UO_1572 (O_1572,N_29924,N_29556);
xor UO_1573 (O_1573,N_29848,N_29424);
nand UO_1574 (O_1574,N_29676,N_29540);
nand UO_1575 (O_1575,N_29637,N_29689);
or UO_1576 (O_1576,N_29686,N_29418);
nor UO_1577 (O_1577,N_29628,N_29638);
nand UO_1578 (O_1578,N_29574,N_29957);
xor UO_1579 (O_1579,N_29867,N_29931);
nand UO_1580 (O_1580,N_29428,N_29966);
nand UO_1581 (O_1581,N_29591,N_29684);
nor UO_1582 (O_1582,N_29928,N_29691);
or UO_1583 (O_1583,N_29501,N_29429);
and UO_1584 (O_1584,N_29720,N_29411);
and UO_1585 (O_1585,N_29635,N_29822);
and UO_1586 (O_1586,N_29940,N_29692);
nand UO_1587 (O_1587,N_29521,N_29675);
xor UO_1588 (O_1588,N_29767,N_29497);
nand UO_1589 (O_1589,N_29473,N_29680);
and UO_1590 (O_1590,N_29914,N_29668);
and UO_1591 (O_1591,N_29963,N_29856);
and UO_1592 (O_1592,N_29929,N_29628);
nand UO_1593 (O_1593,N_29877,N_29485);
nand UO_1594 (O_1594,N_29417,N_29960);
nor UO_1595 (O_1595,N_29692,N_29562);
nand UO_1596 (O_1596,N_29804,N_29862);
nor UO_1597 (O_1597,N_29828,N_29802);
or UO_1598 (O_1598,N_29482,N_29844);
nor UO_1599 (O_1599,N_29759,N_29565);
or UO_1600 (O_1600,N_29731,N_29899);
and UO_1601 (O_1601,N_29537,N_29503);
or UO_1602 (O_1602,N_29483,N_29935);
xnor UO_1603 (O_1603,N_29793,N_29787);
nor UO_1604 (O_1604,N_29446,N_29626);
or UO_1605 (O_1605,N_29736,N_29413);
and UO_1606 (O_1606,N_29528,N_29477);
xnor UO_1607 (O_1607,N_29972,N_29985);
and UO_1608 (O_1608,N_29583,N_29466);
xor UO_1609 (O_1609,N_29899,N_29627);
nor UO_1610 (O_1610,N_29910,N_29987);
or UO_1611 (O_1611,N_29887,N_29646);
or UO_1612 (O_1612,N_29487,N_29463);
nor UO_1613 (O_1613,N_29931,N_29479);
xor UO_1614 (O_1614,N_29803,N_29541);
xor UO_1615 (O_1615,N_29966,N_29602);
and UO_1616 (O_1616,N_29474,N_29972);
nor UO_1617 (O_1617,N_29809,N_29748);
xnor UO_1618 (O_1618,N_29756,N_29665);
xor UO_1619 (O_1619,N_29604,N_29566);
or UO_1620 (O_1620,N_29803,N_29919);
and UO_1621 (O_1621,N_29985,N_29996);
or UO_1622 (O_1622,N_29769,N_29440);
or UO_1623 (O_1623,N_29780,N_29537);
nand UO_1624 (O_1624,N_29786,N_29748);
and UO_1625 (O_1625,N_29742,N_29709);
xor UO_1626 (O_1626,N_29466,N_29699);
nand UO_1627 (O_1627,N_29455,N_29553);
and UO_1628 (O_1628,N_29549,N_29805);
or UO_1629 (O_1629,N_29773,N_29556);
nor UO_1630 (O_1630,N_29620,N_29409);
xor UO_1631 (O_1631,N_29999,N_29861);
nand UO_1632 (O_1632,N_29994,N_29526);
or UO_1633 (O_1633,N_29545,N_29689);
and UO_1634 (O_1634,N_29665,N_29583);
and UO_1635 (O_1635,N_29841,N_29949);
or UO_1636 (O_1636,N_29775,N_29484);
or UO_1637 (O_1637,N_29575,N_29426);
xnor UO_1638 (O_1638,N_29928,N_29693);
nor UO_1639 (O_1639,N_29909,N_29607);
xor UO_1640 (O_1640,N_29704,N_29502);
nand UO_1641 (O_1641,N_29980,N_29866);
xor UO_1642 (O_1642,N_29750,N_29507);
or UO_1643 (O_1643,N_29419,N_29852);
and UO_1644 (O_1644,N_29879,N_29999);
or UO_1645 (O_1645,N_29516,N_29968);
xor UO_1646 (O_1646,N_29763,N_29968);
xnor UO_1647 (O_1647,N_29721,N_29603);
and UO_1648 (O_1648,N_29627,N_29799);
and UO_1649 (O_1649,N_29562,N_29473);
xnor UO_1650 (O_1650,N_29465,N_29436);
or UO_1651 (O_1651,N_29876,N_29927);
or UO_1652 (O_1652,N_29934,N_29488);
xnor UO_1653 (O_1653,N_29439,N_29981);
nand UO_1654 (O_1654,N_29677,N_29528);
xor UO_1655 (O_1655,N_29476,N_29930);
and UO_1656 (O_1656,N_29931,N_29848);
and UO_1657 (O_1657,N_29724,N_29517);
nor UO_1658 (O_1658,N_29761,N_29679);
nor UO_1659 (O_1659,N_29693,N_29955);
nor UO_1660 (O_1660,N_29640,N_29567);
or UO_1661 (O_1661,N_29809,N_29514);
nor UO_1662 (O_1662,N_29631,N_29541);
nand UO_1663 (O_1663,N_29648,N_29735);
or UO_1664 (O_1664,N_29874,N_29748);
xor UO_1665 (O_1665,N_29524,N_29903);
nor UO_1666 (O_1666,N_29773,N_29757);
nor UO_1667 (O_1667,N_29786,N_29536);
nor UO_1668 (O_1668,N_29558,N_29803);
or UO_1669 (O_1669,N_29659,N_29619);
or UO_1670 (O_1670,N_29633,N_29754);
nand UO_1671 (O_1671,N_29817,N_29857);
xnor UO_1672 (O_1672,N_29575,N_29935);
and UO_1673 (O_1673,N_29404,N_29911);
or UO_1674 (O_1674,N_29760,N_29894);
nor UO_1675 (O_1675,N_29512,N_29949);
xor UO_1676 (O_1676,N_29528,N_29967);
or UO_1677 (O_1677,N_29985,N_29611);
or UO_1678 (O_1678,N_29870,N_29781);
nor UO_1679 (O_1679,N_29973,N_29719);
or UO_1680 (O_1680,N_29782,N_29570);
nand UO_1681 (O_1681,N_29454,N_29476);
and UO_1682 (O_1682,N_29538,N_29794);
xor UO_1683 (O_1683,N_29882,N_29419);
or UO_1684 (O_1684,N_29635,N_29429);
nor UO_1685 (O_1685,N_29933,N_29643);
xor UO_1686 (O_1686,N_29475,N_29848);
nand UO_1687 (O_1687,N_29623,N_29689);
and UO_1688 (O_1688,N_29409,N_29489);
nor UO_1689 (O_1689,N_29555,N_29989);
nand UO_1690 (O_1690,N_29612,N_29861);
nand UO_1691 (O_1691,N_29417,N_29743);
nor UO_1692 (O_1692,N_29760,N_29542);
or UO_1693 (O_1693,N_29898,N_29723);
and UO_1694 (O_1694,N_29739,N_29885);
nand UO_1695 (O_1695,N_29404,N_29813);
xor UO_1696 (O_1696,N_29531,N_29870);
or UO_1697 (O_1697,N_29859,N_29689);
and UO_1698 (O_1698,N_29563,N_29656);
nor UO_1699 (O_1699,N_29655,N_29738);
or UO_1700 (O_1700,N_29722,N_29971);
nand UO_1701 (O_1701,N_29943,N_29443);
and UO_1702 (O_1702,N_29471,N_29962);
nor UO_1703 (O_1703,N_29613,N_29931);
xnor UO_1704 (O_1704,N_29446,N_29669);
nand UO_1705 (O_1705,N_29815,N_29620);
nand UO_1706 (O_1706,N_29590,N_29521);
and UO_1707 (O_1707,N_29569,N_29618);
and UO_1708 (O_1708,N_29550,N_29707);
and UO_1709 (O_1709,N_29609,N_29616);
or UO_1710 (O_1710,N_29458,N_29506);
and UO_1711 (O_1711,N_29937,N_29604);
and UO_1712 (O_1712,N_29553,N_29745);
and UO_1713 (O_1713,N_29908,N_29436);
and UO_1714 (O_1714,N_29574,N_29412);
and UO_1715 (O_1715,N_29878,N_29485);
or UO_1716 (O_1716,N_29738,N_29413);
or UO_1717 (O_1717,N_29556,N_29874);
nand UO_1718 (O_1718,N_29985,N_29846);
xnor UO_1719 (O_1719,N_29838,N_29663);
nand UO_1720 (O_1720,N_29660,N_29933);
xor UO_1721 (O_1721,N_29403,N_29440);
xnor UO_1722 (O_1722,N_29437,N_29800);
nand UO_1723 (O_1723,N_29963,N_29679);
nor UO_1724 (O_1724,N_29921,N_29744);
and UO_1725 (O_1725,N_29467,N_29903);
or UO_1726 (O_1726,N_29566,N_29791);
or UO_1727 (O_1727,N_29930,N_29717);
nor UO_1728 (O_1728,N_29676,N_29769);
or UO_1729 (O_1729,N_29648,N_29891);
and UO_1730 (O_1730,N_29691,N_29716);
nor UO_1731 (O_1731,N_29884,N_29579);
nor UO_1732 (O_1732,N_29978,N_29890);
and UO_1733 (O_1733,N_29774,N_29754);
nor UO_1734 (O_1734,N_29666,N_29585);
xnor UO_1735 (O_1735,N_29696,N_29573);
nand UO_1736 (O_1736,N_29474,N_29799);
and UO_1737 (O_1737,N_29724,N_29872);
nand UO_1738 (O_1738,N_29740,N_29956);
or UO_1739 (O_1739,N_29948,N_29849);
nor UO_1740 (O_1740,N_29629,N_29727);
nor UO_1741 (O_1741,N_29766,N_29761);
nor UO_1742 (O_1742,N_29834,N_29810);
nor UO_1743 (O_1743,N_29598,N_29979);
nor UO_1744 (O_1744,N_29650,N_29757);
or UO_1745 (O_1745,N_29936,N_29951);
xnor UO_1746 (O_1746,N_29636,N_29565);
nor UO_1747 (O_1747,N_29870,N_29747);
and UO_1748 (O_1748,N_29470,N_29415);
and UO_1749 (O_1749,N_29729,N_29993);
nor UO_1750 (O_1750,N_29598,N_29949);
nor UO_1751 (O_1751,N_29427,N_29887);
nand UO_1752 (O_1752,N_29603,N_29631);
and UO_1753 (O_1753,N_29948,N_29863);
xnor UO_1754 (O_1754,N_29532,N_29540);
and UO_1755 (O_1755,N_29714,N_29821);
or UO_1756 (O_1756,N_29622,N_29648);
nor UO_1757 (O_1757,N_29710,N_29712);
nand UO_1758 (O_1758,N_29728,N_29873);
nor UO_1759 (O_1759,N_29492,N_29962);
xor UO_1760 (O_1760,N_29411,N_29960);
and UO_1761 (O_1761,N_29989,N_29717);
and UO_1762 (O_1762,N_29734,N_29411);
and UO_1763 (O_1763,N_29633,N_29571);
and UO_1764 (O_1764,N_29435,N_29520);
xnor UO_1765 (O_1765,N_29955,N_29431);
nand UO_1766 (O_1766,N_29671,N_29963);
nor UO_1767 (O_1767,N_29427,N_29416);
nor UO_1768 (O_1768,N_29957,N_29795);
or UO_1769 (O_1769,N_29867,N_29725);
nand UO_1770 (O_1770,N_29925,N_29550);
nand UO_1771 (O_1771,N_29742,N_29740);
xor UO_1772 (O_1772,N_29653,N_29625);
nor UO_1773 (O_1773,N_29498,N_29893);
and UO_1774 (O_1774,N_29984,N_29937);
and UO_1775 (O_1775,N_29668,N_29890);
or UO_1776 (O_1776,N_29559,N_29979);
or UO_1777 (O_1777,N_29815,N_29630);
and UO_1778 (O_1778,N_29927,N_29834);
nand UO_1779 (O_1779,N_29419,N_29626);
nor UO_1780 (O_1780,N_29617,N_29540);
or UO_1781 (O_1781,N_29656,N_29585);
nand UO_1782 (O_1782,N_29428,N_29557);
xnor UO_1783 (O_1783,N_29712,N_29843);
xor UO_1784 (O_1784,N_29935,N_29807);
nand UO_1785 (O_1785,N_29706,N_29944);
nor UO_1786 (O_1786,N_29789,N_29807);
nor UO_1787 (O_1787,N_29998,N_29764);
nand UO_1788 (O_1788,N_29800,N_29629);
nor UO_1789 (O_1789,N_29525,N_29510);
nor UO_1790 (O_1790,N_29424,N_29911);
and UO_1791 (O_1791,N_29983,N_29442);
or UO_1792 (O_1792,N_29927,N_29583);
nor UO_1793 (O_1793,N_29506,N_29846);
nand UO_1794 (O_1794,N_29770,N_29805);
or UO_1795 (O_1795,N_29776,N_29995);
xnor UO_1796 (O_1796,N_29499,N_29470);
or UO_1797 (O_1797,N_29719,N_29484);
nor UO_1798 (O_1798,N_29826,N_29670);
nand UO_1799 (O_1799,N_29826,N_29908);
and UO_1800 (O_1800,N_29462,N_29467);
and UO_1801 (O_1801,N_29687,N_29409);
and UO_1802 (O_1802,N_29491,N_29556);
or UO_1803 (O_1803,N_29597,N_29803);
xor UO_1804 (O_1804,N_29551,N_29724);
and UO_1805 (O_1805,N_29581,N_29763);
nor UO_1806 (O_1806,N_29821,N_29739);
nor UO_1807 (O_1807,N_29585,N_29958);
and UO_1808 (O_1808,N_29608,N_29996);
xnor UO_1809 (O_1809,N_29437,N_29934);
and UO_1810 (O_1810,N_29826,N_29825);
and UO_1811 (O_1811,N_29926,N_29589);
and UO_1812 (O_1812,N_29449,N_29644);
xor UO_1813 (O_1813,N_29428,N_29805);
nor UO_1814 (O_1814,N_29797,N_29918);
and UO_1815 (O_1815,N_29413,N_29452);
xor UO_1816 (O_1816,N_29882,N_29859);
and UO_1817 (O_1817,N_29421,N_29912);
or UO_1818 (O_1818,N_29916,N_29455);
nand UO_1819 (O_1819,N_29494,N_29456);
nand UO_1820 (O_1820,N_29520,N_29577);
and UO_1821 (O_1821,N_29551,N_29822);
nand UO_1822 (O_1822,N_29860,N_29551);
xor UO_1823 (O_1823,N_29766,N_29616);
or UO_1824 (O_1824,N_29439,N_29835);
xor UO_1825 (O_1825,N_29735,N_29447);
or UO_1826 (O_1826,N_29931,N_29784);
or UO_1827 (O_1827,N_29906,N_29824);
nor UO_1828 (O_1828,N_29980,N_29474);
and UO_1829 (O_1829,N_29637,N_29621);
nor UO_1830 (O_1830,N_29907,N_29524);
or UO_1831 (O_1831,N_29657,N_29816);
nor UO_1832 (O_1832,N_29488,N_29926);
xor UO_1833 (O_1833,N_29585,N_29838);
nor UO_1834 (O_1834,N_29792,N_29590);
xor UO_1835 (O_1835,N_29799,N_29889);
xnor UO_1836 (O_1836,N_29669,N_29761);
xor UO_1837 (O_1837,N_29957,N_29811);
and UO_1838 (O_1838,N_29433,N_29805);
nand UO_1839 (O_1839,N_29663,N_29808);
xor UO_1840 (O_1840,N_29638,N_29929);
nand UO_1841 (O_1841,N_29452,N_29623);
or UO_1842 (O_1842,N_29524,N_29690);
xor UO_1843 (O_1843,N_29961,N_29747);
nand UO_1844 (O_1844,N_29493,N_29400);
and UO_1845 (O_1845,N_29732,N_29820);
or UO_1846 (O_1846,N_29645,N_29724);
nor UO_1847 (O_1847,N_29807,N_29743);
and UO_1848 (O_1848,N_29463,N_29773);
xnor UO_1849 (O_1849,N_29807,N_29430);
nand UO_1850 (O_1850,N_29725,N_29955);
or UO_1851 (O_1851,N_29579,N_29434);
nand UO_1852 (O_1852,N_29807,N_29462);
or UO_1853 (O_1853,N_29902,N_29938);
nand UO_1854 (O_1854,N_29503,N_29509);
xnor UO_1855 (O_1855,N_29655,N_29874);
xor UO_1856 (O_1856,N_29700,N_29695);
or UO_1857 (O_1857,N_29610,N_29700);
nor UO_1858 (O_1858,N_29598,N_29694);
nand UO_1859 (O_1859,N_29523,N_29440);
nand UO_1860 (O_1860,N_29463,N_29868);
nand UO_1861 (O_1861,N_29723,N_29604);
xor UO_1862 (O_1862,N_29991,N_29614);
nor UO_1863 (O_1863,N_29931,N_29990);
and UO_1864 (O_1864,N_29996,N_29776);
nor UO_1865 (O_1865,N_29416,N_29934);
nand UO_1866 (O_1866,N_29980,N_29736);
and UO_1867 (O_1867,N_29681,N_29696);
or UO_1868 (O_1868,N_29607,N_29957);
nor UO_1869 (O_1869,N_29773,N_29545);
nor UO_1870 (O_1870,N_29878,N_29927);
and UO_1871 (O_1871,N_29774,N_29448);
xor UO_1872 (O_1872,N_29813,N_29779);
and UO_1873 (O_1873,N_29837,N_29772);
nor UO_1874 (O_1874,N_29652,N_29644);
nor UO_1875 (O_1875,N_29878,N_29774);
nand UO_1876 (O_1876,N_29431,N_29726);
nor UO_1877 (O_1877,N_29494,N_29507);
xor UO_1878 (O_1878,N_29806,N_29743);
or UO_1879 (O_1879,N_29719,N_29464);
nor UO_1880 (O_1880,N_29455,N_29679);
or UO_1881 (O_1881,N_29760,N_29873);
nand UO_1882 (O_1882,N_29967,N_29519);
and UO_1883 (O_1883,N_29943,N_29920);
nor UO_1884 (O_1884,N_29702,N_29876);
xor UO_1885 (O_1885,N_29803,N_29679);
or UO_1886 (O_1886,N_29715,N_29463);
nand UO_1887 (O_1887,N_29937,N_29423);
nand UO_1888 (O_1888,N_29928,N_29631);
and UO_1889 (O_1889,N_29736,N_29983);
nor UO_1890 (O_1890,N_29867,N_29886);
nor UO_1891 (O_1891,N_29695,N_29973);
nor UO_1892 (O_1892,N_29536,N_29573);
and UO_1893 (O_1893,N_29665,N_29864);
xnor UO_1894 (O_1894,N_29638,N_29485);
nor UO_1895 (O_1895,N_29749,N_29547);
and UO_1896 (O_1896,N_29706,N_29947);
nand UO_1897 (O_1897,N_29603,N_29766);
and UO_1898 (O_1898,N_29845,N_29781);
and UO_1899 (O_1899,N_29960,N_29708);
and UO_1900 (O_1900,N_29516,N_29510);
xnor UO_1901 (O_1901,N_29543,N_29619);
nand UO_1902 (O_1902,N_29589,N_29929);
or UO_1903 (O_1903,N_29981,N_29921);
nor UO_1904 (O_1904,N_29428,N_29561);
nand UO_1905 (O_1905,N_29983,N_29786);
nand UO_1906 (O_1906,N_29942,N_29815);
xnor UO_1907 (O_1907,N_29460,N_29924);
xor UO_1908 (O_1908,N_29405,N_29443);
nor UO_1909 (O_1909,N_29725,N_29595);
xnor UO_1910 (O_1910,N_29438,N_29653);
and UO_1911 (O_1911,N_29756,N_29642);
nor UO_1912 (O_1912,N_29814,N_29755);
and UO_1913 (O_1913,N_29502,N_29977);
nor UO_1914 (O_1914,N_29634,N_29884);
or UO_1915 (O_1915,N_29731,N_29864);
nand UO_1916 (O_1916,N_29500,N_29973);
or UO_1917 (O_1917,N_29557,N_29907);
nor UO_1918 (O_1918,N_29971,N_29484);
or UO_1919 (O_1919,N_29550,N_29447);
and UO_1920 (O_1920,N_29621,N_29524);
nand UO_1921 (O_1921,N_29463,N_29913);
nand UO_1922 (O_1922,N_29812,N_29736);
xor UO_1923 (O_1923,N_29680,N_29448);
and UO_1924 (O_1924,N_29659,N_29834);
nor UO_1925 (O_1925,N_29609,N_29728);
nand UO_1926 (O_1926,N_29416,N_29670);
nand UO_1927 (O_1927,N_29981,N_29982);
and UO_1928 (O_1928,N_29578,N_29526);
xnor UO_1929 (O_1929,N_29772,N_29608);
or UO_1930 (O_1930,N_29442,N_29704);
nand UO_1931 (O_1931,N_29685,N_29729);
nor UO_1932 (O_1932,N_29946,N_29571);
or UO_1933 (O_1933,N_29892,N_29641);
nand UO_1934 (O_1934,N_29589,N_29872);
xor UO_1935 (O_1935,N_29731,N_29902);
and UO_1936 (O_1936,N_29997,N_29831);
nor UO_1937 (O_1937,N_29714,N_29532);
and UO_1938 (O_1938,N_29771,N_29541);
nor UO_1939 (O_1939,N_29832,N_29731);
and UO_1940 (O_1940,N_29544,N_29590);
or UO_1941 (O_1941,N_29890,N_29681);
and UO_1942 (O_1942,N_29430,N_29641);
nor UO_1943 (O_1943,N_29491,N_29924);
nand UO_1944 (O_1944,N_29694,N_29548);
or UO_1945 (O_1945,N_29642,N_29904);
nand UO_1946 (O_1946,N_29838,N_29923);
xnor UO_1947 (O_1947,N_29422,N_29459);
or UO_1948 (O_1948,N_29571,N_29993);
and UO_1949 (O_1949,N_29998,N_29441);
nand UO_1950 (O_1950,N_29900,N_29591);
xor UO_1951 (O_1951,N_29879,N_29754);
or UO_1952 (O_1952,N_29585,N_29804);
nor UO_1953 (O_1953,N_29761,N_29521);
nor UO_1954 (O_1954,N_29427,N_29614);
and UO_1955 (O_1955,N_29862,N_29865);
nor UO_1956 (O_1956,N_29768,N_29756);
or UO_1957 (O_1957,N_29609,N_29491);
and UO_1958 (O_1958,N_29795,N_29467);
xor UO_1959 (O_1959,N_29726,N_29871);
or UO_1960 (O_1960,N_29578,N_29890);
and UO_1961 (O_1961,N_29612,N_29854);
or UO_1962 (O_1962,N_29623,N_29559);
nor UO_1963 (O_1963,N_29678,N_29990);
or UO_1964 (O_1964,N_29444,N_29471);
and UO_1965 (O_1965,N_29633,N_29812);
or UO_1966 (O_1966,N_29862,N_29481);
nor UO_1967 (O_1967,N_29836,N_29833);
xor UO_1968 (O_1968,N_29886,N_29701);
xnor UO_1969 (O_1969,N_29721,N_29824);
xor UO_1970 (O_1970,N_29821,N_29803);
or UO_1971 (O_1971,N_29596,N_29565);
nand UO_1972 (O_1972,N_29615,N_29454);
xnor UO_1973 (O_1973,N_29587,N_29889);
and UO_1974 (O_1974,N_29740,N_29567);
and UO_1975 (O_1975,N_29467,N_29878);
xnor UO_1976 (O_1976,N_29536,N_29687);
nor UO_1977 (O_1977,N_29614,N_29997);
and UO_1978 (O_1978,N_29590,N_29463);
or UO_1979 (O_1979,N_29689,N_29754);
xnor UO_1980 (O_1980,N_29838,N_29646);
or UO_1981 (O_1981,N_29479,N_29823);
nand UO_1982 (O_1982,N_29541,N_29889);
or UO_1983 (O_1983,N_29742,N_29880);
nor UO_1984 (O_1984,N_29417,N_29687);
xor UO_1985 (O_1985,N_29596,N_29597);
xnor UO_1986 (O_1986,N_29897,N_29628);
nand UO_1987 (O_1987,N_29719,N_29873);
and UO_1988 (O_1988,N_29787,N_29969);
and UO_1989 (O_1989,N_29939,N_29618);
or UO_1990 (O_1990,N_29818,N_29463);
xor UO_1991 (O_1991,N_29724,N_29704);
xor UO_1992 (O_1992,N_29490,N_29770);
and UO_1993 (O_1993,N_29438,N_29961);
xnor UO_1994 (O_1994,N_29904,N_29865);
nor UO_1995 (O_1995,N_29888,N_29703);
nand UO_1996 (O_1996,N_29611,N_29715);
nand UO_1997 (O_1997,N_29682,N_29643);
and UO_1998 (O_1998,N_29845,N_29849);
xor UO_1999 (O_1999,N_29424,N_29498);
nor UO_2000 (O_2000,N_29742,N_29460);
or UO_2001 (O_2001,N_29614,N_29910);
nor UO_2002 (O_2002,N_29868,N_29523);
xor UO_2003 (O_2003,N_29842,N_29895);
nor UO_2004 (O_2004,N_29848,N_29502);
and UO_2005 (O_2005,N_29911,N_29839);
nand UO_2006 (O_2006,N_29546,N_29559);
and UO_2007 (O_2007,N_29529,N_29913);
and UO_2008 (O_2008,N_29542,N_29791);
xor UO_2009 (O_2009,N_29500,N_29896);
nor UO_2010 (O_2010,N_29488,N_29779);
xnor UO_2011 (O_2011,N_29966,N_29460);
or UO_2012 (O_2012,N_29428,N_29886);
xor UO_2013 (O_2013,N_29598,N_29954);
nor UO_2014 (O_2014,N_29459,N_29685);
or UO_2015 (O_2015,N_29514,N_29824);
xnor UO_2016 (O_2016,N_29683,N_29488);
or UO_2017 (O_2017,N_29412,N_29976);
xnor UO_2018 (O_2018,N_29932,N_29835);
and UO_2019 (O_2019,N_29567,N_29711);
and UO_2020 (O_2020,N_29692,N_29503);
or UO_2021 (O_2021,N_29458,N_29688);
xor UO_2022 (O_2022,N_29759,N_29504);
nor UO_2023 (O_2023,N_29927,N_29728);
or UO_2024 (O_2024,N_29860,N_29818);
nand UO_2025 (O_2025,N_29723,N_29736);
nand UO_2026 (O_2026,N_29730,N_29408);
or UO_2027 (O_2027,N_29752,N_29867);
xnor UO_2028 (O_2028,N_29831,N_29786);
nand UO_2029 (O_2029,N_29897,N_29640);
xor UO_2030 (O_2030,N_29879,N_29643);
nor UO_2031 (O_2031,N_29923,N_29719);
or UO_2032 (O_2032,N_29583,N_29889);
nand UO_2033 (O_2033,N_29473,N_29414);
nand UO_2034 (O_2034,N_29964,N_29580);
nor UO_2035 (O_2035,N_29934,N_29756);
and UO_2036 (O_2036,N_29485,N_29502);
xor UO_2037 (O_2037,N_29899,N_29933);
nand UO_2038 (O_2038,N_29403,N_29494);
or UO_2039 (O_2039,N_29505,N_29710);
nor UO_2040 (O_2040,N_29979,N_29760);
nor UO_2041 (O_2041,N_29974,N_29836);
and UO_2042 (O_2042,N_29871,N_29958);
nor UO_2043 (O_2043,N_29461,N_29464);
nor UO_2044 (O_2044,N_29400,N_29477);
nand UO_2045 (O_2045,N_29573,N_29798);
nor UO_2046 (O_2046,N_29506,N_29655);
nand UO_2047 (O_2047,N_29465,N_29421);
nand UO_2048 (O_2048,N_29423,N_29655);
or UO_2049 (O_2049,N_29639,N_29706);
nand UO_2050 (O_2050,N_29465,N_29666);
and UO_2051 (O_2051,N_29637,N_29403);
xnor UO_2052 (O_2052,N_29753,N_29781);
xor UO_2053 (O_2053,N_29908,N_29861);
nor UO_2054 (O_2054,N_29623,N_29581);
or UO_2055 (O_2055,N_29915,N_29675);
xnor UO_2056 (O_2056,N_29646,N_29516);
nand UO_2057 (O_2057,N_29739,N_29633);
nand UO_2058 (O_2058,N_29502,N_29828);
nand UO_2059 (O_2059,N_29461,N_29627);
xnor UO_2060 (O_2060,N_29878,N_29742);
nor UO_2061 (O_2061,N_29612,N_29643);
xor UO_2062 (O_2062,N_29697,N_29430);
xor UO_2063 (O_2063,N_29511,N_29619);
or UO_2064 (O_2064,N_29545,N_29857);
and UO_2065 (O_2065,N_29656,N_29917);
or UO_2066 (O_2066,N_29406,N_29400);
xnor UO_2067 (O_2067,N_29483,N_29487);
nand UO_2068 (O_2068,N_29817,N_29402);
or UO_2069 (O_2069,N_29842,N_29727);
and UO_2070 (O_2070,N_29555,N_29804);
nand UO_2071 (O_2071,N_29807,N_29470);
and UO_2072 (O_2072,N_29988,N_29891);
nand UO_2073 (O_2073,N_29606,N_29662);
nor UO_2074 (O_2074,N_29555,N_29410);
nor UO_2075 (O_2075,N_29528,N_29507);
nor UO_2076 (O_2076,N_29761,N_29584);
nand UO_2077 (O_2077,N_29528,N_29914);
nand UO_2078 (O_2078,N_29529,N_29560);
nor UO_2079 (O_2079,N_29754,N_29977);
and UO_2080 (O_2080,N_29728,N_29720);
xor UO_2081 (O_2081,N_29965,N_29545);
and UO_2082 (O_2082,N_29478,N_29613);
xor UO_2083 (O_2083,N_29853,N_29909);
and UO_2084 (O_2084,N_29843,N_29567);
nand UO_2085 (O_2085,N_29645,N_29508);
nor UO_2086 (O_2086,N_29787,N_29490);
and UO_2087 (O_2087,N_29469,N_29996);
xor UO_2088 (O_2088,N_29859,N_29648);
xnor UO_2089 (O_2089,N_29488,N_29532);
nor UO_2090 (O_2090,N_29426,N_29605);
nand UO_2091 (O_2091,N_29710,N_29959);
and UO_2092 (O_2092,N_29995,N_29848);
nor UO_2093 (O_2093,N_29673,N_29561);
nor UO_2094 (O_2094,N_29681,N_29952);
nor UO_2095 (O_2095,N_29681,N_29828);
xnor UO_2096 (O_2096,N_29777,N_29759);
xor UO_2097 (O_2097,N_29924,N_29405);
nand UO_2098 (O_2098,N_29863,N_29956);
nor UO_2099 (O_2099,N_29540,N_29976);
xor UO_2100 (O_2100,N_29956,N_29526);
or UO_2101 (O_2101,N_29788,N_29619);
nor UO_2102 (O_2102,N_29477,N_29999);
nor UO_2103 (O_2103,N_29801,N_29580);
nand UO_2104 (O_2104,N_29855,N_29906);
nor UO_2105 (O_2105,N_29778,N_29870);
nor UO_2106 (O_2106,N_29625,N_29745);
nand UO_2107 (O_2107,N_29411,N_29664);
or UO_2108 (O_2108,N_29620,N_29796);
nor UO_2109 (O_2109,N_29979,N_29482);
or UO_2110 (O_2110,N_29659,N_29713);
nor UO_2111 (O_2111,N_29536,N_29704);
or UO_2112 (O_2112,N_29624,N_29893);
nand UO_2113 (O_2113,N_29977,N_29989);
xor UO_2114 (O_2114,N_29792,N_29874);
nor UO_2115 (O_2115,N_29874,N_29523);
nor UO_2116 (O_2116,N_29727,N_29862);
or UO_2117 (O_2117,N_29451,N_29640);
and UO_2118 (O_2118,N_29723,N_29490);
xor UO_2119 (O_2119,N_29670,N_29682);
or UO_2120 (O_2120,N_29710,N_29932);
nand UO_2121 (O_2121,N_29726,N_29708);
nand UO_2122 (O_2122,N_29718,N_29875);
nand UO_2123 (O_2123,N_29588,N_29749);
nand UO_2124 (O_2124,N_29708,N_29572);
or UO_2125 (O_2125,N_29690,N_29978);
or UO_2126 (O_2126,N_29886,N_29919);
nor UO_2127 (O_2127,N_29968,N_29420);
and UO_2128 (O_2128,N_29835,N_29479);
or UO_2129 (O_2129,N_29420,N_29602);
or UO_2130 (O_2130,N_29892,N_29508);
nand UO_2131 (O_2131,N_29620,N_29457);
or UO_2132 (O_2132,N_29927,N_29450);
xor UO_2133 (O_2133,N_29933,N_29615);
nand UO_2134 (O_2134,N_29412,N_29962);
or UO_2135 (O_2135,N_29445,N_29698);
or UO_2136 (O_2136,N_29605,N_29693);
and UO_2137 (O_2137,N_29927,N_29509);
and UO_2138 (O_2138,N_29486,N_29828);
nand UO_2139 (O_2139,N_29804,N_29719);
nor UO_2140 (O_2140,N_29584,N_29957);
xnor UO_2141 (O_2141,N_29927,N_29757);
nand UO_2142 (O_2142,N_29876,N_29517);
and UO_2143 (O_2143,N_29664,N_29662);
and UO_2144 (O_2144,N_29498,N_29639);
and UO_2145 (O_2145,N_29977,N_29580);
nand UO_2146 (O_2146,N_29499,N_29724);
or UO_2147 (O_2147,N_29835,N_29559);
and UO_2148 (O_2148,N_29910,N_29919);
or UO_2149 (O_2149,N_29607,N_29928);
or UO_2150 (O_2150,N_29714,N_29661);
and UO_2151 (O_2151,N_29857,N_29894);
xnor UO_2152 (O_2152,N_29468,N_29639);
and UO_2153 (O_2153,N_29620,N_29941);
xor UO_2154 (O_2154,N_29863,N_29703);
xor UO_2155 (O_2155,N_29902,N_29738);
or UO_2156 (O_2156,N_29754,N_29875);
or UO_2157 (O_2157,N_29560,N_29766);
nor UO_2158 (O_2158,N_29957,N_29562);
nand UO_2159 (O_2159,N_29477,N_29879);
nor UO_2160 (O_2160,N_29753,N_29826);
or UO_2161 (O_2161,N_29434,N_29450);
xnor UO_2162 (O_2162,N_29934,N_29484);
nor UO_2163 (O_2163,N_29431,N_29927);
nand UO_2164 (O_2164,N_29932,N_29813);
xnor UO_2165 (O_2165,N_29871,N_29837);
and UO_2166 (O_2166,N_29855,N_29451);
nand UO_2167 (O_2167,N_29765,N_29450);
and UO_2168 (O_2168,N_29556,N_29454);
xnor UO_2169 (O_2169,N_29653,N_29576);
nand UO_2170 (O_2170,N_29602,N_29871);
nor UO_2171 (O_2171,N_29416,N_29943);
and UO_2172 (O_2172,N_29915,N_29474);
xnor UO_2173 (O_2173,N_29881,N_29667);
and UO_2174 (O_2174,N_29483,N_29823);
and UO_2175 (O_2175,N_29483,N_29708);
nor UO_2176 (O_2176,N_29974,N_29473);
and UO_2177 (O_2177,N_29626,N_29616);
nor UO_2178 (O_2178,N_29462,N_29444);
xnor UO_2179 (O_2179,N_29800,N_29806);
nand UO_2180 (O_2180,N_29643,N_29868);
nand UO_2181 (O_2181,N_29830,N_29891);
or UO_2182 (O_2182,N_29816,N_29476);
or UO_2183 (O_2183,N_29481,N_29863);
or UO_2184 (O_2184,N_29964,N_29717);
nand UO_2185 (O_2185,N_29897,N_29670);
and UO_2186 (O_2186,N_29741,N_29474);
nor UO_2187 (O_2187,N_29938,N_29709);
nor UO_2188 (O_2188,N_29851,N_29706);
nor UO_2189 (O_2189,N_29423,N_29469);
xnor UO_2190 (O_2190,N_29687,N_29601);
or UO_2191 (O_2191,N_29974,N_29965);
nand UO_2192 (O_2192,N_29901,N_29977);
nand UO_2193 (O_2193,N_29401,N_29849);
nand UO_2194 (O_2194,N_29823,N_29915);
or UO_2195 (O_2195,N_29779,N_29660);
and UO_2196 (O_2196,N_29910,N_29495);
xnor UO_2197 (O_2197,N_29815,N_29786);
nor UO_2198 (O_2198,N_29768,N_29739);
or UO_2199 (O_2199,N_29507,N_29449);
and UO_2200 (O_2200,N_29883,N_29707);
nor UO_2201 (O_2201,N_29973,N_29873);
and UO_2202 (O_2202,N_29810,N_29645);
nor UO_2203 (O_2203,N_29875,N_29751);
or UO_2204 (O_2204,N_29662,N_29502);
and UO_2205 (O_2205,N_29494,N_29948);
xor UO_2206 (O_2206,N_29578,N_29975);
nand UO_2207 (O_2207,N_29723,N_29444);
nor UO_2208 (O_2208,N_29437,N_29742);
and UO_2209 (O_2209,N_29461,N_29864);
and UO_2210 (O_2210,N_29842,N_29645);
nor UO_2211 (O_2211,N_29906,N_29966);
nand UO_2212 (O_2212,N_29644,N_29939);
or UO_2213 (O_2213,N_29461,N_29639);
or UO_2214 (O_2214,N_29909,N_29919);
xnor UO_2215 (O_2215,N_29506,N_29697);
xnor UO_2216 (O_2216,N_29496,N_29802);
nor UO_2217 (O_2217,N_29915,N_29669);
nand UO_2218 (O_2218,N_29893,N_29964);
and UO_2219 (O_2219,N_29681,N_29557);
or UO_2220 (O_2220,N_29947,N_29540);
nor UO_2221 (O_2221,N_29438,N_29755);
nand UO_2222 (O_2222,N_29897,N_29745);
and UO_2223 (O_2223,N_29624,N_29475);
nor UO_2224 (O_2224,N_29696,N_29997);
nor UO_2225 (O_2225,N_29860,N_29611);
nor UO_2226 (O_2226,N_29728,N_29703);
nand UO_2227 (O_2227,N_29967,N_29963);
or UO_2228 (O_2228,N_29812,N_29634);
nor UO_2229 (O_2229,N_29409,N_29647);
or UO_2230 (O_2230,N_29795,N_29505);
and UO_2231 (O_2231,N_29837,N_29902);
xnor UO_2232 (O_2232,N_29657,N_29687);
xor UO_2233 (O_2233,N_29983,N_29437);
and UO_2234 (O_2234,N_29671,N_29683);
nand UO_2235 (O_2235,N_29717,N_29439);
xor UO_2236 (O_2236,N_29440,N_29514);
and UO_2237 (O_2237,N_29728,N_29409);
or UO_2238 (O_2238,N_29582,N_29957);
nand UO_2239 (O_2239,N_29963,N_29932);
nand UO_2240 (O_2240,N_29505,N_29400);
nand UO_2241 (O_2241,N_29593,N_29817);
xor UO_2242 (O_2242,N_29418,N_29732);
xor UO_2243 (O_2243,N_29418,N_29969);
xor UO_2244 (O_2244,N_29449,N_29547);
xnor UO_2245 (O_2245,N_29992,N_29965);
or UO_2246 (O_2246,N_29614,N_29655);
xnor UO_2247 (O_2247,N_29523,N_29771);
or UO_2248 (O_2248,N_29527,N_29419);
or UO_2249 (O_2249,N_29846,N_29925);
and UO_2250 (O_2250,N_29960,N_29741);
nor UO_2251 (O_2251,N_29677,N_29903);
nor UO_2252 (O_2252,N_29629,N_29713);
and UO_2253 (O_2253,N_29569,N_29630);
nand UO_2254 (O_2254,N_29589,N_29804);
nor UO_2255 (O_2255,N_29704,N_29956);
nor UO_2256 (O_2256,N_29553,N_29885);
and UO_2257 (O_2257,N_29515,N_29883);
xor UO_2258 (O_2258,N_29845,N_29861);
xor UO_2259 (O_2259,N_29406,N_29709);
nor UO_2260 (O_2260,N_29541,N_29436);
xnor UO_2261 (O_2261,N_29508,N_29601);
xnor UO_2262 (O_2262,N_29655,N_29446);
nor UO_2263 (O_2263,N_29565,N_29674);
nand UO_2264 (O_2264,N_29601,N_29910);
xor UO_2265 (O_2265,N_29545,N_29578);
nor UO_2266 (O_2266,N_29890,N_29903);
or UO_2267 (O_2267,N_29516,N_29605);
nor UO_2268 (O_2268,N_29675,N_29931);
nand UO_2269 (O_2269,N_29824,N_29472);
and UO_2270 (O_2270,N_29439,N_29634);
or UO_2271 (O_2271,N_29911,N_29595);
nor UO_2272 (O_2272,N_29559,N_29603);
nor UO_2273 (O_2273,N_29533,N_29661);
xor UO_2274 (O_2274,N_29723,N_29638);
xnor UO_2275 (O_2275,N_29793,N_29584);
xnor UO_2276 (O_2276,N_29864,N_29529);
nor UO_2277 (O_2277,N_29803,N_29891);
or UO_2278 (O_2278,N_29526,N_29742);
or UO_2279 (O_2279,N_29837,N_29840);
nor UO_2280 (O_2280,N_29829,N_29571);
nand UO_2281 (O_2281,N_29577,N_29513);
and UO_2282 (O_2282,N_29955,N_29600);
xnor UO_2283 (O_2283,N_29482,N_29778);
xnor UO_2284 (O_2284,N_29791,N_29675);
and UO_2285 (O_2285,N_29898,N_29944);
and UO_2286 (O_2286,N_29611,N_29549);
xor UO_2287 (O_2287,N_29785,N_29775);
or UO_2288 (O_2288,N_29563,N_29741);
and UO_2289 (O_2289,N_29652,N_29781);
and UO_2290 (O_2290,N_29795,N_29551);
or UO_2291 (O_2291,N_29502,N_29703);
nor UO_2292 (O_2292,N_29721,N_29745);
or UO_2293 (O_2293,N_29776,N_29993);
and UO_2294 (O_2294,N_29871,N_29710);
nand UO_2295 (O_2295,N_29687,N_29654);
and UO_2296 (O_2296,N_29466,N_29881);
or UO_2297 (O_2297,N_29531,N_29596);
or UO_2298 (O_2298,N_29790,N_29659);
nand UO_2299 (O_2299,N_29523,N_29590);
xor UO_2300 (O_2300,N_29419,N_29587);
and UO_2301 (O_2301,N_29590,N_29763);
and UO_2302 (O_2302,N_29466,N_29764);
nor UO_2303 (O_2303,N_29447,N_29471);
xor UO_2304 (O_2304,N_29571,N_29550);
xnor UO_2305 (O_2305,N_29436,N_29964);
nor UO_2306 (O_2306,N_29579,N_29597);
or UO_2307 (O_2307,N_29721,N_29514);
xnor UO_2308 (O_2308,N_29677,N_29445);
and UO_2309 (O_2309,N_29917,N_29673);
xor UO_2310 (O_2310,N_29513,N_29499);
nand UO_2311 (O_2311,N_29418,N_29463);
or UO_2312 (O_2312,N_29624,N_29428);
or UO_2313 (O_2313,N_29834,N_29703);
nand UO_2314 (O_2314,N_29547,N_29565);
and UO_2315 (O_2315,N_29634,N_29591);
and UO_2316 (O_2316,N_29479,N_29724);
nor UO_2317 (O_2317,N_29845,N_29455);
and UO_2318 (O_2318,N_29589,N_29717);
xor UO_2319 (O_2319,N_29983,N_29925);
xnor UO_2320 (O_2320,N_29591,N_29809);
or UO_2321 (O_2321,N_29583,N_29414);
nand UO_2322 (O_2322,N_29661,N_29850);
nand UO_2323 (O_2323,N_29536,N_29602);
nor UO_2324 (O_2324,N_29727,N_29459);
or UO_2325 (O_2325,N_29977,N_29464);
xor UO_2326 (O_2326,N_29850,N_29703);
or UO_2327 (O_2327,N_29641,N_29667);
or UO_2328 (O_2328,N_29596,N_29861);
nor UO_2329 (O_2329,N_29861,N_29865);
nor UO_2330 (O_2330,N_29655,N_29660);
and UO_2331 (O_2331,N_29712,N_29511);
and UO_2332 (O_2332,N_29894,N_29575);
nand UO_2333 (O_2333,N_29506,N_29918);
and UO_2334 (O_2334,N_29485,N_29814);
nor UO_2335 (O_2335,N_29947,N_29414);
xnor UO_2336 (O_2336,N_29827,N_29869);
nand UO_2337 (O_2337,N_29941,N_29912);
nor UO_2338 (O_2338,N_29439,N_29446);
nand UO_2339 (O_2339,N_29585,N_29639);
and UO_2340 (O_2340,N_29807,N_29719);
xnor UO_2341 (O_2341,N_29593,N_29582);
nor UO_2342 (O_2342,N_29683,N_29739);
or UO_2343 (O_2343,N_29411,N_29939);
nor UO_2344 (O_2344,N_29831,N_29790);
and UO_2345 (O_2345,N_29457,N_29934);
and UO_2346 (O_2346,N_29701,N_29717);
or UO_2347 (O_2347,N_29736,N_29860);
nand UO_2348 (O_2348,N_29646,N_29562);
or UO_2349 (O_2349,N_29968,N_29823);
nand UO_2350 (O_2350,N_29750,N_29522);
and UO_2351 (O_2351,N_29438,N_29628);
nand UO_2352 (O_2352,N_29905,N_29574);
nor UO_2353 (O_2353,N_29478,N_29406);
nand UO_2354 (O_2354,N_29580,N_29873);
and UO_2355 (O_2355,N_29517,N_29615);
or UO_2356 (O_2356,N_29518,N_29856);
nor UO_2357 (O_2357,N_29781,N_29928);
nand UO_2358 (O_2358,N_29582,N_29552);
nor UO_2359 (O_2359,N_29512,N_29424);
or UO_2360 (O_2360,N_29642,N_29704);
nor UO_2361 (O_2361,N_29770,N_29800);
or UO_2362 (O_2362,N_29494,N_29523);
and UO_2363 (O_2363,N_29487,N_29610);
nor UO_2364 (O_2364,N_29405,N_29474);
nand UO_2365 (O_2365,N_29950,N_29918);
or UO_2366 (O_2366,N_29720,N_29673);
xor UO_2367 (O_2367,N_29697,N_29775);
xor UO_2368 (O_2368,N_29588,N_29493);
nand UO_2369 (O_2369,N_29568,N_29418);
xnor UO_2370 (O_2370,N_29539,N_29632);
or UO_2371 (O_2371,N_29516,N_29515);
xor UO_2372 (O_2372,N_29863,N_29940);
nand UO_2373 (O_2373,N_29910,N_29515);
and UO_2374 (O_2374,N_29465,N_29897);
nor UO_2375 (O_2375,N_29902,N_29570);
xnor UO_2376 (O_2376,N_29919,N_29971);
nor UO_2377 (O_2377,N_29658,N_29714);
nor UO_2378 (O_2378,N_29791,N_29594);
xnor UO_2379 (O_2379,N_29589,N_29874);
or UO_2380 (O_2380,N_29795,N_29911);
xnor UO_2381 (O_2381,N_29601,N_29602);
xor UO_2382 (O_2382,N_29655,N_29889);
nand UO_2383 (O_2383,N_29949,N_29798);
nor UO_2384 (O_2384,N_29466,N_29826);
or UO_2385 (O_2385,N_29805,N_29616);
nand UO_2386 (O_2386,N_29631,N_29830);
and UO_2387 (O_2387,N_29620,N_29486);
and UO_2388 (O_2388,N_29879,N_29430);
or UO_2389 (O_2389,N_29673,N_29918);
nor UO_2390 (O_2390,N_29436,N_29996);
and UO_2391 (O_2391,N_29967,N_29925);
xor UO_2392 (O_2392,N_29945,N_29886);
nand UO_2393 (O_2393,N_29592,N_29640);
or UO_2394 (O_2394,N_29426,N_29620);
or UO_2395 (O_2395,N_29968,N_29493);
and UO_2396 (O_2396,N_29448,N_29800);
nor UO_2397 (O_2397,N_29783,N_29649);
or UO_2398 (O_2398,N_29740,N_29728);
or UO_2399 (O_2399,N_29838,N_29778);
xnor UO_2400 (O_2400,N_29682,N_29970);
and UO_2401 (O_2401,N_29735,N_29905);
nor UO_2402 (O_2402,N_29830,N_29644);
and UO_2403 (O_2403,N_29537,N_29544);
nor UO_2404 (O_2404,N_29919,N_29699);
xnor UO_2405 (O_2405,N_29557,N_29668);
nor UO_2406 (O_2406,N_29999,N_29731);
nor UO_2407 (O_2407,N_29908,N_29893);
and UO_2408 (O_2408,N_29703,N_29451);
or UO_2409 (O_2409,N_29687,N_29656);
nand UO_2410 (O_2410,N_29652,N_29645);
nor UO_2411 (O_2411,N_29804,N_29916);
nand UO_2412 (O_2412,N_29579,N_29590);
and UO_2413 (O_2413,N_29553,N_29542);
nor UO_2414 (O_2414,N_29562,N_29506);
or UO_2415 (O_2415,N_29753,N_29995);
and UO_2416 (O_2416,N_29606,N_29936);
nand UO_2417 (O_2417,N_29674,N_29776);
and UO_2418 (O_2418,N_29792,N_29803);
or UO_2419 (O_2419,N_29495,N_29967);
and UO_2420 (O_2420,N_29882,N_29785);
nand UO_2421 (O_2421,N_29905,N_29737);
and UO_2422 (O_2422,N_29630,N_29438);
nand UO_2423 (O_2423,N_29454,N_29604);
or UO_2424 (O_2424,N_29573,N_29590);
nand UO_2425 (O_2425,N_29620,N_29557);
and UO_2426 (O_2426,N_29897,N_29982);
xor UO_2427 (O_2427,N_29873,N_29995);
nand UO_2428 (O_2428,N_29922,N_29472);
xor UO_2429 (O_2429,N_29887,N_29569);
and UO_2430 (O_2430,N_29657,N_29720);
and UO_2431 (O_2431,N_29881,N_29807);
xnor UO_2432 (O_2432,N_29910,N_29762);
and UO_2433 (O_2433,N_29572,N_29939);
and UO_2434 (O_2434,N_29863,N_29898);
xnor UO_2435 (O_2435,N_29973,N_29759);
and UO_2436 (O_2436,N_29666,N_29997);
and UO_2437 (O_2437,N_29680,N_29541);
nor UO_2438 (O_2438,N_29477,N_29467);
and UO_2439 (O_2439,N_29768,N_29931);
or UO_2440 (O_2440,N_29878,N_29968);
and UO_2441 (O_2441,N_29605,N_29893);
nor UO_2442 (O_2442,N_29470,N_29862);
and UO_2443 (O_2443,N_29457,N_29481);
or UO_2444 (O_2444,N_29489,N_29987);
nor UO_2445 (O_2445,N_29854,N_29402);
nand UO_2446 (O_2446,N_29928,N_29582);
nand UO_2447 (O_2447,N_29520,N_29632);
nand UO_2448 (O_2448,N_29420,N_29642);
and UO_2449 (O_2449,N_29753,N_29829);
nor UO_2450 (O_2450,N_29900,N_29431);
nor UO_2451 (O_2451,N_29729,N_29949);
or UO_2452 (O_2452,N_29928,N_29469);
nor UO_2453 (O_2453,N_29552,N_29414);
nor UO_2454 (O_2454,N_29420,N_29515);
nor UO_2455 (O_2455,N_29595,N_29981);
xnor UO_2456 (O_2456,N_29435,N_29759);
and UO_2457 (O_2457,N_29483,N_29424);
and UO_2458 (O_2458,N_29846,N_29920);
and UO_2459 (O_2459,N_29611,N_29683);
or UO_2460 (O_2460,N_29735,N_29567);
xnor UO_2461 (O_2461,N_29405,N_29983);
nor UO_2462 (O_2462,N_29424,N_29676);
or UO_2463 (O_2463,N_29619,N_29930);
or UO_2464 (O_2464,N_29457,N_29890);
or UO_2465 (O_2465,N_29583,N_29531);
and UO_2466 (O_2466,N_29914,N_29662);
xnor UO_2467 (O_2467,N_29865,N_29724);
and UO_2468 (O_2468,N_29867,N_29506);
and UO_2469 (O_2469,N_29990,N_29754);
and UO_2470 (O_2470,N_29406,N_29426);
and UO_2471 (O_2471,N_29930,N_29977);
xor UO_2472 (O_2472,N_29771,N_29776);
nor UO_2473 (O_2473,N_29937,N_29572);
nand UO_2474 (O_2474,N_29907,N_29402);
nand UO_2475 (O_2475,N_29627,N_29851);
xor UO_2476 (O_2476,N_29761,N_29975);
nor UO_2477 (O_2477,N_29986,N_29994);
nor UO_2478 (O_2478,N_29620,N_29447);
and UO_2479 (O_2479,N_29825,N_29578);
xnor UO_2480 (O_2480,N_29980,N_29437);
nand UO_2481 (O_2481,N_29963,N_29616);
or UO_2482 (O_2482,N_29711,N_29686);
nand UO_2483 (O_2483,N_29827,N_29455);
nand UO_2484 (O_2484,N_29757,N_29954);
and UO_2485 (O_2485,N_29815,N_29923);
nor UO_2486 (O_2486,N_29694,N_29629);
or UO_2487 (O_2487,N_29773,N_29449);
nand UO_2488 (O_2488,N_29963,N_29599);
xor UO_2489 (O_2489,N_29520,N_29953);
nand UO_2490 (O_2490,N_29979,N_29929);
or UO_2491 (O_2491,N_29821,N_29751);
xnor UO_2492 (O_2492,N_29873,N_29821);
nand UO_2493 (O_2493,N_29908,N_29788);
nand UO_2494 (O_2494,N_29411,N_29529);
and UO_2495 (O_2495,N_29656,N_29619);
or UO_2496 (O_2496,N_29468,N_29644);
or UO_2497 (O_2497,N_29659,N_29773);
or UO_2498 (O_2498,N_29831,N_29866);
or UO_2499 (O_2499,N_29783,N_29874);
nor UO_2500 (O_2500,N_29608,N_29954);
nand UO_2501 (O_2501,N_29552,N_29491);
xor UO_2502 (O_2502,N_29586,N_29933);
and UO_2503 (O_2503,N_29686,N_29901);
nor UO_2504 (O_2504,N_29583,N_29856);
nand UO_2505 (O_2505,N_29891,N_29994);
xor UO_2506 (O_2506,N_29602,N_29951);
xnor UO_2507 (O_2507,N_29682,N_29968);
xnor UO_2508 (O_2508,N_29907,N_29805);
xnor UO_2509 (O_2509,N_29523,N_29768);
and UO_2510 (O_2510,N_29954,N_29434);
and UO_2511 (O_2511,N_29770,N_29543);
xor UO_2512 (O_2512,N_29572,N_29776);
and UO_2513 (O_2513,N_29848,N_29471);
xor UO_2514 (O_2514,N_29436,N_29770);
or UO_2515 (O_2515,N_29547,N_29745);
nand UO_2516 (O_2516,N_29875,N_29777);
or UO_2517 (O_2517,N_29747,N_29885);
nand UO_2518 (O_2518,N_29923,N_29795);
nor UO_2519 (O_2519,N_29499,N_29531);
nor UO_2520 (O_2520,N_29791,N_29913);
and UO_2521 (O_2521,N_29784,N_29976);
xor UO_2522 (O_2522,N_29694,N_29599);
nor UO_2523 (O_2523,N_29525,N_29977);
nor UO_2524 (O_2524,N_29820,N_29548);
nand UO_2525 (O_2525,N_29936,N_29499);
nand UO_2526 (O_2526,N_29978,N_29833);
nor UO_2527 (O_2527,N_29813,N_29545);
xnor UO_2528 (O_2528,N_29506,N_29430);
nand UO_2529 (O_2529,N_29436,N_29923);
nand UO_2530 (O_2530,N_29512,N_29683);
or UO_2531 (O_2531,N_29707,N_29492);
or UO_2532 (O_2532,N_29847,N_29537);
or UO_2533 (O_2533,N_29485,N_29415);
or UO_2534 (O_2534,N_29703,N_29407);
and UO_2535 (O_2535,N_29934,N_29935);
xor UO_2536 (O_2536,N_29622,N_29754);
and UO_2537 (O_2537,N_29842,N_29427);
nor UO_2538 (O_2538,N_29530,N_29747);
nor UO_2539 (O_2539,N_29740,N_29431);
and UO_2540 (O_2540,N_29582,N_29470);
nand UO_2541 (O_2541,N_29813,N_29850);
xor UO_2542 (O_2542,N_29983,N_29915);
or UO_2543 (O_2543,N_29662,N_29700);
or UO_2544 (O_2544,N_29551,N_29505);
nand UO_2545 (O_2545,N_29880,N_29563);
nor UO_2546 (O_2546,N_29773,N_29735);
or UO_2547 (O_2547,N_29425,N_29887);
nand UO_2548 (O_2548,N_29820,N_29978);
xor UO_2549 (O_2549,N_29590,N_29822);
and UO_2550 (O_2550,N_29400,N_29727);
and UO_2551 (O_2551,N_29867,N_29696);
or UO_2552 (O_2552,N_29550,N_29944);
nand UO_2553 (O_2553,N_29948,N_29810);
xor UO_2554 (O_2554,N_29613,N_29418);
nand UO_2555 (O_2555,N_29919,N_29756);
nor UO_2556 (O_2556,N_29706,N_29718);
xnor UO_2557 (O_2557,N_29780,N_29661);
nor UO_2558 (O_2558,N_29720,N_29828);
nor UO_2559 (O_2559,N_29931,N_29805);
nand UO_2560 (O_2560,N_29678,N_29903);
or UO_2561 (O_2561,N_29465,N_29874);
nand UO_2562 (O_2562,N_29723,N_29787);
nor UO_2563 (O_2563,N_29967,N_29504);
nand UO_2564 (O_2564,N_29586,N_29719);
xor UO_2565 (O_2565,N_29844,N_29548);
nand UO_2566 (O_2566,N_29534,N_29727);
nor UO_2567 (O_2567,N_29905,N_29786);
or UO_2568 (O_2568,N_29984,N_29448);
nor UO_2569 (O_2569,N_29424,N_29964);
and UO_2570 (O_2570,N_29817,N_29425);
nand UO_2571 (O_2571,N_29879,N_29500);
nor UO_2572 (O_2572,N_29497,N_29647);
nand UO_2573 (O_2573,N_29912,N_29786);
and UO_2574 (O_2574,N_29456,N_29780);
xnor UO_2575 (O_2575,N_29658,N_29495);
nand UO_2576 (O_2576,N_29844,N_29683);
nand UO_2577 (O_2577,N_29614,N_29973);
xnor UO_2578 (O_2578,N_29701,N_29944);
or UO_2579 (O_2579,N_29729,N_29568);
and UO_2580 (O_2580,N_29945,N_29470);
xor UO_2581 (O_2581,N_29605,N_29828);
or UO_2582 (O_2582,N_29835,N_29436);
nor UO_2583 (O_2583,N_29569,N_29860);
or UO_2584 (O_2584,N_29570,N_29453);
xnor UO_2585 (O_2585,N_29960,N_29523);
and UO_2586 (O_2586,N_29773,N_29895);
nand UO_2587 (O_2587,N_29586,N_29873);
nand UO_2588 (O_2588,N_29914,N_29656);
nand UO_2589 (O_2589,N_29793,N_29606);
and UO_2590 (O_2590,N_29818,N_29539);
nand UO_2591 (O_2591,N_29798,N_29637);
nand UO_2592 (O_2592,N_29766,N_29788);
or UO_2593 (O_2593,N_29904,N_29896);
xnor UO_2594 (O_2594,N_29620,N_29591);
xnor UO_2595 (O_2595,N_29612,N_29447);
and UO_2596 (O_2596,N_29916,N_29742);
xor UO_2597 (O_2597,N_29480,N_29815);
xnor UO_2598 (O_2598,N_29759,N_29884);
or UO_2599 (O_2599,N_29628,N_29957);
xnor UO_2600 (O_2600,N_29569,N_29787);
nand UO_2601 (O_2601,N_29939,N_29843);
or UO_2602 (O_2602,N_29518,N_29776);
nand UO_2603 (O_2603,N_29767,N_29433);
nor UO_2604 (O_2604,N_29883,N_29765);
or UO_2605 (O_2605,N_29556,N_29726);
or UO_2606 (O_2606,N_29722,N_29887);
nor UO_2607 (O_2607,N_29612,N_29498);
or UO_2608 (O_2608,N_29858,N_29778);
nand UO_2609 (O_2609,N_29761,N_29767);
and UO_2610 (O_2610,N_29471,N_29461);
and UO_2611 (O_2611,N_29866,N_29614);
or UO_2612 (O_2612,N_29429,N_29490);
and UO_2613 (O_2613,N_29508,N_29478);
nand UO_2614 (O_2614,N_29974,N_29568);
nor UO_2615 (O_2615,N_29425,N_29412);
and UO_2616 (O_2616,N_29948,N_29443);
nor UO_2617 (O_2617,N_29880,N_29754);
xnor UO_2618 (O_2618,N_29976,N_29545);
nand UO_2619 (O_2619,N_29931,N_29789);
nor UO_2620 (O_2620,N_29480,N_29983);
nand UO_2621 (O_2621,N_29480,N_29443);
xnor UO_2622 (O_2622,N_29538,N_29982);
nand UO_2623 (O_2623,N_29838,N_29952);
nor UO_2624 (O_2624,N_29408,N_29594);
or UO_2625 (O_2625,N_29440,N_29749);
xnor UO_2626 (O_2626,N_29733,N_29708);
xnor UO_2627 (O_2627,N_29659,N_29748);
nor UO_2628 (O_2628,N_29408,N_29947);
and UO_2629 (O_2629,N_29821,N_29695);
nand UO_2630 (O_2630,N_29837,N_29543);
nand UO_2631 (O_2631,N_29855,N_29429);
nor UO_2632 (O_2632,N_29997,N_29719);
and UO_2633 (O_2633,N_29515,N_29703);
or UO_2634 (O_2634,N_29600,N_29456);
nand UO_2635 (O_2635,N_29535,N_29791);
nand UO_2636 (O_2636,N_29981,N_29487);
xor UO_2637 (O_2637,N_29741,N_29783);
and UO_2638 (O_2638,N_29884,N_29858);
or UO_2639 (O_2639,N_29700,N_29517);
or UO_2640 (O_2640,N_29945,N_29819);
nor UO_2641 (O_2641,N_29645,N_29978);
and UO_2642 (O_2642,N_29651,N_29694);
nor UO_2643 (O_2643,N_29997,N_29411);
and UO_2644 (O_2644,N_29764,N_29755);
and UO_2645 (O_2645,N_29442,N_29894);
nand UO_2646 (O_2646,N_29483,N_29401);
or UO_2647 (O_2647,N_29969,N_29413);
nand UO_2648 (O_2648,N_29732,N_29546);
or UO_2649 (O_2649,N_29912,N_29716);
and UO_2650 (O_2650,N_29538,N_29806);
or UO_2651 (O_2651,N_29675,N_29540);
or UO_2652 (O_2652,N_29680,N_29728);
or UO_2653 (O_2653,N_29888,N_29854);
and UO_2654 (O_2654,N_29418,N_29788);
and UO_2655 (O_2655,N_29652,N_29959);
nand UO_2656 (O_2656,N_29511,N_29800);
or UO_2657 (O_2657,N_29896,N_29787);
and UO_2658 (O_2658,N_29535,N_29953);
and UO_2659 (O_2659,N_29932,N_29427);
nand UO_2660 (O_2660,N_29638,N_29927);
nor UO_2661 (O_2661,N_29932,N_29584);
xnor UO_2662 (O_2662,N_29986,N_29911);
and UO_2663 (O_2663,N_29761,N_29452);
nor UO_2664 (O_2664,N_29813,N_29790);
or UO_2665 (O_2665,N_29766,N_29430);
nand UO_2666 (O_2666,N_29465,N_29501);
xnor UO_2667 (O_2667,N_29839,N_29863);
xnor UO_2668 (O_2668,N_29627,N_29607);
or UO_2669 (O_2669,N_29916,N_29983);
nor UO_2670 (O_2670,N_29795,N_29869);
or UO_2671 (O_2671,N_29796,N_29856);
nand UO_2672 (O_2672,N_29501,N_29849);
nand UO_2673 (O_2673,N_29420,N_29848);
nor UO_2674 (O_2674,N_29710,N_29477);
and UO_2675 (O_2675,N_29671,N_29552);
or UO_2676 (O_2676,N_29654,N_29783);
nand UO_2677 (O_2677,N_29561,N_29844);
nand UO_2678 (O_2678,N_29445,N_29936);
xor UO_2679 (O_2679,N_29914,N_29758);
nand UO_2680 (O_2680,N_29725,N_29869);
xnor UO_2681 (O_2681,N_29460,N_29619);
nand UO_2682 (O_2682,N_29762,N_29916);
nor UO_2683 (O_2683,N_29991,N_29673);
nor UO_2684 (O_2684,N_29657,N_29659);
and UO_2685 (O_2685,N_29448,N_29999);
or UO_2686 (O_2686,N_29859,N_29875);
xnor UO_2687 (O_2687,N_29410,N_29994);
or UO_2688 (O_2688,N_29641,N_29899);
nand UO_2689 (O_2689,N_29613,N_29402);
and UO_2690 (O_2690,N_29827,N_29666);
or UO_2691 (O_2691,N_29967,N_29958);
nor UO_2692 (O_2692,N_29843,N_29959);
xor UO_2693 (O_2693,N_29435,N_29807);
xor UO_2694 (O_2694,N_29594,N_29406);
or UO_2695 (O_2695,N_29423,N_29493);
xnor UO_2696 (O_2696,N_29800,N_29719);
nand UO_2697 (O_2697,N_29941,N_29964);
nor UO_2698 (O_2698,N_29568,N_29749);
and UO_2699 (O_2699,N_29484,N_29581);
nor UO_2700 (O_2700,N_29493,N_29448);
nor UO_2701 (O_2701,N_29544,N_29547);
nand UO_2702 (O_2702,N_29457,N_29474);
or UO_2703 (O_2703,N_29520,N_29940);
and UO_2704 (O_2704,N_29979,N_29637);
nand UO_2705 (O_2705,N_29488,N_29574);
or UO_2706 (O_2706,N_29559,N_29810);
nor UO_2707 (O_2707,N_29921,N_29488);
xnor UO_2708 (O_2708,N_29642,N_29743);
or UO_2709 (O_2709,N_29583,N_29851);
nand UO_2710 (O_2710,N_29788,N_29824);
nand UO_2711 (O_2711,N_29890,N_29992);
or UO_2712 (O_2712,N_29663,N_29687);
nor UO_2713 (O_2713,N_29648,N_29719);
or UO_2714 (O_2714,N_29615,N_29731);
or UO_2715 (O_2715,N_29830,N_29780);
xor UO_2716 (O_2716,N_29509,N_29609);
and UO_2717 (O_2717,N_29969,N_29482);
nand UO_2718 (O_2718,N_29718,N_29638);
nand UO_2719 (O_2719,N_29633,N_29977);
or UO_2720 (O_2720,N_29831,N_29887);
and UO_2721 (O_2721,N_29797,N_29427);
nand UO_2722 (O_2722,N_29417,N_29888);
nand UO_2723 (O_2723,N_29945,N_29871);
xor UO_2724 (O_2724,N_29955,N_29901);
and UO_2725 (O_2725,N_29930,N_29934);
xor UO_2726 (O_2726,N_29713,N_29798);
and UO_2727 (O_2727,N_29575,N_29971);
nor UO_2728 (O_2728,N_29467,N_29517);
and UO_2729 (O_2729,N_29814,N_29859);
and UO_2730 (O_2730,N_29408,N_29547);
or UO_2731 (O_2731,N_29484,N_29537);
or UO_2732 (O_2732,N_29680,N_29656);
or UO_2733 (O_2733,N_29580,N_29569);
and UO_2734 (O_2734,N_29678,N_29849);
and UO_2735 (O_2735,N_29791,N_29793);
nor UO_2736 (O_2736,N_29708,N_29430);
nand UO_2737 (O_2737,N_29880,N_29914);
nand UO_2738 (O_2738,N_29525,N_29814);
or UO_2739 (O_2739,N_29466,N_29625);
nand UO_2740 (O_2740,N_29541,N_29894);
or UO_2741 (O_2741,N_29933,N_29789);
nor UO_2742 (O_2742,N_29434,N_29768);
xor UO_2743 (O_2743,N_29646,N_29823);
nor UO_2744 (O_2744,N_29609,N_29918);
or UO_2745 (O_2745,N_29609,N_29803);
or UO_2746 (O_2746,N_29789,N_29909);
nand UO_2747 (O_2747,N_29938,N_29457);
and UO_2748 (O_2748,N_29443,N_29780);
nand UO_2749 (O_2749,N_29442,N_29673);
nor UO_2750 (O_2750,N_29964,N_29839);
nand UO_2751 (O_2751,N_29940,N_29637);
or UO_2752 (O_2752,N_29851,N_29902);
nand UO_2753 (O_2753,N_29444,N_29685);
or UO_2754 (O_2754,N_29912,N_29935);
nor UO_2755 (O_2755,N_29864,N_29557);
nand UO_2756 (O_2756,N_29843,N_29543);
xor UO_2757 (O_2757,N_29590,N_29676);
or UO_2758 (O_2758,N_29604,N_29676);
and UO_2759 (O_2759,N_29617,N_29819);
and UO_2760 (O_2760,N_29569,N_29785);
xnor UO_2761 (O_2761,N_29955,N_29570);
nand UO_2762 (O_2762,N_29463,N_29875);
nand UO_2763 (O_2763,N_29526,N_29771);
or UO_2764 (O_2764,N_29552,N_29805);
nor UO_2765 (O_2765,N_29493,N_29835);
xnor UO_2766 (O_2766,N_29591,N_29813);
nor UO_2767 (O_2767,N_29763,N_29743);
nor UO_2768 (O_2768,N_29977,N_29452);
nand UO_2769 (O_2769,N_29487,N_29843);
nand UO_2770 (O_2770,N_29722,N_29975);
nand UO_2771 (O_2771,N_29649,N_29941);
nand UO_2772 (O_2772,N_29801,N_29982);
nor UO_2773 (O_2773,N_29546,N_29668);
nor UO_2774 (O_2774,N_29851,N_29960);
xnor UO_2775 (O_2775,N_29595,N_29683);
nand UO_2776 (O_2776,N_29666,N_29835);
nor UO_2777 (O_2777,N_29654,N_29588);
nand UO_2778 (O_2778,N_29713,N_29628);
nand UO_2779 (O_2779,N_29568,N_29595);
and UO_2780 (O_2780,N_29937,N_29804);
and UO_2781 (O_2781,N_29518,N_29764);
or UO_2782 (O_2782,N_29881,N_29441);
and UO_2783 (O_2783,N_29483,N_29402);
nand UO_2784 (O_2784,N_29486,N_29481);
and UO_2785 (O_2785,N_29841,N_29864);
or UO_2786 (O_2786,N_29733,N_29694);
xnor UO_2787 (O_2787,N_29948,N_29868);
or UO_2788 (O_2788,N_29791,N_29520);
and UO_2789 (O_2789,N_29950,N_29891);
nand UO_2790 (O_2790,N_29888,N_29976);
nor UO_2791 (O_2791,N_29969,N_29864);
nand UO_2792 (O_2792,N_29587,N_29488);
and UO_2793 (O_2793,N_29652,N_29469);
and UO_2794 (O_2794,N_29822,N_29798);
nand UO_2795 (O_2795,N_29923,N_29605);
or UO_2796 (O_2796,N_29654,N_29421);
xor UO_2797 (O_2797,N_29946,N_29755);
and UO_2798 (O_2798,N_29759,N_29933);
or UO_2799 (O_2799,N_29783,N_29689);
nand UO_2800 (O_2800,N_29732,N_29432);
xor UO_2801 (O_2801,N_29713,N_29960);
and UO_2802 (O_2802,N_29620,N_29915);
xnor UO_2803 (O_2803,N_29739,N_29594);
xnor UO_2804 (O_2804,N_29802,N_29850);
xor UO_2805 (O_2805,N_29909,N_29652);
and UO_2806 (O_2806,N_29949,N_29615);
nor UO_2807 (O_2807,N_29876,N_29640);
xnor UO_2808 (O_2808,N_29685,N_29902);
nor UO_2809 (O_2809,N_29695,N_29952);
xor UO_2810 (O_2810,N_29553,N_29999);
nor UO_2811 (O_2811,N_29763,N_29979);
or UO_2812 (O_2812,N_29999,N_29412);
and UO_2813 (O_2813,N_29413,N_29999);
xor UO_2814 (O_2814,N_29918,N_29937);
or UO_2815 (O_2815,N_29506,N_29421);
or UO_2816 (O_2816,N_29823,N_29866);
and UO_2817 (O_2817,N_29491,N_29738);
and UO_2818 (O_2818,N_29669,N_29562);
xnor UO_2819 (O_2819,N_29884,N_29514);
or UO_2820 (O_2820,N_29545,N_29433);
nor UO_2821 (O_2821,N_29717,N_29668);
nand UO_2822 (O_2822,N_29951,N_29644);
nand UO_2823 (O_2823,N_29567,N_29537);
or UO_2824 (O_2824,N_29535,N_29948);
or UO_2825 (O_2825,N_29520,N_29459);
nand UO_2826 (O_2826,N_29601,N_29651);
nor UO_2827 (O_2827,N_29483,N_29808);
xnor UO_2828 (O_2828,N_29559,N_29536);
xnor UO_2829 (O_2829,N_29500,N_29627);
or UO_2830 (O_2830,N_29781,N_29561);
nand UO_2831 (O_2831,N_29814,N_29530);
or UO_2832 (O_2832,N_29852,N_29412);
and UO_2833 (O_2833,N_29636,N_29474);
and UO_2834 (O_2834,N_29606,N_29986);
nor UO_2835 (O_2835,N_29857,N_29541);
or UO_2836 (O_2836,N_29915,N_29482);
or UO_2837 (O_2837,N_29438,N_29868);
and UO_2838 (O_2838,N_29447,N_29785);
nor UO_2839 (O_2839,N_29467,N_29412);
nand UO_2840 (O_2840,N_29467,N_29986);
and UO_2841 (O_2841,N_29627,N_29480);
xor UO_2842 (O_2842,N_29600,N_29740);
xnor UO_2843 (O_2843,N_29667,N_29788);
nand UO_2844 (O_2844,N_29646,N_29731);
or UO_2845 (O_2845,N_29635,N_29584);
or UO_2846 (O_2846,N_29996,N_29762);
xor UO_2847 (O_2847,N_29981,N_29612);
nand UO_2848 (O_2848,N_29770,N_29689);
or UO_2849 (O_2849,N_29630,N_29871);
nor UO_2850 (O_2850,N_29613,N_29612);
nor UO_2851 (O_2851,N_29406,N_29603);
xor UO_2852 (O_2852,N_29467,N_29704);
and UO_2853 (O_2853,N_29779,N_29723);
and UO_2854 (O_2854,N_29462,N_29537);
or UO_2855 (O_2855,N_29478,N_29976);
or UO_2856 (O_2856,N_29933,N_29572);
or UO_2857 (O_2857,N_29766,N_29422);
nor UO_2858 (O_2858,N_29762,N_29665);
and UO_2859 (O_2859,N_29516,N_29630);
and UO_2860 (O_2860,N_29770,N_29451);
nor UO_2861 (O_2861,N_29829,N_29460);
xnor UO_2862 (O_2862,N_29951,N_29661);
or UO_2863 (O_2863,N_29881,N_29494);
nand UO_2864 (O_2864,N_29910,N_29619);
or UO_2865 (O_2865,N_29894,N_29423);
and UO_2866 (O_2866,N_29474,N_29691);
nand UO_2867 (O_2867,N_29530,N_29789);
xnor UO_2868 (O_2868,N_29855,N_29791);
and UO_2869 (O_2869,N_29405,N_29827);
or UO_2870 (O_2870,N_29820,N_29817);
nand UO_2871 (O_2871,N_29605,N_29892);
or UO_2872 (O_2872,N_29569,N_29706);
xnor UO_2873 (O_2873,N_29956,N_29626);
nand UO_2874 (O_2874,N_29414,N_29870);
xnor UO_2875 (O_2875,N_29453,N_29589);
xnor UO_2876 (O_2876,N_29943,N_29689);
and UO_2877 (O_2877,N_29400,N_29424);
nor UO_2878 (O_2878,N_29942,N_29606);
xor UO_2879 (O_2879,N_29525,N_29868);
nor UO_2880 (O_2880,N_29586,N_29945);
nand UO_2881 (O_2881,N_29588,N_29913);
nor UO_2882 (O_2882,N_29913,N_29998);
nand UO_2883 (O_2883,N_29715,N_29748);
nor UO_2884 (O_2884,N_29984,N_29876);
nor UO_2885 (O_2885,N_29649,N_29560);
and UO_2886 (O_2886,N_29759,N_29561);
nor UO_2887 (O_2887,N_29926,N_29426);
nand UO_2888 (O_2888,N_29694,N_29517);
or UO_2889 (O_2889,N_29995,N_29414);
xnor UO_2890 (O_2890,N_29873,N_29801);
nand UO_2891 (O_2891,N_29871,N_29975);
nor UO_2892 (O_2892,N_29453,N_29607);
and UO_2893 (O_2893,N_29480,N_29556);
xnor UO_2894 (O_2894,N_29898,N_29742);
or UO_2895 (O_2895,N_29492,N_29641);
nand UO_2896 (O_2896,N_29758,N_29675);
or UO_2897 (O_2897,N_29722,N_29555);
xnor UO_2898 (O_2898,N_29991,N_29578);
nand UO_2899 (O_2899,N_29859,N_29825);
nand UO_2900 (O_2900,N_29680,N_29476);
nand UO_2901 (O_2901,N_29878,N_29619);
nand UO_2902 (O_2902,N_29703,N_29649);
or UO_2903 (O_2903,N_29752,N_29644);
xor UO_2904 (O_2904,N_29596,N_29504);
nand UO_2905 (O_2905,N_29930,N_29520);
xor UO_2906 (O_2906,N_29846,N_29672);
xnor UO_2907 (O_2907,N_29575,N_29918);
and UO_2908 (O_2908,N_29517,N_29984);
or UO_2909 (O_2909,N_29898,N_29999);
nand UO_2910 (O_2910,N_29576,N_29522);
xor UO_2911 (O_2911,N_29716,N_29988);
nor UO_2912 (O_2912,N_29878,N_29656);
xor UO_2913 (O_2913,N_29541,N_29799);
nand UO_2914 (O_2914,N_29963,N_29970);
nor UO_2915 (O_2915,N_29432,N_29599);
xor UO_2916 (O_2916,N_29616,N_29428);
nand UO_2917 (O_2917,N_29592,N_29715);
and UO_2918 (O_2918,N_29825,N_29920);
and UO_2919 (O_2919,N_29663,N_29661);
nand UO_2920 (O_2920,N_29662,N_29636);
nand UO_2921 (O_2921,N_29493,N_29457);
nor UO_2922 (O_2922,N_29875,N_29610);
or UO_2923 (O_2923,N_29772,N_29607);
nor UO_2924 (O_2924,N_29407,N_29919);
or UO_2925 (O_2925,N_29631,N_29983);
and UO_2926 (O_2926,N_29568,N_29685);
and UO_2927 (O_2927,N_29510,N_29739);
nor UO_2928 (O_2928,N_29860,N_29480);
nor UO_2929 (O_2929,N_29825,N_29959);
or UO_2930 (O_2930,N_29864,N_29649);
xnor UO_2931 (O_2931,N_29787,N_29922);
nor UO_2932 (O_2932,N_29731,N_29818);
nor UO_2933 (O_2933,N_29587,N_29637);
and UO_2934 (O_2934,N_29489,N_29676);
xnor UO_2935 (O_2935,N_29722,N_29683);
and UO_2936 (O_2936,N_29746,N_29811);
xor UO_2937 (O_2937,N_29545,N_29609);
nor UO_2938 (O_2938,N_29598,N_29977);
nand UO_2939 (O_2939,N_29864,N_29420);
nand UO_2940 (O_2940,N_29939,N_29946);
xor UO_2941 (O_2941,N_29974,N_29402);
nand UO_2942 (O_2942,N_29615,N_29787);
nor UO_2943 (O_2943,N_29714,N_29869);
nor UO_2944 (O_2944,N_29985,N_29873);
xor UO_2945 (O_2945,N_29802,N_29958);
and UO_2946 (O_2946,N_29719,N_29660);
xnor UO_2947 (O_2947,N_29481,N_29962);
and UO_2948 (O_2948,N_29868,N_29548);
or UO_2949 (O_2949,N_29748,N_29922);
nor UO_2950 (O_2950,N_29409,N_29715);
xor UO_2951 (O_2951,N_29824,N_29572);
nand UO_2952 (O_2952,N_29639,N_29413);
nor UO_2953 (O_2953,N_29757,N_29675);
or UO_2954 (O_2954,N_29801,N_29429);
nor UO_2955 (O_2955,N_29470,N_29992);
xnor UO_2956 (O_2956,N_29566,N_29888);
and UO_2957 (O_2957,N_29956,N_29452);
and UO_2958 (O_2958,N_29904,N_29758);
nand UO_2959 (O_2959,N_29601,N_29526);
xor UO_2960 (O_2960,N_29497,N_29651);
nor UO_2961 (O_2961,N_29855,N_29729);
nand UO_2962 (O_2962,N_29921,N_29421);
nor UO_2963 (O_2963,N_29561,N_29562);
nand UO_2964 (O_2964,N_29920,N_29519);
nand UO_2965 (O_2965,N_29602,N_29815);
nor UO_2966 (O_2966,N_29581,N_29585);
nand UO_2967 (O_2967,N_29671,N_29829);
nand UO_2968 (O_2968,N_29418,N_29690);
nand UO_2969 (O_2969,N_29415,N_29587);
or UO_2970 (O_2970,N_29628,N_29919);
and UO_2971 (O_2971,N_29854,N_29817);
nand UO_2972 (O_2972,N_29998,N_29721);
xor UO_2973 (O_2973,N_29427,N_29612);
xnor UO_2974 (O_2974,N_29626,N_29671);
and UO_2975 (O_2975,N_29895,N_29527);
xnor UO_2976 (O_2976,N_29534,N_29839);
or UO_2977 (O_2977,N_29929,N_29740);
or UO_2978 (O_2978,N_29828,N_29509);
nand UO_2979 (O_2979,N_29838,N_29699);
or UO_2980 (O_2980,N_29764,N_29458);
or UO_2981 (O_2981,N_29568,N_29631);
nor UO_2982 (O_2982,N_29953,N_29813);
nor UO_2983 (O_2983,N_29950,N_29618);
nor UO_2984 (O_2984,N_29647,N_29485);
nor UO_2985 (O_2985,N_29401,N_29524);
nor UO_2986 (O_2986,N_29707,N_29443);
nor UO_2987 (O_2987,N_29557,N_29418);
nor UO_2988 (O_2988,N_29503,N_29486);
nor UO_2989 (O_2989,N_29515,N_29485);
and UO_2990 (O_2990,N_29735,N_29760);
nand UO_2991 (O_2991,N_29482,N_29745);
nor UO_2992 (O_2992,N_29901,N_29572);
xnor UO_2993 (O_2993,N_29836,N_29561);
nor UO_2994 (O_2994,N_29853,N_29473);
nand UO_2995 (O_2995,N_29743,N_29518);
and UO_2996 (O_2996,N_29880,N_29773);
nor UO_2997 (O_2997,N_29464,N_29857);
nor UO_2998 (O_2998,N_29889,N_29786);
nand UO_2999 (O_2999,N_29795,N_29671);
nor UO_3000 (O_3000,N_29925,N_29870);
nor UO_3001 (O_3001,N_29581,N_29639);
or UO_3002 (O_3002,N_29476,N_29470);
nand UO_3003 (O_3003,N_29434,N_29431);
and UO_3004 (O_3004,N_29596,N_29640);
nor UO_3005 (O_3005,N_29619,N_29844);
xor UO_3006 (O_3006,N_29619,N_29879);
or UO_3007 (O_3007,N_29433,N_29715);
or UO_3008 (O_3008,N_29842,N_29777);
xor UO_3009 (O_3009,N_29823,N_29514);
or UO_3010 (O_3010,N_29826,N_29913);
nor UO_3011 (O_3011,N_29975,N_29512);
xor UO_3012 (O_3012,N_29552,N_29989);
xor UO_3013 (O_3013,N_29980,N_29855);
nand UO_3014 (O_3014,N_29578,N_29855);
xnor UO_3015 (O_3015,N_29496,N_29816);
xor UO_3016 (O_3016,N_29858,N_29780);
xnor UO_3017 (O_3017,N_29620,N_29583);
and UO_3018 (O_3018,N_29951,N_29811);
and UO_3019 (O_3019,N_29637,N_29853);
or UO_3020 (O_3020,N_29517,N_29937);
nor UO_3021 (O_3021,N_29752,N_29513);
xor UO_3022 (O_3022,N_29404,N_29830);
nor UO_3023 (O_3023,N_29986,N_29510);
nor UO_3024 (O_3024,N_29408,N_29567);
and UO_3025 (O_3025,N_29959,N_29459);
nand UO_3026 (O_3026,N_29903,N_29671);
and UO_3027 (O_3027,N_29547,N_29648);
nor UO_3028 (O_3028,N_29436,N_29962);
nand UO_3029 (O_3029,N_29887,N_29938);
and UO_3030 (O_3030,N_29698,N_29604);
xor UO_3031 (O_3031,N_29659,N_29985);
nand UO_3032 (O_3032,N_29643,N_29663);
nor UO_3033 (O_3033,N_29703,N_29848);
xnor UO_3034 (O_3034,N_29724,N_29476);
or UO_3035 (O_3035,N_29949,N_29744);
xor UO_3036 (O_3036,N_29422,N_29517);
and UO_3037 (O_3037,N_29643,N_29794);
or UO_3038 (O_3038,N_29826,N_29452);
nand UO_3039 (O_3039,N_29706,N_29673);
or UO_3040 (O_3040,N_29403,N_29831);
nor UO_3041 (O_3041,N_29880,N_29562);
or UO_3042 (O_3042,N_29865,N_29850);
nor UO_3043 (O_3043,N_29715,N_29805);
and UO_3044 (O_3044,N_29607,N_29732);
or UO_3045 (O_3045,N_29981,N_29743);
nand UO_3046 (O_3046,N_29979,N_29460);
nor UO_3047 (O_3047,N_29826,N_29616);
nor UO_3048 (O_3048,N_29827,N_29618);
nand UO_3049 (O_3049,N_29506,N_29581);
xnor UO_3050 (O_3050,N_29763,N_29406);
and UO_3051 (O_3051,N_29928,N_29589);
nand UO_3052 (O_3052,N_29797,N_29493);
xnor UO_3053 (O_3053,N_29484,N_29571);
and UO_3054 (O_3054,N_29498,N_29600);
xnor UO_3055 (O_3055,N_29673,N_29705);
xor UO_3056 (O_3056,N_29926,N_29799);
nor UO_3057 (O_3057,N_29778,N_29774);
xnor UO_3058 (O_3058,N_29653,N_29645);
xor UO_3059 (O_3059,N_29604,N_29910);
and UO_3060 (O_3060,N_29609,N_29947);
xnor UO_3061 (O_3061,N_29464,N_29506);
nor UO_3062 (O_3062,N_29418,N_29929);
or UO_3063 (O_3063,N_29917,N_29914);
or UO_3064 (O_3064,N_29469,N_29844);
nor UO_3065 (O_3065,N_29924,N_29511);
nand UO_3066 (O_3066,N_29446,N_29406);
and UO_3067 (O_3067,N_29944,N_29867);
or UO_3068 (O_3068,N_29770,N_29505);
xor UO_3069 (O_3069,N_29620,N_29982);
nand UO_3070 (O_3070,N_29858,N_29916);
nand UO_3071 (O_3071,N_29702,N_29753);
or UO_3072 (O_3072,N_29466,N_29409);
xnor UO_3073 (O_3073,N_29911,N_29918);
xnor UO_3074 (O_3074,N_29505,N_29665);
or UO_3075 (O_3075,N_29773,N_29992);
xnor UO_3076 (O_3076,N_29542,N_29764);
nand UO_3077 (O_3077,N_29512,N_29482);
nor UO_3078 (O_3078,N_29535,N_29806);
and UO_3079 (O_3079,N_29447,N_29739);
xnor UO_3080 (O_3080,N_29906,N_29859);
nor UO_3081 (O_3081,N_29418,N_29657);
and UO_3082 (O_3082,N_29765,N_29829);
or UO_3083 (O_3083,N_29856,N_29800);
nor UO_3084 (O_3084,N_29539,N_29600);
or UO_3085 (O_3085,N_29931,N_29423);
nor UO_3086 (O_3086,N_29708,N_29993);
nor UO_3087 (O_3087,N_29645,N_29496);
nor UO_3088 (O_3088,N_29631,N_29964);
and UO_3089 (O_3089,N_29909,N_29821);
and UO_3090 (O_3090,N_29890,N_29685);
and UO_3091 (O_3091,N_29583,N_29623);
or UO_3092 (O_3092,N_29967,N_29478);
nand UO_3093 (O_3093,N_29911,N_29509);
and UO_3094 (O_3094,N_29703,N_29606);
or UO_3095 (O_3095,N_29629,N_29464);
nand UO_3096 (O_3096,N_29885,N_29627);
xor UO_3097 (O_3097,N_29803,N_29665);
nor UO_3098 (O_3098,N_29612,N_29687);
nand UO_3099 (O_3099,N_29860,N_29486);
nand UO_3100 (O_3100,N_29980,N_29983);
nor UO_3101 (O_3101,N_29911,N_29587);
nor UO_3102 (O_3102,N_29426,N_29711);
or UO_3103 (O_3103,N_29894,N_29985);
xor UO_3104 (O_3104,N_29868,N_29753);
nand UO_3105 (O_3105,N_29891,N_29990);
xnor UO_3106 (O_3106,N_29964,N_29576);
and UO_3107 (O_3107,N_29466,N_29494);
and UO_3108 (O_3108,N_29857,N_29415);
or UO_3109 (O_3109,N_29937,N_29885);
xnor UO_3110 (O_3110,N_29922,N_29652);
xor UO_3111 (O_3111,N_29865,N_29798);
xnor UO_3112 (O_3112,N_29714,N_29533);
or UO_3113 (O_3113,N_29912,N_29473);
nand UO_3114 (O_3114,N_29513,N_29673);
xor UO_3115 (O_3115,N_29823,N_29709);
nor UO_3116 (O_3116,N_29985,N_29925);
xnor UO_3117 (O_3117,N_29928,N_29513);
and UO_3118 (O_3118,N_29659,N_29442);
nand UO_3119 (O_3119,N_29854,N_29833);
or UO_3120 (O_3120,N_29979,N_29798);
and UO_3121 (O_3121,N_29778,N_29990);
xor UO_3122 (O_3122,N_29881,N_29601);
nand UO_3123 (O_3123,N_29482,N_29949);
and UO_3124 (O_3124,N_29600,N_29556);
and UO_3125 (O_3125,N_29736,N_29887);
and UO_3126 (O_3126,N_29953,N_29554);
nor UO_3127 (O_3127,N_29839,N_29722);
nor UO_3128 (O_3128,N_29641,N_29521);
xor UO_3129 (O_3129,N_29769,N_29570);
nand UO_3130 (O_3130,N_29422,N_29972);
xnor UO_3131 (O_3131,N_29656,N_29824);
nor UO_3132 (O_3132,N_29409,N_29579);
and UO_3133 (O_3133,N_29766,N_29556);
or UO_3134 (O_3134,N_29935,N_29880);
nor UO_3135 (O_3135,N_29634,N_29958);
nand UO_3136 (O_3136,N_29749,N_29488);
nor UO_3137 (O_3137,N_29886,N_29913);
and UO_3138 (O_3138,N_29844,N_29875);
nor UO_3139 (O_3139,N_29470,N_29496);
nor UO_3140 (O_3140,N_29594,N_29821);
or UO_3141 (O_3141,N_29882,N_29665);
and UO_3142 (O_3142,N_29861,N_29679);
xnor UO_3143 (O_3143,N_29643,N_29401);
or UO_3144 (O_3144,N_29965,N_29795);
nand UO_3145 (O_3145,N_29967,N_29804);
and UO_3146 (O_3146,N_29972,N_29624);
nand UO_3147 (O_3147,N_29627,N_29755);
nand UO_3148 (O_3148,N_29551,N_29896);
xnor UO_3149 (O_3149,N_29604,N_29981);
or UO_3150 (O_3150,N_29668,N_29408);
xnor UO_3151 (O_3151,N_29476,N_29606);
and UO_3152 (O_3152,N_29452,N_29884);
and UO_3153 (O_3153,N_29600,N_29915);
or UO_3154 (O_3154,N_29905,N_29728);
xor UO_3155 (O_3155,N_29727,N_29908);
nand UO_3156 (O_3156,N_29931,N_29481);
and UO_3157 (O_3157,N_29998,N_29962);
nor UO_3158 (O_3158,N_29783,N_29912);
or UO_3159 (O_3159,N_29857,N_29722);
nand UO_3160 (O_3160,N_29792,N_29918);
or UO_3161 (O_3161,N_29631,N_29814);
nor UO_3162 (O_3162,N_29841,N_29722);
xor UO_3163 (O_3163,N_29580,N_29876);
nand UO_3164 (O_3164,N_29595,N_29423);
and UO_3165 (O_3165,N_29463,N_29683);
xnor UO_3166 (O_3166,N_29719,N_29937);
xnor UO_3167 (O_3167,N_29741,N_29615);
nor UO_3168 (O_3168,N_29829,N_29476);
xor UO_3169 (O_3169,N_29961,N_29483);
nor UO_3170 (O_3170,N_29817,N_29948);
nor UO_3171 (O_3171,N_29528,N_29743);
nor UO_3172 (O_3172,N_29810,N_29760);
or UO_3173 (O_3173,N_29565,N_29988);
nor UO_3174 (O_3174,N_29703,N_29548);
nor UO_3175 (O_3175,N_29401,N_29671);
xnor UO_3176 (O_3176,N_29902,N_29495);
and UO_3177 (O_3177,N_29614,N_29925);
nor UO_3178 (O_3178,N_29519,N_29962);
or UO_3179 (O_3179,N_29694,N_29791);
or UO_3180 (O_3180,N_29632,N_29621);
and UO_3181 (O_3181,N_29626,N_29602);
xnor UO_3182 (O_3182,N_29831,N_29427);
nor UO_3183 (O_3183,N_29585,N_29482);
xnor UO_3184 (O_3184,N_29911,N_29568);
xnor UO_3185 (O_3185,N_29480,N_29607);
or UO_3186 (O_3186,N_29812,N_29843);
xor UO_3187 (O_3187,N_29990,N_29760);
or UO_3188 (O_3188,N_29609,N_29834);
nand UO_3189 (O_3189,N_29978,N_29494);
nand UO_3190 (O_3190,N_29958,N_29532);
and UO_3191 (O_3191,N_29817,N_29809);
or UO_3192 (O_3192,N_29782,N_29895);
nand UO_3193 (O_3193,N_29915,N_29810);
nand UO_3194 (O_3194,N_29905,N_29776);
nand UO_3195 (O_3195,N_29719,N_29642);
nand UO_3196 (O_3196,N_29616,N_29423);
and UO_3197 (O_3197,N_29649,N_29469);
xnor UO_3198 (O_3198,N_29715,N_29991);
nand UO_3199 (O_3199,N_29779,N_29979);
nand UO_3200 (O_3200,N_29752,N_29579);
and UO_3201 (O_3201,N_29919,N_29946);
nand UO_3202 (O_3202,N_29936,N_29452);
xnor UO_3203 (O_3203,N_29784,N_29971);
and UO_3204 (O_3204,N_29854,N_29418);
nand UO_3205 (O_3205,N_29477,N_29689);
xnor UO_3206 (O_3206,N_29406,N_29826);
and UO_3207 (O_3207,N_29532,N_29803);
and UO_3208 (O_3208,N_29829,N_29405);
xor UO_3209 (O_3209,N_29731,N_29613);
or UO_3210 (O_3210,N_29945,N_29496);
nor UO_3211 (O_3211,N_29898,N_29635);
xnor UO_3212 (O_3212,N_29926,N_29813);
xnor UO_3213 (O_3213,N_29903,N_29742);
xor UO_3214 (O_3214,N_29487,N_29707);
nor UO_3215 (O_3215,N_29787,N_29439);
nand UO_3216 (O_3216,N_29466,N_29782);
nor UO_3217 (O_3217,N_29519,N_29972);
xor UO_3218 (O_3218,N_29597,N_29618);
and UO_3219 (O_3219,N_29844,N_29511);
nor UO_3220 (O_3220,N_29885,N_29813);
and UO_3221 (O_3221,N_29707,N_29571);
or UO_3222 (O_3222,N_29685,N_29743);
and UO_3223 (O_3223,N_29563,N_29889);
nand UO_3224 (O_3224,N_29716,N_29441);
xor UO_3225 (O_3225,N_29869,N_29743);
nor UO_3226 (O_3226,N_29886,N_29467);
and UO_3227 (O_3227,N_29718,N_29724);
or UO_3228 (O_3228,N_29436,N_29551);
and UO_3229 (O_3229,N_29822,N_29408);
nand UO_3230 (O_3230,N_29510,N_29505);
xor UO_3231 (O_3231,N_29696,N_29965);
or UO_3232 (O_3232,N_29410,N_29901);
nor UO_3233 (O_3233,N_29695,N_29546);
xnor UO_3234 (O_3234,N_29773,N_29857);
nand UO_3235 (O_3235,N_29608,N_29526);
or UO_3236 (O_3236,N_29845,N_29702);
nor UO_3237 (O_3237,N_29614,N_29433);
xor UO_3238 (O_3238,N_29622,N_29918);
nor UO_3239 (O_3239,N_29806,N_29615);
nor UO_3240 (O_3240,N_29601,N_29519);
nor UO_3241 (O_3241,N_29756,N_29501);
nor UO_3242 (O_3242,N_29899,N_29828);
nor UO_3243 (O_3243,N_29797,N_29757);
nor UO_3244 (O_3244,N_29997,N_29987);
nor UO_3245 (O_3245,N_29447,N_29722);
nand UO_3246 (O_3246,N_29721,N_29786);
nand UO_3247 (O_3247,N_29965,N_29878);
nor UO_3248 (O_3248,N_29611,N_29622);
or UO_3249 (O_3249,N_29760,N_29896);
xnor UO_3250 (O_3250,N_29930,N_29554);
nor UO_3251 (O_3251,N_29997,N_29618);
or UO_3252 (O_3252,N_29795,N_29714);
xnor UO_3253 (O_3253,N_29818,N_29460);
nor UO_3254 (O_3254,N_29532,N_29985);
or UO_3255 (O_3255,N_29430,N_29608);
or UO_3256 (O_3256,N_29966,N_29566);
nor UO_3257 (O_3257,N_29662,N_29638);
or UO_3258 (O_3258,N_29885,N_29511);
nor UO_3259 (O_3259,N_29514,N_29752);
nand UO_3260 (O_3260,N_29479,N_29826);
nor UO_3261 (O_3261,N_29465,N_29671);
xor UO_3262 (O_3262,N_29935,N_29999);
or UO_3263 (O_3263,N_29440,N_29948);
xnor UO_3264 (O_3264,N_29482,N_29688);
nand UO_3265 (O_3265,N_29433,N_29970);
and UO_3266 (O_3266,N_29850,N_29489);
nand UO_3267 (O_3267,N_29617,N_29910);
nor UO_3268 (O_3268,N_29511,N_29467);
nor UO_3269 (O_3269,N_29551,N_29934);
xor UO_3270 (O_3270,N_29656,N_29766);
nand UO_3271 (O_3271,N_29781,N_29837);
and UO_3272 (O_3272,N_29808,N_29599);
or UO_3273 (O_3273,N_29690,N_29740);
or UO_3274 (O_3274,N_29439,N_29606);
xor UO_3275 (O_3275,N_29570,N_29788);
nor UO_3276 (O_3276,N_29657,N_29989);
and UO_3277 (O_3277,N_29742,N_29652);
nor UO_3278 (O_3278,N_29919,N_29733);
or UO_3279 (O_3279,N_29825,N_29405);
nand UO_3280 (O_3280,N_29644,N_29787);
nor UO_3281 (O_3281,N_29634,N_29840);
nor UO_3282 (O_3282,N_29547,N_29704);
and UO_3283 (O_3283,N_29927,N_29447);
xor UO_3284 (O_3284,N_29648,N_29706);
xor UO_3285 (O_3285,N_29418,N_29987);
nand UO_3286 (O_3286,N_29488,N_29809);
and UO_3287 (O_3287,N_29698,N_29425);
or UO_3288 (O_3288,N_29829,N_29731);
nor UO_3289 (O_3289,N_29490,N_29637);
and UO_3290 (O_3290,N_29870,N_29807);
nor UO_3291 (O_3291,N_29671,N_29573);
and UO_3292 (O_3292,N_29699,N_29842);
and UO_3293 (O_3293,N_29493,N_29891);
nor UO_3294 (O_3294,N_29498,N_29992);
and UO_3295 (O_3295,N_29703,N_29720);
xor UO_3296 (O_3296,N_29472,N_29656);
nor UO_3297 (O_3297,N_29672,N_29815);
nand UO_3298 (O_3298,N_29801,N_29694);
nor UO_3299 (O_3299,N_29869,N_29913);
xor UO_3300 (O_3300,N_29875,N_29584);
nand UO_3301 (O_3301,N_29725,N_29833);
and UO_3302 (O_3302,N_29709,N_29986);
or UO_3303 (O_3303,N_29444,N_29793);
or UO_3304 (O_3304,N_29460,N_29853);
xor UO_3305 (O_3305,N_29427,N_29455);
and UO_3306 (O_3306,N_29612,N_29421);
nand UO_3307 (O_3307,N_29891,N_29653);
xnor UO_3308 (O_3308,N_29738,N_29817);
nand UO_3309 (O_3309,N_29792,N_29824);
and UO_3310 (O_3310,N_29480,N_29779);
xnor UO_3311 (O_3311,N_29971,N_29679);
nand UO_3312 (O_3312,N_29872,N_29506);
nor UO_3313 (O_3313,N_29895,N_29968);
xnor UO_3314 (O_3314,N_29551,N_29942);
or UO_3315 (O_3315,N_29944,N_29676);
xor UO_3316 (O_3316,N_29665,N_29670);
nor UO_3317 (O_3317,N_29838,N_29489);
and UO_3318 (O_3318,N_29451,N_29698);
and UO_3319 (O_3319,N_29882,N_29560);
or UO_3320 (O_3320,N_29954,N_29951);
xor UO_3321 (O_3321,N_29649,N_29461);
and UO_3322 (O_3322,N_29771,N_29673);
nor UO_3323 (O_3323,N_29449,N_29679);
or UO_3324 (O_3324,N_29759,N_29969);
or UO_3325 (O_3325,N_29568,N_29979);
nand UO_3326 (O_3326,N_29674,N_29836);
nand UO_3327 (O_3327,N_29761,N_29580);
and UO_3328 (O_3328,N_29419,N_29534);
nor UO_3329 (O_3329,N_29418,N_29628);
xnor UO_3330 (O_3330,N_29502,N_29429);
and UO_3331 (O_3331,N_29574,N_29690);
nor UO_3332 (O_3332,N_29826,N_29728);
xnor UO_3333 (O_3333,N_29400,N_29823);
xnor UO_3334 (O_3334,N_29627,N_29667);
xnor UO_3335 (O_3335,N_29770,N_29737);
nand UO_3336 (O_3336,N_29770,N_29776);
nor UO_3337 (O_3337,N_29533,N_29885);
nand UO_3338 (O_3338,N_29802,N_29597);
or UO_3339 (O_3339,N_29716,N_29672);
or UO_3340 (O_3340,N_29614,N_29717);
and UO_3341 (O_3341,N_29439,N_29986);
nand UO_3342 (O_3342,N_29631,N_29490);
nor UO_3343 (O_3343,N_29830,N_29702);
nand UO_3344 (O_3344,N_29730,N_29934);
or UO_3345 (O_3345,N_29694,N_29896);
nand UO_3346 (O_3346,N_29819,N_29826);
nand UO_3347 (O_3347,N_29681,N_29923);
xnor UO_3348 (O_3348,N_29879,N_29595);
or UO_3349 (O_3349,N_29744,N_29640);
nand UO_3350 (O_3350,N_29807,N_29584);
xor UO_3351 (O_3351,N_29599,N_29860);
nor UO_3352 (O_3352,N_29534,N_29725);
or UO_3353 (O_3353,N_29894,N_29547);
nand UO_3354 (O_3354,N_29954,N_29796);
nand UO_3355 (O_3355,N_29545,N_29828);
nor UO_3356 (O_3356,N_29696,N_29912);
nand UO_3357 (O_3357,N_29873,N_29983);
xor UO_3358 (O_3358,N_29550,N_29661);
xor UO_3359 (O_3359,N_29929,N_29463);
xnor UO_3360 (O_3360,N_29961,N_29768);
nor UO_3361 (O_3361,N_29990,N_29548);
nand UO_3362 (O_3362,N_29739,N_29604);
nand UO_3363 (O_3363,N_29824,N_29490);
nor UO_3364 (O_3364,N_29762,N_29821);
nand UO_3365 (O_3365,N_29857,N_29569);
nand UO_3366 (O_3366,N_29410,N_29433);
or UO_3367 (O_3367,N_29445,N_29862);
xor UO_3368 (O_3368,N_29606,N_29639);
xnor UO_3369 (O_3369,N_29766,N_29845);
or UO_3370 (O_3370,N_29713,N_29717);
xor UO_3371 (O_3371,N_29697,N_29653);
nor UO_3372 (O_3372,N_29872,N_29928);
or UO_3373 (O_3373,N_29650,N_29792);
nor UO_3374 (O_3374,N_29998,N_29689);
or UO_3375 (O_3375,N_29655,N_29992);
xnor UO_3376 (O_3376,N_29635,N_29534);
xnor UO_3377 (O_3377,N_29890,N_29568);
xor UO_3378 (O_3378,N_29639,N_29417);
nor UO_3379 (O_3379,N_29427,N_29525);
nand UO_3380 (O_3380,N_29426,N_29843);
xnor UO_3381 (O_3381,N_29729,N_29866);
nor UO_3382 (O_3382,N_29679,N_29919);
and UO_3383 (O_3383,N_29863,N_29908);
and UO_3384 (O_3384,N_29691,N_29786);
nor UO_3385 (O_3385,N_29420,N_29689);
nor UO_3386 (O_3386,N_29406,N_29842);
nor UO_3387 (O_3387,N_29902,N_29811);
nor UO_3388 (O_3388,N_29873,N_29872);
and UO_3389 (O_3389,N_29620,N_29571);
and UO_3390 (O_3390,N_29961,N_29627);
nor UO_3391 (O_3391,N_29841,N_29789);
nand UO_3392 (O_3392,N_29510,N_29451);
or UO_3393 (O_3393,N_29683,N_29925);
nor UO_3394 (O_3394,N_29812,N_29607);
nor UO_3395 (O_3395,N_29673,N_29610);
and UO_3396 (O_3396,N_29577,N_29985);
xor UO_3397 (O_3397,N_29815,N_29675);
or UO_3398 (O_3398,N_29536,N_29515);
nor UO_3399 (O_3399,N_29785,N_29581);
nor UO_3400 (O_3400,N_29856,N_29961);
nand UO_3401 (O_3401,N_29886,N_29431);
xor UO_3402 (O_3402,N_29651,N_29756);
nor UO_3403 (O_3403,N_29861,N_29867);
nor UO_3404 (O_3404,N_29991,N_29724);
nand UO_3405 (O_3405,N_29649,N_29650);
and UO_3406 (O_3406,N_29830,N_29673);
nor UO_3407 (O_3407,N_29920,N_29874);
nor UO_3408 (O_3408,N_29564,N_29410);
or UO_3409 (O_3409,N_29435,N_29740);
xor UO_3410 (O_3410,N_29587,N_29917);
xor UO_3411 (O_3411,N_29520,N_29870);
xor UO_3412 (O_3412,N_29973,N_29936);
or UO_3413 (O_3413,N_29653,N_29542);
xor UO_3414 (O_3414,N_29813,N_29423);
xnor UO_3415 (O_3415,N_29746,N_29801);
and UO_3416 (O_3416,N_29596,N_29486);
nor UO_3417 (O_3417,N_29978,N_29698);
nor UO_3418 (O_3418,N_29542,N_29709);
xor UO_3419 (O_3419,N_29889,N_29602);
or UO_3420 (O_3420,N_29686,N_29544);
and UO_3421 (O_3421,N_29773,N_29426);
nor UO_3422 (O_3422,N_29731,N_29909);
nand UO_3423 (O_3423,N_29545,N_29956);
xnor UO_3424 (O_3424,N_29893,N_29805);
nor UO_3425 (O_3425,N_29945,N_29480);
or UO_3426 (O_3426,N_29522,N_29730);
nand UO_3427 (O_3427,N_29992,N_29638);
and UO_3428 (O_3428,N_29531,N_29912);
nor UO_3429 (O_3429,N_29703,N_29806);
or UO_3430 (O_3430,N_29506,N_29815);
and UO_3431 (O_3431,N_29746,N_29884);
and UO_3432 (O_3432,N_29598,N_29654);
nor UO_3433 (O_3433,N_29806,N_29537);
xor UO_3434 (O_3434,N_29694,N_29406);
xnor UO_3435 (O_3435,N_29539,N_29954);
nor UO_3436 (O_3436,N_29596,N_29403);
and UO_3437 (O_3437,N_29901,N_29940);
and UO_3438 (O_3438,N_29751,N_29447);
or UO_3439 (O_3439,N_29686,N_29501);
nand UO_3440 (O_3440,N_29951,N_29764);
nor UO_3441 (O_3441,N_29900,N_29784);
nor UO_3442 (O_3442,N_29678,N_29636);
nand UO_3443 (O_3443,N_29613,N_29784);
nor UO_3444 (O_3444,N_29562,N_29695);
nor UO_3445 (O_3445,N_29475,N_29928);
xnor UO_3446 (O_3446,N_29709,N_29592);
xor UO_3447 (O_3447,N_29609,N_29548);
nand UO_3448 (O_3448,N_29545,N_29625);
xnor UO_3449 (O_3449,N_29509,N_29540);
or UO_3450 (O_3450,N_29813,N_29652);
nand UO_3451 (O_3451,N_29762,N_29673);
nor UO_3452 (O_3452,N_29717,N_29673);
xnor UO_3453 (O_3453,N_29862,N_29710);
and UO_3454 (O_3454,N_29661,N_29741);
nand UO_3455 (O_3455,N_29476,N_29942);
and UO_3456 (O_3456,N_29609,N_29568);
nor UO_3457 (O_3457,N_29980,N_29634);
xor UO_3458 (O_3458,N_29894,N_29973);
nand UO_3459 (O_3459,N_29546,N_29859);
nor UO_3460 (O_3460,N_29775,N_29459);
and UO_3461 (O_3461,N_29907,N_29736);
and UO_3462 (O_3462,N_29973,N_29956);
and UO_3463 (O_3463,N_29641,N_29781);
nand UO_3464 (O_3464,N_29487,N_29845);
or UO_3465 (O_3465,N_29594,N_29551);
xnor UO_3466 (O_3466,N_29560,N_29996);
and UO_3467 (O_3467,N_29602,N_29983);
xnor UO_3468 (O_3468,N_29628,N_29706);
xnor UO_3469 (O_3469,N_29698,N_29703);
or UO_3470 (O_3470,N_29474,N_29460);
xnor UO_3471 (O_3471,N_29998,N_29790);
nor UO_3472 (O_3472,N_29639,N_29412);
nor UO_3473 (O_3473,N_29726,N_29445);
nand UO_3474 (O_3474,N_29743,N_29771);
nor UO_3475 (O_3475,N_29565,N_29413);
xnor UO_3476 (O_3476,N_29881,N_29770);
and UO_3477 (O_3477,N_29876,N_29926);
xor UO_3478 (O_3478,N_29403,N_29920);
and UO_3479 (O_3479,N_29437,N_29689);
xor UO_3480 (O_3480,N_29820,N_29673);
nand UO_3481 (O_3481,N_29854,N_29869);
xnor UO_3482 (O_3482,N_29755,N_29573);
nor UO_3483 (O_3483,N_29506,N_29590);
nor UO_3484 (O_3484,N_29697,N_29443);
or UO_3485 (O_3485,N_29413,N_29774);
xnor UO_3486 (O_3486,N_29809,N_29983);
nand UO_3487 (O_3487,N_29718,N_29622);
nand UO_3488 (O_3488,N_29856,N_29881);
nand UO_3489 (O_3489,N_29713,N_29729);
and UO_3490 (O_3490,N_29664,N_29811);
and UO_3491 (O_3491,N_29709,N_29514);
nor UO_3492 (O_3492,N_29669,N_29763);
nand UO_3493 (O_3493,N_29471,N_29662);
or UO_3494 (O_3494,N_29571,N_29607);
or UO_3495 (O_3495,N_29739,N_29708);
xor UO_3496 (O_3496,N_29753,N_29586);
and UO_3497 (O_3497,N_29562,N_29512);
and UO_3498 (O_3498,N_29934,N_29983);
and UO_3499 (O_3499,N_29925,N_29618);
endmodule