module basic_1500_15000_2000_100_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
xor U0 (N_0,In_1464,In_1167);
or U1 (N_1,In_242,In_1321);
or U2 (N_2,In_1082,In_1488);
or U3 (N_3,In_400,In_798);
xor U4 (N_4,In_962,In_308);
nand U5 (N_5,In_142,In_854);
nand U6 (N_6,In_443,In_673);
or U7 (N_7,In_964,In_1411);
and U8 (N_8,In_374,In_508);
xor U9 (N_9,In_956,In_1415);
nor U10 (N_10,In_605,In_1124);
or U11 (N_11,In_594,In_728);
nand U12 (N_12,In_74,In_1423);
nand U13 (N_13,In_992,In_106);
and U14 (N_14,In_205,In_586);
nor U15 (N_15,In_1192,In_395);
and U16 (N_16,In_1177,In_872);
nor U17 (N_17,In_700,In_104);
or U18 (N_18,In_628,In_689);
nor U19 (N_19,In_1202,In_567);
and U20 (N_20,In_321,In_705);
xor U21 (N_21,In_161,In_289);
nand U22 (N_22,In_917,In_758);
nor U23 (N_23,In_709,In_760);
nor U24 (N_24,In_1190,In_265);
or U25 (N_25,In_723,In_47);
xnor U26 (N_26,In_1022,In_1311);
nand U27 (N_27,In_555,In_550);
xnor U28 (N_28,In_561,In_1199);
nand U29 (N_29,In_422,In_152);
nand U30 (N_30,In_816,In_488);
and U31 (N_31,In_973,In_46);
and U32 (N_32,In_721,In_1323);
or U33 (N_33,In_473,In_952);
nand U34 (N_34,In_1481,In_1032);
nand U35 (N_35,In_295,In_41);
xnor U36 (N_36,In_989,In_1000);
and U37 (N_37,In_100,In_1383);
and U38 (N_38,In_334,In_82);
xor U39 (N_39,In_680,In_189);
or U40 (N_40,In_571,In_984);
xor U41 (N_41,In_252,In_12);
nand U42 (N_42,In_1368,In_359);
nand U43 (N_43,In_426,In_707);
and U44 (N_44,In_512,In_271);
and U45 (N_45,In_339,In_472);
nand U46 (N_46,In_736,In_183);
nor U47 (N_47,In_95,In_1157);
or U48 (N_48,In_195,In_479);
nor U49 (N_49,In_887,In_725);
and U50 (N_50,In_1286,In_1444);
nor U51 (N_51,In_1017,In_968);
and U52 (N_52,In_1136,In_314);
nor U53 (N_53,In_873,In_1008);
and U54 (N_54,In_68,In_52);
nand U55 (N_55,In_955,In_622);
nand U56 (N_56,In_196,In_909);
xnor U57 (N_57,In_53,In_625);
nor U58 (N_58,In_766,In_1088);
or U59 (N_59,In_480,In_1206);
and U60 (N_60,In_171,In_1332);
nand U61 (N_61,In_696,In_1356);
nand U62 (N_62,In_893,In_869);
xnor U63 (N_63,In_897,In_1033);
nor U64 (N_64,In_800,In_1009);
nand U65 (N_65,In_1341,In_540);
nand U66 (N_66,In_1319,In_724);
nand U67 (N_67,In_1402,In_1163);
and U68 (N_68,In_115,In_1492);
xnor U69 (N_69,In_1456,In_1059);
or U70 (N_70,In_578,In_225);
or U71 (N_71,In_838,In_665);
xnor U72 (N_72,In_948,In_911);
and U73 (N_73,In_965,In_806);
xor U74 (N_74,In_509,In_783);
nand U75 (N_75,In_312,In_457);
xor U76 (N_76,In_484,In_388);
or U77 (N_77,In_1426,In_1230);
or U78 (N_78,In_967,In_716);
xor U79 (N_79,In_1123,In_497);
nor U80 (N_80,In_1361,In_1495);
and U81 (N_81,In_356,In_603);
or U82 (N_82,In_895,In_519);
xor U83 (N_83,In_785,In_37);
xnor U84 (N_84,In_293,In_514);
nand U85 (N_85,In_1300,In_849);
nand U86 (N_86,In_268,In_902);
nand U87 (N_87,In_391,In_582);
nor U88 (N_88,In_1493,In_450);
nand U89 (N_89,In_524,In_1148);
xnor U90 (N_90,In_1340,In_20);
nor U91 (N_91,In_1364,In_33);
or U92 (N_92,In_796,In_1197);
or U93 (N_93,In_270,In_362);
and U94 (N_94,In_498,In_1299);
xor U95 (N_95,In_311,In_1486);
nor U96 (N_96,In_194,In_1469);
nor U97 (N_97,In_1186,In_392);
or U98 (N_98,In_1246,In_1098);
and U99 (N_99,In_1019,In_584);
nor U100 (N_100,In_1066,In_454);
or U101 (N_101,In_1086,In_1331);
and U102 (N_102,In_536,In_291);
nor U103 (N_103,In_1229,In_495);
nand U104 (N_104,In_1362,In_879);
nor U105 (N_105,In_589,In_31);
and U106 (N_106,In_89,In_912);
xnor U107 (N_107,In_1371,In_939);
or U108 (N_108,In_1035,In_633);
nand U109 (N_109,In_1475,In_1304);
or U110 (N_110,In_674,In_544);
nor U111 (N_111,In_62,In_565);
nor U112 (N_112,In_1313,In_562);
xor U113 (N_113,In_1328,In_537);
and U114 (N_114,In_1222,In_640);
nand U115 (N_115,In_44,In_847);
and U116 (N_116,In_1428,In_373);
nand U117 (N_117,In_292,In_1373);
nand U118 (N_118,In_652,In_23);
nand U119 (N_119,In_1350,In_735);
or U120 (N_120,In_837,In_1215);
or U121 (N_121,In_344,In_126);
nand U122 (N_122,In_699,In_803);
xnor U123 (N_123,In_963,In_79);
and U124 (N_124,In_814,In_315);
or U125 (N_125,In_198,In_330);
or U126 (N_126,In_502,In_752);
nand U127 (N_127,In_780,In_1380);
xnor U128 (N_128,In_1291,In_842);
nor U129 (N_129,In_431,In_539);
and U130 (N_130,In_990,In_1182);
or U131 (N_131,In_220,In_1139);
nor U132 (N_132,In_207,In_279);
nand U133 (N_133,In_98,In_925);
and U134 (N_134,In_483,In_178);
and U135 (N_135,In_831,In_135);
or U136 (N_136,In_1450,In_13);
nor U137 (N_137,In_453,In_1422);
xor U138 (N_138,In_868,In_1375);
xor U139 (N_139,In_923,In_212);
and U140 (N_140,In_995,In_254);
nor U141 (N_141,In_210,In_610);
nor U142 (N_142,In_193,In_1121);
nand U143 (N_143,In_883,In_181);
xor U144 (N_144,In_935,In_713);
or U145 (N_145,In_844,In_69);
and U146 (N_146,In_1218,In_1471);
xor U147 (N_147,In_117,In_597);
xnor U148 (N_148,In_366,In_261);
or U149 (N_149,In_718,In_943);
or U150 (N_150,In_1477,N_41);
nand U151 (N_151,In_1354,In_1155);
xnor U152 (N_152,In_493,N_103);
or U153 (N_153,In_123,In_475);
or U154 (N_154,In_503,In_316);
and U155 (N_155,In_49,In_980);
and U156 (N_156,N_148,N_63);
or U157 (N_157,In_1327,In_99);
xor U158 (N_158,In_1168,In_1478);
xnor U159 (N_159,In_667,In_1317);
and U160 (N_160,In_165,In_86);
or U161 (N_161,In_48,In_157);
or U162 (N_162,In_996,In_947);
and U163 (N_163,In_1016,In_927);
or U164 (N_164,In_953,In_1381);
xnor U165 (N_165,In_826,In_32);
or U166 (N_166,In_1133,In_702);
xnor U167 (N_167,N_121,In_307);
and U168 (N_168,N_19,In_1487);
or U169 (N_169,In_170,In_349);
nand U170 (N_170,In_1257,In_835);
or U171 (N_171,In_148,In_609);
xor U172 (N_172,In_1287,In_75);
nand U173 (N_173,In_146,In_458);
or U174 (N_174,In_136,In_671);
or U175 (N_175,N_22,In_787);
xor U176 (N_176,N_11,In_620);
nor U177 (N_177,In_442,In_749);
xnor U178 (N_178,N_82,In_579);
nand U179 (N_179,In_1179,In_336);
xor U180 (N_180,In_21,In_1093);
and U181 (N_181,In_865,In_863);
or U182 (N_182,In_398,In_282);
and U183 (N_183,In_1164,In_1250);
nand U184 (N_184,In_160,In_581);
or U185 (N_185,In_602,In_1048);
nand U186 (N_186,In_45,In_429);
nor U187 (N_187,In_1106,In_158);
nor U188 (N_188,N_144,In_1258);
nor U189 (N_189,In_1151,In_1346);
nand U190 (N_190,In_1062,In_1290);
and U191 (N_191,In_950,In_677);
nor U192 (N_192,In_738,In_1302);
and U193 (N_193,In_1314,In_1355);
nand U194 (N_194,In_1446,In_466);
xor U195 (N_195,N_79,In_96);
and U196 (N_196,In_1070,In_60);
nor U197 (N_197,In_385,In_1462);
and U198 (N_198,In_245,In_1071);
nand U199 (N_199,In_1343,In_1284);
nor U200 (N_200,In_1391,In_1134);
and U201 (N_201,N_110,N_67);
xor U202 (N_202,In_685,In_1154);
nand U203 (N_203,In_1260,In_1309);
nand U204 (N_204,In_1185,In_830);
nor U205 (N_205,In_938,In_1397);
nand U206 (N_206,In_211,In_256);
or U207 (N_207,In_382,In_345);
xor U208 (N_208,In_520,In_1010);
nand U209 (N_209,In_173,N_42);
and U210 (N_210,In_1376,N_27);
or U211 (N_211,In_1280,In_1173);
and U212 (N_212,In_1102,In_1057);
nand U213 (N_213,In_1254,In_348);
or U214 (N_214,In_972,In_1269);
and U215 (N_215,In_1347,In_1208);
nand U216 (N_216,In_930,In_169);
nor U217 (N_217,In_545,N_131);
nor U218 (N_218,In_1491,In_159);
xnor U219 (N_219,In_632,In_478);
and U220 (N_220,In_525,In_839);
nand U221 (N_221,In_156,In_703);
nor U222 (N_222,In_411,In_1403);
nor U223 (N_223,N_132,N_124);
or U224 (N_224,In_103,In_260);
xnor U225 (N_225,In_648,In_432);
and U226 (N_226,In_175,In_43);
or U227 (N_227,In_592,In_369);
xnor U228 (N_228,In_91,In_1195);
and U229 (N_229,In_1073,In_906);
xnor U230 (N_230,In_435,In_467);
xor U231 (N_231,In_1234,In_1069);
and U232 (N_232,In_19,In_303);
nor U233 (N_233,In_1484,In_1092);
and U234 (N_234,In_836,In_487);
nand U235 (N_235,In_986,In_900);
nand U236 (N_236,In_660,In_805);
nand U237 (N_237,In_1238,In_188);
and U238 (N_238,In_333,In_1103);
or U239 (N_239,In_1494,In_322);
or U240 (N_240,In_401,In_469);
and U241 (N_241,In_215,In_102);
or U242 (N_242,In_732,In_1095);
and U243 (N_243,In_918,N_128);
and U244 (N_244,In_639,In_1334);
and U245 (N_245,In_110,In_283);
nor U246 (N_246,In_777,In_386);
or U247 (N_247,In_1387,In_16);
xor U248 (N_248,In_507,In_881);
nor U249 (N_249,N_77,In_203);
nor U250 (N_250,In_1303,In_249);
or U251 (N_251,N_113,In_247);
xnor U252 (N_252,In_1360,In_720);
or U253 (N_253,In_276,In_494);
xor U254 (N_254,In_802,In_199);
nor U255 (N_255,In_1285,In_223);
and U256 (N_256,In_87,In_961);
nand U257 (N_257,In_238,In_1074);
xnor U258 (N_258,In_1085,In_1409);
nand U259 (N_259,In_1485,In_663);
or U260 (N_260,In_378,In_885);
xor U261 (N_261,In_978,In_569);
or U262 (N_262,In_945,In_1396);
or U263 (N_263,In_1204,In_1147);
xnor U264 (N_264,N_136,In_966);
or U265 (N_265,In_1081,In_482);
and U266 (N_266,In_449,In_987);
nor U267 (N_267,N_17,In_1452);
or U268 (N_268,In_666,In_187);
or U269 (N_269,In_852,N_101);
nor U270 (N_270,In_1169,In_190);
or U271 (N_271,In_1289,N_80);
nand U272 (N_272,In_662,In_884);
nand U273 (N_273,In_1051,In_786);
or U274 (N_274,In_874,In_687);
nand U275 (N_275,In_414,In_682);
or U276 (N_276,N_8,N_69);
nor U277 (N_277,In_614,In_1266);
nand U278 (N_278,In_1233,In_876);
or U279 (N_279,In_1316,In_528);
or U280 (N_280,In_1251,N_71);
nand U281 (N_281,In_1114,In_1413);
xnor U282 (N_282,In_1282,In_1278);
xor U283 (N_283,In_1330,N_140);
nor U284 (N_284,In_1050,In_793);
or U285 (N_285,In_285,In_856);
nand U286 (N_286,In_1454,In_858);
nor U287 (N_287,In_774,In_14);
xnor U288 (N_288,N_138,In_337);
nand U289 (N_289,In_1296,In_983);
or U290 (N_290,In_932,In_988);
and U291 (N_291,In_364,In_598);
nand U292 (N_292,In_745,In_794);
nor U293 (N_293,In_532,In_792);
or U294 (N_294,In_556,In_613);
nand U295 (N_295,In_1089,In_1273);
xnor U296 (N_296,N_44,In_1359);
nand U297 (N_297,In_1305,In_1398);
or U298 (N_298,In_179,In_363);
and U299 (N_299,In_250,In_318);
or U300 (N_300,In_924,In_960);
and U301 (N_301,In_1207,N_187);
nand U302 (N_302,In_486,N_297);
nor U303 (N_303,In_1108,In_755);
nand U304 (N_304,In_1227,In_153);
and U305 (N_305,In_1006,In_167);
and U306 (N_306,In_763,N_24);
or U307 (N_307,N_141,In_834);
nand U308 (N_308,In_120,In_595);
and U309 (N_309,In_815,In_1439);
nand U310 (N_310,N_97,In_58);
nor U311 (N_311,N_236,In_731);
xnor U312 (N_312,In_11,In_1324);
and U313 (N_313,N_200,In_1038);
and U314 (N_314,In_1460,In_908);
or U315 (N_315,In_704,In_1239);
nor U316 (N_316,In_574,In_221);
nor U317 (N_317,N_206,In_191);
nor U318 (N_318,In_197,N_20);
or U319 (N_319,N_275,In_1249);
nand U320 (N_320,In_1193,In_390);
and U321 (N_321,In_1128,In_672);
and U322 (N_322,In_756,In_717);
nand U323 (N_323,In_1120,In_1063);
nor U324 (N_324,In_1420,In_1440);
xor U325 (N_325,N_133,In_737);
and U326 (N_326,In_1165,In_829);
xor U327 (N_327,In_940,N_219);
xor U328 (N_328,In_559,N_231);
nor U329 (N_329,In_575,In_931);
or U330 (N_330,In_1110,In_1277);
nand U331 (N_331,In_470,In_88);
nand U332 (N_332,In_825,In_174);
nand U333 (N_333,In_441,In_751);
nor U334 (N_334,In_1344,In_566);
and U335 (N_335,In_656,In_433);
xor U336 (N_336,In_361,N_4);
or U337 (N_337,N_250,In_402);
xnor U338 (N_338,In_107,In_371);
or U339 (N_339,In_812,In_1472);
xnor U340 (N_340,N_243,In_1205);
or U341 (N_341,N_58,N_48);
nand U342 (N_342,In_66,In_29);
or U343 (N_343,In_331,In_1252);
or U344 (N_344,In_910,In_1122);
and U345 (N_345,In_693,N_130);
nor U346 (N_346,In_649,In_306);
nor U347 (N_347,In_1039,In_857);
and U348 (N_348,In_129,In_25);
nand U349 (N_349,N_86,In_1490);
xnor U350 (N_350,N_93,In_1187);
xor U351 (N_351,In_1281,N_232);
or U352 (N_352,In_287,N_279);
nand U353 (N_353,In_324,In_286);
nand U354 (N_354,N_95,In_1237);
xor U355 (N_355,N_92,In_894);
and U356 (N_356,N_254,N_298);
xor U357 (N_357,In_530,In_809);
or U358 (N_358,In_1220,N_234);
or U359 (N_359,N_245,N_246);
nand U360 (N_360,N_106,In_1067);
nand U361 (N_361,In_1184,In_1437);
and U362 (N_362,In_28,In_1053);
xor U363 (N_363,N_51,In_76);
and U364 (N_364,In_646,In_959);
nor U365 (N_365,In_801,In_1131);
xor U366 (N_366,N_199,In_355);
nor U367 (N_367,In_358,In_1421);
nor U368 (N_368,In_320,N_278);
nand U369 (N_369,In_90,N_56);
nor U370 (N_370,In_241,In_998);
nand U371 (N_371,In_813,In_531);
or U372 (N_372,In_186,In_1363);
and U373 (N_373,In_1209,In_747);
and U374 (N_374,In_396,In_694);
or U375 (N_375,In_1153,In_1339);
and U376 (N_376,In_919,In_1389);
nand U377 (N_377,In_1024,In_420);
nand U378 (N_378,N_115,In_3);
and U379 (N_379,In_529,N_76);
nand U380 (N_380,In_1253,In_243);
and U381 (N_381,In_266,In_1127);
or U382 (N_382,N_126,In_1322);
or U383 (N_383,In_108,In_784);
or U384 (N_384,In_554,In_116);
nor U385 (N_385,In_1366,In_384);
nand U386 (N_386,In_985,In_1283);
nor U387 (N_387,In_1293,In_1467);
xnor U388 (N_388,In_1451,In_119);
or U389 (N_389,In_828,N_226);
nor U390 (N_390,In_213,In_4);
nor U391 (N_391,In_1210,In_50);
or U392 (N_392,In_430,In_1274);
nor U393 (N_393,In_889,In_481);
xnor U394 (N_394,In_740,In_109);
nand U395 (N_395,In_1028,In_867);
nand U396 (N_396,In_714,N_194);
xnor U397 (N_397,In_1497,In_549);
nor U398 (N_398,In_1142,N_129);
xnor U399 (N_399,In_903,In_1457);
and U400 (N_400,In_659,In_501);
xnor U401 (N_401,N_114,In_1453);
xnor U402 (N_402,In_969,In_615);
nand U403 (N_403,N_107,In_1152);
and U404 (N_404,In_172,In_541);
and U405 (N_405,N_185,N_213);
xnor U406 (N_406,In_754,In_608);
and U407 (N_407,In_201,In_1160);
nor U408 (N_408,In_684,In_1441);
and U409 (N_409,In_782,In_1111);
nand U410 (N_410,In_71,In_10);
xor U411 (N_411,In_214,N_3);
and U412 (N_412,N_258,In_779);
nor U413 (N_413,N_36,In_1431);
xor U414 (N_414,In_977,In_819);
and U415 (N_415,In_59,In_1395);
or U416 (N_416,In_821,N_293);
and U417 (N_417,In_730,In_122);
xnor U418 (N_418,N_5,N_192);
nand U419 (N_419,In_1007,In_853);
nand U420 (N_420,N_125,In_790);
nand U421 (N_421,In_8,N_21);
xnor U422 (N_422,In_572,In_1026);
or U423 (N_423,N_251,In_504);
and U424 (N_424,In_216,In_1476);
or U425 (N_425,In_93,In_1447);
xor U426 (N_426,In_645,N_74);
xor U427 (N_427,N_268,In_1270);
nand U428 (N_428,In_1056,In_1052);
or U429 (N_429,In_1196,In_891);
and U430 (N_430,In_657,In_1267);
nor U431 (N_431,In_1117,In_39);
xor U432 (N_432,In_255,In_1166);
nor U433 (N_433,In_417,N_55);
and U434 (N_434,In_412,N_183);
xnor U435 (N_435,In_1012,In_1348);
or U436 (N_436,N_256,N_255);
and U437 (N_437,In_599,N_81);
nor U438 (N_438,In_971,In_1143);
and U439 (N_439,In_421,In_612);
or U440 (N_440,In_368,N_225);
and U441 (N_441,In_642,N_83);
xor U442 (N_442,In_302,In_606);
nand U443 (N_443,In_1259,In_1394);
and U444 (N_444,In_523,In_140);
or U445 (N_445,In_1003,In_1374);
and U446 (N_446,In_1109,In_403);
or U447 (N_447,In_818,In_1276);
nand U448 (N_448,In_1401,In_1406);
xor U449 (N_449,In_177,In_6);
xnor U450 (N_450,In_850,N_338);
xor U451 (N_451,In_463,In_1023);
or U452 (N_452,In_288,In_413);
xnor U453 (N_453,N_330,In_708);
nor U454 (N_454,In_1345,In_1264);
nand U455 (N_455,In_899,N_409);
nor U456 (N_456,In_621,In_1482);
nand U457 (N_457,N_168,In_1393);
or U458 (N_458,N_64,In_1473);
and U459 (N_459,N_259,In_1104);
or U460 (N_460,N_224,In_80);
xnor U461 (N_461,In_410,In_1100);
xnor U462 (N_462,In_1342,In_851);
xnor U463 (N_463,N_377,In_305);
nor U464 (N_464,In_1219,N_160);
or U465 (N_465,N_413,In_1318);
nand U466 (N_466,N_173,N_318);
and U467 (N_467,N_260,In_1146);
and U468 (N_468,N_431,N_156);
xor U469 (N_469,In_974,In_465);
nand U470 (N_470,In_133,In_1336);
and U471 (N_471,In_1004,N_421);
nor U472 (N_472,In_1247,N_379);
nor U473 (N_473,In_105,In_1310);
and U474 (N_474,In_1094,In_590);
nor U475 (N_475,N_283,N_257);
xnor U476 (N_476,In_877,In_299);
xnor U477 (N_477,N_414,In_15);
nor U478 (N_478,N_145,N_274);
and U479 (N_479,In_518,In_1079);
xor U480 (N_480,In_444,N_347);
or U481 (N_481,In_675,N_439);
nand U482 (N_482,In_9,In_1001);
nor U483 (N_483,In_81,In_248);
or U484 (N_484,In_1045,N_50);
nor U485 (N_485,N_122,In_84);
or U486 (N_486,N_390,N_301);
or U487 (N_487,In_244,In_1235);
and U488 (N_488,N_449,In_778);
and U489 (N_489,N_367,In_1194);
xnor U490 (N_490,In_145,In_357);
nor U491 (N_491,In_601,In_451);
xnor U492 (N_492,N_176,In_1174);
nor U493 (N_493,In_750,In_128);
and U494 (N_494,In_695,N_429);
or U495 (N_495,N_87,In_452);
or U496 (N_496,N_262,N_123);
and U497 (N_497,N_209,In_1271);
xor U498 (N_498,In_335,In_1436);
or U499 (N_499,N_385,N_159);
and U500 (N_500,In_997,In_797);
and U501 (N_501,In_769,N_357);
and U502 (N_502,In_799,N_369);
xor U503 (N_503,In_143,N_33);
and U504 (N_504,N_32,In_933);
and U505 (N_505,In_1025,N_350);
nor U506 (N_506,N_389,N_428);
xnor U507 (N_507,N_228,In_630);
nor U508 (N_508,In_325,N_117);
or U509 (N_509,In_773,In_150);
nor U510 (N_510,In_394,N_370);
or U511 (N_511,In_1435,In_139);
nor U512 (N_512,In_1263,In_1407);
or U513 (N_513,In_719,In_729);
nor U514 (N_514,In_710,In_538);
and U515 (N_515,In_65,In_1084);
and U516 (N_516,In_416,N_52);
nand U517 (N_517,In_697,In_227);
xor U518 (N_518,In_623,N_374);
and U519 (N_519,In_1132,In_1382);
nand U520 (N_520,N_31,In_92);
nor U521 (N_521,N_170,In_328);
nand U522 (N_522,In_604,In_499);
xnor U523 (N_523,In_534,In_1211);
xor U524 (N_524,N_142,In_1226);
and U525 (N_525,N_402,In_1113);
nor U526 (N_526,In_97,N_334);
and U527 (N_527,In_1466,In_669);
nand U528 (N_528,In_329,N_443);
and U529 (N_529,N_204,In_166);
nor U530 (N_530,In_807,N_363);
nor U531 (N_531,N_437,N_269);
or U532 (N_532,N_175,N_337);
or U533 (N_533,In_26,N_382);
nor U534 (N_534,In_678,In_1337);
xor U535 (N_535,In_949,N_433);
xnor U536 (N_536,In_1357,In_397);
nor U537 (N_537,In_593,In_946);
and U538 (N_538,N_102,In_164);
nand U539 (N_539,N_47,In_1378);
nor U540 (N_540,N_342,In_1306);
nor U541 (N_541,In_1115,In_114);
or U542 (N_542,In_1096,In_1315);
nand U543 (N_543,In_17,In_1170);
nand U544 (N_544,In_496,In_1301);
nor U545 (N_545,In_1390,In_871);
and U546 (N_546,N_373,In_447);
nor U547 (N_547,N_13,N_394);
and U548 (N_548,In_880,In_1107);
or U549 (N_549,In_1216,N_94);
or U550 (N_550,In_224,N_99);
nand U551 (N_551,In_163,N_18);
and U552 (N_552,In_600,In_1031);
nor U553 (N_553,In_981,N_16);
or U554 (N_554,In_434,N_358);
or U555 (N_555,In_131,In_1042);
and U556 (N_556,In_618,In_1499);
nor U557 (N_557,In_111,N_35);
and U558 (N_558,In_741,In_301);
and U559 (N_559,In_827,N_184);
xnor U560 (N_560,In_1369,N_150);
and U561 (N_561,In_896,N_100);
nor U562 (N_562,N_38,In_905);
nand U563 (N_563,In_548,In_1125);
or U564 (N_564,N_420,In_419);
or U565 (N_565,In_1116,In_1443);
or U566 (N_566,In_423,In_1149);
or U567 (N_567,In_991,N_165);
nor U568 (N_568,N_205,In_901);
nor U569 (N_569,N_440,N_91);
xor U570 (N_570,In_1240,N_57);
nand U571 (N_571,In_343,N_271);
and U572 (N_572,N_25,In_1279);
and U573 (N_573,N_221,In_405);
xnor U574 (N_574,In_1183,In_281);
nor U575 (N_575,N_45,In_437);
nand U576 (N_576,In_1144,In_688);
xnor U577 (N_577,In_898,N_127);
nor U578 (N_578,In_1424,In_775);
or U579 (N_579,In_471,In_393);
nand U580 (N_580,In_272,In_263);
nand U581 (N_581,N_359,N_354);
nand U582 (N_582,In_654,In_1018);
nand U583 (N_583,N_432,In_1430);
or U584 (N_584,In_1030,N_137);
or U585 (N_585,N_120,In_607);
and U586 (N_586,N_248,N_418);
xor U587 (N_587,In_824,In_274);
xor U588 (N_588,N_410,N_376);
nor U589 (N_589,In_218,In_326);
nor U590 (N_590,N_177,In_273);
or U591 (N_591,In_490,In_712);
or U592 (N_592,N_167,In_1231);
nor U593 (N_593,In_347,N_364);
and U594 (N_594,In_229,In_1265);
or U595 (N_595,N_240,N_261);
and U596 (N_596,In_560,In_149);
or U597 (N_597,In_690,In_1126);
and U598 (N_598,N_346,In_1400);
nand U599 (N_599,In_655,N_381);
xnor U600 (N_600,In_125,N_579);
nor U601 (N_601,In_1064,In_1129);
xnor U602 (N_602,In_1445,In_926);
nor U603 (N_603,N_445,N_588);
xnor U604 (N_604,N_284,In_744);
or U605 (N_605,In_500,In_1061);
nor U606 (N_606,In_55,N_332);
nand U607 (N_607,In_715,In_1135);
nand U608 (N_608,N_474,In_185);
nand U609 (N_609,In_733,N_352);
nand U610 (N_610,N_116,In_112);
nand U611 (N_611,In_154,In_144);
and U612 (N_612,In_438,In_1140);
or U613 (N_613,N_340,N_507);
nor U614 (N_614,N_263,In_882);
and U615 (N_615,In_1465,N_188);
xor U616 (N_616,In_251,In_1118);
nand U617 (N_617,N_223,N_496);
xor U618 (N_618,In_808,N_400);
nor U619 (N_619,N_527,In_200);
nor U620 (N_620,In_277,N_203);
nand U621 (N_621,N_49,In_533);
xor U622 (N_622,N_442,In_1002);
xor U623 (N_623,N_457,N_89);
and U624 (N_624,In_1320,N_405);
nor U625 (N_625,N_399,N_384);
or U626 (N_626,In_557,In_588);
nand U627 (N_627,N_387,N_344);
or U628 (N_628,N_201,N_155);
nor U629 (N_629,In_234,In_596);
or U630 (N_630,In_817,In_1405);
or U631 (N_631,In_78,N_191);
and U632 (N_632,N_589,N_302);
or U633 (N_633,N_584,N_554);
nand U634 (N_634,In_958,In_1297);
nand U635 (N_635,N_451,N_522);
nor U636 (N_636,In_861,N_478);
nor U637 (N_637,In_1141,In_576);
or U638 (N_638,N_244,N_595);
xor U639 (N_639,In_643,In_230);
xor U640 (N_640,In_1191,In_1176);
xnor U641 (N_641,N_375,In_776);
and U642 (N_642,In_222,N_85);
or U643 (N_643,In_564,In_1458);
xnor U644 (N_644,In_543,In_1262);
nand U645 (N_645,In_1474,In_408);
nand U646 (N_646,N_172,In_664);
or U647 (N_647,In_1087,N_267);
and U648 (N_648,N_592,In_313);
nor U649 (N_649,N_12,N_537);
or U650 (N_650,In_130,N_90);
nand U651 (N_651,In_1410,In_944);
and U652 (N_652,In_94,N_467);
nand U653 (N_653,In_653,In_351);
or U654 (N_654,In_846,In_54);
and U655 (N_655,In_1434,N_178);
xor U656 (N_656,N_161,In_1172);
or U657 (N_657,N_490,In_36);
xnor U658 (N_658,In_791,N_465);
xor U659 (N_659,In_1217,In_975);
nor U660 (N_660,N_435,In_418);
xnor U661 (N_661,In_278,In_1161);
nor U662 (N_662,N_417,In_921);
nand U663 (N_663,N_135,In_1333);
or U664 (N_664,In_380,N_198);
or U665 (N_665,N_553,In_591);
nand U666 (N_666,N_247,In_297);
nand U667 (N_667,In_352,In_914);
or U668 (N_668,In_155,In_7);
xor U669 (N_669,N_563,In_661);
xor U670 (N_670,In_1275,In_635);
nand U671 (N_671,In_771,In_407);
nor U672 (N_672,N_307,N_543);
or U673 (N_673,In_1461,In_860);
xnor U674 (N_674,In_338,In_379);
xnor U675 (N_675,N_524,N_146);
and U676 (N_676,In_298,N_351);
and U677 (N_677,N_513,N_485);
nand U678 (N_678,In_670,N_109);
and U679 (N_679,In_67,In_1245);
nand U680 (N_680,In_1483,In_888);
xnor U681 (N_681,In_521,N_345);
nand U682 (N_682,N_174,N_530);
xnor U683 (N_683,N_570,In_1438);
nand U684 (N_684,In_1188,N_422);
nor U685 (N_685,In_810,In_262);
nor U686 (N_686,In_206,N_72);
and U687 (N_687,N_599,N_550);
or U688 (N_688,In_1090,N_587);
and U689 (N_689,In_770,N_575);
xor U690 (N_690,N_164,N_336);
and U691 (N_691,In_941,In_77);
and U692 (N_692,In_1256,N_586);
and U693 (N_693,N_419,N_324);
xnor U694 (N_694,N_516,N_6);
or U695 (N_695,In_1075,In_280);
nand U696 (N_696,N_61,In_424);
xor U697 (N_697,In_1414,In_1171);
nand U698 (N_698,N_310,N_574);
nand U699 (N_699,N_10,N_483);
nand U700 (N_700,N_40,N_415);
and U701 (N_701,N_134,In_300);
xnor U702 (N_702,In_788,N_551);
nand U703 (N_703,In_513,In_647);
and U704 (N_704,In_1077,In_583);
nand U705 (N_705,In_552,In_118);
or U706 (N_706,N_216,N_578);
xor U707 (N_707,N_555,N_458);
xnor U708 (N_708,In_1221,N_542);
nor U709 (N_709,N_66,N_386);
nor U710 (N_710,In_406,N_393);
or U711 (N_711,N_327,In_346);
and U712 (N_712,In_477,N_597);
nand U713 (N_713,N_572,In_209);
nand U714 (N_714,N_207,N_500);
nand U715 (N_715,In_459,N_493);
nor U716 (N_716,N_329,In_929);
or U717 (N_717,N_9,In_811);
nand U718 (N_718,N_406,In_425);
nor U719 (N_719,N_237,N_108);
nor U720 (N_720,N_463,N_482);
and U721 (N_721,In_676,In_1158);
or U722 (N_722,N_452,In_317);
or U723 (N_723,In_619,In_1384);
nand U724 (N_724,In_644,In_1181);
nand U725 (N_725,N_407,N_480);
xor U726 (N_726,N_147,In_168);
nand U727 (N_727,N_270,In_226);
nand U728 (N_728,N_538,N_403);
xor U729 (N_729,In_878,N_576);
nor U730 (N_730,In_1386,In_63);
xnor U731 (N_731,In_506,In_768);
and U732 (N_732,N_593,N_499);
or U733 (N_733,N_436,In_1020);
xor U734 (N_734,N_560,N_535);
and U735 (N_735,N_544,In_526);
nand U736 (N_736,In_804,In_370);
nor U737 (N_737,In_626,In_1399);
nor U738 (N_738,In_124,In_1288);
and U739 (N_739,N_179,N_65);
xor U740 (N_740,In_757,N_151);
nand U741 (N_741,In_753,In_820);
nand U742 (N_742,N_280,In_742);
nor U743 (N_743,In_1433,In_1034);
nor U744 (N_744,In_1429,N_580);
or U745 (N_745,N_596,N_37);
nor U746 (N_746,N_395,In_1365);
or U747 (N_747,N_398,N_378);
and U748 (N_748,In_957,In_527);
nand U749 (N_749,In_637,In_1294);
and U750 (N_750,N_692,N_469);
xnor U751 (N_751,In_409,N_96);
nor U752 (N_752,In_1076,N_717);
nand U753 (N_753,In_1099,In_445);
nor U754 (N_754,N_372,In_147);
or U755 (N_755,In_1223,In_1463);
xnor U756 (N_756,In_151,N_249);
nor U757 (N_757,N_652,N_713);
nand U758 (N_758,In_1379,In_1244);
and U759 (N_759,N_656,N_640);
and U760 (N_760,N_111,N_468);
nand U761 (N_761,N_272,In_1449);
or U762 (N_762,In_1225,N_497);
nor U763 (N_763,In_235,N_46);
nand U764 (N_764,In_377,N_654);
nand U765 (N_765,In_1083,In_517);
nand U766 (N_766,In_1308,N_612);
or U767 (N_767,N_660,N_309);
or U768 (N_768,N_546,In_859);
or U769 (N_769,N_470,In_580);
nand U770 (N_770,In_246,N_607);
xor U771 (N_771,In_1200,In_489);
nor U772 (N_772,N_171,In_1370);
or U773 (N_773,N_211,In_176);
and U774 (N_774,N_401,In_722);
nand U775 (N_775,In_309,N_558);
nand U776 (N_776,N_602,N_645);
nand U777 (N_777,N_392,N_627);
xor U778 (N_778,In_461,In_999);
or U779 (N_779,N_475,N_637);
nand U780 (N_780,In_462,N_649);
or U781 (N_781,In_1312,N_636);
nor U782 (N_782,N_313,In_734);
or U783 (N_783,N_677,N_210);
nor U784 (N_784,N_688,In_440);
and U785 (N_785,N_361,In_1377);
or U786 (N_786,N_28,In_296);
xnor U787 (N_787,N_139,N_635);
nor U788 (N_788,In_913,N_195);
xnor U789 (N_789,In_381,N_300);
nor U790 (N_790,N_720,N_642);
nor U791 (N_791,N_448,In_1480);
nor U792 (N_792,N_447,In_1325);
and U793 (N_793,In_795,In_389);
nand U794 (N_794,N_657,N_362);
xor U795 (N_795,In_1432,In_1417);
and U796 (N_796,N_239,N_634);
nor U797 (N_797,In_208,N_532);
nand U798 (N_798,In_1479,In_915);
xnor U799 (N_799,In_658,In_1425);
xor U800 (N_800,In_240,In_764);
nand U801 (N_801,In_1055,N_222);
nor U802 (N_802,N_630,In_253);
or U803 (N_803,N_738,N_529);
nor U804 (N_804,N_323,In_934);
nor U805 (N_805,N_719,N_696);
xor U806 (N_806,In_1072,N_504);
nor U807 (N_807,N_512,In_323);
nand U808 (N_808,N_557,N_647);
nand U809 (N_809,N_748,In_42);
nand U810 (N_810,N_711,In_340);
nor U811 (N_811,N_743,In_510);
nor U812 (N_812,N_722,In_994);
xor U813 (N_813,N_489,In_83);
xor U814 (N_814,In_1358,N_112);
and U815 (N_815,In_61,N_491);
or U816 (N_816,N_556,In_726);
and U817 (N_817,N_118,In_765);
or U818 (N_818,In_870,N_471);
nand U819 (N_819,In_1203,N_582);
nand U820 (N_820,N_631,N_541);
and U821 (N_821,N_119,N_411);
or U822 (N_822,In_558,N_287);
nand U823 (N_823,In_491,In_516);
nor U824 (N_824,In_1352,In_585);
nand U825 (N_825,N_565,N_321);
nor U826 (N_826,N_633,N_289);
or U827 (N_827,In_427,N_671);
nand U828 (N_828,N_545,In_698);
or U829 (N_829,N_208,In_886);
nand U830 (N_830,N_727,N_583);
nand U831 (N_831,N_320,In_137);
xor U832 (N_832,In_1175,In_232);
nand U833 (N_833,N_663,In_236);
nand U834 (N_834,In_85,In_1388);
or U835 (N_835,N_365,In_1021);
or U836 (N_836,In_651,N_477);
and U837 (N_837,N_189,In_73);
or U838 (N_838,N_739,N_526);
and U839 (N_839,N_157,N_88);
nand U840 (N_840,In_1335,N_314);
and U841 (N_841,In_304,N_326);
nand U842 (N_842,N_253,N_646);
and U843 (N_843,N_667,In_138);
nor U844 (N_844,N_650,In_383);
and U845 (N_845,N_430,N_653);
nand U846 (N_846,In_1041,N_721);
xor U847 (N_847,N_598,In_1404);
or U848 (N_848,In_202,N_644);
nor U849 (N_849,N_34,N_153);
xnor U850 (N_850,N_143,N_655);
xnor U851 (N_851,In_1198,N_679);
and U852 (N_852,N_105,In_1418);
xor U853 (N_853,N_355,In_823);
nor U854 (N_854,In_1455,N_651);
and U855 (N_855,In_1178,N_697);
and U856 (N_856,In_1416,N_476);
nor U857 (N_857,N_715,N_0);
xor U858 (N_858,N_517,In_743);
xor U859 (N_859,N_730,N_158);
and U860 (N_860,In_35,In_907);
xor U861 (N_861,In_217,N_495);
nand U862 (N_862,N_238,N_712);
nor U863 (N_863,N_661,N_408);
xor U864 (N_864,N_585,N_299);
nor U865 (N_865,N_624,In_310);
nand U866 (N_866,In_1489,N_368);
nand U867 (N_867,N_514,In_1013);
nand U868 (N_868,N_626,N_577);
xor U869 (N_869,N_230,In_617);
nor U870 (N_870,N_639,N_14);
and U871 (N_871,N_698,In_650);
or U872 (N_872,In_1298,N_594);
xor U873 (N_873,In_1080,In_542);
xnor U874 (N_874,N_723,N_525);
xor U875 (N_875,N_304,N_745);
or U876 (N_876,In_1036,In_1459);
and U877 (N_877,N_412,In_1078);
nand U878 (N_878,In_1,In_1496);
nor U879 (N_879,N_506,N_562);
nor U880 (N_880,In_759,N_60);
nor U881 (N_881,N_328,In_1272);
xnor U882 (N_882,N_423,In_404);
xnor U883 (N_883,N_462,In_892);
xor U884 (N_884,In_267,N_26);
nand U885 (N_885,In_360,N_424);
xor U886 (N_886,N_335,N_341);
and U887 (N_887,In_1372,In_72);
or U888 (N_888,In_762,N_193);
or U889 (N_889,N_39,N_252);
or U890 (N_890,In_979,In_27);
xor U891 (N_891,In_1268,In_162);
nor U892 (N_892,In_38,N_643);
and U893 (N_893,In_1214,N_734);
nor U894 (N_894,N_196,N_685);
and U895 (N_895,N_724,In_767);
nand U896 (N_896,In_456,N_687);
xnor U897 (N_897,In_319,N_43);
and U898 (N_898,In_976,N_59);
nand U899 (N_899,In_474,N_669);
nand U900 (N_900,N_515,N_30);
nor U901 (N_901,In_342,N_775);
xnor U902 (N_902,N_866,In_875);
and U903 (N_903,In_573,In_1448);
nand U904 (N_904,N_308,In_1498);
nor U905 (N_905,In_30,N_163);
nor U906 (N_906,N_750,In_937);
nor U907 (N_907,In_634,N_847);
and U908 (N_908,N_510,N_349);
xor U909 (N_909,In_1040,N_886);
xnor U910 (N_910,N_763,N_519);
or U911 (N_911,N_783,In_843);
and U912 (N_912,N_441,In_121);
nor U913 (N_913,N_735,In_1027);
and U914 (N_914,N_214,N_809);
nand U915 (N_915,N_528,N_862);
xor U916 (N_916,N_397,N_699);
and U917 (N_917,In_1047,In_1005);
and U918 (N_918,N_658,In_638);
or U919 (N_919,N_885,N_707);
nand U920 (N_920,N_695,In_570);
and U921 (N_921,N_804,N_678);
and U922 (N_922,In_629,N_852);
nor U923 (N_923,N_573,N_800);
or U924 (N_924,N_319,N_867);
nand U925 (N_925,N_152,In_1213);
or U926 (N_926,N_893,N_461);
and U927 (N_927,In_789,In_113);
nand U928 (N_928,N_533,In_1392);
and U929 (N_929,N_446,N_479);
and U930 (N_930,N_628,N_540);
nor U931 (N_931,In_1242,N_898);
nand U932 (N_932,N_737,N_670);
nand U933 (N_933,N_753,N_356);
and U934 (N_934,N_786,N_632);
or U935 (N_935,In_468,N_863);
or U936 (N_936,N_281,N_459);
nand U937 (N_937,In_864,N_241);
and U938 (N_938,In_1065,In_706);
nand U939 (N_939,In_415,N_625);
nor U940 (N_940,In_577,N_779);
nand U941 (N_941,N_68,N_825);
nand U942 (N_942,In_1145,N_831);
or U943 (N_943,N_566,N_166);
xor U944 (N_944,N_666,N_780);
and U945 (N_945,N_427,In_387);
xnor U946 (N_946,In_446,In_546);
and U947 (N_947,N_846,N_836);
nand U948 (N_948,N_896,In_683);
nand U949 (N_949,In_951,N_851);
nand U950 (N_950,In_439,N_870);
and U951 (N_951,N_860,N_149);
xnor U952 (N_952,In_627,N_772);
xnor U953 (N_953,In_399,N_778);
and U954 (N_954,N_787,N_371);
nand U955 (N_955,N_539,N_391);
nand U956 (N_956,N_684,In_180);
xor U957 (N_957,N_2,N_531);
nor U958 (N_958,N_600,In_563);
nor U959 (N_959,N_705,In_1385);
and U960 (N_960,N_444,In_1060);
or U961 (N_961,N_197,N_808);
or U962 (N_962,N_648,N_703);
nand U963 (N_963,In_631,N_759);
xnor U964 (N_964,In_954,N_826);
or U965 (N_965,N_841,In_1338);
and U966 (N_966,N_689,N_848);
nand U967 (N_967,N_186,N_850);
nor U968 (N_968,N_732,N_888);
nor U969 (N_969,In_1029,In_464);
nor U970 (N_970,N_590,In_476);
or U971 (N_971,In_840,N_857);
xnor U972 (N_972,N_162,N_868);
or U973 (N_973,N_686,N_810);
or U974 (N_974,N_736,In_56);
and U975 (N_975,N_726,N_315);
and U976 (N_976,In_822,In_681);
nor U977 (N_977,N_488,In_1419);
and U978 (N_978,N_606,N_294);
or U979 (N_979,N_460,In_22);
and U980 (N_980,N_815,N_521);
and U981 (N_981,N_548,In_993);
nand U982 (N_982,In_341,N_830);
and U983 (N_983,N_728,N_854);
or U984 (N_984,N_331,In_781);
nor U985 (N_985,N_523,N_455);
and U986 (N_986,N_725,N_789);
nor U987 (N_987,In_258,N_861);
nand U988 (N_988,N_871,N_1);
and U989 (N_989,N_892,N_807);
nand U990 (N_990,N_603,N_212);
xnor U991 (N_991,In_1248,In_1367);
or U992 (N_992,N_552,N_741);
and U993 (N_993,N_856,N_821);
and U994 (N_994,In_294,N_700);
nor U995 (N_995,N_561,In_184);
nand U996 (N_996,N_571,N_773);
nor U997 (N_997,In_127,N_305);
nand U998 (N_998,In_922,N_218);
or U999 (N_999,N_29,N_874);
nor U1000 (N_1000,N_858,N_306);
or U1001 (N_1001,In_916,N_822);
xnor U1002 (N_1002,N_348,N_708);
nand U1003 (N_1003,In_692,In_1137);
or U1004 (N_1004,N_761,N_615);
and U1005 (N_1005,N_680,N_784);
nor U1006 (N_1006,N_894,N_755);
nand U1007 (N_1007,N_774,N_758);
xor U1008 (N_1008,In_24,N_492);
nand U1009 (N_1009,In_1470,N_73);
and U1010 (N_1010,N_756,N_791);
nand U1011 (N_1011,In_436,N_292);
nand U1012 (N_1012,N_793,In_686);
nand U1013 (N_1013,In_1112,In_845);
and U1014 (N_1014,N_838,N_438);
and U1015 (N_1015,N_877,N_285);
nand U1016 (N_1016,N_675,N_731);
and U1017 (N_1017,N_54,N_383);
and U1018 (N_1018,In_1326,N_770);
and U1019 (N_1019,N_303,In_1412);
nand U1020 (N_1020,N_623,In_233);
or U1021 (N_1021,In_1255,In_134);
nor U1022 (N_1022,In_727,N_757);
or U1023 (N_1023,N_843,N_84);
xor U1024 (N_1024,In_1468,In_1189);
xnor U1025 (N_1025,In_327,N_505);
xor U1026 (N_1026,N_494,N_729);
nor U1027 (N_1027,In_568,N_353);
nand U1028 (N_1028,N_277,N_806);
or U1029 (N_1029,N_672,N_855);
nand U1030 (N_1030,In_1228,In_141);
and U1031 (N_1031,In_936,N_456);
nand U1032 (N_1032,In_1068,In_701);
nand U1033 (N_1033,N_62,In_761);
xnor U1034 (N_1034,N_805,N_508);
or U1035 (N_1035,In_259,In_1427);
nand U1036 (N_1036,In_0,N_618);
nand U1037 (N_1037,N_880,N_276);
or U1038 (N_1038,In_1101,N_534);
and U1039 (N_1039,N_747,N_875);
and U1040 (N_1040,N_266,N_690);
xor U1041 (N_1041,In_1138,In_1044);
or U1042 (N_1042,In_1349,N_288);
or U1043 (N_1043,In_1261,In_1353);
xnor U1044 (N_1044,N_453,N_454);
and U1045 (N_1045,In_772,N_742);
and U1046 (N_1046,N_853,In_535);
xnor U1047 (N_1047,N_714,In_833);
nand U1048 (N_1048,In_57,N_683);
or U1049 (N_1049,N_837,N_817);
or U1050 (N_1050,N_718,N_733);
nor U1051 (N_1051,N_933,N_1007);
and U1052 (N_1052,N_704,N_604);
and U1053 (N_1053,N_1021,N_1028);
or U1054 (N_1054,N_1002,N_1032);
nor U1055 (N_1055,N_937,N_920);
and U1056 (N_1056,N_501,N_339);
nand U1057 (N_1057,N_816,N_709);
nor U1058 (N_1058,N_864,N_946);
nand U1059 (N_1059,N_434,N_620);
nand U1060 (N_1060,N_1025,N_824);
nor U1061 (N_1061,N_569,N_662);
nor U1062 (N_1062,N_486,In_231);
or U1063 (N_1063,N_487,N_941);
nor U1064 (N_1064,In_51,N_963);
nand U1065 (N_1065,In_284,N_953);
xnor U1066 (N_1066,N_785,N_1035);
and U1067 (N_1067,N_609,N_991);
nand U1068 (N_1068,N_1004,N_986);
xnor U1069 (N_1069,In_547,N_1012);
nor U1070 (N_1070,In_372,In_1241);
nor U1071 (N_1071,N_601,N_619);
xnor U1072 (N_1072,N_999,N_547);
nand U1073 (N_1073,N_845,N_1037);
xor U1074 (N_1074,N_608,N_803);
or U1075 (N_1075,N_873,N_872);
or U1076 (N_1076,N_777,In_290);
xor U1077 (N_1077,N_360,N_882);
xnor U1078 (N_1078,In_1091,N_927);
nor U1079 (N_1079,N_520,N_273);
xnor U1080 (N_1080,In_624,N_1005);
and U1081 (N_1081,N_912,N_918);
and U1082 (N_1082,N_265,In_522);
nor U1083 (N_1083,N_682,In_848);
and U1084 (N_1084,N_1001,In_1224);
or U1085 (N_1085,In_132,N_790);
nor U1086 (N_1086,N_518,N_1011);
nor U1087 (N_1087,N_78,In_1351);
nor U1088 (N_1088,N_988,N_311);
nor U1089 (N_1089,N_629,N_316);
nand U1090 (N_1090,N_1017,In_428);
xnor U1091 (N_1091,N_70,N_884);
xnor U1092 (N_1092,N_23,N_290);
or U1093 (N_1093,In_553,N_827);
or U1094 (N_1094,N_814,In_1156);
xnor U1095 (N_1095,N_614,N_1008);
or U1096 (N_1096,N_952,N_1039);
xnor U1097 (N_1097,N_954,N_881);
or U1098 (N_1098,In_1201,In_70);
xnor U1099 (N_1099,N_710,N_818);
nand U1100 (N_1100,N_559,N_992);
nand U1101 (N_1101,N_844,N_749);
nor U1102 (N_1102,N_691,In_455);
and U1103 (N_1103,N_1014,N_1047);
nor U1104 (N_1104,N_878,N_53);
xor U1105 (N_1105,N_940,N_865);
nor U1106 (N_1106,In_1408,In_691);
nor U1107 (N_1107,N_902,In_2);
nand U1108 (N_1108,N_1024,N_802);
and U1109 (N_1109,N_776,In_485);
nand U1110 (N_1110,N_829,N_1029);
nand U1111 (N_1111,N_1033,N_969);
xor U1112 (N_1112,In_101,In_367);
nor U1113 (N_1113,In_1046,N_674);
or U1114 (N_1114,N_1016,In_841);
and U1115 (N_1115,N_928,N_970);
or U1116 (N_1116,N_922,N_976);
nor U1117 (N_1117,N_1044,N_1034);
nor U1118 (N_1118,N_233,In_350);
nor U1119 (N_1119,N_956,N_484);
or U1120 (N_1120,In_204,N_766);
and U1121 (N_1121,N_503,N_1049);
nor U1122 (N_1122,N_549,N_978);
xnor U1123 (N_1123,N_693,N_910);
xor U1124 (N_1124,N_621,N_75);
nor U1125 (N_1125,N_1015,N_799);
nor U1126 (N_1126,N_968,N_229);
nand U1127 (N_1127,N_989,N_380);
and U1128 (N_1128,N_1042,N_765);
xor U1129 (N_1129,N_931,N_312);
xor U1130 (N_1130,N_904,N_502);
nor U1131 (N_1131,N_819,In_855);
or U1132 (N_1132,N_744,N_955);
nor U1133 (N_1133,In_1329,N_202);
and U1134 (N_1134,N_796,N_716);
xnor U1135 (N_1135,In_219,In_1119);
nand U1136 (N_1136,N_794,N_567);
nand U1137 (N_1137,N_833,N_426);
and U1138 (N_1138,N_974,N_938);
and U1139 (N_1139,N_917,N_664);
and U1140 (N_1140,N_1020,N_1010);
and U1141 (N_1141,N_915,N_769);
nand U1142 (N_1142,N_859,N_820);
nand U1143 (N_1143,N_767,N_668);
nand U1144 (N_1144,N_181,N_842);
nand U1145 (N_1145,In_970,N_983);
or U1146 (N_1146,N_591,In_636);
or U1147 (N_1147,N_887,In_587);
nand U1148 (N_1148,N_98,N_936);
nand U1149 (N_1149,N_581,N_984);
nor U1150 (N_1150,N_975,N_616);
and U1151 (N_1151,N_925,N_900);
and U1152 (N_1152,N_388,N_665);
or U1153 (N_1153,N_638,In_890);
and U1154 (N_1154,N_1048,N_673);
and U1155 (N_1155,In_1037,N_169);
nand U1156 (N_1156,In_1150,N_641);
xnor U1157 (N_1157,In_376,N_985);
nor U1158 (N_1158,N_932,N_811);
or U1159 (N_1159,In_505,N_264);
and U1160 (N_1160,N_1031,N_1013);
xnor U1161 (N_1161,In_711,N_994);
and U1162 (N_1162,N_1026,In_375);
nor U1163 (N_1163,N_322,N_869);
nor U1164 (N_1164,N_823,N_1023);
xnor U1165 (N_1165,N_568,N_622);
and U1166 (N_1166,In_832,In_1054);
nor U1167 (N_1167,In_668,N_472);
nand U1168 (N_1168,N_180,In_18);
and U1169 (N_1169,In_942,N_325);
or U1170 (N_1170,N_182,N_740);
nand U1171 (N_1171,N_950,In_448);
or U1172 (N_1172,N_934,In_1097);
nand U1173 (N_1173,N_366,N_1030);
and U1174 (N_1174,N_1018,N_849);
and U1175 (N_1175,In_1014,In_1015);
xor U1176 (N_1176,N_1019,N_981);
nor U1177 (N_1177,N_1040,N_286);
and U1178 (N_1178,N_295,N_966);
nand U1179 (N_1179,N_1006,N_813);
xnor U1180 (N_1180,In_1043,N_980);
and U1181 (N_1181,N_960,N_993);
xor U1182 (N_1182,N_235,N_909);
and U1183 (N_1183,N_1009,N_746);
or U1184 (N_1184,N_701,N_903);
or U1185 (N_1185,In_353,N_923);
or U1186 (N_1186,N_883,In_40);
and U1187 (N_1187,N_613,N_990);
or U1188 (N_1188,N_1038,N_425);
nand U1189 (N_1189,In_1292,N_997);
and U1190 (N_1190,In_679,N_943);
and U1191 (N_1191,In_904,In_1236);
xnor U1192 (N_1192,N_466,N_536);
and U1193 (N_1193,N_876,N_901);
xor U1194 (N_1194,N_924,N_752);
or U1195 (N_1195,N_1027,N_1036);
nor U1196 (N_1196,N_771,N_899);
or U1197 (N_1197,N_220,N_913);
xor U1198 (N_1198,N_919,N_788);
xnor U1199 (N_1199,N_908,N_926);
or U1200 (N_1200,N_1051,N_1111);
xnor U1201 (N_1201,N_1052,N_1136);
nor U1202 (N_1202,N_1119,N_959);
and U1203 (N_1203,N_1122,N_1058);
xnor U1204 (N_1204,N_481,N_1130);
and U1205 (N_1205,N_1169,N_751);
xor U1206 (N_1206,N_1197,N_1066);
xor U1207 (N_1207,N_1022,N_916);
nor U1208 (N_1208,N_1061,N_450);
xnor U1209 (N_1209,N_982,N_1141);
xor U1210 (N_1210,N_1182,N_1164);
xor U1211 (N_1211,N_702,N_1153);
or U1212 (N_1212,N_971,N_1163);
xnor U1213 (N_1213,In_257,In_1130);
xnor U1214 (N_1214,In_982,N_1134);
nand U1215 (N_1215,In_551,N_1112);
nor U1216 (N_1216,N_1188,N_929);
nand U1217 (N_1217,In_34,N_828);
nand U1218 (N_1218,In_928,N_935);
nor U1219 (N_1219,N_681,N_1177);
or U1220 (N_1220,N_972,N_1181);
xor U1221 (N_1221,N_1180,N_832);
and U1222 (N_1222,N_1059,N_1057);
nor U1223 (N_1223,N_1062,N_1093);
xor U1224 (N_1224,N_1077,N_812);
nor U1225 (N_1225,N_1199,N_1135);
nand U1226 (N_1226,N_1102,N_1100);
and U1227 (N_1227,N_1192,N_768);
xor U1228 (N_1228,N_1138,In_1105);
and U1229 (N_1229,N_227,N_798);
nor U1230 (N_1230,N_948,N_659);
nand U1231 (N_1231,N_1137,N_1157);
or U1232 (N_1232,N_676,N_1127);
and U1233 (N_1233,In_1180,In_275);
xnor U1234 (N_1234,N_343,N_905);
nor U1235 (N_1235,N_1056,N_1091);
nand U1236 (N_1236,In_1243,In_1049);
xor U1237 (N_1237,N_404,In_1058);
and U1238 (N_1238,N_1098,N_754);
nor U1239 (N_1239,N_694,N_1184);
nor U1240 (N_1240,N_416,N_792);
nand U1241 (N_1241,In_354,N_762);
xnor U1242 (N_1242,N_511,N_1145);
or U1243 (N_1243,N_942,N_1089);
or U1244 (N_1244,N_1106,N_1174);
and U1245 (N_1245,N_965,N_1160);
nand U1246 (N_1246,N_1190,N_242);
nor U1247 (N_1247,In_1442,N_977);
or U1248 (N_1248,N_1120,N_706);
nor U1249 (N_1249,N_879,N_215);
nand U1250 (N_1250,In_746,N_944);
nor U1251 (N_1251,In_511,N_1083);
or U1252 (N_1252,In_862,In_1307);
or U1253 (N_1253,N_949,N_961);
or U1254 (N_1254,N_396,N_797);
and U1255 (N_1255,N_760,N_1079);
and U1256 (N_1256,N_1173,N_104);
xor U1257 (N_1257,N_1139,N_1183);
or U1258 (N_1258,N_1176,N_1069);
nand U1259 (N_1259,N_1175,N_1196);
xnor U1260 (N_1260,N_610,In_641);
nand U1261 (N_1261,In_5,N_979);
nand U1262 (N_1262,N_1150,In_1162);
xnor U1263 (N_1263,N_1148,N_1179);
and U1264 (N_1264,N_1115,N_1156);
nand U1265 (N_1265,N_1178,N_795);
xnor U1266 (N_1266,N_1114,In_1212);
nor U1267 (N_1267,N_1159,N_1082);
nor U1268 (N_1268,N_1113,N_1118);
nor U1269 (N_1269,N_1107,N_1152);
nand U1270 (N_1270,N_1073,N_964);
and U1271 (N_1271,N_1129,N_890);
or U1272 (N_1272,N_1084,N_1158);
and U1273 (N_1273,N_906,N_1165);
nor U1274 (N_1274,N_1124,N_1195);
or U1275 (N_1275,N_835,N_914);
and U1276 (N_1276,N_317,N_1000);
and U1277 (N_1277,N_1123,N_1076);
nor U1278 (N_1278,N_1090,N_1101);
and U1279 (N_1279,N_1104,N_1094);
and U1280 (N_1280,In_1295,N_1133);
and U1281 (N_1281,N_1168,N_1193);
xor U1282 (N_1282,N_15,N_564);
and U1283 (N_1283,In_492,N_190);
and U1284 (N_1284,N_895,N_1041);
nand U1285 (N_1285,N_1161,N_1063);
or U1286 (N_1286,N_1096,N_154);
xnor U1287 (N_1287,N_1045,N_1085);
nor U1288 (N_1288,N_840,N_1110);
and U1289 (N_1289,N_945,N_1053);
xnor U1290 (N_1290,N_781,N_1081);
xor U1291 (N_1291,N_1054,N_967);
xnor U1292 (N_1292,In_182,N_1172);
and U1293 (N_1293,N_1167,N_907);
or U1294 (N_1294,In_365,N_1087);
and U1295 (N_1295,N_1055,In_515);
nor U1296 (N_1296,N_1171,In_269);
xnor U1297 (N_1297,In_264,N_973);
xnor U1298 (N_1298,N_611,N_1060);
or U1299 (N_1299,N_1185,N_509);
and U1300 (N_1300,N_473,N_1108);
nand U1301 (N_1301,N_1128,N_1154);
xnor U1302 (N_1302,N_1003,N_217);
xnor U1303 (N_1303,N_782,N_995);
xnor U1304 (N_1304,In_192,N_1065);
nand U1305 (N_1305,N_801,N_957);
xor U1306 (N_1306,N_962,N_1099);
nor U1307 (N_1307,N_921,N_1149);
and U1308 (N_1308,N_1071,N_891);
and U1309 (N_1309,N_291,In_1159);
and U1310 (N_1310,N_1125,In_332);
or U1311 (N_1311,N_1068,N_1050);
and U1312 (N_1312,N_1078,N_839);
nand U1313 (N_1313,N_1103,N_1126);
xnor U1314 (N_1314,N_951,N_1043);
or U1315 (N_1315,N_958,N_7);
xnor U1316 (N_1316,In_460,N_1070);
or U1317 (N_1317,In_748,In_616);
xnor U1318 (N_1318,N_1086,N_1121);
nor U1319 (N_1319,N_764,N_617);
and U1320 (N_1320,N_1155,N_1074);
nand U1321 (N_1321,N_1166,N_498);
or U1322 (N_1322,N_1191,N_282);
nor U1323 (N_1323,N_1170,N_1186);
and U1324 (N_1324,N_1046,N_1143);
nand U1325 (N_1325,N_930,N_1189);
or U1326 (N_1326,In_866,N_889);
and U1327 (N_1327,N_1095,N_1151);
and U1328 (N_1328,N_939,N_911);
xnor U1329 (N_1329,N_1080,In_228);
nand U1330 (N_1330,N_1144,In_920);
xnor U1331 (N_1331,N_1146,N_1075);
nor U1332 (N_1332,In_239,N_1117);
or U1333 (N_1333,N_1198,N_1067);
xnor U1334 (N_1334,N_1140,N_1109);
or U1335 (N_1335,N_998,In_1011);
and U1336 (N_1336,In_611,N_1116);
nand U1337 (N_1337,N_1147,N_996);
xnor U1338 (N_1338,N_464,N_1092);
and U1339 (N_1339,In_739,N_1142);
or U1340 (N_1340,N_296,N_1194);
or U1341 (N_1341,N_1088,N_1072);
nand U1342 (N_1342,In_237,N_1097);
or U1343 (N_1343,N_1064,N_1132);
nand U1344 (N_1344,N_1131,N_1187);
nor U1345 (N_1345,In_64,N_987);
and U1346 (N_1346,N_897,N_834);
and U1347 (N_1347,N_1162,N_605);
xor U1348 (N_1348,N_333,In_1232);
nor U1349 (N_1349,N_1105,N_947);
or U1350 (N_1350,N_1206,N_1339);
or U1351 (N_1351,N_1228,N_1313);
nand U1352 (N_1352,N_1265,N_1215);
and U1353 (N_1353,N_1260,N_1242);
nor U1354 (N_1354,N_1305,N_1200);
nand U1355 (N_1355,N_1327,N_1315);
or U1356 (N_1356,N_1311,N_1272);
or U1357 (N_1357,N_1329,N_1271);
or U1358 (N_1358,N_1309,N_1322);
nand U1359 (N_1359,N_1247,N_1273);
xnor U1360 (N_1360,N_1253,N_1285);
and U1361 (N_1361,N_1238,N_1204);
or U1362 (N_1362,N_1258,N_1331);
or U1363 (N_1363,N_1297,N_1347);
nand U1364 (N_1364,N_1320,N_1341);
nor U1365 (N_1365,N_1240,N_1230);
xnor U1366 (N_1366,N_1284,N_1303);
and U1367 (N_1367,N_1274,N_1223);
nand U1368 (N_1368,N_1268,N_1301);
or U1369 (N_1369,N_1296,N_1254);
nand U1370 (N_1370,N_1278,N_1318);
and U1371 (N_1371,N_1293,N_1333);
nor U1372 (N_1372,N_1244,N_1257);
nor U1373 (N_1373,N_1289,N_1344);
xor U1374 (N_1374,N_1335,N_1226);
or U1375 (N_1375,N_1312,N_1263);
nand U1376 (N_1376,N_1340,N_1342);
and U1377 (N_1377,N_1276,N_1245);
and U1378 (N_1378,N_1207,N_1237);
and U1379 (N_1379,N_1270,N_1349);
or U1380 (N_1380,N_1234,N_1299);
nand U1381 (N_1381,N_1222,N_1279);
nand U1382 (N_1382,N_1203,N_1323);
or U1383 (N_1383,N_1255,N_1298);
nor U1384 (N_1384,N_1235,N_1209);
nor U1385 (N_1385,N_1307,N_1211);
nand U1386 (N_1386,N_1267,N_1231);
nor U1387 (N_1387,N_1283,N_1214);
or U1388 (N_1388,N_1287,N_1261);
or U1389 (N_1389,N_1337,N_1256);
xor U1390 (N_1390,N_1308,N_1330);
and U1391 (N_1391,N_1205,N_1275);
xor U1392 (N_1392,N_1219,N_1332);
or U1393 (N_1393,N_1325,N_1227);
xor U1394 (N_1394,N_1236,N_1233);
nand U1395 (N_1395,N_1225,N_1294);
xor U1396 (N_1396,N_1282,N_1251);
nand U1397 (N_1397,N_1232,N_1210);
xnor U1398 (N_1398,N_1201,N_1280);
and U1399 (N_1399,N_1224,N_1262);
nor U1400 (N_1400,N_1310,N_1212);
nor U1401 (N_1401,N_1292,N_1248);
or U1402 (N_1402,N_1213,N_1288);
xor U1403 (N_1403,N_1259,N_1345);
nand U1404 (N_1404,N_1250,N_1269);
xor U1405 (N_1405,N_1295,N_1338);
nor U1406 (N_1406,N_1202,N_1208);
nand U1407 (N_1407,N_1328,N_1334);
and U1408 (N_1408,N_1321,N_1348);
or U1409 (N_1409,N_1252,N_1302);
nor U1410 (N_1410,N_1317,N_1304);
xor U1411 (N_1411,N_1343,N_1220);
and U1412 (N_1412,N_1286,N_1221);
or U1413 (N_1413,N_1249,N_1239);
nand U1414 (N_1414,N_1336,N_1319);
or U1415 (N_1415,N_1216,N_1229);
nor U1416 (N_1416,N_1324,N_1314);
and U1417 (N_1417,N_1241,N_1266);
and U1418 (N_1418,N_1277,N_1217);
nand U1419 (N_1419,N_1300,N_1306);
nand U1420 (N_1420,N_1326,N_1316);
xnor U1421 (N_1421,N_1264,N_1218);
nor U1422 (N_1422,N_1281,N_1346);
nand U1423 (N_1423,N_1290,N_1291);
nor U1424 (N_1424,N_1246,N_1243);
or U1425 (N_1425,N_1201,N_1238);
nor U1426 (N_1426,N_1206,N_1215);
or U1427 (N_1427,N_1348,N_1313);
and U1428 (N_1428,N_1272,N_1324);
xnor U1429 (N_1429,N_1306,N_1258);
nor U1430 (N_1430,N_1325,N_1204);
xor U1431 (N_1431,N_1230,N_1250);
nand U1432 (N_1432,N_1224,N_1246);
nand U1433 (N_1433,N_1320,N_1204);
or U1434 (N_1434,N_1231,N_1219);
xnor U1435 (N_1435,N_1282,N_1315);
xnor U1436 (N_1436,N_1340,N_1204);
nand U1437 (N_1437,N_1269,N_1323);
nor U1438 (N_1438,N_1290,N_1263);
and U1439 (N_1439,N_1296,N_1321);
and U1440 (N_1440,N_1319,N_1291);
and U1441 (N_1441,N_1290,N_1304);
and U1442 (N_1442,N_1342,N_1208);
and U1443 (N_1443,N_1307,N_1305);
and U1444 (N_1444,N_1305,N_1293);
nand U1445 (N_1445,N_1263,N_1315);
and U1446 (N_1446,N_1330,N_1269);
and U1447 (N_1447,N_1249,N_1225);
or U1448 (N_1448,N_1233,N_1280);
and U1449 (N_1449,N_1337,N_1218);
xor U1450 (N_1450,N_1226,N_1308);
nor U1451 (N_1451,N_1263,N_1208);
xor U1452 (N_1452,N_1221,N_1328);
and U1453 (N_1453,N_1329,N_1254);
xor U1454 (N_1454,N_1304,N_1231);
or U1455 (N_1455,N_1235,N_1236);
nand U1456 (N_1456,N_1299,N_1247);
or U1457 (N_1457,N_1277,N_1251);
xor U1458 (N_1458,N_1262,N_1348);
xor U1459 (N_1459,N_1325,N_1282);
and U1460 (N_1460,N_1291,N_1343);
nand U1461 (N_1461,N_1301,N_1256);
or U1462 (N_1462,N_1295,N_1320);
and U1463 (N_1463,N_1217,N_1310);
and U1464 (N_1464,N_1201,N_1307);
or U1465 (N_1465,N_1218,N_1227);
xnor U1466 (N_1466,N_1256,N_1343);
xnor U1467 (N_1467,N_1346,N_1304);
or U1468 (N_1468,N_1260,N_1325);
nor U1469 (N_1469,N_1305,N_1209);
nor U1470 (N_1470,N_1212,N_1272);
or U1471 (N_1471,N_1337,N_1204);
nor U1472 (N_1472,N_1269,N_1284);
and U1473 (N_1473,N_1289,N_1253);
nor U1474 (N_1474,N_1294,N_1232);
xor U1475 (N_1475,N_1232,N_1345);
nor U1476 (N_1476,N_1205,N_1242);
nand U1477 (N_1477,N_1200,N_1339);
and U1478 (N_1478,N_1209,N_1310);
xnor U1479 (N_1479,N_1303,N_1236);
or U1480 (N_1480,N_1285,N_1232);
and U1481 (N_1481,N_1283,N_1269);
and U1482 (N_1482,N_1205,N_1265);
xnor U1483 (N_1483,N_1247,N_1274);
nor U1484 (N_1484,N_1274,N_1291);
xor U1485 (N_1485,N_1299,N_1295);
or U1486 (N_1486,N_1274,N_1345);
nand U1487 (N_1487,N_1333,N_1265);
and U1488 (N_1488,N_1274,N_1303);
nand U1489 (N_1489,N_1337,N_1275);
xnor U1490 (N_1490,N_1306,N_1270);
and U1491 (N_1491,N_1279,N_1344);
or U1492 (N_1492,N_1237,N_1229);
xor U1493 (N_1493,N_1336,N_1238);
xnor U1494 (N_1494,N_1261,N_1219);
or U1495 (N_1495,N_1328,N_1243);
and U1496 (N_1496,N_1324,N_1266);
and U1497 (N_1497,N_1214,N_1303);
or U1498 (N_1498,N_1277,N_1339);
or U1499 (N_1499,N_1325,N_1222);
xor U1500 (N_1500,N_1365,N_1367);
and U1501 (N_1501,N_1428,N_1379);
nand U1502 (N_1502,N_1497,N_1462);
nor U1503 (N_1503,N_1363,N_1362);
xnor U1504 (N_1504,N_1454,N_1413);
nor U1505 (N_1505,N_1381,N_1404);
xnor U1506 (N_1506,N_1374,N_1449);
nor U1507 (N_1507,N_1376,N_1409);
nand U1508 (N_1508,N_1364,N_1419);
and U1509 (N_1509,N_1373,N_1470);
and U1510 (N_1510,N_1429,N_1453);
xnor U1511 (N_1511,N_1397,N_1478);
nand U1512 (N_1512,N_1475,N_1441);
nor U1513 (N_1513,N_1358,N_1405);
nor U1514 (N_1514,N_1448,N_1480);
or U1515 (N_1515,N_1436,N_1439);
nor U1516 (N_1516,N_1458,N_1468);
nor U1517 (N_1517,N_1489,N_1457);
or U1518 (N_1518,N_1420,N_1482);
or U1519 (N_1519,N_1402,N_1494);
nor U1520 (N_1520,N_1401,N_1463);
or U1521 (N_1521,N_1407,N_1387);
nand U1522 (N_1522,N_1432,N_1385);
nor U1523 (N_1523,N_1447,N_1398);
nor U1524 (N_1524,N_1424,N_1491);
nor U1525 (N_1525,N_1459,N_1384);
nand U1526 (N_1526,N_1493,N_1380);
nor U1527 (N_1527,N_1389,N_1430);
nand U1528 (N_1528,N_1438,N_1456);
nand U1529 (N_1529,N_1464,N_1446);
or U1530 (N_1530,N_1486,N_1390);
xor U1531 (N_1531,N_1375,N_1484);
xnor U1532 (N_1532,N_1495,N_1366);
and U1533 (N_1533,N_1396,N_1411);
nand U1534 (N_1534,N_1477,N_1426);
or U1535 (N_1535,N_1455,N_1377);
and U1536 (N_1536,N_1435,N_1452);
or U1537 (N_1537,N_1487,N_1415);
nand U1538 (N_1538,N_1444,N_1394);
nor U1539 (N_1539,N_1417,N_1490);
and U1540 (N_1540,N_1492,N_1421);
or U1541 (N_1541,N_1434,N_1423);
nor U1542 (N_1542,N_1408,N_1354);
and U1543 (N_1543,N_1460,N_1361);
xor U1544 (N_1544,N_1469,N_1416);
nor U1545 (N_1545,N_1488,N_1400);
nor U1546 (N_1546,N_1393,N_1399);
or U1547 (N_1547,N_1382,N_1481);
nand U1548 (N_1548,N_1445,N_1414);
xor U1549 (N_1549,N_1425,N_1410);
or U1550 (N_1550,N_1479,N_1360);
and U1551 (N_1551,N_1383,N_1483);
nor U1552 (N_1552,N_1352,N_1471);
or U1553 (N_1553,N_1472,N_1355);
or U1554 (N_1554,N_1451,N_1412);
nor U1555 (N_1555,N_1386,N_1388);
nor U1556 (N_1556,N_1371,N_1496);
nor U1557 (N_1557,N_1450,N_1418);
xnor U1558 (N_1558,N_1442,N_1395);
or U1559 (N_1559,N_1350,N_1370);
nor U1560 (N_1560,N_1443,N_1467);
or U1561 (N_1561,N_1465,N_1403);
and U1562 (N_1562,N_1499,N_1372);
nand U1563 (N_1563,N_1498,N_1431);
xor U1564 (N_1564,N_1357,N_1392);
nand U1565 (N_1565,N_1406,N_1461);
xnor U1566 (N_1566,N_1485,N_1422);
and U1567 (N_1567,N_1476,N_1359);
xor U1568 (N_1568,N_1466,N_1391);
or U1569 (N_1569,N_1440,N_1473);
or U1570 (N_1570,N_1368,N_1433);
nand U1571 (N_1571,N_1369,N_1474);
nor U1572 (N_1572,N_1437,N_1427);
nor U1573 (N_1573,N_1351,N_1378);
or U1574 (N_1574,N_1356,N_1353);
nand U1575 (N_1575,N_1432,N_1374);
or U1576 (N_1576,N_1452,N_1362);
xnor U1577 (N_1577,N_1491,N_1455);
nand U1578 (N_1578,N_1390,N_1469);
or U1579 (N_1579,N_1424,N_1466);
nor U1580 (N_1580,N_1400,N_1388);
xnor U1581 (N_1581,N_1422,N_1421);
xnor U1582 (N_1582,N_1398,N_1438);
xor U1583 (N_1583,N_1482,N_1484);
nor U1584 (N_1584,N_1460,N_1364);
nand U1585 (N_1585,N_1454,N_1358);
xor U1586 (N_1586,N_1415,N_1470);
nand U1587 (N_1587,N_1474,N_1464);
or U1588 (N_1588,N_1369,N_1456);
xor U1589 (N_1589,N_1364,N_1397);
nand U1590 (N_1590,N_1434,N_1439);
or U1591 (N_1591,N_1392,N_1474);
nor U1592 (N_1592,N_1387,N_1356);
and U1593 (N_1593,N_1441,N_1482);
nor U1594 (N_1594,N_1372,N_1493);
or U1595 (N_1595,N_1485,N_1397);
nor U1596 (N_1596,N_1379,N_1477);
and U1597 (N_1597,N_1418,N_1465);
and U1598 (N_1598,N_1461,N_1470);
nor U1599 (N_1599,N_1390,N_1386);
and U1600 (N_1600,N_1352,N_1411);
and U1601 (N_1601,N_1446,N_1421);
or U1602 (N_1602,N_1355,N_1405);
or U1603 (N_1603,N_1425,N_1433);
or U1604 (N_1604,N_1492,N_1495);
nor U1605 (N_1605,N_1416,N_1420);
nor U1606 (N_1606,N_1366,N_1358);
or U1607 (N_1607,N_1399,N_1479);
and U1608 (N_1608,N_1473,N_1382);
xnor U1609 (N_1609,N_1416,N_1428);
xnor U1610 (N_1610,N_1490,N_1464);
nor U1611 (N_1611,N_1472,N_1372);
or U1612 (N_1612,N_1404,N_1382);
nand U1613 (N_1613,N_1431,N_1413);
or U1614 (N_1614,N_1366,N_1469);
nand U1615 (N_1615,N_1452,N_1472);
nor U1616 (N_1616,N_1466,N_1382);
xnor U1617 (N_1617,N_1463,N_1488);
and U1618 (N_1618,N_1387,N_1461);
and U1619 (N_1619,N_1422,N_1437);
nor U1620 (N_1620,N_1437,N_1429);
and U1621 (N_1621,N_1407,N_1465);
or U1622 (N_1622,N_1360,N_1399);
xor U1623 (N_1623,N_1385,N_1417);
nor U1624 (N_1624,N_1376,N_1419);
or U1625 (N_1625,N_1389,N_1462);
and U1626 (N_1626,N_1420,N_1410);
xor U1627 (N_1627,N_1381,N_1496);
or U1628 (N_1628,N_1482,N_1365);
nor U1629 (N_1629,N_1442,N_1389);
or U1630 (N_1630,N_1378,N_1377);
xor U1631 (N_1631,N_1434,N_1464);
xnor U1632 (N_1632,N_1448,N_1496);
or U1633 (N_1633,N_1422,N_1469);
xnor U1634 (N_1634,N_1421,N_1491);
or U1635 (N_1635,N_1392,N_1351);
nor U1636 (N_1636,N_1418,N_1456);
or U1637 (N_1637,N_1370,N_1367);
or U1638 (N_1638,N_1403,N_1411);
and U1639 (N_1639,N_1474,N_1445);
nand U1640 (N_1640,N_1464,N_1463);
nand U1641 (N_1641,N_1471,N_1489);
xnor U1642 (N_1642,N_1459,N_1371);
xnor U1643 (N_1643,N_1484,N_1370);
or U1644 (N_1644,N_1424,N_1350);
or U1645 (N_1645,N_1457,N_1421);
nor U1646 (N_1646,N_1448,N_1413);
nor U1647 (N_1647,N_1451,N_1390);
nand U1648 (N_1648,N_1404,N_1473);
nand U1649 (N_1649,N_1359,N_1407);
and U1650 (N_1650,N_1569,N_1501);
nand U1651 (N_1651,N_1628,N_1632);
xor U1652 (N_1652,N_1504,N_1541);
nand U1653 (N_1653,N_1557,N_1614);
nand U1654 (N_1654,N_1538,N_1624);
nand U1655 (N_1655,N_1563,N_1556);
and U1656 (N_1656,N_1546,N_1559);
nand U1657 (N_1657,N_1516,N_1599);
nor U1658 (N_1658,N_1529,N_1593);
or U1659 (N_1659,N_1608,N_1631);
nand U1660 (N_1660,N_1519,N_1505);
nand U1661 (N_1661,N_1540,N_1583);
nor U1662 (N_1662,N_1513,N_1566);
nand U1663 (N_1663,N_1645,N_1509);
nor U1664 (N_1664,N_1567,N_1520);
xnor U1665 (N_1665,N_1502,N_1542);
nor U1666 (N_1666,N_1617,N_1573);
xnor U1667 (N_1667,N_1606,N_1572);
nand U1668 (N_1668,N_1536,N_1640);
nand U1669 (N_1669,N_1649,N_1588);
xnor U1670 (N_1670,N_1568,N_1543);
xor U1671 (N_1671,N_1630,N_1591);
or U1672 (N_1672,N_1545,N_1648);
nand U1673 (N_1673,N_1561,N_1511);
nand U1674 (N_1674,N_1636,N_1643);
and U1675 (N_1675,N_1549,N_1621);
nand U1676 (N_1676,N_1535,N_1598);
and U1677 (N_1677,N_1531,N_1577);
xor U1678 (N_1678,N_1618,N_1639);
or U1679 (N_1679,N_1604,N_1578);
nor U1680 (N_1680,N_1602,N_1500);
or U1681 (N_1681,N_1601,N_1551);
xor U1682 (N_1682,N_1587,N_1510);
or U1683 (N_1683,N_1633,N_1539);
nor U1684 (N_1684,N_1533,N_1503);
xnor U1685 (N_1685,N_1646,N_1575);
or U1686 (N_1686,N_1515,N_1638);
xnor U1687 (N_1687,N_1611,N_1605);
or U1688 (N_1688,N_1574,N_1571);
and U1689 (N_1689,N_1514,N_1527);
or U1690 (N_1690,N_1595,N_1619);
nand U1691 (N_1691,N_1647,N_1562);
and U1692 (N_1692,N_1550,N_1623);
nand U1693 (N_1693,N_1625,N_1560);
nand U1694 (N_1694,N_1635,N_1555);
xor U1695 (N_1695,N_1523,N_1544);
nor U1696 (N_1696,N_1553,N_1525);
and U1697 (N_1697,N_1558,N_1641);
and U1698 (N_1698,N_1596,N_1534);
xnor U1699 (N_1699,N_1530,N_1634);
or U1700 (N_1700,N_1594,N_1622);
nand U1701 (N_1701,N_1642,N_1532);
or U1702 (N_1702,N_1586,N_1627);
nor U1703 (N_1703,N_1564,N_1644);
and U1704 (N_1704,N_1508,N_1629);
nor U1705 (N_1705,N_1518,N_1537);
nand U1706 (N_1706,N_1612,N_1615);
nand U1707 (N_1707,N_1626,N_1580);
nand U1708 (N_1708,N_1526,N_1610);
and U1709 (N_1709,N_1584,N_1528);
or U1710 (N_1710,N_1579,N_1570);
and U1711 (N_1711,N_1590,N_1613);
and U1712 (N_1712,N_1522,N_1607);
nor U1713 (N_1713,N_1512,N_1616);
or U1714 (N_1714,N_1547,N_1597);
or U1715 (N_1715,N_1585,N_1620);
nor U1716 (N_1716,N_1554,N_1576);
and U1717 (N_1717,N_1524,N_1517);
xnor U1718 (N_1718,N_1589,N_1507);
xnor U1719 (N_1719,N_1609,N_1552);
or U1720 (N_1720,N_1548,N_1582);
nor U1721 (N_1721,N_1581,N_1521);
xnor U1722 (N_1722,N_1637,N_1603);
nor U1723 (N_1723,N_1506,N_1592);
or U1724 (N_1724,N_1600,N_1565);
or U1725 (N_1725,N_1564,N_1553);
and U1726 (N_1726,N_1640,N_1625);
xor U1727 (N_1727,N_1614,N_1591);
and U1728 (N_1728,N_1602,N_1615);
or U1729 (N_1729,N_1618,N_1620);
nand U1730 (N_1730,N_1552,N_1587);
nor U1731 (N_1731,N_1584,N_1616);
nor U1732 (N_1732,N_1539,N_1575);
or U1733 (N_1733,N_1514,N_1563);
nor U1734 (N_1734,N_1544,N_1535);
or U1735 (N_1735,N_1624,N_1604);
or U1736 (N_1736,N_1628,N_1635);
nand U1737 (N_1737,N_1501,N_1610);
or U1738 (N_1738,N_1610,N_1618);
nor U1739 (N_1739,N_1633,N_1601);
or U1740 (N_1740,N_1618,N_1605);
or U1741 (N_1741,N_1517,N_1647);
nand U1742 (N_1742,N_1602,N_1640);
nor U1743 (N_1743,N_1572,N_1636);
or U1744 (N_1744,N_1595,N_1577);
or U1745 (N_1745,N_1569,N_1581);
nand U1746 (N_1746,N_1562,N_1616);
nor U1747 (N_1747,N_1621,N_1587);
nor U1748 (N_1748,N_1564,N_1569);
xnor U1749 (N_1749,N_1524,N_1612);
xnor U1750 (N_1750,N_1649,N_1548);
nor U1751 (N_1751,N_1564,N_1522);
nor U1752 (N_1752,N_1531,N_1649);
nor U1753 (N_1753,N_1511,N_1646);
xor U1754 (N_1754,N_1520,N_1547);
and U1755 (N_1755,N_1544,N_1500);
or U1756 (N_1756,N_1601,N_1583);
and U1757 (N_1757,N_1629,N_1649);
or U1758 (N_1758,N_1583,N_1599);
nand U1759 (N_1759,N_1527,N_1590);
nor U1760 (N_1760,N_1588,N_1612);
and U1761 (N_1761,N_1592,N_1554);
nand U1762 (N_1762,N_1554,N_1637);
nor U1763 (N_1763,N_1508,N_1597);
nor U1764 (N_1764,N_1585,N_1617);
or U1765 (N_1765,N_1561,N_1547);
and U1766 (N_1766,N_1506,N_1639);
or U1767 (N_1767,N_1622,N_1544);
and U1768 (N_1768,N_1585,N_1610);
or U1769 (N_1769,N_1539,N_1527);
and U1770 (N_1770,N_1557,N_1641);
nand U1771 (N_1771,N_1644,N_1617);
nand U1772 (N_1772,N_1534,N_1521);
xnor U1773 (N_1773,N_1568,N_1584);
and U1774 (N_1774,N_1569,N_1597);
nand U1775 (N_1775,N_1606,N_1577);
or U1776 (N_1776,N_1621,N_1644);
xnor U1777 (N_1777,N_1531,N_1558);
or U1778 (N_1778,N_1551,N_1559);
or U1779 (N_1779,N_1558,N_1621);
nor U1780 (N_1780,N_1637,N_1619);
or U1781 (N_1781,N_1528,N_1506);
nor U1782 (N_1782,N_1629,N_1513);
xor U1783 (N_1783,N_1648,N_1584);
nor U1784 (N_1784,N_1527,N_1546);
nand U1785 (N_1785,N_1562,N_1635);
or U1786 (N_1786,N_1550,N_1532);
nor U1787 (N_1787,N_1542,N_1500);
xnor U1788 (N_1788,N_1523,N_1555);
and U1789 (N_1789,N_1521,N_1543);
xor U1790 (N_1790,N_1627,N_1576);
and U1791 (N_1791,N_1551,N_1550);
xnor U1792 (N_1792,N_1525,N_1597);
nor U1793 (N_1793,N_1643,N_1580);
nor U1794 (N_1794,N_1525,N_1639);
xor U1795 (N_1795,N_1610,N_1581);
and U1796 (N_1796,N_1567,N_1522);
xnor U1797 (N_1797,N_1501,N_1618);
nand U1798 (N_1798,N_1612,N_1551);
nor U1799 (N_1799,N_1526,N_1569);
or U1800 (N_1800,N_1741,N_1660);
nand U1801 (N_1801,N_1715,N_1699);
or U1802 (N_1802,N_1698,N_1781);
xor U1803 (N_1803,N_1795,N_1655);
and U1804 (N_1804,N_1790,N_1667);
nor U1805 (N_1805,N_1745,N_1783);
xnor U1806 (N_1806,N_1776,N_1784);
or U1807 (N_1807,N_1742,N_1739);
nor U1808 (N_1808,N_1716,N_1704);
nand U1809 (N_1809,N_1688,N_1793);
nor U1810 (N_1810,N_1749,N_1683);
nor U1811 (N_1811,N_1737,N_1738);
nor U1812 (N_1812,N_1798,N_1762);
nand U1813 (N_1813,N_1725,N_1756);
nand U1814 (N_1814,N_1734,N_1751);
nand U1815 (N_1815,N_1730,N_1799);
and U1816 (N_1816,N_1712,N_1706);
nand U1817 (N_1817,N_1674,N_1746);
and U1818 (N_1818,N_1720,N_1695);
xnor U1819 (N_1819,N_1797,N_1714);
nand U1820 (N_1820,N_1687,N_1778);
or U1821 (N_1821,N_1753,N_1789);
nand U1822 (N_1822,N_1752,N_1669);
or U1823 (N_1823,N_1766,N_1777);
and U1824 (N_1824,N_1728,N_1703);
nor U1825 (N_1825,N_1772,N_1775);
nand U1826 (N_1826,N_1765,N_1711);
or U1827 (N_1827,N_1710,N_1694);
nand U1828 (N_1828,N_1785,N_1740);
nor U1829 (N_1829,N_1693,N_1701);
nand U1830 (N_1830,N_1782,N_1702);
xnor U1831 (N_1831,N_1653,N_1767);
xnor U1832 (N_1832,N_1657,N_1686);
or U1833 (N_1833,N_1689,N_1676);
and U1834 (N_1834,N_1774,N_1773);
xnor U1835 (N_1835,N_1675,N_1757);
xor U1836 (N_1836,N_1659,N_1684);
xor U1837 (N_1837,N_1652,N_1786);
nand U1838 (N_1838,N_1729,N_1743);
nor U1839 (N_1839,N_1733,N_1780);
xor U1840 (N_1840,N_1692,N_1665);
and U1841 (N_1841,N_1691,N_1650);
and U1842 (N_1842,N_1673,N_1754);
nand U1843 (N_1843,N_1763,N_1705);
nor U1844 (N_1844,N_1685,N_1656);
nor U1845 (N_1845,N_1681,N_1791);
xnor U1846 (N_1846,N_1721,N_1758);
and U1847 (N_1847,N_1727,N_1663);
nor U1848 (N_1848,N_1748,N_1661);
and U1849 (N_1849,N_1690,N_1744);
nand U1850 (N_1850,N_1779,N_1726);
nand U1851 (N_1851,N_1787,N_1735);
nand U1852 (N_1852,N_1732,N_1700);
nand U1853 (N_1853,N_1682,N_1708);
nand U1854 (N_1854,N_1719,N_1654);
or U1855 (N_1855,N_1718,N_1671);
nand U1856 (N_1856,N_1672,N_1696);
nor U1857 (N_1857,N_1792,N_1731);
or U1858 (N_1858,N_1724,N_1760);
and U1859 (N_1859,N_1670,N_1717);
or U1860 (N_1860,N_1658,N_1736);
xor U1861 (N_1861,N_1668,N_1664);
nand U1862 (N_1862,N_1794,N_1769);
and U1863 (N_1863,N_1722,N_1713);
and U1864 (N_1864,N_1768,N_1759);
nand U1865 (N_1865,N_1761,N_1679);
xnor U1866 (N_1866,N_1755,N_1764);
nand U1867 (N_1867,N_1770,N_1709);
xnor U1868 (N_1868,N_1723,N_1707);
nand U1869 (N_1869,N_1677,N_1680);
or U1870 (N_1870,N_1747,N_1788);
nor U1871 (N_1871,N_1697,N_1651);
xnor U1872 (N_1872,N_1666,N_1771);
or U1873 (N_1873,N_1750,N_1796);
nand U1874 (N_1874,N_1678,N_1662);
or U1875 (N_1875,N_1750,N_1730);
nor U1876 (N_1876,N_1744,N_1735);
or U1877 (N_1877,N_1778,N_1786);
or U1878 (N_1878,N_1708,N_1678);
xor U1879 (N_1879,N_1780,N_1731);
nand U1880 (N_1880,N_1655,N_1765);
or U1881 (N_1881,N_1795,N_1711);
and U1882 (N_1882,N_1778,N_1728);
nor U1883 (N_1883,N_1771,N_1784);
xnor U1884 (N_1884,N_1713,N_1668);
xor U1885 (N_1885,N_1657,N_1796);
xnor U1886 (N_1886,N_1741,N_1705);
nor U1887 (N_1887,N_1799,N_1779);
nor U1888 (N_1888,N_1707,N_1736);
xor U1889 (N_1889,N_1750,N_1758);
or U1890 (N_1890,N_1753,N_1717);
xnor U1891 (N_1891,N_1708,N_1733);
and U1892 (N_1892,N_1741,N_1784);
and U1893 (N_1893,N_1686,N_1754);
and U1894 (N_1894,N_1693,N_1793);
and U1895 (N_1895,N_1667,N_1678);
and U1896 (N_1896,N_1710,N_1766);
and U1897 (N_1897,N_1733,N_1774);
nor U1898 (N_1898,N_1757,N_1687);
nor U1899 (N_1899,N_1780,N_1695);
or U1900 (N_1900,N_1747,N_1664);
nand U1901 (N_1901,N_1743,N_1741);
nor U1902 (N_1902,N_1731,N_1664);
nand U1903 (N_1903,N_1788,N_1695);
nor U1904 (N_1904,N_1796,N_1662);
or U1905 (N_1905,N_1687,N_1717);
or U1906 (N_1906,N_1679,N_1782);
nand U1907 (N_1907,N_1658,N_1777);
and U1908 (N_1908,N_1667,N_1740);
and U1909 (N_1909,N_1753,N_1750);
or U1910 (N_1910,N_1705,N_1745);
and U1911 (N_1911,N_1785,N_1683);
or U1912 (N_1912,N_1658,N_1672);
nor U1913 (N_1913,N_1736,N_1691);
nor U1914 (N_1914,N_1789,N_1709);
nand U1915 (N_1915,N_1758,N_1760);
xnor U1916 (N_1916,N_1720,N_1729);
and U1917 (N_1917,N_1722,N_1742);
and U1918 (N_1918,N_1748,N_1675);
or U1919 (N_1919,N_1685,N_1715);
nor U1920 (N_1920,N_1688,N_1681);
or U1921 (N_1921,N_1694,N_1754);
xnor U1922 (N_1922,N_1707,N_1728);
xor U1923 (N_1923,N_1662,N_1713);
nor U1924 (N_1924,N_1682,N_1688);
nor U1925 (N_1925,N_1661,N_1795);
xor U1926 (N_1926,N_1668,N_1767);
nand U1927 (N_1927,N_1730,N_1761);
nand U1928 (N_1928,N_1657,N_1763);
nor U1929 (N_1929,N_1775,N_1791);
or U1930 (N_1930,N_1703,N_1696);
xor U1931 (N_1931,N_1689,N_1713);
and U1932 (N_1932,N_1790,N_1654);
and U1933 (N_1933,N_1791,N_1703);
xnor U1934 (N_1934,N_1747,N_1716);
nor U1935 (N_1935,N_1695,N_1728);
nor U1936 (N_1936,N_1684,N_1744);
and U1937 (N_1937,N_1720,N_1745);
or U1938 (N_1938,N_1675,N_1658);
xnor U1939 (N_1939,N_1667,N_1747);
nor U1940 (N_1940,N_1729,N_1740);
nor U1941 (N_1941,N_1708,N_1657);
nand U1942 (N_1942,N_1714,N_1665);
or U1943 (N_1943,N_1659,N_1721);
xnor U1944 (N_1944,N_1737,N_1731);
xnor U1945 (N_1945,N_1763,N_1655);
xor U1946 (N_1946,N_1737,N_1665);
nand U1947 (N_1947,N_1725,N_1697);
and U1948 (N_1948,N_1662,N_1793);
nand U1949 (N_1949,N_1694,N_1675);
nor U1950 (N_1950,N_1892,N_1826);
nand U1951 (N_1951,N_1866,N_1915);
nor U1952 (N_1952,N_1804,N_1914);
and U1953 (N_1953,N_1818,N_1832);
nand U1954 (N_1954,N_1881,N_1810);
or U1955 (N_1955,N_1886,N_1827);
nor U1956 (N_1956,N_1943,N_1836);
xor U1957 (N_1957,N_1942,N_1903);
and U1958 (N_1958,N_1839,N_1837);
xor U1959 (N_1959,N_1910,N_1946);
xor U1960 (N_1960,N_1927,N_1940);
xnor U1961 (N_1961,N_1851,N_1803);
xnor U1962 (N_1962,N_1842,N_1843);
nand U1963 (N_1963,N_1852,N_1805);
xnor U1964 (N_1964,N_1868,N_1876);
or U1965 (N_1965,N_1816,N_1934);
or U1966 (N_1966,N_1922,N_1885);
nand U1967 (N_1967,N_1874,N_1801);
and U1968 (N_1968,N_1905,N_1854);
and U1969 (N_1969,N_1841,N_1879);
xnor U1970 (N_1970,N_1902,N_1898);
and U1971 (N_1971,N_1880,N_1821);
and U1972 (N_1972,N_1928,N_1916);
and U1973 (N_1973,N_1800,N_1864);
nor U1974 (N_1974,N_1812,N_1840);
nand U1975 (N_1975,N_1877,N_1925);
nor U1976 (N_1976,N_1937,N_1814);
nor U1977 (N_1977,N_1893,N_1856);
nand U1978 (N_1978,N_1887,N_1918);
xor U1979 (N_1979,N_1859,N_1863);
or U1980 (N_1980,N_1917,N_1857);
nand U1981 (N_1981,N_1947,N_1890);
nor U1982 (N_1982,N_1846,N_1936);
nor U1983 (N_1983,N_1822,N_1929);
or U1984 (N_1984,N_1948,N_1853);
nand U1985 (N_1985,N_1931,N_1889);
and U1986 (N_1986,N_1921,N_1867);
or U1987 (N_1987,N_1825,N_1847);
nor U1988 (N_1988,N_1923,N_1884);
nand U1989 (N_1989,N_1811,N_1913);
and U1990 (N_1990,N_1869,N_1838);
nor U1991 (N_1991,N_1834,N_1862);
or U1992 (N_1992,N_1829,N_1807);
nor U1993 (N_1993,N_1932,N_1938);
and U1994 (N_1994,N_1909,N_1870);
or U1995 (N_1995,N_1849,N_1872);
nor U1996 (N_1996,N_1802,N_1824);
xor U1997 (N_1997,N_1945,N_1919);
nand U1998 (N_1998,N_1930,N_1820);
nand U1999 (N_1999,N_1858,N_1809);
nor U2000 (N_2000,N_1896,N_1835);
nand U2001 (N_2001,N_1897,N_1941);
and U2002 (N_2002,N_1873,N_1926);
nor U2003 (N_2003,N_1860,N_1823);
or U2004 (N_2004,N_1895,N_1907);
nor U2005 (N_2005,N_1935,N_1828);
xor U2006 (N_2006,N_1815,N_1806);
and U2007 (N_2007,N_1882,N_1861);
xnor U2008 (N_2008,N_1908,N_1906);
nor U2009 (N_2009,N_1899,N_1949);
nand U2010 (N_2010,N_1871,N_1813);
and U2011 (N_2011,N_1891,N_1894);
xnor U2012 (N_2012,N_1878,N_1904);
and U2013 (N_2013,N_1808,N_1831);
nand U2014 (N_2014,N_1944,N_1901);
nor U2015 (N_2015,N_1933,N_1855);
nor U2016 (N_2016,N_1883,N_1875);
or U2017 (N_2017,N_1920,N_1911);
xnor U2018 (N_2018,N_1939,N_1924);
and U2019 (N_2019,N_1848,N_1833);
xnor U2020 (N_2020,N_1900,N_1817);
or U2021 (N_2021,N_1888,N_1845);
xor U2022 (N_2022,N_1865,N_1830);
or U2023 (N_2023,N_1912,N_1850);
nand U2024 (N_2024,N_1819,N_1844);
xor U2025 (N_2025,N_1909,N_1815);
nand U2026 (N_2026,N_1929,N_1940);
or U2027 (N_2027,N_1812,N_1847);
nor U2028 (N_2028,N_1941,N_1920);
or U2029 (N_2029,N_1905,N_1878);
nor U2030 (N_2030,N_1829,N_1851);
nor U2031 (N_2031,N_1932,N_1867);
nand U2032 (N_2032,N_1899,N_1892);
xnor U2033 (N_2033,N_1830,N_1947);
xor U2034 (N_2034,N_1873,N_1944);
nand U2035 (N_2035,N_1896,N_1891);
and U2036 (N_2036,N_1938,N_1887);
nand U2037 (N_2037,N_1844,N_1841);
and U2038 (N_2038,N_1878,N_1897);
nor U2039 (N_2039,N_1889,N_1898);
nand U2040 (N_2040,N_1853,N_1906);
and U2041 (N_2041,N_1842,N_1936);
or U2042 (N_2042,N_1939,N_1933);
nand U2043 (N_2043,N_1877,N_1893);
nor U2044 (N_2044,N_1850,N_1825);
xnor U2045 (N_2045,N_1890,N_1880);
or U2046 (N_2046,N_1818,N_1803);
and U2047 (N_2047,N_1841,N_1905);
or U2048 (N_2048,N_1931,N_1882);
xor U2049 (N_2049,N_1848,N_1846);
or U2050 (N_2050,N_1948,N_1927);
xor U2051 (N_2051,N_1948,N_1854);
nand U2052 (N_2052,N_1939,N_1893);
and U2053 (N_2053,N_1813,N_1876);
or U2054 (N_2054,N_1939,N_1810);
or U2055 (N_2055,N_1882,N_1908);
and U2056 (N_2056,N_1862,N_1809);
xor U2057 (N_2057,N_1824,N_1806);
and U2058 (N_2058,N_1940,N_1943);
or U2059 (N_2059,N_1887,N_1900);
xnor U2060 (N_2060,N_1817,N_1864);
nor U2061 (N_2061,N_1929,N_1872);
nand U2062 (N_2062,N_1948,N_1894);
or U2063 (N_2063,N_1936,N_1911);
nor U2064 (N_2064,N_1944,N_1908);
nand U2065 (N_2065,N_1869,N_1820);
xnor U2066 (N_2066,N_1937,N_1840);
and U2067 (N_2067,N_1889,N_1922);
nor U2068 (N_2068,N_1907,N_1845);
and U2069 (N_2069,N_1826,N_1862);
nor U2070 (N_2070,N_1922,N_1944);
nor U2071 (N_2071,N_1934,N_1942);
nor U2072 (N_2072,N_1854,N_1802);
nand U2073 (N_2073,N_1809,N_1926);
xor U2074 (N_2074,N_1839,N_1892);
or U2075 (N_2075,N_1841,N_1921);
nand U2076 (N_2076,N_1909,N_1947);
nor U2077 (N_2077,N_1894,N_1827);
nand U2078 (N_2078,N_1807,N_1827);
nand U2079 (N_2079,N_1907,N_1920);
and U2080 (N_2080,N_1880,N_1937);
nor U2081 (N_2081,N_1856,N_1801);
and U2082 (N_2082,N_1898,N_1925);
xnor U2083 (N_2083,N_1887,N_1837);
nand U2084 (N_2084,N_1809,N_1928);
nand U2085 (N_2085,N_1879,N_1865);
and U2086 (N_2086,N_1825,N_1826);
nor U2087 (N_2087,N_1812,N_1809);
or U2088 (N_2088,N_1865,N_1924);
and U2089 (N_2089,N_1949,N_1894);
or U2090 (N_2090,N_1905,N_1861);
nor U2091 (N_2091,N_1928,N_1903);
and U2092 (N_2092,N_1824,N_1864);
and U2093 (N_2093,N_1802,N_1855);
or U2094 (N_2094,N_1846,N_1929);
xnor U2095 (N_2095,N_1942,N_1840);
nand U2096 (N_2096,N_1878,N_1891);
or U2097 (N_2097,N_1885,N_1911);
or U2098 (N_2098,N_1911,N_1818);
and U2099 (N_2099,N_1923,N_1925);
nor U2100 (N_2100,N_2035,N_1953);
nand U2101 (N_2101,N_2005,N_1968);
nor U2102 (N_2102,N_1967,N_2017);
or U2103 (N_2103,N_2031,N_2004);
or U2104 (N_2104,N_1955,N_2090);
nand U2105 (N_2105,N_2054,N_1966);
nand U2106 (N_2106,N_2095,N_1950);
nor U2107 (N_2107,N_2050,N_2043);
and U2108 (N_2108,N_2069,N_2087);
or U2109 (N_2109,N_1982,N_1972);
and U2110 (N_2110,N_1986,N_1969);
and U2111 (N_2111,N_2047,N_2070);
or U2112 (N_2112,N_1962,N_1983);
or U2113 (N_2113,N_2091,N_2098);
xor U2114 (N_2114,N_2071,N_2057);
nand U2115 (N_2115,N_2086,N_2073);
nor U2116 (N_2116,N_2074,N_2018);
nand U2117 (N_2117,N_2033,N_2099);
and U2118 (N_2118,N_1988,N_1990);
nor U2119 (N_2119,N_1956,N_1996);
or U2120 (N_2120,N_2058,N_2042);
or U2121 (N_2121,N_2038,N_1963);
nor U2122 (N_2122,N_1998,N_2001);
nor U2123 (N_2123,N_2093,N_2076);
or U2124 (N_2124,N_2063,N_2048);
nor U2125 (N_2125,N_2077,N_2060);
xor U2126 (N_2126,N_1977,N_2036);
nand U2127 (N_2127,N_2006,N_2085);
and U2128 (N_2128,N_2023,N_2009);
or U2129 (N_2129,N_2064,N_2052);
nor U2130 (N_2130,N_1984,N_2041);
xor U2131 (N_2131,N_1952,N_2046);
or U2132 (N_2132,N_2025,N_1981);
or U2133 (N_2133,N_2066,N_1992);
nor U2134 (N_2134,N_2061,N_2062);
nor U2135 (N_2135,N_1975,N_1995);
xnor U2136 (N_2136,N_1993,N_1989);
nand U2137 (N_2137,N_2026,N_2089);
xor U2138 (N_2138,N_1987,N_2088);
nor U2139 (N_2139,N_1985,N_2092);
and U2140 (N_2140,N_2003,N_1994);
and U2141 (N_2141,N_2084,N_2024);
nand U2142 (N_2142,N_2078,N_2051);
nor U2143 (N_2143,N_1971,N_2040);
xnor U2144 (N_2144,N_1965,N_2014);
nand U2145 (N_2145,N_2083,N_2067);
nor U2146 (N_2146,N_2008,N_1979);
nor U2147 (N_2147,N_2012,N_2028);
nand U2148 (N_2148,N_2096,N_2097);
nand U2149 (N_2149,N_2029,N_1991);
nand U2150 (N_2150,N_1976,N_1954);
nand U2151 (N_2151,N_1961,N_2072);
and U2152 (N_2152,N_2037,N_2016);
or U2153 (N_2153,N_2059,N_2075);
or U2154 (N_2154,N_1973,N_2056);
nor U2155 (N_2155,N_1974,N_2015);
nor U2156 (N_2156,N_1958,N_2068);
xor U2157 (N_2157,N_2030,N_2053);
nand U2158 (N_2158,N_2065,N_1980);
nor U2159 (N_2159,N_2020,N_1999);
nand U2160 (N_2160,N_2027,N_2019);
or U2161 (N_2161,N_1959,N_2007);
or U2162 (N_2162,N_2002,N_2034);
nand U2163 (N_2163,N_1978,N_2011);
or U2164 (N_2164,N_2055,N_2010);
nand U2165 (N_2165,N_2021,N_2013);
nand U2166 (N_2166,N_2039,N_2049);
nand U2167 (N_2167,N_1951,N_2079);
nand U2168 (N_2168,N_2022,N_2094);
nand U2169 (N_2169,N_2081,N_1997);
nand U2170 (N_2170,N_2032,N_2000);
or U2171 (N_2171,N_2082,N_2045);
and U2172 (N_2172,N_2080,N_1957);
nor U2173 (N_2173,N_1964,N_2044);
xnor U2174 (N_2174,N_1970,N_1960);
or U2175 (N_2175,N_2014,N_1978);
and U2176 (N_2176,N_2080,N_2072);
or U2177 (N_2177,N_1977,N_1969);
nor U2178 (N_2178,N_1952,N_1950);
or U2179 (N_2179,N_1993,N_2097);
and U2180 (N_2180,N_2058,N_2048);
or U2181 (N_2181,N_1993,N_2054);
xnor U2182 (N_2182,N_2014,N_2025);
or U2183 (N_2183,N_1995,N_2090);
nor U2184 (N_2184,N_2066,N_2023);
or U2185 (N_2185,N_2007,N_2092);
xnor U2186 (N_2186,N_2015,N_2028);
and U2187 (N_2187,N_2036,N_1960);
and U2188 (N_2188,N_1999,N_2067);
nand U2189 (N_2189,N_2071,N_1991);
and U2190 (N_2190,N_1984,N_2045);
nand U2191 (N_2191,N_2023,N_1981);
nor U2192 (N_2192,N_2085,N_2026);
and U2193 (N_2193,N_1986,N_2005);
xor U2194 (N_2194,N_2058,N_2014);
nor U2195 (N_2195,N_2018,N_1954);
and U2196 (N_2196,N_1988,N_2073);
or U2197 (N_2197,N_2076,N_1990);
or U2198 (N_2198,N_2073,N_2015);
nand U2199 (N_2199,N_2041,N_1978);
or U2200 (N_2200,N_2022,N_2064);
xnor U2201 (N_2201,N_2041,N_2084);
xnor U2202 (N_2202,N_1975,N_2096);
nor U2203 (N_2203,N_1964,N_2006);
or U2204 (N_2204,N_1975,N_1996);
and U2205 (N_2205,N_2006,N_2083);
or U2206 (N_2206,N_1979,N_2088);
nor U2207 (N_2207,N_2006,N_2067);
nor U2208 (N_2208,N_1956,N_1959);
and U2209 (N_2209,N_2078,N_2074);
nand U2210 (N_2210,N_1968,N_1960);
and U2211 (N_2211,N_2059,N_2057);
and U2212 (N_2212,N_2032,N_1969);
nor U2213 (N_2213,N_2062,N_1999);
xor U2214 (N_2214,N_2005,N_2003);
and U2215 (N_2215,N_2065,N_2026);
xor U2216 (N_2216,N_2088,N_1996);
nor U2217 (N_2217,N_2085,N_1997);
nor U2218 (N_2218,N_2015,N_2006);
and U2219 (N_2219,N_2035,N_2094);
nor U2220 (N_2220,N_2036,N_2087);
xor U2221 (N_2221,N_2077,N_2092);
nand U2222 (N_2222,N_2058,N_2064);
nand U2223 (N_2223,N_1953,N_1975);
xnor U2224 (N_2224,N_2090,N_2072);
nor U2225 (N_2225,N_2035,N_2015);
or U2226 (N_2226,N_1966,N_2006);
or U2227 (N_2227,N_2051,N_2016);
nand U2228 (N_2228,N_1980,N_2035);
or U2229 (N_2229,N_1978,N_2087);
nor U2230 (N_2230,N_2083,N_2068);
or U2231 (N_2231,N_2034,N_2068);
or U2232 (N_2232,N_1983,N_2060);
or U2233 (N_2233,N_1963,N_2010);
or U2234 (N_2234,N_2083,N_1975);
and U2235 (N_2235,N_1959,N_1965);
and U2236 (N_2236,N_2098,N_2092);
nand U2237 (N_2237,N_1997,N_2078);
nand U2238 (N_2238,N_2069,N_2061);
or U2239 (N_2239,N_1997,N_2059);
nor U2240 (N_2240,N_2040,N_2087);
xnor U2241 (N_2241,N_2029,N_2022);
and U2242 (N_2242,N_2023,N_2088);
xnor U2243 (N_2243,N_2034,N_2007);
xnor U2244 (N_2244,N_2078,N_2011);
nor U2245 (N_2245,N_2098,N_1970);
or U2246 (N_2246,N_2036,N_2079);
xnor U2247 (N_2247,N_1998,N_1954);
nor U2248 (N_2248,N_2034,N_2037);
and U2249 (N_2249,N_2069,N_2098);
and U2250 (N_2250,N_2240,N_2202);
nand U2251 (N_2251,N_2116,N_2181);
nand U2252 (N_2252,N_2186,N_2162);
xnor U2253 (N_2253,N_2132,N_2208);
or U2254 (N_2254,N_2158,N_2184);
or U2255 (N_2255,N_2229,N_2189);
xnor U2256 (N_2256,N_2179,N_2129);
xnor U2257 (N_2257,N_2243,N_2159);
xor U2258 (N_2258,N_2225,N_2236);
and U2259 (N_2259,N_2241,N_2111);
xor U2260 (N_2260,N_2102,N_2238);
or U2261 (N_2261,N_2115,N_2231);
nor U2262 (N_2262,N_2217,N_2148);
nand U2263 (N_2263,N_2237,N_2170);
and U2264 (N_2264,N_2196,N_2141);
nand U2265 (N_2265,N_2137,N_2163);
xnor U2266 (N_2266,N_2191,N_2212);
or U2267 (N_2267,N_2232,N_2108);
and U2268 (N_2268,N_2226,N_2112);
nor U2269 (N_2269,N_2194,N_2228);
nand U2270 (N_2270,N_2140,N_2185);
or U2271 (N_2271,N_2104,N_2220);
xor U2272 (N_2272,N_2248,N_2244);
and U2273 (N_2273,N_2143,N_2166);
and U2274 (N_2274,N_2134,N_2207);
and U2275 (N_2275,N_2172,N_2147);
or U2276 (N_2276,N_2110,N_2205);
and U2277 (N_2277,N_2201,N_2164);
nand U2278 (N_2278,N_2203,N_2101);
nor U2279 (N_2279,N_2157,N_2178);
nand U2280 (N_2280,N_2105,N_2188);
nor U2281 (N_2281,N_2119,N_2210);
and U2282 (N_2282,N_2180,N_2171);
xnor U2283 (N_2283,N_2204,N_2154);
nor U2284 (N_2284,N_2249,N_2136);
nand U2285 (N_2285,N_2224,N_2214);
or U2286 (N_2286,N_2197,N_2133);
and U2287 (N_2287,N_2218,N_2161);
or U2288 (N_2288,N_2230,N_2174);
xnor U2289 (N_2289,N_2160,N_2177);
xor U2290 (N_2290,N_2187,N_2247);
nand U2291 (N_2291,N_2200,N_2146);
xor U2292 (N_2292,N_2139,N_2100);
or U2293 (N_2293,N_2193,N_2168);
or U2294 (N_2294,N_2213,N_2128);
nand U2295 (N_2295,N_2221,N_2150);
xor U2296 (N_2296,N_2138,N_2227);
nor U2297 (N_2297,N_2109,N_2211);
nand U2298 (N_2298,N_2144,N_2245);
or U2299 (N_2299,N_2167,N_2176);
nor U2300 (N_2300,N_2169,N_2131);
nand U2301 (N_2301,N_2235,N_2121);
xnor U2302 (N_2302,N_2183,N_2223);
xor U2303 (N_2303,N_2222,N_2242);
and U2304 (N_2304,N_2182,N_2216);
xnor U2305 (N_2305,N_2234,N_2165);
nor U2306 (N_2306,N_2153,N_2151);
nand U2307 (N_2307,N_2190,N_2175);
xnor U2308 (N_2308,N_2206,N_2233);
xor U2309 (N_2309,N_2173,N_2122);
or U2310 (N_2310,N_2113,N_2114);
nor U2311 (N_2311,N_2103,N_2149);
nor U2312 (N_2312,N_2126,N_2239);
nand U2313 (N_2313,N_2199,N_2156);
and U2314 (N_2314,N_2123,N_2219);
nor U2315 (N_2315,N_2127,N_2120);
and U2316 (N_2316,N_2106,N_2155);
or U2317 (N_2317,N_2192,N_2118);
nand U2318 (N_2318,N_2246,N_2195);
xor U2319 (N_2319,N_2124,N_2135);
nor U2320 (N_2320,N_2209,N_2215);
xor U2321 (N_2321,N_2198,N_2142);
nand U2322 (N_2322,N_2107,N_2152);
or U2323 (N_2323,N_2130,N_2145);
or U2324 (N_2324,N_2117,N_2125);
and U2325 (N_2325,N_2157,N_2102);
nand U2326 (N_2326,N_2242,N_2186);
or U2327 (N_2327,N_2242,N_2138);
and U2328 (N_2328,N_2225,N_2196);
nor U2329 (N_2329,N_2169,N_2212);
xnor U2330 (N_2330,N_2222,N_2100);
xnor U2331 (N_2331,N_2102,N_2231);
nor U2332 (N_2332,N_2243,N_2242);
xnor U2333 (N_2333,N_2241,N_2233);
xor U2334 (N_2334,N_2189,N_2161);
or U2335 (N_2335,N_2183,N_2201);
nor U2336 (N_2336,N_2241,N_2171);
nand U2337 (N_2337,N_2211,N_2182);
and U2338 (N_2338,N_2200,N_2124);
or U2339 (N_2339,N_2116,N_2188);
or U2340 (N_2340,N_2143,N_2169);
xnor U2341 (N_2341,N_2116,N_2242);
nand U2342 (N_2342,N_2136,N_2231);
nor U2343 (N_2343,N_2134,N_2246);
nand U2344 (N_2344,N_2112,N_2159);
nor U2345 (N_2345,N_2194,N_2179);
nor U2346 (N_2346,N_2193,N_2116);
nand U2347 (N_2347,N_2103,N_2154);
and U2348 (N_2348,N_2145,N_2207);
nor U2349 (N_2349,N_2249,N_2163);
and U2350 (N_2350,N_2193,N_2122);
nor U2351 (N_2351,N_2232,N_2165);
or U2352 (N_2352,N_2206,N_2139);
xnor U2353 (N_2353,N_2210,N_2129);
and U2354 (N_2354,N_2169,N_2200);
nand U2355 (N_2355,N_2148,N_2231);
nor U2356 (N_2356,N_2110,N_2114);
xor U2357 (N_2357,N_2129,N_2146);
or U2358 (N_2358,N_2236,N_2114);
nand U2359 (N_2359,N_2234,N_2143);
nand U2360 (N_2360,N_2123,N_2238);
nand U2361 (N_2361,N_2238,N_2237);
and U2362 (N_2362,N_2178,N_2176);
nand U2363 (N_2363,N_2122,N_2181);
and U2364 (N_2364,N_2115,N_2166);
nor U2365 (N_2365,N_2115,N_2204);
nand U2366 (N_2366,N_2126,N_2246);
and U2367 (N_2367,N_2112,N_2105);
and U2368 (N_2368,N_2175,N_2224);
and U2369 (N_2369,N_2188,N_2219);
and U2370 (N_2370,N_2242,N_2119);
nor U2371 (N_2371,N_2167,N_2232);
or U2372 (N_2372,N_2119,N_2137);
xnor U2373 (N_2373,N_2109,N_2206);
or U2374 (N_2374,N_2176,N_2169);
nor U2375 (N_2375,N_2116,N_2103);
and U2376 (N_2376,N_2108,N_2130);
or U2377 (N_2377,N_2175,N_2179);
or U2378 (N_2378,N_2224,N_2215);
and U2379 (N_2379,N_2115,N_2144);
xor U2380 (N_2380,N_2189,N_2249);
nand U2381 (N_2381,N_2124,N_2127);
nor U2382 (N_2382,N_2146,N_2191);
and U2383 (N_2383,N_2237,N_2103);
or U2384 (N_2384,N_2243,N_2149);
nand U2385 (N_2385,N_2184,N_2135);
or U2386 (N_2386,N_2152,N_2168);
nand U2387 (N_2387,N_2166,N_2189);
or U2388 (N_2388,N_2245,N_2137);
xor U2389 (N_2389,N_2145,N_2124);
xor U2390 (N_2390,N_2241,N_2136);
xor U2391 (N_2391,N_2232,N_2155);
and U2392 (N_2392,N_2171,N_2161);
nand U2393 (N_2393,N_2213,N_2142);
or U2394 (N_2394,N_2152,N_2202);
nand U2395 (N_2395,N_2141,N_2109);
and U2396 (N_2396,N_2181,N_2102);
xor U2397 (N_2397,N_2153,N_2183);
xnor U2398 (N_2398,N_2219,N_2205);
or U2399 (N_2399,N_2103,N_2179);
nor U2400 (N_2400,N_2275,N_2259);
nor U2401 (N_2401,N_2313,N_2305);
xnor U2402 (N_2402,N_2357,N_2395);
nand U2403 (N_2403,N_2276,N_2355);
and U2404 (N_2404,N_2381,N_2293);
xnor U2405 (N_2405,N_2348,N_2336);
nor U2406 (N_2406,N_2374,N_2251);
and U2407 (N_2407,N_2302,N_2287);
and U2408 (N_2408,N_2391,N_2271);
or U2409 (N_2409,N_2361,N_2325);
nand U2410 (N_2410,N_2254,N_2345);
or U2411 (N_2411,N_2353,N_2387);
or U2412 (N_2412,N_2252,N_2289);
xnor U2413 (N_2413,N_2378,N_2328);
xnor U2414 (N_2414,N_2301,N_2322);
xor U2415 (N_2415,N_2333,N_2268);
nand U2416 (N_2416,N_2292,N_2369);
nand U2417 (N_2417,N_2320,N_2250);
and U2418 (N_2418,N_2299,N_2380);
and U2419 (N_2419,N_2282,N_2396);
nor U2420 (N_2420,N_2356,N_2274);
and U2421 (N_2421,N_2388,N_2281);
nand U2422 (N_2422,N_2359,N_2319);
nor U2423 (N_2423,N_2330,N_2354);
and U2424 (N_2424,N_2277,N_2331);
nand U2425 (N_2425,N_2340,N_2266);
nand U2426 (N_2426,N_2335,N_2365);
nor U2427 (N_2427,N_2257,N_2308);
nor U2428 (N_2428,N_2338,N_2253);
nor U2429 (N_2429,N_2290,N_2306);
nand U2430 (N_2430,N_2360,N_2273);
nand U2431 (N_2431,N_2364,N_2342);
and U2432 (N_2432,N_2346,N_2379);
nand U2433 (N_2433,N_2368,N_2260);
nand U2434 (N_2434,N_2362,N_2397);
and U2435 (N_2435,N_2270,N_2264);
nor U2436 (N_2436,N_2310,N_2341);
nand U2437 (N_2437,N_2377,N_2385);
xnor U2438 (N_2438,N_2337,N_2329);
xnor U2439 (N_2439,N_2372,N_2332);
or U2440 (N_2440,N_2291,N_2286);
or U2441 (N_2441,N_2351,N_2280);
or U2442 (N_2442,N_2288,N_2358);
or U2443 (N_2443,N_2383,N_2326);
nor U2444 (N_2444,N_2370,N_2297);
xor U2445 (N_2445,N_2386,N_2284);
nand U2446 (N_2446,N_2296,N_2373);
xor U2447 (N_2447,N_2344,N_2309);
or U2448 (N_2448,N_2375,N_2256);
xor U2449 (N_2449,N_2399,N_2334);
xor U2450 (N_2450,N_2303,N_2262);
and U2451 (N_2451,N_2315,N_2279);
nand U2452 (N_2452,N_2352,N_2283);
nor U2453 (N_2453,N_2255,N_2295);
and U2454 (N_2454,N_2265,N_2269);
and U2455 (N_2455,N_2321,N_2371);
and U2456 (N_2456,N_2304,N_2285);
and U2457 (N_2457,N_2261,N_2272);
and U2458 (N_2458,N_2258,N_2339);
nor U2459 (N_2459,N_2347,N_2317);
nand U2460 (N_2460,N_2350,N_2323);
nand U2461 (N_2461,N_2316,N_2394);
nor U2462 (N_2462,N_2389,N_2367);
nand U2463 (N_2463,N_2311,N_2278);
nor U2464 (N_2464,N_2300,N_2363);
xor U2465 (N_2465,N_2298,N_2349);
nor U2466 (N_2466,N_2366,N_2263);
xor U2467 (N_2467,N_2398,N_2314);
nor U2468 (N_2468,N_2307,N_2390);
nor U2469 (N_2469,N_2393,N_2392);
and U2470 (N_2470,N_2384,N_2294);
xnor U2471 (N_2471,N_2312,N_2382);
xor U2472 (N_2472,N_2324,N_2327);
or U2473 (N_2473,N_2343,N_2267);
nand U2474 (N_2474,N_2376,N_2318);
nand U2475 (N_2475,N_2330,N_2369);
nand U2476 (N_2476,N_2376,N_2268);
nor U2477 (N_2477,N_2322,N_2381);
or U2478 (N_2478,N_2306,N_2252);
or U2479 (N_2479,N_2370,N_2267);
or U2480 (N_2480,N_2258,N_2394);
or U2481 (N_2481,N_2337,N_2280);
and U2482 (N_2482,N_2390,N_2299);
or U2483 (N_2483,N_2324,N_2336);
or U2484 (N_2484,N_2396,N_2275);
xor U2485 (N_2485,N_2301,N_2326);
and U2486 (N_2486,N_2375,N_2323);
nand U2487 (N_2487,N_2277,N_2314);
nor U2488 (N_2488,N_2341,N_2292);
nor U2489 (N_2489,N_2395,N_2298);
nor U2490 (N_2490,N_2367,N_2276);
nor U2491 (N_2491,N_2370,N_2292);
xor U2492 (N_2492,N_2269,N_2270);
and U2493 (N_2493,N_2382,N_2280);
xor U2494 (N_2494,N_2389,N_2388);
nor U2495 (N_2495,N_2342,N_2326);
and U2496 (N_2496,N_2319,N_2273);
nand U2497 (N_2497,N_2389,N_2382);
nand U2498 (N_2498,N_2380,N_2309);
and U2499 (N_2499,N_2373,N_2252);
nor U2500 (N_2500,N_2324,N_2297);
and U2501 (N_2501,N_2256,N_2355);
nand U2502 (N_2502,N_2285,N_2364);
nand U2503 (N_2503,N_2300,N_2253);
xnor U2504 (N_2504,N_2280,N_2309);
or U2505 (N_2505,N_2303,N_2254);
or U2506 (N_2506,N_2341,N_2278);
or U2507 (N_2507,N_2322,N_2303);
nor U2508 (N_2508,N_2381,N_2341);
nor U2509 (N_2509,N_2340,N_2270);
nand U2510 (N_2510,N_2274,N_2277);
xnor U2511 (N_2511,N_2386,N_2273);
nor U2512 (N_2512,N_2321,N_2317);
and U2513 (N_2513,N_2336,N_2388);
nor U2514 (N_2514,N_2344,N_2335);
and U2515 (N_2515,N_2286,N_2362);
and U2516 (N_2516,N_2288,N_2265);
or U2517 (N_2517,N_2387,N_2285);
xnor U2518 (N_2518,N_2360,N_2399);
or U2519 (N_2519,N_2365,N_2362);
xor U2520 (N_2520,N_2307,N_2379);
nand U2521 (N_2521,N_2277,N_2363);
xor U2522 (N_2522,N_2349,N_2369);
or U2523 (N_2523,N_2329,N_2265);
and U2524 (N_2524,N_2369,N_2353);
xor U2525 (N_2525,N_2257,N_2293);
and U2526 (N_2526,N_2259,N_2258);
nand U2527 (N_2527,N_2344,N_2269);
and U2528 (N_2528,N_2395,N_2334);
nor U2529 (N_2529,N_2318,N_2346);
xor U2530 (N_2530,N_2374,N_2303);
nand U2531 (N_2531,N_2298,N_2264);
and U2532 (N_2532,N_2331,N_2338);
or U2533 (N_2533,N_2296,N_2293);
nand U2534 (N_2534,N_2289,N_2358);
or U2535 (N_2535,N_2256,N_2357);
and U2536 (N_2536,N_2267,N_2374);
nor U2537 (N_2537,N_2343,N_2251);
and U2538 (N_2538,N_2273,N_2283);
and U2539 (N_2539,N_2363,N_2274);
xnor U2540 (N_2540,N_2330,N_2375);
or U2541 (N_2541,N_2336,N_2290);
xnor U2542 (N_2542,N_2367,N_2266);
nor U2543 (N_2543,N_2259,N_2365);
nor U2544 (N_2544,N_2258,N_2322);
and U2545 (N_2545,N_2326,N_2250);
nor U2546 (N_2546,N_2341,N_2284);
or U2547 (N_2547,N_2295,N_2286);
xor U2548 (N_2548,N_2271,N_2293);
and U2549 (N_2549,N_2391,N_2281);
nand U2550 (N_2550,N_2500,N_2412);
nand U2551 (N_2551,N_2514,N_2477);
or U2552 (N_2552,N_2526,N_2441);
or U2553 (N_2553,N_2525,N_2509);
and U2554 (N_2554,N_2415,N_2442);
nor U2555 (N_2555,N_2437,N_2427);
and U2556 (N_2556,N_2444,N_2537);
xor U2557 (N_2557,N_2403,N_2485);
nand U2558 (N_2558,N_2533,N_2404);
or U2559 (N_2559,N_2425,N_2445);
nand U2560 (N_2560,N_2481,N_2453);
nor U2561 (N_2561,N_2498,N_2476);
nand U2562 (N_2562,N_2527,N_2470);
and U2563 (N_2563,N_2455,N_2434);
or U2564 (N_2564,N_2497,N_2504);
and U2565 (N_2565,N_2432,N_2417);
xor U2566 (N_2566,N_2420,N_2436);
nand U2567 (N_2567,N_2462,N_2465);
nor U2568 (N_2568,N_2494,N_2402);
and U2569 (N_2569,N_2535,N_2435);
nand U2570 (N_2570,N_2493,N_2474);
nand U2571 (N_2571,N_2548,N_2539);
and U2572 (N_2572,N_2523,N_2456);
or U2573 (N_2573,N_2433,N_2407);
nand U2574 (N_2574,N_2520,N_2515);
or U2575 (N_2575,N_2511,N_2458);
xnor U2576 (N_2576,N_2447,N_2422);
xor U2577 (N_2577,N_2409,N_2506);
or U2578 (N_2578,N_2475,N_2540);
nor U2579 (N_2579,N_2424,N_2516);
xor U2580 (N_2580,N_2521,N_2469);
xor U2581 (N_2581,N_2438,N_2471);
nor U2582 (N_2582,N_2513,N_2489);
nand U2583 (N_2583,N_2418,N_2426);
nor U2584 (N_2584,N_2541,N_2491);
xor U2585 (N_2585,N_2414,N_2510);
or U2586 (N_2586,N_2487,N_2495);
nor U2587 (N_2587,N_2478,N_2542);
xor U2588 (N_2588,N_2423,N_2543);
nor U2589 (N_2589,N_2463,N_2483);
nor U2590 (N_2590,N_2428,N_2466);
xnor U2591 (N_2591,N_2518,N_2501);
and U2592 (N_2592,N_2486,N_2460);
xnor U2593 (N_2593,N_2545,N_2488);
and U2594 (N_2594,N_2400,N_2490);
xnor U2595 (N_2595,N_2429,N_2411);
xor U2596 (N_2596,N_2536,N_2405);
nor U2597 (N_2597,N_2534,N_2502);
xor U2598 (N_2598,N_2484,N_2496);
xor U2599 (N_2599,N_2410,N_2529);
nand U2600 (N_2600,N_2503,N_2452);
or U2601 (N_2601,N_2492,N_2448);
or U2602 (N_2602,N_2482,N_2439);
nand U2603 (N_2603,N_2468,N_2528);
nor U2604 (N_2604,N_2499,N_2532);
nand U2605 (N_2605,N_2467,N_2419);
nand U2606 (N_2606,N_2507,N_2408);
or U2607 (N_2607,N_2430,N_2538);
and U2608 (N_2608,N_2547,N_2479);
xnor U2609 (N_2609,N_2546,N_2472);
nand U2610 (N_2610,N_2443,N_2524);
nor U2611 (N_2611,N_2473,N_2451);
xor U2612 (N_2612,N_2450,N_2401);
nand U2613 (N_2613,N_2480,N_2464);
nor U2614 (N_2614,N_2449,N_2522);
nand U2615 (N_2615,N_2421,N_2519);
nor U2616 (N_2616,N_2457,N_2431);
nand U2617 (N_2617,N_2549,N_2406);
and U2618 (N_2618,N_2530,N_2544);
or U2619 (N_2619,N_2459,N_2440);
xor U2620 (N_2620,N_2454,N_2446);
and U2621 (N_2621,N_2416,N_2508);
and U2622 (N_2622,N_2531,N_2461);
nor U2623 (N_2623,N_2413,N_2517);
or U2624 (N_2624,N_2505,N_2512);
xor U2625 (N_2625,N_2522,N_2469);
or U2626 (N_2626,N_2403,N_2535);
or U2627 (N_2627,N_2499,N_2491);
xor U2628 (N_2628,N_2431,N_2488);
nor U2629 (N_2629,N_2464,N_2448);
xor U2630 (N_2630,N_2426,N_2449);
or U2631 (N_2631,N_2465,N_2501);
or U2632 (N_2632,N_2401,N_2507);
or U2633 (N_2633,N_2478,N_2436);
or U2634 (N_2634,N_2441,N_2404);
nand U2635 (N_2635,N_2404,N_2412);
xor U2636 (N_2636,N_2400,N_2493);
xnor U2637 (N_2637,N_2502,N_2435);
nand U2638 (N_2638,N_2451,N_2449);
and U2639 (N_2639,N_2415,N_2422);
nor U2640 (N_2640,N_2436,N_2415);
and U2641 (N_2641,N_2442,N_2446);
and U2642 (N_2642,N_2445,N_2456);
and U2643 (N_2643,N_2476,N_2459);
xnor U2644 (N_2644,N_2482,N_2496);
nand U2645 (N_2645,N_2429,N_2495);
and U2646 (N_2646,N_2414,N_2469);
nand U2647 (N_2647,N_2480,N_2402);
and U2648 (N_2648,N_2524,N_2428);
and U2649 (N_2649,N_2437,N_2447);
nand U2650 (N_2650,N_2406,N_2449);
and U2651 (N_2651,N_2408,N_2532);
or U2652 (N_2652,N_2489,N_2436);
and U2653 (N_2653,N_2499,N_2503);
or U2654 (N_2654,N_2508,N_2533);
and U2655 (N_2655,N_2441,N_2483);
and U2656 (N_2656,N_2409,N_2518);
xor U2657 (N_2657,N_2494,N_2423);
nand U2658 (N_2658,N_2472,N_2501);
or U2659 (N_2659,N_2541,N_2502);
xnor U2660 (N_2660,N_2532,N_2450);
nor U2661 (N_2661,N_2549,N_2473);
nor U2662 (N_2662,N_2446,N_2431);
and U2663 (N_2663,N_2473,N_2456);
and U2664 (N_2664,N_2426,N_2406);
and U2665 (N_2665,N_2465,N_2526);
or U2666 (N_2666,N_2528,N_2514);
and U2667 (N_2667,N_2426,N_2501);
or U2668 (N_2668,N_2426,N_2508);
xor U2669 (N_2669,N_2488,N_2526);
or U2670 (N_2670,N_2534,N_2463);
xor U2671 (N_2671,N_2540,N_2401);
and U2672 (N_2672,N_2412,N_2427);
nand U2673 (N_2673,N_2487,N_2478);
and U2674 (N_2674,N_2532,N_2545);
nand U2675 (N_2675,N_2548,N_2440);
nand U2676 (N_2676,N_2515,N_2457);
xor U2677 (N_2677,N_2544,N_2503);
xnor U2678 (N_2678,N_2533,N_2509);
and U2679 (N_2679,N_2501,N_2484);
nor U2680 (N_2680,N_2526,N_2402);
and U2681 (N_2681,N_2437,N_2525);
nand U2682 (N_2682,N_2541,N_2532);
nand U2683 (N_2683,N_2435,N_2530);
and U2684 (N_2684,N_2413,N_2414);
xnor U2685 (N_2685,N_2478,N_2528);
nor U2686 (N_2686,N_2480,N_2448);
nand U2687 (N_2687,N_2471,N_2417);
nor U2688 (N_2688,N_2492,N_2538);
nor U2689 (N_2689,N_2521,N_2459);
or U2690 (N_2690,N_2401,N_2490);
nand U2691 (N_2691,N_2450,N_2546);
and U2692 (N_2692,N_2531,N_2544);
nor U2693 (N_2693,N_2422,N_2445);
nor U2694 (N_2694,N_2464,N_2453);
and U2695 (N_2695,N_2400,N_2429);
or U2696 (N_2696,N_2546,N_2531);
xnor U2697 (N_2697,N_2434,N_2511);
nand U2698 (N_2698,N_2509,N_2438);
or U2699 (N_2699,N_2429,N_2437);
nor U2700 (N_2700,N_2656,N_2637);
nor U2701 (N_2701,N_2560,N_2636);
xnor U2702 (N_2702,N_2667,N_2671);
nand U2703 (N_2703,N_2570,N_2592);
xor U2704 (N_2704,N_2629,N_2673);
and U2705 (N_2705,N_2664,N_2666);
nor U2706 (N_2706,N_2643,N_2670);
nand U2707 (N_2707,N_2680,N_2558);
or U2708 (N_2708,N_2630,N_2686);
xor U2709 (N_2709,N_2665,N_2655);
nor U2710 (N_2710,N_2650,N_2617);
xnor U2711 (N_2711,N_2627,N_2619);
xnor U2712 (N_2712,N_2674,N_2632);
or U2713 (N_2713,N_2618,N_2648);
xnor U2714 (N_2714,N_2660,N_2572);
nand U2715 (N_2715,N_2596,N_2698);
xnor U2716 (N_2716,N_2564,N_2669);
or U2717 (N_2717,N_2687,N_2692);
xor U2718 (N_2718,N_2641,N_2672);
and U2719 (N_2719,N_2590,N_2591);
nor U2720 (N_2720,N_2647,N_2603);
nor U2721 (N_2721,N_2616,N_2678);
or U2722 (N_2722,N_2638,N_2695);
xnor U2723 (N_2723,N_2694,N_2658);
nor U2724 (N_2724,N_2557,N_2697);
nand U2725 (N_2725,N_2693,N_2550);
xor U2726 (N_2726,N_2690,N_2657);
and U2727 (N_2727,N_2566,N_2649);
or U2728 (N_2728,N_2654,N_2587);
nor U2729 (N_2729,N_2579,N_2679);
xor U2730 (N_2730,N_2615,N_2668);
and U2731 (N_2731,N_2645,N_2659);
nand U2732 (N_2732,N_2639,N_2661);
and U2733 (N_2733,N_2553,N_2633);
or U2734 (N_2734,N_2689,N_2577);
and U2735 (N_2735,N_2682,N_2663);
or U2736 (N_2736,N_2677,N_2588);
or U2737 (N_2737,N_2582,N_2613);
xnor U2738 (N_2738,N_2635,N_2621);
xnor U2739 (N_2739,N_2681,N_2699);
nand U2740 (N_2740,N_2688,N_2585);
and U2741 (N_2741,N_2562,N_2563);
nor U2742 (N_2742,N_2598,N_2554);
xor U2743 (N_2743,N_2675,N_2584);
and U2744 (N_2744,N_2662,N_2640);
or U2745 (N_2745,N_2606,N_2568);
xor U2746 (N_2746,N_2623,N_2676);
or U2747 (N_2747,N_2607,N_2593);
nand U2748 (N_2748,N_2628,N_2576);
or U2749 (N_2749,N_2594,N_2624);
and U2750 (N_2750,N_2691,N_2575);
xor U2751 (N_2751,N_2652,N_2601);
xor U2752 (N_2752,N_2644,N_2620);
nand U2753 (N_2753,N_2565,N_2578);
nor U2754 (N_2754,N_2631,N_2556);
nor U2755 (N_2755,N_2614,N_2622);
xnor U2756 (N_2756,N_2612,N_2574);
nor U2757 (N_2757,N_2605,N_2684);
xnor U2758 (N_2758,N_2696,N_2625);
or U2759 (N_2759,N_2653,N_2651);
xor U2760 (N_2760,N_2551,N_2561);
xnor U2761 (N_2761,N_2642,N_2599);
xor U2762 (N_2762,N_2626,N_2567);
nand U2763 (N_2763,N_2569,N_2604);
nor U2764 (N_2764,N_2602,N_2581);
and U2765 (N_2765,N_2597,N_2571);
nor U2766 (N_2766,N_2580,N_2600);
or U2767 (N_2767,N_2609,N_2595);
nand U2768 (N_2768,N_2586,N_2611);
or U2769 (N_2769,N_2634,N_2608);
nand U2770 (N_2770,N_2555,N_2610);
xor U2771 (N_2771,N_2559,N_2583);
or U2772 (N_2772,N_2683,N_2646);
nand U2773 (N_2773,N_2573,N_2552);
xnor U2774 (N_2774,N_2589,N_2685);
or U2775 (N_2775,N_2692,N_2660);
and U2776 (N_2776,N_2652,N_2621);
nor U2777 (N_2777,N_2565,N_2659);
or U2778 (N_2778,N_2601,N_2599);
and U2779 (N_2779,N_2657,N_2609);
or U2780 (N_2780,N_2572,N_2640);
xor U2781 (N_2781,N_2638,N_2605);
or U2782 (N_2782,N_2643,N_2645);
xor U2783 (N_2783,N_2644,N_2562);
xor U2784 (N_2784,N_2650,N_2669);
nor U2785 (N_2785,N_2588,N_2691);
or U2786 (N_2786,N_2635,N_2607);
nor U2787 (N_2787,N_2694,N_2620);
xor U2788 (N_2788,N_2635,N_2618);
or U2789 (N_2789,N_2633,N_2643);
or U2790 (N_2790,N_2682,N_2564);
xor U2791 (N_2791,N_2657,N_2558);
xnor U2792 (N_2792,N_2627,N_2584);
nor U2793 (N_2793,N_2607,N_2566);
xor U2794 (N_2794,N_2614,N_2570);
and U2795 (N_2795,N_2607,N_2600);
nand U2796 (N_2796,N_2654,N_2570);
nand U2797 (N_2797,N_2643,N_2577);
nand U2798 (N_2798,N_2652,N_2638);
and U2799 (N_2799,N_2646,N_2629);
and U2800 (N_2800,N_2596,N_2574);
xor U2801 (N_2801,N_2645,N_2697);
and U2802 (N_2802,N_2600,N_2561);
and U2803 (N_2803,N_2591,N_2644);
nor U2804 (N_2804,N_2592,N_2593);
nand U2805 (N_2805,N_2685,N_2650);
and U2806 (N_2806,N_2603,N_2602);
or U2807 (N_2807,N_2558,N_2620);
xor U2808 (N_2808,N_2613,N_2668);
nor U2809 (N_2809,N_2698,N_2674);
or U2810 (N_2810,N_2623,N_2633);
xnor U2811 (N_2811,N_2596,N_2672);
and U2812 (N_2812,N_2559,N_2649);
xnor U2813 (N_2813,N_2617,N_2592);
xnor U2814 (N_2814,N_2697,N_2637);
nand U2815 (N_2815,N_2555,N_2564);
or U2816 (N_2816,N_2587,N_2626);
nand U2817 (N_2817,N_2607,N_2554);
and U2818 (N_2818,N_2590,N_2588);
nor U2819 (N_2819,N_2646,N_2588);
xor U2820 (N_2820,N_2687,N_2680);
and U2821 (N_2821,N_2570,N_2575);
nand U2822 (N_2822,N_2626,N_2683);
xor U2823 (N_2823,N_2628,N_2683);
nor U2824 (N_2824,N_2586,N_2617);
xnor U2825 (N_2825,N_2597,N_2653);
nand U2826 (N_2826,N_2598,N_2650);
and U2827 (N_2827,N_2645,N_2585);
or U2828 (N_2828,N_2571,N_2611);
xnor U2829 (N_2829,N_2565,N_2605);
nand U2830 (N_2830,N_2606,N_2586);
nand U2831 (N_2831,N_2628,N_2595);
xnor U2832 (N_2832,N_2569,N_2611);
and U2833 (N_2833,N_2592,N_2576);
nor U2834 (N_2834,N_2562,N_2651);
nor U2835 (N_2835,N_2698,N_2586);
or U2836 (N_2836,N_2571,N_2696);
nor U2837 (N_2837,N_2674,N_2697);
nand U2838 (N_2838,N_2636,N_2661);
and U2839 (N_2839,N_2550,N_2553);
nor U2840 (N_2840,N_2553,N_2649);
nand U2841 (N_2841,N_2618,N_2604);
and U2842 (N_2842,N_2561,N_2669);
nand U2843 (N_2843,N_2652,N_2661);
or U2844 (N_2844,N_2631,N_2583);
and U2845 (N_2845,N_2690,N_2605);
and U2846 (N_2846,N_2568,N_2646);
and U2847 (N_2847,N_2585,N_2690);
and U2848 (N_2848,N_2669,N_2612);
or U2849 (N_2849,N_2569,N_2575);
nor U2850 (N_2850,N_2720,N_2784);
and U2851 (N_2851,N_2743,N_2739);
xnor U2852 (N_2852,N_2849,N_2832);
or U2853 (N_2853,N_2771,N_2819);
xor U2854 (N_2854,N_2728,N_2715);
nand U2855 (N_2855,N_2736,N_2763);
xor U2856 (N_2856,N_2778,N_2790);
and U2857 (N_2857,N_2751,N_2809);
nand U2858 (N_2858,N_2812,N_2823);
and U2859 (N_2859,N_2818,N_2805);
and U2860 (N_2860,N_2710,N_2702);
nand U2861 (N_2861,N_2811,N_2744);
nor U2862 (N_2862,N_2735,N_2802);
xnor U2863 (N_2863,N_2772,N_2803);
nor U2864 (N_2864,N_2714,N_2724);
nor U2865 (N_2865,N_2755,N_2733);
or U2866 (N_2866,N_2748,N_2793);
and U2867 (N_2867,N_2775,N_2796);
xnor U2868 (N_2868,N_2709,N_2711);
nor U2869 (N_2869,N_2749,N_2829);
xor U2870 (N_2870,N_2825,N_2788);
or U2871 (N_2871,N_2700,N_2773);
and U2872 (N_2872,N_2729,N_2722);
and U2873 (N_2873,N_2701,N_2770);
nand U2874 (N_2874,N_2726,N_2753);
or U2875 (N_2875,N_2703,N_2712);
xnor U2876 (N_2876,N_2727,N_2835);
xor U2877 (N_2877,N_2836,N_2830);
or U2878 (N_2878,N_2756,N_2828);
and U2879 (N_2879,N_2741,N_2801);
and U2880 (N_2880,N_2837,N_2774);
nor U2881 (N_2881,N_2766,N_2732);
and U2882 (N_2882,N_2740,N_2731);
nand U2883 (N_2883,N_2780,N_2704);
and U2884 (N_2884,N_2846,N_2708);
or U2885 (N_2885,N_2795,N_2844);
and U2886 (N_2886,N_2705,N_2838);
or U2887 (N_2887,N_2806,N_2848);
xor U2888 (N_2888,N_2794,N_2734);
nand U2889 (N_2889,N_2831,N_2779);
or U2890 (N_2890,N_2777,N_2843);
nor U2891 (N_2891,N_2808,N_2821);
and U2892 (N_2892,N_2826,N_2759);
and U2893 (N_2893,N_2761,N_2776);
and U2894 (N_2894,N_2827,N_2719);
nand U2895 (N_2895,N_2797,N_2765);
and U2896 (N_2896,N_2817,N_2814);
nor U2897 (N_2897,N_2800,N_2816);
xnor U2898 (N_2898,N_2820,N_2730);
and U2899 (N_2899,N_2750,N_2787);
nand U2900 (N_2900,N_2721,N_2768);
xnor U2901 (N_2901,N_2785,N_2717);
or U2902 (N_2902,N_2782,N_2810);
or U2903 (N_2903,N_2747,N_2760);
or U2904 (N_2904,N_2842,N_2769);
xnor U2905 (N_2905,N_2833,N_2745);
and U2906 (N_2906,N_2783,N_2742);
or U2907 (N_2907,N_2791,N_2758);
nor U2908 (N_2908,N_2840,N_2767);
xor U2909 (N_2909,N_2804,N_2716);
nor U2910 (N_2910,N_2764,N_2752);
nor U2911 (N_2911,N_2839,N_2786);
or U2912 (N_2912,N_2822,N_2737);
nand U2913 (N_2913,N_2792,N_2824);
or U2914 (N_2914,N_2789,N_2781);
or U2915 (N_2915,N_2799,N_2841);
xor U2916 (N_2916,N_2813,N_2762);
xor U2917 (N_2917,N_2713,N_2757);
and U2918 (N_2918,N_2723,N_2815);
and U2919 (N_2919,N_2834,N_2725);
or U2920 (N_2920,N_2718,N_2738);
or U2921 (N_2921,N_2746,N_2847);
nor U2922 (N_2922,N_2845,N_2754);
xor U2923 (N_2923,N_2807,N_2706);
xor U2924 (N_2924,N_2707,N_2798);
nand U2925 (N_2925,N_2802,N_2777);
nor U2926 (N_2926,N_2833,N_2751);
xnor U2927 (N_2927,N_2760,N_2825);
xnor U2928 (N_2928,N_2817,N_2754);
or U2929 (N_2929,N_2748,N_2833);
and U2930 (N_2930,N_2779,N_2794);
and U2931 (N_2931,N_2842,N_2803);
xnor U2932 (N_2932,N_2797,N_2774);
nor U2933 (N_2933,N_2739,N_2710);
nand U2934 (N_2934,N_2768,N_2789);
nand U2935 (N_2935,N_2815,N_2783);
and U2936 (N_2936,N_2752,N_2769);
and U2937 (N_2937,N_2835,N_2846);
xor U2938 (N_2938,N_2797,N_2776);
or U2939 (N_2939,N_2765,N_2712);
nand U2940 (N_2940,N_2769,N_2750);
or U2941 (N_2941,N_2769,N_2801);
and U2942 (N_2942,N_2805,N_2744);
nor U2943 (N_2943,N_2806,N_2845);
or U2944 (N_2944,N_2846,N_2748);
or U2945 (N_2945,N_2799,N_2758);
or U2946 (N_2946,N_2722,N_2801);
nand U2947 (N_2947,N_2745,N_2717);
or U2948 (N_2948,N_2784,N_2764);
or U2949 (N_2949,N_2828,N_2795);
and U2950 (N_2950,N_2701,N_2847);
nand U2951 (N_2951,N_2819,N_2802);
or U2952 (N_2952,N_2701,N_2802);
and U2953 (N_2953,N_2810,N_2771);
nor U2954 (N_2954,N_2823,N_2729);
xnor U2955 (N_2955,N_2702,N_2739);
nand U2956 (N_2956,N_2706,N_2751);
or U2957 (N_2957,N_2819,N_2783);
or U2958 (N_2958,N_2816,N_2725);
nand U2959 (N_2959,N_2846,N_2717);
or U2960 (N_2960,N_2834,N_2760);
nand U2961 (N_2961,N_2734,N_2769);
and U2962 (N_2962,N_2709,N_2734);
and U2963 (N_2963,N_2771,N_2805);
and U2964 (N_2964,N_2725,N_2711);
xnor U2965 (N_2965,N_2722,N_2718);
nor U2966 (N_2966,N_2779,N_2834);
nand U2967 (N_2967,N_2809,N_2750);
and U2968 (N_2968,N_2738,N_2835);
and U2969 (N_2969,N_2848,N_2758);
or U2970 (N_2970,N_2840,N_2810);
nand U2971 (N_2971,N_2800,N_2730);
and U2972 (N_2972,N_2842,N_2753);
xor U2973 (N_2973,N_2724,N_2813);
xnor U2974 (N_2974,N_2829,N_2723);
nor U2975 (N_2975,N_2714,N_2823);
nor U2976 (N_2976,N_2720,N_2729);
or U2977 (N_2977,N_2807,N_2758);
nor U2978 (N_2978,N_2804,N_2773);
nand U2979 (N_2979,N_2836,N_2837);
xor U2980 (N_2980,N_2753,N_2793);
and U2981 (N_2981,N_2833,N_2815);
nor U2982 (N_2982,N_2747,N_2846);
nor U2983 (N_2983,N_2769,N_2751);
xnor U2984 (N_2984,N_2710,N_2830);
nand U2985 (N_2985,N_2820,N_2816);
nor U2986 (N_2986,N_2800,N_2741);
and U2987 (N_2987,N_2773,N_2735);
xor U2988 (N_2988,N_2728,N_2834);
nand U2989 (N_2989,N_2807,N_2716);
nor U2990 (N_2990,N_2794,N_2760);
nor U2991 (N_2991,N_2812,N_2822);
nand U2992 (N_2992,N_2821,N_2826);
nor U2993 (N_2993,N_2835,N_2740);
nor U2994 (N_2994,N_2824,N_2821);
and U2995 (N_2995,N_2776,N_2770);
or U2996 (N_2996,N_2709,N_2824);
or U2997 (N_2997,N_2794,N_2840);
and U2998 (N_2998,N_2848,N_2818);
or U2999 (N_2999,N_2767,N_2808);
nand U3000 (N_3000,N_2853,N_2928);
nand U3001 (N_3001,N_2935,N_2925);
and U3002 (N_3002,N_2970,N_2983);
and U3003 (N_3003,N_2886,N_2878);
nor U3004 (N_3004,N_2936,N_2915);
and U3005 (N_3005,N_2999,N_2978);
nand U3006 (N_3006,N_2974,N_2982);
and U3007 (N_3007,N_2892,N_2857);
and U3008 (N_3008,N_2998,N_2876);
or U3009 (N_3009,N_2950,N_2901);
nor U3010 (N_3010,N_2949,N_2855);
nand U3011 (N_3011,N_2986,N_2956);
and U3012 (N_3012,N_2906,N_2866);
nand U3013 (N_3013,N_2984,N_2941);
xnor U3014 (N_3014,N_2882,N_2902);
nand U3015 (N_3015,N_2851,N_2969);
nand U3016 (N_3016,N_2993,N_2959);
nand U3017 (N_3017,N_2887,N_2944);
and U3018 (N_3018,N_2923,N_2960);
nor U3019 (N_3019,N_2904,N_2896);
xnor U3020 (N_3020,N_2962,N_2933);
nand U3021 (N_3021,N_2918,N_2958);
and U3022 (N_3022,N_2893,N_2979);
nor U3023 (N_3023,N_2852,N_2955);
xnor U3024 (N_3024,N_2879,N_2860);
nor U3025 (N_3025,N_2854,N_2920);
nand U3026 (N_3026,N_2895,N_2943);
xnor U3027 (N_3027,N_2903,N_2953);
nor U3028 (N_3028,N_2899,N_2964);
nor U3029 (N_3029,N_2913,N_2890);
nor U3030 (N_3030,N_2988,N_2973);
or U3031 (N_3031,N_2880,N_2939);
nand U3032 (N_3032,N_2872,N_2865);
or U3033 (N_3033,N_2965,N_2907);
nor U3034 (N_3034,N_2968,N_2931);
nand U3035 (N_3035,N_2884,N_2908);
or U3036 (N_3036,N_2861,N_2946);
or U3037 (N_3037,N_2930,N_2971);
or U3038 (N_3038,N_2859,N_2991);
and U3039 (N_3039,N_2985,N_2975);
xnor U3040 (N_3040,N_2911,N_2924);
xnor U3041 (N_3041,N_2862,N_2850);
xor U3042 (N_3042,N_2864,N_2910);
and U3043 (N_3043,N_2881,N_2891);
and U3044 (N_3044,N_2980,N_2967);
xnor U3045 (N_3045,N_2929,N_2877);
xnor U3046 (N_3046,N_2938,N_2858);
and U3047 (N_3047,N_2868,N_2869);
nand U3048 (N_3048,N_2957,N_2875);
xor U3049 (N_3049,N_2873,N_2863);
nor U3050 (N_3050,N_2927,N_2952);
or U3051 (N_3051,N_2909,N_2919);
nand U3052 (N_3052,N_2994,N_2989);
or U3053 (N_3053,N_2981,N_2937);
and U3054 (N_3054,N_2932,N_2966);
nor U3055 (N_3055,N_2914,N_2997);
xnor U3056 (N_3056,N_2954,N_2996);
xnor U3057 (N_3057,N_2916,N_2922);
and U3058 (N_3058,N_2972,N_2948);
nand U3059 (N_3059,N_2894,N_2926);
xnor U3060 (N_3060,N_2990,N_2905);
and U3061 (N_3061,N_2870,N_2898);
and U3062 (N_3062,N_2900,N_2897);
xor U3063 (N_3063,N_2987,N_2889);
or U3064 (N_3064,N_2856,N_2934);
and U3065 (N_3065,N_2874,N_2951);
nand U3066 (N_3066,N_2871,N_2888);
and U3067 (N_3067,N_2995,N_2942);
nor U3068 (N_3068,N_2885,N_2977);
and U3069 (N_3069,N_2921,N_2883);
xor U3070 (N_3070,N_2976,N_2940);
xor U3071 (N_3071,N_2947,N_2945);
and U3072 (N_3072,N_2961,N_2917);
nor U3073 (N_3073,N_2992,N_2963);
and U3074 (N_3074,N_2912,N_2867);
nor U3075 (N_3075,N_2991,N_2941);
nand U3076 (N_3076,N_2959,N_2904);
nor U3077 (N_3077,N_2868,N_2906);
nand U3078 (N_3078,N_2999,N_2961);
xor U3079 (N_3079,N_2864,N_2993);
or U3080 (N_3080,N_2877,N_2899);
and U3081 (N_3081,N_2863,N_2995);
xnor U3082 (N_3082,N_2977,N_2959);
xor U3083 (N_3083,N_2892,N_2906);
xor U3084 (N_3084,N_2876,N_2908);
nand U3085 (N_3085,N_2862,N_2857);
xnor U3086 (N_3086,N_2867,N_2980);
or U3087 (N_3087,N_2993,N_2989);
nor U3088 (N_3088,N_2883,N_2925);
nand U3089 (N_3089,N_2955,N_2892);
nor U3090 (N_3090,N_2951,N_2857);
or U3091 (N_3091,N_2944,N_2951);
and U3092 (N_3092,N_2856,N_2889);
xnor U3093 (N_3093,N_2907,N_2874);
or U3094 (N_3094,N_2868,N_2944);
nor U3095 (N_3095,N_2970,N_2888);
and U3096 (N_3096,N_2852,N_2970);
nor U3097 (N_3097,N_2962,N_2973);
xnor U3098 (N_3098,N_2981,N_2955);
and U3099 (N_3099,N_2864,N_2981);
xnor U3100 (N_3100,N_2887,N_2901);
and U3101 (N_3101,N_2960,N_2901);
nand U3102 (N_3102,N_2925,N_2988);
nor U3103 (N_3103,N_2909,N_2862);
and U3104 (N_3104,N_2994,N_2899);
and U3105 (N_3105,N_2997,N_2913);
nor U3106 (N_3106,N_2934,N_2872);
xnor U3107 (N_3107,N_2941,N_2957);
or U3108 (N_3108,N_2931,N_2984);
nor U3109 (N_3109,N_2925,N_2957);
xnor U3110 (N_3110,N_2939,N_2857);
nor U3111 (N_3111,N_2996,N_2964);
or U3112 (N_3112,N_2894,N_2936);
nand U3113 (N_3113,N_2976,N_2968);
and U3114 (N_3114,N_2892,N_2919);
nand U3115 (N_3115,N_2951,N_2966);
xor U3116 (N_3116,N_2892,N_2851);
or U3117 (N_3117,N_2908,N_2917);
nand U3118 (N_3118,N_2973,N_2995);
xor U3119 (N_3119,N_2998,N_2861);
and U3120 (N_3120,N_2984,N_2867);
nor U3121 (N_3121,N_2953,N_2963);
xor U3122 (N_3122,N_2977,N_2908);
and U3123 (N_3123,N_2881,N_2956);
nor U3124 (N_3124,N_2948,N_2918);
nor U3125 (N_3125,N_2859,N_2976);
xnor U3126 (N_3126,N_2966,N_2883);
nor U3127 (N_3127,N_2856,N_2919);
or U3128 (N_3128,N_2903,N_2934);
or U3129 (N_3129,N_2855,N_2918);
and U3130 (N_3130,N_2967,N_2911);
or U3131 (N_3131,N_2959,N_2888);
xor U3132 (N_3132,N_2859,N_2897);
or U3133 (N_3133,N_2868,N_2983);
or U3134 (N_3134,N_2904,N_2863);
nand U3135 (N_3135,N_2858,N_2996);
nor U3136 (N_3136,N_2912,N_2869);
nand U3137 (N_3137,N_2920,N_2957);
nand U3138 (N_3138,N_2948,N_2962);
or U3139 (N_3139,N_2872,N_2867);
xor U3140 (N_3140,N_2935,N_2867);
xnor U3141 (N_3141,N_2869,N_2941);
and U3142 (N_3142,N_2885,N_2974);
xnor U3143 (N_3143,N_2858,N_2991);
and U3144 (N_3144,N_2936,N_2873);
and U3145 (N_3145,N_2990,N_2867);
xor U3146 (N_3146,N_2911,N_2906);
xnor U3147 (N_3147,N_2965,N_2982);
nand U3148 (N_3148,N_2861,N_2995);
nand U3149 (N_3149,N_2898,N_2978);
or U3150 (N_3150,N_3093,N_3030);
and U3151 (N_3151,N_3149,N_3078);
or U3152 (N_3152,N_3115,N_3135);
nand U3153 (N_3153,N_3025,N_3107);
nand U3154 (N_3154,N_3142,N_3101);
nor U3155 (N_3155,N_3081,N_3146);
nand U3156 (N_3156,N_3064,N_3011);
nor U3157 (N_3157,N_3027,N_3007);
xor U3158 (N_3158,N_3041,N_3092);
xnor U3159 (N_3159,N_3066,N_3130);
nor U3160 (N_3160,N_3074,N_3087);
xor U3161 (N_3161,N_3047,N_3144);
or U3162 (N_3162,N_3037,N_3004);
and U3163 (N_3163,N_3109,N_3126);
nor U3164 (N_3164,N_3127,N_3063);
or U3165 (N_3165,N_3108,N_3094);
nand U3166 (N_3166,N_3039,N_3133);
nand U3167 (N_3167,N_3040,N_3091);
xnor U3168 (N_3168,N_3015,N_3019);
and U3169 (N_3169,N_3117,N_3140);
nor U3170 (N_3170,N_3067,N_3137);
xnor U3171 (N_3171,N_3114,N_3124);
nor U3172 (N_3172,N_3042,N_3009);
and U3173 (N_3173,N_3033,N_3089);
and U3174 (N_3174,N_3029,N_3008);
nand U3175 (N_3175,N_3060,N_3084);
xnor U3176 (N_3176,N_3077,N_3131);
xor U3177 (N_3177,N_3032,N_3028);
nand U3178 (N_3178,N_3003,N_3075);
or U3179 (N_3179,N_3106,N_3006);
nor U3180 (N_3180,N_3110,N_3082);
and U3181 (N_3181,N_3129,N_3013);
and U3182 (N_3182,N_3070,N_3098);
nor U3183 (N_3183,N_3050,N_3053);
xor U3184 (N_3184,N_3112,N_3148);
nand U3185 (N_3185,N_3034,N_3125);
and U3186 (N_3186,N_3022,N_3086);
nor U3187 (N_3187,N_3016,N_3044);
nand U3188 (N_3188,N_3031,N_3145);
nor U3189 (N_3189,N_3071,N_3069);
nand U3190 (N_3190,N_3141,N_3134);
xor U3191 (N_3191,N_3072,N_3096);
or U3192 (N_3192,N_3113,N_3116);
or U3193 (N_3193,N_3100,N_3083);
nor U3194 (N_3194,N_3061,N_3080);
or U3195 (N_3195,N_3095,N_3017);
and U3196 (N_3196,N_3020,N_3000);
xnor U3197 (N_3197,N_3085,N_3036);
nand U3198 (N_3198,N_3076,N_3046);
or U3199 (N_3199,N_3024,N_3005);
nand U3200 (N_3200,N_3139,N_3065);
xor U3201 (N_3201,N_3054,N_3048);
or U3202 (N_3202,N_3097,N_3055);
or U3203 (N_3203,N_3049,N_3021);
or U3204 (N_3204,N_3128,N_3023);
and U3205 (N_3205,N_3088,N_3122);
nor U3206 (N_3206,N_3103,N_3014);
nor U3207 (N_3207,N_3111,N_3010);
or U3208 (N_3208,N_3132,N_3038);
nor U3209 (N_3209,N_3012,N_3068);
and U3210 (N_3210,N_3073,N_3136);
xor U3211 (N_3211,N_3057,N_3002);
nor U3212 (N_3212,N_3090,N_3026);
nand U3213 (N_3213,N_3056,N_3105);
xnor U3214 (N_3214,N_3035,N_3059);
or U3215 (N_3215,N_3018,N_3104);
or U3216 (N_3216,N_3051,N_3001);
xnor U3217 (N_3217,N_3062,N_3043);
or U3218 (N_3218,N_3121,N_3102);
or U3219 (N_3219,N_3099,N_3138);
and U3220 (N_3220,N_3079,N_3123);
xor U3221 (N_3221,N_3045,N_3143);
nor U3222 (N_3222,N_3119,N_3118);
and U3223 (N_3223,N_3120,N_3147);
xnor U3224 (N_3224,N_3052,N_3058);
or U3225 (N_3225,N_3038,N_3015);
nand U3226 (N_3226,N_3110,N_3122);
or U3227 (N_3227,N_3028,N_3095);
nor U3228 (N_3228,N_3143,N_3090);
nor U3229 (N_3229,N_3023,N_3019);
nor U3230 (N_3230,N_3118,N_3057);
or U3231 (N_3231,N_3135,N_3119);
and U3232 (N_3232,N_3132,N_3011);
and U3233 (N_3233,N_3146,N_3052);
and U3234 (N_3234,N_3089,N_3141);
and U3235 (N_3235,N_3026,N_3147);
xor U3236 (N_3236,N_3129,N_3066);
and U3237 (N_3237,N_3133,N_3053);
nand U3238 (N_3238,N_3105,N_3021);
and U3239 (N_3239,N_3082,N_3143);
nor U3240 (N_3240,N_3141,N_3013);
nor U3241 (N_3241,N_3001,N_3085);
xnor U3242 (N_3242,N_3046,N_3102);
and U3243 (N_3243,N_3145,N_3093);
nor U3244 (N_3244,N_3021,N_3100);
or U3245 (N_3245,N_3071,N_3037);
nand U3246 (N_3246,N_3005,N_3030);
and U3247 (N_3247,N_3045,N_3121);
nor U3248 (N_3248,N_3005,N_3046);
nand U3249 (N_3249,N_3141,N_3015);
or U3250 (N_3250,N_3046,N_3011);
and U3251 (N_3251,N_3011,N_3122);
xnor U3252 (N_3252,N_3045,N_3147);
nand U3253 (N_3253,N_3087,N_3002);
nand U3254 (N_3254,N_3060,N_3049);
xor U3255 (N_3255,N_3021,N_3068);
or U3256 (N_3256,N_3005,N_3137);
xor U3257 (N_3257,N_3061,N_3054);
nand U3258 (N_3258,N_3050,N_3006);
nand U3259 (N_3259,N_3004,N_3066);
and U3260 (N_3260,N_3143,N_3111);
and U3261 (N_3261,N_3133,N_3074);
and U3262 (N_3262,N_3145,N_3050);
or U3263 (N_3263,N_3117,N_3019);
nor U3264 (N_3264,N_3057,N_3075);
or U3265 (N_3265,N_3117,N_3006);
nand U3266 (N_3266,N_3091,N_3037);
xor U3267 (N_3267,N_3064,N_3054);
nand U3268 (N_3268,N_3076,N_3032);
nor U3269 (N_3269,N_3138,N_3008);
and U3270 (N_3270,N_3034,N_3059);
or U3271 (N_3271,N_3052,N_3053);
and U3272 (N_3272,N_3064,N_3137);
and U3273 (N_3273,N_3106,N_3051);
and U3274 (N_3274,N_3049,N_3144);
xnor U3275 (N_3275,N_3111,N_3130);
and U3276 (N_3276,N_3093,N_3059);
nor U3277 (N_3277,N_3108,N_3054);
and U3278 (N_3278,N_3032,N_3106);
nor U3279 (N_3279,N_3042,N_3073);
xnor U3280 (N_3280,N_3001,N_3026);
and U3281 (N_3281,N_3033,N_3097);
or U3282 (N_3282,N_3031,N_3063);
or U3283 (N_3283,N_3009,N_3059);
or U3284 (N_3284,N_3030,N_3127);
or U3285 (N_3285,N_3101,N_3044);
nor U3286 (N_3286,N_3090,N_3116);
and U3287 (N_3287,N_3129,N_3133);
and U3288 (N_3288,N_3030,N_3056);
nand U3289 (N_3289,N_3136,N_3110);
and U3290 (N_3290,N_3024,N_3119);
and U3291 (N_3291,N_3038,N_3109);
and U3292 (N_3292,N_3028,N_3127);
and U3293 (N_3293,N_3131,N_3079);
nand U3294 (N_3294,N_3062,N_3013);
xor U3295 (N_3295,N_3127,N_3141);
and U3296 (N_3296,N_3076,N_3117);
or U3297 (N_3297,N_3010,N_3100);
or U3298 (N_3298,N_3018,N_3057);
or U3299 (N_3299,N_3042,N_3113);
or U3300 (N_3300,N_3279,N_3219);
and U3301 (N_3301,N_3170,N_3214);
nor U3302 (N_3302,N_3181,N_3159);
and U3303 (N_3303,N_3224,N_3260);
xor U3304 (N_3304,N_3245,N_3221);
and U3305 (N_3305,N_3242,N_3211);
xnor U3306 (N_3306,N_3276,N_3246);
nand U3307 (N_3307,N_3266,N_3286);
nor U3308 (N_3308,N_3180,N_3281);
or U3309 (N_3309,N_3204,N_3161);
or U3310 (N_3310,N_3241,N_3201);
and U3311 (N_3311,N_3202,N_3230);
or U3312 (N_3312,N_3178,N_3155);
nand U3313 (N_3313,N_3207,N_3174);
or U3314 (N_3314,N_3233,N_3243);
or U3315 (N_3315,N_3272,N_3226);
or U3316 (N_3316,N_3259,N_3195);
or U3317 (N_3317,N_3191,N_3256);
nand U3318 (N_3318,N_3165,N_3196);
nor U3319 (N_3319,N_3283,N_3203);
nand U3320 (N_3320,N_3213,N_3265);
and U3321 (N_3321,N_3289,N_3227);
nand U3322 (N_3322,N_3229,N_3263);
nand U3323 (N_3323,N_3199,N_3277);
and U3324 (N_3324,N_3220,N_3215);
nor U3325 (N_3325,N_3291,N_3194);
xnor U3326 (N_3326,N_3231,N_3162);
and U3327 (N_3327,N_3298,N_3236);
nand U3328 (N_3328,N_3257,N_3206);
xor U3329 (N_3329,N_3189,N_3280);
nand U3330 (N_3330,N_3182,N_3158);
xor U3331 (N_3331,N_3152,N_3274);
nor U3332 (N_3332,N_3160,N_3288);
nor U3333 (N_3333,N_3252,N_3200);
or U3334 (N_3334,N_3166,N_3173);
nand U3335 (N_3335,N_3212,N_3228);
nor U3336 (N_3336,N_3264,N_3175);
and U3337 (N_3337,N_3187,N_3208);
nor U3338 (N_3338,N_3234,N_3153);
nor U3339 (N_3339,N_3254,N_3251);
xor U3340 (N_3340,N_3225,N_3240);
or U3341 (N_3341,N_3297,N_3258);
xnor U3342 (N_3342,N_3275,N_3296);
xor U3343 (N_3343,N_3271,N_3185);
and U3344 (N_3344,N_3190,N_3235);
nor U3345 (N_3345,N_3232,N_3284);
nor U3346 (N_3346,N_3249,N_3223);
or U3347 (N_3347,N_3216,N_3154);
nor U3348 (N_3348,N_3278,N_3217);
and U3349 (N_3349,N_3262,N_3177);
xnor U3350 (N_3350,N_3292,N_3237);
xnor U3351 (N_3351,N_3184,N_3295);
nand U3352 (N_3352,N_3163,N_3157);
xnor U3353 (N_3353,N_3169,N_3167);
or U3354 (N_3354,N_3255,N_3268);
or U3355 (N_3355,N_3172,N_3250);
and U3356 (N_3356,N_3171,N_3151);
xnor U3357 (N_3357,N_3253,N_3197);
or U3358 (N_3358,N_3168,N_3294);
xnor U3359 (N_3359,N_3205,N_3244);
or U3360 (N_3360,N_3218,N_3164);
and U3361 (N_3361,N_3179,N_3248);
and U3362 (N_3362,N_3282,N_3285);
nor U3363 (N_3363,N_3193,N_3287);
and U3364 (N_3364,N_3222,N_3239);
nor U3365 (N_3365,N_3238,N_3156);
or U3366 (N_3366,N_3209,N_3188);
xor U3367 (N_3367,N_3270,N_3176);
or U3368 (N_3368,N_3150,N_3290);
and U3369 (N_3369,N_3269,N_3186);
xnor U3370 (N_3370,N_3267,N_3299);
nand U3371 (N_3371,N_3198,N_3210);
nand U3372 (N_3372,N_3293,N_3273);
xor U3373 (N_3373,N_3192,N_3183);
or U3374 (N_3374,N_3261,N_3247);
nand U3375 (N_3375,N_3281,N_3162);
or U3376 (N_3376,N_3239,N_3211);
nor U3377 (N_3377,N_3299,N_3245);
nand U3378 (N_3378,N_3253,N_3202);
or U3379 (N_3379,N_3230,N_3187);
nand U3380 (N_3380,N_3217,N_3232);
nand U3381 (N_3381,N_3201,N_3223);
and U3382 (N_3382,N_3189,N_3173);
xor U3383 (N_3383,N_3204,N_3173);
nor U3384 (N_3384,N_3212,N_3221);
xor U3385 (N_3385,N_3239,N_3233);
xor U3386 (N_3386,N_3296,N_3185);
or U3387 (N_3387,N_3192,N_3272);
nor U3388 (N_3388,N_3180,N_3164);
or U3389 (N_3389,N_3229,N_3259);
nand U3390 (N_3390,N_3241,N_3220);
nor U3391 (N_3391,N_3184,N_3225);
nor U3392 (N_3392,N_3292,N_3239);
or U3393 (N_3393,N_3240,N_3206);
and U3394 (N_3394,N_3216,N_3159);
nor U3395 (N_3395,N_3239,N_3209);
and U3396 (N_3396,N_3226,N_3258);
nand U3397 (N_3397,N_3164,N_3217);
and U3398 (N_3398,N_3272,N_3278);
and U3399 (N_3399,N_3284,N_3285);
or U3400 (N_3400,N_3158,N_3277);
nand U3401 (N_3401,N_3195,N_3248);
xor U3402 (N_3402,N_3270,N_3256);
nand U3403 (N_3403,N_3150,N_3234);
or U3404 (N_3404,N_3178,N_3156);
or U3405 (N_3405,N_3255,N_3233);
or U3406 (N_3406,N_3169,N_3235);
xor U3407 (N_3407,N_3184,N_3234);
and U3408 (N_3408,N_3186,N_3161);
or U3409 (N_3409,N_3213,N_3224);
nor U3410 (N_3410,N_3257,N_3168);
xnor U3411 (N_3411,N_3218,N_3228);
and U3412 (N_3412,N_3261,N_3231);
xor U3413 (N_3413,N_3166,N_3163);
or U3414 (N_3414,N_3204,N_3252);
or U3415 (N_3415,N_3219,N_3275);
or U3416 (N_3416,N_3256,N_3171);
and U3417 (N_3417,N_3186,N_3206);
nand U3418 (N_3418,N_3295,N_3272);
xor U3419 (N_3419,N_3166,N_3190);
or U3420 (N_3420,N_3214,N_3268);
or U3421 (N_3421,N_3226,N_3229);
or U3422 (N_3422,N_3191,N_3225);
or U3423 (N_3423,N_3235,N_3221);
and U3424 (N_3424,N_3256,N_3258);
xor U3425 (N_3425,N_3271,N_3210);
nand U3426 (N_3426,N_3167,N_3236);
nand U3427 (N_3427,N_3257,N_3266);
or U3428 (N_3428,N_3244,N_3162);
and U3429 (N_3429,N_3229,N_3195);
and U3430 (N_3430,N_3166,N_3183);
and U3431 (N_3431,N_3152,N_3182);
or U3432 (N_3432,N_3254,N_3256);
xnor U3433 (N_3433,N_3224,N_3254);
nor U3434 (N_3434,N_3243,N_3160);
nand U3435 (N_3435,N_3203,N_3271);
and U3436 (N_3436,N_3277,N_3183);
nand U3437 (N_3437,N_3282,N_3293);
or U3438 (N_3438,N_3210,N_3179);
and U3439 (N_3439,N_3167,N_3287);
and U3440 (N_3440,N_3247,N_3273);
nor U3441 (N_3441,N_3222,N_3196);
and U3442 (N_3442,N_3239,N_3258);
nand U3443 (N_3443,N_3257,N_3254);
or U3444 (N_3444,N_3281,N_3194);
nand U3445 (N_3445,N_3287,N_3177);
xor U3446 (N_3446,N_3213,N_3219);
nor U3447 (N_3447,N_3227,N_3261);
nand U3448 (N_3448,N_3231,N_3281);
nand U3449 (N_3449,N_3228,N_3156);
nand U3450 (N_3450,N_3324,N_3369);
nand U3451 (N_3451,N_3339,N_3378);
xor U3452 (N_3452,N_3326,N_3446);
or U3453 (N_3453,N_3437,N_3314);
nand U3454 (N_3454,N_3439,N_3405);
nand U3455 (N_3455,N_3387,N_3331);
nor U3456 (N_3456,N_3409,N_3365);
nor U3457 (N_3457,N_3301,N_3367);
xor U3458 (N_3458,N_3370,N_3356);
or U3459 (N_3459,N_3375,N_3337);
xnor U3460 (N_3460,N_3410,N_3377);
or U3461 (N_3461,N_3380,N_3350);
or U3462 (N_3462,N_3388,N_3421);
or U3463 (N_3463,N_3354,N_3342);
nor U3464 (N_3464,N_3353,N_3442);
and U3465 (N_3465,N_3392,N_3319);
xnor U3466 (N_3466,N_3418,N_3344);
or U3467 (N_3467,N_3368,N_3399);
xor U3468 (N_3468,N_3389,N_3438);
nand U3469 (N_3469,N_3321,N_3335);
nor U3470 (N_3470,N_3414,N_3362);
nand U3471 (N_3471,N_3341,N_3376);
nor U3472 (N_3472,N_3309,N_3436);
xor U3473 (N_3473,N_3352,N_3360);
nor U3474 (N_3474,N_3310,N_3374);
and U3475 (N_3475,N_3325,N_3312);
xor U3476 (N_3476,N_3379,N_3385);
nand U3477 (N_3477,N_3359,N_3334);
and U3478 (N_3478,N_3364,N_3347);
xnor U3479 (N_3479,N_3402,N_3413);
nand U3480 (N_3480,N_3386,N_3373);
xnor U3481 (N_3481,N_3333,N_3419);
xor U3482 (N_3482,N_3403,N_3435);
xor U3483 (N_3483,N_3423,N_3441);
nor U3484 (N_3484,N_3431,N_3328);
xnor U3485 (N_3485,N_3327,N_3427);
nor U3486 (N_3486,N_3448,N_3434);
nand U3487 (N_3487,N_3306,N_3396);
nor U3488 (N_3488,N_3398,N_3372);
nor U3489 (N_3489,N_3322,N_3307);
or U3490 (N_3490,N_3323,N_3346);
or U3491 (N_3491,N_3336,N_3393);
and U3492 (N_3492,N_3440,N_3351);
and U3493 (N_3493,N_3308,N_3361);
or U3494 (N_3494,N_3381,N_3422);
nor U3495 (N_3495,N_3363,N_3340);
xor U3496 (N_3496,N_3444,N_3343);
or U3497 (N_3497,N_3330,N_3383);
nand U3498 (N_3498,N_3404,N_3411);
or U3499 (N_3499,N_3305,N_3428);
or U3500 (N_3500,N_3345,N_3420);
xnor U3501 (N_3501,N_3366,N_3394);
nand U3502 (N_3502,N_3449,N_3430);
xnor U3503 (N_3503,N_3315,N_3445);
xnor U3504 (N_3504,N_3417,N_3429);
or U3505 (N_3505,N_3432,N_3406);
xnor U3506 (N_3506,N_3400,N_3443);
or U3507 (N_3507,N_3303,N_3416);
xnor U3508 (N_3508,N_3302,N_3357);
nor U3509 (N_3509,N_3329,N_3397);
nor U3510 (N_3510,N_3425,N_3318);
nor U3511 (N_3511,N_3433,N_3316);
and U3512 (N_3512,N_3355,N_3408);
nor U3513 (N_3513,N_3395,N_3407);
nor U3514 (N_3514,N_3415,N_3384);
xor U3515 (N_3515,N_3300,N_3390);
nand U3516 (N_3516,N_3426,N_3382);
nand U3517 (N_3517,N_3304,N_3391);
nor U3518 (N_3518,N_3311,N_3317);
nor U3519 (N_3519,N_3401,N_3332);
and U3520 (N_3520,N_3412,N_3358);
nand U3521 (N_3521,N_3349,N_3338);
nand U3522 (N_3522,N_3447,N_3313);
nand U3523 (N_3523,N_3371,N_3320);
nor U3524 (N_3524,N_3424,N_3348);
nand U3525 (N_3525,N_3371,N_3439);
xnor U3526 (N_3526,N_3309,N_3333);
nor U3527 (N_3527,N_3432,N_3378);
nor U3528 (N_3528,N_3363,N_3373);
and U3529 (N_3529,N_3400,N_3385);
nor U3530 (N_3530,N_3397,N_3443);
and U3531 (N_3531,N_3338,N_3302);
or U3532 (N_3532,N_3347,N_3376);
and U3533 (N_3533,N_3349,N_3306);
or U3534 (N_3534,N_3323,N_3381);
or U3535 (N_3535,N_3440,N_3335);
and U3536 (N_3536,N_3359,N_3362);
nor U3537 (N_3537,N_3315,N_3310);
or U3538 (N_3538,N_3400,N_3344);
xnor U3539 (N_3539,N_3327,N_3344);
xor U3540 (N_3540,N_3379,N_3433);
nor U3541 (N_3541,N_3408,N_3339);
and U3542 (N_3542,N_3333,N_3410);
and U3543 (N_3543,N_3440,N_3448);
nor U3544 (N_3544,N_3349,N_3316);
nand U3545 (N_3545,N_3358,N_3307);
and U3546 (N_3546,N_3429,N_3432);
or U3547 (N_3547,N_3435,N_3421);
or U3548 (N_3548,N_3388,N_3358);
nand U3549 (N_3549,N_3440,N_3422);
or U3550 (N_3550,N_3400,N_3446);
nor U3551 (N_3551,N_3329,N_3392);
nor U3552 (N_3552,N_3374,N_3386);
xor U3553 (N_3553,N_3400,N_3306);
or U3554 (N_3554,N_3423,N_3399);
or U3555 (N_3555,N_3322,N_3399);
xor U3556 (N_3556,N_3388,N_3310);
and U3557 (N_3557,N_3304,N_3413);
xor U3558 (N_3558,N_3320,N_3425);
and U3559 (N_3559,N_3417,N_3394);
xor U3560 (N_3560,N_3351,N_3341);
xor U3561 (N_3561,N_3309,N_3328);
nor U3562 (N_3562,N_3368,N_3331);
nand U3563 (N_3563,N_3399,N_3372);
nor U3564 (N_3564,N_3374,N_3439);
and U3565 (N_3565,N_3392,N_3308);
xnor U3566 (N_3566,N_3394,N_3413);
xor U3567 (N_3567,N_3422,N_3322);
xnor U3568 (N_3568,N_3353,N_3307);
nand U3569 (N_3569,N_3448,N_3340);
or U3570 (N_3570,N_3364,N_3409);
nor U3571 (N_3571,N_3303,N_3430);
and U3572 (N_3572,N_3331,N_3380);
or U3573 (N_3573,N_3384,N_3354);
nor U3574 (N_3574,N_3433,N_3374);
and U3575 (N_3575,N_3317,N_3419);
nand U3576 (N_3576,N_3346,N_3306);
nand U3577 (N_3577,N_3370,N_3448);
and U3578 (N_3578,N_3426,N_3341);
xor U3579 (N_3579,N_3442,N_3302);
or U3580 (N_3580,N_3334,N_3378);
nand U3581 (N_3581,N_3399,N_3309);
and U3582 (N_3582,N_3382,N_3323);
or U3583 (N_3583,N_3318,N_3449);
and U3584 (N_3584,N_3376,N_3322);
nor U3585 (N_3585,N_3396,N_3310);
nor U3586 (N_3586,N_3444,N_3346);
nand U3587 (N_3587,N_3333,N_3358);
xor U3588 (N_3588,N_3341,N_3326);
xnor U3589 (N_3589,N_3434,N_3402);
nand U3590 (N_3590,N_3406,N_3390);
and U3591 (N_3591,N_3415,N_3315);
or U3592 (N_3592,N_3392,N_3390);
xnor U3593 (N_3593,N_3336,N_3408);
and U3594 (N_3594,N_3388,N_3390);
xnor U3595 (N_3595,N_3344,N_3364);
nor U3596 (N_3596,N_3328,N_3381);
or U3597 (N_3597,N_3411,N_3307);
nand U3598 (N_3598,N_3304,N_3306);
nand U3599 (N_3599,N_3445,N_3311);
nand U3600 (N_3600,N_3536,N_3463);
nand U3601 (N_3601,N_3503,N_3506);
or U3602 (N_3602,N_3585,N_3543);
or U3603 (N_3603,N_3470,N_3471);
xnor U3604 (N_3604,N_3532,N_3542);
nand U3605 (N_3605,N_3514,N_3566);
and U3606 (N_3606,N_3581,N_3509);
xor U3607 (N_3607,N_3592,N_3531);
nand U3608 (N_3608,N_3571,N_3504);
or U3609 (N_3609,N_3549,N_3553);
or U3610 (N_3610,N_3593,N_3483);
or U3611 (N_3611,N_3507,N_3526);
xnor U3612 (N_3612,N_3467,N_3584);
nand U3613 (N_3613,N_3573,N_3493);
nor U3614 (N_3614,N_3473,N_3569);
or U3615 (N_3615,N_3591,N_3494);
or U3616 (N_3616,N_3530,N_3466);
nor U3617 (N_3617,N_3484,N_3599);
and U3618 (N_3618,N_3598,N_3563);
xor U3619 (N_3619,N_3588,N_3562);
nand U3620 (N_3620,N_3476,N_3464);
xnor U3621 (N_3621,N_3469,N_3545);
xor U3622 (N_3622,N_3492,N_3564);
nand U3623 (N_3623,N_3512,N_3567);
nor U3624 (N_3624,N_3458,N_3583);
nand U3625 (N_3625,N_3475,N_3565);
xor U3626 (N_3626,N_3489,N_3570);
and U3627 (N_3627,N_3548,N_3559);
or U3628 (N_3628,N_3577,N_3544);
nand U3629 (N_3629,N_3534,N_3488);
nor U3630 (N_3630,N_3459,N_3552);
and U3631 (N_3631,N_3482,N_3537);
or U3632 (N_3632,N_3491,N_3462);
nor U3633 (N_3633,N_3511,N_3575);
xor U3634 (N_3634,N_3515,N_3551);
xnor U3635 (N_3635,N_3461,N_3500);
nand U3636 (N_3636,N_3510,N_3460);
xor U3637 (N_3637,N_3529,N_3582);
nor U3638 (N_3638,N_3453,N_3538);
nand U3639 (N_3639,N_3472,N_3596);
and U3640 (N_3640,N_3499,N_3540);
xnor U3641 (N_3641,N_3578,N_3521);
nand U3642 (N_3642,N_3527,N_3508);
and U3643 (N_3643,N_3525,N_3465);
and U3644 (N_3644,N_3502,N_3568);
or U3645 (N_3645,N_3523,N_3590);
nand U3646 (N_3646,N_3539,N_3541);
xor U3647 (N_3647,N_3496,N_3556);
nor U3648 (N_3648,N_3522,N_3478);
nand U3649 (N_3649,N_3513,N_3535);
nor U3650 (N_3650,N_3490,N_3477);
nand U3651 (N_3651,N_3474,N_3597);
or U3652 (N_3652,N_3457,N_3516);
xnor U3653 (N_3653,N_3547,N_3519);
nor U3654 (N_3654,N_3520,N_3524);
and U3655 (N_3655,N_3580,N_3586);
xor U3656 (N_3656,N_3572,N_3505);
or U3657 (N_3657,N_3550,N_3479);
xnor U3658 (N_3658,N_3451,N_3594);
nor U3659 (N_3659,N_3574,N_3558);
nand U3660 (N_3660,N_3554,N_3498);
nand U3661 (N_3661,N_3561,N_3487);
and U3662 (N_3662,N_3517,N_3454);
nor U3663 (N_3663,N_3555,N_3576);
nand U3664 (N_3664,N_3501,N_3495);
nand U3665 (N_3665,N_3589,N_3579);
xor U3666 (N_3666,N_3485,N_3557);
nand U3667 (N_3667,N_3533,N_3546);
and U3668 (N_3668,N_3486,N_3480);
or U3669 (N_3669,N_3595,N_3497);
nand U3670 (N_3670,N_3468,N_3481);
nand U3671 (N_3671,N_3452,N_3450);
xnor U3672 (N_3672,N_3528,N_3587);
or U3673 (N_3673,N_3560,N_3455);
xor U3674 (N_3674,N_3518,N_3456);
nand U3675 (N_3675,N_3467,N_3516);
nor U3676 (N_3676,N_3551,N_3595);
or U3677 (N_3677,N_3593,N_3463);
and U3678 (N_3678,N_3507,N_3584);
or U3679 (N_3679,N_3515,N_3595);
nor U3680 (N_3680,N_3559,N_3563);
and U3681 (N_3681,N_3497,N_3558);
nand U3682 (N_3682,N_3585,N_3466);
xnor U3683 (N_3683,N_3455,N_3554);
xnor U3684 (N_3684,N_3547,N_3584);
xnor U3685 (N_3685,N_3582,N_3514);
nand U3686 (N_3686,N_3508,N_3531);
nand U3687 (N_3687,N_3523,N_3525);
nand U3688 (N_3688,N_3537,N_3459);
xnor U3689 (N_3689,N_3578,N_3516);
xor U3690 (N_3690,N_3451,N_3457);
or U3691 (N_3691,N_3551,N_3470);
or U3692 (N_3692,N_3559,N_3573);
nor U3693 (N_3693,N_3481,N_3494);
xor U3694 (N_3694,N_3531,N_3570);
nor U3695 (N_3695,N_3494,N_3598);
nand U3696 (N_3696,N_3598,N_3490);
nand U3697 (N_3697,N_3561,N_3463);
or U3698 (N_3698,N_3497,N_3509);
nand U3699 (N_3699,N_3568,N_3516);
and U3700 (N_3700,N_3583,N_3547);
or U3701 (N_3701,N_3450,N_3587);
and U3702 (N_3702,N_3575,N_3460);
xor U3703 (N_3703,N_3522,N_3457);
and U3704 (N_3704,N_3533,N_3516);
or U3705 (N_3705,N_3454,N_3462);
nand U3706 (N_3706,N_3522,N_3463);
and U3707 (N_3707,N_3509,N_3594);
nand U3708 (N_3708,N_3575,N_3556);
nor U3709 (N_3709,N_3452,N_3556);
or U3710 (N_3710,N_3508,N_3574);
and U3711 (N_3711,N_3536,N_3540);
and U3712 (N_3712,N_3538,N_3504);
nor U3713 (N_3713,N_3507,N_3561);
nor U3714 (N_3714,N_3464,N_3473);
nor U3715 (N_3715,N_3599,N_3456);
xor U3716 (N_3716,N_3583,N_3534);
xor U3717 (N_3717,N_3453,N_3532);
nor U3718 (N_3718,N_3589,N_3486);
nand U3719 (N_3719,N_3494,N_3584);
nor U3720 (N_3720,N_3553,N_3490);
and U3721 (N_3721,N_3493,N_3556);
and U3722 (N_3722,N_3528,N_3450);
xor U3723 (N_3723,N_3507,N_3552);
and U3724 (N_3724,N_3459,N_3543);
or U3725 (N_3725,N_3582,N_3478);
nand U3726 (N_3726,N_3551,N_3482);
and U3727 (N_3727,N_3513,N_3525);
xnor U3728 (N_3728,N_3546,N_3475);
nand U3729 (N_3729,N_3487,N_3542);
nand U3730 (N_3730,N_3509,N_3513);
nor U3731 (N_3731,N_3481,N_3523);
nand U3732 (N_3732,N_3565,N_3499);
nand U3733 (N_3733,N_3469,N_3511);
or U3734 (N_3734,N_3459,N_3538);
or U3735 (N_3735,N_3562,N_3552);
or U3736 (N_3736,N_3587,N_3459);
xor U3737 (N_3737,N_3571,N_3529);
and U3738 (N_3738,N_3481,N_3502);
nand U3739 (N_3739,N_3511,N_3465);
nor U3740 (N_3740,N_3470,N_3506);
nand U3741 (N_3741,N_3490,N_3492);
nor U3742 (N_3742,N_3558,N_3545);
xor U3743 (N_3743,N_3554,N_3562);
or U3744 (N_3744,N_3572,N_3524);
or U3745 (N_3745,N_3596,N_3456);
nor U3746 (N_3746,N_3506,N_3550);
and U3747 (N_3747,N_3577,N_3510);
or U3748 (N_3748,N_3589,N_3468);
nand U3749 (N_3749,N_3549,N_3545);
and U3750 (N_3750,N_3647,N_3669);
or U3751 (N_3751,N_3741,N_3690);
nand U3752 (N_3752,N_3710,N_3682);
or U3753 (N_3753,N_3622,N_3630);
and U3754 (N_3754,N_3655,N_3617);
and U3755 (N_3755,N_3629,N_3715);
or U3756 (N_3756,N_3628,N_3624);
xnor U3757 (N_3757,N_3729,N_3658);
or U3758 (N_3758,N_3613,N_3651);
xor U3759 (N_3759,N_3625,N_3619);
nor U3760 (N_3760,N_3683,N_3616);
xor U3761 (N_3761,N_3699,N_3650);
or U3762 (N_3762,N_3737,N_3662);
or U3763 (N_3763,N_3640,N_3621);
and U3764 (N_3764,N_3646,N_3738);
nand U3765 (N_3765,N_3603,N_3745);
xnor U3766 (N_3766,N_3660,N_3703);
nand U3767 (N_3767,N_3749,N_3678);
xnor U3768 (N_3768,N_3709,N_3644);
nor U3769 (N_3769,N_3679,N_3702);
nor U3770 (N_3770,N_3673,N_3637);
and U3771 (N_3771,N_3747,N_3688);
nor U3772 (N_3772,N_3627,N_3611);
nor U3773 (N_3773,N_3674,N_3743);
nand U3774 (N_3774,N_3687,N_3689);
or U3775 (N_3775,N_3670,N_3663);
nand U3776 (N_3776,N_3618,N_3686);
or U3777 (N_3777,N_3626,N_3711);
nand U3778 (N_3778,N_3739,N_3634);
xnor U3779 (N_3779,N_3607,N_3666);
or U3780 (N_3780,N_3609,N_3684);
or U3781 (N_3781,N_3677,N_3615);
nor U3782 (N_3782,N_3604,N_3730);
or U3783 (N_3783,N_3631,N_3704);
nand U3784 (N_3784,N_3698,N_3659);
xnor U3785 (N_3785,N_3740,N_3692);
xnor U3786 (N_3786,N_3748,N_3693);
nand U3787 (N_3787,N_3671,N_3722);
xnor U3788 (N_3788,N_3732,N_3657);
nor U3789 (N_3789,N_3723,N_3742);
or U3790 (N_3790,N_3633,N_3705);
xnor U3791 (N_3791,N_3707,N_3665);
or U3792 (N_3792,N_3708,N_3733);
xor U3793 (N_3793,N_3717,N_3691);
nor U3794 (N_3794,N_3638,N_3639);
and U3795 (N_3795,N_3731,N_3721);
or U3796 (N_3796,N_3719,N_3680);
nor U3797 (N_3797,N_3701,N_3606);
and U3798 (N_3798,N_3668,N_3675);
or U3799 (N_3799,N_3696,N_3685);
nand U3800 (N_3800,N_3667,N_3661);
or U3801 (N_3801,N_3681,N_3720);
or U3802 (N_3802,N_3648,N_3713);
or U3803 (N_3803,N_3623,N_3605);
nor U3804 (N_3804,N_3718,N_3642);
or U3805 (N_3805,N_3727,N_3620);
xor U3806 (N_3806,N_3697,N_3716);
or U3807 (N_3807,N_3744,N_3734);
xor U3808 (N_3808,N_3712,N_3635);
nor U3809 (N_3809,N_3714,N_3700);
nor U3810 (N_3810,N_3724,N_3601);
or U3811 (N_3811,N_3608,N_3735);
nor U3812 (N_3812,N_3664,N_3652);
nor U3813 (N_3813,N_3672,N_3636);
or U3814 (N_3814,N_3641,N_3654);
and U3815 (N_3815,N_3649,N_3653);
xnor U3816 (N_3816,N_3725,N_3600);
xnor U3817 (N_3817,N_3695,N_3645);
nor U3818 (N_3818,N_3632,N_3643);
nor U3819 (N_3819,N_3676,N_3706);
nand U3820 (N_3820,N_3694,N_3736);
xor U3821 (N_3821,N_3610,N_3602);
and U3822 (N_3822,N_3656,N_3746);
xor U3823 (N_3823,N_3728,N_3612);
and U3824 (N_3824,N_3614,N_3726);
nor U3825 (N_3825,N_3736,N_3657);
nor U3826 (N_3826,N_3703,N_3608);
or U3827 (N_3827,N_3687,N_3600);
and U3828 (N_3828,N_3665,N_3619);
nand U3829 (N_3829,N_3673,N_3612);
nor U3830 (N_3830,N_3630,N_3707);
and U3831 (N_3831,N_3616,N_3725);
xnor U3832 (N_3832,N_3684,N_3668);
nor U3833 (N_3833,N_3696,N_3719);
and U3834 (N_3834,N_3719,N_3643);
nor U3835 (N_3835,N_3690,N_3725);
xor U3836 (N_3836,N_3702,N_3673);
and U3837 (N_3837,N_3629,N_3705);
and U3838 (N_3838,N_3694,N_3698);
and U3839 (N_3839,N_3680,N_3625);
nor U3840 (N_3840,N_3705,N_3605);
and U3841 (N_3841,N_3698,N_3669);
xnor U3842 (N_3842,N_3700,N_3628);
nor U3843 (N_3843,N_3740,N_3626);
nand U3844 (N_3844,N_3713,N_3691);
or U3845 (N_3845,N_3734,N_3624);
and U3846 (N_3846,N_3702,N_3648);
and U3847 (N_3847,N_3655,N_3611);
nor U3848 (N_3848,N_3745,N_3747);
or U3849 (N_3849,N_3605,N_3603);
nand U3850 (N_3850,N_3639,N_3704);
and U3851 (N_3851,N_3645,N_3659);
xor U3852 (N_3852,N_3632,N_3702);
nand U3853 (N_3853,N_3682,N_3640);
xnor U3854 (N_3854,N_3700,N_3650);
nand U3855 (N_3855,N_3736,N_3655);
and U3856 (N_3856,N_3731,N_3690);
or U3857 (N_3857,N_3602,N_3615);
xnor U3858 (N_3858,N_3649,N_3665);
nand U3859 (N_3859,N_3649,N_3678);
and U3860 (N_3860,N_3748,N_3603);
nand U3861 (N_3861,N_3705,N_3632);
or U3862 (N_3862,N_3647,N_3731);
and U3863 (N_3863,N_3741,N_3652);
or U3864 (N_3864,N_3686,N_3701);
and U3865 (N_3865,N_3645,N_3678);
nor U3866 (N_3866,N_3627,N_3616);
nand U3867 (N_3867,N_3647,N_3620);
or U3868 (N_3868,N_3731,N_3635);
nor U3869 (N_3869,N_3731,N_3703);
or U3870 (N_3870,N_3636,N_3712);
nand U3871 (N_3871,N_3610,N_3708);
or U3872 (N_3872,N_3719,N_3662);
or U3873 (N_3873,N_3630,N_3608);
xor U3874 (N_3874,N_3621,N_3722);
nor U3875 (N_3875,N_3701,N_3749);
and U3876 (N_3876,N_3724,N_3638);
nand U3877 (N_3877,N_3630,N_3746);
or U3878 (N_3878,N_3610,N_3624);
nor U3879 (N_3879,N_3675,N_3648);
xor U3880 (N_3880,N_3666,N_3609);
nand U3881 (N_3881,N_3639,N_3656);
or U3882 (N_3882,N_3650,N_3683);
or U3883 (N_3883,N_3607,N_3688);
and U3884 (N_3884,N_3695,N_3681);
or U3885 (N_3885,N_3727,N_3716);
nand U3886 (N_3886,N_3747,N_3608);
xnor U3887 (N_3887,N_3672,N_3716);
and U3888 (N_3888,N_3678,N_3625);
and U3889 (N_3889,N_3718,N_3720);
nor U3890 (N_3890,N_3614,N_3722);
or U3891 (N_3891,N_3743,N_3719);
xnor U3892 (N_3892,N_3653,N_3741);
xnor U3893 (N_3893,N_3727,N_3659);
and U3894 (N_3894,N_3630,N_3667);
and U3895 (N_3895,N_3724,N_3715);
nand U3896 (N_3896,N_3640,N_3668);
nor U3897 (N_3897,N_3707,N_3710);
nor U3898 (N_3898,N_3723,N_3735);
nand U3899 (N_3899,N_3671,N_3681);
nand U3900 (N_3900,N_3856,N_3866);
and U3901 (N_3901,N_3789,N_3784);
xnor U3902 (N_3902,N_3788,N_3799);
xnor U3903 (N_3903,N_3889,N_3793);
nor U3904 (N_3904,N_3800,N_3867);
xnor U3905 (N_3905,N_3781,N_3865);
xnor U3906 (N_3906,N_3824,N_3817);
or U3907 (N_3907,N_3869,N_3841);
and U3908 (N_3908,N_3887,N_3852);
xnor U3909 (N_3909,N_3755,N_3837);
xor U3910 (N_3910,N_3826,N_3830);
nor U3911 (N_3911,N_3884,N_3750);
nand U3912 (N_3912,N_3802,N_3758);
or U3913 (N_3913,N_3882,N_3779);
nand U3914 (N_3914,N_3792,N_3823);
and U3915 (N_3915,N_3893,N_3771);
or U3916 (N_3916,N_3829,N_3795);
nor U3917 (N_3917,N_3875,N_3871);
or U3918 (N_3918,N_3776,N_3854);
nand U3919 (N_3919,N_3870,N_3783);
nand U3920 (N_3920,N_3820,N_3818);
xnor U3921 (N_3921,N_3765,N_3896);
nand U3922 (N_3922,N_3751,N_3885);
nand U3923 (N_3923,N_3848,N_3801);
nor U3924 (N_3924,N_3874,N_3873);
nand U3925 (N_3925,N_3775,N_3844);
nor U3926 (N_3926,N_3794,N_3857);
xor U3927 (N_3927,N_3754,N_3862);
nor U3928 (N_3928,N_3768,N_3888);
xnor U3929 (N_3929,N_3787,N_3756);
nor U3930 (N_3930,N_3883,N_3859);
xnor U3931 (N_3931,N_3769,N_3813);
and U3932 (N_3932,N_3861,N_3809);
or U3933 (N_3933,N_3766,N_3786);
xnor U3934 (N_3934,N_3816,N_3880);
and U3935 (N_3935,N_3806,N_3827);
xnor U3936 (N_3936,N_3819,N_3894);
nand U3937 (N_3937,N_3855,N_3833);
and U3938 (N_3938,N_3782,N_3767);
or U3939 (N_3939,N_3890,N_3810);
xnor U3940 (N_3940,N_3835,N_3860);
and U3941 (N_3941,N_3847,N_3780);
or U3942 (N_3942,N_3778,N_3803);
nand U3943 (N_3943,N_3814,N_3838);
and U3944 (N_3944,N_3876,N_3853);
and U3945 (N_3945,N_3760,N_3864);
or U3946 (N_3946,N_3858,N_3834);
nand U3947 (N_3947,N_3851,N_3777);
or U3948 (N_3948,N_3831,N_3815);
or U3949 (N_3949,N_3822,N_3774);
and U3950 (N_3950,N_3761,N_3791);
and U3951 (N_3951,N_3821,N_3773);
nand U3952 (N_3952,N_3805,N_3899);
or U3953 (N_3953,N_3879,N_3886);
nand U3954 (N_3954,N_3849,N_3759);
nand U3955 (N_3955,N_3812,N_3763);
and U3956 (N_3956,N_3757,N_3846);
nand U3957 (N_3957,N_3796,N_3807);
and U3958 (N_3958,N_3877,N_3785);
nand U3959 (N_3959,N_3891,N_3762);
nand U3960 (N_3960,N_3811,N_3764);
and U3961 (N_3961,N_3878,N_3797);
and U3962 (N_3962,N_3842,N_3798);
nand U3963 (N_3963,N_3843,N_3825);
or U3964 (N_3964,N_3839,N_3898);
nand U3965 (N_3965,N_3863,N_3895);
or U3966 (N_3966,N_3881,N_3770);
and U3967 (N_3967,N_3808,N_3840);
xor U3968 (N_3968,N_3872,N_3828);
xnor U3969 (N_3969,N_3868,N_3804);
nand U3970 (N_3970,N_3892,N_3753);
or U3971 (N_3971,N_3850,N_3832);
or U3972 (N_3972,N_3845,N_3772);
nor U3973 (N_3973,N_3836,N_3752);
or U3974 (N_3974,N_3897,N_3790);
and U3975 (N_3975,N_3797,N_3888);
xor U3976 (N_3976,N_3893,N_3831);
xor U3977 (N_3977,N_3816,N_3779);
or U3978 (N_3978,N_3781,N_3764);
or U3979 (N_3979,N_3871,N_3803);
xnor U3980 (N_3980,N_3826,N_3765);
xnor U3981 (N_3981,N_3865,N_3760);
and U3982 (N_3982,N_3767,N_3798);
xor U3983 (N_3983,N_3801,N_3898);
xnor U3984 (N_3984,N_3787,N_3780);
and U3985 (N_3985,N_3869,N_3802);
nor U3986 (N_3986,N_3792,N_3764);
nor U3987 (N_3987,N_3852,N_3811);
or U3988 (N_3988,N_3778,N_3829);
nand U3989 (N_3989,N_3777,N_3874);
nor U3990 (N_3990,N_3771,N_3800);
and U3991 (N_3991,N_3895,N_3791);
and U3992 (N_3992,N_3837,N_3768);
xnor U3993 (N_3993,N_3877,N_3821);
nor U3994 (N_3994,N_3798,N_3861);
xnor U3995 (N_3995,N_3853,N_3784);
nand U3996 (N_3996,N_3798,N_3823);
xor U3997 (N_3997,N_3838,N_3899);
xnor U3998 (N_3998,N_3831,N_3760);
or U3999 (N_3999,N_3755,N_3761);
nor U4000 (N_4000,N_3852,N_3897);
and U4001 (N_4001,N_3761,N_3811);
nor U4002 (N_4002,N_3890,N_3796);
nor U4003 (N_4003,N_3899,N_3832);
nor U4004 (N_4004,N_3756,N_3814);
nor U4005 (N_4005,N_3886,N_3853);
nor U4006 (N_4006,N_3797,N_3753);
or U4007 (N_4007,N_3861,N_3836);
nor U4008 (N_4008,N_3884,N_3866);
or U4009 (N_4009,N_3855,N_3762);
and U4010 (N_4010,N_3884,N_3898);
nand U4011 (N_4011,N_3783,N_3856);
xnor U4012 (N_4012,N_3856,N_3775);
nand U4013 (N_4013,N_3831,N_3889);
xnor U4014 (N_4014,N_3825,N_3794);
or U4015 (N_4015,N_3829,N_3897);
or U4016 (N_4016,N_3894,N_3794);
and U4017 (N_4017,N_3868,N_3852);
nor U4018 (N_4018,N_3832,N_3785);
xor U4019 (N_4019,N_3775,N_3886);
nor U4020 (N_4020,N_3765,N_3875);
xnor U4021 (N_4021,N_3764,N_3789);
nor U4022 (N_4022,N_3858,N_3852);
xor U4023 (N_4023,N_3750,N_3752);
nor U4024 (N_4024,N_3753,N_3826);
xnor U4025 (N_4025,N_3850,N_3847);
or U4026 (N_4026,N_3768,N_3845);
and U4027 (N_4027,N_3786,N_3772);
xor U4028 (N_4028,N_3819,N_3886);
and U4029 (N_4029,N_3831,N_3757);
or U4030 (N_4030,N_3847,N_3808);
or U4031 (N_4031,N_3840,N_3761);
nand U4032 (N_4032,N_3867,N_3791);
and U4033 (N_4033,N_3785,N_3765);
nor U4034 (N_4034,N_3868,N_3837);
xnor U4035 (N_4035,N_3829,N_3871);
xor U4036 (N_4036,N_3812,N_3831);
or U4037 (N_4037,N_3876,N_3837);
xor U4038 (N_4038,N_3894,N_3776);
and U4039 (N_4039,N_3768,N_3834);
nor U4040 (N_4040,N_3753,N_3771);
and U4041 (N_4041,N_3801,N_3779);
nor U4042 (N_4042,N_3870,N_3899);
or U4043 (N_4043,N_3780,N_3821);
and U4044 (N_4044,N_3777,N_3857);
nand U4045 (N_4045,N_3787,N_3862);
nor U4046 (N_4046,N_3876,N_3764);
nor U4047 (N_4047,N_3882,N_3876);
nand U4048 (N_4048,N_3804,N_3797);
and U4049 (N_4049,N_3875,N_3873);
nand U4050 (N_4050,N_3975,N_3998);
or U4051 (N_4051,N_3923,N_3965);
or U4052 (N_4052,N_3929,N_3931);
nor U4053 (N_4053,N_3952,N_3963);
nand U4054 (N_4054,N_3984,N_4014);
nor U4055 (N_4055,N_4044,N_3964);
nor U4056 (N_4056,N_4031,N_3913);
nor U4057 (N_4057,N_4022,N_3976);
and U4058 (N_4058,N_3908,N_3907);
xnor U4059 (N_4059,N_3972,N_3999);
nand U4060 (N_4060,N_3971,N_4034);
or U4061 (N_4061,N_3902,N_3906);
and U4062 (N_4062,N_3943,N_4024);
and U4063 (N_4063,N_3916,N_4012);
or U4064 (N_4064,N_4042,N_4043);
xnor U4065 (N_4065,N_3977,N_3942);
nor U4066 (N_4066,N_4028,N_3918);
or U4067 (N_4067,N_4021,N_3949);
and U4068 (N_4068,N_3983,N_4049);
xnor U4069 (N_4069,N_3950,N_3982);
and U4070 (N_4070,N_3968,N_3980);
nor U4071 (N_4071,N_3930,N_4037);
and U4072 (N_4072,N_4036,N_4032);
or U4073 (N_4073,N_3910,N_3936);
and U4074 (N_4074,N_3961,N_3941);
nor U4075 (N_4075,N_3915,N_4001);
xor U4076 (N_4076,N_4041,N_3978);
and U4077 (N_4077,N_4008,N_4033);
and U4078 (N_4078,N_3917,N_4025);
xor U4079 (N_4079,N_3985,N_3997);
or U4080 (N_4080,N_4029,N_3945);
nor U4081 (N_4081,N_4035,N_3947);
nand U4082 (N_4082,N_3900,N_4010);
or U4083 (N_4083,N_3990,N_4047);
or U4084 (N_4084,N_3996,N_4023);
or U4085 (N_4085,N_3987,N_4048);
and U4086 (N_4086,N_3970,N_3932);
xnor U4087 (N_4087,N_3955,N_3909);
or U4088 (N_4088,N_4026,N_3925);
nand U4089 (N_4089,N_3911,N_3974);
and U4090 (N_4090,N_3979,N_3928);
nor U4091 (N_4091,N_4011,N_3921);
or U4092 (N_4092,N_3988,N_4039);
or U4093 (N_4093,N_4045,N_4018);
and U4094 (N_4094,N_3927,N_4000);
or U4095 (N_4095,N_4004,N_3994);
nor U4096 (N_4096,N_4020,N_3956);
nor U4097 (N_4097,N_3934,N_4009);
nor U4098 (N_4098,N_3926,N_3914);
xnor U4099 (N_4099,N_4016,N_4013);
or U4100 (N_4100,N_3937,N_3924);
xnor U4101 (N_4101,N_3940,N_3981);
or U4102 (N_4102,N_3957,N_4006);
or U4103 (N_4103,N_3986,N_3962);
xnor U4104 (N_4104,N_3944,N_3901);
nand U4105 (N_4105,N_3948,N_4046);
nand U4106 (N_4106,N_3935,N_3959);
nor U4107 (N_4107,N_3903,N_3933);
and U4108 (N_4108,N_3905,N_4019);
nand U4109 (N_4109,N_4038,N_3991);
and U4110 (N_4110,N_3993,N_3912);
nor U4111 (N_4111,N_4015,N_3960);
nand U4112 (N_4112,N_4040,N_3966);
or U4113 (N_4113,N_4017,N_3904);
and U4114 (N_4114,N_3919,N_3967);
xor U4115 (N_4115,N_3954,N_3939);
xor U4116 (N_4116,N_4003,N_3953);
or U4117 (N_4117,N_3920,N_4002);
and U4118 (N_4118,N_4005,N_3922);
or U4119 (N_4119,N_3951,N_3938);
and U4120 (N_4120,N_4027,N_3958);
xnor U4121 (N_4121,N_3989,N_3995);
or U4122 (N_4122,N_3992,N_4007);
and U4123 (N_4123,N_3969,N_4030);
xnor U4124 (N_4124,N_3973,N_3946);
or U4125 (N_4125,N_3980,N_3937);
and U4126 (N_4126,N_3912,N_3999);
and U4127 (N_4127,N_3937,N_3999);
or U4128 (N_4128,N_3972,N_3933);
and U4129 (N_4129,N_4003,N_4005);
xor U4130 (N_4130,N_4012,N_3989);
and U4131 (N_4131,N_3968,N_4025);
xnor U4132 (N_4132,N_3973,N_3952);
and U4133 (N_4133,N_3966,N_3911);
xnor U4134 (N_4134,N_3967,N_3916);
or U4135 (N_4135,N_4040,N_3953);
nand U4136 (N_4136,N_3992,N_3958);
xnor U4137 (N_4137,N_3971,N_4023);
xor U4138 (N_4138,N_3966,N_3930);
xor U4139 (N_4139,N_3961,N_4026);
xor U4140 (N_4140,N_3940,N_4007);
and U4141 (N_4141,N_4014,N_4022);
nand U4142 (N_4142,N_4011,N_4034);
or U4143 (N_4143,N_4036,N_3926);
or U4144 (N_4144,N_3905,N_4009);
nand U4145 (N_4145,N_4015,N_3994);
and U4146 (N_4146,N_3934,N_3939);
xor U4147 (N_4147,N_3933,N_4020);
nand U4148 (N_4148,N_3928,N_4049);
xnor U4149 (N_4149,N_4037,N_3915);
nor U4150 (N_4150,N_3934,N_3919);
and U4151 (N_4151,N_3956,N_4018);
or U4152 (N_4152,N_3905,N_4036);
nor U4153 (N_4153,N_3941,N_3982);
nand U4154 (N_4154,N_4012,N_4027);
or U4155 (N_4155,N_3905,N_4045);
xnor U4156 (N_4156,N_3980,N_3961);
and U4157 (N_4157,N_4022,N_3956);
xnor U4158 (N_4158,N_3900,N_4049);
and U4159 (N_4159,N_3927,N_4019);
nand U4160 (N_4160,N_3916,N_3953);
or U4161 (N_4161,N_4040,N_3904);
xnor U4162 (N_4162,N_3969,N_3945);
xnor U4163 (N_4163,N_3959,N_3982);
nand U4164 (N_4164,N_3980,N_4032);
xor U4165 (N_4165,N_3986,N_3984);
and U4166 (N_4166,N_3919,N_4001);
or U4167 (N_4167,N_3924,N_3930);
and U4168 (N_4168,N_3985,N_4018);
xor U4169 (N_4169,N_3979,N_3943);
and U4170 (N_4170,N_3938,N_3901);
xor U4171 (N_4171,N_4033,N_3940);
or U4172 (N_4172,N_3925,N_3938);
xor U4173 (N_4173,N_3987,N_3943);
xnor U4174 (N_4174,N_3937,N_4026);
xnor U4175 (N_4175,N_3955,N_3957);
nand U4176 (N_4176,N_3971,N_3904);
nor U4177 (N_4177,N_3992,N_3948);
and U4178 (N_4178,N_3962,N_3998);
or U4179 (N_4179,N_3933,N_3917);
nand U4180 (N_4180,N_3909,N_3951);
and U4181 (N_4181,N_3919,N_4000);
or U4182 (N_4182,N_3953,N_3974);
or U4183 (N_4183,N_3968,N_3991);
nand U4184 (N_4184,N_3962,N_3929);
nor U4185 (N_4185,N_3978,N_3923);
nand U4186 (N_4186,N_4006,N_4034);
or U4187 (N_4187,N_4038,N_3972);
or U4188 (N_4188,N_4037,N_3919);
nand U4189 (N_4189,N_4014,N_4032);
nor U4190 (N_4190,N_3968,N_3958);
and U4191 (N_4191,N_3944,N_3983);
xor U4192 (N_4192,N_3947,N_3914);
nand U4193 (N_4193,N_3905,N_3914);
nor U4194 (N_4194,N_4004,N_3932);
nor U4195 (N_4195,N_3970,N_3900);
and U4196 (N_4196,N_3999,N_3982);
and U4197 (N_4197,N_4013,N_4031);
xnor U4198 (N_4198,N_3986,N_3914);
nor U4199 (N_4199,N_3954,N_3970);
nand U4200 (N_4200,N_4069,N_4079);
nand U4201 (N_4201,N_4161,N_4170);
and U4202 (N_4202,N_4075,N_4142);
nand U4203 (N_4203,N_4095,N_4154);
xnor U4204 (N_4204,N_4087,N_4121);
and U4205 (N_4205,N_4058,N_4099);
nor U4206 (N_4206,N_4183,N_4110);
and U4207 (N_4207,N_4074,N_4061);
nor U4208 (N_4208,N_4175,N_4182);
xor U4209 (N_4209,N_4134,N_4130);
and U4210 (N_4210,N_4153,N_4186);
or U4211 (N_4211,N_4173,N_4148);
and U4212 (N_4212,N_4111,N_4135);
xor U4213 (N_4213,N_4125,N_4167);
nand U4214 (N_4214,N_4184,N_4191);
and U4215 (N_4215,N_4198,N_4098);
and U4216 (N_4216,N_4185,N_4193);
xor U4217 (N_4217,N_4101,N_4080);
and U4218 (N_4218,N_4179,N_4053);
nor U4219 (N_4219,N_4070,N_4122);
and U4220 (N_4220,N_4165,N_4078);
or U4221 (N_4221,N_4107,N_4196);
and U4222 (N_4222,N_4166,N_4199);
nand U4223 (N_4223,N_4155,N_4068);
or U4224 (N_4224,N_4190,N_4131);
nand U4225 (N_4225,N_4093,N_4141);
nor U4226 (N_4226,N_4092,N_4126);
or U4227 (N_4227,N_4137,N_4160);
xnor U4228 (N_4228,N_4120,N_4174);
xnor U4229 (N_4229,N_4071,N_4172);
nand U4230 (N_4230,N_4082,N_4117);
or U4231 (N_4231,N_4143,N_4089);
nor U4232 (N_4232,N_4189,N_4194);
or U4233 (N_4233,N_4171,N_4114);
nand U4234 (N_4234,N_4077,N_4139);
or U4235 (N_4235,N_4119,N_4138);
nand U4236 (N_4236,N_4094,N_4059);
nand U4237 (N_4237,N_4158,N_4106);
or U4238 (N_4238,N_4197,N_4133);
and U4239 (N_4239,N_4112,N_4109);
nor U4240 (N_4240,N_4064,N_4118);
and U4241 (N_4241,N_4067,N_4051);
or U4242 (N_4242,N_4123,N_4054);
xor U4243 (N_4243,N_4090,N_4084);
nor U4244 (N_4244,N_4105,N_4144);
and U4245 (N_4245,N_4124,N_4136);
xnor U4246 (N_4246,N_4177,N_4066);
nor U4247 (N_4247,N_4188,N_4086);
and U4248 (N_4248,N_4063,N_4073);
nand U4249 (N_4249,N_4147,N_4052);
xor U4250 (N_4250,N_4176,N_4163);
nand U4251 (N_4251,N_4088,N_4057);
and U4252 (N_4252,N_4178,N_4076);
or U4253 (N_4253,N_4091,N_4151);
or U4254 (N_4254,N_4162,N_4192);
nor U4255 (N_4255,N_4181,N_4157);
nor U4256 (N_4256,N_4168,N_4103);
nand U4257 (N_4257,N_4156,N_4146);
and U4258 (N_4258,N_4072,N_4060);
and U4259 (N_4259,N_4083,N_4104);
nand U4260 (N_4260,N_4100,N_4132);
nand U4261 (N_4261,N_4129,N_4164);
and U4262 (N_4262,N_4062,N_4127);
nor U4263 (N_4263,N_4097,N_4056);
xnor U4264 (N_4264,N_4145,N_4096);
and U4265 (N_4265,N_4115,N_4140);
xnor U4266 (N_4266,N_4108,N_4081);
or U4267 (N_4267,N_4065,N_4180);
xnor U4268 (N_4268,N_4195,N_4152);
nand U4269 (N_4269,N_4116,N_4050);
nand U4270 (N_4270,N_4113,N_4128);
nand U4271 (N_4271,N_4149,N_4102);
nor U4272 (N_4272,N_4187,N_4085);
and U4273 (N_4273,N_4169,N_4055);
nor U4274 (N_4274,N_4150,N_4159);
and U4275 (N_4275,N_4085,N_4138);
or U4276 (N_4276,N_4139,N_4198);
xor U4277 (N_4277,N_4086,N_4130);
nor U4278 (N_4278,N_4090,N_4063);
or U4279 (N_4279,N_4060,N_4183);
xnor U4280 (N_4280,N_4130,N_4162);
or U4281 (N_4281,N_4186,N_4095);
nor U4282 (N_4282,N_4140,N_4098);
and U4283 (N_4283,N_4175,N_4093);
and U4284 (N_4284,N_4125,N_4078);
nor U4285 (N_4285,N_4106,N_4183);
nor U4286 (N_4286,N_4080,N_4059);
xor U4287 (N_4287,N_4109,N_4158);
and U4288 (N_4288,N_4112,N_4187);
nor U4289 (N_4289,N_4185,N_4127);
nor U4290 (N_4290,N_4154,N_4090);
nand U4291 (N_4291,N_4110,N_4052);
and U4292 (N_4292,N_4199,N_4131);
nor U4293 (N_4293,N_4127,N_4074);
or U4294 (N_4294,N_4072,N_4138);
and U4295 (N_4295,N_4141,N_4073);
xnor U4296 (N_4296,N_4165,N_4054);
nor U4297 (N_4297,N_4164,N_4182);
xor U4298 (N_4298,N_4195,N_4111);
nor U4299 (N_4299,N_4152,N_4134);
nand U4300 (N_4300,N_4170,N_4147);
and U4301 (N_4301,N_4150,N_4099);
xor U4302 (N_4302,N_4063,N_4086);
or U4303 (N_4303,N_4080,N_4122);
or U4304 (N_4304,N_4175,N_4116);
and U4305 (N_4305,N_4162,N_4092);
and U4306 (N_4306,N_4189,N_4156);
nand U4307 (N_4307,N_4175,N_4090);
nor U4308 (N_4308,N_4185,N_4068);
nand U4309 (N_4309,N_4183,N_4087);
nand U4310 (N_4310,N_4108,N_4059);
nor U4311 (N_4311,N_4110,N_4126);
xor U4312 (N_4312,N_4109,N_4055);
nor U4313 (N_4313,N_4153,N_4162);
and U4314 (N_4314,N_4075,N_4091);
nor U4315 (N_4315,N_4075,N_4134);
or U4316 (N_4316,N_4138,N_4091);
nor U4317 (N_4317,N_4122,N_4104);
or U4318 (N_4318,N_4096,N_4132);
or U4319 (N_4319,N_4191,N_4174);
xnor U4320 (N_4320,N_4138,N_4090);
nand U4321 (N_4321,N_4132,N_4164);
nand U4322 (N_4322,N_4130,N_4059);
and U4323 (N_4323,N_4172,N_4079);
and U4324 (N_4324,N_4062,N_4069);
xnor U4325 (N_4325,N_4089,N_4111);
or U4326 (N_4326,N_4183,N_4178);
and U4327 (N_4327,N_4078,N_4172);
nand U4328 (N_4328,N_4170,N_4071);
nor U4329 (N_4329,N_4151,N_4121);
nand U4330 (N_4330,N_4111,N_4077);
and U4331 (N_4331,N_4054,N_4163);
or U4332 (N_4332,N_4156,N_4169);
nor U4333 (N_4333,N_4168,N_4092);
nand U4334 (N_4334,N_4134,N_4064);
xor U4335 (N_4335,N_4172,N_4099);
nand U4336 (N_4336,N_4175,N_4055);
nand U4337 (N_4337,N_4091,N_4144);
and U4338 (N_4338,N_4101,N_4062);
nand U4339 (N_4339,N_4138,N_4083);
and U4340 (N_4340,N_4146,N_4149);
xor U4341 (N_4341,N_4070,N_4114);
or U4342 (N_4342,N_4180,N_4061);
and U4343 (N_4343,N_4191,N_4062);
or U4344 (N_4344,N_4111,N_4121);
xor U4345 (N_4345,N_4132,N_4056);
xor U4346 (N_4346,N_4059,N_4141);
or U4347 (N_4347,N_4188,N_4183);
or U4348 (N_4348,N_4064,N_4107);
and U4349 (N_4349,N_4068,N_4119);
nor U4350 (N_4350,N_4212,N_4214);
nor U4351 (N_4351,N_4269,N_4310);
nand U4352 (N_4352,N_4288,N_4312);
nand U4353 (N_4353,N_4264,N_4235);
nand U4354 (N_4354,N_4309,N_4238);
xnor U4355 (N_4355,N_4254,N_4299);
nor U4356 (N_4356,N_4329,N_4341);
and U4357 (N_4357,N_4291,N_4272);
xnor U4358 (N_4358,N_4339,N_4227);
nor U4359 (N_4359,N_4328,N_4346);
and U4360 (N_4360,N_4295,N_4249);
xnor U4361 (N_4361,N_4278,N_4216);
and U4362 (N_4362,N_4266,N_4302);
nand U4363 (N_4363,N_4300,N_4226);
xnor U4364 (N_4364,N_4204,N_4298);
nand U4365 (N_4365,N_4247,N_4200);
or U4366 (N_4366,N_4338,N_4289);
nor U4367 (N_4367,N_4306,N_4316);
nor U4368 (N_4368,N_4228,N_4245);
and U4369 (N_4369,N_4262,N_4275);
nand U4370 (N_4370,N_4243,N_4286);
nor U4371 (N_4371,N_4342,N_4336);
or U4372 (N_4372,N_4301,N_4236);
xnor U4373 (N_4373,N_4280,N_4232);
and U4374 (N_4374,N_4274,N_4250);
or U4375 (N_4375,N_4209,N_4284);
and U4376 (N_4376,N_4206,N_4322);
xnor U4377 (N_4377,N_4282,N_4205);
nand U4378 (N_4378,N_4308,N_4317);
and U4379 (N_4379,N_4244,N_4315);
nor U4380 (N_4380,N_4305,N_4287);
and U4381 (N_4381,N_4268,N_4265);
nor U4382 (N_4382,N_4248,N_4340);
xor U4383 (N_4383,N_4290,N_4337);
nor U4384 (N_4384,N_4331,N_4324);
nor U4385 (N_4385,N_4241,N_4217);
nor U4386 (N_4386,N_4332,N_4321);
xor U4387 (N_4387,N_4230,N_4325);
nand U4388 (N_4388,N_4323,N_4258);
nand U4389 (N_4389,N_4320,N_4344);
and U4390 (N_4390,N_4314,N_4240);
xnor U4391 (N_4391,N_4257,N_4237);
or U4392 (N_4392,N_4319,N_4256);
and U4393 (N_4393,N_4273,N_4239);
and U4394 (N_4394,N_4215,N_4219);
or U4395 (N_4395,N_4267,N_4297);
and U4396 (N_4396,N_4277,N_4220);
nand U4397 (N_4397,N_4234,N_4279);
and U4398 (N_4398,N_4229,N_4221);
nor U4399 (N_4399,N_4311,N_4307);
or U4400 (N_4400,N_4296,N_4222);
nand U4401 (N_4401,N_4313,N_4276);
nand U4402 (N_4402,N_4218,N_4255);
or U4403 (N_4403,N_4292,N_4202);
or U4404 (N_4404,N_4330,N_4260);
and U4405 (N_4405,N_4259,N_4285);
or U4406 (N_4406,N_4203,N_4263);
and U4407 (N_4407,N_4345,N_4211);
nor U4408 (N_4408,N_4343,N_4294);
xor U4409 (N_4409,N_4270,N_4246);
or U4410 (N_4410,N_4261,N_4210);
xor U4411 (N_4411,N_4348,N_4347);
nor U4412 (N_4412,N_4253,N_4303);
nand U4413 (N_4413,N_4333,N_4349);
or U4414 (N_4414,N_4293,N_4326);
or U4415 (N_4415,N_4281,N_4208);
nor U4416 (N_4416,N_4242,N_4252);
xnor U4417 (N_4417,N_4201,N_4318);
nand U4418 (N_4418,N_4335,N_4251);
and U4419 (N_4419,N_4327,N_4231);
xnor U4420 (N_4420,N_4213,N_4334);
or U4421 (N_4421,N_4224,N_4225);
and U4422 (N_4422,N_4283,N_4304);
or U4423 (N_4423,N_4223,N_4207);
and U4424 (N_4424,N_4233,N_4271);
xor U4425 (N_4425,N_4312,N_4310);
and U4426 (N_4426,N_4271,N_4220);
nand U4427 (N_4427,N_4219,N_4297);
nor U4428 (N_4428,N_4254,N_4218);
or U4429 (N_4429,N_4326,N_4299);
nor U4430 (N_4430,N_4261,N_4332);
nand U4431 (N_4431,N_4341,N_4228);
or U4432 (N_4432,N_4234,N_4245);
nor U4433 (N_4433,N_4258,N_4209);
xnor U4434 (N_4434,N_4298,N_4308);
or U4435 (N_4435,N_4221,N_4336);
xnor U4436 (N_4436,N_4274,N_4349);
xor U4437 (N_4437,N_4206,N_4234);
and U4438 (N_4438,N_4220,N_4218);
xor U4439 (N_4439,N_4235,N_4281);
xor U4440 (N_4440,N_4313,N_4346);
nand U4441 (N_4441,N_4306,N_4313);
and U4442 (N_4442,N_4249,N_4236);
nand U4443 (N_4443,N_4271,N_4218);
and U4444 (N_4444,N_4292,N_4338);
nor U4445 (N_4445,N_4335,N_4343);
nand U4446 (N_4446,N_4294,N_4230);
and U4447 (N_4447,N_4332,N_4202);
and U4448 (N_4448,N_4310,N_4283);
or U4449 (N_4449,N_4266,N_4297);
and U4450 (N_4450,N_4260,N_4207);
and U4451 (N_4451,N_4347,N_4252);
nor U4452 (N_4452,N_4265,N_4341);
nand U4453 (N_4453,N_4324,N_4252);
xnor U4454 (N_4454,N_4328,N_4326);
or U4455 (N_4455,N_4288,N_4297);
and U4456 (N_4456,N_4301,N_4347);
and U4457 (N_4457,N_4336,N_4309);
nor U4458 (N_4458,N_4274,N_4324);
nor U4459 (N_4459,N_4277,N_4215);
nand U4460 (N_4460,N_4216,N_4264);
and U4461 (N_4461,N_4311,N_4346);
xor U4462 (N_4462,N_4325,N_4249);
and U4463 (N_4463,N_4282,N_4216);
nand U4464 (N_4464,N_4284,N_4294);
and U4465 (N_4465,N_4209,N_4243);
or U4466 (N_4466,N_4227,N_4323);
nor U4467 (N_4467,N_4251,N_4266);
and U4468 (N_4468,N_4335,N_4264);
nand U4469 (N_4469,N_4308,N_4295);
nor U4470 (N_4470,N_4256,N_4331);
and U4471 (N_4471,N_4273,N_4277);
nand U4472 (N_4472,N_4269,N_4203);
and U4473 (N_4473,N_4220,N_4302);
xnor U4474 (N_4474,N_4242,N_4220);
nor U4475 (N_4475,N_4260,N_4301);
nor U4476 (N_4476,N_4238,N_4276);
or U4477 (N_4477,N_4330,N_4285);
nand U4478 (N_4478,N_4327,N_4296);
nand U4479 (N_4479,N_4346,N_4227);
and U4480 (N_4480,N_4254,N_4335);
nand U4481 (N_4481,N_4201,N_4295);
and U4482 (N_4482,N_4267,N_4309);
or U4483 (N_4483,N_4208,N_4239);
xor U4484 (N_4484,N_4235,N_4203);
and U4485 (N_4485,N_4211,N_4256);
or U4486 (N_4486,N_4304,N_4326);
xnor U4487 (N_4487,N_4240,N_4299);
xor U4488 (N_4488,N_4301,N_4267);
or U4489 (N_4489,N_4329,N_4236);
nand U4490 (N_4490,N_4332,N_4293);
or U4491 (N_4491,N_4342,N_4229);
and U4492 (N_4492,N_4256,N_4299);
nor U4493 (N_4493,N_4345,N_4200);
and U4494 (N_4494,N_4295,N_4242);
nand U4495 (N_4495,N_4254,N_4340);
nand U4496 (N_4496,N_4234,N_4230);
nand U4497 (N_4497,N_4222,N_4333);
nor U4498 (N_4498,N_4231,N_4213);
nand U4499 (N_4499,N_4307,N_4248);
or U4500 (N_4500,N_4360,N_4403);
nor U4501 (N_4501,N_4420,N_4463);
or U4502 (N_4502,N_4369,N_4353);
nand U4503 (N_4503,N_4477,N_4481);
or U4504 (N_4504,N_4386,N_4478);
nor U4505 (N_4505,N_4475,N_4370);
or U4506 (N_4506,N_4492,N_4457);
nor U4507 (N_4507,N_4367,N_4355);
and U4508 (N_4508,N_4452,N_4398);
nand U4509 (N_4509,N_4377,N_4372);
xnor U4510 (N_4510,N_4381,N_4467);
or U4511 (N_4511,N_4497,N_4417);
xnor U4512 (N_4512,N_4416,N_4412);
nor U4513 (N_4513,N_4484,N_4418);
nor U4514 (N_4514,N_4451,N_4486);
xor U4515 (N_4515,N_4405,N_4365);
or U4516 (N_4516,N_4401,N_4385);
nor U4517 (N_4517,N_4395,N_4436);
nor U4518 (N_4518,N_4495,N_4356);
nand U4519 (N_4519,N_4430,N_4396);
or U4520 (N_4520,N_4358,N_4421);
and U4521 (N_4521,N_4474,N_4460);
and U4522 (N_4522,N_4489,N_4465);
xor U4523 (N_4523,N_4456,N_4482);
xor U4524 (N_4524,N_4399,N_4350);
nand U4525 (N_4525,N_4422,N_4490);
nand U4526 (N_4526,N_4472,N_4443);
nor U4527 (N_4527,N_4373,N_4404);
xor U4528 (N_4528,N_4476,N_4409);
xor U4529 (N_4529,N_4487,N_4485);
and U4530 (N_4530,N_4442,N_4455);
nand U4531 (N_4531,N_4471,N_4454);
nor U4532 (N_4532,N_4453,N_4480);
or U4533 (N_4533,N_4473,N_4446);
xnor U4534 (N_4534,N_4419,N_4364);
nor U4535 (N_4535,N_4359,N_4352);
xor U4536 (N_4536,N_4444,N_4408);
or U4537 (N_4537,N_4423,N_4392);
and U4538 (N_4538,N_4391,N_4464);
nand U4539 (N_4539,N_4429,N_4382);
and U4540 (N_4540,N_4461,N_4435);
xor U4541 (N_4541,N_4491,N_4438);
or U4542 (N_4542,N_4431,N_4397);
and U4543 (N_4543,N_4388,N_4493);
or U4544 (N_4544,N_4368,N_4494);
and U4545 (N_4545,N_4439,N_4499);
and U4546 (N_4546,N_4462,N_4387);
or U4547 (N_4547,N_4406,N_4378);
and U4548 (N_4548,N_4410,N_4459);
xnor U4549 (N_4549,N_4374,N_4483);
xnor U4550 (N_4550,N_4432,N_4414);
and U4551 (N_4551,N_4424,N_4402);
and U4552 (N_4552,N_4389,N_4411);
nor U4553 (N_4553,N_4447,N_4470);
and U4554 (N_4554,N_4498,N_4362);
or U4555 (N_4555,N_4357,N_4415);
and U4556 (N_4556,N_4383,N_4466);
nand U4557 (N_4557,N_4390,N_4400);
or U4558 (N_4558,N_4394,N_4380);
xnor U4559 (N_4559,N_4363,N_4448);
xnor U4560 (N_4560,N_4441,N_4427);
xnor U4561 (N_4561,N_4407,N_4440);
or U4562 (N_4562,N_4393,N_4428);
nor U4563 (N_4563,N_4426,N_4437);
nand U4564 (N_4564,N_4445,N_4434);
nand U4565 (N_4565,N_4361,N_4458);
or U4566 (N_4566,N_4371,N_4413);
nor U4567 (N_4567,N_4425,N_4354);
or U4568 (N_4568,N_4375,N_4379);
nor U4569 (N_4569,N_4488,N_4496);
xnor U4570 (N_4570,N_4376,N_4449);
and U4571 (N_4571,N_4469,N_4366);
nor U4572 (N_4572,N_4384,N_4433);
or U4573 (N_4573,N_4479,N_4468);
or U4574 (N_4574,N_4450,N_4351);
and U4575 (N_4575,N_4433,N_4372);
nand U4576 (N_4576,N_4463,N_4390);
nor U4577 (N_4577,N_4360,N_4475);
xor U4578 (N_4578,N_4356,N_4435);
nand U4579 (N_4579,N_4471,N_4391);
or U4580 (N_4580,N_4489,N_4475);
xnor U4581 (N_4581,N_4418,N_4478);
nor U4582 (N_4582,N_4465,N_4451);
and U4583 (N_4583,N_4418,N_4400);
nor U4584 (N_4584,N_4467,N_4370);
nand U4585 (N_4585,N_4414,N_4393);
nor U4586 (N_4586,N_4395,N_4355);
or U4587 (N_4587,N_4481,N_4412);
or U4588 (N_4588,N_4381,N_4442);
xor U4589 (N_4589,N_4378,N_4358);
nand U4590 (N_4590,N_4396,N_4458);
nand U4591 (N_4591,N_4381,N_4418);
xnor U4592 (N_4592,N_4419,N_4456);
and U4593 (N_4593,N_4354,N_4390);
or U4594 (N_4594,N_4435,N_4416);
or U4595 (N_4595,N_4455,N_4392);
and U4596 (N_4596,N_4392,N_4453);
xor U4597 (N_4597,N_4452,N_4451);
xnor U4598 (N_4598,N_4370,N_4355);
or U4599 (N_4599,N_4441,N_4354);
nor U4600 (N_4600,N_4353,N_4413);
nand U4601 (N_4601,N_4430,N_4463);
nand U4602 (N_4602,N_4394,N_4389);
or U4603 (N_4603,N_4465,N_4480);
or U4604 (N_4604,N_4422,N_4467);
or U4605 (N_4605,N_4423,N_4353);
and U4606 (N_4606,N_4467,N_4475);
or U4607 (N_4607,N_4426,N_4451);
nor U4608 (N_4608,N_4351,N_4426);
nand U4609 (N_4609,N_4422,N_4445);
nand U4610 (N_4610,N_4365,N_4400);
or U4611 (N_4611,N_4435,N_4388);
nand U4612 (N_4612,N_4356,N_4440);
xor U4613 (N_4613,N_4499,N_4399);
nand U4614 (N_4614,N_4457,N_4437);
nand U4615 (N_4615,N_4398,N_4378);
and U4616 (N_4616,N_4394,N_4493);
xnor U4617 (N_4617,N_4468,N_4395);
and U4618 (N_4618,N_4451,N_4467);
nor U4619 (N_4619,N_4446,N_4438);
and U4620 (N_4620,N_4415,N_4423);
xnor U4621 (N_4621,N_4498,N_4378);
nand U4622 (N_4622,N_4398,N_4429);
xnor U4623 (N_4623,N_4472,N_4370);
xor U4624 (N_4624,N_4477,N_4379);
or U4625 (N_4625,N_4477,N_4409);
or U4626 (N_4626,N_4444,N_4461);
and U4627 (N_4627,N_4491,N_4486);
and U4628 (N_4628,N_4494,N_4387);
or U4629 (N_4629,N_4405,N_4473);
nand U4630 (N_4630,N_4387,N_4471);
or U4631 (N_4631,N_4471,N_4426);
and U4632 (N_4632,N_4410,N_4455);
and U4633 (N_4633,N_4359,N_4435);
nor U4634 (N_4634,N_4392,N_4463);
nand U4635 (N_4635,N_4367,N_4429);
xnor U4636 (N_4636,N_4395,N_4414);
or U4637 (N_4637,N_4491,N_4350);
nand U4638 (N_4638,N_4435,N_4358);
or U4639 (N_4639,N_4410,N_4432);
nor U4640 (N_4640,N_4489,N_4498);
or U4641 (N_4641,N_4376,N_4350);
nor U4642 (N_4642,N_4393,N_4484);
nor U4643 (N_4643,N_4455,N_4440);
nand U4644 (N_4644,N_4446,N_4375);
nand U4645 (N_4645,N_4451,N_4447);
and U4646 (N_4646,N_4494,N_4498);
nor U4647 (N_4647,N_4369,N_4453);
xor U4648 (N_4648,N_4447,N_4480);
and U4649 (N_4649,N_4497,N_4403);
or U4650 (N_4650,N_4525,N_4605);
nand U4651 (N_4651,N_4595,N_4563);
xor U4652 (N_4652,N_4533,N_4539);
nand U4653 (N_4653,N_4526,N_4542);
xnor U4654 (N_4654,N_4543,N_4639);
nand U4655 (N_4655,N_4597,N_4648);
or U4656 (N_4656,N_4570,N_4553);
and U4657 (N_4657,N_4540,N_4504);
nor U4658 (N_4658,N_4623,N_4562);
or U4659 (N_4659,N_4555,N_4557);
nor U4660 (N_4660,N_4637,N_4567);
and U4661 (N_4661,N_4590,N_4512);
nor U4662 (N_4662,N_4642,N_4560);
xor U4663 (N_4663,N_4524,N_4589);
nand U4664 (N_4664,N_4518,N_4582);
xor U4665 (N_4665,N_4551,N_4592);
and U4666 (N_4666,N_4596,N_4606);
nand U4667 (N_4667,N_4644,N_4600);
xnor U4668 (N_4668,N_4584,N_4618);
nor U4669 (N_4669,N_4558,N_4588);
nand U4670 (N_4670,N_4576,N_4507);
or U4671 (N_4671,N_4566,N_4635);
nand U4672 (N_4672,N_4641,N_4523);
nor U4673 (N_4673,N_4591,N_4501);
and U4674 (N_4674,N_4536,N_4556);
nand U4675 (N_4675,N_4636,N_4578);
nor U4676 (N_4676,N_4601,N_4564);
or U4677 (N_4677,N_4569,N_4506);
nor U4678 (N_4678,N_4520,N_4500);
nor U4679 (N_4679,N_4528,N_4568);
nand U4680 (N_4680,N_4634,N_4534);
nor U4681 (N_4681,N_4628,N_4538);
or U4682 (N_4682,N_4633,N_4517);
nand U4683 (N_4683,N_4544,N_4640);
xor U4684 (N_4684,N_4530,N_4647);
and U4685 (N_4685,N_4552,N_4624);
and U4686 (N_4686,N_4577,N_4535);
nand U4687 (N_4687,N_4549,N_4608);
xnor U4688 (N_4688,N_4522,N_4554);
and U4689 (N_4689,N_4529,N_4585);
nand U4690 (N_4690,N_4546,N_4643);
xnor U4691 (N_4691,N_4509,N_4631);
nand U4692 (N_4692,N_4531,N_4583);
xnor U4693 (N_4693,N_4629,N_4513);
nor U4694 (N_4694,N_4610,N_4580);
xnor U4695 (N_4695,N_4620,N_4649);
nor U4696 (N_4696,N_4511,N_4598);
nand U4697 (N_4697,N_4616,N_4622);
and U4698 (N_4698,N_4614,N_4547);
and U4699 (N_4699,N_4575,N_4645);
nor U4700 (N_4700,N_4532,N_4548);
nand U4701 (N_4701,N_4646,N_4502);
and U4702 (N_4702,N_4516,N_4574);
nor U4703 (N_4703,N_4527,N_4515);
xnor U4704 (N_4704,N_4541,N_4632);
and U4705 (N_4705,N_4612,N_4599);
and U4706 (N_4706,N_4514,N_4508);
and U4707 (N_4707,N_4561,N_4503);
nand U4708 (N_4708,N_4572,N_4587);
nand U4709 (N_4709,N_4586,N_4609);
xor U4710 (N_4710,N_4604,N_4537);
xor U4711 (N_4711,N_4565,N_4621);
or U4712 (N_4712,N_4545,N_4638);
and U4713 (N_4713,N_4603,N_4617);
nor U4714 (N_4714,N_4559,N_4510);
and U4715 (N_4715,N_4607,N_4521);
nor U4716 (N_4716,N_4594,N_4593);
nand U4717 (N_4717,N_4505,N_4550);
or U4718 (N_4718,N_4613,N_4571);
xor U4719 (N_4719,N_4625,N_4602);
xor U4720 (N_4720,N_4519,N_4627);
and U4721 (N_4721,N_4630,N_4611);
or U4722 (N_4722,N_4573,N_4579);
or U4723 (N_4723,N_4619,N_4626);
or U4724 (N_4724,N_4581,N_4615);
and U4725 (N_4725,N_4554,N_4642);
or U4726 (N_4726,N_4551,N_4587);
and U4727 (N_4727,N_4532,N_4561);
nand U4728 (N_4728,N_4531,N_4561);
nand U4729 (N_4729,N_4506,N_4566);
nand U4730 (N_4730,N_4628,N_4542);
and U4731 (N_4731,N_4606,N_4633);
xor U4732 (N_4732,N_4619,N_4560);
or U4733 (N_4733,N_4629,N_4508);
xor U4734 (N_4734,N_4600,N_4550);
or U4735 (N_4735,N_4576,N_4516);
or U4736 (N_4736,N_4561,N_4606);
nor U4737 (N_4737,N_4547,N_4536);
xnor U4738 (N_4738,N_4543,N_4576);
nor U4739 (N_4739,N_4641,N_4556);
nor U4740 (N_4740,N_4619,N_4552);
nor U4741 (N_4741,N_4516,N_4596);
nor U4742 (N_4742,N_4543,N_4646);
nand U4743 (N_4743,N_4593,N_4602);
nor U4744 (N_4744,N_4568,N_4587);
and U4745 (N_4745,N_4645,N_4576);
nor U4746 (N_4746,N_4568,N_4503);
nor U4747 (N_4747,N_4606,N_4541);
xnor U4748 (N_4748,N_4639,N_4539);
or U4749 (N_4749,N_4551,N_4531);
xnor U4750 (N_4750,N_4623,N_4508);
xor U4751 (N_4751,N_4572,N_4645);
and U4752 (N_4752,N_4514,N_4563);
and U4753 (N_4753,N_4632,N_4518);
and U4754 (N_4754,N_4505,N_4570);
nor U4755 (N_4755,N_4557,N_4609);
xnor U4756 (N_4756,N_4605,N_4595);
or U4757 (N_4757,N_4515,N_4551);
nor U4758 (N_4758,N_4625,N_4553);
xor U4759 (N_4759,N_4607,N_4567);
xor U4760 (N_4760,N_4543,N_4601);
xor U4761 (N_4761,N_4577,N_4647);
nor U4762 (N_4762,N_4534,N_4599);
nand U4763 (N_4763,N_4597,N_4589);
xnor U4764 (N_4764,N_4623,N_4585);
nand U4765 (N_4765,N_4648,N_4521);
xor U4766 (N_4766,N_4596,N_4571);
nor U4767 (N_4767,N_4590,N_4560);
or U4768 (N_4768,N_4568,N_4647);
or U4769 (N_4769,N_4646,N_4534);
and U4770 (N_4770,N_4580,N_4569);
nor U4771 (N_4771,N_4603,N_4543);
or U4772 (N_4772,N_4613,N_4531);
xnor U4773 (N_4773,N_4615,N_4638);
nor U4774 (N_4774,N_4604,N_4564);
nor U4775 (N_4775,N_4524,N_4501);
xor U4776 (N_4776,N_4543,N_4566);
and U4777 (N_4777,N_4645,N_4561);
nand U4778 (N_4778,N_4579,N_4511);
nor U4779 (N_4779,N_4553,N_4590);
xor U4780 (N_4780,N_4517,N_4649);
or U4781 (N_4781,N_4604,N_4585);
and U4782 (N_4782,N_4509,N_4645);
or U4783 (N_4783,N_4528,N_4545);
xnor U4784 (N_4784,N_4587,N_4617);
or U4785 (N_4785,N_4533,N_4541);
nand U4786 (N_4786,N_4593,N_4546);
xnor U4787 (N_4787,N_4590,N_4640);
and U4788 (N_4788,N_4622,N_4585);
nor U4789 (N_4789,N_4577,N_4571);
nor U4790 (N_4790,N_4520,N_4576);
and U4791 (N_4791,N_4592,N_4522);
nor U4792 (N_4792,N_4524,N_4527);
xor U4793 (N_4793,N_4586,N_4614);
xor U4794 (N_4794,N_4559,N_4511);
nor U4795 (N_4795,N_4587,N_4626);
nand U4796 (N_4796,N_4609,N_4633);
xor U4797 (N_4797,N_4539,N_4587);
xor U4798 (N_4798,N_4613,N_4541);
or U4799 (N_4799,N_4588,N_4581);
nand U4800 (N_4800,N_4779,N_4684);
or U4801 (N_4801,N_4758,N_4700);
and U4802 (N_4802,N_4749,N_4785);
and U4803 (N_4803,N_4663,N_4764);
and U4804 (N_4804,N_4709,N_4723);
xnor U4805 (N_4805,N_4671,N_4761);
nor U4806 (N_4806,N_4740,N_4745);
nor U4807 (N_4807,N_4790,N_4672);
xnor U4808 (N_4808,N_4772,N_4755);
and U4809 (N_4809,N_4652,N_4746);
nor U4810 (N_4810,N_4660,N_4774);
or U4811 (N_4811,N_4752,N_4795);
and U4812 (N_4812,N_4767,N_4703);
and U4813 (N_4813,N_4653,N_4670);
nand U4814 (N_4814,N_4760,N_4701);
or U4815 (N_4815,N_4694,N_4702);
or U4816 (N_4816,N_4708,N_4750);
or U4817 (N_4817,N_4783,N_4770);
and U4818 (N_4818,N_4724,N_4748);
or U4819 (N_4819,N_4654,N_4683);
or U4820 (N_4820,N_4714,N_4682);
or U4821 (N_4821,N_4679,N_4693);
nand U4822 (N_4822,N_4747,N_4674);
nand U4823 (N_4823,N_4728,N_4754);
nand U4824 (N_4824,N_4696,N_4689);
or U4825 (N_4825,N_4718,N_4778);
or U4826 (N_4826,N_4743,N_4707);
xnor U4827 (N_4827,N_4713,N_4725);
nand U4828 (N_4828,N_4662,N_4791);
or U4829 (N_4829,N_4768,N_4676);
xnor U4830 (N_4830,N_4782,N_4729);
nand U4831 (N_4831,N_4726,N_4675);
nand U4832 (N_4832,N_4688,N_4650);
and U4833 (N_4833,N_4757,N_4794);
nor U4834 (N_4834,N_4734,N_4780);
and U4835 (N_4835,N_4756,N_4658);
or U4836 (N_4836,N_4705,N_4711);
and U4837 (N_4837,N_4744,N_4776);
nor U4838 (N_4838,N_4687,N_4735);
xor U4839 (N_4839,N_4781,N_4690);
and U4840 (N_4840,N_4715,N_4680);
or U4841 (N_4841,N_4739,N_4667);
and U4842 (N_4842,N_4730,N_4775);
or U4843 (N_4843,N_4664,N_4759);
nor U4844 (N_4844,N_4685,N_4668);
nor U4845 (N_4845,N_4796,N_4769);
nand U4846 (N_4846,N_4712,N_4793);
nand U4847 (N_4847,N_4697,N_4742);
nor U4848 (N_4848,N_4771,N_4698);
and U4849 (N_4849,N_4784,N_4704);
or U4850 (N_4850,N_4717,N_4737);
and U4851 (N_4851,N_4765,N_4699);
or U4852 (N_4852,N_4741,N_4727);
and U4853 (N_4853,N_4657,N_4738);
nand U4854 (N_4854,N_4787,N_4786);
xnor U4855 (N_4855,N_4656,N_4721);
xor U4856 (N_4856,N_4692,N_4673);
nand U4857 (N_4857,N_4799,N_4731);
nor U4858 (N_4858,N_4733,N_4797);
and U4859 (N_4859,N_4677,N_4716);
nor U4860 (N_4860,N_4678,N_4695);
or U4861 (N_4861,N_4661,N_4681);
xnor U4862 (N_4862,N_4753,N_4719);
nor U4863 (N_4863,N_4691,N_4736);
and U4864 (N_4864,N_4651,N_4666);
or U4865 (N_4865,N_4792,N_4669);
xor U4866 (N_4866,N_4665,N_4789);
xnor U4867 (N_4867,N_4655,N_4720);
xnor U4868 (N_4868,N_4763,N_4766);
xnor U4869 (N_4869,N_4686,N_4722);
and U4870 (N_4870,N_4777,N_4751);
and U4871 (N_4871,N_4788,N_4762);
xnor U4872 (N_4872,N_4798,N_4659);
xor U4873 (N_4873,N_4710,N_4773);
nor U4874 (N_4874,N_4706,N_4732);
nand U4875 (N_4875,N_4737,N_4684);
xnor U4876 (N_4876,N_4758,N_4792);
nand U4877 (N_4877,N_4704,N_4799);
nor U4878 (N_4878,N_4704,N_4765);
nor U4879 (N_4879,N_4756,N_4740);
or U4880 (N_4880,N_4659,N_4666);
and U4881 (N_4881,N_4752,N_4745);
xor U4882 (N_4882,N_4708,N_4713);
or U4883 (N_4883,N_4735,N_4713);
xnor U4884 (N_4884,N_4718,N_4771);
xor U4885 (N_4885,N_4722,N_4731);
or U4886 (N_4886,N_4688,N_4783);
and U4887 (N_4887,N_4658,N_4752);
and U4888 (N_4888,N_4667,N_4704);
nand U4889 (N_4889,N_4662,N_4713);
xnor U4890 (N_4890,N_4672,N_4690);
and U4891 (N_4891,N_4739,N_4758);
or U4892 (N_4892,N_4673,N_4738);
nor U4893 (N_4893,N_4792,N_4683);
nor U4894 (N_4894,N_4736,N_4734);
and U4895 (N_4895,N_4743,N_4731);
nand U4896 (N_4896,N_4713,N_4758);
and U4897 (N_4897,N_4766,N_4710);
xor U4898 (N_4898,N_4731,N_4652);
xnor U4899 (N_4899,N_4653,N_4721);
nand U4900 (N_4900,N_4779,N_4711);
and U4901 (N_4901,N_4775,N_4739);
or U4902 (N_4902,N_4751,N_4723);
xnor U4903 (N_4903,N_4733,N_4781);
nor U4904 (N_4904,N_4745,N_4734);
xnor U4905 (N_4905,N_4654,N_4738);
xnor U4906 (N_4906,N_4753,N_4667);
nor U4907 (N_4907,N_4748,N_4760);
nor U4908 (N_4908,N_4655,N_4651);
nor U4909 (N_4909,N_4698,N_4719);
nor U4910 (N_4910,N_4680,N_4693);
or U4911 (N_4911,N_4735,N_4797);
xnor U4912 (N_4912,N_4775,N_4759);
nand U4913 (N_4913,N_4673,N_4693);
or U4914 (N_4914,N_4748,N_4753);
nor U4915 (N_4915,N_4700,N_4747);
nand U4916 (N_4916,N_4799,N_4785);
nor U4917 (N_4917,N_4792,N_4662);
nor U4918 (N_4918,N_4743,N_4792);
nand U4919 (N_4919,N_4692,N_4782);
nand U4920 (N_4920,N_4717,N_4725);
nor U4921 (N_4921,N_4728,N_4715);
xor U4922 (N_4922,N_4661,N_4777);
xor U4923 (N_4923,N_4677,N_4749);
or U4924 (N_4924,N_4776,N_4787);
xor U4925 (N_4925,N_4683,N_4782);
xnor U4926 (N_4926,N_4720,N_4753);
and U4927 (N_4927,N_4717,N_4799);
xnor U4928 (N_4928,N_4660,N_4748);
nand U4929 (N_4929,N_4672,N_4698);
nand U4930 (N_4930,N_4687,N_4710);
xor U4931 (N_4931,N_4798,N_4684);
nor U4932 (N_4932,N_4741,N_4771);
nand U4933 (N_4933,N_4650,N_4791);
nand U4934 (N_4934,N_4726,N_4661);
or U4935 (N_4935,N_4684,N_4751);
nand U4936 (N_4936,N_4673,N_4793);
nand U4937 (N_4937,N_4798,N_4687);
nand U4938 (N_4938,N_4689,N_4687);
nor U4939 (N_4939,N_4654,N_4741);
nand U4940 (N_4940,N_4716,N_4773);
nor U4941 (N_4941,N_4682,N_4752);
nand U4942 (N_4942,N_4798,N_4772);
xnor U4943 (N_4943,N_4749,N_4652);
nor U4944 (N_4944,N_4724,N_4655);
and U4945 (N_4945,N_4771,N_4790);
nand U4946 (N_4946,N_4728,N_4654);
nor U4947 (N_4947,N_4668,N_4701);
xnor U4948 (N_4948,N_4764,N_4799);
xor U4949 (N_4949,N_4793,N_4740);
xor U4950 (N_4950,N_4889,N_4885);
or U4951 (N_4951,N_4827,N_4925);
or U4952 (N_4952,N_4820,N_4874);
nand U4953 (N_4953,N_4895,N_4880);
or U4954 (N_4954,N_4816,N_4801);
nor U4955 (N_4955,N_4902,N_4881);
and U4956 (N_4956,N_4910,N_4924);
and U4957 (N_4957,N_4920,N_4863);
and U4958 (N_4958,N_4918,N_4821);
nor U4959 (N_4959,N_4855,N_4848);
nor U4960 (N_4960,N_4931,N_4804);
and U4961 (N_4961,N_4892,N_4847);
or U4962 (N_4962,N_4861,N_4948);
xor U4963 (N_4963,N_4834,N_4823);
or U4964 (N_4964,N_4870,N_4846);
nand U4965 (N_4965,N_4935,N_4900);
nor U4966 (N_4966,N_4916,N_4914);
xor U4967 (N_4967,N_4907,N_4901);
or U4968 (N_4968,N_4840,N_4852);
xor U4969 (N_4969,N_4825,N_4937);
nand U4970 (N_4970,N_4854,N_4831);
or U4971 (N_4971,N_4845,N_4807);
nor U4972 (N_4972,N_4946,N_4815);
nand U4973 (N_4973,N_4832,N_4802);
nand U4974 (N_4974,N_4873,N_4819);
nand U4975 (N_4975,N_4877,N_4883);
or U4976 (N_4976,N_4886,N_4933);
and U4977 (N_4977,N_4806,N_4926);
xnor U4978 (N_4978,N_4865,N_4919);
or U4979 (N_4979,N_4894,N_4884);
nand U4980 (N_4980,N_4800,N_4811);
nand U4981 (N_4981,N_4842,N_4936);
xor U4982 (N_4982,N_4882,N_4913);
nand U4983 (N_4983,N_4837,N_4909);
nor U4984 (N_4984,N_4803,N_4839);
and U4985 (N_4985,N_4938,N_4888);
or U4986 (N_4986,N_4878,N_4887);
xnor U4987 (N_4987,N_4947,N_4923);
xor U4988 (N_4988,N_4856,N_4922);
or U4989 (N_4989,N_4844,N_4808);
nor U4990 (N_4990,N_4945,N_4896);
and U4991 (N_4991,N_4859,N_4934);
nand U4992 (N_4992,N_4812,N_4876);
xnor U4993 (N_4993,N_4862,N_4904);
or U4994 (N_4994,N_4908,N_4829);
nand U4995 (N_4995,N_4891,N_4813);
nor U4996 (N_4996,N_4941,N_4814);
nand U4997 (N_4997,N_4869,N_4949);
or U4998 (N_4998,N_4860,N_4868);
and U4999 (N_4999,N_4940,N_4875);
xnor U5000 (N_5000,N_4850,N_4898);
and U5001 (N_5001,N_4838,N_4932);
nand U5002 (N_5002,N_4912,N_4805);
nand U5003 (N_5003,N_4944,N_4939);
and U5004 (N_5004,N_4917,N_4897);
and U5005 (N_5005,N_4835,N_4942);
nor U5006 (N_5006,N_4929,N_4903);
and U5007 (N_5007,N_4871,N_4864);
and U5008 (N_5008,N_4867,N_4810);
or U5009 (N_5009,N_4826,N_4858);
and U5010 (N_5010,N_4824,N_4943);
xnor U5011 (N_5011,N_4872,N_4849);
and U5012 (N_5012,N_4893,N_4830);
nand U5013 (N_5013,N_4851,N_4921);
and U5014 (N_5014,N_4853,N_4833);
nand U5015 (N_5015,N_4927,N_4906);
xnor U5016 (N_5016,N_4809,N_4841);
nor U5017 (N_5017,N_4866,N_4899);
xnor U5018 (N_5018,N_4836,N_4911);
or U5019 (N_5019,N_4828,N_4822);
nand U5020 (N_5020,N_4857,N_4905);
and U5021 (N_5021,N_4843,N_4915);
nand U5022 (N_5022,N_4817,N_4879);
or U5023 (N_5023,N_4928,N_4890);
nor U5024 (N_5024,N_4930,N_4818);
nand U5025 (N_5025,N_4817,N_4839);
nor U5026 (N_5026,N_4808,N_4801);
and U5027 (N_5027,N_4819,N_4860);
and U5028 (N_5028,N_4892,N_4858);
nor U5029 (N_5029,N_4856,N_4928);
xnor U5030 (N_5030,N_4934,N_4905);
xor U5031 (N_5031,N_4933,N_4836);
xnor U5032 (N_5032,N_4937,N_4860);
xnor U5033 (N_5033,N_4855,N_4849);
and U5034 (N_5034,N_4935,N_4916);
or U5035 (N_5035,N_4833,N_4854);
nand U5036 (N_5036,N_4938,N_4947);
or U5037 (N_5037,N_4919,N_4929);
or U5038 (N_5038,N_4820,N_4928);
and U5039 (N_5039,N_4876,N_4938);
or U5040 (N_5040,N_4889,N_4918);
xnor U5041 (N_5041,N_4811,N_4931);
xnor U5042 (N_5042,N_4867,N_4856);
nand U5043 (N_5043,N_4912,N_4896);
and U5044 (N_5044,N_4881,N_4839);
nand U5045 (N_5045,N_4840,N_4896);
xnor U5046 (N_5046,N_4921,N_4932);
nand U5047 (N_5047,N_4939,N_4933);
nand U5048 (N_5048,N_4871,N_4806);
nand U5049 (N_5049,N_4947,N_4897);
nand U5050 (N_5050,N_4825,N_4938);
and U5051 (N_5051,N_4849,N_4911);
xnor U5052 (N_5052,N_4820,N_4810);
nand U5053 (N_5053,N_4905,N_4861);
or U5054 (N_5054,N_4835,N_4920);
nor U5055 (N_5055,N_4846,N_4859);
nor U5056 (N_5056,N_4893,N_4848);
xnor U5057 (N_5057,N_4879,N_4823);
and U5058 (N_5058,N_4804,N_4827);
xor U5059 (N_5059,N_4861,N_4940);
nand U5060 (N_5060,N_4832,N_4929);
or U5061 (N_5061,N_4947,N_4889);
nor U5062 (N_5062,N_4844,N_4944);
nand U5063 (N_5063,N_4889,N_4811);
and U5064 (N_5064,N_4821,N_4807);
and U5065 (N_5065,N_4869,N_4913);
nor U5066 (N_5066,N_4855,N_4874);
nand U5067 (N_5067,N_4905,N_4911);
and U5068 (N_5068,N_4849,N_4803);
nand U5069 (N_5069,N_4897,N_4920);
nor U5070 (N_5070,N_4917,N_4859);
nor U5071 (N_5071,N_4940,N_4914);
xor U5072 (N_5072,N_4936,N_4876);
or U5073 (N_5073,N_4804,N_4810);
or U5074 (N_5074,N_4859,N_4834);
and U5075 (N_5075,N_4829,N_4883);
nor U5076 (N_5076,N_4890,N_4813);
or U5077 (N_5077,N_4831,N_4840);
and U5078 (N_5078,N_4911,N_4933);
nand U5079 (N_5079,N_4836,N_4847);
nand U5080 (N_5080,N_4863,N_4875);
or U5081 (N_5081,N_4885,N_4901);
nand U5082 (N_5082,N_4835,N_4863);
xnor U5083 (N_5083,N_4837,N_4844);
or U5084 (N_5084,N_4844,N_4857);
and U5085 (N_5085,N_4895,N_4831);
or U5086 (N_5086,N_4924,N_4876);
and U5087 (N_5087,N_4943,N_4935);
xor U5088 (N_5088,N_4901,N_4912);
or U5089 (N_5089,N_4808,N_4861);
nand U5090 (N_5090,N_4912,N_4856);
and U5091 (N_5091,N_4807,N_4802);
or U5092 (N_5092,N_4803,N_4907);
xnor U5093 (N_5093,N_4859,N_4883);
nor U5094 (N_5094,N_4819,N_4826);
xor U5095 (N_5095,N_4862,N_4811);
xor U5096 (N_5096,N_4832,N_4923);
or U5097 (N_5097,N_4831,N_4878);
and U5098 (N_5098,N_4844,N_4937);
nor U5099 (N_5099,N_4838,N_4924);
or U5100 (N_5100,N_5054,N_5005);
or U5101 (N_5101,N_4981,N_5004);
nor U5102 (N_5102,N_5058,N_4983);
nand U5103 (N_5103,N_5019,N_4955);
nor U5104 (N_5104,N_5070,N_5088);
nand U5105 (N_5105,N_4996,N_5085);
or U5106 (N_5106,N_5090,N_5065);
nand U5107 (N_5107,N_5044,N_5018);
nor U5108 (N_5108,N_5040,N_5022);
or U5109 (N_5109,N_5008,N_4979);
nor U5110 (N_5110,N_5092,N_4958);
nand U5111 (N_5111,N_5093,N_5036);
or U5112 (N_5112,N_5015,N_5042);
nor U5113 (N_5113,N_5049,N_5079);
nor U5114 (N_5114,N_4952,N_4957);
nand U5115 (N_5115,N_4972,N_5026);
or U5116 (N_5116,N_5097,N_5076);
and U5117 (N_5117,N_4987,N_5045);
nand U5118 (N_5118,N_4961,N_5075);
nand U5119 (N_5119,N_5078,N_5053);
nor U5120 (N_5120,N_5051,N_4967);
nor U5121 (N_5121,N_5064,N_5002);
and U5122 (N_5122,N_4960,N_5094);
nor U5123 (N_5123,N_4950,N_5037);
nor U5124 (N_5124,N_5077,N_4982);
nor U5125 (N_5125,N_5060,N_4994);
and U5126 (N_5126,N_5021,N_4985);
or U5127 (N_5127,N_5010,N_4992);
nor U5128 (N_5128,N_4963,N_4968);
or U5129 (N_5129,N_4977,N_5095);
xor U5130 (N_5130,N_5028,N_5096);
nand U5131 (N_5131,N_5011,N_5001);
xnor U5132 (N_5132,N_5043,N_5067);
nand U5133 (N_5133,N_4971,N_5048);
or U5134 (N_5134,N_5057,N_4997);
nor U5135 (N_5135,N_5023,N_5069);
xnor U5136 (N_5136,N_5027,N_5081);
or U5137 (N_5137,N_5087,N_5080);
or U5138 (N_5138,N_4973,N_5072);
xor U5139 (N_5139,N_4959,N_5038);
nand U5140 (N_5140,N_4976,N_4953);
nand U5141 (N_5141,N_5091,N_5071);
or U5142 (N_5142,N_5089,N_5062);
nor U5143 (N_5143,N_4988,N_4995);
or U5144 (N_5144,N_4978,N_5052);
or U5145 (N_5145,N_5034,N_4964);
nand U5146 (N_5146,N_5000,N_4991);
xnor U5147 (N_5147,N_5033,N_5063);
nand U5148 (N_5148,N_5017,N_5068);
nor U5149 (N_5149,N_4984,N_4974);
or U5150 (N_5150,N_4986,N_5032);
and U5151 (N_5151,N_4962,N_5029);
nand U5152 (N_5152,N_4954,N_5083);
and U5153 (N_5153,N_5086,N_5016);
nor U5154 (N_5154,N_5014,N_4980);
xnor U5155 (N_5155,N_5056,N_5039);
xnor U5156 (N_5156,N_5013,N_4965);
and U5157 (N_5157,N_5055,N_5006);
xor U5158 (N_5158,N_5003,N_5050);
xor U5159 (N_5159,N_5084,N_5024);
and U5160 (N_5160,N_5082,N_5025);
and U5161 (N_5161,N_5009,N_5066);
or U5162 (N_5162,N_4966,N_4993);
or U5163 (N_5163,N_5030,N_4990);
nor U5164 (N_5164,N_5031,N_5035);
or U5165 (N_5165,N_4970,N_5099);
or U5166 (N_5166,N_5020,N_5012);
xnor U5167 (N_5167,N_4956,N_4989);
or U5168 (N_5168,N_5098,N_5007);
and U5169 (N_5169,N_5061,N_4999);
and U5170 (N_5170,N_4998,N_5074);
or U5171 (N_5171,N_5041,N_5047);
nand U5172 (N_5172,N_4951,N_5046);
nor U5173 (N_5173,N_5059,N_4969);
or U5174 (N_5174,N_4975,N_5073);
nand U5175 (N_5175,N_5066,N_5015);
nand U5176 (N_5176,N_5087,N_5054);
xnor U5177 (N_5177,N_5006,N_5020);
and U5178 (N_5178,N_5079,N_4960);
nor U5179 (N_5179,N_5042,N_5053);
and U5180 (N_5180,N_5071,N_5024);
nor U5181 (N_5181,N_5016,N_4952);
or U5182 (N_5182,N_4983,N_5064);
xor U5183 (N_5183,N_4991,N_4971);
nor U5184 (N_5184,N_5089,N_4954);
nand U5185 (N_5185,N_5049,N_5073);
nand U5186 (N_5186,N_5095,N_5027);
and U5187 (N_5187,N_4955,N_4960);
nor U5188 (N_5188,N_5029,N_5004);
xnor U5189 (N_5189,N_4983,N_5023);
nor U5190 (N_5190,N_5010,N_5044);
xnor U5191 (N_5191,N_5026,N_4950);
xor U5192 (N_5192,N_5020,N_5082);
nand U5193 (N_5193,N_4953,N_4962);
nor U5194 (N_5194,N_5005,N_4981);
or U5195 (N_5195,N_5026,N_4998);
and U5196 (N_5196,N_5072,N_5075);
and U5197 (N_5197,N_5024,N_4959);
and U5198 (N_5198,N_4993,N_5018);
or U5199 (N_5199,N_4995,N_5013);
or U5200 (N_5200,N_5076,N_5067);
nand U5201 (N_5201,N_4997,N_5085);
and U5202 (N_5202,N_5078,N_4998);
xnor U5203 (N_5203,N_5035,N_5081);
xnor U5204 (N_5204,N_5070,N_4969);
nor U5205 (N_5205,N_4965,N_4993);
or U5206 (N_5206,N_5050,N_5082);
xor U5207 (N_5207,N_5031,N_5054);
nand U5208 (N_5208,N_5082,N_5058);
and U5209 (N_5209,N_4975,N_4974);
or U5210 (N_5210,N_5044,N_4998);
and U5211 (N_5211,N_4999,N_5068);
and U5212 (N_5212,N_5084,N_5077);
and U5213 (N_5213,N_4970,N_5045);
and U5214 (N_5214,N_5027,N_4983);
nor U5215 (N_5215,N_5048,N_4976);
nor U5216 (N_5216,N_4974,N_5052);
nand U5217 (N_5217,N_5086,N_4989);
nand U5218 (N_5218,N_5085,N_5028);
nor U5219 (N_5219,N_5031,N_4981);
xor U5220 (N_5220,N_5000,N_5084);
nand U5221 (N_5221,N_5026,N_4974);
nand U5222 (N_5222,N_4981,N_5078);
nand U5223 (N_5223,N_4985,N_5059);
and U5224 (N_5224,N_5025,N_4960);
nand U5225 (N_5225,N_5012,N_5096);
and U5226 (N_5226,N_5012,N_5071);
nand U5227 (N_5227,N_5052,N_5059);
or U5228 (N_5228,N_4982,N_5000);
xor U5229 (N_5229,N_5041,N_4977);
nor U5230 (N_5230,N_5053,N_5070);
and U5231 (N_5231,N_5034,N_5043);
nand U5232 (N_5232,N_4984,N_5083);
nand U5233 (N_5233,N_5017,N_5013);
xnor U5234 (N_5234,N_5058,N_4970);
or U5235 (N_5235,N_5081,N_4972);
nand U5236 (N_5236,N_5048,N_5010);
nor U5237 (N_5237,N_5071,N_5030);
and U5238 (N_5238,N_5027,N_5018);
nor U5239 (N_5239,N_4990,N_5093);
nor U5240 (N_5240,N_5098,N_4951);
or U5241 (N_5241,N_5080,N_4988);
and U5242 (N_5242,N_5061,N_5050);
nor U5243 (N_5243,N_5012,N_5057);
nand U5244 (N_5244,N_5046,N_5037);
and U5245 (N_5245,N_5001,N_4974);
or U5246 (N_5246,N_5003,N_5055);
xnor U5247 (N_5247,N_5004,N_5067);
xor U5248 (N_5248,N_5053,N_5033);
xor U5249 (N_5249,N_4999,N_5047);
xor U5250 (N_5250,N_5246,N_5144);
and U5251 (N_5251,N_5113,N_5114);
or U5252 (N_5252,N_5170,N_5131);
nand U5253 (N_5253,N_5228,N_5128);
xor U5254 (N_5254,N_5165,N_5150);
and U5255 (N_5255,N_5211,N_5105);
and U5256 (N_5256,N_5248,N_5197);
or U5257 (N_5257,N_5196,N_5109);
or U5258 (N_5258,N_5188,N_5205);
or U5259 (N_5259,N_5193,N_5181);
xnor U5260 (N_5260,N_5224,N_5146);
nor U5261 (N_5261,N_5120,N_5244);
or U5262 (N_5262,N_5198,N_5187);
xnor U5263 (N_5263,N_5191,N_5243);
nand U5264 (N_5264,N_5200,N_5174);
nor U5265 (N_5265,N_5151,N_5241);
and U5266 (N_5266,N_5119,N_5117);
xnor U5267 (N_5267,N_5210,N_5185);
xnor U5268 (N_5268,N_5129,N_5125);
and U5269 (N_5269,N_5158,N_5132);
nor U5270 (N_5270,N_5160,N_5111);
nand U5271 (N_5271,N_5177,N_5141);
or U5272 (N_5272,N_5122,N_5207);
nor U5273 (N_5273,N_5218,N_5137);
nor U5274 (N_5274,N_5178,N_5123);
or U5275 (N_5275,N_5219,N_5232);
and U5276 (N_5276,N_5199,N_5172);
or U5277 (N_5277,N_5209,N_5226);
xor U5278 (N_5278,N_5216,N_5135);
nor U5279 (N_5279,N_5201,N_5153);
or U5280 (N_5280,N_5190,N_5202);
or U5281 (N_5281,N_5204,N_5149);
xnor U5282 (N_5282,N_5104,N_5222);
or U5283 (N_5283,N_5145,N_5169);
and U5284 (N_5284,N_5133,N_5139);
and U5285 (N_5285,N_5107,N_5136);
nand U5286 (N_5286,N_5183,N_5116);
xor U5287 (N_5287,N_5237,N_5213);
or U5288 (N_5288,N_5159,N_5245);
nor U5289 (N_5289,N_5240,N_5176);
and U5290 (N_5290,N_5194,N_5155);
or U5291 (N_5291,N_5152,N_5127);
nand U5292 (N_5292,N_5164,N_5242);
or U5293 (N_5293,N_5108,N_5156);
nor U5294 (N_5294,N_5195,N_5247);
nor U5295 (N_5295,N_5163,N_5189);
xor U5296 (N_5296,N_5225,N_5212);
xnor U5297 (N_5297,N_5184,N_5220);
nor U5298 (N_5298,N_5115,N_5234);
and U5299 (N_5299,N_5121,N_5171);
and U5300 (N_5300,N_5186,N_5233);
and U5301 (N_5301,N_5236,N_5173);
and U5302 (N_5302,N_5106,N_5167);
xor U5303 (N_5303,N_5126,N_5168);
xnor U5304 (N_5304,N_5142,N_5147);
nand U5305 (N_5305,N_5217,N_5206);
xor U5306 (N_5306,N_5124,N_5249);
or U5307 (N_5307,N_5235,N_5179);
or U5308 (N_5308,N_5143,N_5134);
nand U5309 (N_5309,N_5182,N_5100);
or U5310 (N_5310,N_5154,N_5215);
nand U5311 (N_5311,N_5230,N_5118);
xor U5312 (N_5312,N_5166,N_5180);
nor U5313 (N_5313,N_5162,N_5238);
or U5314 (N_5314,N_5231,N_5101);
xnor U5315 (N_5315,N_5161,N_5157);
and U5316 (N_5316,N_5203,N_5208);
and U5317 (N_5317,N_5239,N_5112);
xnor U5318 (N_5318,N_5227,N_5110);
nand U5319 (N_5319,N_5103,N_5214);
xnor U5320 (N_5320,N_5140,N_5192);
nor U5321 (N_5321,N_5175,N_5138);
nand U5322 (N_5322,N_5223,N_5148);
nor U5323 (N_5323,N_5221,N_5102);
xor U5324 (N_5324,N_5229,N_5130);
nand U5325 (N_5325,N_5132,N_5209);
nand U5326 (N_5326,N_5135,N_5241);
xor U5327 (N_5327,N_5123,N_5170);
and U5328 (N_5328,N_5191,N_5227);
or U5329 (N_5329,N_5225,N_5236);
or U5330 (N_5330,N_5187,N_5176);
nand U5331 (N_5331,N_5240,N_5154);
xnor U5332 (N_5332,N_5204,N_5183);
nand U5333 (N_5333,N_5204,N_5115);
xnor U5334 (N_5334,N_5121,N_5144);
and U5335 (N_5335,N_5110,N_5117);
nand U5336 (N_5336,N_5227,N_5120);
or U5337 (N_5337,N_5142,N_5161);
xnor U5338 (N_5338,N_5207,N_5107);
and U5339 (N_5339,N_5136,N_5213);
and U5340 (N_5340,N_5186,N_5182);
nand U5341 (N_5341,N_5208,N_5122);
xnor U5342 (N_5342,N_5167,N_5228);
nand U5343 (N_5343,N_5162,N_5165);
nand U5344 (N_5344,N_5229,N_5140);
or U5345 (N_5345,N_5213,N_5186);
and U5346 (N_5346,N_5135,N_5233);
nand U5347 (N_5347,N_5178,N_5137);
or U5348 (N_5348,N_5247,N_5212);
and U5349 (N_5349,N_5197,N_5163);
nor U5350 (N_5350,N_5228,N_5180);
nor U5351 (N_5351,N_5138,N_5171);
xnor U5352 (N_5352,N_5233,N_5168);
and U5353 (N_5353,N_5165,N_5202);
and U5354 (N_5354,N_5172,N_5216);
nand U5355 (N_5355,N_5110,N_5219);
and U5356 (N_5356,N_5149,N_5213);
or U5357 (N_5357,N_5130,N_5227);
and U5358 (N_5358,N_5243,N_5133);
xor U5359 (N_5359,N_5185,N_5139);
or U5360 (N_5360,N_5120,N_5121);
and U5361 (N_5361,N_5105,N_5209);
xor U5362 (N_5362,N_5240,N_5145);
nand U5363 (N_5363,N_5143,N_5206);
or U5364 (N_5364,N_5170,N_5177);
xor U5365 (N_5365,N_5169,N_5200);
or U5366 (N_5366,N_5238,N_5178);
nor U5367 (N_5367,N_5159,N_5201);
and U5368 (N_5368,N_5202,N_5137);
nor U5369 (N_5369,N_5132,N_5218);
xor U5370 (N_5370,N_5128,N_5216);
nand U5371 (N_5371,N_5113,N_5206);
or U5372 (N_5372,N_5222,N_5113);
or U5373 (N_5373,N_5118,N_5102);
and U5374 (N_5374,N_5160,N_5166);
nand U5375 (N_5375,N_5187,N_5119);
nand U5376 (N_5376,N_5150,N_5249);
and U5377 (N_5377,N_5167,N_5160);
nand U5378 (N_5378,N_5238,N_5102);
xor U5379 (N_5379,N_5159,N_5202);
or U5380 (N_5380,N_5233,N_5211);
xor U5381 (N_5381,N_5229,N_5219);
xnor U5382 (N_5382,N_5100,N_5208);
and U5383 (N_5383,N_5158,N_5108);
xnor U5384 (N_5384,N_5177,N_5171);
and U5385 (N_5385,N_5138,N_5186);
and U5386 (N_5386,N_5226,N_5223);
or U5387 (N_5387,N_5218,N_5158);
xnor U5388 (N_5388,N_5188,N_5212);
or U5389 (N_5389,N_5121,N_5161);
or U5390 (N_5390,N_5159,N_5144);
nor U5391 (N_5391,N_5196,N_5198);
and U5392 (N_5392,N_5181,N_5168);
nand U5393 (N_5393,N_5249,N_5173);
nor U5394 (N_5394,N_5185,N_5110);
or U5395 (N_5395,N_5153,N_5181);
nor U5396 (N_5396,N_5209,N_5221);
nor U5397 (N_5397,N_5208,N_5127);
or U5398 (N_5398,N_5243,N_5195);
nand U5399 (N_5399,N_5150,N_5207);
xnor U5400 (N_5400,N_5313,N_5379);
nor U5401 (N_5401,N_5268,N_5325);
nor U5402 (N_5402,N_5384,N_5376);
xnor U5403 (N_5403,N_5284,N_5367);
nor U5404 (N_5404,N_5345,N_5368);
nand U5405 (N_5405,N_5389,N_5337);
nand U5406 (N_5406,N_5286,N_5288);
and U5407 (N_5407,N_5298,N_5255);
nor U5408 (N_5408,N_5358,N_5270);
or U5409 (N_5409,N_5381,N_5302);
nand U5410 (N_5410,N_5252,N_5387);
nor U5411 (N_5411,N_5280,N_5394);
nor U5412 (N_5412,N_5362,N_5330);
nor U5413 (N_5413,N_5261,N_5262);
or U5414 (N_5414,N_5277,N_5392);
and U5415 (N_5415,N_5361,N_5304);
nand U5416 (N_5416,N_5316,N_5321);
and U5417 (N_5417,N_5258,N_5357);
xor U5418 (N_5418,N_5253,N_5297);
nor U5419 (N_5419,N_5354,N_5353);
and U5420 (N_5420,N_5303,N_5349);
nand U5421 (N_5421,N_5256,N_5269);
xor U5422 (N_5422,N_5274,N_5343);
or U5423 (N_5423,N_5254,N_5364);
nand U5424 (N_5424,N_5374,N_5378);
xnor U5425 (N_5425,N_5275,N_5356);
nand U5426 (N_5426,N_5293,N_5309);
and U5427 (N_5427,N_5299,N_5292);
nand U5428 (N_5428,N_5273,N_5315);
or U5429 (N_5429,N_5319,N_5264);
nand U5430 (N_5430,N_5370,N_5366);
nand U5431 (N_5431,N_5329,N_5398);
nand U5432 (N_5432,N_5373,N_5263);
nand U5433 (N_5433,N_5351,N_5352);
and U5434 (N_5434,N_5311,N_5265);
or U5435 (N_5435,N_5342,N_5295);
or U5436 (N_5436,N_5271,N_5338);
xnor U5437 (N_5437,N_5346,N_5344);
nand U5438 (N_5438,N_5322,N_5396);
nand U5439 (N_5439,N_5386,N_5257);
xor U5440 (N_5440,N_5347,N_5290);
xor U5441 (N_5441,N_5375,N_5296);
and U5442 (N_5442,N_5336,N_5266);
or U5443 (N_5443,N_5323,N_5380);
and U5444 (N_5444,N_5300,N_5377);
and U5445 (N_5445,N_5260,N_5339);
nor U5446 (N_5446,N_5272,N_5388);
xnor U5447 (N_5447,N_5365,N_5278);
or U5448 (N_5448,N_5301,N_5251);
or U5449 (N_5449,N_5331,N_5283);
or U5450 (N_5450,N_5308,N_5391);
nand U5451 (N_5451,N_5267,N_5332);
nand U5452 (N_5452,N_5397,N_5276);
or U5453 (N_5453,N_5385,N_5399);
and U5454 (N_5454,N_5318,N_5390);
xnor U5455 (N_5455,N_5305,N_5372);
and U5456 (N_5456,N_5289,N_5334);
and U5457 (N_5457,N_5371,N_5317);
or U5458 (N_5458,N_5326,N_5355);
nand U5459 (N_5459,N_5340,N_5310);
nand U5460 (N_5460,N_5333,N_5327);
or U5461 (N_5461,N_5348,N_5324);
or U5462 (N_5462,N_5393,N_5282);
nand U5463 (N_5463,N_5341,N_5285);
nor U5464 (N_5464,N_5350,N_5312);
xor U5465 (N_5465,N_5281,N_5291);
xnor U5466 (N_5466,N_5383,N_5382);
or U5467 (N_5467,N_5369,N_5395);
and U5468 (N_5468,N_5363,N_5306);
and U5469 (N_5469,N_5359,N_5314);
nor U5470 (N_5470,N_5307,N_5294);
nor U5471 (N_5471,N_5328,N_5320);
nand U5472 (N_5472,N_5250,N_5360);
xnor U5473 (N_5473,N_5287,N_5279);
or U5474 (N_5474,N_5335,N_5259);
and U5475 (N_5475,N_5299,N_5337);
nor U5476 (N_5476,N_5263,N_5358);
nor U5477 (N_5477,N_5348,N_5384);
xnor U5478 (N_5478,N_5374,N_5345);
nor U5479 (N_5479,N_5271,N_5368);
xnor U5480 (N_5480,N_5314,N_5353);
and U5481 (N_5481,N_5268,N_5254);
and U5482 (N_5482,N_5375,N_5374);
and U5483 (N_5483,N_5341,N_5283);
or U5484 (N_5484,N_5362,N_5384);
xnor U5485 (N_5485,N_5281,N_5377);
or U5486 (N_5486,N_5365,N_5289);
or U5487 (N_5487,N_5345,N_5399);
nor U5488 (N_5488,N_5260,N_5381);
and U5489 (N_5489,N_5386,N_5344);
nand U5490 (N_5490,N_5379,N_5299);
and U5491 (N_5491,N_5360,N_5301);
and U5492 (N_5492,N_5368,N_5376);
or U5493 (N_5493,N_5315,N_5373);
and U5494 (N_5494,N_5289,N_5383);
xnor U5495 (N_5495,N_5252,N_5371);
and U5496 (N_5496,N_5356,N_5313);
xor U5497 (N_5497,N_5373,N_5377);
xnor U5498 (N_5498,N_5280,N_5355);
nand U5499 (N_5499,N_5364,N_5252);
and U5500 (N_5500,N_5346,N_5332);
nor U5501 (N_5501,N_5275,N_5287);
xnor U5502 (N_5502,N_5357,N_5371);
nand U5503 (N_5503,N_5314,N_5266);
nand U5504 (N_5504,N_5371,N_5397);
or U5505 (N_5505,N_5276,N_5343);
nand U5506 (N_5506,N_5311,N_5261);
xnor U5507 (N_5507,N_5399,N_5312);
or U5508 (N_5508,N_5294,N_5308);
and U5509 (N_5509,N_5262,N_5327);
xor U5510 (N_5510,N_5290,N_5375);
or U5511 (N_5511,N_5380,N_5383);
or U5512 (N_5512,N_5315,N_5356);
and U5513 (N_5513,N_5336,N_5257);
and U5514 (N_5514,N_5335,N_5350);
nor U5515 (N_5515,N_5386,N_5280);
xor U5516 (N_5516,N_5277,N_5365);
nand U5517 (N_5517,N_5353,N_5278);
or U5518 (N_5518,N_5339,N_5270);
or U5519 (N_5519,N_5260,N_5372);
nand U5520 (N_5520,N_5341,N_5370);
xor U5521 (N_5521,N_5314,N_5332);
and U5522 (N_5522,N_5304,N_5350);
xor U5523 (N_5523,N_5349,N_5389);
or U5524 (N_5524,N_5391,N_5390);
and U5525 (N_5525,N_5324,N_5331);
or U5526 (N_5526,N_5287,N_5384);
nor U5527 (N_5527,N_5267,N_5349);
nand U5528 (N_5528,N_5330,N_5321);
and U5529 (N_5529,N_5266,N_5329);
nor U5530 (N_5530,N_5361,N_5300);
nand U5531 (N_5531,N_5261,N_5253);
and U5532 (N_5532,N_5374,N_5273);
nor U5533 (N_5533,N_5330,N_5315);
nand U5534 (N_5534,N_5259,N_5312);
nand U5535 (N_5535,N_5258,N_5365);
nor U5536 (N_5536,N_5385,N_5299);
nand U5537 (N_5537,N_5336,N_5367);
nand U5538 (N_5538,N_5295,N_5326);
xor U5539 (N_5539,N_5347,N_5279);
xor U5540 (N_5540,N_5388,N_5302);
nand U5541 (N_5541,N_5398,N_5311);
nor U5542 (N_5542,N_5356,N_5293);
xor U5543 (N_5543,N_5383,N_5322);
and U5544 (N_5544,N_5328,N_5284);
or U5545 (N_5545,N_5252,N_5316);
nand U5546 (N_5546,N_5399,N_5383);
nand U5547 (N_5547,N_5354,N_5317);
xor U5548 (N_5548,N_5304,N_5385);
xnor U5549 (N_5549,N_5352,N_5268);
and U5550 (N_5550,N_5409,N_5468);
nand U5551 (N_5551,N_5519,N_5457);
and U5552 (N_5552,N_5433,N_5439);
nor U5553 (N_5553,N_5512,N_5465);
xor U5554 (N_5554,N_5510,N_5540);
nand U5555 (N_5555,N_5420,N_5482);
nor U5556 (N_5556,N_5514,N_5506);
nor U5557 (N_5557,N_5546,N_5511);
or U5558 (N_5558,N_5494,N_5531);
and U5559 (N_5559,N_5483,N_5407);
nor U5560 (N_5560,N_5523,N_5455);
or U5561 (N_5561,N_5452,N_5426);
nand U5562 (N_5562,N_5538,N_5470);
and U5563 (N_5563,N_5481,N_5487);
nand U5564 (N_5564,N_5529,N_5497);
xnor U5565 (N_5565,N_5537,N_5499);
nand U5566 (N_5566,N_5411,N_5460);
nand U5567 (N_5567,N_5456,N_5418);
and U5568 (N_5568,N_5535,N_5525);
nor U5569 (N_5569,N_5548,N_5417);
nand U5570 (N_5570,N_5521,N_5400);
nand U5571 (N_5571,N_5508,N_5416);
nor U5572 (N_5572,N_5527,N_5459);
and U5573 (N_5573,N_5545,N_5415);
nand U5574 (N_5574,N_5422,N_5524);
xnor U5575 (N_5575,N_5427,N_5475);
nor U5576 (N_5576,N_5466,N_5450);
nand U5577 (N_5577,N_5408,N_5463);
nand U5578 (N_5578,N_5493,N_5484);
or U5579 (N_5579,N_5443,N_5479);
xor U5580 (N_5580,N_5515,N_5402);
nand U5581 (N_5581,N_5442,N_5403);
nor U5582 (N_5582,N_5448,N_5447);
xor U5583 (N_5583,N_5485,N_5477);
or U5584 (N_5584,N_5489,N_5528);
or U5585 (N_5585,N_5476,N_5478);
nor U5586 (N_5586,N_5539,N_5464);
nor U5587 (N_5587,N_5405,N_5440);
nand U5588 (N_5588,N_5441,N_5530);
and U5589 (N_5589,N_5505,N_5504);
nor U5590 (N_5590,N_5509,N_5517);
nand U5591 (N_5591,N_5516,N_5532);
xnor U5592 (N_5592,N_5549,N_5412);
nand U5593 (N_5593,N_5496,N_5480);
and U5594 (N_5594,N_5469,N_5437);
or U5595 (N_5595,N_5488,N_5471);
xor U5596 (N_5596,N_5503,N_5458);
and U5597 (N_5597,N_5522,N_5401);
xnor U5598 (N_5598,N_5423,N_5453);
or U5599 (N_5599,N_5495,N_5472);
nor U5600 (N_5600,N_5541,N_5436);
nor U5601 (N_5601,N_5547,N_5534);
nor U5602 (N_5602,N_5431,N_5424);
nand U5603 (N_5603,N_5507,N_5518);
nand U5604 (N_5604,N_5490,N_5543);
nand U5605 (N_5605,N_5520,N_5533);
xnor U5606 (N_5606,N_5542,N_5414);
or U5607 (N_5607,N_5501,N_5486);
and U5608 (N_5608,N_5498,N_5445);
nor U5609 (N_5609,N_5526,N_5429);
nand U5610 (N_5610,N_5446,N_5435);
nand U5611 (N_5611,N_5444,N_5474);
nand U5612 (N_5612,N_5461,N_5434);
and U5613 (N_5613,N_5404,N_5544);
nand U5614 (N_5614,N_5410,N_5425);
nand U5615 (N_5615,N_5421,N_5438);
nor U5616 (N_5616,N_5462,N_5454);
or U5617 (N_5617,N_5513,N_5536);
or U5618 (N_5618,N_5492,N_5432);
xor U5619 (N_5619,N_5430,N_5428);
nand U5620 (N_5620,N_5473,N_5449);
xnor U5621 (N_5621,N_5467,N_5419);
and U5622 (N_5622,N_5500,N_5491);
or U5623 (N_5623,N_5413,N_5451);
nor U5624 (N_5624,N_5502,N_5406);
or U5625 (N_5625,N_5518,N_5461);
xor U5626 (N_5626,N_5483,N_5499);
nand U5627 (N_5627,N_5499,N_5488);
xnor U5628 (N_5628,N_5444,N_5462);
xnor U5629 (N_5629,N_5432,N_5483);
or U5630 (N_5630,N_5500,N_5415);
or U5631 (N_5631,N_5460,N_5429);
nand U5632 (N_5632,N_5494,N_5405);
nand U5633 (N_5633,N_5417,N_5509);
nand U5634 (N_5634,N_5529,N_5473);
xnor U5635 (N_5635,N_5448,N_5500);
or U5636 (N_5636,N_5488,N_5460);
nor U5637 (N_5637,N_5503,N_5531);
and U5638 (N_5638,N_5449,N_5415);
nand U5639 (N_5639,N_5506,N_5418);
nor U5640 (N_5640,N_5480,N_5534);
nand U5641 (N_5641,N_5490,N_5409);
and U5642 (N_5642,N_5496,N_5478);
or U5643 (N_5643,N_5481,N_5443);
xnor U5644 (N_5644,N_5484,N_5516);
nand U5645 (N_5645,N_5496,N_5437);
and U5646 (N_5646,N_5538,N_5524);
nand U5647 (N_5647,N_5454,N_5502);
or U5648 (N_5648,N_5400,N_5479);
nor U5649 (N_5649,N_5478,N_5504);
and U5650 (N_5650,N_5470,N_5466);
nor U5651 (N_5651,N_5520,N_5535);
nor U5652 (N_5652,N_5455,N_5494);
nor U5653 (N_5653,N_5546,N_5476);
xor U5654 (N_5654,N_5461,N_5504);
xnor U5655 (N_5655,N_5411,N_5541);
and U5656 (N_5656,N_5415,N_5520);
nor U5657 (N_5657,N_5402,N_5514);
and U5658 (N_5658,N_5438,N_5522);
nand U5659 (N_5659,N_5427,N_5498);
nor U5660 (N_5660,N_5458,N_5444);
nand U5661 (N_5661,N_5401,N_5508);
nor U5662 (N_5662,N_5525,N_5416);
nand U5663 (N_5663,N_5545,N_5494);
nand U5664 (N_5664,N_5442,N_5505);
nand U5665 (N_5665,N_5526,N_5543);
or U5666 (N_5666,N_5400,N_5524);
or U5667 (N_5667,N_5496,N_5477);
nand U5668 (N_5668,N_5479,N_5549);
and U5669 (N_5669,N_5420,N_5410);
xnor U5670 (N_5670,N_5453,N_5455);
nand U5671 (N_5671,N_5527,N_5450);
and U5672 (N_5672,N_5461,N_5512);
xor U5673 (N_5673,N_5485,N_5427);
or U5674 (N_5674,N_5401,N_5498);
nor U5675 (N_5675,N_5449,N_5532);
nand U5676 (N_5676,N_5451,N_5454);
nand U5677 (N_5677,N_5403,N_5468);
and U5678 (N_5678,N_5495,N_5517);
or U5679 (N_5679,N_5491,N_5484);
and U5680 (N_5680,N_5428,N_5535);
nor U5681 (N_5681,N_5524,N_5522);
or U5682 (N_5682,N_5494,N_5511);
or U5683 (N_5683,N_5442,N_5464);
and U5684 (N_5684,N_5486,N_5434);
and U5685 (N_5685,N_5491,N_5460);
or U5686 (N_5686,N_5534,N_5425);
or U5687 (N_5687,N_5478,N_5492);
nand U5688 (N_5688,N_5414,N_5498);
and U5689 (N_5689,N_5541,N_5506);
nor U5690 (N_5690,N_5520,N_5526);
and U5691 (N_5691,N_5533,N_5504);
and U5692 (N_5692,N_5548,N_5431);
nand U5693 (N_5693,N_5496,N_5514);
nor U5694 (N_5694,N_5406,N_5404);
xnor U5695 (N_5695,N_5445,N_5452);
or U5696 (N_5696,N_5544,N_5470);
and U5697 (N_5697,N_5442,N_5407);
xor U5698 (N_5698,N_5425,N_5485);
nand U5699 (N_5699,N_5539,N_5512);
or U5700 (N_5700,N_5562,N_5639);
nor U5701 (N_5701,N_5618,N_5597);
or U5702 (N_5702,N_5690,N_5669);
xor U5703 (N_5703,N_5647,N_5564);
nand U5704 (N_5704,N_5572,N_5590);
and U5705 (N_5705,N_5699,N_5698);
xnor U5706 (N_5706,N_5687,N_5579);
or U5707 (N_5707,N_5633,N_5644);
nand U5708 (N_5708,N_5688,N_5552);
and U5709 (N_5709,N_5568,N_5640);
and U5710 (N_5710,N_5580,N_5569);
or U5711 (N_5711,N_5682,N_5575);
xor U5712 (N_5712,N_5595,N_5660);
nand U5713 (N_5713,N_5620,N_5646);
and U5714 (N_5714,N_5630,N_5599);
or U5715 (N_5715,N_5631,N_5592);
and U5716 (N_5716,N_5654,N_5606);
and U5717 (N_5717,N_5655,N_5675);
nor U5718 (N_5718,N_5604,N_5672);
nand U5719 (N_5719,N_5612,N_5574);
nor U5720 (N_5720,N_5673,N_5679);
and U5721 (N_5721,N_5670,N_5615);
and U5722 (N_5722,N_5676,N_5627);
or U5723 (N_5723,N_5634,N_5591);
or U5724 (N_5724,N_5628,N_5653);
nor U5725 (N_5725,N_5645,N_5567);
nand U5726 (N_5726,N_5658,N_5680);
or U5727 (N_5727,N_5608,N_5617);
xnor U5728 (N_5728,N_5603,N_5684);
xor U5729 (N_5729,N_5555,N_5593);
nand U5730 (N_5730,N_5689,N_5588);
xor U5731 (N_5731,N_5600,N_5616);
nand U5732 (N_5732,N_5661,N_5561);
nor U5733 (N_5733,N_5678,N_5641);
or U5734 (N_5734,N_5621,N_5659);
or U5735 (N_5735,N_5611,N_5551);
and U5736 (N_5736,N_5586,N_5582);
and U5737 (N_5737,N_5666,N_5554);
or U5738 (N_5738,N_5607,N_5570);
or U5739 (N_5739,N_5576,N_5565);
nand U5740 (N_5740,N_5587,N_5610);
nand U5741 (N_5741,N_5692,N_5636);
and U5742 (N_5742,N_5671,N_5663);
nor U5743 (N_5743,N_5697,N_5695);
or U5744 (N_5744,N_5667,N_5609);
and U5745 (N_5745,N_5638,N_5553);
or U5746 (N_5746,N_5559,N_5683);
nand U5747 (N_5747,N_5601,N_5623);
nor U5748 (N_5748,N_5557,N_5693);
or U5749 (N_5749,N_5665,N_5598);
nand U5750 (N_5750,N_5668,N_5625);
and U5751 (N_5751,N_5556,N_5632);
nor U5752 (N_5752,N_5581,N_5573);
nand U5753 (N_5753,N_5691,N_5635);
nand U5754 (N_5754,N_5614,N_5657);
xor U5755 (N_5755,N_5578,N_5594);
xor U5756 (N_5756,N_5681,N_5677);
nand U5757 (N_5757,N_5651,N_5696);
nor U5758 (N_5758,N_5649,N_5656);
or U5759 (N_5759,N_5566,N_5642);
and U5760 (N_5760,N_5605,N_5626);
and U5761 (N_5761,N_5685,N_5662);
or U5762 (N_5762,N_5560,N_5613);
or U5763 (N_5763,N_5674,N_5652);
and U5764 (N_5764,N_5629,N_5637);
nand U5765 (N_5765,N_5694,N_5686);
nor U5766 (N_5766,N_5622,N_5571);
or U5767 (N_5767,N_5577,N_5648);
nor U5768 (N_5768,N_5602,N_5584);
or U5769 (N_5769,N_5589,N_5624);
nor U5770 (N_5770,N_5550,N_5585);
xor U5771 (N_5771,N_5583,N_5650);
and U5772 (N_5772,N_5558,N_5619);
xor U5773 (N_5773,N_5664,N_5596);
xnor U5774 (N_5774,N_5563,N_5643);
nand U5775 (N_5775,N_5557,N_5597);
xnor U5776 (N_5776,N_5664,N_5670);
and U5777 (N_5777,N_5636,N_5560);
or U5778 (N_5778,N_5563,N_5672);
xor U5779 (N_5779,N_5608,N_5578);
nor U5780 (N_5780,N_5626,N_5629);
nor U5781 (N_5781,N_5686,N_5665);
or U5782 (N_5782,N_5576,N_5610);
or U5783 (N_5783,N_5587,N_5646);
or U5784 (N_5784,N_5634,N_5571);
nand U5785 (N_5785,N_5615,N_5626);
nand U5786 (N_5786,N_5575,N_5689);
or U5787 (N_5787,N_5618,N_5646);
nand U5788 (N_5788,N_5694,N_5647);
nor U5789 (N_5789,N_5648,N_5576);
or U5790 (N_5790,N_5569,N_5699);
xnor U5791 (N_5791,N_5601,N_5615);
xnor U5792 (N_5792,N_5565,N_5695);
and U5793 (N_5793,N_5591,N_5602);
nor U5794 (N_5794,N_5632,N_5625);
nor U5795 (N_5795,N_5647,N_5667);
xor U5796 (N_5796,N_5639,N_5626);
or U5797 (N_5797,N_5634,N_5605);
and U5798 (N_5798,N_5687,N_5581);
nand U5799 (N_5799,N_5575,N_5645);
nand U5800 (N_5800,N_5556,N_5637);
nor U5801 (N_5801,N_5568,N_5635);
xnor U5802 (N_5802,N_5596,N_5629);
and U5803 (N_5803,N_5696,N_5614);
or U5804 (N_5804,N_5699,N_5597);
nand U5805 (N_5805,N_5654,N_5662);
nor U5806 (N_5806,N_5565,N_5659);
xnor U5807 (N_5807,N_5681,N_5619);
nand U5808 (N_5808,N_5697,N_5676);
xor U5809 (N_5809,N_5565,N_5637);
or U5810 (N_5810,N_5587,N_5687);
xor U5811 (N_5811,N_5604,N_5611);
and U5812 (N_5812,N_5589,N_5616);
xnor U5813 (N_5813,N_5645,N_5631);
nand U5814 (N_5814,N_5617,N_5669);
nand U5815 (N_5815,N_5602,N_5660);
or U5816 (N_5816,N_5629,N_5589);
xnor U5817 (N_5817,N_5667,N_5639);
xnor U5818 (N_5818,N_5670,N_5661);
and U5819 (N_5819,N_5610,N_5698);
or U5820 (N_5820,N_5657,N_5673);
nand U5821 (N_5821,N_5552,N_5671);
or U5822 (N_5822,N_5609,N_5652);
nor U5823 (N_5823,N_5561,N_5573);
xnor U5824 (N_5824,N_5588,N_5662);
nand U5825 (N_5825,N_5587,N_5699);
and U5826 (N_5826,N_5688,N_5598);
or U5827 (N_5827,N_5565,N_5550);
or U5828 (N_5828,N_5566,N_5652);
nor U5829 (N_5829,N_5640,N_5654);
or U5830 (N_5830,N_5680,N_5617);
and U5831 (N_5831,N_5573,N_5623);
nand U5832 (N_5832,N_5689,N_5692);
or U5833 (N_5833,N_5587,N_5618);
nor U5834 (N_5834,N_5676,N_5668);
or U5835 (N_5835,N_5696,N_5670);
or U5836 (N_5836,N_5638,N_5682);
nor U5837 (N_5837,N_5622,N_5568);
nand U5838 (N_5838,N_5672,N_5688);
nor U5839 (N_5839,N_5616,N_5662);
and U5840 (N_5840,N_5568,N_5684);
xor U5841 (N_5841,N_5669,N_5563);
and U5842 (N_5842,N_5591,N_5697);
nand U5843 (N_5843,N_5676,N_5643);
and U5844 (N_5844,N_5577,N_5651);
nor U5845 (N_5845,N_5580,N_5637);
nor U5846 (N_5846,N_5686,N_5584);
xor U5847 (N_5847,N_5554,N_5609);
nor U5848 (N_5848,N_5648,N_5665);
nand U5849 (N_5849,N_5625,N_5609);
and U5850 (N_5850,N_5792,N_5772);
or U5851 (N_5851,N_5821,N_5709);
xor U5852 (N_5852,N_5779,N_5769);
nand U5853 (N_5853,N_5719,N_5740);
and U5854 (N_5854,N_5758,N_5711);
xor U5855 (N_5855,N_5754,N_5773);
or U5856 (N_5856,N_5729,N_5759);
or U5857 (N_5857,N_5734,N_5753);
or U5858 (N_5858,N_5789,N_5733);
nand U5859 (N_5859,N_5712,N_5785);
xnor U5860 (N_5860,N_5846,N_5768);
nor U5861 (N_5861,N_5722,N_5765);
xor U5862 (N_5862,N_5700,N_5715);
xnor U5863 (N_5863,N_5757,N_5732);
and U5864 (N_5864,N_5811,N_5836);
and U5865 (N_5865,N_5707,N_5763);
nor U5866 (N_5866,N_5752,N_5832);
nand U5867 (N_5867,N_5831,N_5736);
nor U5868 (N_5868,N_5805,N_5749);
nand U5869 (N_5869,N_5844,N_5784);
nand U5870 (N_5870,N_5822,N_5783);
or U5871 (N_5871,N_5841,N_5760);
xnor U5872 (N_5872,N_5848,N_5817);
nor U5873 (N_5873,N_5737,N_5816);
xnor U5874 (N_5874,N_5703,N_5721);
nor U5875 (N_5875,N_5748,N_5750);
nor U5876 (N_5876,N_5835,N_5812);
nor U5877 (N_5877,N_5714,N_5786);
xor U5878 (N_5878,N_5813,N_5744);
xor U5879 (N_5879,N_5826,N_5718);
xnor U5880 (N_5880,N_5825,N_5807);
nand U5881 (N_5881,N_5771,N_5837);
and U5882 (N_5882,N_5818,N_5815);
nand U5883 (N_5883,N_5770,N_5782);
xnor U5884 (N_5884,N_5702,N_5706);
or U5885 (N_5885,N_5775,N_5761);
or U5886 (N_5886,N_5746,N_5777);
nand U5887 (N_5887,N_5845,N_5730);
nor U5888 (N_5888,N_5767,N_5745);
nor U5889 (N_5889,N_5728,N_5755);
or U5890 (N_5890,N_5781,N_5849);
or U5891 (N_5891,N_5738,N_5796);
nor U5892 (N_5892,N_5791,N_5814);
and U5893 (N_5893,N_5806,N_5833);
xnor U5894 (N_5894,N_5823,N_5820);
and U5895 (N_5895,N_5762,N_5801);
and U5896 (N_5896,N_5838,N_5751);
or U5897 (N_5897,N_5793,N_5809);
xor U5898 (N_5898,N_5827,N_5705);
xor U5899 (N_5899,N_5834,N_5704);
nor U5900 (N_5900,N_5735,N_5724);
xnor U5901 (N_5901,N_5778,N_5725);
xor U5902 (N_5902,N_5799,N_5808);
and U5903 (N_5903,N_5731,N_5824);
xnor U5904 (N_5904,N_5787,N_5743);
nand U5905 (N_5905,N_5830,N_5804);
and U5906 (N_5906,N_5795,N_5739);
nand U5907 (N_5907,N_5747,N_5726);
nor U5908 (N_5908,N_5766,N_5727);
or U5909 (N_5909,N_5829,N_5794);
nor U5910 (N_5910,N_5840,N_5847);
or U5911 (N_5911,N_5716,N_5828);
xnor U5912 (N_5912,N_5810,N_5776);
and U5913 (N_5913,N_5774,N_5741);
or U5914 (N_5914,N_5710,N_5788);
nand U5915 (N_5915,N_5764,N_5839);
nor U5916 (N_5916,N_5797,N_5803);
nand U5917 (N_5917,N_5842,N_5701);
and U5918 (N_5918,N_5819,N_5742);
or U5919 (N_5919,N_5723,N_5780);
or U5920 (N_5920,N_5802,N_5713);
xnor U5921 (N_5921,N_5720,N_5800);
xor U5922 (N_5922,N_5798,N_5790);
nor U5923 (N_5923,N_5756,N_5717);
or U5924 (N_5924,N_5708,N_5843);
nor U5925 (N_5925,N_5756,N_5791);
nand U5926 (N_5926,N_5844,N_5713);
nor U5927 (N_5927,N_5760,N_5706);
nand U5928 (N_5928,N_5768,N_5804);
or U5929 (N_5929,N_5778,N_5728);
nand U5930 (N_5930,N_5723,N_5787);
nand U5931 (N_5931,N_5759,N_5827);
xor U5932 (N_5932,N_5713,N_5798);
xnor U5933 (N_5933,N_5700,N_5797);
or U5934 (N_5934,N_5808,N_5718);
xnor U5935 (N_5935,N_5755,N_5749);
or U5936 (N_5936,N_5730,N_5795);
nor U5937 (N_5937,N_5731,N_5753);
xor U5938 (N_5938,N_5702,N_5786);
nand U5939 (N_5939,N_5784,N_5811);
and U5940 (N_5940,N_5791,N_5701);
nand U5941 (N_5941,N_5756,N_5731);
xor U5942 (N_5942,N_5723,N_5841);
nor U5943 (N_5943,N_5831,N_5730);
and U5944 (N_5944,N_5769,N_5777);
or U5945 (N_5945,N_5766,N_5776);
or U5946 (N_5946,N_5831,N_5742);
or U5947 (N_5947,N_5839,N_5759);
or U5948 (N_5948,N_5704,N_5805);
nor U5949 (N_5949,N_5813,N_5843);
nor U5950 (N_5950,N_5837,N_5778);
nor U5951 (N_5951,N_5758,N_5780);
nand U5952 (N_5952,N_5766,N_5809);
nor U5953 (N_5953,N_5751,N_5761);
and U5954 (N_5954,N_5803,N_5770);
and U5955 (N_5955,N_5715,N_5749);
nor U5956 (N_5956,N_5739,N_5809);
nor U5957 (N_5957,N_5813,N_5721);
nand U5958 (N_5958,N_5802,N_5765);
and U5959 (N_5959,N_5703,N_5724);
or U5960 (N_5960,N_5713,N_5748);
nand U5961 (N_5961,N_5766,N_5724);
nand U5962 (N_5962,N_5846,N_5710);
nand U5963 (N_5963,N_5776,N_5830);
nor U5964 (N_5964,N_5776,N_5783);
or U5965 (N_5965,N_5817,N_5725);
nor U5966 (N_5966,N_5732,N_5731);
nand U5967 (N_5967,N_5818,N_5763);
nor U5968 (N_5968,N_5769,N_5826);
and U5969 (N_5969,N_5708,N_5775);
xnor U5970 (N_5970,N_5759,N_5772);
nor U5971 (N_5971,N_5839,N_5760);
and U5972 (N_5972,N_5767,N_5837);
nor U5973 (N_5973,N_5796,N_5777);
xnor U5974 (N_5974,N_5757,N_5820);
or U5975 (N_5975,N_5768,N_5786);
and U5976 (N_5976,N_5712,N_5811);
nand U5977 (N_5977,N_5845,N_5822);
or U5978 (N_5978,N_5700,N_5728);
and U5979 (N_5979,N_5713,N_5797);
nor U5980 (N_5980,N_5815,N_5827);
and U5981 (N_5981,N_5773,N_5726);
xnor U5982 (N_5982,N_5784,N_5794);
nand U5983 (N_5983,N_5771,N_5815);
nor U5984 (N_5984,N_5740,N_5717);
nor U5985 (N_5985,N_5804,N_5798);
and U5986 (N_5986,N_5800,N_5795);
nand U5987 (N_5987,N_5720,N_5792);
nor U5988 (N_5988,N_5771,N_5709);
nand U5989 (N_5989,N_5726,N_5775);
xor U5990 (N_5990,N_5783,N_5816);
and U5991 (N_5991,N_5763,N_5781);
or U5992 (N_5992,N_5794,N_5772);
or U5993 (N_5993,N_5706,N_5816);
or U5994 (N_5994,N_5792,N_5789);
nand U5995 (N_5995,N_5838,N_5770);
or U5996 (N_5996,N_5792,N_5821);
nor U5997 (N_5997,N_5745,N_5709);
nor U5998 (N_5998,N_5736,N_5792);
xnor U5999 (N_5999,N_5746,N_5775);
or U6000 (N_6000,N_5902,N_5928);
nor U6001 (N_6001,N_5964,N_5852);
and U6002 (N_6002,N_5882,N_5944);
nand U6003 (N_6003,N_5867,N_5985);
xnor U6004 (N_6004,N_5924,N_5983);
and U6005 (N_6005,N_5996,N_5977);
and U6006 (N_6006,N_5901,N_5949);
nor U6007 (N_6007,N_5921,N_5961);
nand U6008 (N_6008,N_5870,N_5969);
or U6009 (N_6009,N_5932,N_5879);
and U6010 (N_6010,N_5945,N_5970);
nand U6011 (N_6011,N_5871,N_5911);
xor U6012 (N_6012,N_5929,N_5873);
xnor U6013 (N_6013,N_5981,N_5965);
and U6014 (N_6014,N_5860,N_5880);
nor U6015 (N_6015,N_5923,N_5994);
and U6016 (N_6016,N_5861,N_5872);
xor U6017 (N_6017,N_5858,N_5973);
and U6018 (N_6018,N_5941,N_5998);
nor U6019 (N_6019,N_5982,N_5884);
or U6020 (N_6020,N_5963,N_5895);
nor U6021 (N_6021,N_5937,N_5933);
nor U6022 (N_6022,N_5952,N_5908);
or U6023 (N_6023,N_5859,N_5905);
or U6024 (N_6024,N_5894,N_5980);
nor U6025 (N_6025,N_5883,N_5925);
or U6026 (N_6026,N_5974,N_5976);
and U6027 (N_6027,N_5966,N_5854);
nand U6028 (N_6028,N_5938,N_5986);
and U6029 (N_6029,N_5865,N_5891);
or U6030 (N_6030,N_5997,N_5857);
nand U6031 (N_6031,N_5907,N_5958);
nor U6032 (N_6032,N_5885,N_5991);
and U6033 (N_6033,N_5878,N_5897);
nor U6034 (N_6034,N_5900,N_5943);
nand U6035 (N_6035,N_5864,N_5990);
xnor U6036 (N_6036,N_5947,N_5868);
xnor U6037 (N_6037,N_5888,N_5971);
nor U6038 (N_6038,N_5934,N_5919);
or U6039 (N_6039,N_5850,N_5893);
xor U6040 (N_6040,N_5851,N_5910);
nor U6041 (N_6041,N_5917,N_5914);
xor U6042 (N_6042,N_5862,N_5909);
or U6043 (N_6043,N_5940,N_5993);
and U6044 (N_6044,N_5877,N_5951);
xor U6045 (N_6045,N_5960,N_5992);
nor U6046 (N_6046,N_5954,N_5922);
nand U6047 (N_6047,N_5984,N_5959);
xor U6048 (N_6048,N_5967,N_5866);
and U6049 (N_6049,N_5892,N_5875);
xor U6050 (N_6050,N_5926,N_5968);
nor U6051 (N_6051,N_5957,N_5989);
nor U6052 (N_6052,N_5913,N_5927);
nor U6053 (N_6053,N_5881,N_5904);
or U6054 (N_6054,N_5979,N_5930);
nor U6055 (N_6055,N_5931,N_5935);
xor U6056 (N_6056,N_5978,N_5950);
nand U6057 (N_6057,N_5918,N_5999);
and U6058 (N_6058,N_5939,N_5874);
and U6059 (N_6059,N_5896,N_5899);
xor U6060 (N_6060,N_5886,N_5987);
nor U6061 (N_6061,N_5876,N_5995);
and U6062 (N_6062,N_5915,N_5863);
or U6063 (N_6063,N_5898,N_5856);
nand U6064 (N_6064,N_5912,N_5948);
xnor U6065 (N_6065,N_5890,N_5920);
xnor U6066 (N_6066,N_5853,N_5906);
xnor U6067 (N_6067,N_5975,N_5855);
nor U6068 (N_6068,N_5936,N_5942);
xnor U6069 (N_6069,N_5903,N_5955);
and U6070 (N_6070,N_5962,N_5916);
xnor U6071 (N_6071,N_5889,N_5946);
nor U6072 (N_6072,N_5956,N_5887);
and U6073 (N_6073,N_5869,N_5972);
and U6074 (N_6074,N_5988,N_5953);
and U6075 (N_6075,N_5949,N_5906);
xnor U6076 (N_6076,N_5896,N_5910);
nor U6077 (N_6077,N_5870,N_5899);
or U6078 (N_6078,N_5930,N_5946);
and U6079 (N_6079,N_5961,N_5881);
xor U6080 (N_6080,N_5867,N_5853);
nor U6081 (N_6081,N_5890,N_5925);
nor U6082 (N_6082,N_5905,N_5975);
nor U6083 (N_6083,N_5897,N_5909);
nor U6084 (N_6084,N_5864,N_5908);
or U6085 (N_6085,N_5884,N_5932);
or U6086 (N_6086,N_5971,N_5988);
and U6087 (N_6087,N_5875,N_5951);
or U6088 (N_6088,N_5906,N_5953);
nor U6089 (N_6089,N_5922,N_5873);
or U6090 (N_6090,N_5956,N_5851);
nand U6091 (N_6091,N_5879,N_5911);
and U6092 (N_6092,N_5977,N_5945);
nand U6093 (N_6093,N_5875,N_5911);
xor U6094 (N_6094,N_5946,N_5873);
nand U6095 (N_6095,N_5987,N_5894);
or U6096 (N_6096,N_5873,N_5866);
xnor U6097 (N_6097,N_5940,N_5851);
nor U6098 (N_6098,N_5864,N_5929);
nand U6099 (N_6099,N_5981,N_5888);
and U6100 (N_6100,N_5992,N_5977);
or U6101 (N_6101,N_5872,N_5978);
or U6102 (N_6102,N_5918,N_5910);
nand U6103 (N_6103,N_5907,N_5997);
nor U6104 (N_6104,N_5881,N_5920);
nand U6105 (N_6105,N_5981,N_5948);
xnor U6106 (N_6106,N_5928,N_5949);
or U6107 (N_6107,N_5853,N_5899);
or U6108 (N_6108,N_5887,N_5884);
and U6109 (N_6109,N_5925,N_5863);
or U6110 (N_6110,N_5982,N_5890);
xnor U6111 (N_6111,N_5948,N_5970);
nor U6112 (N_6112,N_5857,N_5859);
or U6113 (N_6113,N_5888,N_5853);
nor U6114 (N_6114,N_5852,N_5884);
xnor U6115 (N_6115,N_5947,N_5864);
xnor U6116 (N_6116,N_5984,N_5919);
nand U6117 (N_6117,N_5904,N_5996);
and U6118 (N_6118,N_5861,N_5941);
and U6119 (N_6119,N_5990,N_5949);
or U6120 (N_6120,N_5929,N_5852);
xnor U6121 (N_6121,N_5982,N_5973);
xor U6122 (N_6122,N_5898,N_5869);
nor U6123 (N_6123,N_5998,N_5909);
xor U6124 (N_6124,N_5997,N_5938);
and U6125 (N_6125,N_5887,N_5983);
nand U6126 (N_6126,N_5869,N_5955);
nand U6127 (N_6127,N_5915,N_5878);
nor U6128 (N_6128,N_5855,N_5950);
xor U6129 (N_6129,N_5932,N_5970);
nand U6130 (N_6130,N_5934,N_5955);
nor U6131 (N_6131,N_5928,N_5867);
nand U6132 (N_6132,N_5874,N_5883);
and U6133 (N_6133,N_5859,N_5987);
nand U6134 (N_6134,N_5881,N_5889);
and U6135 (N_6135,N_5945,N_5926);
or U6136 (N_6136,N_5902,N_5959);
and U6137 (N_6137,N_5989,N_5917);
nand U6138 (N_6138,N_5888,N_5942);
and U6139 (N_6139,N_5962,N_5917);
or U6140 (N_6140,N_5994,N_5943);
and U6141 (N_6141,N_5994,N_5946);
and U6142 (N_6142,N_5953,N_5966);
xor U6143 (N_6143,N_5953,N_5998);
nor U6144 (N_6144,N_5928,N_5885);
xor U6145 (N_6145,N_5951,N_5904);
nor U6146 (N_6146,N_5960,N_5854);
or U6147 (N_6147,N_5973,N_5953);
nand U6148 (N_6148,N_5957,N_5927);
nand U6149 (N_6149,N_5922,N_5912);
and U6150 (N_6150,N_6100,N_6065);
or U6151 (N_6151,N_6058,N_6128);
nand U6152 (N_6152,N_6105,N_6042);
nand U6153 (N_6153,N_6020,N_6034);
xor U6154 (N_6154,N_6113,N_6007);
nand U6155 (N_6155,N_6006,N_6102);
xnor U6156 (N_6156,N_6135,N_6056);
and U6157 (N_6157,N_6032,N_6000);
and U6158 (N_6158,N_6131,N_6144);
nor U6159 (N_6159,N_6112,N_6103);
nand U6160 (N_6160,N_6010,N_6090);
and U6161 (N_6161,N_6035,N_6141);
or U6162 (N_6162,N_6067,N_6149);
and U6163 (N_6163,N_6108,N_6088);
nand U6164 (N_6164,N_6138,N_6059);
xnor U6165 (N_6165,N_6029,N_6092);
and U6166 (N_6166,N_6040,N_6075);
nor U6167 (N_6167,N_6147,N_6039);
and U6168 (N_6168,N_6097,N_6051);
xnor U6169 (N_6169,N_6085,N_6049);
and U6170 (N_6170,N_6081,N_6120);
and U6171 (N_6171,N_6046,N_6036);
nand U6172 (N_6172,N_6134,N_6025);
and U6173 (N_6173,N_6122,N_6133);
nor U6174 (N_6174,N_6082,N_6142);
nand U6175 (N_6175,N_6004,N_6009);
xnor U6176 (N_6176,N_6139,N_6084);
nand U6177 (N_6177,N_6037,N_6143);
or U6178 (N_6178,N_6031,N_6012);
or U6179 (N_6179,N_6048,N_6132);
nor U6180 (N_6180,N_6109,N_6117);
or U6181 (N_6181,N_6096,N_6123);
xnor U6182 (N_6182,N_6064,N_6001);
nand U6183 (N_6183,N_6045,N_6083);
nor U6184 (N_6184,N_6003,N_6060);
and U6185 (N_6185,N_6079,N_6073);
nand U6186 (N_6186,N_6129,N_6107);
nor U6187 (N_6187,N_6118,N_6137);
xor U6188 (N_6188,N_6019,N_6023);
or U6189 (N_6189,N_6005,N_6057);
nand U6190 (N_6190,N_6070,N_6086);
xnor U6191 (N_6191,N_6115,N_6033);
and U6192 (N_6192,N_6047,N_6018);
nor U6193 (N_6193,N_6078,N_6026);
or U6194 (N_6194,N_6013,N_6072);
and U6195 (N_6195,N_6024,N_6061);
or U6196 (N_6196,N_6095,N_6038);
xnor U6197 (N_6197,N_6021,N_6077);
and U6198 (N_6198,N_6146,N_6098);
or U6199 (N_6199,N_6053,N_6022);
or U6200 (N_6200,N_6080,N_6099);
xnor U6201 (N_6201,N_6041,N_6114);
nor U6202 (N_6202,N_6027,N_6148);
nor U6203 (N_6203,N_6011,N_6101);
or U6204 (N_6204,N_6028,N_6126);
or U6205 (N_6205,N_6044,N_6014);
xnor U6206 (N_6206,N_6091,N_6069);
and U6207 (N_6207,N_6136,N_6050);
nor U6208 (N_6208,N_6062,N_6110);
and U6209 (N_6209,N_6043,N_6055);
nand U6210 (N_6210,N_6130,N_6016);
or U6211 (N_6211,N_6093,N_6119);
xor U6212 (N_6212,N_6104,N_6017);
or U6213 (N_6213,N_6052,N_6071);
nor U6214 (N_6214,N_6106,N_6111);
nand U6215 (N_6215,N_6066,N_6127);
xnor U6216 (N_6216,N_6015,N_6125);
xnor U6217 (N_6217,N_6124,N_6068);
nand U6218 (N_6218,N_6087,N_6145);
xor U6219 (N_6219,N_6116,N_6074);
and U6220 (N_6220,N_6094,N_6054);
nor U6221 (N_6221,N_6008,N_6089);
xnor U6222 (N_6222,N_6140,N_6002);
or U6223 (N_6223,N_6076,N_6063);
nand U6224 (N_6224,N_6030,N_6121);
or U6225 (N_6225,N_6012,N_6136);
nor U6226 (N_6226,N_6083,N_6095);
or U6227 (N_6227,N_6057,N_6089);
nor U6228 (N_6228,N_6126,N_6045);
or U6229 (N_6229,N_6000,N_6001);
xor U6230 (N_6230,N_6061,N_6056);
nor U6231 (N_6231,N_6111,N_6142);
or U6232 (N_6232,N_6107,N_6111);
and U6233 (N_6233,N_6122,N_6008);
nand U6234 (N_6234,N_6080,N_6059);
nand U6235 (N_6235,N_6004,N_6124);
nor U6236 (N_6236,N_6107,N_6025);
and U6237 (N_6237,N_6074,N_6050);
or U6238 (N_6238,N_6020,N_6146);
or U6239 (N_6239,N_6039,N_6000);
nor U6240 (N_6240,N_6139,N_6134);
xnor U6241 (N_6241,N_6068,N_6006);
and U6242 (N_6242,N_6067,N_6001);
or U6243 (N_6243,N_6018,N_6091);
and U6244 (N_6244,N_6133,N_6145);
xor U6245 (N_6245,N_6081,N_6030);
nand U6246 (N_6246,N_6064,N_6040);
and U6247 (N_6247,N_6062,N_6094);
nand U6248 (N_6248,N_6045,N_6027);
and U6249 (N_6249,N_6056,N_6031);
or U6250 (N_6250,N_6067,N_6037);
nand U6251 (N_6251,N_6053,N_6091);
or U6252 (N_6252,N_6103,N_6114);
nand U6253 (N_6253,N_6112,N_6138);
nand U6254 (N_6254,N_6090,N_6101);
nand U6255 (N_6255,N_6136,N_6101);
nand U6256 (N_6256,N_6122,N_6125);
and U6257 (N_6257,N_6110,N_6081);
and U6258 (N_6258,N_6117,N_6122);
or U6259 (N_6259,N_6031,N_6075);
nand U6260 (N_6260,N_6145,N_6146);
and U6261 (N_6261,N_6000,N_6085);
and U6262 (N_6262,N_6116,N_6001);
and U6263 (N_6263,N_6124,N_6023);
nand U6264 (N_6264,N_6045,N_6110);
nand U6265 (N_6265,N_6129,N_6090);
xnor U6266 (N_6266,N_6145,N_6137);
xnor U6267 (N_6267,N_6009,N_6139);
nor U6268 (N_6268,N_6113,N_6104);
or U6269 (N_6269,N_6032,N_6057);
xor U6270 (N_6270,N_6004,N_6138);
or U6271 (N_6271,N_6119,N_6085);
nor U6272 (N_6272,N_6004,N_6018);
nor U6273 (N_6273,N_6077,N_6018);
and U6274 (N_6274,N_6057,N_6098);
nor U6275 (N_6275,N_6060,N_6019);
nand U6276 (N_6276,N_6035,N_6025);
or U6277 (N_6277,N_6058,N_6067);
and U6278 (N_6278,N_6124,N_6055);
or U6279 (N_6279,N_6006,N_6031);
nor U6280 (N_6280,N_6106,N_6135);
nand U6281 (N_6281,N_6131,N_6114);
and U6282 (N_6282,N_6012,N_6026);
and U6283 (N_6283,N_6045,N_6012);
and U6284 (N_6284,N_6002,N_6118);
and U6285 (N_6285,N_6026,N_6089);
and U6286 (N_6286,N_6145,N_6132);
xnor U6287 (N_6287,N_6026,N_6008);
nor U6288 (N_6288,N_6076,N_6050);
nand U6289 (N_6289,N_6143,N_6049);
and U6290 (N_6290,N_6072,N_6083);
xor U6291 (N_6291,N_6068,N_6055);
xnor U6292 (N_6292,N_6013,N_6038);
and U6293 (N_6293,N_6128,N_6045);
nor U6294 (N_6294,N_6066,N_6083);
nor U6295 (N_6295,N_6010,N_6116);
nor U6296 (N_6296,N_6092,N_6106);
and U6297 (N_6297,N_6140,N_6107);
or U6298 (N_6298,N_6139,N_6108);
or U6299 (N_6299,N_6098,N_6020);
and U6300 (N_6300,N_6187,N_6198);
nor U6301 (N_6301,N_6202,N_6270);
and U6302 (N_6302,N_6190,N_6163);
nor U6303 (N_6303,N_6218,N_6257);
nand U6304 (N_6304,N_6228,N_6231);
nor U6305 (N_6305,N_6237,N_6253);
or U6306 (N_6306,N_6211,N_6291);
or U6307 (N_6307,N_6289,N_6244);
nand U6308 (N_6308,N_6246,N_6293);
nor U6309 (N_6309,N_6220,N_6241);
xor U6310 (N_6310,N_6155,N_6171);
and U6311 (N_6311,N_6267,N_6297);
and U6312 (N_6312,N_6227,N_6156);
or U6313 (N_6313,N_6199,N_6154);
xnor U6314 (N_6314,N_6252,N_6200);
or U6315 (N_6315,N_6229,N_6217);
or U6316 (N_6316,N_6185,N_6181);
nor U6317 (N_6317,N_6260,N_6197);
xor U6318 (N_6318,N_6283,N_6168);
nor U6319 (N_6319,N_6150,N_6159);
or U6320 (N_6320,N_6207,N_6284);
or U6321 (N_6321,N_6261,N_6295);
nand U6322 (N_6322,N_6279,N_6161);
nor U6323 (N_6323,N_6194,N_6269);
nor U6324 (N_6324,N_6235,N_6255);
and U6325 (N_6325,N_6280,N_6292);
nor U6326 (N_6326,N_6205,N_6240);
and U6327 (N_6327,N_6184,N_6183);
and U6328 (N_6328,N_6273,N_6251);
nor U6329 (N_6329,N_6214,N_6243);
or U6330 (N_6330,N_6151,N_6296);
nand U6331 (N_6331,N_6285,N_6272);
or U6332 (N_6332,N_6271,N_6264);
nor U6333 (N_6333,N_6206,N_6233);
and U6334 (N_6334,N_6204,N_6176);
nand U6335 (N_6335,N_6274,N_6172);
nand U6336 (N_6336,N_6212,N_6188);
and U6337 (N_6337,N_6278,N_6238);
nor U6338 (N_6338,N_6234,N_6216);
and U6339 (N_6339,N_6262,N_6173);
xnor U6340 (N_6340,N_6175,N_6281);
nand U6341 (N_6341,N_6203,N_6258);
xnor U6342 (N_6342,N_6230,N_6288);
nor U6343 (N_6343,N_6165,N_6208);
or U6344 (N_6344,N_6196,N_6282);
xnor U6345 (N_6345,N_6191,N_6213);
xor U6346 (N_6346,N_6201,N_6223);
xnor U6347 (N_6347,N_6286,N_6167);
and U6348 (N_6348,N_6265,N_6169);
nor U6349 (N_6349,N_6189,N_6226);
or U6350 (N_6350,N_6178,N_6225);
and U6351 (N_6351,N_6298,N_6290);
and U6352 (N_6352,N_6254,N_6209);
and U6353 (N_6353,N_6236,N_6164);
nor U6354 (N_6354,N_6166,N_6256);
nor U6355 (N_6355,N_6268,N_6222);
nand U6356 (N_6356,N_6250,N_6245);
and U6357 (N_6357,N_6275,N_6186);
nand U6358 (N_6358,N_6180,N_6259);
nand U6359 (N_6359,N_6210,N_6294);
and U6360 (N_6360,N_6239,N_6193);
xor U6361 (N_6361,N_6263,N_6224);
xnor U6362 (N_6362,N_6221,N_6299);
and U6363 (N_6363,N_6174,N_6287);
or U6364 (N_6364,N_6162,N_6153);
nand U6365 (N_6365,N_6219,N_6232);
and U6366 (N_6366,N_6215,N_6157);
and U6367 (N_6367,N_6242,N_6160);
or U6368 (N_6368,N_6249,N_6158);
xnor U6369 (N_6369,N_6247,N_6266);
or U6370 (N_6370,N_6248,N_6179);
xor U6371 (N_6371,N_6177,N_6276);
xor U6372 (N_6372,N_6182,N_6277);
and U6373 (N_6373,N_6192,N_6170);
and U6374 (N_6374,N_6152,N_6195);
xor U6375 (N_6375,N_6235,N_6153);
nor U6376 (N_6376,N_6289,N_6268);
or U6377 (N_6377,N_6196,N_6179);
and U6378 (N_6378,N_6216,N_6261);
xor U6379 (N_6379,N_6203,N_6249);
xnor U6380 (N_6380,N_6231,N_6201);
nand U6381 (N_6381,N_6251,N_6252);
nand U6382 (N_6382,N_6267,N_6190);
xor U6383 (N_6383,N_6216,N_6232);
xnor U6384 (N_6384,N_6221,N_6286);
nor U6385 (N_6385,N_6229,N_6173);
and U6386 (N_6386,N_6259,N_6172);
nor U6387 (N_6387,N_6225,N_6268);
xor U6388 (N_6388,N_6219,N_6165);
nand U6389 (N_6389,N_6260,N_6188);
nand U6390 (N_6390,N_6297,N_6152);
or U6391 (N_6391,N_6248,N_6293);
nor U6392 (N_6392,N_6161,N_6260);
nand U6393 (N_6393,N_6183,N_6169);
nand U6394 (N_6394,N_6299,N_6286);
or U6395 (N_6395,N_6151,N_6222);
or U6396 (N_6396,N_6166,N_6237);
or U6397 (N_6397,N_6164,N_6188);
nor U6398 (N_6398,N_6267,N_6175);
nand U6399 (N_6399,N_6172,N_6237);
nor U6400 (N_6400,N_6251,N_6177);
or U6401 (N_6401,N_6240,N_6263);
and U6402 (N_6402,N_6266,N_6166);
nand U6403 (N_6403,N_6160,N_6298);
nor U6404 (N_6404,N_6174,N_6221);
nor U6405 (N_6405,N_6236,N_6222);
nor U6406 (N_6406,N_6275,N_6237);
nor U6407 (N_6407,N_6180,N_6286);
xnor U6408 (N_6408,N_6277,N_6291);
nor U6409 (N_6409,N_6255,N_6205);
nand U6410 (N_6410,N_6258,N_6193);
or U6411 (N_6411,N_6292,N_6241);
or U6412 (N_6412,N_6198,N_6211);
or U6413 (N_6413,N_6293,N_6232);
and U6414 (N_6414,N_6165,N_6238);
nor U6415 (N_6415,N_6167,N_6226);
and U6416 (N_6416,N_6158,N_6232);
or U6417 (N_6417,N_6228,N_6245);
nor U6418 (N_6418,N_6235,N_6184);
nand U6419 (N_6419,N_6289,N_6293);
nand U6420 (N_6420,N_6195,N_6215);
and U6421 (N_6421,N_6182,N_6158);
nand U6422 (N_6422,N_6172,N_6298);
nor U6423 (N_6423,N_6196,N_6194);
xor U6424 (N_6424,N_6185,N_6282);
and U6425 (N_6425,N_6231,N_6272);
and U6426 (N_6426,N_6150,N_6235);
and U6427 (N_6427,N_6153,N_6198);
nand U6428 (N_6428,N_6262,N_6224);
nand U6429 (N_6429,N_6265,N_6177);
nor U6430 (N_6430,N_6167,N_6233);
or U6431 (N_6431,N_6291,N_6157);
nand U6432 (N_6432,N_6164,N_6221);
xnor U6433 (N_6433,N_6170,N_6199);
or U6434 (N_6434,N_6172,N_6151);
nor U6435 (N_6435,N_6289,N_6176);
and U6436 (N_6436,N_6150,N_6274);
and U6437 (N_6437,N_6278,N_6171);
and U6438 (N_6438,N_6259,N_6238);
nor U6439 (N_6439,N_6184,N_6245);
nand U6440 (N_6440,N_6257,N_6150);
and U6441 (N_6441,N_6218,N_6151);
nand U6442 (N_6442,N_6249,N_6248);
xor U6443 (N_6443,N_6168,N_6243);
and U6444 (N_6444,N_6247,N_6274);
or U6445 (N_6445,N_6179,N_6198);
nor U6446 (N_6446,N_6165,N_6159);
nor U6447 (N_6447,N_6294,N_6226);
nor U6448 (N_6448,N_6183,N_6259);
nand U6449 (N_6449,N_6265,N_6224);
xnor U6450 (N_6450,N_6398,N_6319);
and U6451 (N_6451,N_6324,N_6350);
or U6452 (N_6452,N_6368,N_6338);
and U6453 (N_6453,N_6417,N_6373);
nor U6454 (N_6454,N_6366,N_6400);
and U6455 (N_6455,N_6335,N_6408);
nand U6456 (N_6456,N_6401,N_6349);
nor U6457 (N_6457,N_6308,N_6395);
or U6458 (N_6458,N_6418,N_6331);
and U6459 (N_6459,N_6414,N_6363);
nand U6460 (N_6460,N_6353,N_6397);
nand U6461 (N_6461,N_6322,N_6409);
and U6462 (N_6462,N_6329,N_6359);
and U6463 (N_6463,N_6421,N_6358);
or U6464 (N_6464,N_6390,N_6413);
or U6465 (N_6465,N_6383,N_6337);
xnor U6466 (N_6466,N_6436,N_6315);
nand U6467 (N_6467,N_6371,N_6344);
nand U6468 (N_6468,N_6310,N_6374);
or U6469 (N_6469,N_6356,N_6419);
xor U6470 (N_6470,N_6440,N_6424);
or U6471 (N_6471,N_6439,N_6399);
nor U6472 (N_6472,N_6354,N_6303);
and U6473 (N_6473,N_6332,N_6449);
and U6474 (N_6474,N_6300,N_6384);
nand U6475 (N_6475,N_6404,N_6375);
xnor U6476 (N_6476,N_6410,N_6361);
and U6477 (N_6477,N_6427,N_6355);
nand U6478 (N_6478,N_6323,N_6412);
xnor U6479 (N_6479,N_6325,N_6444);
xnor U6480 (N_6480,N_6317,N_6447);
xor U6481 (N_6481,N_6334,N_6362);
and U6482 (N_6482,N_6352,N_6387);
and U6483 (N_6483,N_6316,N_6382);
xor U6484 (N_6484,N_6326,N_6430);
nor U6485 (N_6485,N_6396,N_6336);
xnor U6486 (N_6486,N_6422,N_6441);
nand U6487 (N_6487,N_6340,N_6341);
nand U6488 (N_6488,N_6431,N_6328);
nor U6489 (N_6489,N_6402,N_6381);
or U6490 (N_6490,N_6392,N_6305);
nor U6491 (N_6491,N_6426,N_6394);
or U6492 (N_6492,N_6314,N_6343);
nand U6493 (N_6493,N_6376,N_6347);
nor U6494 (N_6494,N_6360,N_6302);
and U6495 (N_6495,N_6415,N_6367);
xor U6496 (N_6496,N_6434,N_6377);
and U6497 (N_6497,N_6429,N_6407);
nand U6498 (N_6498,N_6345,N_6388);
nor U6499 (N_6499,N_6416,N_6391);
xor U6500 (N_6500,N_6301,N_6357);
or U6501 (N_6501,N_6446,N_6432);
and U6502 (N_6502,N_6420,N_6403);
and U6503 (N_6503,N_6386,N_6342);
and U6504 (N_6504,N_6365,N_6312);
nor U6505 (N_6505,N_6442,N_6306);
or U6506 (N_6506,N_6364,N_6346);
xor U6507 (N_6507,N_6438,N_6313);
nand U6508 (N_6508,N_6372,N_6309);
and U6509 (N_6509,N_6425,N_6369);
nor U6510 (N_6510,N_6443,N_6389);
or U6511 (N_6511,N_6339,N_6318);
nand U6512 (N_6512,N_6320,N_6304);
xnor U6513 (N_6513,N_6437,N_6448);
nor U6514 (N_6514,N_6393,N_6378);
and U6515 (N_6515,N_6406,N_6428);
nand U6516 (N_6516,N_6370,N_6311);
or U6517 (N_6517,N_6385,N_6307);
and U6518 (N_6518,N_6380,N_6433);
or U6519 (N_6519,N_6321,N_6333);
xnor U6520 (N_6520,N_6411,N_6330);
nand U6521 (N_6521,N_6351,N_6423);
and U6522 (N_6522,N_6405,N_6435);
xor U6523 (N_6523,N_6379,N_6445);
xor U6524 (N_6524,N_6348,N_6327);
and U6525 (N_6525,N_6326,N_6423);
nand U6526 (N_6526,N_6349,N_6319);
and U6527 (N_6527,N_6384,N_6333);
xnor U6528 (N_6528,N_6360,N_6330);
nand U6529 (N_6529,N_6411,N_6429);
nor U6530 (N_6530,N_6341,N_6319);
xnor U6531 (N_6531,N_6347,N_6361);
xor U6532 (N_6532,N_6354,N_6329);
or U6533 (N_6533,N_6410,N_6397);
and U6534 (N_6534,N_6347,N_6410);
and U6535 (N_6535,N_6379,N_6356);
nor U6536 (N_6536,N_6398,N_6330);
nor U6537 (N_6537,N_6360,N_6357);
and U6538 (N_6538,N_6365,N_6382);
and U6539 (N_6539,N_6361,N_6345);
xnor U6540 (N_6540,N_6330,N_6447);
and U6541 (N_6541,N_6373,N_6338);
nand U6542 (N_6542,N_6375,N_6374);
or U6543 (N_6543,N_6403,N_6328);
nor U6544 (N_6544,N_6312,N_6301);
nand U6545 (N_6545,N_6391,N_6301);
and U6546 (N_6546,N_6422,N_6310);
nand U6547 (N_6547,N_6331,N_6357);
and U6548 (N_6548,N_6303,N_6315);
xnor U6549 (N_6549,N_6428,N_6421);
xnor U6550 (N_6550,N_6374,N_6307);
and U6551 (N_6551,N_6409,N_6386);
or U6552 (N_6552,N_6336,N_6390);
or U6553 (N_6553,N_6416,N_6448);
nand U6554 (N_6554,N_6333,N_6338);
or U6555 (N_6555,N_6418,N_6374);
nand U6556 (N_6556,N_6391,N_6411);
or U6557 (N_6557,N_6426,N_6397);
nor U6558 (N_6558,N_6427,N_6443);
xor U6559 (N_6559,N_6403,N_6344);
nand U6560 (N_6560,N_6359,N_6423);
nand U6561 (N_6561,N_6353,N_6323);
nor U6562 (N_6562,N_6418,N_6315);
and U6563 (N_6563,N_6415,N_6356);
nand U6564 (N_6564,N_6424,N_6369);
and U6565 (N_6565,N_6408,N_6422);
or U6566 (N_6566,N_6439,N_6403);
and U6567 (N_6567,N_6309,N_6315);
nand U6568 (N_6568,N_6305,N_6345);
xor U6569 (N_6569,N_6317,N_6432);
xnor U6570 (N_6570,N_6433,N_6354);
nand U6571 (N_6571,N_6437,N_6314);
nor U6572 (N_6572,N_6389,N_6393);
and U6573 (N_6573,N_6383,N_6315);
xnor U6574 (N_6574,N_6315,N_6390);
nor U6575 (N_6575,N_6339,N_6400);
nand U6576 (N_6576,N_6361,N_6409);
and U6577 (N_6577,N_6361,N_6421);
nor U6578 (N_6578,N_6334,N_6364);
or U6579 (N_6579,N_6400,N_6300);
nor U6580 (N_6580,N_6313,N_6440);
nand U6581 (N_6581,N_6346,N_6306);
or U6582 (N_6582,N_6421,N_6399);
nor U6583 (N_6583,N_6386,N_6309);
xnor U6584 (N_6584,N_6399,N_6347);
xor U6585 (N_6585,N_6371,N_6445);
and U6586 (N_6586,N_6411,N_6318);
nand U6587 (N_6587,N_6315,N_6347);
nand U6588 (N_6588,N_6389,N_6361);
or U6589 (N_6589,N_6347,N_6448);
nand U6590 (N_6590,N_6400,N_6320);
and U6591 (N_6591,N_6394,N_6445);
xor U6592 (N_6592,N_6440,N_6310);
or U6593 (N_6593,N_6410,N_6305);
nor U6594 (N_6594,N_6317,N_6444);
nor U6595 (N_6595,N_6329,N_6336);
or U6596 (N_6596,N_6372,N_6342);
nand U6597 (N_6597,N_6428,N_6356);
and U6598 (N_6598,N_6351,N_6372);
nand U6599 (N_6599,N_6312,N_6376);
nand U6600 (N_6600,N_6573,N_6451);
or U6601 (N_6601,N_6526,N_6559);
and U6602 (N_6602,N_6547,N_6538);
nor U6603 (N_6603,N_6578,N_6474);
nor U6604 (N_6604,N_6485,N_6531);
nand U6605 (N_6605,N_6576,N_6524);
or U6606 (N_6606,N_6516,N_6472);
nand U6607 (N_6607,N_6490,N_6528);
nand U6608 (N_6608,N_6487,N_6501);
nand U6609 (N_6609,N_6565,N_6536);
or U6610 (N_6610,N_6457,N_6585);
and U6611 (N_6611,N_6458,N_6508);
xor U6612 (N_6612,N_6455,N_6461);
nand U6613 (N_6613,N_6552,N_6479);
and U6614 (N_6614,N_6475,N_6544);
and U6615 (N_6615,N_6583,N_6556);
xnor U6616 (N_6616,N_6555,N_6577);
and U6617 (N_6617,N_6486,N_6465);
or U6618 (N_6618,N_6504,N_6480);
and U6619 (N_6619,N_6594,N_6586);
and U6620 (N_6620,N_6534,N_6581);
or U6621 (N_6621,N_6575,N_6463);
nand U6622 (N_6622,N_6590,N_6499);
xor U6623 (N_6623,N_6533,N_6537);
xor U6624 (N_6624,N_6453,N_6529);
nor U6625 (N_6625,N_6502,N_6493);
xor U6626 (N_6626,N_6469,N_6542);
or U6627 (N_6627,N_6473,N_6492);
or U6628 (N_6628,N_6591,N_6541);
nand U6629 (N_6629,N_6478,N_6553);
nand U6630 (N_6630,N_6456,N_6574);
and U6631 (N_6631,N_6484,N_6539);
nor U6632 (N_6632,N_6584,N_6561);
xor U6633 (N_6633,N_6557,N_6535);
xor U6634 (N_6634,N_6500,N_6572);
or U6635 (N_6635,N_6496,N_6519);
nor U6636 (N_6636,N_6546,N_6599);
xor U6637 (N_6637,N_6580,N_6593);
and U6638 (N_6638,N_6530,N_6568);
or U6639 (N_6639,N_6468,N_6532);
nor U6640 (N_6640,N_6558,N_6505);
xnor U6641 (N_6641,N_6596,N_6554);
and U6642 (N_6642,N_6460,N_6549);
and U6643 (N_6643,N_6507,N_6582);
or U6644 (N_6644,N_6571,N_6452);
and U6645 (N_6645,N_6462,N_6515);
or U6646 (N_6646,N_6522,N_6514);
xor U6647 (N_6647,N_6476,N_6521);
or U6648 (N_6648,N_6471,N_6592);
and U6649 (N_6649,N_6509,N_6564);
nand U6650 (N_6650,N_6567,N_6477);
and U6651 (N_6651,N_6481,N_6454);
nand U6652 (N_6652,N_6488,N_6525);
nor U6653 (N_6653,N_6513,N_6498);
and U6654 (N_6654,N_6598,N_6588);
nor U6655 (N_6655,N_6497,N_6587);
nand U6656 (N_6656,N_6518,N_6520);
xor U6657 (N_6657,N_6569,N_6527);
nand U6658 (N_6658,N_6450,N_6550);
and U6659 (N_6659,N_6510,N_6545);
xor U6660 (N_6660,N_6566,N_6548);
xor U6661 (N_6661,N_6562,N_6595);
or U6662 (N_6662,N_6540,N_6512);
nor U6663 (N_6663,N_6483,N_6489);
or U6664 (N_6664,N_6589,N_6495);
nand U6665 (N_6665,N_6523,N_6503);
and U6666 (N_6666,N_6570,N_6579);
nor U6667 (N_6667,N_6560,N_6543);
nand U6668 (N_6668,N_6517,N_6464);
or U6669 (N_6669,N_6470,N_6551);
nor U6670 (N_6670,N_6494,N_6466);
xnor U6671 (N_6671,N_6459,N_6506);
nor U6672 (N_6672,N_6467,N_6511);
xor U6673 (N_6673,N_6491,N_6482);
xor U6674 (N_6674,N_6597,N_6563);
nand U6675 (N_6675,N_6563,N_6499);
or U6676 (N_6676,N_6576,N_6572);
and U6677 (N_6677,N_6528,N_6474);
nor U6678 (N_6678,N_6560,N_6495);
nor U6679 (N_6679,N_6579,N_6521);
or U6680 (N_6680,N_6562,N_6505);
nand U6681 (N_6681,N_6547,N_6459);
and U6682 (N_6682,N_6453,N_6514);
and U6683 (N_6683,N_6562,N_6454);
and U6684 (N_6684,N_6548,N_6544);
and U6685 (N_6685,N_6470,N_6474);
nor U6686 (N_6686,N_6505,N_6525);
or U6687 (N_6687,N_6506,N_6595);
xnor U6688 (N_6688,N_6576,N_6512);
nor U6689 (N_6689,N_6478,N_6547);
and U6690 (N_6690,N_6462,N_6481);
nor U6691 (N_6691,N_6466,N_6457);
xnor U6692 (N_6692,N_6572,N_6484);
nand U6693 (N_6693,N_6533,N_6584);
nand U6694 (N_6694,N_6579,N_6524);
nor U6695 (N_6695,N_6521,N_6580);
and U6696 (N_6696,N_6490,N_6562);
or U6697 (N_6697,N_6589,N_6538);
or U6698 (N_6698,N_6524,N_6575);
and U6699 (N_6699,N_6513,N_6533);
xor U6700 (N_6700,N_6498,N_6486);
or U6701 (N_6701,N_6540,N_6532);
xor U6702 (N_6702,N_6584,N_6496);
nor U6703 (N_6703,N_6451,N_6566);
nand U6704 (N_6704,N_6508,N_6514);
nor U6705 (N_6705,N_6484,N_6584);
nor U6706 (N_6706,N_6455,N_6572);
nand U6707 (N_6707,N_6582,N_6571);
and U6708 (N_6708,N_6526,N_6471);
or U6709 (N_6709,N_6464,N_6528);
and U6710 (N_6710,N_6496,N_6596);
nor U6711 (N_6711,N_6510,N_6495);
or U6712 (N_6712,N_6490,N_6586);
and U6713 (N_6713,N_6460,N_6565);
or U6714 (N_6714,N_6565,N_6570);
or U6715 (N_6715,N_6554,N_6526);
nor U6716 (N_6716,N_6561,N_6560);
or U6717 (N_6717,N_6483,N_6543);
xnor U6718 (N_6718,N_6589,N_6572);
xor U6719 (N_6719,N_6505,N_6529);
and U6720 (N_6720,N_6550,N_6539);
or U6721 (N_6721,N_6559,N_6560);
or U6722 (N_6722,N_6494,N_6492);
nand U6723 (N_6723,N_6464,N_6454);
xnor U6724 (N_6724,N_6489,N_6491);
and U6725 (N_6725,N_6515,N_6542);
and U6726 (N_6726,N_6588,N_6573);
xnor U6727 (N_6727,N_6500,N_6509);
xor U6728 (N_6728,N_6466,N_6521);
nor U6729 (N_6729,N_6487,N_6477);
or U6730 (N_6730,N_6547,N_6494);
nor U6731 (N_6731,N_6479,N_6543);
or U6732 (N_6732,N_6479,N_6569);
nand U6733 (N_6733,N_6535,N_6516);
xor U6734 (N_6734,N_6465,N_6495);
nor U6735 (N_6735,N_6583,N_6471);
xor U6736 (N_6736,N_6501,N_6457);
and U6737 (N_6737,N_6547,N_6529);
nand U6738 (N_6738,N_6594,N_6574);
nand U6739 (N_6739,N_6522,N_6508);
nor U6740 (N_6740,N_6521,N_6505);
or U6741 (N_6741,N_6451,N_6591);
nand U6742 (N_6742,N_6575,N_6583);
xor U6743 (N_6743,N_6531,N_6520);
nor U6744 (N_6744,N_6516,N_6583);
nor U6745 (N_6745,N_6500,N_6577);
xor U6746 (N_6746,N_6519,N_6582);
nand U6747 (N_6747,N_6572,N_6464);
xnor U6748 (N_6748,N_6518,N_6511);
and U6749 (N_6749,N_6543,N_6490);
and U6750 (N_6750,N_6674,N_6685);
nor U6751 (N_6751,N_6709,N_6657);
or U6752 (N_6752,N_6673,N_6706);
nand U6753 (N_6753,N_6741,N_6737);
and U6754 (N_6754,N_6647,N_6622);
nor U6755 (N_6755,N_6632,N_6693);
or U6756 (N_6756,N_6636,N_6637);
nor U6757 (N_6757,N_6671,N_6700);
xor U6758 (N_6758,N_6601,N_6654);
nand U6759 (N_6759,N_6658,N_6716);
and U6760 (N_6760,N_6627,N_6688);
or U6761 (N_6761,N_6613,N_6666);
nand U6762 (N_6762,N_6603,N_6662);
and U6763 (N_6763,N_6602,N_6672);
and U6764 (N_6764,N_6682,N_6626);
nor U6765 (N_6765,N_6664,N_6677);
nor U6766 (N_6766,N_6661,N_6656);
and U6767 (N_6767,N_6696,N_6634);
nor U6768 (N_6768,N_6701,N_6623);
nor U6769 (N_6769,N_6631,N_6722);
xnor U6770 (N_6770,N_6618,N_6718);
nand U6771 (N_6771,N_6689,N_6625);
and U6772 (N_6772,N_6745,N_6630);
xnor U6773 (N_6773,N_6621,N_6644);
nor U6774 (N_6774,N_6686,N_6619);
nand U6775 (N_6775,N_6740,N_6733);
xor U6776 (N_6776,N_6746,N_6684);
nand U6777 (N_6777,N_6702,N_6600);
xor U6778 (N_6778,N_6663,N_6680);
nand U6779 (N_6779,N_6679,N_6707);
nand U6780 (N_6780,N_6628,N_6669);
or U6781 (N_6781,N_6749,N_6649);
or U6782 (N_6782,N_6641,N_6725);
or U6783 (N_6783,N_6606,N_6727);
nor U6784 (N_6784,N_6608,N_6748);
and U6785 (N_6785,N_6610,N_6726);
xnor U6786 (N_6786,N_6711,N_6744);
xnor U6787 (N_6787,N_6735,N_6692);
nor U6788 (N_6788,N_6670,N_6724);
nand U6789 (N_6789,N_6616,N_6640);
nor U6790 (N_6790,N_6730,N_6650);
or U6791 (N_6791,N_6604,N_6667);
or U6792 (N_6792,N_6660,N_6624);
or U6793 (N_6793,N_6609,N_6714);
and U6794 (N_6794,N_6612,N_6683);
xor U6795 (N_6795,N_6738,N_6678);
or U6796 (N_6796,N_6703,N_6695);
xor U6797 (N_6797,N_6620,N_6708);
xnor U6798 (N_6798,N_6723,N_6747);
nand U6799 (N_6799,N_6742,N_6648);
nand U6800 (N_6800,N_6651,N_6665);
xor U6801 (N_6801,N_6687,N_6638);
nor U6802 (N_6802,N_6643,N_6715);
or U6803 (N_6803,N_6713,N_6633);
xor U6804 (N_6804,N_6614,N_6698);
nand U6805 (N_6805,N_6739,N_6611);
and U6806 (N_6806,N_6699,N_6635);
nand U6807 (N_6807,N_6645,N_6694);
and U6808 (N_6808,N_6655,N_6729);
nor U6809 (N_6809,N_6732,N_6717);
and U6810 (N_6810,N_6642,N_6675);
and U6811 (N_6811,N_6653,N_6736);
nor U6812 (N_6812,N_6728,N_6607);
nor U6813 (N_6813,N_6639,N_6710);
and U6814 (N_6814,N_6719,N_6697);
nor U6815 (N_6815,N_6743,N_6646);
and U6816 (N_6816,N_6731,N_6615);
and U6817 (N_6817,N_6734,N_6720);
xor U6818 (N_6818,N_6712,N_6617);
or U6819 (N_6819,N_6705,N_6629);
and U6820 (N_6820,N_6605,N_6681);
xnor U6821 (N_6821,N_6721,N_6676);
nor U6822 (N_6822,N_6690,N_6659);
nor U6823 (N_6823,N_6704,N_6652);
or U6824 (N_6824,N_6668,N_6691);
nand U6825 (N_6825,N_6610,N_6650);
or U6826 (N_6826,N_6636,N_6616);
nand U6827 (N_6827,N_6602,N_6645);
nor U6828 (N_6828,N_6634,N_6682);
and U6829 (N_6829,N_6608,N_6654);
xnor U6830 (N_6830,N_6679,N_6634);
nor U6831 (N_6831,N_6715,N_6654);
nand U6832 (N_6832,N_6743,N_6710);
xnor U6833 (N_6833,N_6715,N_6613);
nor U6834 (N_6834,N_6718,N_6634);
and U6835 (N_6835,N_6710,N_6708);
nor U6836 (N_6836,N_6638,N_6748);
or U6837 (N_6837,N_6617,N_6685);
xor U6838 (N_6838,N_6729,N_6630);
and U6839 (N_6839,N_6664,N_6743);
nor U6840 (N_6840,N_6680,N_6646);
nand U6841 (N_6841,N_6736,N_6737);
or U6842 (N_6842,N_6701,N_6670);
nand U6843 (N_6843,N_6640,N_6655);
xor U6844 (N_6844,N_6703,N_6713);
and U6845 (N_6845,N_6642,N_6620);
nand U6846 (N_6846,N_6668,N_6649);
nand U6847 (N_6847,N_6627,N_6644);
nand U6848 (N_6848,N_6746,N_6605);
or U6849 (N_6849,N_6715,N_6662);
xnor U6850 (N_6850,N_6625,N_6693);
xor U6851 (N_6851,N_6643,N_6622);
nand U6852 (N_6852,N_6745,N_6640);
or U6853 (N_6853,N_6633,N_6619);
or U6854 (N_6854,N_6696,N_6726);
and U6855 (N_6855,N_6696,N_6692);
or U6856 (N_6856,N_6604,N_6713);
nor U6857 (N_6857,N_6661,N_6667);
or U6858 (N_6858,N_6607,N_6652);
xnor U6859 (N_6859,N_6734,N_6662);
or U6860 (N_6860,N_6610,N_6699);
and U6861 (N_6861,N_6658,N_6724);
and U6862 (N_6862,N_6702,N_6721);
nor U6863 (N_6863,N_6648,N_6612);
nand U6864 (N_6864,N_6626,N_6604);
and U6865 (N_6865,N_6640,N_6671);
and U6866 (N_6866,N_6662,N_6631);
nor U6867 (N_6867,N_6671,N_6706);
nor U6868 (N_6868,N_6728,N_6738);
xnor U6869 (N_6869,N_6643,N_6701);
nand U6870 (N_6870,N_6609,N_6605);
and U6871 (N_6871,N_6627,N_6741);
or U6872 (N_6872,N_6663,N_6716);
or U6873 (N_6873,N_6621,N_6733);
nor U6874 (N_6874,N_6680,N_6631);
nand U6875 (N_6875,N_6607,N_6616);
nor U6876 (N_6876,N_6714,N_6659);
nor U6877 (N_6877,N_6722,N_6699);
and U6878 (N_6878,N_6671,N_6710);
and U6879 (N_6879,N_6645,N_6630);
nor U6880 (N_6880,N_6724,N_6655);
nor U6881 (N_6881,N_6700,N_6668);
or U6882 (N_6882,N_6736,N_6717);
and U6883 (N_6883,N_6655,N_6734);
nand U6884 (N_6884,N_6749,N_6731);
or U6885 (N_6885,N_6614,N_6625);
nor U6886 (N_6886,N_6605,N_6694);
nor U6887 (N_6887,N_6661,N_6703);
and U6888 (N_6888,N_6626,N_6723);
xnor U6889 (N_6889,N_6605,N_6642);
nor U6890 (N_6890,N_6740,N_6679);
and U6891 (N_6891,N_6699,N_6614);
nand U6892 (N_6892,N_6606,N_6671);
xor U6893 (N_6893,N_6683,N_6679);
and U6894 (N_6894,N_6640,N_6666);
nor U6895 (N_6895,N_6691,N_6602);
or U6896 (N_6896,N_6676,N_6727);
nor U6897 (N_6897,N_6692,N_6625);
or U6898 (N_6898,N_6741,N_6666);
or U6899 (N_6899,N_6619,N_6694);
xor U6900 (N_6900,N_6858,N_6873);
and U6901 (N_6901,N_6890,N_6760);
xor U6902 (N_6902,N_6787,N_6762);
nor U6903 (N_6903,N_6816,N_6875);
or U6904 (N_6904,N_6750,N_6857);
xnor U6905 (N_6905,N_6829,N_6870);
nor U6906 (N_6906,N_6791,N_6796);
xnor U6907 (N_6907,N_6758,N_6889);
nor U6908 (N_6908,N_6801,N_6833);
or U6909 (N_6909,N_6754,N_6826);
and U6910 (N_6910,N_6770,N_6761);
nand U6911 (N_6911,N_6877,N_6756);
nand U6912 (N_6912,N_6855,N_6896);
xnor U6913 (N_6913,N_6764,N_6869);
xor U6914 (N_6914,N_6895,N_6794);
xnor U6915 (N_6915,N_6864,N_6848);
or U6916 (N_6916,N_6824,N_6850);
and U6917 (N_6917,N_6798,N_6755);
or U6918 (N_6918,N_6753,N_6835);
xor U6919 (N_6919,N_6795,N_6776);
xnor U6920 (N_6920,N_6840,N_6884);
xor U6921 (N_6921,N_6847,N_6831);
nor U6922 (N_6922,N_6853,N_6821);
and U6923 (N_6923,N_6894,N_6856);
nor U6924 (N_6924,N_6780,N_6839);
nor U6925 (N_6925,N_6888,N_6837);
xnor U6926 (N_6926,N_6867,N_6752);
xor U6927 (N_6927,N_6846,N_6772);
and U6928 (N_6928,N_6767,N_6825);
and U6929 (N_6929,N_6893,N_6879);
nor U6930 (N_6930,N_6782,N_6834);
or U6931 (N_6931,N_6852,N_6865);
nor U6932 (N_6932,N_6818,N_6851);
xor U6933 (N_6933,N_6766,N_6866);
and U6934 (N_6934,N_6786,N_6792);
nand U6935 (N_6935,N_6808,N_6803);
xnor U6936 (N_6936,N_6859,N_6815);
or U6937 (N_6937,N_6775,N_6807);
nor U6938 (N_6938,N_6759,N_6854);
nor U6939 (N_6939,N_6874,N_6830);
xor U6940 (N_6940,N_6823,N_6885);
xor U6941 (N_6941,N_6778,N_6891);
nor U6942 (N_6942,N_6789,N_6810);
xnor U6943 (N_6943,N_6868,N_6842);
nor U6944 (N_6944,N_6876,N_6836);
nand U6945 (N_6945,N_6841,N_6881);
and U6946 (N_6946,N_6799,N_6883);
and U6947 (N_6947,N_6880,N_6899);
nor U6948 (N_6948,N_6763,N_6805);
nand U6949 (N_6949,N_6809,N_6860);
nor U6950 (N_6950,N_6827,N_6800);
or U6951 (N_6951,N_6804,N_6882);
nor U6952 (N_6952,N_6774,N_6765);
and U6953 (N_6953,N_6813,N_6898);
nand U6954 (N_6954,N_6802,N_6783);
xor U6955 (N_6955,N_6781,N_6838);
and U6956 (N_6956,N_6843,N_6822);
and U6957 (N_6957,N_6871,N_6814);
and U6958 (N_6958,N_6806,N_6773);
xnor U6959 (N_6959,N_6768,N_6845);
xor U6960 (N_6960,N_6863,N_6892);
nor U6961 (N_6961,N_6817,N_6819);
or U6962 (N_6962,N_6862,N_6878);
and U6963 (N_6963,N_6887,N_6812);
or U6964 (N_6964,N_6872,N_6757);
nor U6965 (N_6965,N_6820,N_6784);
nand U6966 (N_6966,N_6779,N_6849);
nand U6967 (N_6967,N_6861,N_6797);
nor U6968 (N_6968,N_6751,N_6828);
nor U6969 (N_6969,N_6771,N_6793);
and U6970 (N_6970,N_6832,N_6811);
and U6971 (N_6971,N_6886,N_6777);
nor U6972 (N_6972,N_6769,N_6785);
or U6973 (N_6973,N_6844,N_6788);
and U6974 (N_6974,N_6790,N_6897);
nand U6975 (N_6975,N_6791,N_6763);
or U6976 (N_6976,N_6878,N_6760);
nand U6977 (N_6977,N_6818,N_6810);
and U6978 (N_6978,N_6812,N_6877);
or U6979 (N_6979,N_6803,N_6832);
and U6980 (N_6980,N_6773,N_6775);
or U6981 (N_6981,N_6844,N_6858);
nor U6982 (N_6982,N_6766,N_6829);
nor U6983 (N_6983,N_6826,N_6831);
and U6984 (N_6984,N_6851,N_6889);
and U6985 (N_6985,N_6804,N_6880);
nor U6986 (N_6986,N_6800,N_6768);
nor U6987 (N_6987,N_6751,N_6786);
and U6988 (N_6988,N_6873,N_6834);
or U6989 (N_6989,N_6767,N_6778);
and U6990 (N_6990,N_6899,N_6779);
nand U6991 (N_6991,N_6800,N_6782);
or U6992 (N_6992,N_6893,N_6766);
nand U6993 (N_6993,N_6780,N_6819);
or U6994 (N_6994,N_6773,N_6890);
xor U6995 (N_6995,N_6822,N_6765);
nand U6996 (N_6996,N_6790,N_6751);
xor U6997 (N_6997,N_6805,N_6765);
and U6998 (N_6998,N_6820,N_6891);
nand U6999 (N_6999,N_6858,N_6768);
xnor U7000 (N_7000,N_6855,N_6782);
or U7001 (N_7001,N_6832,N_6796);
nand U7002 (N_7002,N_6777,N_6855);
nand U7003 (N_7003,N_6759,N_6770);
nor U7004 (N_7004,N_6850,N_6851);
or U7005 (N_7005,N_6821,N_6772);
nor U7006 (N_7006,N_6894,N_6789);
nand U7007 (N_7007,N_6833,N_6897);
nand U7008 (N_7008,N_6819,N_6772);
or U7009 (N_7009,N_6830,N_6822);
nor U7010 (N_7010,N_6798,N_6835);
nand U7011 (N_7011,N_6811,N_6827);
or U7012 (N_7012,N_6753,N_6887);
or U7013 (N_7013,N_6875,N_6821);
xor U7014 (N_7014,N_6820,N_6854);
nand U7015 (N_7015,N_6766,N_6896);
and U7016 (N_7016,N_6798,N_6852);
or U7017 (N_7017,N_6814,N_6816);
and U7018 (N_7018,N_6817,N_6771);
nor U7019 (N_7019,N_6771,N_6785);
xnor U7020 (N_7020,N_6861,N_6835);
nand U7021 (N_7021,N_6796,N_6814);
nand U7022 (N_7022,N_6804,N_6836);
or U7023 (N_7023,N_6757,N_6855);
nand U7024 (N_7024,N_6786,N_6868);
nand U7025 (N_7025,N_6815,N_6813);
nor U7026 (N_7026,N_6762,N_6854);
and U7027 (N_7027,N_6877,N_6789);
nor U7028 (N_7028,N_6813,N_6777);
or U7029 (N_7029,N_6876,N_6863);
nor U7030 (N_7030,N_6877,N_6803);
or U7031 (N_7031,N_6899,N_6861);
nor U7032 (N_7032,N_6790,N_6807);
nor U7033 (N_7033,N_6758,N_6772);
nand U7034 (N_7034,N_6751,N_6811);
nand U7035 (N_7035,N_6759,N_6822);
or U7036 (N_7036,N_6860,N_6785);
nand U7037 (N_7037,N_6815,N_6755);
or U7038 (N_7038,N_6753,N_6847);
xnor U7039 (N_7039,N_6781,N_6800);
nor U7040 (N_7040,N_6751,N_6883);
nor U7041 (N_7041,N_6771,N_6797);
nor U7042 (N_7042,N_6878,N_6897);
nand U7043 (N_7043,N_6872,N_6764);
and U7044 (N_7044,N_6766,N_6884);
nand U7045 (N_7045,N_6782,N_6899);
or U7046 (N_7046,N_6831,N_6812);
xor U7047 (N_7047,N_6841,N_6893);
xor U7048 (N_7048,N_6778,N_6836);
xnor U7049 (N_7049,N_6895,N_6758);
nand U7050 (N_7050,N_6980,N_7007);
or U7051 (N_7051,N_6912,N_6931);
xnor U7052 (N_7052,N_6993,N_6932);
or U7053 (N_7053,N_6994,N_7041);
or U7054 (N_7054,N_6973,N_7011);
xnor U7055 (N_7055,N_6940,N_6933);
and U7056 (N_7056,N_6958,N_6904);
nand U7057 (N_7057,N_6984,N_6986);
or U7058 (N_7058,N_7009,N_6996);
nand U7059 (N_7059,N_7037,N_7047);
xnor U7060 (N_7060,N_6938,N_7040);
nand U7061 (N_7061,N_7033,N_6916);
or U7062 (N_7062,N_6967,N_7042);
nand U7063 (N_7063,N_6957,N_6965);
or U7064 (N_7064,N_6928,N_6970);
nand U7065 (N_7065,N_6947,N_6939);
and U7066 (N_7066,N_7016,N_6909);
xor U7067 (N_7067,N_6978,N_7026);
or U7068 (N_7068,N_6926,N_6966);
nor U7069 (N_7069,N_7029,N_6948);
and U7070 (N_7070,N_7013,N_6976);
and U7071 (N_7071,N_6953,N_7038);
nor U7072 (N_7072,N_6989,N_6963);
nand U7073 (N_7073,N_6964,N_6979);
nand U7074 (N_7074,N_6922,N_6919);
nand U7075 (N_7075,N_6988,N_6936);
and U7076 (N_7076,N_6907,N_7021);
xnor U7077 (N_7077,N_6992,N_7005);
xnor U7078 (N_7078,N_6915,N_6937);
xor U7079 (N_7079,N_7049,N_7039);
xnor U7080 (N_7080,N_7008,N_6900);
or U7081 (N_7081,N_7024,N_6962);
nand U7082 (N_7082,N_7001,N_7010);
xor U7083 (N_7083,N_6943,N_6914);
nand U7084 (N_7084,N_7031,N_7002);
xnor U7085 (N_7085,N_6918,N_6910);
or U7086 (N_7086,N_6929,N_7017);
or U7087 (N_7087,N_6969,N_6955);
and U7088 (N_7088,N_6954,N_6960);
nor U7089 (N_7089,N_6906,N_6923);
xor U7090 (N_7090,N_6952,N_6946);
or U7091 (N_7091,N_6944,N_6971);
nor U7092 (N_7092,N_6991,N_7018);
xnor U7093 (N_7093,N_6905,N_7035);
xor U7094 (N_7094,N_7027,N_6968);
and U7095 (N_7095,N_6945,N_6902);
xor U7096 (N_7096,N_6920,N_7003);
nor U7097 (N_7097,N_7020,N_7044);
xnor U7098 (N_7098,N_6942,N_7028);
nor U7099 (N_7099,N_7036,N_7043);
and U7100 (N_7100,N_6998,N_6961);
or U7101 (N_7101,N_6941,N_6924);
nand U7102 (N_7102,N_6927,N_7045);
xnor U7103 (N_7103,N_6950,N_6903);
nor U7104 (N_7104,N_6972,N_6959);
and U7105 (N_7105,N_6983,N_6974);
or U7106 (N_7106,N_6956,N_6951);
nor U7107 (N_7107,N_7048,N_6990);
xnor U7108 (N_7108,N_7012,N_7014);
xnor U7109 (N_7109,N_6913,N_7015);
nand U7110 (N_7110,N_7006,N_7023);
nand U7111 (N_7111,N_6975,N_7034);
or U7112 (N_7112,N_6901,N_6908);
nor U7113 (N_7113,N_7046,N_6921);
nor U7114 (N_7114,N_6949,N_6925);
xnor U7115 (N_7115,N_6982,N_7000);
nand U7116 (N_7116,N_7019,N_7032);
nand U7117 (N_7117,N_6934,N_6995);
nor U7118 (N_7118,N_6911,N_6985);
or U7119 (N_7119,N_7030,N_6917);
nor U7120 (N_7120,N_6935,N_6987);
xnor U7121 (N_7121,N_6999,N_6930);
xor U7122 (N_7122,N_7022,N_6997);
or U7123 (N_7123,N_7004,N_6981);
nor U7124 (N_7124,N_6977,N_7025);
xor U7125 (N_7125,N_6963,N_6926);
nor U7126 (N_7126,N_7004,N_6977);
or U7127 (N_7127,N_6969,N_6945);
nand U7128 (N_7128,N_6957,N_6905);
nor U7129 (N_7129,N_7029,N_7040);
xor U7130 (N_7130,N_6925,N_7030);
or U7131 (N_7131,N_7026,N_6972);
or U7132 (N_7132,N_6958,N_6946);
nand U7133 (N_7133,N_6908,N_7011);
or U7134 (N_7134,N_7019,N_6923);
or U7135 (N_7135,N_6900,N_6988);
or U7136 (N_7136,N_7035,N_7026);
nor U7137 (N_7137,N_7004,N_6931);
nor U7138 (N_7138,N_7049,N_7029);
and U7139 (N_7139,N_7045,N_7018);
or U7140 (N_7140,N_6943,N_7030);
and U7141 (N_7141,N_7014,N_7024);
or U7142 (N_7142,N_6911,N_7036);
and U7143 (N_7143,N_7049,N_6956);
nand U7144 (N_7144,N_6996,N_6972);
or U7145 (N_7145,N_6966,N_7037);
nand U7146 (N_7146,N_6989,N_6940);
nand U7147 (N_7147,N_7043,N_6939);
or U7148 (N_7148,N_7010,N_6962);
or U7149 (N_7149,N_7012,N_7034);
or U7150 (N_7150,N_7029,N_6962);
or U7151 (N_7151,N_7041,N_6983);
nor U7152 (N_7152,N_6968,N_7012);
nor U7153 (N_7153,N_6997,N_7030);
or U7154 (N_7154,N_6900,N_6981);
nand U7155 (N_7155,N_6996,N_6997);
xnor U7156 (N_7156,N_7032,N_6994);
nand U7157 (N_7157,N_6940,N_6949);
and U7158 (N_7158,N_7034,N_6933);
nor U7159 (N_7159,N_6942,N_7008);
nor U7160 (N_7160,N_6967,N_7004);
or U7161 (N_7161,N_6937,N_6903);
and U7162 (N_7162,N_6979,N_6966);
xnor U7163 (N_7163,N_6969,N_7032);
xor U7164 (N_7164,N_6962,N_6907);
and U7165 (N_7165,N_6943,N_6927);
nor U7166 (N_7166,N_7032,N_7046);
nor U7167 (N_7167,N_6989,N_7026);
and U7168 (N_7168,N_6988,N_6980);
nand U7169 (N_7169,N_6926,N_6970);
and U7170 (N_7170,N_6981,N_6934);
and U7171 (N_7171,N_6965,N_7034);
xnor U7172 (N_7172,N_7012,N_7015);
nand U7173 (N_7173,N_6948,N_6959);
nor U7174 (N_7174,N_6997,N_6988);
nor U7175 (N_7175,N_6928,N_7010);
nor U7176 (N_7176,N_6941,N_7004);
nand U7177 (N_7177,N_7038,N_6991);
or U7178 (N_7178,N_6997,N_6962);
and U7179 (N_7179,N_6917,N_6957);
xnor U7180 (N_7180,N_7033,N_6904);
or U7181 (N_7181,N_6911,N_7030);
or U7182 (N_7182,N_6933,N_6997);
and U7183 (N_7183,N_6966,N_6995);
and U7184 (N_7184,N_7003,N_6902);
or U7185 (N_7185,N_6977,N_7040);
nor U7186 (N_7186,N_7041,N_7039);
or U7187 (N_7187,N_6946,N_7043);
or U7188 (N_7188,N_6962,N_6947);
xor U7189 (N_7189,N_6985,N_7042);
nor U7190 (N_7190,N_6977,N_6949);
or U7191 (N_7191,N_6987,N_6951);
nand U7192 (N_7192,N_7030,N_7022);
or U7193 (N_7193,N_6960,N_7035);
nand U7194 (N_7194,N_6910,N_6921);
nor U7195 (N_7195,N_6992,N_7026);
or U7196 (N_7196,N_6943,N_6966);
nor U7197 (N_7197,N_7021,N_7004);
nor U7198 (N_7198,N_6943,N_6991);
xor U7199 (N_7199,N_6913,N_6943);
and U7200 (N_7200,N_7054,N_7146);
and U7201 (N_7201,N_7088,N_7166);
xnor U7202 (N_7202,N_7174,N_7134);
or U7203 (N_7203,N_7190,N_7171);
and U7204 (N_7204,N_7085,N_7197);
and U7205 (N_7205,N_7102,N_7090);
nor U7206 (N_7206,N_7060,N_7176);
nand U7207 (N_7207,N_7184,N_7139);
nand U7208 (N_7208,N_7121,N_7066);
nor U7209 (N_7209,N_7059,N_7109);
and U7210 (N_7210,N_7132,N_7141);
nand U7211 (N_7211,N_7131,N_7079);
nor U7212 (N_7212,N_7160,N_7101);
xnor U7213 (N_7213,N_7147,N_7155);
and U7214 (N_7214,N_7063,N_7145);
nand U7215 (N_7215,N_7072,N_7196);
nand U7216 (N_7216,N_7086,N_7050);
or U7217 (N_7217,N_7157,N_7077);
or U7218 (N_7218,N_7119,N_7181);
and U7219 (N_7219,N_7186,N_7083);
nand U7220 (N_7220,N_7076,N_7152);
or U7221 (N_7221,N_7055,N_7180);
or U7222 (N_7222,N_7053,N_7168);
or U7223 (N_7223,N_7099,N_7082);
or U7224 (N_7224,N_7069,N_7189);
nor U7225 (N_7225,N_7110,N_7100);
xnor U7226 (N_7226,N_7104,N_7092);
or U7227 (N_7227,N_7096,N_7169);
xnor U7228 (N_7228,N_7192,N_7129);
or U7229 (N_7229,N_7095,N_7106);
nor U7230 (N_7230,N_7093,N_7073);
xor U7231 (N_7231,N_7194,N_7162);
or U7232 (N_7232,N_7065,N_7108);
nor U7233 (N_7233,N_7097,N_7051);
xnor U7234 (N_7234,N_7173,N_7105);
nor U7235 (N_7235,N_7136,N_7172);
nor U7236 (N_7236,N_7130,N_7061);
nand U7237 (N_7237,N_7144,N_7124);
nor U7238 (N_7238,N_7058,N_7164);
xor U7239 (N_7239,N_7071,N_7154);
nor U7240 (N_7240,N_7127,N_7133);
and U7241 (N_7241,N_7081,N_7199);
or U7242 (N_7242,N_7089,N_7159);
or U7243 (N_7243,N_7149,N_7087);
and U7244 (N_7244,N_7150,N_7116);
and U7245 (N_7245,N_7178,N_7193);
nand U7246 (N_7246,N_7128,N_7182);
nor U7247 (N_7247,N_7179,N_7153);
or U7248 (N_7248,N_7113,N_7111);
nand U7249 (N_7249,N_7191,N_7122);
or U7250 (N_7250,N_7080,N_7188);
and U7251 (N_7251,N_7167,N_7057);
xor U7252 (N_7252,N_7123,N_7175);
and U7253 (N_7253,N_7177,N_7126);
nor U7254 (N_7254,N_7107,N_7115);
nor U7255 (N_7255,N_7075,N_7135);
nor U7256 (N_7256,N_7185,N_7056);
nand U7257 (N_7257,N_7137,N_7183);
or U7258 (N_7258,N_7163,N_7078);
or U7259 (N_7259,N_7070,N_7195);
or U7260 (N_7260,N_7074,N_7068);
and U7261 (N_7261,N_7112,N_7062);
and U7262 (N_7262,N_7052,N_7158);
and U7263 (N_7263,N_7148,N_7120);
xor U7264 (N_7264,N_7103,N_7143);
nor U7265 (N_7265,N_7067,N_7187);
and U7266 (N_7266,N_7117,N_7198);
or U7267 (N_7267,N_7142,N_7084);
xor U7268 (N_7268,N_7125,N_7091);
nand U7269 (N_7269,N_7118,N_7064);
nor U7270 (N_7270,N_7140,N_7138);
nand U7271 (N_7271,N_7094,N_7114);
xnor U7272 (N_7272,N_7165,N_7156);
and U7273 (N_7273,N_7170,N_7151);
and U7274 (N_7274,N_7098,N_7161);
or U7275 (N_7275,N_7176,N_7166);
nor U7276 (N_7276,N_7119,N_7198);
nand U7277 (N_7277,N_7093,N_7107);
nor U7278 (N_7278,N_7197,N_7182);
nand U7279 (N_7279,N_7105,N_7157);
nor U7280 (N_7280,N_7051,N_7123);
nor U7281 (N_7281,N_7167,N_7111);
nand U7282 (N_7282,N_7108,N_7162);
nor U7283 (N_7283,N_7158,N_7126);
xnor U7284 (N_7284,N_7128,N_7198);
or U7285 (N_7285,N_7102,N_7094);
nor U7286 (N_7286,N_7059,N_7072);
xnor U7287 (N_7287,N_7069,N_7181);
and U7288 (N_7288,N_7131,N_7143);
or U7289 (N_7289,N_7185,N_7098);
or U7290 (N_7290,N_7155,N_7174);
xor U7291 (N_7291,N_7101,N_7187);
and U7292 (N_7292,N_7179,N_7131);
nor U7293 (N_7293,N_7132,N_7053);
nand U7294 (N_7294,N_7161,N_7155);
nand U7295 (N_7295,N_7136,N_7190);
nor U7296 (N_7296,N_7170,N_7123);
nor U7297 (N_7297,N_7054,N_7073);
or U7298 (N_7298,N_7060,N_7076);
nor U7299 (N_7299,N_7149,N_7055);
nor U7300 (N_7300,N_7057,N_7148);
or U7301 (N_7301,N_7131,N_7177);
xor U7302 (N_7302,N_7168,N_7091);
xnor U7303 (N_7303,N_7160,N_7083);
or U7304 (N_7304,N_7192,N_7156);
xor U7305 (N_7305,N_7177,N_7173);
and U7306 (N_7306,N_7124,N_7166);
or U7307 (N_7307,N_7079,N_7069);
nand U7308 (N_7308,N_7139,N_7187);
or U7309 (N_7309,N_7116,N_7054);
xor U7310 (N_7310,N_7145,N_7180);
or U7311 (N_7311,N_7073,N_7156);
and U7312 (N_7312,N_7106,N_7069);
xor U7313 (N_7313,N_7097,N_7118);
and U7314 (N_7314,N_7088,N_7171);
xor U7315 (N_7315,N_7186,N_7095);
or U7316 (N_7316,N_7110,N_7133);
xor U7317 (N_7317,N_7168,N_7180);
xnor U7318 (N_7318,N_7157,N_7162);
or U7319 (N_7319,N_7070,N_7191);
or U7320 (N_7320,N_7118,N_7071);
and U7321 (N_7321,N_7110,N_7072);
xnor U7322 (N_7322,N_7084,N_7195);
or U7323 (N_7323,N_7105,N_7136);
xnor U7324 (N_7324,N_7121,N_7105);
or U7325 (N_7325,N_7142,N_7098);
nand U7326 (N_7326,N_7162,N_7077);
or U7327 (N_7327,N_7130,N_7172);
or U7328 (N_7328,N_7101,N_7054);
or U7329 (N_7329,N_7054,N_7189);
nor U7330 (N_7330,N_7135,N_7177);
or U7331 (N_7331,N_7160,N_7081);
and U7332 (N_7332,N_7098,N_7183);
and U7333 (N_7333,N_7175,N_7171);
xnor U7334 (N_7334,N_7194,N_7115);
or U7335 (N_7335,N_7081,N_7100);
or U7336 (N_7336,N_7079,N_7138);
nand U7337 (N_7337,N_7131,N_7096);
and U7338 (N_7338,N_7169,N_7191);
nand U7339 (N_7339,N_7111,N_7180);
or U7340 (N_7340,N_7050,N_7154);
nand U7341 (N_7341,N_7166,N_7115);
and U7342 (N_7342,N_7053,N_7054);
or U7343 (N_7343,N_7108,N_7086);
nand U7344 (N_7344,N_7101,N_7064);
nand U7345 (N_7345,N_7189,N_7085);
nand U7346 (N_7346,N_7094,N_7171);
xor U7347 (N_7347,N_7136,N_7184);
nand U7348 (N_7348,N_7114,N_7189);
nor U7349 (N_7349,N_7181,N_7122);
and U7350 (N_7350,N_7276,N_7230);
and U7351 (N_7351,N_7292,N_7326);
nand U7352 (N_7352,N_7320,N_7226);
nand U7353 (N_7353,N_7234,N_7330);
nand U7354 (N_7354,N_7344,N_7281);
and U7355 (N_7355,N_7218,N_7256);
and U7356 (N_7356,N_7268,N_7346);
nand U7357 (N_7357,N_7274,N_7202);
and U7358 (N_7358,N_7242,N_7291);
or U7359 (N_7359,N_7325,N_7200);
nor U7360 (N_7360,N_7251,N_7259);
or U7361 (N_7361,N_7209,N_7253);
or U7362 (N_7362,N_7214,N_7252);
and U7363 (N_7363,N_7248,N_7269);
nor U7364 (N_7364,N_7337,N_7254);
nand U7365 (N_7365,N_7342,N_7316);
nand U7366 (N_7366,N_7213,N_7308);
or U7367 (N_7367,N_7302,N_7310);
nand U7368 (N_7368,N_7287,N_7227);
and U7369 (N_7369,N_7279,N_7306);
or U7370 (N_7370,N_7266,N_7289);
nand U7371 (N_7371,N_7272,N_7241);
nand U7372 (N_7372,N_7283,N_7347);
nor U7373 (N_7373,N_7317,N_7305);
nand U7374 (N_7374,N_7312,N_7225);
and U7375 (N_7375,N_7212,N_7270);
nor U7376 (N_7376,N_7282,N_7294);
nand U7377 (N_7377,N_7300,N_7247);
or U7378 (N_7378,N_7329,N_7298);
nor U7379 (N_7379,N_7203,N_7206);
and U7380 (N_7380,N_7246,N_7334);
or U7381 (N_7381,N_7275,N_7339);
nor U7382 (N_7382,N_7273,N_7290);
nand U7383 (N_7383,N_7219,N_7249);
nor U7384 (N_7384,N_7299,N_7315);
or U7385 (N_7385,N_7224,N_7208);
or U7386 (N_7386,N_7245,N_7221);
and U7387 (N_7387,N_7336,N_7265);
and U7388 (N_7388,N_7324,N_7288);
nor U7389 (N_7389,N_7318,N_7328);
or U7390 (N_7390,N_7237,N_7223);
or U7391 (N_7391,N_7240,N_7255);
nor U7392 (N_7392,N_7228,N_7232);
nor U7393 (N_7393,N_7211,N_7301);
nand U7394 (N_7394,N_7201,N_7321);
or U7395 (N_7395,N_7271,N_7322);
nor U7396 (N_7396,N_7331,N_7338);
xnor U7397 (N_7397,N_7229,N_7348);
nor U7398 (N_7398,N_7296,N_7238);
xnor U7399 (N_7399,N_7319,N_7231);
nand U7400 (N_7400,N_7235,N_7314);
and U7401 (N_7401,N_7327,N_7343);
and U7402 (N_7402,N_7204,N_7280);
or U7403 (N_7403,N_7335,N_7278);
and U7404 (N_7404,N_7216,N_7333);
and U7405 (N_7405,N_7293,N_7332);
nand U7406 (N_7406,N_7262,N_7297);
nand U7407 (N_7407,N_7250,N_7267);
or U7408 (N_7408,N_7263,N_7261);
or U7409 (N_7409,N_7341,N_7349);
xnor U7410 (N_7410,N_7222,N_7236);
nand U7411 (N_7411,N_7284,N_7233);
and U7412 (N_7412,N_7309,N_7264);
and U7413 (N_7413,N_7285,N_7295);
and U7414 (N_7414,N_7244,N_7311);
and U7415 (N_7415,N_7258,N_7303);
or U7416 (N_7416,N_7307,N_7260);
xor U7417 (N_7417,N_7207,N_7277);
nor U7418 (N_7418,N_7304,N_7205);
nor U7419 (N_7419,N_7210,N_7345);
nand U7420 (N_7420,N_7323,N_7239);
or U7421 (N_7421,N_7217,N_7286);
nand U7422 (N_7422,N_7215,N_7257);
or U7423 (N_7423,N_7313,N_7243);
or U7424 (N_7424,N_7220,N_7340);
nand U7425 (N_7425,N_7264,N_7325);
and U7426 (N_7426,N_7290,N_7318);
nand U7427 (N_7427,N_7246,N_7305);
or U7428 (N_7428,N_7202,N_7221);
xor U7429 (N_7429,N_7324,N_7211);
xor U7430 (N_7430,N_7205,N_7329);
xnor U7431 (N_7431,N_7266,N_7252);
nand U7432 (N_7432,N_7317,N_7345);
xnor U7433 (N_7433,N_7209,N_7283);
xnor U7434 (N_7434,N_7347,N_7241);
xor U7435 (N_7435,N_7267,N_7292);
and U7436 (N_7436,N_7292,N_7320);
nand U7437 (N_7437,N_7212,N_7268);
nor U7438 (N_7438,N_7257,N_7337);
or U7439 (N_7439,N_7264,N_7280);
xnor U7440 (N_7440,N_7282,N_7228);
nor U7441 (N_7441,N_7322,N_7331);
nor U7442 (N_7442,N_7274,N_7233);
nand U7443 (N_7443,N_7329,N_7273);
xor U7444 (N_7444,N_7256,N_7323);
nor U7445 (N_7445,N_7243,N_7348);
nor U7446 (N_7446,N_7301,N_7244);
xor U7447 (N_7447,N_7314,N_7248);
nor U7448 (N_7448,N_7330,N_7343);
nor U7449 (N_7449,N_7326,N_7231);
nand U7450 (N_7450,N_7322,N_7344);
or U7451 (N_7451,N_7201,N_7262);
xnor U7452 (N_7452,N_7226,N_7323);
or U7453 (N_7453,N_7319,N_7323);
or U7454 (N_7454,N_7262,N_7214);
nand U7455 (N_7455,N_7300,N_7243);
or U7456 (N_7456,N_7212,N_7234);
xor U7457 (N_7457,N_7209,N_7340);
xor U7458 (N_7458,N_7208,N_7269);
nand U7459 (N_7459,N_7298,N_7238);
or U7460 (N_7460,N_7295,N_7323);
xnor U7461 (N_7461,N_7229,N_7238);
or U7462 (N_7462,N_7312,N_7298);
nand U7463 (N_7463,N_7308,N_7219);
xnor U7464 (N_7464,N_7223,N_7242);
or U7465 (N_7465,N_7245,N_7268);
nand U7466 (N_7466,N_7311,N_7234);
and U7467 (N_7467,N_7270,N_7316);
nor U7468 (N_7468,N_7222,N_7336);
or U7469 (N_7469,N_7304,N_7298);
xnor U7470 (N_7470,N_7275,N_7298);
or U7471 (N_7471,N_7214,N_7345);
nor U7472 (N_7472,N_7234,N_7283);
or U7473 (N_7473,N_7306,N_7281);
nand U7474 (N_7474,N_7217,N_7253);
and U7475 (N_7475,N_7289,N_7227);
nor U7476 (N_7476,N_7318,N_7235);
and U7477 (N_7477,N_7260,N_7319);
xor U7478 (N_7478,N_7316,N_7264);
xnor U7479 (N_7479,N_7264,N_7317);
nand U7480 (N_7480,N_7242,N_7273);
and U7481 (N_7481,N_7314,N_7303);
nand U7482 (N_7482,N_7321,N_7226);
xnor U7483 (N_7483,N_7269,N_7250);
nor U7484 (N_7484,N_7228,N_7316);
nand U7485 (N_7485,N_7259,N_7341);
and U7486 (N_7486,N_7261,N_7231);
xor U7487 (N_7487,N_7293,N_7229);
xnor U7488 (N_7488,N_7272,N_7233);
or U7489 (N_7489,N_7227,N_7214);
or U7490 (N_7490,N_7212,N_7251);
nor U7491 (N_7491,N_7349,N_7301);
nand U7492 (N_7492,N_7238,N_7308);
and U7493 (N_7493,N_7225,N_7221);
and U7494 (N_7494,N_7207,N_7253);
and U7495 (N_7495,N_7245,N_7311);
nand U7496 (N_7496,N_7256,N_7219);
or U7497 (N_7497,N_7340,N_7324);
xor U7498 (N_7498,N_7332,N_7264);
or U7499 (N_7499,N_7338,N_7336);
nand U7500 (N_7500,N_7423,N_7355);
xor U7501 (N_7501,N_7409,N_7419);
nor U7502 (N_7502,N_7424,N_7410);
xnor U7503 (N_7503,N_7405,N_7493);
xor U7504 (N_7504,N_7356,N_7458);
nor U7505 (N_7505,N_7432,N_7364);
nor U7506 (N_7506,N_7380,N_7495);
or U7507 (N_7507,N_7441,N_7459);
or U7508 (N_7508,N_7491,N_7487);
xor U7509 (N_7509,N_7494,N_7442);
or U7510 (N_7510,N_7427,N_7414);
nand U7511 (N_7511,N_7381,N_7430);
and U7512 (N_7512,N_7499,N_7476);
nand U7513 (N_7513,N_7383,N_7351);
nor U7514 (N_7514,N_7376,N_7392);
nand U7515 (N_7515,N_7363,N_7452);
or U7516 (N_7516,N_7471,N_7375);
and U7517 (N_7517,N_7426,N_7420);
nand U7518 (N_7518,N_7475,N_7418);
nor U7519 (N_7519,N_7443,N_7438);
or U7520 (N_7520,N_7439,N_7388);
and U7521 (N_7521,N_7367,N_7454);
and U7522 (N_7522,N_7444,N_7455);
or U7523 (N_7523,N_7398,N_7449);
nor U7524 (N_7524,N_7384,N_7387);
nand U7525 (N_7525,N_7389,N_7372);
xnor U7526 (N_7526,N_7377,N_7433);
xor U7527 (N_7527,N_7357,N_7391);
nand U7528 (N_7528,N_7353,N_7369);
and U7529 (N_7529,N_7378,N_7415);
and U7530 (N_7530,N_7373,N_7404);
and U7531 (N_7531,N_7397,N_7436);
nor U7532 (N_7532,N_7362,N_7462);
and U7533 (N_7533,N_7411,N_7457);
xor U7534 (N_7534,N_7401,N_7370);
nor U7535 (N_7535,N_7498,N_7456);
or U7536 (N_7536,N_7407,N_7483);
nor U7537 (N_7537,N_7406,N_7361);
xnor U7538 (N_7538,N_7421,N_7359);
xor U7539 (N_7539,N_7393,N_7431);
and U7540 (N_7540,N_7402,N_7446);
or U7541 (N_7541,N_7451,N_7408);
and U7542 (N_7542,N_7394,N_7396);
nand U7543 (N_7543,N_7467,N_7360);
nor U7544 (N_7544,N_7478,N_7497);
and U7545 (N_7545,N_7482,N_7486);
nand U7546 (N_7546,N_7435,N_7358);
and U7547 (N_7547,N_7465,N_7385);
and U7548 (N_7548,N_7400,N_7447);
and U7549 (N_7549,N_7490,N_7479);
xnor U7550 (N_7550,N_7464,N_7468);
nor U7551 (N_7551,N_7445,N_7469);
nor U7552 (N_7552,N_7417,N_7382);
nor U7553 (N_7553,N_7488,N_7480);
xnor U7554 (N_7554,N_7473,N_7448);
nor U7555 (N_7555,N_7428,N_7354);
nand U7556 (N_7556,N_7350,N_7496);
and U7557 (N_7557,N_7365,N_7463);
xnor U7558 (N_7558,N_7472,N_7395);
xor U7559 (N_7559,N_7485,N_7470);
nand U7560 (N_7560,N_7450,N_7390);
and U7561 (N_7561,N_7440,N_7412);
xor U7562 (N_7562,N_7489,N_7481);
or U7563 (N_7563,N_7399,N_7422);
or U7564 (N_7564,N_7379,N_7477);
nor U7565 (N_7565,N_7466,N_7374);
and U7566 (N_7566,N_7492,N_7461);
or U7567 (N_7567,N_7413,N_7386);
or U7568 (N_7568,N_7474,N_7403);
xor U7569 (N_7569,N_7429,N_7453);
or U7570 (N_7570,N_7484,N_7460);
and U7571 (N_7571,N_7437,N_7352);
or U7572 (N_7572,N_7368,N_7425);
xor U7573 (N_7573,N_7434,N_7416);
xnor U7574 (N_7574,N_7366,N_7371);
xnor U7575 (N_7575,N_7432,N_7433);
or U7576 (N_7576,N_7452,N_7422);
or U7577 (N_7577,N_7399,N_7388);
or U7578 (N_7578,N_7422,N_7448);
and U7579 (N_7579,N_7439,N_7459);
and U7580 (N_7580,N_7364,N_7405);
or U7581 (N_7581,N_7422,N_7386);
and U7582 (N_7582,N_7487,N_7395);
nand U7583 (N_7583,N_7458,N_7456);
or U7584 (N_7584,N_7483,N_7403);
xor U7585 (N_7585,N_7382,N_7432);
or U7586 (N_7586,N_7401,N_7447);
or U7587 (N_7587,N_7469,N_7434);
and U7588 (N_7588,N_7452,N_7353);
or U7589 (N_7589,N_7352,N_7442);
xnor U7590 (N_7590,N_7401,N_7475);
or U7591 (N_7591,N_7419,N_7415);
and U7592 (N_7592,N_7360,N_7494);
nand U7593 (N_7593,N_7374,N_7400);
nor U7594 (N_7594,N_7384,N_7477);
and U7595 (N_7595,N_7427,N_7410);
and U7596 (N_7596,N_7403,N_7424);
nor U7597 (N_7597,N_7383,N_7453);
or U7598 (N_7598,N_7409,N_7438);
nor U7599 (N_7599,N_7449,N_7473);
nor U7600 (N_7600,N_7401,N_7405);
and U7601 (N_7601,N_7426,N_7485);
and U7602 (N_7602,N_7443,N_7363);
nor U7603 (N_7603,N_7470,N_7373);
nand U7604 (N_7604,N_7353,N_7386);
xor U7605 (N_7605,N_7453,N_7387);
nor U7606 (N_7606,N_7352,N_7372);
nand U7607 (N_7607,N_7424,N_7385);
xor U7608 (N_7608,N_7437,N_7472);
or U7609 (N_7609,N_7380,N_7371);
nand U7610 (N_7610,N_7488,N_7472);
or U7611 (N_7611,N_7480,N_7427);
and U7612 (N_7612,N_7447,N_7410);
or U7613 (N_7613,N_7376,N_7403);
xnor U7614 (N_7614,N_7418,N_7451);
nor U7615 (N_7615,N_7367,N_7352);
and U7616 (N_7616,N_7404,N_7490);
xor U7617 (N_7617,N_7444,N_7364);
and U7618 (N_7618,N_7394,N_7492);
xor U7619 (N_7619,N_7358,N_7422);
or U7620 (N_7620,N_7399,N_7468);
nor U7621 (N_7621,N_7379,N_7479);
xnor U7622 (N_7622,N_7368,N_7376);
nor U7623 (N_7623,N_7473,N_7392);
and U7624 (N_7624,N_7410,N_7442);
nand U7625 (N_7625,N_7373,N_7401);
nor U7626 (N_7626,N_7371,N_7496);
nor U7627 (N_7627,N_7459,N_7447);
nor U7628 (N_7628,N_7371,N_7447);
or U7629 (N_7629,N_7355,N_7457);
nand U7630 (N_7630,N_7440,N_7415);
xor U7631 (N_7631,N_7472,N_7379);
nand U7632 (N_7632,N_7476,N_7437);
nor U7633 (N_7633,N_7472,N_7430);
nand U7634 (N_7634,N_7478,N_7377);
nand U7635 (N_7635,N_7383,N_7378);
nand U7636 (N_7636,N_7488,N_7458);
and U7637 (N_7637,N_7392,N_7440);
nand U7638 (N_7638,N_7446,N_7470);
xnor U7639 (N_7639,N_7405,N_7425);
nor U7640 (N_7640,N_7396,N_7413);
xor U7641 (N_7641,N_7491,N_7471);
nand U7642 (N_7642,N_7479,N_7491);
and U7643 (N_7643,N_7490,N_7499);
nor U7644 (N_7644,N_7367,N_7483);
and U7645 (N_7645,N_7414,N_7438);
and U7646 (N_7646,N_7397,N_7389);
or U7647 (N_7647,N_7411,N_7440);
and U7648 (N_7648,N_7454,N_7399);
nor U7649 (N_7649,N_7399,N_7413);
and U7650 (N_7650,N_7517,N_7645);
nor U7651 (N_7651,N_7640,N_7647);
nor U7652 (N_7652,N_7613,N_7624);
nor U7653 (N_7653,N_7593,N_7579);
xor U7654 (N_7654,N_7556,N_7509);
and U7655 (N_7655,N_7564,N_7574);
nor U7656 (N_7656,N_7614,N_7559);
nor U7657 (N_7657,N_7534,N_7523);
or U7658 (N_7658,N_7605,N_7529);
nor U7659 (N_7659,N_7589,N_7567);
xnor U7660 (N_7660,N_7618,N_7586);
xnor U7661 (N_7661,N_7508,N_7615);
xnor U7662 (N_7662,N_7583,N_7533);
xor U7663 (N_7663,N_7638,N_7535);
nor U7664 (N_7664,N_7643,N_7541);
nand U7665 (N_7665,N_7538,N_7561);
or U7666 (N_7666,N_7565,N_7552);
nor U7667 (N_7667,N_7555,N_7536);
or U7668 (N_7668,N_7609,N_7560);
xnor U7669 (N_7669,N_7633,N_7620);
nor U7670 (N_7670,N_7627,N_7596);
or U7671 (N_7671,N_7641,N_7521);
and U7672 (N_7672,N_7500,N_7634);
xnor U7673 (N_7673,N_7557,N_7577);
nor U7674 (N_7674,N_7527,N_7522);
xor U7675 (N_7675,N_7612,N_7606);
nand U7676 (N_7676,N_7562,N_7602);
and U7677 (N_7677,N_7591,N_7511);
nor U7678 (N_7678,N_7642,N_7506);
and U7679 (N_7679,N_7520,N_7510);
and U7680 (N_7680,N_7531,N_7553);
nor U7681 (N_7681,N_7543,N_7570);
and U7682 (N_7682,N_7537,N_7649);
xor U7683 (N_7683,N_7549,N_7547);
nor U7684 (N_7684,N_7544,N_7554);
xnor U7685 (N_7685,N_7550,N_7611);
nand U7686 (N_7686,N_7571,N_7578);
nor U7687 (N_7687,N_7617,N_7558);
nor U7688 (N_7688,N_7539,N_7646);
nand U7689 (N_7689,N_7639,N_7588);
nand U7690 (N_7690,N_7505,N_7607);
and U7691 (N_7691,N_7501,N_7623);
xor U7692 (N_7692,N_7525,N_7604);
xnor U7693 (N_7693,N_7528,N_7626);
nand U7694 (N_7694,N_7518,N_7568);
and U7695 (N_7695,N_7519,N_7622);
and U7696 (N_7696,N_7530,N_7594);
and U7697 (N_7697,N_7542,N_7636);
nor U7698 (N_7698,N_7630,N_7619);
nor U7699 (N_7699,N_7503,N_7603);
xnor U7700 (N_7700,N_7540,N_7601);
nand U7701 (N_7701,N_7644,N_7637);
nor U7702 (N_7702,N_7631,N_7616);
nand U7703 (N_7703,N_7526,N_7580);
and U7704 (N_7704,N_7648,N_7581);
and U7705 (N_7705,N_7507,N_7572);
nand U7706 (N_7706,N_7610,N_7576);
or U7707 (N_7707,N_7582,N_7516);
and U7708 (N_7708,N_7629,N_7546);
nand U7709 (N_7709,N_7597,N_7595);
or U7710 (N_7710,N_7575,N_7628);
and U7711 (N_7711,N_7608,N_7532);
or U7712 (N_7712,N_7504,N_7632);
or U7713 (N_7713,N_7598,N_7524);
xor U7714 (N_7714,N_7621,N_7551);
xor U7715 (N_7715,N_7569,N_7548);
or U7716 (N_7716,N_7566,N_7599);
and U7717 (N_7717,N_7635,N_7600);
or U7718 (N_7718,N_7592,N_7563);
nor U7719 (N_7719,N_7585,N_7584);
and U7720 (N_7720,N_7514,N_7587);
or U7721 (N_7721,N_7512,N_7590);
xnor U7722 (N_7722,N_7545,N_7573);
and U7723 (N_7723,N_7625,N_7502);
nor U7724 (N_7724,N_7513,N_7515);
nor U7725 (N_7725,N_7641,N_7626);
nand U7726 (N_7726,N_7574,N_7588);
nand U7727 (N_7727,N_7597,N_7541);
or U7728 (N_7728,N_7621,N_7556);
or U7729 (N_7729,N_7559,N_7513);
and U7730 (N_7730,N_7504,N_7594);
and U7731 (N_7731,N_7607,N_7638);
and U7732 (N_7732,N_7510,N_7544);
xnor U7733 (N_7733,N_7644,N_7580);
xor U7734 (N_7734,N_7593,N_7538);
or U7735 (N_7735,N_7550,N_7591);
nand U7736 (N_7736,N_7503,N_7531);
and U7737 (N_7737,N_7524,N_7622);
xor U7738 (N_7738,N_7574,N_7560);
or U7739 (N_7739,N_7544,N_7619);
nor U7740 (N_7740,N_7527,N_7520);
xor U7741 (N_7741,N_7573,N_7504);
nand U7742 (N_7742,N_7517,N_7597);
or U7743 (N_7743,N_7570,N_7646);
and U7744 (N_7744,N_7518,N_7537);
xor U7745 (N_7745,N_7513,N_7610);
nand U7746 (N_7746,N_7628,N_7604);
nor U7747 (N_7747,N_7649,N_7548);
xor U7748 (N_7748,N_7584,N_7601);
nand U7749 (N_7749,N_7627,N_7548);
nor U7750 (N_7750,N_7607,N_7572);
xor U7751 (N_7751,N_7526,N_7643);
nand U7752 (N_7752,N_7501,N_7581);
or U7753 (N_7753,N_7602,N_7581);
or U7754 (N_7754,N_7581,N_7517);
and U7755 (N_7755,N_7503,N_7572);
nor U7756 (N_7756,N_7595,N_7591);
or U7757 (N_7757,N_7516,N_7601);
and U7758 (N_7758,N_7512,N_7534);
nand U7759 (N_7759,N_7594,N_7593);
or U7760 (N_7760,N_7530,N_7524);
xor U7761 (N_7761,N_7577,N_7527);
nand U7762 (N_7762,N_7573,N_7523);
or U7763 (N_7763,N_7524,N_7502);
xnor U7764 (N_7764,N_7607,N_7536);
xnor U7765 (N_7765,N_7616,N_7563);
xnor U7766 (N_7766,N_7516,N_7564);
or U7767 (N_7767,N_7604,N_7527);
xnor U7768 (N_7768,N_7509,N_7527);
nor U7769 (N_7769,N_7576,N_7589);
nand U7770 (N_7770,N_7540,N_7565);
nor U7771 (N_7771,N_7620,N_7548);
and U7772 (N_7772,N_7580,N_7605);
nand U7773 (N_7773,N_7507,N_7607);
nand U7774 (N_7774,N_7639,N_7594);
or U7775 (N_7775,N_7582,N_7615);
xor U7776 (N_7776,N_7544,N_7519);
xnor U7777 (N_7777,N_7646,N_7648);
and U7778 (N_7778,N_7607,N_7568);
or U7779 (N_7779,N_7519,N_7531);
nor U7780 (N_7780,N_7515,N_7616);
nor U7781 (N_7781,N_7584,N_7605);
nand U7782 (N_7782,N_7608,N_7627);
nor U7783 (N_7783,N_7580,N_7624);
or U7784 (N_7784,N_7510,N_7576);
or U7785 (N_7785,N_7642,N_7529);
and U7786 (N_7786,N_7589,N_7522);
or U7787 (N_7787,N_7558,N_7536);
and U7788 (N_7788,N_7500,N_7604);
nand U7789 (N_7789,N_7640,N_7643);
and U7790 (N_7790,N_7612,N_7523);
and U7791 (N_7791,N_7624,N_7644);
nor U7792 (N_7792,N_7618,N_7510);
xor U7793 (N_7793,N_7541,N_7501);
nor U7794 (N_7794,N_7549,N_7556);
nand U7795 (N_7795,N_7572,N_7512);
xnor U7796 (N_7796,N_7612,N_7546);
and U7797 (N_7797,N_7633,N_7563);
nand U7798 (N_7798,N_7638,N_7512);
nand U7799 (N_7799,N_7601,N_7520);
xor U7800 (N_7800,N_7658,N_7756);
nand U7801 (N_7801,N_7674,N_7741);
nand U7802 (N_7802,N_7737,N_7773);
nand U7803 (N_7803,N_7766,N_7664);
or U7804 (N_7804,N_7725,N_7769);
nand U7805 (N_7805,N_7679,N_7764);
and U7806 (N_7806,N_7767,N_7788);
nand U7807 (N_7807,N_7673,N_7666);
xor U7808 (N_7808,N_7786,N_7738);
nor U7809 (N_7809,N_7789,N_7659);
nand U7810 (N_7810,N_7670,N_7746);
nor U7811 (N_7811,N_7677,N_7742);
or U7812 (N_7812,N_7791,N_7689);
and U7813 (N_7813,N_7694,N_7703);
or U7814 (N_7814,N_7716,N_7693);
nand U7815 (N_7815,N_7721,N_7794);
or U7816 (N_7816,N_7713,N_7663);
or U7817 (N_7817,N_7672,N_7757);
nand U7818 (N_7818,N_7692,N_7739);
nor U7819 (N_7819,N_7701,N_7686);
nor U7820 (N_7820,N_7730,N_7775);
nor U7821 (N_7821,N_7743,N_7657);
xnor U7822 (N_7822,N_7785,N_7710);
nand U7823 (N_7823,N_7750,N_7724);
nor U7824 (N_7824,N_7774,N_7690);
nor U7825 (N_7825,N_7798,N_7723);
xnor U7826 (N_7826,N_7697,N_7676);
nand U7827 (N_7827,N_7667,N_7688);
and U7828 (N_7828,N_7772,N_7700);
and U7829 (N_7829,N_7790,N_7782);
and U7830 (N_7830,N_7732,N_7762);
xnor U7831 (N_7831,N_7660,N_7675);
nand U7832 (N_7832,N_7662,N_7656);
and U7833 (N_7833,N_7705,N_7678);
and U7834 (N_7834,N_7708,N_7793);
nand U7835 (N_7835,N_7755,N_7749);
and U7836 (N_7836,N_7685,N_7681);
and U7837 (N_7837,N_7714,N_7780);
or U7838 (N_7838,N_7735,N_7748);
nand U7839 (N_7839,N_7744,N_7728);
nand U7840 (N_7840,N_7650,N_7654);
and U7841 (N_7841,N_7759,N_7751);
xnor U7842 (N_7842,N_7792,N_7661);
or U7843 (N_7843,N_7696,N_7695);
or U7844 (N_7844,N_7731,N_7795);
nand U7845 (N_7845,N_7655,N_7722);
xnor U7846 (N_7846,N_7758,N_7719);
nor U7847 (N_7847,N_7718,N_7712);
or U7848 (N_7848,N_7711,N_7682);
nand U7849 (N_7849,N_7776,N_7698);
nor U7850 (N_7850,N_7752,N_7736);
nor U7851 (N_7851,N_7707,N_7726);
nand U7852 (N_7852,N_7652,N_7770);
or U7853 (N_7853,N_7734,N_7733);
and U7854 (N_7854,N_7699,N_7702);
nand U7855 (N_7855,N_7753,N_7720);
xor U7856 (N_7856,N_7799,N_7784);
or U7857 (N_7857,N_7796,N_7777);
and U7858 (N_7858,N_7691,N_7779);
or U7859 (N_7859,N_7653,N_7665);
and U7860 (N_7860,N_7778,N_7783);
nand U7861 (N_7861,N_7765,N_7651);
nand U7862 (N_7862,N_7763,N_7671);
nand U7863 (N_7863,N_7717,N_7781);
xor U7864 (N_7864,N_7797,N_7683);
and U7865 (N_7865,N_7740,N_7729);
nand U7866 (N_7866,N_7709,N_7669);
nor U7867 (N_7867,N_7768,N_7715);
xnor U7868 (N_7868,N_7680,N_7745);
and U7869 (N_7869,N_7771,N_7704);
nor U7870 (N_7870,N_7687,N_7761);
xnor U7871 (N_7871,N_7760,N_7684);
nor U7872 (N_7872,N_7787,N_7727);
or U7873 (N_7873,N_7706,N_7747);
xnor U7874 (N_7874,N_7754,N_7668);
xor U7875 (N_7875,N_7686,N_7757);
or U7876 (N_7876,N_7751,N_7690);
xor U7877 (N_7877,N_7759,N_7735);
or U7878 (N_7878,N_7735,N_7722);
and U7879 (N_7879,N_7667,N_7795);
nor U7880 (N_7880,N_7720,N_7731);
nor U7881 (N_7881,N_7674,N_7783);
xor U7882 (N_7882,N_7720,N_7716);
nor U7883 (N_7883,N_7688,N_7778);
nor U7884 (N_7884,N_7739,N_7710);
xnor U7885 (N_7885,N_7781,N_7777);
and U7886 (N_7886,N_7687,N_7725);
or U7887 (N_7887,N_7730,N_7685);
or U7888 (N_7888,N_7684,N_7695);
xor U7889 (N_7889,N_7746,N_7795);
or U7890 (N_7890,N_7761,N_7652);
or U7891 (N_7891,N_7683,N_7675);
and U7892 (N_7892,N_7741,N_7738);
or U7893 (N_7893,N_7717,N_7682);
and U7894 (N_7894,N_7760,N_7742);
xnor U7895 (N_7895,N_7686,N_7773);
xor U7896 (N_7896,N_7685,N_7789);
xnor U7897 (N_7897,N_7792,N_7771);
nor U7898 (N_7898,N_7726,N_7717);
and U7899 (N_7899,N_7791,N_7717);
xnor U7900 (N_7900,N_7762,N_7794);
or U7901 (N_7901,N_7794,N_7654);
or U7902 (N_7902,N_7722,N_7767);
nor U7903 (N_7903,N_7677,N_7683);
or U7904 (N_7904,N_7797,N_7735);
and U7905 (N_7905,N_7758,N_7732);
xor U7906 (N_7906,N_7737,N_7787);
xnor U7907 (N_7907,N_7779,N_7753);
nand U7908 (N_7908,N_7781,N_7753);
nand U7909 (N_7909,N_7697,N_7783);
or U7910 (N_7910,N_7751,N_7674);
xor U7911 (N_7911,N_7769,N_7664);
or U7912 (N_7912,N_7782,N_7659);
and U7913 (N_7913,N_7765,N_7784);
xnor U7914 (N_7914,N_7688,N_7701);
xor U7915 (N_7915,N_7709,N_7772);
and U7916 (N_7916,N_7650,N_7762);
nand U7917 (N_7917,N_7776,N_7750);
or U7918 (N_7918,N_7740,N_7725);
nand U7919 (N_7919,N_7751,N_7669);
xnor U7920 (N_7920,N_7667,N_7687);
xor U7921 (N_7921,N_7738,N_7663);
xnor U7922 (N_7922,N_7659,N_7716);
or U7923 (N_7923,N_7741,N_7746);
nor U7924 (N_7924,N_7674,N_7700);
and U7925 (N_7925,N_7750,N_7744);
xor U7926 (N_7926,N_7683,N_7771);
xnor U7927 (N_7927,N_7773,N_7721);
and U7928 (N_7928,N_7794,N_7691);
nand U7929 (N_7929,N_7766,N_7724);
or U7930 (N_7930,N_7675,N_7776);
xnor U7931 (N_7931,N_7689,N_7768);
and U7932 (N_7932,N_7743,N_7713);
and U7933 (N_7933,N_7683,N_7687);
xor U7934 (N_7934,N_7659,N_7728);
and U7935 (N_7935,N_7770,N_7796);
and U7936 (N_7936,N_7695,N_7783);
nand U7937 (N_7937,N_7741,N_7745);
nand U7938 (N_7938,N_7663,N_7736);
or U7939 (N_7939,N_7715,N_7785);
and U7940 (N_7940,N_7787,N_7797);
or U7941 (N_7941,N_7676,N_7656);
nor U7942 (N_7942,N_7759,N_7661);
nor U7943 (N_7943,N_7652,N_7756);
nand U7944 (N_7944,N_7787,N_7764);
xnor U7945 (N_7945,N_7721,N_7793);
xnor U7946 (N_7946,N_7678,N_7650);
or U7947 (N_7947,N_7682,N_7678);
nor U7948 (N_7948,N_7752,N_7683);
and U7949 (N_7949,N_7650,N_7655);
and U7950 (N_7950,N_7838,N_7913);
xor U7951 (N_7951,N_7870,N_7866);
nand U7952 (N_7952,N_7875,N_7939);
nor U7953 (N_7953,N_7807,N_7827);
or U7954 (N_7954,N_7850,N_7868);
and U7955 (N_7955,N_7847,N_7934);
nor U7956 (N_7956,N_7809,N_7890);
or U7957 (N_7957,N_7942,N_7873);
xnor U7958 (N_7958,N_7872,N_7918);
xor U7959 (N_7959,N_7898,N_7948);
and U7960 (N_7960,N_7940,N_7917);
nor U7961 (N_7961,N_7865,N_7846);
nand U7962 (N_7962,N_7857,N_7810);
nand U7963 (N_7963,N_7830,N_7831);
and U7964 (N_7964,N_7935,N_7931);
and U7965 (N_7965,N_7878,N_7819);
xnor U7966 (N_7966,N_7910,N_7906);
nor U7967 (N_7967,N_7837,N_7901);
nand U7968 (N_7968,N_7818,N_7888);
xnor U7969 (N_7969,N_7927,N_7909);
xnor U7970 (N_7970,N_7876,N_7922);
xnor U7971 (N_7971,N_7843,N_7801);
nor U7972 (N_7972,N_7928,N_7916);
nor U7973 (N_7973,N_7829,N_7854);
nor U7974 (N_7974,N_7895,N_7826);
nor U7975 (N_7975,N_7880,N_7840);
nor U7976 (N_7976,N_7947,N_7921);
xnor U7977 (N_7977,N_7896,N_7902);
nor U7978 (N_7978,N_7943,N_7937);
xnor U7979 (N_7979,N_7930,N_7856);
and U7980 (N_7980,N_7885,N_7825);
nand U7981 (N_7981,N_7897,N_7822);
xnor U7982 (N_7982,N_7849,N_7874);
xnor U7983 (N_7983,N_7852,N_7811);
nor U7984 (N_7984,N_7851,N_7899);
xnor U7985 (N_7985,N_7813,N_7848);
nand U7986 (N_7986,N_7867,N_7889);
nor U7987 (N_7987,N_7824,N_7853);
or U7988 (N_7988,N_7861,N_7859);
nand U7989 (N_7989,N_7863,N_7805);
and U7990 (N_7990,N_7871,N_7834);
nand U7991 (N_7991,N_7803,N_7891);
xor U7992 (N_7992,N_7932,N_7814);
xnor U7993 (N_7993,N_7938,N_7893);
nand U7994 (N_7994,N_7862,N_7925);
nor U7995 (N_7995,N_7894,N_7912);
and U7996 (N_7996,N_7903,N_7836);
nor U7997 (N_7997,N_7879,N_7883);
and U7998 (N_7998,N_7915,N_7923);
and U7999 (N_7999,N_7933,N_7820);
or U8000 (N_8000,N_7860,N_7842);
and U8001 (N_8001,N_7828,N_7946);
or U8002 (N_8002,N_7926,N_7833);
or U8003 (N_8003,N_7907,N_7941);
or U8004 (N_8004,N_7816,N_7841);
xnor U8005 (N_8005,N_7821,N_7845);
nor U8006 (N_8006,N_7900,N_7904);
and U8007 (N_8007,N_7835,N_7877);
or U8008 (N_8008,N_7949,N_7844);
xor U8009 (N_8009,N_7869,N_7892);
nand U8010 (N_8010,N_7812,N_7864);
nor U8011 (N_8011,N_7815,N_7855);
and U8012 (N_8012,N_7802,N_7911);
nor U8013 (N_8013,N_7808,N_7823);
xor U8014 (N_8014,N_7858,N_7914);
nor U8015 (N_8015,N_7905,N_7945);
or U8016 (N_8016,N_7817,N_7881);
or U8017 (N_8017,N_7806,N_7884);
xor U8018 (N_8018,N_7886,N_7887);
xnor U8019 (N_8019,N_7839,N_7804);
xnor U8020 (N_8020,N_7936,N_7882);
or U8021 (N_8021,N_7944,N_7920);
nor U8022 (N_8022,N_7908,N_7832);
xnor U8023 (N_8023,N_7800,N_7929);
xnor U8024 (N_8024,N_7924,N_7919);
or U8025 (N_8025,N_7882,N_7862);
nor U8026 (N_8026,N_7829,N_7949);
nand U8027 (N_8027,N_7939,N_7854);
nand U8028 (N_8028,N_7867,N_7824);
xnor U8029 (N_8029,N_7932,N_7853);
nand U8030 (N_8030,N_7903,N_7898);
or U8031 (N_8031,N_7897,N_7912);
xor U8032 (N_8032,N_7930,N_7825);
xor U8033 (N_8033,N_7947,N_7855);
nand U8034 (N_8034,N_7848,N_7905);
or U8035 (N_8035,N_7800,N_7867);
and U8036 (N_8036,N_7944,N_7861);
nor U8037 (N_8037,N_7853,N_7827);
xor U8038 (N_8038,N_7943,N_7946);
nor U8039 (N_8039,N_7899,N_7818);
or U8040 (N_8040,N_7875,N_7863);
nand U8041 (N_8041,N_7854,N_7884);
nor U8042 (N_8042,N_7947,N_7930);
or U8043 (N_8043,N_7947,N_7890);
and U8044 (N_8044,N_7807,N_7890);
nor U8045 (N_8045,N_7857,N_7867);
nor U8046 (N_8046,N_7870,N_7878);
or U8047 (N_8047,N_7823,N_7876);
and U8048 (N_8048,N_7919,N_7812);
xor U8049 (N_8049,N_7895,N_7832);
and U8050 (N_8050,N_7889,N_7926);
nor U8051 (N_8051,N_7915,N_7931);
nor U8052 (N_8052,N_7937,N_7885);
or U8053 (N_8053,N_7808,N_7851);
nand U8054 (N_8054,N_7931,N_7844);
xnor U8055 (N_8055,N_7921,N_7931);
xnor U8056 (N_8056,N_7940,N_7832);
nand U8057 (N_8057,N_7942,N_7888);
nor U8058 (N_8058,N_7849,N_7830);
xor U8059 (N_8059,N_7905,N_7837);
xor U8060 (N_8060,N_7884,N_7816);
xor U8061 (N_8061,N_7910,N_7886);
nand U8062 (N_8062,N_7899,N_7929);
xnor U8063 (N_8063,N_7938,N_7905);
nand U8064 (N_8064,N_7828,N_7864);
nor U8065 (N_8065,N_7931,N_7919);
and U8066 (N_8066,N_7852,N_7939);
xnor U8067 (N_8067,N_7840,N_7837);
xnor U8068 (N_8068,N_7922,N_7909);
nor U8069 (N_8069,N_7855,N_7879);
nor U8070 (N_8070,N_7934,N_7826);
nor U8071 (N_8071,N_7945,N_7889);
nor U8072 (N_8072,N_7905,N_7846);
nand U8073 (N_8073,N_7847,N_7879);
nand U8074 (N_8074,N_7861,N_7819);
nor U8075 (N_8075,N_7822,N_7839);
and U8076 (N_8076,N_7808,N_7802);
and U8077 (N_8077,N_7895,N_7802);
or U8078 (N_8078,N_7866,N_7935);
nor U8079 (N_8079,N_7920,N_7897);
nand U8080 (N_8080,N_7876,N_7892);
nor U8081 (N_8081,N_7889,N_7804);
or U8082 (N_8082,N_7940,N_7939);
xnor U8083 (N_8083,N_7867,N_7875);
xnor U8084 (N_8084,N_7803,N_7932);
or U8085 (N_8085,N_7855,N_7899);
or U8086 (N_8086,N_7914,N_7915);
nor U8087 (N_8087,N_7909,N_7948);
and U8088 (N_8088,N_7818,N_7921);
nand U8089 (N_8089,N_7866,N_7910);
and U8090 (N_8090,N_7936,N_7911);
xnor U8091 (N_8091,N_7939,N_7868);
and U8092 (N_8092,N_7841,N_7826);
nor U8093 (N_8093,N_7804,N_7929);
and U8094 (N_8094,N_7923,N_7934);
and U8095 (N_8095,N_7860,N_7879);
xnor U8096 (N_8096,N_7858,N_7826);
and U8097 (N_8097,N_7887,N_7915);
nor U8098 (N_8098,N_7940,N_7837);
nor U8099 (N_8099,N_7842,N_7935);
and U8100 (N_8100,N_8001,N_7984);
or U8101 (N_8101,N_8007,N_8089);
or U8102 (N_8102,N_8085,N_8010);
xnor U8103 (N_8103,N_8038,N_8070);
or U8104 (N_8104,N_8017,N_7992);
and U8105 (N_8105,N_7970,N_7965);
or U8106 (N_8106,N_8061,N_8059);
nand U8107 (N_8107,N_8063,N_7959);
or U8108 (N_8108,N_8024,N_8035);
and U8109 (N_8109,N_7967,N_8069);
xnor U8110 (N_8110,N_8034,N_8033);
xnor U8111 (N_8111,N_8012,N_8067);
nor U8112 (N_8112,N_7974,N_7954);
and U8113 (N_8113,N_7985,N_8040);
or U8114 (N_8114,N_8075,N_8073);
nand U8115 (N_8115,N_7994,N_8049);
nor U8116 (N_8116,N_8051,N_8030);
nand U8117 (N_8117,N_8068,N_8037);
and U8118 (N_8118,N_7955,N_8018);
and U8119 (N_8119,N_7968,N_8020);
xor U8120 (N_8120,N_7979,N_7972);
nand U8121 (N_8121,N_8099,N_8002);
nand U8122 (N_8122,N_8029,N_8013);
nor U8123 (N_8123,N_8021,N_8052);
nor U8124 (N_8124,N_8076,N_8026);
nand U8125 (N_8125,N_7988,N_7991);
xor U8126 (N_8126,N_7996,N_8084);
nand U8127 (N_8127,N_8036,N_7961);
and U8128 (N_8128,N_8009,N_8004);
nand U8129 (N_8129,N_8078,N_7962);
and U8130 (N_8130,N_7998,N_7957);
nor U8131 (N_8131,N_8048,N_7976);
nor U8132 (N_8132,N_7980,N_8066);
nand U8133 (N_8133,N_8005,N_7993);
or U8134 (N_8134,N_7977,N_7971);
nand U8135 (N_8135,N_8091,N_8016);
nand U8136 (N_8136,N_8093,N_8050);
or U8137 (N_8137,N_8080,N_7964);
nand U8138 (N_8138,N_7995,N_8081);
or U8139 (N_8139,N_8047,N_8065);
nor U8140 (N_8140,N_8041,N_7986);
nand U8141 (N_8141,N_8025,N_8071);
xnor U8142 (N_8142,N_8056,N_7953);
xor U8143 (N_8143,N_7982,N_7983);
xor U8144 (N_8144,N_7981,N_8045);
nand U8145 (N_8145,N_7973,N_7999);
xnor U8146 (N_8146,N_8032,N_8000);
nor U8147 (N_8147,N_8060,N_8011);
nand U8148 (N_8148,N_7958,N_8023);
or U8149 (N_8149,N_8088,N_7987);
and U8150 (N_8150,N_8097,N_7950);
nand U8151 (N_8151,N_8077,N_8072);
xor U8152 (N_8152,N_8074,N_7960);
or U8153 (N_8153,N_7989,N_8079);
nand U8154 (N_8154,N_8031,N_8003);
xnor U8155 (N_8155,N_8022,N_8042);
and U8156 (N_8156,N_8086,N_8019);
and U8157 (N_8157,N_8039,N_8057);
and U8158 (N_8158,N_8082,N_8054);
and U8159 (N_8159,N_8044,N_8027);
xor U8160 (N_8160,N_8046,N_8062);
or U8161 (N_8161,N_7975,N_8015);
xnor U8162 (N_8162,N_7952,N_8006);
and U8163 (N_8163,N_7963,N_8090);
and U8164 (N_8164,N_8098,N_8008);
xor U8165 (N_8165,N_7978,N_7997);
or U8166 (N_8166,N_8083,N_8095);
nand U8167 (N_8167,N_8064,N_7966);
nor U8168 (N_8168,N_7990,N_8043);
and U8169 (N_8169,N_8053,N_8055);
xor U8170 (N_8170,N_7951,N_8028);
nand U8171 (N_8171,N_7969,N_7956);
and U8172 (N_8172,N_8087,N_8014);
or U8173 (N_8173,N_8094,N_8092);
nand U8174 (N_8174,N_8096,N_8058);
and U8175 (N_8175,N_7961,N_8084);
xnor U8176 (N_8176,N_7986,N_8012);
nor U8177 (N_8177,N_7998,N_8084);
and U8178 (N_8178,N_8096,N_8030);
or U8179 (N_8179,N_8047,N_8075);
nor U8180 (N_8180,N_8007,N_7999);
and U8181 (N_8181,N_7999,N_8042);
and U8182 (N_8182,N_7959,N_8037);
nand U8183 (N_8183,N_7961,N_8051);
and U8184 (N_8184,N_8026,N_7976);
xnor U8185 (N_8185,N_8020,N_7978);
nor U8186 (N_8186,N_7986,N_7955);
nor U8187 (N_8187,N_8068,N_7996);
nand U8188 (N_8188,N_7993,N_7981);
or U8189 (N_8189,N_7962,N_7987);
nand U8190 (N_8190,N_7956,N_8001);
nand U8191 (N_8191,N_8016,N_8060);
and U8192 (N_8192,N_8007,N_8042);
or U8193 (N_8193,N_7989,N_8042);
xor U8194 (N_8194,N_8057,N_8042);
nor U8195 (N_8195,N_7989,N_7994);
nand U8196 (N_8196,N_8073,N_8025);
nand U8197 (N_8197,N_7972,N_7962);
xnor U8198 (N_8198,N_8043,N_8092);
nor U8199 (N_8199,N_7962,N_8076);
nor U8200 (N_8200,N_7969,N_7972);
xnor U8201 (N_8201,N_8026,N_7987);
or U8202 (N_8202,N_8038,N_7965);
nor U8203 (N_8203,N_7972,N_8026);
nand U8204 (N_8204,N_7975,N_7951);
nand U8205 (N_8205,N_8003,N_7990);
and U8206 (N_8206,N_7951,N_8003);
and U8207 (N_8207,N_8086,N_8054);
nand U8208 (N_8208,N_8019,N_7974);
nand U8209 (N_8209,N_8079,N_8010);
or U8210 (N_8210,N_8001,N_7957);
or U8211 (N_8211,N_7995,N_8037);
nand U8212 (N_8212,N_8079,N_7973);
xor U8213 (N_8213,N_7989,N_8011);
nor U8214 (N_8214,N_7977,N_8072);
nand U8215 (N_8215,N_8005,N_8001);
xnor U8216 (N_8216,N_7998,N_8079);
nor U8217 (N_8217,N_7965,N_7995);
xnor U8218 (N_8218,N_8009,N_8097);
xor U8219 (N_8219,N_8039,N_8064);
and U8220 (N_8220,N_7996,N_7959);
nor U8221 (N_8221,N_7982,N_7952);
xor U8222 (N_8222,N_8057,N_7990);
nor U8223 (N_8223,N_8099,N_8039);
xor U8224 (N_8224,N_7979,N_8015);
nand U8225 (N_8225,N_8086,N_8047);
nand U8226 (N_8226,N_8054,N_7959);
or U8227 (N_8227,N_8073,N_8012);
or U8228 (N_8228,N_8022,N_8063);
and U8229 (N_8229,N_7955,N_8002);
or U8230 (N_8230,N_7974,N_8061);
nor U8231 (N_8231,N_7974,N_7975);
nand U8232 (N_8232,N_8005,N_8065);
nor U8233 (N_8233,N_7956,N_8076);
nand U8234 (N_8234,N_8091,N_7962);
or U8235 (N_8235,N_8014,N_8069);
nand U8236 (N_8236,N_8035,N_8013);
xor U8237 (N_8237,N_7997,N_7983);
or U8238 (N_8238,N_8072,N_8025);
nand U8239 (N_8239,N_8060,N_8035);
nor U8240 (N_8240,N_8023,N_7973);
and U8241 (N_8241,N_7991,N_8006);
and U8242 (N_8242,N_8059,N_7975);
nor U8243 (N_8243,N_8037,N_8001);
xnor U8244 (N_8244,N_8002,N_8081);
xor U8245 (N_8245,N_8041,N_8070);
and U8246 (N_8246,N_7984,N_8000);
or U8247 (N_8247,N_7986,N_8099);
or U8248 (N_8248,N_8072,N_8082);
or U8249 (N_8249,N_7962,N_8005);
or U8250 (N_8250,N_8243,N_8191);
or U8251 (N_8251,N_8106,N_8216);
nor U8252 (N_8252,N_8100,N_8160);
and U8253 (N_8253,N_8228,N_8174);
and U8254 (N_8254,N_8169,N_8193);
xnor U8255 (N_8255,N_8171,N_8199);
xnor U8256 (N_8256,N_8224,N_8144);
or U8257 (N_8257,N_8143,N_8234);
nor U8258 (N_8258,N_8103,N_8212);
and U8259 (N_8259,N_8131,N_8196);
xnor U8260 (N_8260,N_8217,N_8248);
nand U8261 (N_8261,N_8222,N_8187);
or U8262 (N_8262,N_8192,N_8226);
xnor U8263 (N_8263,N_8215,N_8130);
xnor U8264 (N_8264,N_8116,N_8161);
or U8265 (N_8265,N_8205,N_8206);
or U8266 (N_8266,N_8190,N_8150);
and U8267 (N_8267,N_8126,N_8133);
nand U8268 (N_8268,N_8105,N_8120);
or U8269 (N_8269,N_8213,N_8180);
nor U8270 (N_8270,N_8127,N_8208);
and U8271 (N_8271,N_8112,N_8227);
or U8272 (N_8272,N_8156,N_8111);
nor U8273 (N_8273,N_8245,N_8157);
xnor U8274 (N_8274,N_8230,N_8207);
and U8275 (N_8275,N_8147,N_8233);
xnor U8276 (N_8276,N_8170,N_8214);
and U8277 (N_8277,N_8241,N_8194);
nand U8278 (N_8278,N_8238,N_8223);
xor U8279 (N_8279,N_8109,N_8183);
or U8280 (N_8280,N_8167,N_8134);
nor U8281 (N_8281,N_8113,N_8165);
xnor U8282 (N_8282,N_8202,N_8151);
and U8283 (N_8283,N_8128,N_8172);
or U8284 (N_8284,N_8110,N_8114);
nand U8285 (N_8285,N_8182,N_8142);
nor U8286 (N_8286,N_8219,N_8201);
xor U8287 (N_8287,N_8249,N_8232);
and U8288 (N_8288,N_8186,N_8218);
xnor U8289 (N_8289,N_8173,N_8239);
nor U8290 (N_8290,N_8139,N_8188);
nand U8291 (N_8291,N_8200,N_8135);
or U8292 (N_8292,N_8185,N_8102);
and U8293 (N_8293,N_8159,N_8119);
or U8294 (N_8294,N_8203,N_8242);
or U8295 (N_8295,N_8124,N_8195);
or U8296 (N_8296,N_8107,N_8198);
and U8297 (N_8297,N_8220,N_8132);
nand U8298 (N_8298,N_8145,N_8225);
xor U8299 (N_8299,N_8168,N_8122);
nor U8300 (N_8300,N_8118,N_8240);
or U8301 (N_8301,N_8247,N_8197);
xor U8302 (N_8302,N_8210,N_8149);
nand U8303 (N_8303,N_8152,N_8177);
or U8304 (N_8304,N_8229,N_8153);
nand U8305 (N_8305,N_8148,N_8231);
nor U8306 (N_8306,N_8236,N_8184);
nand U8307 (N_8307,N_8246,N_8244);
nor U8308 (N_8308,N_8158,N_8140);
or U8309 (N_8309,N_8146,N_8235);
nor U8310 (N_8310,N_8179,N_8125);
nand U8311 (N_8311,N_8178,N_8121);
xor U8312 (N_8312,N_8115,N_8108);
and U8313 (N_8313,N_8221,N_8117);
or U8314 (N_8314,N_8211,N_8136);
xnor U8315 (N_8315,N_8175,N_8155);
and U8316 (N_8316,N_8164,N_8162);
or U8317 (N_8317,N_8101,N_8138);
and U8318 (N_8318,N_8204,N_8104);
nand U8319 (N_8319,N_8176,N_8163);
nor U8320 (N_8320,N_8129,N_8209);
nor U8321 (N_8321,N_8237,N_8181);
and U8322 (N_8322,N_8154,N_8123);
nor U8323 (N_8323,N_8137,N_8166);
nand U8324 (N_8324,N_8141,N_8189);
nor U8325 (N_8325,N_8153,N_8103);
or U8326 (N_8326,N_8132,N_8174);
xnor U8327 (N_8327,N_8238,N_8196);
or U8328 (N_8328,N_8131,N_8137);
or U8329 (N_8329,N_8105,N_8102);
xnor U8330 (N_8330,N_8148,N_8210);
nor U8331 (N_8331,N_8140,N_8142);
xnor U8332 (N_8332,N_8221,N_8125);
and U8333 (N_8333,N_8171,N_8114);
xor U8334 (N_8334,N_8213,N_8220);
or U8335 (N_8335,N_8237,N_8145);
or U8336 (N_8336,N_8115,N_8249);
nor U8337 (N_8337,N_8140,N_8162);
nand U8338 (N_8338,N_8127,N_8140);
and U8339 (N_8339,N_8167,N_8126);
and U8340 (N_8340,N_8183,N_8175);
and U8341 (N_8341,N_8242,N_8113);
nand U8342 (N_8342,N_8124,N_8228);
xnor U8343 (N_8343,N_8182,N_8107);
and U8344 (N_8344,N_8246,N_8158);
nand U8345 (N_8345,N_8220,N_8232);
xnor U8346 (N_8346,N_8244,N_8220);
xnor U8347 (N_8347,N_8132,N_8173);
nor U8348 (N_8348,N_8189,N_8107);
or U8349 (N_8349,N_8173,N_8192);
xnor U8350 (N_8350,N_8150,N_8180);
or U8351 (N_8351,N_8129,N_8130);
or U8352 (N_8352,N_8171,N_8214);
nand U8353 (N_8353,N_8109,N_8215);
nand U8354 (N_8354,N_8113,N_8134);
nor U8355 (N_8355,N_8191,N_8166);
nand U8356 (N_8356,N_8122,N_8203);
or U8357 (N_8357,N_8104,N_8198);
nor U8358 (N_8358,N_8183,N_8141);
and U8359 (N_8359,N_8245,N_8228);
nor U8360 (N_8360,N_8247,N_8181);
nand U8361 (N_8361,N_8137,N_8212);
xnor U8362 (N_8362,N_8192,N_8184);
nor U8363 (N_8363,N_8233,N_8201);
xnor U8364 (N_8364,N_8115,N_8167);
and U8365 (N_8365,N_8215,N_8221);
xnor U8366 (N_8366,N_8203,N_8116);
or U8367 (N_8367,N_8223,N_8209);
xnor U8368 (N_8368,N_8247,N_8248);
nor U8369 (N_8369,N_8234,N_8136);
and U8370 (N_8370,N_8135,N_8249);
nand U8371 (N_8371,N_8137,N_8205);
or U8372 (N_8372,N_8122,N_8130);
xnor U8373 (N_8373,N_8234,N_8230);
nor U8374 (N_8374,N_8100,N_8109);
and U8375 (N_8375,N_8231,N_8135);
or U8376 (N_8376,N_8239,N_8192);
nand U8377 (N_8377,N_8201,N_8108);
or U8378 (N_8378,N_8120,N_8111);
and U8379 (N_8379,N_8193,N_8232);
nor U8380 (N_8380,N_8244,N_8214);
or U8381 (N_8381,N_8108,N_8248);
nand U8382 (N_8382,N_8214,N_8148);
nand U8383 (N_8383,N_8188,N_8154);
and U8384 (N_8384,N_8238,N_8171);
and U8385 (N_8385,N_8232,N_8175);
and U8386 (N_8386,N_8172,N_8173);
nor U8387 (N_8387,N_8114,N_8155);
nor U8388 (N_8388,N_8123,N_8187);
nand U8389 (N_8389,N_8216,N_8228);
or U8390 (N_8390,N_8224,N_8195);
nand U8391 (N_8391,N_8121,N_8160);
nand U8392 (N_8392,N_8111,N_8148);
nor U8393 (N_8393,N_8102,N_8195);
or U8394 (N_8394,N_8204,N_8102);
nand U8395 (N_8395,N_8142,N_8187);
nor U8396 (N_8396,N_8180,N_8168);
and U8397 (N_8397,N_8188,N_8197);
or U8398 (N_8398,N_8223,N_8197);
and U8399 (N_8399,N_8238,N_8188);
or U8400 (N_8400,N_8304,N_8254);
nand U8401 (N_8401,N_8259,N_8273);
nand U8402 (N_8402,N_8302,N_8334);
xor U8403 (N_8403,N_8368,N_8293);
and U8404 (N_8404,N_8319,N_8395);
or U8405 (N_8405,N_8356,N_8391);
nor U8406 (N_8406,N_8382,N_8326);
nor U8407 (N_8407,N_8397,N_8286);
and U8408 (N_8408,N_8301,N_8392);
nand U8409 (N_8409,N_8399,N_8353);
nor U8410 (N_8410,N_8369,N_8384);
and U8411 (N_8411,N_8388,N_8346);
nor U8412 (N_8412,N_8367,N_8372);
and U8413 (N_8413,N_8300,N_8398);
nand U8414 (N_8414,N_8295,N_8276);
or U8415 (N_8415,N_8299,N_8298);
nand U8416 (N_8416,N_8364,N_8283);
nand U8417 (N_8417,N_8269,N_8306);
nor U8418 (N_8418,N_8393,N_8282);
nand U8419 (N_8419,N_8387,N_8296);
or U8420 (N_8420,N_8379,N_8284);
nand U8421 (N_8421,N_8290,N_8362);
nor U8422 (N_8422,N_8294,N_8385);
nor U8423 (N_8423,N_8331,N_8263);
nor U8424 (N_8424,N_8349,N_8297);
and U8425 (N_8425,N_8303,N_8328);
or U8426 (N_8426,N_8355,N_8317);
nor U8427 (N_8427,N_8322,N_8352);
or U8428 (N_8428,N_8390,N_8321);
nand U8429 (N_8429,N_8255,N_8291);
or U8430 (N_8430,N_8377,N_8345);
nor U8431 (N_8431,N_8380,N_8309);
or U8432 (N_8432,N_8261,N_8361);
or U8433 (N_8433,N_8370,N_8251);
xor U8434 (N_8434,N_8280,N_8337);
or U8435 (N_8435,N_8262,N_8347);
and U8436 (N_8436,N_8376,N_8320);
or U8437 (N_8437,N_8308,N_8325);
or U8438 (N_8438,N_8310,N_8373);
nor U8439 (N_8439,N_8396,N_8252);
xor U8440 (N_8440,N_8365,N_8250);
nand U8441 (N_8441,N_8386,N_8332);
nand U8442 (N_8442,N_8289,N_8351);
or U8443 (N_8443,N_8335,N_8375);
xnor U8444 (N_8444,N_8358,N_8277);
and U8445 (N_8445,N_8339,N_8343);
or U8446 (N_8446,N_8312,N_8316);
nand U8447 (N_8447,N_8354,N_8260);
xnor U8448 (N_8448,N_8333,N_8287);
nand U8449 (N_8449,N_8253,N_8272);
nand U8450 (N_8450,N_8359,N_8265);
and U8451 (N_8451,N_8342,N_8275);
nand U8452 (N_8452,N_8281,N_8267);
or U8453 (N_8453,N_8271,N_8341);
and U8454 (N_8454,N_8338,N_8305);
and U8455 (N_8455,N_8315,N_8383);
nor U8456 (N_8456,N_8360,N_8381);
xnor U8457 (N_8457,N_8366,N_8274);
nand U8458 (N_8458,N_8266,N_8258);
nand U8459 (N_8459,N_8329,N_8314);
nor U8460 (N_8460,N_8371,N_8363);
nor U8461 (N_8461,N_8378,N_8327);
and U8462 (N_8462,N_8256,N_8279);
and U8463 (N_8463,N_8340,N_8285);
nand U8464 (N_8464,N_8278,N_8357);
nand U8465 (N_8465,N_8344,N_8313);
nand U8466 (N_8466,N_8270,N_8330);
and U8467 (N_8467,N_8311,N_8318);
xor U8468 (N_8468,N_8288,N_8394);
or U8469 (N_8469,N_8389,N_8348);
xor U8470 (N_8470,N_8324,N_8292);
and U8471 (N_8471,N_8257,N_8336);
xor U8472 (N_8472,N_8264,N_8350);
and U8473 (N_8473,N_8268,N_8374);
or U8474 (N_8474,N_8307,N_8323);
nand U8475 (N_8475,N_8397,N_8335);
or U8476 (N_8476,N_8327,N_8370);
and U8477 (N_8477,N_8385,N_8391);
and U8478 (N_8478,N_8292,N_8313);
xor U8479 (N_8479,N_8399,N_8264);
or U8480 (N_8480,N_8380,N_8297);
nand U8481 (N_8481,N_8251,N_8311);
and U8482 (N_8482,N_8317,N_8270);
nand U8483 (N_8483,N_8391,N_8363);
or U8484 (N_8484,N_8303,N_8381);
nand U8485 (N_8485,N_8281,N_8311);
nand U8486 (N_8486,N_8270,N_8354);
nand U8487 (N_8487,N_8371,N_8374);
nor U8488 (N_8488,N_8322,N_8275);
nand U8489 (N_8489,N_8372,N_8340);
or U8490 (N_8490,N_8355,N_8398);
or U8491 (N_8491,N_8282,N_8388);
and U8492 (N_8492,N_8316,N_8275);
nor U8493 (N_8493,N_8306,N_8341);
xnor U8494 (N_8494,N_8380,N_8307);
or U8495 (N_8495,N_8373,N_8348);
nor U8496 (N_8496,N_8325,N_8282);
or U8497 (N_8497,N_8317,N_8268);
or U8498 (N_8498,N_8348,N_8326);
xor U8499 (N_8499,N_8292,N_8317);
xnor U8500 (N_8500,N_8357,N_8337);
nand U8501 (N_8501,N_8253,N_8378);
nand U8502 (N_8502,N_8322,N_8268);
or U8503 (N_8503,N_8385,N_8267);
or U8504 (N_8504,N_8335,N_8253);
or U8505 (N_8505,N_8383,N_8364);
nand U8506 (N_8506,N_8349,N_8395);
nor U8507 (N_8507,N_8334,N_8303);
nor U8508 (N_8508,N_8378,N_8390);
and U8509 (N_8509,N_8305,N_8337);
nand U8510 (N_8510,N_8289,N_8304);
nor U8511 (N_8511,N_8337,N_8269);
and U8512 (N_8512,N_8314,N_8273);
nor U8513 (N_8513,N_8261,N_8319);
and U8514 (N_8514,N_8256,N_8369);
or U8515 (N_8515,N_8394,N_8261);
or U8516 (N_8516,N_8356,N_8336);
nand U8517 (N_8517,N_8296,N_8374);
xor U8518 (N_8518,N_8360,N_8261);
and U8519 (N_8519,N_8313,N_8254);
nor U8520 (N_8520,N_8374,N_8252);
nand U8521 (N_8521,N_8281,N_8252);
and U8522 (N_8522,N_8326,N_8398);
nor U8523 (N_8523,N_8317,N_8261);
xnor U8524 (N_8524,N_8305,N_8280);
xnor U8525 (N_8525,N_8366,N_8252);
xnor U8526 (N_8526,N_8293,N_8272);
and U8527 (N_8527,N_8287,N_8340);
and U8528 (N_8528,N_8312,N_8299);
nand U8529 (N_8529,N_8352,N_8324);
and U8530 (N_8530,N_8330,N_8313);
and U8531 (N_8531,N_8295,N_8361);
and U8532 (N_8532,N_8368,N_8342);
nor U8533 (N_8533,N_8252,N_8325);
and U8534 (N_8534,N_8359,N_8251);
and U8535 (N_8535,N_8350,N_8322);
and U8536 (N_8536,N_8389,N_8375);
nand U8537 (N_8537,N_8278,N_8250);
and U8538 (N_8538,N_8278,N_8388);
nand U8539 (N_8539,N_8304,N_8255);
or U8540 (N_8540,N_8269,N_8397);
nand U8541 (N_8541,N_8315,N_8374);
and U8542 (N_8542,N_8269,N_8348);
xor U8543 (N_8543,N_8372,N_8273);
nor U8544 (N_8544,N_8260,N_8329);
or U8545 (N_8545,N_8357,N_8388);
nand U8546 (N_8546,N_8306,N_8303);
and U8547 (N_8547,N_8377,N_8388);
and U8548 (N_8548,N_8337,N_8322);
nand U8549 (N_8549,N_8370,N_8362);
nor U8550 (N_8550,N_8491,N_8417);
or U8551 (N_8551,N_8523,N_8490);
or U8552 (N_8552,N_8487,N_8424);
nor U8553 (N_8553,N_8459,N_8460);
or U8554 (N_8554,N_8534,N_8464);
nand U8555 (N_8555,N_8405,N_8499);
and U8556 (N_8556,N_8429,N_8537);
xnor U8557 (N_8557,N_8481,N_8469);
or U8558 (N_8558,N_8532,N_8531);
nand U8559 (N_8559,N_8444,N_8522);
nand U8560 (N_8560,N_8435,N_8497);
xnor U8561 (N_8561,N_8547,N_8495);
nand U8562 (N_8562,N_8451,N_8529);
nand U8563 (N_8563,N_8488,N_8541);
xnor U8564 (N_8564,N_8479,N_8519);
nor U8565 (N_8565,N_8434,N_8473);
or U8566 (N_8566,N_8536,N_8420);
or U8567 (N_8567,N_8494,N_8516);
nor U8568 (N_8568,N_8507,N_8535);
nor U8569 (N_8569,N_8401,N_8442);
or U8570 (N_8570,N_8506,N_8478);
nand U8571 (N_8571,N_8440,N_8530);
or U8572 (N_8572,N_8456,N_8423);
and U8573 (N_8573,N_8482,N_8453);
and U8574 (N_8574,N_8528,N_8408);
or U8575 (N_8575,N_8533,N_8492);
or U8576 (N_8576,N_8496,N_8465);
xnor U8577 (N_8577,N_8443,N_8544);
and U8578 (N_8578,N_8433,N_8513);
xnor U8579 (N_8579,N_8437,N_8466);
and U8580 (N_8580,N_8501,N_8414);
xor U8581 (N_8581,N_8450,N_8505);
and U8582 (N_8582,N_8489,N_8483);
xor U8583 (N_8583,N_8455,N_8521);
xor U8584 (N_8584,N_8504,N_8503);
or U8585 (N_8585,N_8514,N_8546);
or U8586 (N_8586,N_8474,N_8421);
xnor U8587 (N_8587,N_8426,N_8549);
and U8588 (N_8588,N_8436,N_8407);
nor U8589 (N_8589,N_8411,N_8480);
xor U8590 (N_8590,N_8409,N_8548);
xor U8591 (N_8591,N_8500,N_8515);
nand U8592 (N_8592,N_8458,N_8502);
nand U8593 (N_8593,N_8454,N_8476);
and U8594 (N_8594,N_8538,N_8471);
xor U8595 (N_8595,N_8446,N_8477);
nor U8596 (N_8596,N_8427,N_8461);
and U8597 (N_8597,N_8509,N_8486);
nand U8598 (N_8598,N_8484,N_8517);
nand U8599 (N_8599,N_8539,N_8524);
and U8600 (N_8600,N_8415,N_8508);
and U8601 (N_8601,N_8425,N_8468);
and U8602 (N_8602,N_8428,N_8498);
xor U8603 (N_8603,N_8448,N_8472);
nand U8604 (N_8604,N_8403,N_8540);
and U8605 (N_8605,N_8430,N_8400);
nor U8606 (N_8606,N_8510,N_8493);
xnor U8607 (N_8607,N_8416,N_8545);
nand U8608 (N_8608,N_8422,N_8527);
xor U8609 (N_8609,N_8470,N_8449);
xor U8610 (N_8610,N_8542,N_8520);
xnor U8611 (N_8611,N_8404,N_8438);
nand U8612 (N_8612,N_8406,N_8485);
nor U8613 (N_8613,N_8410,N_8447);
nor U8614 (N_8614,N_8475,N_8445);
xor U8615 (N_8615,N_8463,N_8402);
xor U8616 (N_8616,N_8452,N_8441);
nor U8617 (N_8617,N_8439,N_8418);
nand U8618 (N_8618,N_8462,N_8467);
and U8619 (N_8619,N_8511,N_8431);
and U8620 (N_8620,N_8526,N_8432);
or U8621 (N_8621,N_8518,N_8525);
or U8622 (N_8622,N_8413,N_8457);
xnor U8623 (N_8623,N_8412,N_8419);
or U8624 (N_8624,N_8512,N_8543);
nand U8625 (N_8625,N_8425,N_8525);
nand U8626 (N_8626,N_8471,N_8411);
and U8627 (N_8627,N_8481,N_8446);
and U8628 (N_8628,N_8481,N_8478);
and U8629 (N_8629,N_8409,N_8473);
xor U8630 (N_8630,N_8466,N_8539);
xor U8631 (N_8631,N_8406,N_8524);
xnor U8632 (N_8632,N_8460,N_8487);
and U8633 (N_8633,N_8451,N_8512);
and U8634 (N_8634,N_8446,N_8403);
or U8635 (N_8635,N_8509,N_8406);
and U8636 (N_8636,N_8511,N_8527);
and U8637 (N_8637,N_8491,N_8527);
nor U8638 (N_8638,N_8442,N_8450);
nor U8639 (N_8639,N_8519,N_8404);
nor U8640 (N_8640,N_8450,N_8451);
or U8641 (N_8641,N_8540,N_8426);
nand U8642 (N_8642,N_8544,N_8517);
nand U8643 (N_8643,N_8500,N_8512);
xnor U8644 (N_8644,N_8444,N_8533);
xnor U8645 (N_8645,N_8545,N_8510);
or U8646 (N_8646,N_8499,N_8518);
nand U8647 (N_8647,N_8479,N_8522);
nor U8648 (N_8648,N_8449,N_8465);
or U8649 (N_8649,N_8423,N_8516);
and U8650 (N_8650,N_8406,N_8470);
nand U8651 (N_8651,N_8436,N_8459);
or U8652 (N_8652,N_8510,N_8517);
or U8653 (N_8653,N_8495,N_8523);
or U8654 (N_8654,N_8408,N_8486);
and U8655 (N_8655,N_8409,N_8485);
and U8656 (N_8656,N_8456,N_8498);
nor U8657 (N_8657,N_8502,N_8494);
nand U8658 (N_8658,N_8546,N_8492);
nand U8659 (N_8659,N_8420,N_8491);
xnor U8660 (N_8660,N_8496,N_8502);
nor U8661 (N_8661,N_8444,N_8528);
and U8662 (N_8662,N_8499,N_8507);
nor U8663 (N_8663,N_8533,N_8536);
and U8664 (N_8664,N_8511,N_8459);
nand U8665 (N_8665,N_8512,N_8417);
and U8666 (N_8666,N_8403,N_8543);
xor U8667 (N_8667,N_8547,N_8446);
nand U8668 (N_8668,N_8533,N_8419);
and U8669 (N_8669,N_8481,N_8427);
or U8670 (N_8670,N_8401,N_8418);
and U8671 (N_8671,N_8429,N_8548);
nor U8672 (N_8672,N_8433,N_8443);
and U8673 (N_8673,N_8476,N_8532);
and U8674 (N_8674,N_8500,N_8403);
or U8675 (N_8675,N_8420,N_8425);
and U8676 (N_8676,N_8490,N_8506);
nor U8677 (N_8677,N_8531,N_8479);
nand U8678 (N_8678,N_8546,N_8487);
or U8679 (N_8679,N_8541,N_8439);
and U8680 (N_8680,N_8410,N_8429);
and U8681 (N_8681,N_8436,N_8491);
and U8682 (N_8682,N_8535,N_8472);
or U8683 (N_8683,N_8512,N_8458);
and U8684 (N_8684,N_8534,N_8517);
or U8685 (N_8685,N_8480,N_8529);
xor U8686 (N_8686,N_8470,N_8429);
xor U8687 (N_8687,N_8415,N_8421);
nor U8688 (N_8688,N_8480,N_8515);
or U8689 (N_8689,N_8518,N_8515);
or U8690 (N_8690,N_8453,N_8473);
xor U8691 (N_8691,N_8538,N_8440);
or U8692 (N_8692,N_8503,N_8500);
and U8693 (N_8693,N_8504,N_8472);
xnor U8694 (N_8694,N_8478,N_8428);
nand U8695 (N_8695,N_8446,N_8540);
nand U8696 (N_8696,N_8402,N_8526);
or U8697 (N_8697,N_8520,N_8536);
nor U8698 (N_8698,N_8504,N_8411);
or U8699 (N_8699,N_8513,N_8483);
nand U8700 (N_8700,N_8688,N_8667);
nor U8701 (N_8701,N_8592,N_8629);
or U8702 (N_8702,N_8671,N_8633);
or U8703 (N_8703,N_8639,N_8643);
and U8704 (N_8704,N_8687,N_8694);
or U8705 (N_8705,N_8673,N_8577);
nand U8706 (N_8706,N_8644,N_8697);
or U8707 (N_8707,N_8576,N_8609);
xor U8708 (N_8708,N_8636,N_8686);
xor U8709 (N_8709,N_8564,N_8675);
nand U8710 (N_8710,N_8693,N_8572);
nand U8711 (N_8711,N_8660,N_8615);
and U8712 (N_8712,N_8678,N_8695);
and U8713 (N_8713,N_8611,N_8603);
nand U8714 (N_8714,N_8631,N_8648);
nor U8715 (N_8715,N_8655,N_8562);
xnor U8716 (N_8716,N_8582,N_8654);
or U8717 (N_8717,N_8612,N_8580);
xnor U8718 (N_8718,N_8657,N_8591);
xnor U8719 (N_8719,N_8550,N_8598);
nor U8720 (N_8720,N_8569,N_8561);
or U8721 (N_8721,N_8610,N_8677);
or U8722 (N_8722,N_8632,N_8627);
nand U8723 (N_8723,N_8696,N_8563);
or U8724 (N_8724,N_8659,N_8670);
nor U8725 (N_8725,N_8679,N_8662);
nor U8726 (N_8726,N_8650,N_8649);
or U8727 (N_8727,N_8668,N_8616);
or U8728 (N_8728,N_8652,N_8680);
nand U8729 (N_8729,N_8588,N_8596);
nor U8730 (N_8730,N_8692,N_8674);
xnor U8731 (N_8731,N_8589,N_8606);
nor U8732 (N_8732,N_8690,N_8607);
nand U8733 (N_8733,N_8663,N_8691);
nand U8734 (N_8734,N_8645,N_8669);
and U8735 (N_8735,N_8630,N_8618);
or U8736 (N_8736,N_8555,N_8658);
or U8737 (N_8737,N_8560,N_8684);
and U8738 (N_8738,N_8698,N_8640);
nand U8739 (N_8739,N_8672,N_8552);
and U8740 (N_8740,N_8614,N_8699);
nor U8741 (N_8741,N_8624,N_8575);
nand U8742 (N_8742,N_8584,N_8590);
or U8743 (N_8743,N_8601,N_8567);
nand U8744 (N_8744,N_8579,N_8571);
xor U8745 (N_8745,N_8634,N_8646);
nor U8746 (N_8746,N_8666,N_8622);
and U8747 (N_8747,N_8585,N_8554);
nand U8748 (N_8748,N_8566,N_8605);
xor U8749 (N_8749,N_8623,N_8638);
and U8750 (N_8750,N_8681,N_8557);
nor U8751 (N_8751,N_8597,N_8685);
nor U8752 (N_8752,N_8661,N_8682);
nor U8753 (N_8753,N_8551,N_8621);
or U8754 (N_8754,N_8613,N_8604);
or U8755 (N_8755,N_8581,N_8586);
or U8756 (N_8756,N_8553,N_8683);
or U8757 (N_8757,N_8573,N_8626);
or U8758 (N_8758,N_8635,N_8642);
xor U8759 (N_8759,N_8574,N_8676);
xnor U8760 (N_8760,N_8570,N_8602);
or U8761 (N_8761,N_8665,N_8628);
or U8762 (N_8762,N_8689,N_8664);
or U8763 (N_8763,N_8656,N_8583);
nand U8764 (N_8764,N_8651,N_8647);
nand U8765 (N_8765,N_8556,N_8620);
nand U8766 (N_8766,N_8617,N_8637);
nor U8767 (N_8767,N_8653,N_8625);
nand U8768 (N_8768,N_8587,N_8559);
and U8769 (N_8769,N_8600,N_8568);
or U8770 (N_8770,N_8565,N_8608);
xor U8771 (N_8771,N_8578,N_8593);
xnor U8772 (N_8772,N_8641,N_8594);
or U8773 (N_8773,N_8599,N_8558);
nor U8774 (N_8774,N_8595,N_8619);
and U8775 (N_8775,N_8691,N_8588);
xnor U8776 (N_8776,N_8629,N_8638);
nand U8777 (N_8777,N_8611,N_8666);
nand U8778 (N_8778,N_8553,N_8616);
nand U8779 (N_8779,N_8666,N_8677);
nor U8780 (N_8780,N_8574,N_8669);
or U8781 (N_8781,N_8583,N_8659);
xnor U8782 (N_8782,N_8599,N_8603);
xnor U8783 (N_8783,N_8642,N_8595);
or U8784 (N_8784,N_8638,N_8673);
nor U8785 (N_8785,N_8556,N_8688);
and U8786 (N_8786,N_8689,N_8602);
and U8787 (N_8787,N_8613,N_8569);
nand U8788 (N_8788,N_8698,N_8561);
nor U8789 (N_8789,N_8571,N_8667);
xnor U8790 (N_8790,N_8653,N_8575);
nor U8791 (N_8791,N_8627,N_8685);
nor U8792 (N_8792,N_8617,N_8656);
xor U8793 (N_8793,N_8627,N_8622);
or U8794 (N_8794,N_8597,N_8588);
nor U8795 (N_8795,N_8606,N_8644);
and U8796 (N_8796,N_8604,N_8594);
and U8797 (N_8797,N_8561,N_8681);
xnor U8798 (N_8798,N_8617,N_8687);
nand U8799 (N_8799,N_8611,N_8612);
xnor U8800 (N_8800,N_8594,N_8687);
xnor U8801 (N_8801,N_8615,N_8647);
nor U8802 (N_8802,N_8657,N_8589);
or U8803 (N_8803,N_8563,N_8585);
nor U8804 (N_8804,N_8611,N_8668);
nor U8805 (N_8805,N_8657,N_8663);
nand U8806 (N_8806,N_8583,N_8608);
or U8807 (N_8807,N_8591,N_8686);
nand U8808 (N_8808,N_8564,N_8577);
xnor U8809 (N_8809,N_8675,N_8572);
nor U8810 (N_8810,N_8596,N_8566);
and U8811 (N_8811,N_8586,N_8645);
nor U8812 (N_8812,N_8654,N_8598);
and U8813 (N_8813,N_8594,N_8572);
nand U8814 (N_8814,N_8697,N_8682);
or U8815 (N_8815,N_8616,N_8661);
and U8816 (N_8816,N_8578,N_8570);
and U8817 (N_8817,N_8649,N_8677);
nor U8818 (N_8818,N_8636,N_8644);
xor U8819 (N_8819,N_8637,N_8648);
and U8820 (N_8820,N_8659,N_8641);
nor U8821 (N_8821,N_8651,N_8551);
xnor U8822 (N_8822,N_8574,N_8675);
nand U8823 (N_8823,N_8588,N_8572);
and U8824 (N_8824,N_8619,N_8638);
and U8825 (N_8825,N_8698,N_8634);
or U8826 (N_8826,N_8659,N_8562);
and U8827 (N_8827,N_8631,N_8690);
and U8828 (N_8828,N_8561,N_8680);
nand U8829 (N_8829,N_8564,N_8578);
or U8830 (N_8830,N_8698,N_8673);
nand U8831 (N_8831,N_8669,N_8572);
and U8832 (N_8832,N_8593,N_8596);
nor U8833 (N_8833,N_8561,N_8604);
nand U8834 (N_8834,N_8617,N_8604);
xnor U8835 (N_8835,N_8697,N_8581);
and U8836 (N_8836,N_8694,N_8607);
nor U8837 (N_8837,N_8663,N_8553);
nand U8838 (N_8838,N_8552,N_8551);
nor U8839 (N_8839,N_8599,N_8653);
nor U8840 (N_8840,N_8647,N_8559);
and U8841 (N_8841,N_8699,N_8610);
xnor U8842 (N_8842,N_8656,N_8592);
xnor U8843 (N_8843,N_8606,N_8600);
and U8844 (N_8844,N_8694,N_8621);
and U8845 (N_8845,N_8557,N_8581);
xnor U8846 (N_8846,N_8630,N_8586);
xor U8847 (N_8847,N_8612,N_8563);
xnor U8848 (N_8848,N_8608,N_8563);
nand U8849 (N_8849,N_8672,N_8562);
nand U8850 (N_8850,N_8705,N_8769);
or U8851 (N_8851,N_8781,N_8805);
nor U8852 (N_8852,N_8842,N_8703);
xor U8853 (N_8853,N_8716,N_8812);
and U8854 (N_8854,N_8770,N_8749);
nor U8855 (N_8855,N_8784,N_8813);
nor U8856 (N_8856,N_8755,N_8829);
nand U8857 (N_8857,N_8789,N_8778);
and U8858 (N_8858,N_8782,N_8771);
or U8859 (N_8859,N_8754,N_8807);
nand U8860 (N_8860,N_8844,N_8794);
xor U8861 (N_8861,N_8840,N_8787);
nor U8862 (N_8862,N_8814,N_8841);
nor U8863 (N_8863,N_8801,N_8713);
and U8864 (N_8864,N_8762,N_8735);
or U8865 (N_8865,N_8779,N_8702);
xor U8866 (N_8866,N_8704,N_8803);
nand U8867 (N_8867,N_8712,N_8811);
or U8868 (N_8868,N_8739,N_8708);
or U8869 (N_8869,N_8768,N_8839);
xnor U8870 (N_8870,N_8791,N_8725);
nand U8871 (N_8871,N_8757,N_8810);
or U8872 (N_8872,N_8726,N_8700);
and U8873 (N_8873,N_8802,N_8847);
and U8874 (N_8874,N_8835,N_8711);
or U8875 (N_8875,N_8833,N_8738);
nand U8876 (N_8876,N_8798,N_8741);
xor U8877 (N_8877,N_8732,N_8720);
nor U8878 (N_8878,N_8743,N_8717);
and U8879 (N_8879,N_8736,N_8817);
and U8880 (N_8880,N_8724,N_8729);
or U8881 (N_8881,N_8848,N_8836);
xnor U8882 (N_8882,N_8828,N_8767);
nor U8883 (N_8883,N_8843,N_8758);
nand U8884 (N_8884,N_8747,N_8790);
xnor U8885 (N_8885,N_8760,N_8819);
xor U8886 (N_8886,N_8796,N_8753);
nand U8887 (N_8887,N_8765,N_8774);
xor U8888 (N_8888,N_8797,N_8837);
nand U8889 (N_8889,N_8746,N_8824);
or U8890 (N_8890,N_8849,N_8723);
nand U8891 (N_8891,N_8737,N_8752);
or U8892 (N_8892,N_8815,N_8709);
and U8893 (N_8893,N_8822,N_8777);
and U8894 (N_8894,N_8763,N_8823);
nand U8895 (N_8895,N_8831,N_8804);
nor U8896 (N_8896,N_8826,N_8845);
xor U8897 (N_8897,N_8728,N_8785);
or U8898 (N_8898,N_8714,N_8780);
nor U8899 (N_8899,N_8745,N_8764);
and U8900 (N_8900,N_8731,N_8775);
nor U8901 (N_8901,N_8821,N_8710);
and U8902 (N_8902,N_8846,N_8786);
xnor U8903 (N_8903,N_8759,N_8792);
or U8904 (N_8904,N_8832,N_8788);
nor U8905 (N_8905,N_8719,N_8806);
or U8906 (N_8906,N_8834,N_8838);
or U8907 (N_8907,N_8783,N_8734);
nor U8908 (N_8908,N_8776,N_8809);
xor U8909 (N_8909,N_8706,N_8816);
xor U8910 (N_8910,N_8800,N_8740);
nand U8911 (N_8911,N_8730,N_8733);
or U8912 (N_8912,N_8808,N_8820);
and U8913 (N_8913,N_8744,N_8830);
or U8914 (N_8914,N_8750,N_8761);
xor U8915 (N_8915,N_8742,N_8827);
or U8916 (N_8916,N_8825,N_8718);
nand U8917 (N_8917,N_8721,N_8818);
xnor U8918 (N_8918,N_8773,N_8766);
and U8919 (N_8919,N_8722,N_8748);
xor U8920 (N_8920,N_8799,N_8793);
xor U8921 (N_8921,N_8701,N_8795);
or U8922 (N_8922,N_8751,N_8756);
and U8923 (N_8923,N_8707,N_8772);
or U8924 (N_8924,N_8727,N_8715);
xor U8925 (N_8925,N_8707,N_8774);
nand U8926 (N_8926,N_8737,N_8809);
xor U8927 (N_8927,N_8811,N_8846);
or U8928 (N_8928,N_8741,N_8794);
or U8929 (N_8929,N_8774,N_8739);
nand U8930 (N_8930,N_8775,N_8776);
or U8931 (N_8931,N_8783,N_8795);
nor U8932 (N_8932,N_8758,N_8749);
and U8933 (N_8933,N_8843,N_8746);
and U8934 (N_8934,N_8845,N_8777);
nand U8935 (N_8935,N_8841,N_8812);
nor U8936 (N_8936,N_8814,N_8759);
xnor U8937 (N_8937,N_8829,N_8841);
nand U8938 (N_8938,N_8847,N_8733);
nor U8939 (N_8939,N_8779,N_8827);
xor U8940 (N_8940,N_8811,N_8731);
nand U8941 (N_8941,N_8798,N_8827);
and U8942 (N_8942,N_8821,N_8838);
nand U8943 (N_8943,N_8787,N_8809);
and U8944 (N_8944,N_8749,N_8804);
or U8945 (N_8945,N_8823,N_8820);
or U8946 (N_8946,N_8793,N_8824);
xor U8947 (N_8947,N_8727,N_8728);
xnor U8948 (N_8948,N_8701,N_8715);
and U8949 (N_8949,N_8830,N_8717);
and U8950 (N_8950,N_8779,N_8819);
and U8951 (N_8951,N_8710,N_8830);
xor U8952 (N_8952,N_8790,N_8716);
and U8953 (N_8953,N_8795,N_8726);
and U8954 (N_8954,N_8725,N_8743);
nand U8955 (N_8955,N_8741,N_8782);
and U8956 (N_8956,N_8827,N_8753);
nor U8957 (N_8957,N_8786,N_8837);
and U8958 (N_8958,N_8750,N_8831);
and U8959 (N_8959,N_8763,N_8843);
nor U8960 (N_8960,N_8785,N_8807);
or U8961 (N_8961,N_8820,N_8708);
or U8962 (N_8962,N_8809,N_8733);
and U8963 (N_8963,N_8731,N_8722);
nor U8964 (N_8964,N_8838,N_8808);
or U8965 (N_8965,N_8722,N_8730);
nand U8966 (N_8966,N_8828,N_8829);
and U8967 (N_8967,N_8760,N_8770);
nor U8968 (N_8968,N_8841,N_8831);
and U8969 (N_8969,N_8748,N_8813);
nand U8970 (N_8970,N_8772,N_8813);
xnor U8971 (N_8971,N_8757,N_8825);
or U8972 (N_8972,N_8735,N_8792);
nor U8973 (N_8973,N_8818,N_8842);
or U8974 (N_8974,N_8768,N_8742);
and U8975 (N_8975,N_8820,N_8775);
or U8976 (N_8976,N_8809,N_8703);
nand U8977 (N_8977,N_8847,N_8707);
xor U8978 (N_8978,N_8836,N_8713);
nand U8979 (N_8979,N_8724,N_8814);
xor U8980 (N_8980,N_8730,N_8841);
nand U8981 (N_8981,N_8736,N_8704);
nand U8982 (N_8982,N_8847,N_8825);
nor U8983 (N_8983,N_8827,N_8746);
nand U8984 (N_8984,N_8780,N_8763);
or U8985 (N_8985,N_8760,N_8777);
xnor U8986 (N_8986,N_8796,N_8736);
or U8987 (N_8987,N_8807,N_8815);
nor U8988 (N_8988,N_8747,N_8796);
xnor U8989 (N_8989,N_8812,N_8790);
nand U8990 (N_8990,N_8725,N_8724);
and U8991 (N_8991,N_8847,N_8796);
or U8992 (N_8992,N_8833,N_8818);
or U8993 (N_8993,N_8808,N_8728);
xor U8994 (N_8994,N_8839,N_8798);
and U8995 (N_8995,N_8717,N_8838);
xor U8996 (N_8996,N_8782,N_8776);
nor U8997 (N_8997,N_8846,N_8726);
xor U8998 (N_8998,N_8793,N_8771);
or U8999 (N_8999,N_8765,N_8755);
nor U9000 (N_9000,N_8888,N_8991);
or U9001 (N_9001,N_8959,N_8910);
or U9002 (N_9002,N_8873,N_8977);
or U9003 (N_9003,N_8972,N_8853);
nor U9004 (N_9004,N_8997,N_8887);
or U9005 (N_9005,N_8957,N_8858);
xnor U9006 (N_9006,N_8978,N_8894);
nand U9007 (N_9007,N_8996,N_8893);
nand U9008 (N_9008,N_8881,N_8979);
or U9009 (N_9009,N_8983,N_8925);
nor U9010 (N_9010,N_8871,N_8967);
nor U9011 (N_9011,N_8913,N_8960);
nor U9012 (N_9012,N_8889,N_8966);
and U9013 (N_9013,N_8902,N_8929);
xnor U9014 (N_9014,N_8980,N_8974);
nor U9015 (N_9015,N_8964,N_8868);
or U9016 (N_9016,N_8956,N_8870);
nand U9017 (N_9017,N_8916,N_8874);
nand U9018 (N_9018,N_8994,N_8914);
xnor U9019 (N_9019,N_8892,N_8990);
or U9020 (N_9020,N_8962,N_8900);
xor U9021 (N_9021,N_8863,N_8985);
nor U9022 (N_9022,N_8952,N_8981);
nand U9023 (N_9023,N_8919,N_8896);
xor U9024 (N_9024,N_8936,N_8989);
nand U9025 (N_9025,N_8884,N_8965);
xor U9026 (N_9026,N_8963,N_8975);
nand U9027 (N_9027,N_8982,N_8999);
or U9028 (N_9028,N_8905,N_8876);
and U9029 (N_9029,N_8854,N_8922);
and U9030 (N_9030,N_8865,N_8950);
nor U9031 (N_9031,N_8941,N_8867);
xnor U9032 (N_9032,N_8866,N_8945);
and U9033 (N_9033,N_8855,N_8992);
nor U9034 (N_9034,N_8882,N_8890);
nand U9035 (N_9035,N_8953,N_8943);
xnor U9036 (N_9036,N_8850,N_8986);
xor U9037 (N_9037,N_8969,N_8949);
or U9038 (N_9038,N_8946,N_8917);
nor U9039 (N_9039,N_8988,N_8880);
or U9040 (N_9040,N_8932,N_8976);
nand U9041 (N_9041,N_8901,N_8906);
or U9042 (N_9042,N_8852,N_8859);
or U9043 (N_9043,N_8973,N_8885);
xor U9044 (N_9044,N_8860,N_8861);
and U9045 (N_9045,N_8869,N_8878);
nand U9046 (N_9046,N_8933,N_8944);
nand U9047 (N_9047,N_8924,N_8899);
or U9048 (N_9048,N_8904,N_8921);
or U9049 (N_9049,N_8984,N_8897);
nand U9050 (N_9050,N_8955,N_8875);
nand U9051 (N_9051,N_8879,N_8909);
nor U9052 (N_9052,N_8864,N_8987);
nor U9053 (N_9053,N_8948,N_8931);
nand U9054 (N_9054,N_8934,N_8851);
or U9055 (N_9055,N_8942,N_8940);
nor U9056 (N_9056,N_8971,N_8939);
xnor U9057 (N_9057,N_8958,N_8995);
and U9058 (N_9058,N_8908,N_8954);
nor U9059 (N_9059,N_8928,N_8912);
nor U9060 (N_9060,N_8935,N_8993);
or U9061 (N_9061,N_8920,N_8961);
nor U9062 (N_9062,N_8947,N_8907);
nand U9063 (N_9063,N_8895,N_8998);
or U9064 (N_9064,N_8930,N_8923);
nand U9065 (N_9065,N_8856,N_8872);
or U9066 (N_9066,N_8898,N_8862);
nor U9067 (N_9067,N_8926,N_8886);
nand U9068 (N_9068,N_8951,N_8927);
or U9069 (N_9069,N_8877,N_8915);
or U9070 (N_9070,N_8903,N_8911);
or U9071 (N_9071,N_8857,N_8938);
and U9072 (N_9072,N_8918,N_8891);
or U9073 (N_9073,N_8937,N_8968);
xnor U9074 (N_9074,N_8883,N_8970);
xnor U9075 (N_9075,N_8954,N_8935);
and U9076 (N_9076,N_8919,N_8946);
xnor U9077 (N_9077,N_8889,N_8912);
xor U9078 (N_9078,N_8860,N_8892);
nor U9079 (N_9079,N_8915,N_8856);
and U9080 (N_9080,N_8998,N_8873);
nor U9081 (N_9081,N_8938,N_8908);
nor U9082 (N_9082,N_8910,N_8981);
nor U9083 (N_9083,N_8948,N_8854);
nand U9084 (N_9084,N_8856,N_8934);
xor U9085 (N_9085,N_8989,N_8877);
or U9086 (N_9086,N_8902,N_8872);
xnor U9087 (N_9087,N_8958,N_8998);
nor U9088 (N_9088,N_8939,N_8968);
and U9089 (N_9089,N_8872,N_8950);
nor U9090 (N_9090,N_8910,N_8935);
nand U9091 (N_9091,N_8941,N_8981);
or U9092 (N_9092,N_8867,N_8909);
nand U9093 (N_9093,N_8982,N_8911);
and U9094 (N_9094,N_8936,N_8919);
nor U9095 (N_9095,N_8937,N_8911);
xnor U9096 (N_9096,N_8971,N_8945);
and U9097 (N_9097,N_8880,N_8969);
nor U9098 (N_9098,N_8924,N_8890);
and U9099 (N_9099,N_8870,N_8980);
xor U9100 (N_9100,N_8990,N_8998);
nand U9101 (N_9101,N_8881,N_8972);
or U9102 (N_9102,N_8907,N_8900);
and U9103 (N_9103,N_8921,N_8962);
or U9104 (N_9104,N_8938,N_8933);
or U9105 (N_9105,N_8861,N_8882);
nand U9106 (N_9106,N_8854,N_8893);
nand U9107 (N_9107,N_8951,N_8855);
xnor U9108 (N_9108,N_8943,N_8904);
nand U9109 (N_9109,N_8946,N_8925);
nor U9110 (N_9110,N_8945,N_8908);
nor U9111 (N_9111,N_8962,N_8867);
xnor U9112 (N_9112,N_8869,N_8901);
nor U9113 (N_9113,N_8975,N_8905);
or U9114 (N_9114,N_8877,N_8894);
xor U9115 (N_9115,N_8961,N_8869);
xnor U9116 (N_9116,N_8859,N_8985);
and U9117 (N_9117,N_8860,N_8875);
and U9118 (N_9118,N_8992,N_8974);
nand U9119 (N_9119,N_8896,N_8851);
xnor U9120 (N_9120,N_8906,N_8937);
xor U9121 (N_9121,N_8965,N_8958);
nand U9122 (N_9122,N_8950,N_8873);
and U9123 (N_9123,N_8958,N_8984);
nand U9124 (N_9124,N_8964,N_8989);
nor U9125 (N_9125,N_8949,N_8866);
nand U9126 (N_9126,N_8992,N_8898);
or U9127 (N_9127,N_8978,N_8898);
or U9128 (N_9128,N_8958,N_8907);
and U9129 (N_9129,N_8986,N_8921);
and U9130 (N_9130,N_8938,N_8924);
and U9131 (N_9131,N_8940,N_8944);
nor U9132 (N_9132,N_8851,N_8947);
nand U9133 (N_9133,N_8969,N_8864);
and U9134 (N_9134,N_8950,N_8879);
nor U9135 (N_9135,N_8880,N_8853);
xnor U9136 (N_9136,N_8980,N_8898);
nor U9137 (N_9137,N_8878,N_8877);
or U9138 (N_9138,N_8866,N_8916);
nor U9139 (N_9139,N_8866,N_8951);
and U9140 (N_9140,N_8882,N_8854);
and U9141 (N_9141,N_8976,N_8875);
and U9142 (N_9142,N_8899,N_8891);
and U9143 (N_9143,N_8869,N_8867);
and U9144 (N_9144,N_8997,N_8954);
xor U9145 (N_9145,N_8890,N_8952);
xnor U9146 (N_9146,N_8918,N_8924);
or U9147 (N_9147,N_8957,N_8976);
nand U9148 (N_9148,N_8879,N_8917);
nand U9149 (N_9149,N_8858,N_8940);
or U9150 (N_9150,N_9041,N_9143);
nand U9151 (N_9151,N_9061,N_9092);
nor U9152 (N_9152,N_9008,N_9138);
or U9153 (N_9153,N_9067,N_9023);
nor U9154 (N_9154,N_9047,N_9050);
and U9155 (N_9155,N_9112,N_9003);
nand U9156 (N_9156,N_9046,N_9146);
nor U9157 (N_9157,N_9139,N_9072);
and U9158 (N_9158,N_9076,N_9000);
nor U9159 (N_9159,N_9094,N_9096);
or U9160 (N_9160,N_9117,N_9021);
and U9161 (N_9161,N_9032,N_9049);
nand U9162 (N_9162,N_9090,N_9005);
nand U9163 (N_9163,N_9101,N_9013);
xnor U9164 (N_9164,N_9051,N_9056);
and U9165 (N_9165,N_9033,N_9048);
and U9166 (N_9166,N_9075,N_9009);
and U9167 (N_9167,N_9016,N_9108);
xnor U9168 (N_9168,N_9135,N_9084);
nor U9169 (N_9169,N_9042,N_9098);
nand U9170 (N_9170,N_9105,N_9071);
nand U9171 (N_9171,N_9093,N_9057);
and U9172 (N_9172,N_9054,N_9040);
xnor U9173 (N_9173,N_9074,N_9118);
or U9174 (N_9174,N_9080,N_9002);
and U9175 (N_9175,N_9011,N_9132);
and U9176 (N_9176,N_9116,N_9022);
nor U9177 (N_9177,N_9095,N_9102);
or U9178 (N_9178,N_9130,N_9088);
nand U9179 (N_9179,N_9129,N_9086);
nor U9180 (N_9180,N_9060,N_9062);
nor U9181 (N_9181,N_9106,N_9128);
nand U9182 (N_9182,N_9030,N_9134);
and U9183 (N_9183,N_9019,N_9052);
nand U9184 (N_9184,N_9149,N_9031);
xor U9185 (N_9185,N_9028,N_9127);
xnor U9186 (N_9186,N_9133,N_9091);
nand U9187 (N_9187,N_9014,N_9079);
xor U9188 (N_9188,N_9007,N_9120);
xnor U9189 (N_9189,N_9073,N_9137);
xnor U9190 (N_9190,N_9126,N_9124);
and U9191 (N_9191,N_9045,N_9148);
nor U9192 (N_9192,N_9109,N_9068);
xnor U9193 (N_9193,N_9026,N_9081);
or U9194 (N_9194,N_9024,N_9037);
or U9195 (N_9195,N_9082,N_9131);
nand U9196 (N_9196,N_9114,N_9125);
xnor U9197 (N_9197,N_9121,N_9064);
and U9198 (N_9198,N_9103,N_9140);
nor U9199 (N_9199,N_9100,N_9053);
nand U9200 (N_9200,N_9069,N_9097);
nand U9201 (N_9201,N_9038,N_9010);
nor U9202 (N_9202,N_9136,N_9115);
or U9203 (N_9203,N_9055,N_9087);
or U9204 (N_9204,N_9029,N_9059);
and U9205 (N_9205,N_9144,N_9044);
or U9206 (N_9206,N_9123,N_9036);
and U9207 (N_9207,N_9020,N_9089);
or U9208 (N_9208,N_9099,N_9017);
and U9209 (N_9209,N_9141,N_9006);
nor U9210 (N_9210,N_9142,N_9066);
or U9211 (N_9211,N_9015,N_9110);
and U9212 (N_9212,N_9058,N_9004);
or U9213 (N_9213,N_9070,N_9147);
nor U9214 (N_9214,N_9085,N_9043);
and U9215 (N_9215,N_9065,N_9113);
nand U9216 (N_9216,N_9012,N_9083);
and U9217 (N_9217,N_9035,N_9107);
and U9218 (N_9218,N_9025,N_9018);
or U9219 (N_9219,N_9111,N_9145);
nand U9220 (N_9220,N_9063,N_9077);
or U9221 (N_9221,N_9039,N_9122);
nand U9222 (N_9222,N_9027,N_9078);
xor U9223 (N_9223,N_9001,N_9119);
nand U9224 (N_9224,N_9034,N_9104);
or U9225 (N_9225,N_9129,N_9108);
nand U9226 (N_9226,N_9128,N_9073);
and U9227 (N_9227,N_9062,N_9090);
nor U9228 (N_9228,N_9036,N_9083);
xor U9229 (N_9229,N_9126,N_9095);
xnor U9230 (N_9230,N_9112,N_9079);
nand U9231 (N_9231,N_9016,N_9038);
and U9232 (N_9232,N_9014,N_9129);
nand U9233 (N_9233,N_9003,N_9117);
or U9234 (N_9234,N_9019,N_9071);
or U9235 (N_9235,N_9146,N_9001);
xnor U9236 (N_9236,N_9066,N_9005);
nor U9237 (N_9237,N_9088,N_9011);
xor U9238 (N_9238,N_9148,N_9103);
xor U9239 (N_9239,N_9067,N_9102);
xor U9240 (N_9240,N_9114,N_9022);
or U9241 (N_9241,N_9088,N_9008);
nand U9242 (N_9242,N_9004,N_9040);
xor U9243 (N_9243,N_9117,N_9124);
or U9244 (N_9244,N_9019,N_9013);
xnor U9245 (N_9245,N_9021,N_9095);
nor U9246 (N_9246,N_9103,N_9055);
nor U9247 (N_9247,N_9148,N_9146);
nand U9248 (N_9248,N_9015,N_9068);
nor U9249 (N_9249,N_9081,N_9013);
or U9250 (N_9250,N_9135,N_9069);
nor U9251 (N_9251,N_9049,N_9118);
xor U9252 (N_9252,N_9048,N_9015);
nand U9253 (N_9253,N_9099,N_9094);
nor U9254 (N_9254,N_9071,N_9045);
nor U9255 (N_9255,N_9068,N_9117);
and U9256 (N_9256,N_9040,N_9134);
xnor U9257 (N_9257,N_9008,N_9062);
and U9258 (N_9258,N_9049,N_9031);
or U9259 (N_9259,N_9089,N_9056);
or U9260 (N_9260,N_9100,N_9119);
and U9261 (N_9261,N_9012,N_9080);
nor U9262 (N_9262,N_9040,N_9137);
xnor U9263 (N_9263,N_9073,N_9038);
nor U9264 (N_9264,N_9115,N_9010);
or U9265 (N_9265,N_9130,N_9095);
xnor U9266 (N_9266,N_9121,N_9011);
nor U9267 (N_9267,N_9148,N_9064);
or U9268 (N_9268,N_9043,N_9099);
or U9269 (N_9269,N_9099,N_9010);
nand U9270 (N_9270,N_9018,N_9013);
or U9271 (N_9271,N_9014,N_9127);
or U9272 (N_9272,N_9148,N_9036);
nand U9273 (N_9273,N_9130,N_9010);
or U9274 (N_9274,N_9114,N_9028);
xor U9275 (N_9275,N_9027,N_9147);
nand U9276 (N_9276,N_9125,N_9096);
and U9277 (N_9277,N_9021,N_9058);
or U9278 (N_9278,N_9114,N_9083);
nand U9279 (N_9279,N_9011,N_9098);
nor U9280 (N_9280,N_9060,N_9089);
nor U9281 (N_9281,N_9119,N_9052);
or U9282 (N_9282,N_9006,N_9113);
and U9283 (N_9283,N_9133,N_9034);
nand U9284 (N_9284,N_9035,N_9044);
nor U9285 (N_9285,N_9056,N_9144);
nor U9286 (N_9286,N_9062,N_9129);
or U9287 (N_9287,N_9097,N_9003);
nor U9288 (N_9288,N_9044,N_9065);
nor U9289 (N_9289,N_9043,N_9134);
nand U9290 (N_9290,N_9103,N_9024);
or U9291 (N_9291,N_9066,N_9035);
and U9292 (N_9292,N_9101,N_9076);
or U9293 (N_9293,N_9021,N_9007);
or U9294 (N_9294,N_9120,N_9016);
or U9295 (N_9295,N_9110,N_9134);
nand U9296 (N_9296,N_9014,N_9091);
nor U9297 (N_9297,N_9013,N_9039);
nand U9298 (N_9298,N_9117,N_9128);
nand U9299 (N_9299,N_9121,N_9131);
and U9300 (N_9300,N_9288,N_9225);
or U9301 (N_9301,N_9290,N_9242);
nand U9302 (N_9302,N_9297,N_9191);
and U9303 (N_9303,N_9292,N_9189);
xnor U9304 (N_9304,N_9190,N_9176);
or U9305 (N_9305,N_9237,N_9230);
nor U9306 (N_9306,N_9259,N_9188);
nand U9307 (N_9307,N_9272,N_9287);
nand U9308 (N_9308,N_9211,N_9204);
and U9309 (N_9309,N_9286,N_9258);
and U9310 (N_9310,N_9218,N_9267);
nand U9311 (N_9311,N_9262,N_9195);
and U9312 (N_9312,N_9260,N_9275);
xor U9313 (N_9313,N_9210,N_9171);
and U9314 (N_9314,N_9165,N_9269);
nand U9315 (N_9315,N_9174,N_9232);
nand U9316 (N_9316,N_9264,N_9213);
and U9317 (N_9317,N_9152,N_9219);
nand U9318 (N_9318,N_9294,N_9257);
or U9319 (N_9319,N_9207,N_9192);
and U9320 (N_9320,N_9157,N_9214);
and U9321 (N_9321,N_9229,N_9185);
and U9322 (N_9322,N_9251,N_9276);
nand U9323 (N_9323,N_9274,N_9180);
xor U9324 (N_9324,N_9293,N_9254);
xnor U9325 (N_9325,N_9239,N_9205);
and U9326 (N_9326,N_9154,N_9158);
xnor U9327 (N_9327,N_9212,N_9209);
or U9328 (N_9328,N_9256,N_9243);
and U9329 (N_9329,N_9271,N_9155);
nor U9330 (N_9330,N_9270,N_9248);
and U9331 (N_9331,N_9238,N_9253);
nor U9332 (N_9332,N_9208,N_9244);
nor U9333 (N_9333,N_9175,N_9181);
nand U9334 (N_9334,N_9217,N_9201);
nor U9335 (N_9335,N_9277,N_9196);
and U9336 (N_9336,N_9227,N_9241);
nand U9337 (N_9337,N_9159,N_9161);
or U9338 (N_9338,N_9178,N_9255);
xor U9339 (N_9339,N_9206,N_9252);
nor U9340 (N_9340,N_9198,N_9250);
nand U9341 (N_9341,N_9279,N_9182);
xor U9342 (N_9342,N_9167,N_9249);
xor U9343 (N_9343,N_9295,N_9202);
nor U9344 (N_9344,N_9298,N_9186);
xor U9345 (N_9345,N_9216,N_9184);
xor U9346 (N_9346,N_9280,N_9197);
and U9347 (N_9347,N_9164,N_9173);
xor U9348 (N_9348,N_9240,N_9215);
and U9349 (N_9349,N_9168,N_9266);
nand U9350 (N_9350,N_9156,N_9299);
and U9351 (N_9351,N_9222,N_9183);
nand U9352 (N_9352,N_9234,N_9224);
xnor U9353 (N_9353,N_9153,N_9235);
and U9354 (N_9354,N_9281,N_9194);
xor U9355 (N_9355,N_9221,N_9245);
nor U9356 (N_9356,N_9246,N_9278);
or U9357 (N_9357,N_9236,N_9169);
xnor U9358 (N_9358,N_9273,N_9231);
nor U9359 (N_9359,N_9282,N_9150);
and U9360 (N_9360,N_9283,N_9223);
nand U9361 (N_9361,N_9170,N_9179);
xnor U9362 (N_9362,N_9263,N_9296);
nor U9363 (N_9363,N_9160,N_9151);
nand U9364 (N_9364,N_9172,N_9193);
and U9365 (N_9365,N_9247,N_9162);
xor U9366 (N_9366,N_9291,N_9289);
or U9367 (N_9367,N_9228,N_9268);
nand U9368 (N_9368,N_9199,N_9285);
nor U9369 (N_9369,N_9226,N_9203);
and U9370 (N_9370,N_9187,N_9177);
nand U9371 (N_9371,N_9284,N_9163);
nor U9372 (N_9372,N_9166,N_9220);
nor U9373 (N_9373,N_9233,N_9261);
nor U9374 (N_9374,N_9200,N_9265);
nand U9375 (N_9375,N_9160,N_9269);
nand U9376 (N_9376,N_9203,N_9261);
and U9377 (N_9377,N_9151,N_9255);
and U9378 (N_9378,N_9287,N_9156);
and U9379 (N_9379,N_9250,N_9298);
nand U9380 (N_9380,N_9159,N_9153);
and U9381 (N_9381,N_9185,N_9271);
nor U9382 (N_9382,N_9195,N_9229);
xor U9383 (N_9383,N_9290,N_9272);
nor U9384 (N_9384,N_9249,N_9257);
nand U9385 (N_9385,N_9168,N_9255);
nand U9386 (N_9386,N_9206,N_9271);
and U9387 (N_9387,N_9156,N_9210);
xor U9388 (N_9388,N_9191,N_9212);
and U9389 (N_9389,N_9167,N_9225);
nand U9390 (N_9390,N_9270,N_9223);
or U9391 (N_9391,N_9284,N_9291);
and U9392 (N_9392,N_9189,N_9287);
and U9393 (N_9393,N_9211,N_9161);
or U9394 (N_9394,N_9170,N_9174);
and U9395 (N_9395,N_9203,N_9217);
xor U9396 (N_9396,N_9240,N_9224);
and U9397 (N_9397,N_9202,N_9296);
and U9398 (N_9398,N_9246,N_9185);
nor U9399 (N_9399,N_9168,N_9215);
and U9400 (N_9400,N_9195,N_9227);
xnor U9401 (N_9401,N_9295,N_9187);
xor U9402 (N_9402,N_9165,N_9160);
or U9403 (N_9403,N_9272,N_9209);
and U9404 (N_9404,N_9216,N_9198);
and U9405 (N_9405,N_9277,N_9289);
or U9406 (N_9406,N_9200,N_9238);
and U9407 (N_9407,N_9233,N_9189);
or U9408 (N_9408,N_9211,N_9208);
nor U9409 (N_9409,N_9159,N_9246);
or U9410 (N_9410,N_9271,N_9181);
xnor U9411 (N_9411,N_9279,N_9265);
nand U9412 (N_9412,N_9164,N_9283);
nand U9413 (N_9413,N_9280,N_9191);
xnor U9414 (N_9414,N_9197,N_9216);
nand U9415 (N_9415,N_9286,N_9194);
nand U9416 (N_9416,N_9170,N_9233);
or U9417 (N_9417,N_9191,N_9214);
or U9418 (N_9418,N_9180,N_9280);
or U9419 (N_9419,N_9277,N_9216);
nand U9420 (N_9420,N_9256,N_9241);
and U9421 (N_9421,N_9233,N_9238);
nand U9422 (N_9422,N_9199,N_9179);
xnor U9423 (N_9423,N_9161,N_9264);
xnor U9424 (N_9424,N_9194,N_9156);
or U9425 (N_9425,N_9151,N_9172);
nand U9426 (N_9426,N_9155,N_9270);
xor U9427 (N_9427,N_9237,N_9291);
nand U9428 (N_9428,N_9161,N_9250);
or U9429 (N_9429,N_9208,N_9284);
nand U9430 (N_9430,N_9166,N_9245);
or U9431 (N_9431,N_9266,N_9295);
xor U9432 (N_9432,N_9152,N_9286);
and U9433 (N_9433,N_9258,N_9172);
nand U9434 (N_9434,N_9230,N_9255);
and U9435 (N_9435,N_9209,N_9218);
or U9436 (N_9436,N_9234,N_9165);
xnor U9437 (N_9437,N_9265,N_9163);
and U9438 (N_9438,N_9233,N_9282);
xnor U9439 (N_9439,N_9292,N_9239);
nor U9440 (N_9440,N_9150,N_9166);
nor U9441 (N_9441,N_9172,N_9208);
or U9442 (N_9442,N_9183,N_9167);
xor U9443 (N_9443,N_9169,N_9221);
xor U9444 (N_9444,N_9198,N_9179);
and U9445 (N_9445,N_9152,N_9243);
nand U9446 (N_9446,N_9199,N_9188);
and U9447 (N_9447,N_9262,N_9253);
nor U9448 (N_9448,N_9275,N_9170);
nand U9449 (N_9449,N_9268,N_9160);
or U9450 (N_9450,N_9323,N_9427);
nor U9451 (N_9451,N_9348,N_9417);
nor U9452 (N_9452,N_9368,N_9446);
nor U9453 (N_9453,N_9349,N_9445);
or U9454 (N_9454,N_9424,N_9364);
nand U9455 (N_9455,N_9377,N_9301);
and U9456 (N_9456,N_9360,N_9322);
xnor U9457 (N_9457,N_9400,N_9350);
nand U9458 (N_9458,N_9394,N_9341);
nand U9459 (N_9459,N_9318,N_9371);
or U9460 (N_9460,N_9311,N_9395);
or U9461 (N_9461,N_9392,N_9338);
nand U9462 (N_9462,N_9387,N_9403);
or U9463 (N_9463,N_9447,N_9416);
nor U9464 (N_9464,N_9367,N_9372);
and U9465 (N_9465,N_9378,N_9342);
or U9466 (N_9466,N_9406,N_9327);
xnor U9467 (N_9467,N_9428,N_9331);
nand U9468 (N_9468,N_9354,N_9319);
and U9469 (N_9469,N_9330,N_9315);
and U9470 (N_9470,N_9312,N_9382);
nor U9471 (N_9471,N_9441,N_9356);
nor U9472 (N_9472,N_9423,N_9429);
xor U9473 (N_9473,N_9376,N_9399);
and U9474 (N_9474,N_9418,N_9339);
or U9475 (N_9475,N_9410,N_9389);
and U9476 (N_9476,N_9321,N_9449);
nand U9477 (N_9477,N_9381,N_9317);
and U9478 (N_9478,N_9396,N_9326);
xnor U9479 (N_9479,N_9357,N_9363);
and U9480 (N_9480,N_9359,N_9352);
nand U9481 (N_9481,N_9370,N_9383);
nand U9482 (N_9482,N_9422,N_9329);
nand U9483 (N_9483,N_9347,N_9306);
nand U9484 (N_9484,N_9385,N_9436);
nor U9485 (N_9485,N_9309,N_9369);
nand U9486 (N_9486,N_9358,N_9345);
nand U9487 (N_9487,N_9413,N_9365);
nor U9488 (N_9488,N_9425,N_9307);
xor U9489 (N_9489,N_9375,N_9435);
or U9490 (N_9490,N_9430,N_9334);
nor U9491 (N_9491,N_9304,N_9398);
xor U9492 (N_9492,N_9366,N_9373);
xnor U9493 (N_9493,N_9407,N_9397);
xor U9494 (N_9494,N_9439,N_9346);
xnor U9495 (N_9495,N_9391,N_9421);
nand U9496 (N_9496,N_9444,N_9401);
xnor U9497 (N_9497,N_9316,N_9328);
or U9498 (N_9498,N_9303,N_9332);
nor U9499 (N_9499,N_9443,N_9340);
or U9500 (N_9500,N_9414,N_9390);
xnor U9501 (N_9501,N_9343,N_9379);
nand U9502 (N_9502,N_9305,N_9412);
and U9503 (N_9503,N_9415,N_9336);
nor U9504 (N_9504,N_9393,N_9448);
xnor U9505 (N_9505,N_9344,N_9437);
or U9506 (N_9506,N_9337,N_9431);
xnor U9507 (N_9507,N_9335,N_9310);
and U9508 (N_9508,N_9300,N_9442);
and U9509 (N_9509,N_9333,N_9432);
xor U9510 (N_9510,N_9433,N_9409);
nor U9511 (N_9511,N_9434,N_9420);
nor U9512 (N_9512,N_9362,N_9384);
nand U9513 (N_9513,N_9405,N_9353);
and U9514 (N_9514,N_9426,N_9314);
nor U9515 (N_9515,N_9411,N_9374);
and U9516 (N_9516,N_9313,N_9351);
nor U9517 (N_9517,N_9308,N_9402);
xor U9518 (N_9518,N_9386,N_9404);
or U9519 (N_9519,N_9438,N_9388);
xor U9520 (N_9520,N_9380,N_9355);
nor U9521 (N_9521,N_9408,N_9361);
and U9522 (N_9522,N_9440,N_9419);
or U9523 (N_9523,N_9325,N_9302);
nand U9524 (N_9524,N_9320,N_9324);
and U9525 (N_9525,N_9369,N_9304);
nand U9526 (N_9526,N_9326,N_9337);
nand U9527 (N_9527,N_9362,N_9342);
nor U9528 (N_9528,N_9377,N_9326);
or U9529 (N_9529,N_9415,N_9337);
nor U9530 (N_9530,N_9364,N_9302);
nor U9531 (N_9531,N_9302,N_9332);
xor U9532 (N_9532,N_9401,N_9402);
and U9533 (N_9533,N_9374,N_9377);
nor U9534 (N_9534,N_9383,N_9417);
and U9535 (N_9535,N_9345,N_9405);
nand U9536 (N_9536,N_9399,N_9365);
or U9537 (N_9537,N_9305,N_9433);
xnor U9538 (N_9538,N_9418,N_9317);
xnor U9539 (N_9539,N_9344,N_9343);
nand U9540 (N_9540,N_9390,N_9417);
and U9541 (N_9541,N_9436,N_9394);
and U9542 (N_9542,N_9377,N_9380);
or U9543 (N_9543,N_9325,N_9394);
or U9544 (N_9544,N_9329,N_9435);
nand U9545 (N_9545,N_9384,N_9370);
and U9546 (N_9546,N_9309,N_9400);
nand U9547 (N_9547,N_9314,N_9447);
nor U9548 (N_9548,N_9420,N_9357);
nand U9549 (N_9549,N_9398,N_9438);
xor U9550 (N_9550,N_9348,N_9442);
xor U9551 (N_9551,N_9371,N_9303);
and U9552 (N_9552,N_9325,N_9411);
nand U9553 (N_9553,N_9441,N_9401);
and U9554 (N_9554,N_9436,N_9313);
xor U9555 (N_9555,N_9301,N_9448);
nand U9556 (N_9556,N_9310,N_9370);
xor U9557 (N_9557,N_9392,N_9448);
nor U9558 (N_9558,N_9317,N_9328);
nand U9559 (N_9559,N_9300,N_9347);
nor U9560 (N_9560,N_9309,N_9361);
nand U9561 (N_9561,N_9444,N_9356);
xor U9562 (N_9562,N_9444,N_9437);
and U9563 (N_9563,N_9367,N_9349);
or U9564 (N_9564,N_9426,N_9422);
and U9565 (N_9565,N_9405,N_9416);
and U9566 (N_9566,N_9338,N_9352);
xor U9567 (N_9567,N_9330,N_9393);
nor U9568 (N_9568,N_9362,N_9302);
xor U9569 (N_9569,N_9353,N_9426);
or U9570 (N_9570,N_9379,N_9414);
nor U9571 (N_9571,N_9320,N_9434);
nor U9572 (N_9572,N_9303,N_9437);
and U9573 (N_9573,N_9445,N_9420);
nor U9574 (N_9574,N_9346,N_9341);
or U9575 (N_9575,N_9414,N_9371);
xnor U9576 (N_9576,N_9327,N_9343);
xnor U9577 (N_9577,N_9353,N_9302);
and U9578 (N_9578,N_9395,N_9394);
or U9579 (N_9579,N_9426,N_9360);
xnor U9580 (N_9580,N_9388,N_9334);
xnor U9581 (N_9581,N_9371,N_9388);
and U9582 (N_9582,N_9358,N_9331);
and U9583 (N_9583,N_9399,N_9406);
nor U9584 (N_9584,N_9332,N_9380);
xor U9585 (N_9585,N_9417,N_9434);
or U9586 (N_9586,N_9444,N_9406);
or U9587 (N_9587,N_9415,N_9306);
nand U9588 (N_9588,N_9333,N_9328);
nand U9589 (N_9589,N_9419,N_9338);
nor U9590 (N_9590,N_9300,N_9305);
or U9591 (N_9591,N_9362,N_9358);
and U9592 (N_9592,N_9320,N_9398);
nor U9593 (N_9593,N_9437,N_9394);
or U9594 (N_9594,N_9318,N_9301);
nor U9595 (N_9595,N_9321,N_9339);
or U9596 (N_9596,N_9346,N_9405);
nor U9597 (N_9597,N_9412,N_9313);
nor U9598 (N_9598,N_9420,N_9406);
nor U9599 (N_9599,N_9398,N_9436);
xor U9600 (N_9600,N_9528,N_9565);
nor U9601 (N_9601,N_9457,N_9476);
nand U9602 (N_9602,N_9500,N_9548);
nand U9603 (N_9603,N_9566,N_9470);
or U9604 (N_9604,N_9533,N_9555);
or U9605 (N_9605,N_9468,N_9502);
nand U9606 (N_9606,N_9567,N_9556);
xnor U9607 (N_9607,N_9462,N_9524);
xnor U9608 (N_9608,N_9529,N_9450);
xor U9609 (N_9609,N_9597,N_9586);
and U9610 (N_9610,N_9509,N_9577);
xnor U9611 (N_9611,N_9497,N_9552);
nand U9612 (N_9612,N_9550,N_9564);
or U9613 (N_9613,N_9543,N_9482);
nor U9614 (N_9614,N_9491,N_9569);
or U9615 (N_9615,N_9469,N_9558);
and U9616 (N_9616,N_9467,N_9589);
or U9617 (N_9617,N_9455,N_9584);
xnor U9618 (N_9618,N_9553,N_9537);
xnor U9619 (N_9619,N_9477,N_9525);
or U9620 (N_9620,N_9501,N_9576);
xor U9621 (N_9621,N_9554,N_9512);
xor U9622 (N_9622,N_9514,N_9560);
nor U9623 (N_9623,N_9474,N_9459);
xor U9624 (N_9624,N_9588,N_9563);
nor U9625 (N_9625,N_9575,N_9580);
or U9626 (N_9626,N_9545,N_9594);
and U9627 (N_9627,N_9549,N_9510);
nand U9628 (N_9628,N_9458,N_9583);
or U9629 (N_9629,N_9492,N_9522);
nand U9630 (N_9630,N_9520,N_9538);
or U9631 (N_9631,N_9519,N_9488);
nand U9632 (N_9632,N_9456,N_9475);
or U9633 (N_9633,N_9485,N_9504);
and U9634 (N_9634,N_9534,N_9572);
xnor U9635 (N_9635,N_9591,N_9532);
or U9636 (N_9636,N_9489,N_9570);
nand U9637 (N_9637,N_9503,N_9511);
xor U9638 (N_9638,N_9579,N_9581);
nand U9639 (N_9639,N_9466,N_9465);
xor U9640 (N_9640,N_9516,N_9592);
and U9641 (N_9641,N_9513,N_9506);
nand U9642 (N_9642,N_9486,N_9453);
nand U9643 (N_9643,N_9578,N_9562);
xnor U9644 (N_9644,N_9451,N_9490);
nor U9645 (N_9645,N_9593,N_9493);
nor U9646 (N_9646,N_9582,N_9471);
nor U9647 (N_9647,N_9452,N_9541);
nor U9648 (N_9648,N_9527,N_9483);
nand U9649 (N_9649,N_9463,N_9517);
xnor U9650 (N_9650,N_9515,N_9599);
nand U9651 (N_9651,N_9590,N_9568);
xnor U9652 (N_9652,N_9546,N_9461);
nand U9653 (N_9653,N_9526,N_9505);
xnor U9654 (N_9654,N_9571,N_9596);
nor U9655 (N_9655,N_9454,N_9508);
or U9656 (N_9656,N_9460,N_9507);
and U9657 (N_9657,N_9540,N_9535);
nor U9658 (N_9658,N_9585,N_9587);
and U9659 (N_9659,N_9478,N_9495);
xnor U9660 (N_9660,N_9536,N_9598);
xnor U9661 (N_9661,N_9473,N_9530);
nand U9662 (N_9662,N_9547,N_9498);
nand U9663 (N_9663,N_9573,N_9484);
and U9664 (N_9664,N_9464,N_9595);
xnor U9665 (N_9665,N_9494,N_9539);
and U9666 (N_9666,N_9542,N_9531);
and U9667 (N_9667,N_9574,N_9496);
or U9668 (N_9668,N_9518,N_9481);
xor U9669 (N_9669,N_9557,N_9472);
and U9670 (N_9670,N_9559,N_9544);
nand U9671 (N_9671,N_9480,N_9479);
and U9672 (N_9672,N_9561,N_9551);
nor U9673 (N_9673,N_9521,N_9523);
or U9674 (N_9674,N_9487,N_9499);
and U9675 (N_9675,N_9476,N_9588);
or U9676 (N_9676,N_9452,N_9583);
nor U9677 (N_9677,N_9518,N_9521);
xor U9678 (N_9678,N_9524,N_9503);
nand U9679 (N_9679,N_9528,N_9495);
and U9680 (N_9680,N_9477,N_9502);
or U9681 (N_9681,N_9502,N_9575);
nor U9682 (N_9682,N_9546,N_9476);
or U9683 (N_9683,N_9504,N_9479);
xor U9684 (N_9684,N_9467,N_9487);
and U9685 (N_9685,N_9500,N_9466);
nand U9686 (N_9686,N_9538,N_9584);
or U9687 (N_9687,N_9458,N_9494);
nor U9688 (N_9688,N_9553,N_9558);
xnor U9689 (N_9689,N_9505,N_9479);
xor U9690 (N_9690,N_9519,N_9483);
nor U9691 (N_9691,N_9566,N_9568);
nand U9692 (N_9692,N_9504,N_9490);
xor U9693 (N_9693,N_9494,N_9544);
nor U9694 (N_9694,N_9494,N_9457);
xnor U9695 (N_9695,N_9559,N_9518);
xnor U9696 (N_9696,N_9467,N_9452);
and U9697 (N_9697,N_9480,N_9567);
and U9698 (N_9698,N_9483,N_9518);
nand U9699 (N_9699,N_9589,N_9477);
xor U9700 (N_9700,N_9577,N_9454);
nand U9701 (N_9701,N_9540,N_9545);
or U9702 (N_9702,N_9477,N_9493);
nor U9703 (N_9703,N_9514,N_9482);
nor U9704 (N_9704,N_9490,N_9531);
and U9705 (N_9705,N_9587,N_9506);
and U9706 (N_9706,N_9504,N_9458);
and U9707 (N_9707,N_9599,N_9474);
nor U9708 (N_9708,N_9453,N_9467);
nor U9709 (N_9709,N_9568,N_9464);
and U9710 (N_9710,N_9477,N_9558);
nor U9711 (N_9711,N_9534,N_9558);
and U9712 (N_9712,N_9553,N_9571);
or U9713 (N_9713,N_9557,N_9480);
and U9714 (N_9714,N_9549,N_9588);
xnor U9715 (N_9715,N_9517,N_9534);
nand U9716 (N_9716,N_9538,N_9555);
nor U9717 (N_9717,N_9516,N_9547);
and U9718 (N_9718,N_9558,N_9597);
xnor U9719 (N_9719,N_9479,N_9467);
and U9720 (N_9720,N_9574,N_9516);
xor U9721 (N_9721,N_9564,N_9593);
xor U9722 (N_9722,N_9509,N_9517);
and U9723 (N_9723,N_9460,N_9493);
nor U9724 (N_9724,N_9484,N_9561);
xnor U9725 (N_9725,N_9587,N_9511);
nand U9726 (N_9726,N_9545,N_9482);
nand U9727 (N_9727,N_9553,N_9459);
or U9728 (N_9728,N_9456,N_9482);
and U9729 (N_9729,N_9471,N_9588);
xnor U9730 (N_9730,N_9576,N_9580);
xnor U9731 (N_9731,N_9544,N_9531);
and U9732 (N_9732,N_9597,N_9458);
or U9733 (N_9733,N_9549,N_9570);
nor U9734 (N_9734,N_9550,N_9584);
or U9735 (N_9735,N_9533,N_9586);
nor U9736 (N_9736,N_9538,N_9470);
xnor U9737 (N_9737,N_9496,N_9461);
xor U9738 (N_9738,N_9560,N_9588);
nor U9739 (N_9739,N_9548,N_9541);
and U9740 (N_9740,N_9502,N_9499);
and U9741 (N_9741,N_9493,N_9598);
nand U9742 (N_9742,N_9542,N_9451);
xnor U9743 (N_9743,N_9460,N_9566);
and U9744 (N_9744,N_9496,N_9531);
nand U9745 (N_9745,N_9462,N_9479);
xor U9746 (N_9746,N_9563,N_9464);
xnor U9747 (N_9747,N_9490,N_9478);
nor U9748 (N_9748,N_9451,N_9504);
or U9749 (N_9749,N_9477,N_9522);
and U9750 (N_9750,N_9723,N_9651);
nor U9751 (N_9751,N_9652,N_9607);
nor U9752 (N_9752,N_9688,N_9636);
xor U9753 (N_9753,N_9670,N_9693);
nor U9754 (N_9754,N_9653,N_9635);
and U9755 (N_9755,N_9620,N_9738);
and U9756 (N_9756,N_9601,N_9669);
and U9757 (N_9757,N_9708,N_9608);
and U9758 (N_9758,N_9614,N_9659);
nor U9759 (N_9759,N_9641,N_9679);
nor U9760 (N_9760,N_9638,N_9649);
nand U9761 (N_9761,N_9713,N_9703);
or U9762 (N_9762,N_9694,N_9735);
nand U9763 (N_9763,N_9700,N_9705);
nand U9764 (N_9764,N_9710,N_9663);
nor U9765 (N_9765,N_9648,N_9678);
nor U9766 (N_9766,N_9642,N_9732);
and U9767 (N_9767,N_9695,N_9685);
or U9768 (N_9768,N_9615,N_9644);
or U9769 (N_9769,N_9726,N_9677);
or U9770 (N_9770,N_9704,N_9633);
nand U9771 (N_9771,N_9602,N_9668);
or U9772 (N_9772,N_9740,N_9680);
and U9773 (N_9773,N_9603,N_9697);
and U9774 (N_9774,N_9600,N_9686);
nor U9775 (N_9775,N_9718,N_9637);
and U9776 (N_9776,N_9717,N_9661);
nand U9777 (N_9777,N_9617,N_9682);
nand U9778 (N_9778,N_9746,N_9736);
nand U9779 (N_9779,N_9612,N_9743);
xor U9780 (N_9780,N_9640,N_9737);
nand U9781 (N_9781,N_9674,N_9673);
or U9782 (N_9782,N_9654,N_9714);
xnor U9783 (N_9783,N_9622,N_9698);
and U9784 (N_9784,N_9631,N_9739);
nand U9785 (N_9785,N_9684,N_9645);
nor U9786 (N_9786,N_9627,N_9683);
or U9787 (N_9787,N_9619,N_9747);
or U9788 (N_9788,N_9616,N_9702);
and U9789 (N_9789,N_9691,N_9634);
xnor U9790 (N_9790,N_9629,N_9662);
or U9791 (N_9791,N_9676,N_9625);
nor U9792 (N_9792,N_9742,N_9639);
nand U9793 (N_9793,N_9647,N_9630);
xor U9794 (N_9794,N_9722,N_9613);
nor U9795 (N_9795,N_9675,N_9727);
and U9796 (N_9796,N_9719,N_9658);
nand U9797 (N_9797,N_9660,N_9626);
xor U9798 (N_9798,N_9699,N_9650);
nor U9799 (N_9799,N_9707,N_9715);
xor U9800 (N_9800,N_9621,N_9748);
and U9801 (N_9801,N_9604,N_9655);
or U9802 (N_9802,N_9706,N_9701);
xor U9803 (N_9803,N_9712,N_9730);
xnor U9804 (N_9804,N_9672,N_9716);
or U9805 (N_9805,N_9696,N_9656);
nor U9806 (N_9806,N_9610,N_9728);
nand U9807 (N_9807,N_9643,N_9709);
xor U9808 (N_9808,N_9720,N_9744);
nor U9809 (N_9809,N_9731,N_9646);
nor U9810 (N_9810,N_9671,N_9618);
or U9811 (N_9811,N_9657,N_9690);
nor U9812 (N_9812,N_9749,N_9687);
nor U9813 (N_9813,N_9606,N_9689);
or U9814 (N_9814,N_9628,N_9605);
nor U9815 (N_9815,N_9733,N_9711);
or U9816 (N_9816,N_9692,N_9721);
nor U9817 (N_9817,N_9632,N_9741);
xnor U9818 (N_9818,N_9667,N_9729);
and U9819 (N_9819,N_9609,N_9664);
or U9820 (N_9820,N_9724,N_9665);
nor U9821 (N_9821,N_9745,N_9624);
nor U9822 (N_9822,N_9666,N_9681);
or U9823 (N_9823,N_9611,N_9725);
and U9824 (N_9824,N_9734,N_9623);
nor U9825 (N_9825,N_9677,N_9657);
or U9826 (N_9826,N_9716,N_9654);
or U9827 (N_9827,N_9667,N_9693);
or U9828 (N_9828,N_9732,N_9631);
xor U9829 (N_9829,N_9712,N_9641);
and U9830 (N_9830,N_9666,N_9642);
nor U9831 (N_9831,N_9692,N_9676);
and U9832 (N_9832,N_9739,N_9614);
or U9833 (N_9833,N_9713,N_9684);
nor U9834 (N_9834,N_9650,N_9673);
nor U9835 (N_9835,N_9688,N_9737);
or U9836 (N_9836,N_9659,N_9630);
xnor U9837 (N_9837,N_9660,N_9743);
nor U9838 (N_9838,N_9746,N_9743);
nor U9839 (N_9839,N_9614,N_9634);
nor U9840 (N_9840,N_9647,N_9671);
and U9841 (N_9841,N_9641,N_9618);
nand U9842 (N_9842,N_9615,N_9718);
xor U9843 (N_9843,N_9727,N_9604);
nand U9844 (N_9844,N_9654,N_9640);
nand U9845 (N_9845,N_9731,N_9664);
nor U9846 (N_9846,N_9643,N_9620);
nand U9847 (N_9847,N_9639,N_9611);
xor U9848 (N_9848,N_9647,N_9605);
xor U9849 (N_9849,N_9717,N_9707);
xnor U9850 (N_9850,N_9705,N_9704);
nand U9851 (N_9851,N_9677,N_9670);
or U9852 (N_9852,N_9653,N_9707);
or U9853 (N_9853,N_9696,N_9677);
nand U9854 (N_9854,N_9704,N_9747);
nor U9855 (N_9855,N_9667,N_9696);
and U9856 (N_9856,N_9668,N_9698);
xnor U9857 (N_9857,N_9647,N_9633);
and U9858 (N_9858,N_9689,N_9724);
nand U9859 (N_9859,N_9720,N_9701);
nand U9860 (N_9860,N_9707,N_9683);
nor U9861 (N_9861,N_9733,N_9700);
and U9862 (N_9862,N_9646,N_9706);
nor U9863 (N_9863,N_9609,N_9630);
and U9864 (N_9864,N_9649,N_9606);
xnor U9865 (N_9865,N_9604,N_9651);
nand U9866 (N_9866,N_9654,N_9649);
xor U9867 (N_9867,N_9748,N_9710);
nand U9868 (N_9868,N_9748,N_9677);
xnor U9869 (N_9869,N_9623,N_9747);
xor U9870 (N_9870,N_9744,N_9739);
nor U9871 (N_9871,N_9691,N_9734);
nand U9872 (N_9872,N_9633,N_9733);
xor U9873 (N_9873,N_9612,N_9697);
and U9874 (N_9874,N_9695,N_9601);
nand U9875 (N_9875,N_9641,N_9690);
and U9876 (N_9876,N_9680,N_9749);
xor U9877 (N_9877,N_9739,N_9671);
xnor U9878 (N_9878,N_9688,N_9662);
nand U9879 (N_9879,N_9686,N_9610);
nor U9880 (N_9880,N_9692,N_9713);
nand U9881 (N_9881,N_9748,N_9723);
or U9882 (N_9882,N_9698,N_9601);
xor U9883 (N_9883,N_9632,N_9713);
nand U9884 (N_9884,N_9613,N_9689);
nor U9885 (N_9885,N_9652,N_9737);
and U9886 (N_9886,N_9717,N_9716);
xnor U9887 (N_9887,N_9664,N_9628);
and U9888 (N_9888,N_9654,N_9661);
xnor U9889 (N_9889,N_9709,N_9675);
or U9890 (N_9890,N_9624,N_9635);
nor U9891 (N_9891,N_9709,N_9625);
nand U9892 (N_9892,N_9676,N_9706);
nor U9893 (N_9893,N_9687,N_9736);
and U9894 (N_9894,N_9737,N_9707);
and U9895 (N_9895,N_9620,N_9626);
and U9896 (N_9896,N_9632,N_9688);
nand U9897 (N_9897,N_9660,N_9698);
and U9898 (N_9898,N_9611,N_9709);
or U9899 (N_9899,N_9699,N_9731);
nand U9900 (N_9900,N_9766,N_9875);
and U9901 (N_9901,N_9860,N_9898);
and U9902 (N_9902,N_9757,N_9897);
or U9903 (N_9903,N_9823,N_9861);
or U9904 (N_9904,N_9863,N_9758);
or U9905 (N_9905,N_9792,N_9856);
or U9906 (N_9906,N_9770,N_9873);
nand U9907 (N_9907,N_9824,N_9814);
and U9908 (N_9908,N_9879,N_9815);
or U9909 (N_9909,N_9869,N_9852);
nor U9910 (N_9910,N_9849,N_9759);
xnor U9911 (N_9911,N_9878,N_9831);
nor U9912 (N_9912,N_9891,N_9884);
nand U9913 (N_9913,N_9754,N_9877);
xor U9914 (N_9914,N_9840,N_9843);
nand U9915 (N_9915,N_9780,N_9858);
nand U9916 (N_9916,N_9881,N_9805);
nand U9917 (N_9917,N_9756,N_9802);
or U9918 (N_9918,N_9784,N_9787);
xor U9919 (N_9919,N_9779,N_9774);
xor U9920 (N_9920,N_9791,N_9855);
or U9921 (N_9921,N_9876,N_9767);
or U9922 (N_9922,N_9854,N_9888);
nor U9923 (N_9923,N_9887,N_9896);
nand U9924 (N_9924,N_9859,N_9844);
and U9925 (N_9925,N_9867,N_9837);
nor U9926 (N_9926,N_9872,N_9786);
nor U9927 (N_9927,N_9807,N_9769);
or U9928 (N_9928,N_9795,N_9817);
or U9929 (N_9929,N_9781,N_9800);
and U9930 (N_9930,N_9808,N_9776);
or U9931 (N_9931,N_9882,N_9894);
and U9932 (N_9932,N_9773,N_9793);
nor U9933 (N_9933,N_9827,N_9760);
nor U9934 (N_9934,N_9783,N_9847);
or U9935 (N_9935,N_9771,N_9803);
nand U9936 (N_9936,N_9857,N_9842);
and U9937 (N_9937,N_9864,N_9886);
nand U9938 (N_9938,N_9789,N_9868);
and U9939 (N_9939,N_9790,N_9865);
nand U9940 (N_9940,N_9895,N_9763);
nand U9941 (N_9941,N_9853,N_9755);
xnor U9942 (N_9942,N_9889,N_9753);
nand U9943 (N_9943,N_9841,N_9832);
xor U9944 (N_9944,N_9830,N_9777);
xnor U9945 (N_9945,N_9833,N_9821);
or U9946 (N_9946,N_9871,N_9838);
nand U9947 (N_9947,N_9778,N_9835);
and U9948 (N_9948,N_9829,N_9870);
nand U9949 (N_9949,N_9883,N_9874);
nor U9950 (N_9950,N_9797,N_9846);
nand U9951 (N_9951,N_9813,N_9806);
or U9952 (N_9952,N_9862,N_9765);
nor U9953 (N_9953,N_9866,N_9839);
nand U9954 (N_9954,N_9768,N_9880);
and U9955 (N_9955,N_9822,N_9785);
xor U9956 (N_9956,N_9850,N_9750);
or U9957 (N_9957,N_9751,N_9818);
nor U9958 (N_9958,N_9834,N_9812);
or U9959 (N_9959,N_9845,N_9890);
nand U9960 (N_9960,N_9819,N_9836);
nor U9961 (N_9961,N_9892,N_9825);
xnor U9962 (N_9962,N_9764,N_9798);
or U9963 (N_9963,N_9801,N_9804);
or U9964 (N_9964,N_9772,N_9796);
xnor U9965 (N_9965,N_9848,N_9820);
or U9966 (N_9966,N_9885,N_9828);
and U9967 (N_9967,N_9788,N_9809);
nor U9968 (N_9968,N_9799,N_9794);
xnor U9969 (N_9969,N_9811,N_9816);
and U9970 (N_9970,N_9851,N_9752);
or U9971 (N_9971,N_9899,N_9826);
and U9972 (N_9972,N_9775,N_9893);
and U9973 (N_9973,N_9761,N_9782);
nor U9974 (N_9974,N_9762,N_9810);
xnor U9975 (N_9975,N_9786,N_9895);
or U9976 (N_9976,N_9831,N_9829);
nand U9977 (N_9977,N_9786,N_9790);
nor U9978 (N_9978,N_9847,N_9897);
xnor U9979 (N_9979,N_9859,N_9808);
nor U9980 (N_9980,N_9770,N_9829);
or U9981 (N_9981,N_9841,N_9806);
nor U9982 (N_9982,N_9766,N_9814);
nor U9983 (N_9983,N_9887,N_9776);
xor U9984 (N_9984,N_9832,N_9807);
xor U9985 (N_9985,N_9868,N_9807);
nor U9986 (N_9986,N_9794,N_9779);
nor U9987 (N_9987,N_9794,N_9754);
nand U9988 (N_9988,N_9824,N_9755);
xnor U9989 (N_9989,N_9856,N_9852);
nor U9990 (N_9990,N_9788,N_9793);
and U9991 (N_9991,N_9884,N_9774);
nor U9992 (N_9992,N_9758,N_9765);
nor U9993 (N_9993,N_9803,N_9770);
or U9994 (N_9994,N_9843,N_9824);
nand U9995 (N_9995,N_9785,N_9781);
nor U9996 (N_9996,N_9885,N_9778);
nand U9997 (N_9997,N_9837,N_9808);
and U9998 (N_9998,N_9850,N_9848);
and U9999 (N_9999,N_9880,N_9861);
nand U10000 (N_10000,N_9803,N_9793);
xor U10001 (N_10001,N_9775,N_9774);
nand U10002 (N_10002,N_9764,N_9866);
nor U10003 (N_10003,N_9761,N_9836);
and U10004 (N_10004,N_9874,N_9781);
xnor U10005 (N_10005,N_9866,N_9755);
nand U10006 (N_10006,N_9787,N_9844);
nor U10007 (N_10007,N_9822,N_9779);
and U10008 (N_10008,N_9884,N_9869);
nand U10009 (N_10009,N_9823,N_9860);
or U10010 (N_10010,N_9850,N_9808);
nand U10011 (N_10011,N_9871,N_9759);
nand U10012 (N_10012,N_9838,N_9762);
or U10013 (N_10013,N_9807,N_9753);
nor U10014 (N_10014,N_9847,N_9786);
xnor U10015 (N_10015,N_9809,N_9863);
or U10016 (N_10016,N_9890,N_9820);
or U10017 (N_10017,N_9835,N_9791);
or U10018 (N_10018,N_9819,N_9803);
or U10019 (N_10019,N_9843,N_9781);
and U10020 (N_10020,N_9799,N_9838);
nor U10021 (N_10021,N_9847,N_9782);
nand U10022 (N_10022,N_9856,N_9782);
xor U10023 (N_10023,N_9835,N_9862);
and U10024 (N_10024,N_9853,N_9867);
and U10025 (N_10025,N_9760,N_9810);
xnor U10026 (N_10026,N_9754,N_9851);
and U10027 (N_10027,N_9826,N_9857);
xnor U10028 (N_10028,N_9761,N_9847);
or U10029 (N_10029,N_9848,N_9819);
nor U10030 (N_10030,N_9857,N_9822);
and U10031 (N_10031,N_9809,N_9751);
nand U10032 (N_10032,N_9770,N_9893);
nand U10033 (N_10033,N_9831,N_9888);
nand U10034 (N_10034,N_9795,N_9779);
or U10035 (N_10035,N_9789,N_9810);
nand U10036 (N_10036,N_9816,N_9753);
xnor U10037 (N_10037,N_9755,N_9780);
nor U10038 (N_10038,N_9825,N_9884);
and U10039 (N_10039,N_9878,N_9837);
nand U10040 (N_10040,N_9799,N_9866);
nor U10041 (N_10041,N_9888,N_9783);
and U10042 (N_10042,N_9766,N_9759);
and U10043 (N_10043,N_9857,N_9765);
nor U10044 (N_10044,N_9835,N_9853);
or U10045 (N_10045,N_9767,N_9750);
nand U10046 (N_10046,N_9829,N_9823);
nand U10047 (N_10047,N_9765,N_9808);
nor U10048 (N_10048,N_9812,N_9833);
and U10049 (N_10049,N_9894,N_9899);
nand U10050 (N_10050,N_9997,N_10028);
xnor U10051 (N_10051,N_9934,N_9910);
xor U10052 (N_10052,N_9999,N_10017);
and U10053 (N_10053,N_9954,N_10047);
nor U10054 (N_10054,N_10036,N_10012);
or U10055 (N_10055,N_9959,N_9928);
or U10056 (N_10056,N_9996,N_10044);
or U10057 (N_10057,N_10021,N_9968);
or U10058 (N_10058,N_9957,N_9964);
or U10059 (N_10059,N_9930,N_9940);
and U10060 (N_10060,N_9967,N_10015);
or U10061 (N_10061,N_9937,N_9914);
nand U10062 (N_10062,N_9931,N_10007);
or U10063 (N_10063,N_9933,N_10025);
nor U10064 (N_10064,N_9976,N_9960);
or U10065 (N_10065,N_9971,N_9925);
nor U10066 (N_10066,N_9991,N_9939);
nand U10067 (N_10067,N_10033,N_9920);
or U10068 (N_10068,N_9998,N_9949);
xor U10069 (N_10069,N_10030,N_10042);
nor U10070 (N_10070,N_9918,N_9944);
nor U10071 (N_10071,N_9919,N_9985);
nand U10072 (N_10072,N_10045,N_10038);
or U10073 (N_10073,N_10016,N_9982);
nand U10074 (N_10074,N_9978,N_9900);
xnor U10075 (N_10075,N_9915,N_10027);
nor U10076 (N_10076,N_9966,N_9921);
or U10077 (N_10077,N_10041,N_9961);
nor U10078 (N_10078,N_9977,N_9962);
nand U10079 (N_10079,N_10004,N_9973);
nand U10080 (N_10080,N_9947,N_10048);
and U10081 (N_10081,N_9917,N_10008);
and U10082 (N_10082,N_9984,N_10014);
and U10083 (N_10083,N_9926,N_9906);
nand U10084 (N_10084,N_10011,N_9943);
and U10085 (N_10085,N_9951,N_9938);
and U10086 (N_10086,N_9993,N_9990);
nor U10087 (N_10087,N_9948,N_9988);
nor U10088 (N_10088,N_9902,N_10018);
or U10089 (N_10089,N_10005,N_10040);
xnor U10090 (N_10090,N_9904,N_9994);
nor U10091 (N_10091,N_10000,N_9942);
xnor U10092 (N_10092,N_10039,N_10013);
nand U10093 (N_10093,N_9953,N_9979);
or U10094 (N_10094,N_9995,N_9956);
nor U10095 (N_10095,N_9935,N_9981);
or U10096 (N_10096,N_9965,N_10002);
xor U10097 (N_10097,N_10020,N_10003);
or U10098 (N_10098,N_9945,N_10029);
xor U10099 (N_10099,N_9989,N_9913);
nand U10100 (N_10100,N_9908,N_10006);
or U10101 (N_10101,N_10024,N_9983);
nand U10102 (N_10102,N_9987,N_9941);
nand U10103 (N_10103,N_9975,N_9924);
nor U10104 (N_10104,N_9909,N_9916);
nor U10105 (N_10105,N_9903,N_9912);
nand U10106 (N_10106,N_9972,N_9936);
nor U10107 (N_10107,N_10026,N_10031);
nand U10108 (N_10108,N_10046,N_10022);
nor U10109 (N_10109,N_10049,N_9974);
nor U10110 (N_10110,N_10034,N_10001);
xor U10111 (N_10111,N_9927,N_9932);
nor U10112 (N_10112,N_10035,N_10037);
nor U10113 (N_10113,N_10009,N_9950);
and U10114 (N_10114,N_10019,N_9955);
nand U10115 (N_10115,N_9922,N_9923);
xnor U10116 (N_10116,N_9980,N_10010);
nor U10117 (N_10117,N_9992,N_9963);
and U10118 (N_10118,N_9905,N_10043);
nand U10119 (N_10119,N_10023,N_9946);
xor U10120 (N_10120,N_10032,N_9907);
nand U10121 (N_10121,N_9969,N_9958);
or U10122 (N_10122,N_9901,N_9970);
or U10123 (N_10123,N_9952,N_9986);
and U10124 (N_10124,N_9911,N_9929);
or U10125 (N_10125,N_10001,N_9914);
or U10126 (N_10126,N_9966,N_9981);
or U10127 (N_10127,N_10001,N_10014);
and U10128 (N_10128,N_10035,N_9998);
or U10129 (N_10129,N_10025,N_9960);
nand U10130 (N_10130,N_9913,N_9946);
nand U10131 (N_10131,N_9996,N_9900);
and U10132 (N_10132,N_9945,N_9946);
or U10133 (N_10133,N_9955,N_10029);
nand U10134 (N_10134,N_10047,N_9965);
and U10135 (N_10135,N_10047,N_9956);
or U10136 (N_10136,N_9939,N_9999);
nor U10137 (N_10137,N_9983,N_9906);
or U10138 (N_10138,N_9987,N_10016);
xnor U10139 (N_10139,N_9924,N_10024);
xnor U10140 (N_10140,N_9961,N_10005);
or U10141 (N_10141,N_9942,N_10020);
xor U10142 (N_10142,N_9933,N_9906);
nand U10143 (N_10143,N_9956,N_9996);
nor U10144 (N_10144,N_9966,N_9904);
and U10145 (N_10145,N_9904,N_10009);
nand U10146 (N_10146,N_10016,N_10041);
or U10147 (N_10147,N_10002,N_10026);
and U10148 (N_10148,N_10000,N_9982);
or U10149 (N_10149,N_9927,N_10020);
nor U10150 (N_10150,N_9961,N_9922);
xor U10151 (N_10151,N_9921,N_9902);
or U10152 (N_10152,N_10029,N_10032);
nor U10153 (N_10153,N_9955,N_9981);
xnor U10154 (N_10154,N_10018,N_10001);
nor U10155 (N_10155,N_9910,N_9950);
nor U10156 (N_10156,N_9948,N_10032);
nand U10157 (N_10157,N_10029,N_9962);
nor U10158 (N_10158,N_9902,N_9906);
xnor U10159 (N_10159,N_9914,N_10039);
nor U10160 (N_10160,N_9979,N_9985);
or U10161 (N_10161,N_9959,N_9996);
nor U10162 (N_10162,N_9926,N_9955);
and U10163 (N_10163,N_9982,N_9947);
xnor U10164 (N_10164,N_9920,N_9942);
xor U10165 (N_10165,N_9901,N_10004);
nand U10166 (N_10166,N_9994,N_9972);
or U10167 (N_10167,N_10040,N_10048);
nor U10168 (N_10168,N_9974,N_9966);
xnor U10169 (N_10169,N_9980,N_9913);
or U10170 (N_10170,N_9979,N_9911);
xor U10171 (N_10171,N_9965,N_10012);
and U10172 (N_10172,N_9963,N_10048);
xor U10173 (N_10173,N_10027,N_10030);
or U10174 (N_10174,N_10006,N_9900);
nor U10175 (N_10175,N_10021,N_9938);
nor U10176 (N_10176,N_9951,N_9917);
nor U10177 (N_10177,N_10035,N_10049);
xor U10178 (N_10178,N_9974,N_10023);
or U10179 (N_10179,N_9945,N_9915);
and U10180 (N_10180,N_9913,N_9909);
nor U10181 (N_10181,N_9986,N_10003);
xnor U10182 (N_10182,N_9998,N_10026);
nor U10183 (N_10183,N_9971,N_9930);
nor U10184 (N_10184,N_10005,N_9914);
or U10185 (N_10185,N_9941,N_9951);
nand U10186 (N_10186,N_9939,N_10001);
or U10187 (N_10187,N_10026,N_9947);
and U10188 (N_10188,N_10040,N_9948);
nor U10189 (N_10189,N_9946,N_9915);
and U10190 (N_10190,N_10019,N_9999);
xnor U10191 (N_10191,N_9917,N_9967);
and U10192 (N_10192,N_9946,N_9932);
xnor U10193 (N_10193,N_9956,N_9946);
nand U10194 (N_10194,N_9988,N_9957);
xnor U10195 (N_10195,N_9900,N_9975);
and U10196 (N_10196,N_10041,N_9913);
nand U10197 (N_10197,N_10038,N_9979);
nor U10198 (N_10198,N_9986,N_9969);
and U10199 (N_10199,N_9985,N_9984);
or U10200 (N_10200,N_10107,N_10118);
xnor U10201 (N_10201,N_10087,N_10144);
xor U10202 (N_10202,N_10154,N_10106);
xor U10203 (N_10203,N_10071,N_10089);
and U10204 (N_10204,N_10140,N_10193);
xor U10205 (N_10205,N_10053,N_10163);
nor U10206 (N_10206,N_10116,N_10103);
xnor U10207 (N_10207,N_10082,N_10079);
xor U10208 (N_10208,N_10156,N_10058);
or U10209 (N_10209,N_10196,N_10182);
and U10210 (N_10210,N_10179,N_10147);
nor U10211 (N_10211,N_10162,N_10199);
xor U10212 (N_10212,N_10148,N_10068);
or U10213 (N_10213,N_10158,N_10113);
xor U10214 (N_10214,N_10090,N_10096);
xnor U10215 (N_10215,N_10124,N_10115);
nand U10216 (N_10216,N_10074,N_10092);
and U10217 (N_10217,N_10131,N_10132);
xnor U10218 (N_10218,N_10095,N_10078);
nor U10219 (N_10219,N_10133,N_10129);
xnor U10220 (N_10220,N_10060,N_10143);
xnor U10221 (N_10221,N_10157,N_10167);
nand U10222 (N_10222,N_10072,N_10097);
and U10223 (N_10223,N_10141,N_10052);
xnor U10224 (N_10224,N_10159,N_10191);
nand U10225 (N_10225,N_10180,N_10102);
or U10226 (N_10226,N_10137,N_10139);
nand U10227 (N_10227,N_10146,N_10117);
nand U10228 (N_10228,N_10083,N_10105);
or U10229 (N_10229,N_10197,N_10055);
or U10230 (N_10230,N_10066,N_10084);
nand U10231 (N_10231,N_10069,N_10100);
or U10232 (N_10232,N_10099,N_10198);
nand U10233 (N_10233,N_10187,N_10150);
nor U10234 (N_10234,N_10057,N_10195);
nor U10235 (N_10235,N_10173,N_10086);
nand U10236 (N_10236,N_10127,N_10135);
nor U10237 (N_10237,N_10123,N_10171);
nor U10238 (N_10238,N_10153,N_10077);
nand U10239 (N_10239,N_10130,N_10142);
nand U10240 (N_10240,N_10166,N_10181);
nand U10241 (N_10241,N_10184,N_10194);
or U10242 (N_10242,N_10098,N_10093);
nor U10243 (N_10243,N_10059,N_10165);
xor U10244 (N_10244,N_10111,N_10178);
and U10245 (N_10245,N_10151,N_10172);
xor U10246 (N_10246,N_10149,N_10070);
or U10247 (N_10247,N_10091,N_10062);
xnor U10248 (N_10248,N_10122,N_10081);
or U10249 (N_10249,N_10168,N_10189);
and U10250 (N_10250,N_10112,N_10155);
xor U10251 (N_10251,N_10161,N_10186);
nand U10252 (N_10252,N_10119,N_10136);
and U10253 (N_10253,N_10160,N_10126);
nor U10254 (N_10254,N_10192,N_10050);
or U10255 (N_10255,N_10094,N_10114);
xnor U10256 (N_10256,N_10177,N_10067);
and U10257 (N_10257,N_10054,N_10170);
and U10258 (N_10258,N_10125,N_10185);
nand U10259 (N_10259,N_10088,N_10051);
nor U10260 (N_10260,N_10075,N_10164);
nor U10261 (N_10261,N_10080,N_10134);
nand U10262 (N_10262,N_10152,N_10175);
nand U10263 (N_10263,N_10128,N_10065);
or U10264 (N_10264,N_10085,N_10064);
nand U10265 (N_10265,N_10076,N_10145);
nor U10266 (N_10266,N_10061,N_10183);
and U10267 (N_10267,N_10190,N_10176);
nand U10268 (N_10268,N_10108,N_10138);
xnor U10269 (N_10269,N_10109,N_10104);
nor U10270 (N_10270,N_10101,N_10121);
and U10271 (N_10271,N_10188,N_10073);
and U10272 (N_10272,N_10120,N_10174);
and U10273 (N_10273,N_10063,N_10056);
or U10274 (N_10274,N_10110,N_10169);
xnor U10275 (N_10275,N_10174,N_10102);
nor U10276 (N_10276,N_10116,N_10162);
and U10277 (N_10277,N_10059,N_10109);
xnor U10278 (N_10278,N_10173,N_10093);
xor U10279 (N_10279,N_10111,N_10055);
or U10280 (N_10280,N_10070,N_10192);
xor U10281 (N_10281,N_10139,N_10085);
or U10282 (N_10282,N_10052,N_10188);
nor U10283 (N_10283,N_10174,N_10107);
and U10284 (N_10284,N_10130,N_10060);
and U10285 (N_10285,N_10172,N_10071);
nor U10286 (N_10286,N_10074,N_10088);
xor U10287 (N_10287,N_10122,N_10129);
nand U10288 (N_10288,N_10078,N_10076);
xnor U10289 (N_10289,N_10161,N_10053);
or U10290 (N_10290,N_10075,N_10138);
and U10291 (N_10291,N_10186,N_10078);
or U10292 (N_10292,N_10065,N_10076);
and U10293 (N_10293,N_10133,N_10184);
xnor U10294 (N_10294,N_10100,N_10192);
or U10295 (N_10295,N_10098,N_10105);
nor U10296 (N_10296,N_10167,N_10185);
nor U10297 (N_10297,N_10191,N_10105);
nand U10298 (N_10298,N_10110,N_10085);
nor U10299 (N_10299,N_10176,N_10098);
nand U10300 (N_10300,N_10118,N_10162);
and U10301 (N_10301,N_10063,N_10109);
nor U10302 (N_10302,N_10150,N_10066);
nor U10303 (N_10303,N_10123,N_10164);
or U10304 (N_10304,N_10198,N_10070);
nor U10305 (N_10305,N_10183,N_10159);
or U10306 (N_10306,N_10163,N_10153);
and U10307 (N_10307,N_10161,N_10051);
and U10308 (N_10308,N_10153,N_10117);
or U10309 (N_10309,N_10175,N_10129);
or U10310 (N_10310,N_10134,N_10161);
and U10311 (N_10311,N_10138,N_10137);
and U10312 (N_10312,N_10179,N_10089);
nor U10313 (N_10313,N_10100,N_10170);
or U10314 (N_10314,N_10086,N_10140);
or U10315 (N_10315,N_10099,N_10178);
xnor U10316 (N_10316,N_10176,N_10109);
xnor U10317 (N_10317,N_10177,N_10143);
nand U10318 (N_10318,N_10173,N_10051);
nor U10319 (N_10319,N_10167,N_10102);
and U10320 (N_10320,N_10172,N_10095);
xor U10321 (N_10321,N_10162,N_10166);
and U10322 (N_10322,N_10139,N_10171);
or U10323 (N_10323,N_10079,N_10199);
and U10324 (N_10324,N_10183,N_10086);
or U10325 (N_10325,N_10079,N_10089);
and U10326 (N_10326,N_10172,N_10150);
nor U10327 (N_10327,N_10097,N_10117);
nor U10328 (N_10328,N_10064,N_10058);
nor U10329 (N_10329,N_10107,N_10062);
and U10330 (N_10330,N_10159,N_10121);
nor U10331 (N_10331,N_10129,N_10142);
or U10332 (N_10332,N_10154,N_10108);
nand U10333 (N_10333,N_10170,N_10141);
xnor U10334 (N_10334,N_10100,N_10146);
nor U10335 (N_10335,N_10073,N_10177);
nor U10336 (N_10336,N_10176,N_10067);
xnor U10337 (N_10337,N_10126,N_10060);
xor U10338 (N_10338,N_10097,N_10124);
nor U10339 (N_10339,N_10193,N_10121);
xor U10340 (N_10340,N_10066,N_10143);
xnor U10341 (N_10341,N_10087,N_10171);
xor U10342 (N_10342,N_10094,N_10122);
nor U10343 (N_10343,N_10175,N_10119);
nor U10344 (N_10344,N_10197,N_10063);
xor U10345 (N_10345,N_10159,N_10087);
nand U10346 (N_10346,N_10053,N_10084);
or U10347 (N_10347,N_10157,N_10114);
nor U10348 (N_10348,N_10073,N_10133);
nor U10349 (N_10349,N_10076,N_10088);
and U10350 (N_10350,N_10225,N_10318);
xnor U10351 (N_10351,N_10287,N_10217);
or U10352 (N_10352,N_10305,N_10315);
or U10353 (N_10353,N_10300,N_10207);
and U10354 (N_10354,N_10321,N_10347);
nor U10355 (N_10355,N_10302,N_10303);
or U10356 (N_10356,N_10316,N_10340);
nor U10357 (N_10357,N_10270,N_10272);
or U10358 (N_10358,N_10249,N_10348);
or U10359 (N_10359,N_10343,N_10210);
or U10360 (N_10360,N_10329,N_10216);
and U10361 (N_10361,N_10241,N_10304);
xnor U10362 (N_10362,N_10232,N_10248);
and U10363 (N_10363,N_10332,N_10271);
nor U10364 (N_10364,N_10284,N_10201);
xor U10365 (N_10365,N_10220,N_10322);
and U10366 (N_10366,N_10238,N_10273);
or U10367 (N_10367,N_10280,N_10336);
nand U10368 (N_10368,N_10298,N_10215);
and U10369 (N_10369,N_10208,N_10247);
nor U10370 (N_10370,N_10267,N_10233);
nor U10371 (N_10371,N_10221,N_10345);
and U10372 (N_10372,N_10240,N_10263);
and U10373 (N_10373,N_10276,N_10229);
nand U10374 (N_10374,N_10330,N_10257);
nand U10375 (N_10375,N_10274,N_10289);
and U10376 (N_10376,N_10312,N_10282);
xor U10377 (N_10377,N_10224,N_10297);
and U10378 (N_10378,N_10211,N_10219);
and U10379 (N_10379,N_10236,N_10346);
nor U10380 (N_10380,N_10261,N_10251);
or U10381 (N_10381,N_10252,N_10325);
nand U10382 (N_10382,N_10254,N_10310);
and U10383 (N_10383,N_10231,N_10235);
nand U10384 (N_10384,N_10227,N_10306);
nand U10385 (N_10385,N_10292,N_10334);
xnor U10386 (N_10386,N_10327,N_10230);
or U10387 (N_10387,N_10202,N_10278);
or U10388 (N_10388,N_10319,N_10275);
nand U10389 (N_10389,N_10307,N_10222);
xnor U10390 (N_10390,N_10255,N_10212);
or U10391 (N_10391,N_10333,N_10344);
or U10392 (N_10392,N_10266,N_10311);
and U10393 (N_10393,N_10269,N_10301);
nor U10394 (N_10394,N_10286,N_10342);
and U10395 (N_10395,N_10242,N_10279);
nand U10396 (N_10396,N_10226,N_10244);
xnor U10397 (N_10397,N_10223,N_10313);
nand U10398 (N_10398,N_10314,N_10205);
nand U10399 (N_10399,N_10328,N_10228);
or U10400 (N_10400,N_10245,N_10326);
and U10401 (N_10401,N_10268,N_10237);
xnor U10402 (N_10402,N_10239,N_10213);
xor U10403 (N_10403,N_10335,N_10295);
and U10404 (N_10404,N_10324,N_10206);
xor U10405 (N_10405,N_10256,N_10323);
xnor U10406 (N_10406,N_10290,N_10259);
nor U10407 (N_10407,N_10294,N_10285);
nand U10408 (N_10408,N_10288,N_10299);
nor U10409 (N_10409,N_10296,N_10204);
nand U10410 (N_10410,N_10339,N_10293);
xnor U10411 (N_10411,N_10320,N_10264);
nand U10412 (N_10412,N_10331,N_10258);
xnor U10413 (N_10413,N_10277,N_10262);
nor U10414 (N_10414,N_10253,N_10341);
or U10415 (N_10415,N_10246,N_10291);
or U10416 (N_10416,N_10283,N_10218);
nor U10417 (N_10417,N_10203,N_10243);
and U10418 (N_10418,N_10214,N_10308);
nor U10419 (N_10419,N_10265,N_10349);
and U10420 (N_10420,N_10309,N_10200);
or U10421 (N_10421,N_10338,N_10234);
or U10422 (N_10422,N_10281,N_10260);
nand U10423 (N_10423,N_10337,N_10317);
xnor U10424 (N_10424,N_10209,N_10250);
xor U10425 (N_10425,N_10302,N_10305);
or U10426 (N_10426,N_10253,N_10239);
nor U10427 (N_10427,N_10237,N_10319);
or U10428 (N_10428,N_10224,N_10341);
and U10429 (N_10429,N_10293,N_10317);
nand U10430 (N_10430,N_10201,N_10347);
nand U10431 (N_10431,N_10253,N_10249);
nand U10432 (N_10432,N_10208,N_10309);
xor U10433 (N_10433,N_10264,N_10246);
nand U10434 (N_10434,N_10320,N_10211);
and U10435 (N_10435,N_10213,N_10346);
or U10436 (N_10436,N_10332,N_10206);
nor U10437 (N_10437,N_10289,N_10343);
or U10438 (N_10438,N_10317,N_10200);
xor U10439 (N_10439,N_10329,N_10286);
or U10440 (N_10440,N_10243,N_10271);
nor U10441 (N_10441,N_10230,N_10232);
xnor U10442 (N_10442,N_10252,N_10345);
nand U10443 (N_10443,N_10264,N_10301);
and U10444 (N_10444,N_10280,N_10242);
xnor U10445 (N_10445,N_10231,N_10344);
nand U10446 (N_10446,N_10285,N_10300);
nand U10447 (N_10447,N_10238,N_10228);
and U10448 (N_10448,N_10261,N_10243);
and U10449 (N_10449,N_10260,N_10207);
nor U10450 (N_10450,N_10285,N_10347);
and U10451 (N_10451,N_10325,N_10314);
and U10452 (N_10452,N_10343,N_10296);
nand U10453 (N_10453,N_10259,N_10251);
xor U10454 (N_10454,N_10260,N_10298);
or U10455 (N_10455,N_10308,N_10226);
nor U10456 (N_10456,N_10211,N_10249);
nand U10457 (N_10457,N_10299,N_10291);
xnor U10458 (N_10458,N_10301,N_10219);
xor U10459 (N_10459,N_10269,N_10335);
nand U10460 (N_10460,N_10206,N_10312);
nor U10461 (N_10461,N_10244,N_10268);
nor U10462 (N_10462,N_10319,N_10337);
or U10463 (N_10463,N_10307,N_10324);
nand U10464 (N_10464,N_10346,N_10275);
or U10465 (N_10465,N_10347,N_10301);
nand U10466 (N_10466,N_10262,N_10313);
and U10467 (N_10467,N_10242,N_10253);
nand U10468 (N_10468,N_10257,N_10249);
xnor U10469 (N_10469,N_10218,N_10232);
and U10470 (N_10470,N_10269,N_10298);
or U10471 (N_10471,N_10277,N_10204);
and U10472 (N_10472,N_10275,N_10215);
nor U10473 (N_10473,N_10316,N_10210);
xnor U10474 (N_10474,N_10217,N_10219);
nor U10475 (N_10475,N_10277,N_10247);
or U10476 (N_10476,N_10239,N_10293);
xor U10477 (N_10477,N_10347,N_10264);
and U10478 (N_10478,N_10213,N_10345);
or U10479 (N_10479,N_10339,N_10236);
nor U10480 (N_10480,N_10309,N_10243);
or U10481 (N_10481,N_10261,N_10252);
or U10482 (N_10482,N_10247,N_10242);
nand U10483 (N_10483,N_10298,N_10250);
or U10484 (N_10484,N_10221,N_10242);
and U10485 (N_10485,N_10349,N_10275);
or U10486 (N_10486,N_10332,N_10312);
nand U10487 (N_10487,N_10321,N_10212);
and U10488 (N_10488,N_10216,N_10293);
xor U10489 (N_10489,N_10317,N_10309);
and U10490 (N_10490,N_10287,N_10319);
or U10491 (N_10491,N_10336,N_10240);
or U10492 (N_10492,N_10296,N_10325);
nand U10493 (N_10493,N_10253,N_10298);
or U10494 (N_10494,N_10227,N_10272);
xnor U10495 (N_10495,N_10245,N_10304);
nand U10496 (N_10496,N_10225,N_10228);
and U10497 (N_10497,N_10274,N_10334);
or U10498 (N_10498,N_10348,N_10315);
nand U10499 (N_10499,N_10221,N_10207);
xnor U10500 (N_10500,N_10466,N_10425);
nor U10501 (N_10501,N_10386,N_10376);
nor U10502 (N_10502,N_10491,N_10465);
and U10503 (N_10503,N_10428,N_10445);
or U10504 (N_10504,N_10498,N_10449);
xor U10505 (N_10505,N_10394,N_10493);
nor U10506 (N_10506,N_10401,N_10487);
or U10507 (N_10507,N_10448,N_10494);
nand U10508 (N_10508,N_10410,N_10483);
nor U10509 (N_10509,N_10464,N_10353);
nand U10510 (N_10510,N_10456,N_10354);
nand U10511 (N_10511,N_10356,N_10367);
nand U10512 (N_10512,N_10358,N_10414);
nand U10513 (N_10513,N_10436,N_10399);
and U10514 (N_10514,N_10489,N_10446);
nor U10515 (N_10515,N_10463,N_10452);
nand U10516 (N_10516,N_10404,N_10460);
nor U10517 (N_10517,N_10373,N_10434);
nand U10518 (N_10518,N_10432,N_10429);
nor U10519 (N_10519,N_10473,N_10488);
xnor U10520 (N_10520,N_10443,N_10486);
xnor U10521 (N_10521,N_10388,N_10475);
and U10522 (N_10522,N_10417,N_10362);
nand U10523 (N_10523,N_10453,N_10467);
or U10524 (N_10524,N_10470,N_10459);
nand U10525 (N_10525,N_10461,N_10372);
or U10526 (N_10526,N_10442,N_10457);
nand U10527 (N_10527,N_10409,N_10398);
or U10528 (N_10528,N_10364,N_10368);
nor U10529 (N_10529,N_10416,N_10468);
or U10530 (N_10530,N_10403,N_10413);
nor U10531 (N_10531,N_10369,N_10482);
and U10532 (N_10532,N_10351,N_10384);
nand U10533 (N_10533,N_10391,N_10390);
nand U10534 (N_10534,N_10471,N_10397);
nand U10535 (N_10535,N_10438,N_10492);
nor U10536 (N_10536,N_10484,N_10497);
or U10537 (N_10537,N_10366,N_10421);
xor U10538 (N_10538,N_10355,N_10393);
and U10539 (N_10539,N_10437,N_10379);
nand U10540 (N_10540,N_10469,N_10444);
and U10541 (N_10541,N_10387,N_10407);
and U10542 (N_10542,N_10481,N_10365);
or U10543 (N_10543,N_10412,N_10480);
or U10544 (N_10544,N_10495,N_10378);
and U10545 (N_10545,N_10499,N_10462);
or U10546 (N_10546,N_10485,N_10440);
or U10547 (N_10547,N_10352,N_10479);
xor U10548 (N_10548,N_10360,N_10383);
xor U10549 (N_10549,N_10439,N_10380);
xor U10550 (N_10550,N_10431,N_10451);
xnor U10551 (N_10551,N_10455,N_10441);
nor U10552 (N_10552,N_10447,N_10405);
and U10553 (N_10553,N_10423,N_10426);
and U10554 (N_10554,N_10363,N_10418);
nor U10555 (N_10555,N_10433,N_10385);
nor U10556 (N_10556,N_10430,N_10458);
and U10557 (N_10557,N_10415,N_10357);
and U10558 (N_10558,N_10422,N_10472);
or U10559 (N_10559,N_10377,N_10424);
and U10560 (N_10560,N_10477,N_10490);
xnor U10561 (N_10561,N_10474,N_10406);
nor U10562 (N_10562,N_10450,N_10496);
nor U10563 (N_10563,N_10381,N_10408);
xor U10564 (N_10564,N_10359,N_10350);
or U10565 (N_10565,N_10396,N_10382);
nor U10566 (N_10566,N_10395,N_10420);
or U10567 (N_10567,N_10375,N_10419);
nor U10568 (N_10568,N_10402,N_10370);
nor U10569 (N_10569,N_10371,N_10389);
xnor U10570 (N_10570,N_10361,N_10411);
xor U10571 (N_10571,N_10374,N_10478);
xnor U10572 (N_10572,N_10476,N_10427);
and U10573 (N_10573,N_10454,N_10392);
nor U10574 (N_10574,N_10400,N_10435);
or U10575 (N_10575,N_10372,N_10361);
nor U10576 (N_10576,N_10386,N_10429);
and U10577 (N_10577,N_10427,N_10373);
nor U10578 (N_10578,N_10430,N_10462);
or U10579 (N_10579,N_10387,N_10375);
and U10580 (N_10580,N_10490,N_10473);
and U10581 (N_10581,N_10499,N_10354);
and U10582 (N_10582,N_10426,N_10371);
nor U10583 (N_10583,N_10437,N_10471);
nand U10584 (N_10584,N_10374,N_10444);
and U10585 (N_10585,N_10432,N_10403);
nor U10586 (N_10586,N_10471,N_10492);
or U10587 (N_10587,N_10455,N_10487);
nor U10588 (N_10588,N_10385,N_10442);
and U10589 (N_10589,N_10437,N_10354);
and U10590 (N_10590,N_10358,N_10428);
xnor U10591 (N_10591,N_10379,N_10459);
or U10592 (N_10592,N_10482,N_10375);
nand U10593 (N_10593,N_10443,N_10485);
or U10594 (N_10594,N_10392,N_10367);
and U10595 (N_10595,N_10429,N_10379);
or U10596 (N_10596,N_10364,N_10452);
and U10597 (N_10597,N_10406,N_10450);
nand U10598 (N_10598,N_10399,N_10357);
nor U10599 (N_10599,N_10428,N_10360);
xor U10600 (N_10600,N_10371,N_10465);
xnor U10601 (N_10601,N_10450,N_10360);
xor U10602 (N_10602,N_10426,N_10365);
or U10603 (N_10603,N_10487,N_10426);
and U10604 (N_10604,N_10460,N_10388);
xnor U10605 (N_10605,N_10380,N_10351);
and U10606 (N_10606,N_10362,N_10413);
nand U10607 (N_10607,N_10442,N_10484);
xor U10608 (N_10608,N_10450,N_10433);
xor U10609 (N_10609,N_10354,N_10388);
nand U10610 (N_10610,N_10467,N_10455);
xnor U10611 (N_10611,N_10406,N_10384);
or U10612 (N_10612,N_10408,N_10470);
nor U10613 (N_10613,N_10403,N_10427);
xnor U10614 (N_10614,N_10451,N_10418);
xnor U10615 (N_10615,N_10487,N_10491);
nor U10616 (N_10616,N_10457,N_10386);
nand U10617 (N_10617,N_10464,N_10428);
xnor U10618 (N_10618,N_10438,N_10382);
nand U10619 (N_10619,N_10476,N_10492);
or U10620 (N_10620,N_10486,N_10469);
and U10621 (N_10621,N_10413,N_10465);
nand U10622 (N_10622,N_10482,N_10404);
nand U10623 (N_10623,N_10435,N_10388);
nor U10624 (N_10624,N_10410,N_10436);
nor U10625 (N_10625,N_10458,N_10489);
nor U10626 (N_10626,N_10369,N_10409);
and U10627 (N_10627,N_10489,N_10475);
nor U10628 (N_10628,N_10435,N_10458);
nand U10629 (N_10629,N_10487,N_10449);
and U10630 (N_10630,N_10377,N_10437);
nand U10631 (N_10631,N_10495,N_10487);
xor U10632 (N_10632,N_10396,N_10381);
and U10633 (N_10633,N_10350,N_10455);
nor U10634 (N_10634,N_10401,N_10483);
nand U10635 (N_10635,N_10428,N_10438);
or U10636 (N_10636,N_10471,N_10353);
nand U10637 (N_10637,N_10398,N_10473);
or U10638 (N_10638,N_10404,N_10376);
xnor U10639 (N_10639,N_10395,N_10390);
nor U10640 (N_10640,N_10450,N_10446);
and U10641 (N_10641,N_10407,N_10450);
and U10642 (N_10642,N_10396,N_10439);
and U10643 (N_10643,N_10364,N_10375);
or U10644 (N_10644,N_10423,N_10467);
nand U10645 (N_10645,N_10439,N_10417);
nor U10646 (N_10646,N_10422,N_10391);
nor U10647 (N_10647,N_10411,N_10403);
xnor U10648 (N_10648,N_10443,N_10389);
or U10649 (N_10649,N_10457,N_10479);
and U10650 (N_10650,N_10535,N_10548);
nor U10651 (N_10651,N_10576,N_10618);
nor U10652 (N_10652,N_10540,N_10620);
nand U10653 (N_10653,N_10533,N_10531);
or U10654 (N_10654,N_10517,N_10514);
xor U10655 (N_10655,N_10532,N_10636);
nand U10656 (N_10656,N_10648,N_10600);
nor U10657 (N_10657,N_10643,N_10556);
or U10658 (N_10658,N_10512,N_10505);
xnor U10659 (N_10659,N_10578,N_10637);
or U10660 (N_10660,N_10501,N_10506);
or U10661 (N_10661,N_10502,N_10622);
nand U10662 (N_10662,N_10536,N_10565);
or U10663 (N_10663,N_10584,N_10573);
nand U10664 (N_10664,N_10617,N_10635);
nor U10665 (N_10665,N_10523,N_10534);
and U10666 (N_10666,N_10549,N_10644);
nand U10667 (N_10667,N_10545,N_10564);
or U10668 (N_10668,N_10553,N_10575);
nand U10669 (N_10669,N_10642,N_10627);
xor U10670 (N_10670,N_10509,N_10537);
nor U10671 (N_10671,N_10515,N_10518);
xor U10672 (N_10672,N_10590,N_10595);
nor U10673 (N_10673,N_10582,N_10615);
and U10674 (N_10674,N_10599,N_10641);
nor U10675 (N_10675,N_10607,N_10592);
nor U10676 (N_10676,N_10561,N_10546);
xor U10677 (N_10677,N_10593,N_10588);
xor U10678 (N_10678,N_10569,N_10554);
and U10679 (N_10679,N_10527,N_10602);
nand U10680 (N_10680,N_10649,N_10528);
or U10681 (N_10681,N_10568,N_10550);
or U10682 (N_10682,N_10596,N_10605);
nand U10683 (N_10683,N_10566,N_10585);
nor U10684 (N_10684,N_10581,N_10598);
nand U10685 (N_10685,N_10604,N_10521);
nand U10686 (N_10686,N_10583,N_10603);
or U10687 (N_10687,N_10629,N_10621);
or U10688 (N_10688,N_10589,N_10520);
nand U10689 (N_10689,N_10544,N_10591);
or U10690 (N_10690,N_10614,N_10547);
xor U10691 (N_10691,N_10555,N_10628);
nand U10692 (N_10692,N_10608,N_10511);
and U10693 (N_10693,N_10508,N_10526);
nand U10694 (N_10694,N_10580,N_10606);
nand U10695 (N_10695,N_10507,N_10571);
nor U10696 (N_10696,N_10625,N_10638);
nor U10697 (N_10697,N_10557,N_10616);
and U10698 (N_10698,N_10624,N_10619);
xor U10699 (N_10699,N_10567,N_10542);
and U10700 (N_10700,N_10586,N_10519);
nor U10701 (N_10701,N_10530,N_10552);
and U10702 (N_10702,N_10633,N_10634);
xnor U10703 (N_10703,N_10631,N_10645);
nor U10704 (N_10704,N_10559,N_10611);
and U10705 (N_10705,N_10504,N_10612);
nor U10706 (N_10706,N_10539,N_10543);
xor U10707 (N_10707,N_10597,N_10587);
nand U10708 (N_10708,N_10594,N_10574);
nor U10709 (N_10709,N_10601,N_10500);
xor U10710 (N_10710,N_10639,N_10647);
or U10711 (N_10711,N_10613,N_10640);
nor U10712 (N_10712,N_10538,N_10632);
nand U10713 (N_10713,N_10572,N_10503);
nand U10714 (N_10714,N_10610,N_10541);
nor U10715 (N_10715,N_10525,N_10551);
and U10716 (N_10716,N_10516,N_10623);
nor U10717 (N_10717,N_10560,N_10630);
nor U10718 (N_10718,N_10646,N_10626);
xor U10719 (N_10719,N_10529,N_10609);
or U10720 (N_10720,N_10579,N_10522);
and U10721 (N_10721,N_10558,N_10570);
nor U10722 (N_10722,N_10513,N_10524);
nor U10723 (N_10723,N_10577,N_10510);
and U10724 (N_10724,N_10563,N_10562);
or U10725 (N_10725,N_10504,N_10607);
nor U10726 (N_10726,N_10570,N_10612);
and U10727 (N_10727,N_10596,N_10553);
xor U10728 (N_10728,N_10528,N_10633);
nand U10729 (N_10729,N_10636,N_10632);
and U10730 (N_10730,N_10562,N_10516);
or U10731 (N_10731,N_10506,N_10553);
nor U10732 (N_10732,N_10509,N_10541);
nor U10733 (N_10733,N_10596,N_10649);
xor U10734 (N_10734,N_10514,N_10545);
or U10735 (N_10735,N_10580,N_10564);
and U10736 (N_10736,N_10580,N_10527);
and U10737 (N_10737,N_10632,N_10631);
or U10738 (N_10738,N_10522,N_10543);
nand U10739 (N_10739,N_10598,N_10502);
nor U10740 (N_10740,N_10577,N_10500);
or U10741 (N_10741,N_10538,N_10621);
nand U10742 (N_10742,N_10524,N_10642);
and U10743 (N_10743,N_10531,N_10567);
or U10744 (N_10744,N_10549,N_10600);
and U10745 (N_10745,N_10501,N_10502);
xnor U10746 (N_10746,N_10613,N_10597);
nor U10747 (N_10747,N_10507,N_10560);
or U10748 (N_10748,N_10607,N_10623);
and U10749 (N_10749,N_10592,N_10553);
nor U10750 (N_10750,N_10636,N_10552);
nand U10751 (N_10751,N_10562,N_10613);
nor U10752 (N_10752,N_10632,N_10647);
nand U10753 (N_10753,N_10607,N_10635);
nand U10754 (N_10754,N_10648,N_10520);
nand U10755 (N_10755,N_10513,N_10543);
nand U10756 (N_10756,N_10536,N_10600);
and U10757 (N_10757,N_10516,N_10600);
nor U10758 (N_10758,N_10584,N_10570);
and U10759 (N_10759,N_10529,N_10647);
nand U10760 (N_10760,N_10521,N_10585);
or U10761 (N_10761,N_10600,N_10628);
or U10762 (N_10762,N_10539,N_10515);
or U10763 (N_10763,N_10598,N_10636);
nand U10764 (N_10764,N_10635,N_10586);
or U10765 (N_10765,N_10619,N_10617);
and U10766 (N_10766,N_10629,N_10631);
and U10767 (N_10767,N_10503,N_10635);
xor U10768 (N_10768,N_10585,N_10522);
and U10769 (N_10769,N_10590,N_10504);
xor U10770 (N_10770,N_10584,N_10586);
nor U10771 (N_10771,N_10552,N_10610);
and U10772 (N_10772,N_10566,N_10602);
xnor U10773 (N_10773,N_10623,N_10619);
xnor U10774 (N_10774,N_10547,N_10519);
or U10775 (N_10775,N_10537,N_10617);
nand U10776 (N_10776,N_10510,N_10505);
nand U10777 (N_10777,N_10547,N_10596);
and U10778 (N_10778,N_10637,N_10617);
or U10779 (N_10779,N_10633,N_10502);
xnor U10780 (N_10780,N_10644,N_10570);
and U10781 (N_10781,N_10619,N_10577);
and U10782 (N_10782,N_10573,N_10644);
nand U10783 (N_10783,N_10509,N_10566);
or U10784 (N_10784,N_10607,N_10598);
xor U10785 (N_10785,N_10574,N_10592);
xor U10786 (N_10786,N_10589,N_10517);
nor U10787 (N_10787,N_10623,N_10590);
or U10788 (N_10788,N_10511,N_10538);
and U10789 (N_10789,N_10615,N_10601);
nor U10790 (N_10790,N_10560,N_10543);
and U10791 (N_10791,N_10513,N_10576);
and U10792 (N_10792,N_10540,N_10642);
and U10793 (N_10793,N_10523,N_10610);
nor U10794 (N_10794,N_10585,N_10545);
nand U10795 (N_10795,N_10535,N_10638);
nand U10796 (N_10796,N_10555,N_10539);
or U10797 (N_10797,N_10530,N_10546);
or U10798 (N_10798,N_10532,N_10619);
nand U10799 (N_10799,N_10527,N_10542);
and U10800 (N_10800,N_10746,N_10785);
xnor U10801 (N_10801,N_10702,N_10776);
xor U10802 (N_10802,N_10666,N_10754);
xor U10803 (N_10803,N_10768,N_10718);
or U10804 (N_10804,N_10739,N_10792);
nand U10805 (N_10805,N_10701,N_10758);
nor U10806 (N_10806,N_10752,N_10766);
nand U10807 (N_10807,N_10659,N_10738);
xnor U10808 (N_10808,N_10760,N_10654);
and U10809 (N_10809,N_10729,N_10767);
and U10810 (N_10810,N_10687,N_10715);
nor U10811 (N_10811,N_10799,N_10781);
nand U10812 (N_10812,N_10740,N_10726);
and U10813 (N_10813,N_10679,N_10663);
and U10814 (N_10814,N_10782,N_10783);
nor U10815 (N_10815,N_10689,N_10751);
nor U10816 (N_10816,N_10677,N_10753);
or U10817 (N_10817,N_10672,N_10728);
xor U10818 (N_10818,N_10712,N_10691);
or U10819 (N_10819,N_10736,N_10731);
and U10820 (N_10820,N_10693,N_10684);
or U10821 (N_10821,N_10720,N_10668);
or U10822 (N_10822,N_10749,N_10723);
and U10823 (N_10823,N_10786,N_10690);
xnor U10824 (N_10824,N_10730,N_10655);
and U10825 (N_10825,N_10657,N_10791);
nor U10826 (N_10826,N_10775,N_10704);
xnor U10827 (N_10827,N_10700,N_10713);
or U10828 (N_10828,N_10793,N_10745);
or U10829 (N_10829,N_10709,N_10722);
xnor U10830 (N_10830,N_10790,N_10737);
xor U10831 (N_10831,N_10763,N_10770);
or U10832 (N_10832,N_10761,N_10673);
and U10833 (N_10833,N_10708,N_10756);
or U10834 (N_10834,N_10676,N_10777);
xor U10835 (N_10835,N_10686,N_10795);
xnor U10836 (N_10836,N_10757,N_10675);
and U10837 (N_10837,N_10710,N_10674);
nor U10838 (N_10838,N_10762,N_10721);
or U10839 (N_10839,N_10716,N_10727);
nand U10840 (N_10840,N_10688,N_10788);
xor U10841 (N_10841,N_10773,N_10741);
xnor U10842 (N_10842,N_10661,N_10759);
xor U10843 (N_10843,N_10765,N_10744);
nor U10844 (N_10844,N_10707,N_10733);
or U10845 (N_10845,N_10724,N_10662);
and U10846 (N_10846,N_10692,N_10695);
or U10847 (N_10847,N_10735,N_10683);
nand U10848 (N_10848,N_10653,N_10769);
and U10849 (N_10849,N_10685,N_10774);
nor U10850 (N_10850,N_10650,N_10711);
nand U10851 (N_10851,N_10678,N_10669);
nand U10852 (N_10852,N_10725,N_10772);
nor U10853 (N_10853,N_10658,N_10699);
nand U10854 (N_10854,N_10656,N_10747);
and U10855 (N_10855,N_10664,N_10755);
nand U10856 (N_10856,N_10706,N_10714);
and U10857 (N_10857,N_10784,N_10796);
nor U10858 (N_10858,N_10734,N_10698);
nor U10859 (N_10859,N_10652,N_10671);
xor U10860 (N_10860,N_10798,N_10680);
nand U10861 (N_10861,N_10748,N_10771);
xnor U10862 (N_10862,N_10743,N_10750);
and U10863 (N_10863,N_10681,N_10670);
xor U10864 (N_10864,N_10667,N_10665);
nand U10865 (N_10865,N_10778,N_10764);
nand U10866 (N_10866,N_10717,N_10787);
xnor U10867 (N_10867,N_10660,N_10780);
nand U10868 (N_10868,N_10696,N_10697);
and U10869 (N_10869,N_10789,N_10694);
and U10870 (N_10870,N_10794,N_10719);
nand U10871 (N_10871,N_10797,N_10682);
nor U10872 (N_10872,N_10651,N_10705);
xor U10873 (N_10873,N_10732,N_10703);
nand U10874 (N_10874,N_10779,N_10742);
xor U10875 (N_10875,N_10794,N_10724);
and U10876 (N_10876,N_10742,N_10678);
nand U10877 (N_10877,N_10786,N_10799);
nor U10878 (N_10878,N_10690,N_10735);
xnor U10879 (N_10879,N_10732,N_10679);
and U10880 (N_10880,N_10778,N_10697);
xnor U10881 (N_10881,N_10681,N_10776);
xnor U10882 (N_10882,N_10730,N_10661);
xor U10883 (N_10883,N_10654,N_10715);
nand U10884 (N_10884,N_10711,N_10678);
nand U10885 (N_10885,N_10694,N_10711);
and U10886 (N_10886,N_10748,N_10730);
nor U10887 (N_10887,N_10671,N_10762);
or U10888 (N_10888,N_10653,N_10701);
xor U10889 (N_10889,N_10779,N_10748);
nor U10890 (N_10890,N_10731,N_10777);
and U10891 (N_10891,N_10672,N_10753);
nand U10892 (N_10892,N_10743,N_10775);
nand U10893 (N_10893,N_10776,N_10704);
nand U10894 (N_10894,N_10659,N_10790);
xor U10895 (N_10895,N_10779,N_10766);
or U10896 (N_10896,N_10698,N_10672);
nor U10897 (N_10897,N_10758,N_10703);
or U10898 (N_10898,N_10666,N_10778);
nand U10899 (N_10899,N_10692,N_10756);
and U10900 (N_10900,N_10691,N_10736);
xor U10901 (N_10901,N_10651,N_10688);
or U10902 (N_10902,N_10790,N_10700);
nor U10903 (N_10903,N_10761,N_10681);
or U10904 (N_10904,N_10670,N_10679);
nand U10905 (N_10905,N_10733,N_10737);
or U10906 (N_10906,N_10707,N_10748);
or U10907 (N_10907,N_10777,N_10670);
nand U10908 (N_10908,N_10669,N_10694);
or U10909 (N_10909,N_10724,N_10739);
nor U10910 (N_10910,N_10680,N_10711);
xor U10911 (N_10911,N_10746,N_10745);
nor U10912 (N_10912,N_10740,N_10776);
xor U10913 (N_10913,N_10784,N_10651);
or U10914 (N_10914,N_10675,N_10716);
nand U10915 (N_10915,N_10664,N_10795);
nor U10916 (N_10916,N_10773,N_10753);
or U10917 (N_10917,N_10758,N_10723);
nor U10918 (N_10918,N_10722,N_10784);
xnor U10919 (N_10919,N_10742,N_10754);
nor U10920 (N_10920,N_10689,N_10752);
or U10921 (N_10921,N_10668,N_10715);
xor U10922 (N_10922,N_10715,N_10694);
xor U10923 (N_10923,N_10668,N_10769);
xor U10924 (N_10924,N_10716,N_10693);
nor U10925 (N_10925,N_10779,N_10789);
nor U10926 (N_10926,N_10699,N_10716);
xnor U10927 (N_10927,N_10689,N_10755);
and U10928 (N_10928,N_10689,N_10742);
and U10929 (N_10929,N_10742,N_10786);
nand U10930 (N_10930,N_10737,N_10756);
or U10931 (N_10931,N_10686,N_10748);
xnor U10932 (N_10932,N_10782,N_10796);
nand U10933 (N_10933,N_10792,N_10712);
or U10934 (N_10934,N_10734,N_10686);
nand U10935 (N_10935,N_10651,N_10716);
or U10936 (N_10936,N_10703,N_10726);
nor U10937 (N_10937,N_10760,N_10670);
xnor U10938 (N_10938,N_10695,N_10749);
or U10939 (N_10939,N_10702,N_10689);
or U10940 (N_10940,N_10653,N_10673);
nand U10941 (N_10941,N_10709,N_10714);
xnor U10942 (N_10942,N_10716,N_10788);
and U10943 (N_10943,N_10690,N_10653);
xor U10944 (N_10944,N_10715,N_10713);
nor U10945 (N_10945,N_10738,N_10687);
or U10946 (N_10946,N_10655,N_10732);
nor U10947 (N_10947,N_10670,N_10738);
or U10948 (N_10948,N_10658,N_10755);
nand U10949 (N_10949,N_10683,N_10744);
or U10950 (N_10950,N_10910,N_10870);
nand U10951 (N_10951,N_10802,N_10871);
nand U10952 (N_10952,N_10810,N_10878);
nor U10953 (N_10953,N_10808,N_10845);
and U10954 (N_10954,N_10809,N_10858);
nor U10955 (N_10955,N_10939,N_10853);
and U10956 (N_10956,N_10839,N_10846);
or U10957 (N_10957,N_10921,N_10840);
nand U10958 (N_10958,N_10805,N_10823);
or U10959 (N_10959,N_10857,N_10913);
nor U10960 (N_10960,N_10822,N_10905);
and U10961 (N_10961,N_10900,N_10886);
xnor U10962 (N_10962,N_10936,N_10942);
nand U10963 (N_10963,N_10836,N_10838);
xnor U10964 (N_10964,N_10875,N_10918);
nand U10965 (N_10965,N_10803,N_10800);
xor U10966 (N_10966,N_10830,N_10880);
and U10967 (N_10967,N_10863,N_10920);
nor U10968 (N_10968,N_10818,N_10841);
and U10969 (N_10969,N_10855,N_10887);
and U10970 (N_10970,N_10860,N_10842);
xor U10971 (N_10971,N_10949,N_10877);
or U10972 (N_10972,N_10931,N_10907);
and U10973 (N_10973,N_10849,N_10806);
nor U10974 (N_10974,N_10843,N_10854);
nand U10975 (N_10975,N_10941,N_10844);
xor U10976 (N_10976,N_10945,N_10820);
nor U10977 (N_10977,N_10885,N_10821);
or U10978 (N_10978,N_10825,N_10874);
or U10979 (N_10979,N_10917,N_10948);
nor U10980 (N_10980,N_10850,N_10816);
nor U10981 (N_10981,N_10893,N_10894);
or U10982 (N_10982,N_10867,N_10851);
or U10983 (N_10983,N_10902,N_10940);
nor U10984 (N_10984,N_10925,N_10888);
nor U10985 (N_10985,N_10909,N_10944);
xnor U10986 (N_10986,N_10938,N_10801);
xor U10987 (N_10987,N_10916,N_10834);
and U10988 (N_10988,N_10911,N_10924);
nand U10989 (N_10989,N_10828,N_10804);
xnor U10990 (N_10990,N_10869,N_10829);
nand U10991 (N_10991,N_10831,N_10837);
and U10992 (N_10992,N_10872,N_10919);
nor U10993 (N_10993,N_10932,N_10832);
or U10994 (N_10994,N_10897,N_10935);
and U10995 (N_10995,N_10906,N_10896);
nor U10996 (N_10996,N_10826,N_10811);
nand U10997 (N_10997,N_10827,N_10813);
xor U10998 (N_10998,N_10817,N_10879);
nand U10999 (N_10999,N_10912,N_10883);
nor U11000 (N_11000,N_10864,N_10891);
or U11001 (N_11001,N_10856,N_10812);
and U11002 (N_11002,N_10852,N_10928);
nor U11003 (N_11003,N_10868,N_10895);
nand U11004 (N_11004,N_10847,N_10833);
or U11005 (N_11005,N_10933,N_10892);
and U11006 (N_11006,N_10943,N_10889);
nor U11007 (N_11007,N_10915,N_10884);
nand U11008 (N_11008,N_10937,N_10901);
nor U11009 (N_11009,N_10861,N_10929);
or U11010 (N_11010,N_10815,N_10904);
xnor U11011 (N_11011,N_10862,N_10882);
xnor U11012 (N_11012,N_10898,N_10814);
nor U11013 (N_11013,N_10881,N_10947);
nor U11014 (N_11014,N_10934,N_10922);
nor U11015 (N_11015,N_10926,N_10866);
nor U11016 (N_11016,N_10930,N_10873);
xor U11017 (N_11017,N_10819,N_10807);
and U11018 (N_11018,N_10927,N_10890);
nand U11019 (N_11019,N_10835,N_10899);
and U11020 (N_11020,N_10848,N_10914);
xnor U11021 (N_11021,N_10824,N_10876);
nand U11022 (N_11022,N_10923,N_10946);
nand U11023 (N_11023,N_10908,N_10903);
nand U11024 (N_11024,N_10859,N_10865);
and U11025 (N_11025,N_10813,N_10825);
xnor U11026 (N_11026,N_10934,N_10895);
xnor U11027 (N_11027,N_10804,N_10905);
or U11028 (N_11028,N_10847,N_10817);
and U11029 (N_11029,N_10870,N_10808);
nor U11030 (N_11030,N_10864,N_10867);
nor U11031 (N_11031,N_10859,N_10947);
and U11032 (N_11032,N_10817,N_10832);
xor U11033 (N_11033,N_10889,N_10922);
nand U11034 (N_11034,N_10932,N_10935);
nand U11035 (N_11035,N_10929,N_10915);
nor U11036 (N_11036,N_10847,N_10826);
nand U11037 (N_11037,N_10816,N_10819);
and U11038 (N_11038,N_10830,N_10814);
nand U11039 (N_11039,N_10930,N_10921);
and U11040 (N_11040,N_10887,N_10916);
nor U11041 (N_11041,N_10930,N_10820);
and U11042 (N_11042,N_10903,N_10912);
nor U11043 (N_11043,N_10919,N_10805);
or U11044 (N_11044,N_10846,N_10927);
or U11045 (N_11045,N_10910,N_10865);
or U11046 (N_11046,N_10811,N_10905);
or U11047 (N_11047,N_10833,N_10800);
xor U11048 (N_11048,N_10843,N_10823);
nor U11049 (N_11049,N_10823,N_10825);
nand U11050 (N_11050,N_10907,N_10867);
nand U11051 (N_11051,N_10861,N_10871);
or U11052 (N_11052,N_10856,N_10923);
xor U11053 (N_11053,N_10830,N_10852);
nor U11054 (N_11054,N_10829,N_10817);
nand U11055 (N_11055,N_10800,N_10859);
and U11056 (N_11056,N_10879,N_10835);
xnor U11057 (N_11057,N_10834,N_10854);
xor U11058 (N_11058,N_10893,N_10824);
nor U11059 (N_11059,N_10930,N_10923);
nor U11060 (N_11060,N_10810,N_10889);
nand U11061 (N_11061,N_10826,N_10883);
and U11062 (N_11062,N_10919,N_10839);
xor U11063 (N_11063,N_10833,N_10935);
or U11064 (N_11064,N_10811,N_10920);
and U11065 (N_11065,N_10846,N_10906);
or U11066 (N_11066,N_10804,N_10833);
and U11067 (N_11067,N_10927,N_10810);
nand U11068 (N_11068,N_10837,N_10809);
nor U11069 (N_11069,N_10939,N_10849);
and U11070 (N_11070,N_10851,N_10825);
or U11071 (N_11071,N_10873,N_10870);
nor U11072 (N_11072,N_10887,N_10939);
nor U11073 (N_11073,N_10899,N_10803);
or U11074 (N_11074,N_10856,N_10857);
or U11075 (N_11075,N_10802,N_10915);
or U11076 (N_11076,N_10829,N_10947);
or U11077 (N_11077,N_10803,N_10880);
nor U11078 (N_11078,N_10815,N_10906);
nand U11079 (N_11079,N_10878,N_10902);
or U11080 (N_11080,N_10847,N_10864);
and U11081 (N_11081,N_10864,N_10802);
and U11082 (N_11082,N_10897,N_10865);
or U11083 (N_11083,N_10922,N_10810);
nor U11084 (N_11084,N_10892,N_10819);
nor U11085 (N_11085,N_10821,N_10835);
nor U11086 (N_11086,N_10893,N_10829);
nor U11087 (N_11087,N_10855,N_10943);
nor U11088 (N_11088,N_10838,N_10811);
and U11089 (N_11089,N_10867,N_10880);
nand U11090 (N_11090,N_10819,N_10844);
and U11091 (N_11091,N_10832,N_10865);
or U11092 (N_11092,N_10904,N_10913);
and U11093 (N_11093,N_10914,N_10838);
xor U11094 (N_11094,N_10942,N_10885);
xnor U11095 (N_11095,N_10879,N_10927);
nor U11096 (N_11096,N_10814,N_10839);
nor U11097 (N_11097,N_10905,N_10906);
xor U11098 (N_11098,N_10832,N_10878);
nor U11099 (N_11099,N_10907,N_10937);
xnor U11100 (N_11100,N_11051,N_11097);
or U11101 (N_11101,N_11096,N_10972);
and U11102 (N_11102,N_10977,N_10971);
and U11103 (N_11103,N_11089,N_11000);
nand U11104 (N_11104,N_11048,N_10976);
or U11105 (N_11105,N_11078,N_11030);
or U11106 (N_11106,N_11095,N_11027);
and U11107 (N_11107,N_10969,N_11090);
nor U11108 (N_11108,N_10978,N_11009);
and U11109 (N_11109,N_11006,N_10956);
nand U11110 (N_11110,N_11018,N_10961);
nor U11111 (N_11111,N_11004,N_11080);
or U11112 (N_11112,N_11024,N_11075);
and U11113 (N_11113,N_10986,N_11028);
and U11114 (N_11114,N_11012,N_11062);
or U11115 (N_11115,N_11003,N_11063);
nor U11116 (N_11116,N_10981,N_11053);
and U11117 (N_11117,N_11025,N_11046);
nor U11118 (N_11118,N_10973,N_10993);
nand U11119 (N_11119,N_11040,N_11047);
xor U11120 (N_11120,N_11098,N_11061);
and U11121 (N_11121,N_11081,N_10982);
nand U11122 (N_11122,N_10995,N_10975);
nor U11123 (N_11123,N_11015,N_11065);
nand U11124 (N_11124,N_10974,N_10985);
or U11125 (N_11125,N_10953,N_11005);
and U11126 (N_11126,N_11079,N_11092);
xnor U11127 (N_11127,N_10954,N_10980);
nand U11128 (N_11128,N_11042,N_10989);
or U11129 (N_11129,N_10983,N_11021);
nor U11130 (N_11130,N_10966,N_11074);
nand U11131 (N_11131,N_10991,N_10994);
nor U11132 (N_11132,N_11059,N_10965);
nor U11133 (N_11133,N_10964,N_11085);
xnor U11134 (N_11134,N_11084,N_11001);
xnor U11135 (N_11135,N_11029,N_11023);
and U11136 (N_11136,N_11044,N_11019);
nand U11137 (N_11137,N_11071,N_10958);
xor U11138 (N_11138,N_11050,N_10988);
or U11139 (N_11139,N_11094,N_11007);
xor U11140 (N_11140,N_11041,N_11013);
xnor U11141 (N_11141,N_11020,N_10950);
xor U11142 (N_11142,N_11087,N_11056);
and U11143 (N_11143,N_11038,N_11036);
xor U11144 (N_11144,N_11039,N_11070);
and U11145 (N_11145,N_11037,N_11086);
nand U11146 (N_11146,N_11069,N_10999);
nor U11147 (N_11147,N_10984,N_11035);
nand U11148 (N_11148,N_10992,N_10997);
nand U11149 (N_11149,N_11049,N_10962);
or U11150 (N_11150,N_10955,N_10990);
xnor U11151 (N_11151,N_11026,N_11083);
and U11152 (N_11152,N_11045,N_11067);
xnor U11153 (N_11153,N_11031,N_11076);
or U11154 (N_11154,N_11064,N_10968);
xor U11155 (N_11155,N_11082,N_11093);
nand U11156 (N_11156,N_10957,N_10951);
nor U11157 (N_11157,N_10952,N_10998);
nand U11158 (N_11158,N_11058,N_11060);
and U11159 (N_11159,N_11010,N_10970);
nand U11160 (N_11160,N_11073,N_11016);
or U11161 (N_11161,N_11043,N_11032);
xnor U11162 (N_11162,N_11077,N_10959);
or U11163 (N_11163,N_11088,N_11055);
xnor U11164 (N_11164,N_10967,N_11033);
nor U11165 (N_11165,N_11011,N_10987);
nand U11166 (N_11166,N_11057,N_11054);
nor U11167 (N_11167,N_11022,N_10996);
xnor U11168 (N_11168,N_11072,N_11014);
xor U11169 (N_11169,N_11002,N_11099);
or U11170 (N_11170,N_11052,N_10963);
or U11171 (N_11171,N_11034,N_11091);
nand U11172 (N_11172,N_10979,N_10960);
nand U11173 (N_11173,N_11066,N_11008);
or U11174 (N_11174,N_11017,N_11068);
and U11175 (N_11175,N_10965,N_11022);
and U11176 (N_11176,N_11071,N_11097);
or U11177 (N_11177,N_11054,N_10997);
or U11178 (N_11178,N_11061,N_11018);
nand U11179 (N_11179,N_10956,N_10951);
nand U11180 (N_11180,N_11021,N_11072);
or U11181 (N_11181,N_11010,N_11004);
nor U11182 (N_11182,N_10999,N_11085);
and U11183 (N_11183,N_11038,N_11089);
and U11184 (N_11184,N_10972,N_11039);
or U11185 (N_11185,N_11020,N_11011);
nand U11186 (N_11186,N_11080,N_11023);
xnor U11187 (N_11187,N_11069,N_10955);
xor U11188 (N_11188,N_11027,N_11066);
nand U11189 (N_11189,N_11004,N_10992);
xnor U11190 (N_11190,N_10972,N_11019);
nor U11191 (N_11191,N_11032,N_11093);
nand U11192 (N_11192,N_11099,N_11074);
xnor U11193 (N_11193,N_11052,N_11017);
or U11194 (N_11194,N_10953,N_11023);
or U11195 (N_11195,N_11042,N_11007);
nand U11196 (N_11196,N_11054,N_10953);
nor U11197 (N_11197,N_10994,N_11077);
xnor U11198 (N_11198,N_10951,N_10960);
and U11199 (N_11199,N_11095,N_11029);
nand U11200 (N_11200,N_11017,N_11062);
nand U11201 (N_11201,N_10979,N_11084);
nor U11202 (N_11202,N_11072,N_10998);
nand U11203 (N_11203,N_11069,N_10962);
and U11204 (N_11204,N_10965,N_11027);
or U11205 (N_11205,N_10990,N_10980);
or U11206 (N_11206,N_11036,N_10994);
or U11207 (N_11207,N_11046,N_11099);
or U11208 (N_11208,N_10972,N_11091);
xnor U11209 (N_11209,N_11011,N_10990);
xor U11210 (N_11210,N_10979,N_11099);
nor U11211 (N_11211,N_11029,N_11046);
and U11212 (N_11212,N_11076,N_11066);
nand U11213 (N_11213,N_11043,N_11072);
and U11214 (N_11214,N_11039,N_10985);
and U11215 (N_11215,N_10994,N_10957);
and U11216 (N_11216,N_11033,N_10978);
nor U11217 (N_11217,N_11090,N_11085);
xor U11218 (N_11218,N_11072,N_11018);
nor U11219 (N_11219,N_11072,N_11049);
nor U11220 (N_11220,N_11004,N_11067);
or U11221 (N_11221,N_10969,N_11093);
and U11222 (N_11222,N_11062,N_11038);
nor U11223 (N_11223,N_10990,N_10994);
nand U11224 (N_11224,N_10961,N_11022);
nand U11225 (N_11225,N_11007,N_11083);
and U11226 (N_11226,N_11023,N_10998);
nand U11227 (N_11227,N_11030,N_11072);
or U11228 (N_11228,N_11073,N_11031);
nand U11229 (N_11229,N_10982,N_11028);
nand U11230 (N_11230,N_11065,N_11017);
nor U11231 (N_11231,N_10998,N_11095);
nand U11232 (N_11232,N_11068,N_11042);
or U11233 (N_11233,N_10957,N_11080);
nor U11234 (N_11234,N_11038,N_11009);
xor U11235 (N_11235,N_11089,N_11039);
nor U11236 (N_11236,N_10964,N_10953);
xnor U11237 (N_11237,N_11078,N_11073);
xor U11238 (N_11238,N_10973,N_11081);
or U11239 (N_11239,N_10950,N_10997);
or U11240 (N_11240,N_10985,N_11056);
xnor U11241 (N_11241,N_11015,N_11035);
and U11242 (N_11242,N_10997,N_10954);
nor U11243 (N_11243,N_10979,N_10990);
and U11244 (N_11244,N_11042,N_10962);
or U11245 (N_11245,N_11085,N_11086);
nor U11246 (N_11246,N_10960,N_10992);
and U11247 (N_11247,N_11066,N_11013);
or U11248 (N_11248,N_11078,N_10998);
nand U11249 (N_11249,N_11057,N_10994);
xor U11250 (N_11250,N_11217,N_11188);
nor U11251 (N_11251,N_11231,N_11145);
nor U11252 (N_11252,N_11183,N_11201);
xor U11253 (N_11253,N_11227,N_11208);
nor U11254 (N_11254,N_11125,N_11216);
nor U11255 (N_11255,N_11211,N_11238);
nor U11256 (N_11256,N_11156,N_11179);
nand U11257 (N_11257,N_11147,N_11166);
nand U11258 (N_11258,N_11234,N_11162);
xnor U11259 (N_11259,N_11213,N_11108);
or U11260 (N_11260,N_11247,N_11109);
or U11261 (N_11261,N_11171,N_11116);
and U11262 (N_11262,N_11221,N_11244);
nor U11263 (N_11263,N_11240,N_11118);
nand U11264 (N_11264,N_11248,N_11105);
nor U11265 (N_11265,N_11161,N_11165);
and U11266 (N_11266,N_11112,N_11160);
nor U11267 (N_11267,N_11167,N_11198);
and U11268 (N_11268,N_11168,N_11215);
nor U11269 (N_11269,N_11134,N_11139);
xor U11270 (N_11270,N_11131,N_11197);
or U11271 (N_11271,N_11140,N_11218);
or U11272 (N_11272,N_11151,N_11192);
nand U11273 (N_11273,N_11203,N_11214);
nor U11274 (N_11274,N_11141,N_11136);
nor U11275 (N_11275,N_11154,N_11194);
nor U11276 (N_11276,N_11103,N_11107);
or U11277 (N_11277,N_11121,N_11178);
nand U11278 (N_11278,N_11126,N_11219);
or U11279 (N_11279,N_11132,N_11129);
nor U11280 (N_11280,N_11128,N_11235);
nor U11281 (N_11281,N_11142,N_11182);
and U11282 (N_11282,N_11209,N_11164);
nand U11283 (N_11283,N_11157,N_11241);
and U11284 (N_11284,N_11133,N_11184);
xor U11285 (N_11285,N_11224,N_11246);
or U11286 (N_11286,N_11102,N_11124);
and U11287 (N_11287,N_11143,N_11239);
and U11288 (N_11288,N_11245,N_11200);
nand U11289 (N_11289,N_11135,N_11137);
xor U11290 (N_11290,N_11196,N_11193);
xnor U11291 (N_11291,N_11220,N_11175);
nor U11292 (N_11292,N_11190,N_11228);
and U11293 (N_11293,N_11104,N_11172);
nand U11294 (N_11294,N_11176,N_11187);
nor U11295 (N_11295,N_11243,N_11101);
nand U11296 (N_11296,N_11229,N_11199);
or U11297 (N_11297,N_11242,N_11195);
nor U11298 (N_11298,N_11115,N_11123);
nor U11299 (N_11299,N_11149,N_11249);
nand U11300 (N_11300,N_11138,N_11113);
nor U11301 (N_11301,N_11127,N_11146);
or U11302 (N_11302,N_11237,N_11236);
nor U11303 (N_11303,N_11174,N_11169);
xnor U11304 (N_11304,N_11226,N_11153);
or U11305 (N_11305,N_11212,N_11148);
and U11306 (N_11306,N_11204,N_11117);
nor U11307 (N_11307,N_11119,N_11158);
nor U11308 (N_11308,N_11170,N_11191);
and U11309 (N_11309,N_11185,N_11120);
nand U11310 (N_11310,N_11223,N_11180);
nand U11311 (N_11311,N_11155,N_11222);
nor U11312 (N_11312,N_11159,N_11163);
or U11313 (N_11313,N_11150,N_11110);
nand U11314 (N_11314,N_11177,N_11230);
nand U11315 (N_11315,N_11202,N_11106);
or U11316 (N_11316,N_11111,N_11181);
and U11317 (N_11317,N_11114,N_11173);
or U11318 (N_11318,N_11186,N_11122);
nor U11319 (N_11319,N_11210,N_11189);
or U11320 (N_11320,N_11232,N_11130);
and U11321 (N_11321,N_11225,N_11206);
nand U11322 (N_11322,N_11233,N_11144);
or U11323 (N_11323,N_11100,N_11152);
or U11324 (N_11324,N_11207,N_11205);
nor U11325 (N_11325,N_11241,N_11126);
nor U11326 (N_11326,N_11107,N_11160);
and U11327 (N_11327,N_11117,N_11172);
or U11328 (N_11328,N_11212,N_11201);
nor U11329 (N_11329,N_11119,N_11173);
nand U11330 (N_11330,N_11235,N_11175);
nand U11331 (N_11331,N_11155,N_11110);
xnor U11332 (N_11332,N_11130,N_11248);
or U11333 (N_11333,N_11116,N_11243);
nand U11334 (N_11334,N_11110,N_11236);
xor U11335 (N_11335,N_11197,N_11146);
nor U11336 (N_11336,N_11191,N_11231);
nor U11337 (N_11337,N_11229,N_11149);
and U11338 (N_11338,N_11190,N_11137);
nand U11339 (N_11339,N_11208,N_11149);
nor U11340 (N_11340,N_11177,N_11108);
or U11341 (N_11341,N_11205,N_11105);
nand U11342 (N_11342,N_11183,N_11206);
nor U11343 (N_11343,N_11186,N_11237);
and U11344 (N_11344,N_11212,N_11174);
and U11345 (N_11345,N_11169,N_11155);
and U11346 (N_11346,N_11114,N_11171);
nand U11347 (N_11347,N_11122,N_11120);
nand U11348 (N_11348,N_11177,N_11225);
nor U11349 (N_11349,N_11249,N_11218);
or U11350 (N_11350,N_11150,N_11186);
and U11351 (N_11351,N_11239,N_11106);
or U11352 (N_11352,N_11180,N_11167);
or U11353 (N_11353,N_11140,N_11136);
nand U11354 (N_11354,N_11101,N_11128);
xor U11355 (N_11355,N_11244,N_11205);
nor U11356 (N_11356,N_11167,N_11203);
or U11357 (N_11357,N_11167,N_11210);
nand U11358 (N_11358,N_11125,N_11213);
or U11359 (N_11359,N_11167,N_11128);
and U11360 (N_11360,N_11167,N_11124);
and U11361 (N_11361,N_11191,N_11212);
xor U11362 (N_11362,N_11102,N_11235);
nand U11363 (N_11363,N_11228,N_11175);
nand U11364 (N_11364,N_11117,N_11176);
nor U11365 (N_11365,N_11175,N_11183);
nand U11366 (N_11366,N_11153,N_11128);
nor U11367 (N_11367,N_11125,N_11178);
and U11368 (N_11368,N_11194,N_11135);
and U11369 (N_11369,N_11116,N_11209);
nor U11370 (N_11370,N_11182,N_11184);
and U11371 (N_11371,N_11197,N_11175);
and U11372 (N_11372,N_11121,N_11157);
or U11373 (N_11373,N_11246,N_11167);
nor U11374 (N_11374,N_11234,N_11220);
xnor U11375 (N_11375,N_11174,N_11197);
and U11376 (N_11376,N_11196,N_11179);
nor U11377 (N_11377,N_11149,N_11185);
and U11378 (N_11378,N_11128,N_11186);
nor U11379 (N_11379,N_11205,N_11170);
and U11380 (N_11380,N_11111,N_11150);
or U11381 (N_11381,N_11219,N_11152);
nor U11382 (N_11382,N_11117,N_11244);
and U11383 (N_11383,N_11193,N_11131);
xnor U11384 (N_11384,N_11220,N_11237);
nor U11385 (N_11385,N_11126,N_11163);
or U11386 (N_11386,N_11114,N_11184);
or U11387 (N_11387,N_11249,N_11169);
nand U11388 (N_11388,N_11168,N_11106);
or U11389 (N_11389,N_11121,N_11237);
nor U11390 (N_11390,N_11172,N_11171);
xor U11391 (N_11391,N_11104,N_11158);
xnor U11392 (N_11392,N_11246,N_11136);
nor U11393 (N_11393,N_11236,N_11114);
or U11394 (N_11394,N_11157,N_11230);
nand U11395 (N_11395,N_11191,N_11141);
or U11396 (N_11396,N_11229,N_11179);
xor U11397 (N_11397,N_11123,N_11160);
nor U11398 (N_11398,N_11114,N_11124);
and U11399 (N_11399,N_11141,N_11164);
nor U11400 (N_11400,N_11265,N_11380);
xor U11401 (N_11401,N_11261,N_11363);
and U11402 (N_11402,N_11358,N_11291);
nand U11403 (N_11403,N_11276,N_11321);
or U11404 (N_11404,N_11369,N_11256);
nand U11405 (N_11405,N_11304,N_11356);
xor U11406 (N_11406,N_11326,N_11340);
and U11407 (N_11407,N_11327,N_11374);
xnor U11408 (N_11408,N_11364,N_11310);
nand U11409 (N_11409,N_11362,N_11320);
nand U11410 (N_11410,N_11395,N_11251);
nand U11411 (N_11411,N_11300,N_11324);
or U11412 (N_11412,N_11336,N_11378);
or U11413 (N_11413,N_11318,N_11302);
and U11414 (N_11414,N_11385,N_11286);
and U11415 (N_11415,N_11383,N_11387);
and U11416 (N_11416,N_11330,N_11294);
xor U11417 (N_11417,N_11386,N_11303);
or U11418 (N_11418,N_11375,N_11257);
and U11419 (N_11419,N_11266,N_11331);
nand U11420 (N_11420,N_11269,N_11317);
nand U11421 (N_11421,N_11264,N_11262);
xor U11422 (N_11422,N_11323,N_11377);
or U11423 (N_11423,N_11360,N_11339);
or U11424 (N_11424,N_11347,N_11287);
and U11425 (N_11425,N_11329,N_11392);
or U11426 (N_11426,N_11384,N_11338);
nor U11427 (N_11427,N_11273,N_11292);
or U11428 (N_11428,N_11350,N_11315);
nor U11429 (N_11429,N_11376,N_11333);
and U11430 (N_11430,N_11370,N_11361);
and U11431 (N_11431,N_11313,N_11296);
or U11432 (N_11432,N_11278,N_11354);
nor U11433 (N_11433,N_11275,N_11373);
xor U11434 (N_11434,N_11306,N_11282);
and U11435 (N_11435,N_11263,N_11393);
or U11436 (N_11436,N_11274,N_11283);
and U11437 (N_11437,N_11258,N_11343);
and U11438 (N_11438,N_11399,N_11382);
or U11439 (N_11439,N_11389,N_11341);
nor U11440 (N_11440,N_11355,N_11367);
xor U11441 (N_11441,N_11365,N_11368);
nor U11442 (N_11442,N_11268,N_11379);
xor U11443 (N_11443,N_11381,N_11398);
and U11444 (N_11444,N_11332,N_11281);
nand U11445 (N_11445,N_11345,N_11295);
or U11446 (N_11446,N_11335,N_11305);
nand U11447 (N_11447,N_11325,N_11372);
and U11448 (N_11448,N_11301,N_11388);
nand U11449 (N_11449,N_11348,N_11316);
or U11450 (N_11450,N_11284,N_11353);
and U11451 (N_11451,N_11308,N_11298);
or U11452 (N_11452,N_11307,N_11297);
xor U11453 (N_11453,N_11259,N_11346);
nand U11454 (N_11454,N_11357,N_11272);
nand U11455 (N_11455,N_11250,N_11311);
and U11456 (N_11456,N_11277,N_11390);
nand U11457 (N_11457,N_11351,N_11289);
nand U11458 (N_11458,N_11397,N_11342);
or U11459 (N_11459,N_11260,N_11253);
nand U11460 (N_11460,N_11352,N_11293);
nor U11461 (N_11461,N_11328,N_11309);
or U11462 (N_11462,N_11394,N_11270);
or U11463 (N_11463,N_11255,N_11337);
and U11464 (N_11464,N_11254,N_11252);
nor U11465 (N_11465,N_11279,N_11312);
xor U11466 (N_11466,N_11359,N_11271);
or U11467 (N_11467,N_11285,N_11267);
nand U11468 (N_11468,N_11322,N_11334);
nand U11469 (N_11469,N_11314,N_11349);
xor U11470 (N_11470,N_11299,N_11396);
nor U11471 (N_11471,N_11391,N_11344);
nor U11472 (N_11472,N_11280,N_11288);
nor U11473 (N_11473,N_11366,N_11319);
nand U11474 (N_11474,N_11290,N_11371);
nand U11475 (N_11475,N_11357,N_11382);
or U11476 (N_11476,N_11398,N_11360);
or U11477 (N_11477,N_11280,N_11296);
nand U11478 (N_11478,N_11359,N_11369);
xnor U11479 (N_11479,N_11260,N_11303);
nand U11480 (N_11480,N_11319,N_11358);
and U11481 (N_11481,N_11330,N_11334);
nand U11482 (N_11482,N_11340,N_11297);
and U11483 (N_11483,N_11265,N_11277);
xor U11484 (N_11484,N_11348,N_11310);
or U11485 (N_11485,N_11277,N_11319);
xnor U11486 (N_11486,N_11276,N_11327);
nor U11487 (N_11487,N_11331,N_11325);
and U11488 (N_11488,N_11319,N_11389);
nor U11489 (N_11489,N_11255,N_11266);
nand U11490 (N_11490,N_11310,N_11278);
and U11491 (N_11491,N_11368,N_11381);
and U11492 (N_11492,N_11318,N_11384);
nor U11493 (N_11493,N_11295,N_11261);
nand U11494 (N_11494,N_11309,N_11275);
nand U11495 (N_11495,N_11376,N_11371);
nor U11496 (N_11496,N_11331,N_11351);
nand U11497 (N_11497,N_11358,N_11277);
and U11498 (N_11498,N_11386,N_11288);
and U11499 (N_11499,N_11307,N_11383);
or U11500 (N_11500,N_11318,N_11376);
nand U11501 (N_11501,N_11301,N_11387);
or U11502 (N_11502,N_11362,N_11274);
nand U11503 (N_11503,N_11358,N_11343);
or U11504 (N_11504,N_11384,N_11386);
and U11505 (N_11505,N_11268,N_11299);
and U11506 (N_11506,N_11326,N_11331);
and U11507 (N_11507,N_11359,N_11342);
nand U11508 (N_11508,N_11364,N_11303);
xnor U11509 (N_11509,N_11378,N_11314);
xnor U11510 (N_11510,N_11299,N_11314);
nor U11511 (N_11511,N_11313,N_11287);
and U11512 (N_11512,N_11365,N_11374);
xor U11513 (N_11513,N_11279,N_11348);
xnor U11514 (N_11514,N_11378,N_11331);
nand U11515 (N_11515,N_11278,N_11379);
nor U11516 (N_11516,N_11274,N_11346);
xor U11517 (N_11517,N_11343,N_11396);
or U11518 (N_11518,N_11303,N_11256);
or U11519 (N_11519,N_11381,N_11294);
nand U11520 (N_11520,N_11334,N_11351);
nor U11521 (N_11521,N_11328,N_11303);
and U11522 (N_11522,N_11307,N_11286);
nor U11523 (N_11523,N_11390,N_11279);
xor U11524 (N_11524,N_11355,N_11374);
and U11525 (N_11525,N_11364,N_11386);
and U11526 (N_11526,N_11379,N_11277);
and U11527 (N_11527,N_11397,N_11303);
and U11528 (N_11528,N_11371,N_11382);
xor U11529 (N_11529,N_11328,N_11375);
xor U11530 (N_11530,N_11270,N_11300);
nor U11531 (N_11531,N_11319,N_11354);
nand U11532 (N_11532,N_11365,N_11253);
xor U11533 (N_11533,N_11261,N_11319);
or U11534 (N_11534,N_11382,N_11370);
nor U11535 (N_11535,N_11297,N_11326);
nand U11536 (N_11536,N_11280,N_11334);
or U11537 (N_11537,N_11347,N_11285);
and U11538 (N_11538,N_11332,N_11376);
nand U11539 (N_11539,N_11321,N_11348);
and U11540 (N_11540,N_11265,N_11336);
xnor U11541 (N_11541,N_11262,N_11377);
and U11542 (N_11542,N_11288,N_11393);
and U11543 (N_11543,N_11293,N_11286);
nand U11544 (N_11544,N_11389,N_11277);
nor U11545 (N_11545,N_11291,N_11296);
nor U11546 (N_11546,N_11279,N_11328);
nor U11547 (N_11547,N_11395,N_11254);
or U11548 (N_11548,N_11265,N_11314);
and U11549 (N_11549,N_11337,N_11275);
xnor U11550 (N_11550,N_11486,N_11406);
or U11551 (N_11551,N_11502,N_11467);
xor U11552 (N_11552,N_11537,N_11470);
nand U11553 (N_11553,N_11455,N_11506);
nand U11554 (N_11554,N_11417,N_11508);
nor U11555 (N_11555,N_11532,N_11405);
nor U11556 (N_11556,N_11438,N_11431);
and U11557 (N_11557,N_11521,N_11453);
xor U11558 (N_11558,N_11426,N_11509);
or U11559 (N_11559,N_11474,N_11473);
nand U11560 (N_11560,N_11476,N_11493);
nor U11561 (N_11561,N_11544,N_11513);
or U11562 (N_11562,N_11535,N_11400);
nand U11563 (N_11563,N_11429,N_11463);
nand U11564 (N_11564,N_11488,N_11549);
or U11565 (N_11565,N_11530,N_11505);
nor U11566 (N_11566,N_11545,N_11539);
xor U11567 (N_11567,N_11531,N_11424);
xnor U11568 (N_11568,N_11495,N_11543);
nor U11569 (N_11569,N_11498,N_11441);
nor U11570 (N_11570,N_11480,N_11496);
and U11571 (N_11571,N_11465,N_11501);
and U11572 (N_11572,N_11415,N_11439);
or U11573 (N_11573,N_11515,N_11477);
xor U11574 (N_11574,N_11443,N_11408);
nor U11575 (N_11575,N_11402,N_11435);
nand U11576 (N_11576,N_11514,N_11466);
xor U11577 (N_11577,N_11425,N_11460);
or U11578 (N_11578,N_11503,N_11533);
xor U11579 (N_11579,N_11540,N_11538);
and U11580 (N_11580,N_11444,N_11412);
and U11581 (N_11581,N_11511,N_11451);
nand U11582 (N_11582,N_11485,N_11418);
xnor U11583 (N_11583,N_11534,N_11423);
or U11584 (N_11584,N_11416,N_11454);
or U11585 (N_11585,N_11469,N_11411);
or U11586 (N_11586,N_11519,N_11437);
xnor U11587 (N_11587,N_11472,N_11475);
nand U11588 (N_11588,N_11548,N_11419);
xnor U11589 (N_11589,N_11432,N_11458);
or U11590 (N_11590,N_11536,N_11524);
and U11591 (N_11591,N_11457,N_11428);
or U11592 (N_11592,N_11430,N_11436);
or U11593 (N_11593,N_11479,N_11445);
or U11594 (N_11594,N_11422,N_11404);
nor U11595 (N_11595,N_11547,N_11522);
xnor U11596 (N_11596,N_11459,N_11525);
nand U11597 (N_11597,N_11403,N_11414);
or U11598 (N_11598,N_11546,N_11464);
or U11599 (N_11599,N_11489,N_11478);
nand U11600 (N_11600,N_11542,N_11484);
or U11601 (N_11601,N_11447,N_11510);
nand U11602 (N_11602,N_11452,N_11491);
nand U11603 (N_11603,N_11494,N_11499);
or U11604 (N_11604,N_11481,N_11456);
nand U11605 (N_11605,N_11462,N_11527);
nand U11606 (N_11606,N_11440,N_11448);
nand U11607 (N_11607,N_11407,N_11520);
nand U11608 (N_11608,N_11492,N_11504);
or U11609 (N_11609,N_11512,N_11517);
or U11610 (N_11610,N_11529,N_11471);
xor U11611 (N_11611,N_11500,N_11442);
xor U11612 (N_11612,N_11516,N_11507);
or U11613 (N_11613,N_11541,N_11518);
or U11614 (N_11614,N_11427,N_11410);
nand U11615 (N_11615,N_11482,N_11483);
nand U11616 (N_11616,N_11523,N_11497);
and U11617 (N_11617,N_11433,N_11421);
nor U11618 (N_11618,N_11526,N_11401);
nor U11619 (N_11619,N_11461,N_11449);
xnor U11620 (N_11620,N_11413,N_11487);
and U11621 (N_11621,N_11468,N_11434);
xor U11622 (N_11622,N_11528,N_11446);
xnor U11623 (N_11623,N_11409,N_11420);
nor U11624 (N_11624,N_11450,N_11490);
or U11625 (N_11625,N_11435,N_11490);
nand U11626 (N_11626,N_11548,N_11408);
or U11627 (N_11627,N_11464,N_11516);
nor U11628 (N_11628,N_11407,N_11492);
and U11629 (N_11629,N_11432,N_11449);
xor U11630 (N_11630,N_11444,N_11408);
or U11631 (N_11631,N_11411,N_11510);
and U11632 (N_11632,N_11501,N_11404);
nand U11633 (N_11633,N_11503,N_11429);
nor U11634 (N_11634,N_11523,N_11432);
and U11635 (N_11635,N_11416,N_11448);
xor U11636 (N_11636,N_11492,N_11541);
xor U11637 (N_11637,N_11439,N_11414);
and U11638 (N_11638,N_11473,N_11450);
and U11639 (N_11639,N_11482,N_11409);
nand U11640 (N_11640,N_11426,N_11461);
and U11641 (N_11641,N_11402,N_11487);
and U11642 (N_11642,N_11410,N_11520);
nand U11643 (N_11643,N_11496,N_11542);
or U11644 (N_11644,N_11458,N_11440);
or U11645 (N_11645,N_11484,N_11490);
xnor U11646 (N_11646,N_11456,N_11509);
or U11647 (N_11647,N_11402,N_11478);
and U11648 (N_11648,N_11541,N_11524);
and U11649 (N_11649,N_11426,N_11518);
and U11650 (N_11650,N_11541,N_11400);
and U11651 (N_11651,N_11476,N_11451);
xor U11652 (N_11652,N_11470,N_11508);
and U11653 (N_11653,N_11433,N_11447);
xnor U11654 (N_11654,N_11431,N_11428);
or U11655 (N_11655,N_11440,N_11453);
nand U11656 (N_11656,N_11494,N_11432);
nand U11657 (N_11657,N_11546,N_11461);
nor U11658 (N_11658,N_11511,N_11423);
or U11659 (N_11659,N_11461,N_11483);
and U11660 (N_11660,N_11465,N_11544);
nor U11661 (N_11661,N_11530,N_11429);
xor U11662 (N_11662,N_11423,N_11482);
or U11663 (N_11663,N_11509,N_11525);
or U11664 (N_11664,N_11464,N_11534);
and U11665 (N_11665,N_11466,N_11436);
xnor U11666 (N_11666,N_11419,N_11459);
or U11667 (N_11667,N_11442,N_11458);
nand U11668 (N_11668,N_11533,N_11506);
nand U11669 (N_11669,N_11463,N_11540);
nand U11670 (N_11670,N_11494,N_11543);
and U11671 (N_11671,N_11460,N_11527);
nand U11672 (N_11672,N_11404,N_11487);
or U11673 (N_11673,N_11483,N_11549);
and U11674 (N_11674,N_11497,N_11540);
and U11675 (N_11675,N_11522,N_11529);
or U11676 (N_11676,N_11473,N_11478);
xor U11677 (N_11677,N_11446,N_11469);
nand U11678 (N_11678,N_11481,N_11431);
and U11679 (N_11679,N_11512,N_11510);
or U11680 (N_11680,N_11530,N_11454);
nor U11681 (N_11681,N_11455,N_11443);
xor U11682 (N_11682,N_11432,N_11435);
or U11683 (N_11683,N_11484,N_11491);
nor U11684 (N_11684,N_11495,N_11530);
nor U11685 (N_11685,N_11412,N_11451);
xnor U11686 (N_11686,N_11535,N_11519);
nor U11687 (N_11687,N_11446,N_11540);
or U11688 (N_11688,N_11433,N_11498);
or U11689 (N_11689,N_11529,N_11417);
nor U11690 (N_11690,N_11492,N_11436);
or U11691 (N_11691,N_11440,N_11452);
or U11692 (N_11692,N_11536,N_11403);
and U11693 (N_11693,N_11538,N_11481);
or U11694 (N_11694,N_11460,N_11403);
xor U11695 (N_11695,N_11494,N_11449);
xnor U11696 (N_11696,N_11412,N_11477);
xor U11697 (N_11697,N_11409,N_11522);
xor U11698 (N_11698,N_11527,N_11453);
and U11699 (N_11699,N_11549,N_11435);
nand U11700 (N_11700,N_11577,N_11579);
or U11701 (N_11701,N_11665,N_11648);
or U11702 (N_11702,N_11682,N_11611);
nand U11703 (N_11703,N_11610,N_11556);
nand U11704 (N_11704,N_11661,N_11681);
xor U11705 (N_11705,N_11573,N_11602);
or U11706 (N_11706,N_11576,N_11569);
or U11707 (N_11707,N_11596,N_11564);
xor U11708 (N_11708,N_11687,N_11571);
xor U11709 (N_11709,N_11679,N_11590);
xor U11710 (N_11710,N_11654,N_11694);
nand U11711 (N_11711,N_11572,N_11696);
nor U11712 (N_11712,N_11608,N_11589);
nand U11713 (N_11713,N_11593,N_11652);
nand U11714 (N_11714,N_11617,N_11616);
and U11715 (N_11715,N_11620,N_11587);
xor U11716 (N_11716,N_11632,N_11680);
xor U11717 (N_11717,N_11603,N_11636);
or U11718 (N_11718,N_11634,N_11685);
nand U11719 (N_11719,N_11689,N_11582);
or U11720 (N_11720,N_11633,N_11618);
or U11721 (N_11721,N_11657,N_11619);
and U11722 (N_11722,N_11683,N_11672);
or U11723 (N_11723,N_11565,N_11669);
nor U11724 (N_11724,N_11660,N_11604);
nor U11725 (N_11725,N_11585,N_11613);
nor U11726 (N_11726,N_11676,N_11686);
nand U11727 (N_11727,N_11625,N_11615);
nand U11728 (N_11728,N_11640,N_11612);
nor U11729 (N_11729,N_11562,N_11626);
nand U11730 (N_11730,N_11688,N_11675);
nand U11731 (N_11731,N_11555,N_11651);
xnor U11732 (N_11732,N_11597,N_11677);
nor U11733 (N_11733,N_11635,N_11639);
nor U11734 (N_11734,N_11666,N_11650);
or U11735 (N_11735,N_11624,N_11638);
and U11736 (N_11736,N_11667,N_11693);
nand U11737 (N_11737,N_11588,N_11559);
nor U11738 (N_11738,N_11691,N_11578);
nand U11739 (N_11739,N_11567,N_11600);
xor U11740 (N_11740,N_11557,N_11697);
and U11741 (N_11741,N_11649,N_11643);
and U11742 (N_11742,N_11553,N_11606);
nor U11743 (N_11743,N_11646,N_11658);
nand U11744 (N_11744,N_11674,N_11629);
and U11745 (N_11745,N_11628,N_11656);
xor U11746 (N_11746,N_11575,N_11598);
xnor U11747 (N_11747,N_11601,N_11614);
nor U11748 (N_11748,N_11570,N_11631);
xor U11749 (N_11749,N_11623,N_11645);
or U11750 (N_11750,N_11695,N_11655);
or U11751 (N_11751,N_11684,N_11690);
and U11752 (N_11752,N_11599,N_11580);
and U11753 (N_11753,N_11698,N_11641);
nor U11754 (N_11754,N_11678,N_11550);
and U11755 (N_11755,N_11692,N_11552);
and U11756 (N_11756,N_11592,N_11568);
nand U11757 (N_11757,N_11595,N_11662);
and U11758 (N_11758,N_11558,N_11607);
nand U11759 (N_11759,N_11581,N_11609);
xnor U11760 (N_11760,N_11594,N_11566);
nand U11761 (N_11761,N_11583,N_11584);
and U11762 (N_11762,N_11591,N_11673);
nor U11763 (N_11763,N_11663,N_11621);
and U11764 (N_11764,N_11670,N_11699);
or U11765 (N_11765,N_11586,N_11653);
nand U11766 (N_11766,N_11561,N_11627);
or U11767 (N_11767,N_11563,N_11642);
and U11768 (N_11768,N_11605,N_11630);
nand U11769 (N_11769,N_11647,N_11644);
and U11770 (N_11770,N_11554,N_11659);
or U11771 (N_11771,N_11664,N_11622);
nand U11772 (N_11772,N_11671,N_11574);
or U11773 (N_11773,N_11551,N_11668);
or U11774 (N_11774,N_11560,N_11637);
nor U11775 (N_11775,N_11642,N_11564);
or U11776 (N_11776,N_11610,N_11613);
nand U11777 (N_11777,N_11617,N_11596);
and U11778 (N_11778,N_11564,N_11698);
xor U11779 (N_11779,N_11677,N_11567);
or U11780 (N_11780,N_11552,N_11619);
nor U11781 (N_11781,N_11642,N_11658);
nor U11782 (N_11782,N_11642,N_11677);
or U11783 (N_11783,N_11682,N_11692);
nand U11784 (N_11784,N_11582,N_11653);
nand U11785 (N_11785,N_11570,N_11554);
and U11786 (N_11786,N_11667,N_11553);
and U11787 (N_11787,N_11691,N_11684);
xnor U11788 (N_11788,N_11615,N_11677);
nor U11789 (N_11789,N_11655,N_11600);
and U11790 (N_11790,N_11598,N_11646);
and U11791 (N_11791,N_11651,N_11551);
nor U11792 (N_11792,N_11571,N_11575);
or U11793 (N_11793,N_11637,N_11605);
nor U11794 (N_11794,N_11676,N_11690);
or U11795 (N_11795,N_11603,N_11668);
nor U11796 (N_11796,N_11652,N_11581);
nor U11797 (N_11797,N_11678,N_11603);
nand U11798 (N_11798,N_11650,N_11633);
or U11799 (N_11799,N_11637,N_11649);
and U11800 (N_11800,N_11593,N_11621);
nand U11801 (N_11801,N_11613,N_11697);
nor U11802 (N_11802,N_11574,N_11621);
nor U11803 (N_11803,N_11656,N_11644);
nand U11804 (N_11804,N_11584,N_11656);
xor U11805 (N_11805,N_11659,N_11677);
nor U11806 (N_11806,N_11667,N_11617);
or U11807 (N_11807,N_11567,N_11580);
or U11808 (N_11808,N_11562,N_11573);
or U11809 (N_11809,N_11697,N_11602);
xnor U11810 (N_11810,N_11683,N_11556);
or U11811 (N_11811,N_11590,N_11585);
and U11812 (N_11812,N_11604,N_11640);
nor U11813 (N_11813,N_11622,N_11620);
nor U11814 (N_11814,N_11610,N_11565);
and U11815 (N_11815,N_11628,N_11665);
xor U11816 (N_11816,N_11699,N_11629);
nand U11817 (N_11817,N_11674,N_11579);
and U11818 (N_11818,N_11609,N_11676);
nor U11819 (N_11819,N_11588,N_11602);
or U11820 (N_11820,N_11699,N_11651);
or U11821 (N_11821,N_11658,N_11577);
nor U11822 (N_11822,N_11602,N_11553);
nor U11823 (N_11823,N_11576,N_11554);
xor U11824 (N_11824,N_11571,N_11698);
nand U11825 (N_11825,N_11668,N_11686);
or U11826 (N_11826,N_11584,N_11552);
or U11827 (N_11827,N_11583,N_11681);
and U11828 (N_11828,N_11607,N_11603);
nor U11829 (N_11829,N_11598,N_11573);
and U11830 (N_11830,N_11619,N_11575);
and U11831 (N_11831,N_11622,N_11685);
and U11832 (N_11832,N_11660,N_11658);
xnor U11833 (N_11833,N_11622,N_11576);
and U11834 (N_11834,N_11573,N_11673);
nand U11835 (N_11835,N_11652,N_11586);
or U11836 (N_11836,N_11604,N_11634);
or U11837 (N_11837,N_11625,N_11596);
or U11838 (N_11838,N_11585,N_11691);
and U11839 (N_11839,N_11563,N_11689);
nand U11840 (N_11840,N_11611,N_11676);
or U11841 (N_11841,N_11589,N_11568);
nand U11842 (N_11842,N_11556,N_11699);
nor U11843 (N_11843,N_11572,N_11653);
nor U11844 (N_11844,N_11697,N_11570);
xnor U11845 (N_11845,N_11596,N_11594);
nand U11846 (N_11846,N_11570,N_11569);
nor U11847 (N_11847,N_11558,N_11672);
nand U11848 (N_11848,N_11594,N_11620);
and U11849 (N_11849,N_11678,N_11632);
xnor U11850 (N_11850,N_11802,N_11809);
nand U11851 (N_11851,N_11738,N_11726);
nor U11852 (N_11852,N_11791,N_11748);
xnor U11853 (N_11853,N_11832,N_11731);
xnor U11854 (N_11854,N_11828,N_11811);
nor U11855 (N_11855,N_11757,N_11778);
nor U11856 (N_11856,N_11849,N_11827);
nor U11857 (N_11857,N_11761,N_11835);
xor U11858 (N_11858,N_11847,N_11739);
nand U11859 (N_11859,N_11705,N_11775);
nand U11860 (N_11860,N_11789,N_11727);
nor U11861 (N_11861,N_11808,N_11725);
nor U11862 (N_11862,N_11829,N_11764);
xnor U11863 (N_11863,N_11821,N_11774);
or U11864 (N_11864,N_11734,N_11711);
nor U11865 (N_11865,N_11744,N_11767);
nand U11866 (N_11866,N_11760,N_11801);
nor U11867 (N_11867,N_11756,N_11784);
and U11868 (N_11868,N_11845,N_11790);
nor U11869 (N_11869,N_11795,N_11842);
or U11870 (N_11870,N_11836,N_11701);
nand U11871 (N_11871,N_11702,N_11735);
nand U11872 (N_11872,N_11742,N_11817);
xnor U11873 (N_11873,N_11839,N_11810);
nand U11874 (N_11874,N_11770,N_11848);
nor U11875 (N_11875,N_11806,N_11723);
nand U11876 (N_11876,N_11834,N_11721);
nor U11877 (N_11877,N_11743,N_11716);
and U11878 (N_11878,N_11754,N_11786);
nor U11879 (N_11879,N_11780,N_11812);
and U11880 (N_11880,N_11749,N_11703);
and U11881 (N_11881,N_11841,N_11814);
nand U11882 (N_11882,N_11793,N_11720);
nand U11883 (N_11883,N_11722,N_11712);
xnor U11884 (N_11884,N_11805,N_11782);
xor U11885 (N_11885,N_11771,N_11838);
and U11886 (N_11886,N_11816,N_11830);
nand U11887 (N_11887,N_11792,N_11718);
nor U11888 (N_11888,N_11755,N_11825);
nor U11889 (N_11889,N_11730,N_11773);
nor U11890 (N_11890,N_11704,N_11788);
nor U11891 (N_11891,N_11762,N_11844);
nand U11892 (N_11892,N_11846,N_11840);
and U11893 (N_11893,N_11803,N_11785);
nor U11894 (N_11894,N_11800,N_11724);
or U11895 (N_11895,N_11750,N_11700);
xor U11896 (N_11896,N_11797,N_11807);
or U11897 (N_11897,N_11719,N_11798);
or U11898 (N_11898,N_11781,N_11787);
xnor U11899 (N_11899,N_11833,N_11729);
or U11900 (N_11900,N_11794,N_11737);
nor U11901 (N_11901,N_11752,N_11713);
nand U11902 (N_11902,N_11824,N_11818);
nand U11903 (N_11903,N_11733,N_11741);
or U11904 (N_11904,N_11768,N_11747);
and U11905 (N_11905,N_11732,N_11769);
nor U11906 (N_11906,N_11815,N_11843);
and U11907 (N_11907,N_11710,N_11709);
and U11908 (N_11908,N_11714,N_11819);
nor U11909 (N_11909,N_11751,N_11779);
nor U11910 (N_11910,N_11783,N_11813);
and U11911 (N_11911,N_11826,N_11822);
xnor U11912 (N_11912,N_11746,N_11776);
nand U11913 (N_11913,N_11708,N_11736);
xor U11914 (N_11914,N_11715,N_11740);
and U11915 (N_11915,N_11758,N_11753);
nor U11916 (N_11916,N_11837,N_11766);
or U11917 (N_11917,N_11759,N_11796);
and U11918 (N_11918,N_11804,N_11717);
or U11919 (N_11919,N_11823,N_11799);
or U11920 (N_11920,N_11707,N_11728);
and U11921 (N_11921,N_11706,N_11820);
xnor U11922 (N_11922,N_11772,N_11763);
or U11923 (N_11923,N_11777,N_11765);
and U11924 (N_11924,N_11831,N_11745);
xor U11925 (N_11925,N_11770,N_11701);
nand U11926 (N_11926,N_11741,N_11785);
nor U11927 (N_11927,N_11786,N_11818);
nor U11928 (N_11928,N_11806,N_11816);
nor U11929 (N_11929,N_11752,N_11842);
and U11930 (N_11930,N_11768,N_11834);
nand U11931 (N_11931,N_11829,N_11837);
or U11932 (N_11932,N_11787,N_11838);
or U11933 (N_11933,N_11734,N_11730);
nor U11934 (N_11934,N_11835,N_11736);
or U11935 (N_11935,N_11797,N_11739);
or U11936 (N_11936,N_11790,N_11726);
or U11937 (N_11937,N_11728,N_11817);
nor U11938 (N_11938,N_11826,N_11760);
xor U11939 (N_11939,N_11824,N_11840);
and U11940 (N_11940,N_11774,N_11768);
nor U11941 (N_11941,N_11815,N_11703);
xor U11942 (N_11942,N_11823,N_11779);
nand U11943 (N_11943,N_11805,N_11729);
nor U11944 (N_11944,N_11836,N_11803);
xnor U11945 (N_11945,N_11830,N_11826);
nand U11946 (N_11946,N_11712,N_11758);
or U11947 (N_11947,N_11810,N_11725);
nand U11948 (N_11948,N_11790,N_11753);
or U11949 (N_11949,N_11747,N_11764);
nor U11950 (N_11950,N_11740,N_11819);
nor U11951 (N_11951,N_11711,N_11733);
or U11952 (N_11952,N_11829,N_11752);
nor U11953 (N_11953,N_11772,N_11802);
or U11954 (N_11954,N_11796,N_11732);
nand U11955 (N_11955,N_11786,N_11819);
xnor U11956 (N_11956,N_11707,N_11846);
and U11957 (N_11957,N_11733,N_11823);
nand U11958 (N_11958,N_11753,N_11784);
nor U11959 (N_11959,N_11750,N_11810);
nor U11960 (N_11960,N_11753,N_11815);
nand U11961 (N_11961,N_11712,N_11704);
and U11962 (N_11962,N_11747,N_11842);
and U11963 (N_11963,N_11709,N_11716);
nor U11964 (N_11964,N_11800,N_11727);
nand U11965 (N_11965,N_11787,N_11770);
nor U11966 (N_11966,N_11776,N_11737);
and U11967 (N_11967,N_11745,N_11735);
nor U11968 (N_11968,N_11818,N_11704);
and U11969 (N_11969,N_11833,N_11762);
xor U11970 (N_11970,N_11742,N_11788);
nor U11971 (N_11971,N_11790,N_11731);
nand U11972 (N_11972,N_11830,N_11736);
and U11973 (N_11973,N_11756,N_11718);
nor U11974 (N_11974,N_11729,N_11807);
and U11975 (N_11975,N_11772,N_11835);
and U11976 (N_11976,N_11728,N_11818);
nor U11977 (N_11977,N_11723,N_11765);
nor U11978 (N_11978,N_11827,N_11793);
or U11979 (N_11979,N_11840,N_11847);
and U11980 (N_11980,N_11738,N_11803);
and U11981 (N_11981,N_11717,N_11774);
and U11982 (N_11982,N_11831,N_11789);
nand U11983 (N_11983,N_11774,N_11772);
nor U11984 (N_11984,N_11758,N_11772);
and U11985 (N_11985,N_11824,N_11795);
nand U11986 (N_11986,N_11727,N_11816);
nand U11987 (N_11987,N_11736,N_11791);
xor U11988 (N_11988,N_11827,N_11805);
xor U11989 (N_11989,N_11830,N_11700);
nor U11990 (N_11990,N_11721,N_11706);
xnor U11991 (N_11991,N_11787,N_11779);
or U11992 (N_11992,N_11758,N_11714);
nor U11993 (N_11993,N_11710,N_11805);
nor U11994 (N_11994,N_11736,N_11834);
nor U11995 (N_11995,N_11847,N_11814);
or U11996 (N_11996,N_11796,N_11794);
and U11997 (N_11997,N_11803,N_11782);
and U11998 (N_11998,N_11774,N_11804);
and U11999 (N_11999,N_11701,N_11793);
or U12000 (N_12000,N_11894,N_11927);
nor U12001 (N_12001,N_11913,N_11867);
nor U12002 (N_12002,N_11854,N_11943);
xnor U12003 (N_12003,N_11874,N_11925);
nand U12004 (N_12004,N_11972,N_11953);
and U12005 (N_12005,N_11862,N_11952);
xnor U12006 (N_12006,N_11858,N_11850);
nor U12007 (N_12007,N_11877,N_11869);
nor U12008 (N_12008,N_11895,N_11965);
nand U12009 (N_12009,N_11963,N_11992);
nand U12010 (N_12010,N_11900,N_11999);
nor U12011 (N_12011,N_11866,N_11890);
or U12012 (N_12012,N_11954,N_11970);
nor U12013 (N_12013,N_11986,N_11923);
xor U12014 (N_12014,N_11956,N_11966);
nand U12015 (N_12015,N_11933,N_11909);
nor U12016 (N_12016,N_11876,N_11915);
and U12017 (N_12017,N_11924,N_11942);
or U12018 (N_12018,N_11980,N_11865);
or U12019 (N_12019,N_11975,N_11961);
xor U12020 (N_12020,N_11872,N_11897);
nor U12021 (N_12021,N_11896,N_11993);
nor U12022 (N_12022,N_11989,N_11930);
xor U12023 (N_12023,N_11902,N_11937);
nor U12024 (N_12024,N_11916,N_11982);
nand U12025 (N_12025,N_11853,N_11983);
xnor U12026 (N_12026,N_11985,N_11957);
nor U12027 (N_12027,N_11950,N_11860);
nand U12028 (N_12028,N_11979,N_11932);
or U12029 (N_12029,N_11978,N_11907);
nor U12030 (N_12030,N_11905,N_11962);
nor U12031 (N_12031,N_11949,N_11922);
xnor U12032 (N_12032,N_11948,N_11868);
xor U12033 (N_12033,N_11873,N_11939);
xnor U12034 (N_12034,N_11852,N_11958);
nor U12035 (N_12035,N_11917,N_11981);
and U12036 (N_12036,N_11946,N_11910);
or U12037 (N_12037,N_11973,N_11855);
nand U12038 (N_12038,N_11964,N_11880);
nor U12039 (N_12039,N_11984,N_11988);
nand U12040 (N_12040,N_11884,N_11908);
or U12041 (N_12041,N_11889,N_11994);
nor U12042 (N_12042,N_11940,N_11934);
nor U12043 (N_12043,N_11903,N_11891);
or U12044 (N_12044,N_11875,N_11959);
nor U12045 (N_12045,N_11945,N_11870);
and U12046 (N_12046,N_11859,N_11995);
nand U12047 (N_12047,N_11861,N_11892);
nor U12048 (N_12048,N_11990,N_11938);
or U12049 (N_12049,N_11914,N_11871);
nand U12050 (N_12050,N_11991,N_11974);
xnor U12051 (N_12051,N_11960,N_11918);
nor U12052 (N_12052,N_11912,N_11882);
nand U12053 (N_12053,N_11967,N_11899);
or U12054 (N_12054,N_11969,N_11951);
xor U12055 (N_12055,N_11863,N_11936);
nor U12056 (N_12056,N_11931,N_11906);
and U12057 (N_12057,N_11935,N_11864);
nor U12058 (N_12058,N_11885,N_11976);
xor U12059 (N_12059,N_11941,N_11997);
xnor U12060 (N_12060,N_11944,N_11883);
or U12061 (N_12061,N_11887,N_11898);
or U12062 (N_12062,N_11921,N_11888);
xnor U12063 (N_12063,N_11987,N_11886);
and U12064 (N_12064,N_11929,N_11851);
xnor U12065 (N_12065,N_11878,N_11881);
xor U12066 (N_12066,N_11968,N_11947);
xor U12067 (N_12067,N_11955,N_11977);
xnor U12068 (N_12068,N_11928,N_11919);
nor U12069 (N_12069,N_11856,N_11893);
and U12070 (N_12070,N_11901,N_11920);
or U12071 (N_12071,N_11857,N_11971);
nand U12072 (N_12072,N_11879,N_11926);
xnor U12073 (N_12073,N_11996,N_11911);
and U12074 (N_12074,N_11904,N_11998);
nor U12075 (N_12075,N_11950,N_11996);
and U12076 (N_12076,N_11875,N_11934);
nand U12077 (N_12077,N_11940,N_11952);
and U12078 (N_12078,N_11997,N_11988);
nor U12079 (N_12079,N_11938,N_11887);
xnor U12080 (N_12080,N_11852,N_11993);
nand U12081 (N_12081,N_11877,N_11921);
nand U12082 (N_12082,N_11866,N_11924);
nor U12083 (N_12083,N_11943,N_11940);
xnor U12084 (N_12084,N_11888,N_11919);
or U12085 (N_12085,N_11912,N_11922);
or U12086 (N_12086,N_11928,N_11872);
nor U12087 (N_12087,N_11965,N_11898);
nand U12088 (N_12088,N_11874,N_11997);
nor U12089 (N_12089,N_11907,N_11944);
xnor U12090 (N_12090,N_11953,N_11891);
xor U12091 (N_12091,N_11883,N_11967);
xnor U12092 (N_12092,N_11909,N_11856);
xnor U12093 (N_12093,N_11996,N_11946);
nand U12094 (N_12094,N_11852,N_11968);
and U12095 (N_12095,N_11855,N_11996);
nor U12096 (N_12096,N_11869,N_11961);
and U12097 (N_12097,N_11906,N_11853);
and U12098 (N_12098,N_11965,N_11917);
xor U12099 (N_12099,N_11889,N_11938);
and U12100 (N_12100,N_11933,N_11924);
or U12101 (N_12101,N_11978,N_11984);
and U12102 (N_12102,N_11915,N_11934);
nand U12103 (N_12103,N_11916,N_11911);
and U12104 (N_12104,N_11928,N_11932);
nand U12105 (N_12105,N_11923,N_11982);
nand U12106 (N_12106,N_11991,N_11853);
and U12107 (N_12107,N_11976,N_11949);
and U12108 (N_12108,N_11916,N_11917);
and U12109 (N_12109,N_11898,N_11941);
and U12110 (N_12110,N_11896,N_11946);
nor U12111 (N_12111,N_11915,N_11887);
or U12112 (N_12112,N_11869,N_11979);
or U12113 (N_12113,N_11857,N_11903);
nand U12114 (N_12114,N_11894,N_11906);
nand U12115 (N_12115,N_11897,N_11891);
nor U12116 (N_12116,N_11960,N_11944);
xnor U12117 (N_12117,N_11894,N_11986);
and U12118 (N_12118,N_11958,N_11893);
and U12119 (N_12119,N_11901,N_11885);
and U12120 (N_12120,N_11940,N_11856);
xnor U12121 (N_12121,N_11977,N_11943);
nand U12122 (N_12122,N_11853,N_11918);
nand U12123 (N_12123,N_11875,N_11937);
nand U12124 (N_12124,N_11952,N_11991);
xnor U12125 (N_12125,N_11873,N_11961);
or U12126 (N_12126,N_11953,N_11979);
xnor U12127 (N_12127,N_11887,N_11903);
nand U12128 (N_12128,N_11885,N_11989);
and U12129 (N_12129,N_11919,N_11885);
xnor U12130 (N_12130,N_11907,N_11885);
xor U12131 (N_12131,N_11956,N_11987);
and U12132 (N_12132,N_11863,N_11897);
nor U12133 (N_12133,N_11890,N_11851);
or U12134 (N_12134,N_11936,N_11962);
nor U12135 (N_12135,N_11903,N_11988);
or U12136 (N_12136,N_11851,N_11861);
or U12137 (N_12137,N_11870,N_11854);
or U12138 (N_12138,N_11918,N_11911);
or U12139 (N_12139,N_11978,N_11908);
nand U12140 (N_12140,N_11973,N_11857);
and U12141 (N_12141,N_11920,N_11863);
nor U12142 (N_12142,N_11855,N_11876);
nor U12143 (N_12143,N_11985,N_11976);
xor U12144 (N_12144,N_11855,N_11907);
or U12145 (N_12145,N_11877,N_11857);
or U12146 (N_12146,N_11868,N_11939);
or U12147 (N_12147,N_11861,N_11873);
xnor U12148 (N_12148,N_11888,N_11913);
or U12149 (N_12149,N_11943,N_11898);
xor U12150 (N_12150,N_12095,N_12082);
xnor U12151 (N_12151,N_12060,N_12106);
xnor U12152 (N_12152,N_12100,N_12023);
or U12153 (N_12153,N_12133,N_12038);
nor U12154 (N_12154,N_12016,N_12053);
or U12155 (N_12155,N_12065,N_12092);
xnor U12156 (N_12156,N_12110,N_12113);
nand U12157 (N_12157,N_12034,N_12037);
nor U12158 (N_12158,N_12003,N_12012);
nor U12159 (N_12159,N_12117,N_12145);
xnor U12160 (N_12160,N_12088,N_12134);
or U12161 (N_12161,N_12099,N_12090);
and U12162 (N_12162,N_12098,N_12124);
nor U12163 (N_12163,N_12131,N_12109);
and U12164 (N_12164,N_12096,N_12148);
nand U12165 (N_12165,N_12043,N_12105);
nand U12166 (N_12166,N_12078,N_12121);
and U12167 (N_12167,N_12130,N_12044);
and U12168 (N_12168,N_12138,N_12141);
nand U12169 (N_12169,N_12135,N_12018);
xor U12170 (N_12170,N_12108,N_12123);
or U12171 (N_12171,N_12027,N_12051);
nand U12172 (N_12172,N_12097,N_12064);
and U12173 (N_12173,N_12102,N_12070);
xor U12174 (N_12174,N_12052,N_12025);
xnor U12175 (N_12175,N_12143,N_12068);
nand U12176 (N_12176,N_12001,N_12031);
nor U12177 (N_12177,N_12040,N_12081);
xnor U12178 (N_12178,N_12146,N_12014);
or U12179 (N_12179,N_12039,N_12072);
nor U12180 (N_12180,N_12029,N_12017);
nand U12181 (N_12181,N_12119,N_12115);
or U12182 (N_12182,N_12036,N_12005);
nand U12183 (N_12183,N_12028,N_12104);
nand U12184 (N_12184,N_12047,N_12076);
or U12185 (N_12185,N_12055,N_12144);
nor U12186 (N_12186,N_12139,N_12042);
or U12187 (N_12187,N_12132,N_12009);
nand U12188 (N_12188,N_12054,N_12136);
and U12189 (N_12189,N_12063,N_12008);
nand U12190 (N_12190,N_12022,N_12007);
nor U12191 (N_12191,N_12061,N_12084);
nand U12192 (N_12192,N_12062,N_12056);
and U12193 (N_12193,N_12066,N_12122);
xor U12194 (N_12194,N_12024,N_12006);
xnor U12195 (N_12195,N_12010,N_12125);
nand U12196 (N_12196,N_12026,N_12067);
nand U12197 (N_12197,N_12118,N_12059);
nand U12198 (N_12198,N_12019,N_12149);
nor U12199 (N_12199,N_12079,N_12000);
or U12200 (N_12200,N_12069,N_12049);
nor U12201 (N_12201,N_12091,N_12058);
nor U12202 (N_12202,N_12041,N_12089);
nand U12203 (N_12203,N_12093,N_12083);
nand U12204 (N_12204,N_12114,N_12004);
nand U12205 (N_12205,N_12075,N_12103);
nor U12206 (N_12206,N_12035,N_12080);
xnor U12207 (N_12207,N_12086,N_12011);
nor U12208 (N_12208,N_12087,N_12046);
nor U12209 (N_12209,N_12073,N_12074);
nand U12210 (N_12210,N_12126,N_12127);
nand U12211 (N_12211,N_12094,N_12013);
and U12212 (N_12212,N_12015,N_12142);
or U12213 (N_12213,N_12116,N_12107);
and U12214 (N_12214,N_12033,N_12101);
nand U12215 (N_12215,N_12057,N_12021);
nand U12216 (N_12216,N_12020,N_12112);
nand U12217 (N_12217,N_12032,N_12140);
xnor U12218 (N_12218,N_12050,N_12030);
nand U12219 (N_12219,N_12085,N_12120);
or U12220 (N_12220,N_12129,N_12147);
nor U12221 (N_12221,N_12045,N_12002);
nand U12222 (N_12222,N_12128,N_12111);
xor U12223 (N_12223,N_12077,N_12048);
or U12224 (N_12224,N_12071,N_12137);
nand U12225 (N_12225,N_12110,N_12103);
and U12226 (N_12226,N_12143,N_12085);
xnor U12227 (N_12227,N_12029,N_12041);
and U12228 (N_12228,N_12064,N_12084);
and U12229 (N_12229,N_12116,N_12023);
nand U12230 (N_12230,N_12149,N_12061);
nand U12231 (N_12231,N_12093,N_12035);
xor U12232 (N_12232,N_12130,N_12067);
nor U12233 (N_12233,N_12075,N_12063);
nor U12234 (N_12234,N_12104,N_12144);
and U12235 (N_12235,N_12144,N_12052);
and U12236 (N_12236,N_12065,N_12126);
and U12237 (N_12237,N_12087,N_12042);
nor U12238 (N_12238,N_12137,N_12088);
nor U12239 (N_12239,N_12002,N_12132);
nor U12240 (N_12240,N_12032,N_12138);
nand U12241 (N_12241,N_12022,N_12112);
and U12242 (N_12242,N_12037,N_12094);
and U12243 (N_12243,N_12006,N_12009);
nand U12244 (N_12244,N_12056,N_12012);
or U12245 (N_12245,N_12148,N_12019);
xor U12246 (N_12246,N_12065,N_12023);
xor U12247 (N_12247,N_12016,N_12081);
nor U12248 (N_12248,N_12085,N_12016);
nand U12249 (N_12249,N_12121,N_12091);
nand U12250 (N_12250,N_12121,N_12097);
nor U12251 (N_12251,N_12065,N_12012);
nor U12252 (N_12252,N_12079,N_12131);
and U12253 (N_12253,N_12000,N_12095);
nand U12254 (N_12254,N_12046,N_12030);
nor U12255 (N_12255,N_12016,N_12026);
nand U12256 (N_12256,N_12022,N_12073);
nand U12257 (N_12257,N_12143,N_12083);
and U12258 (N_12258,N_12093,N_12119);
and U12259 (N_12259,N_12135,N_12022);
or U12260 (N_12260,N_12111,N_12109);
xor U12261 (N_12261,N_12006,N_12081);
xor U12262 (N_12262,N_12034,N_12005);
nor U12263 (N_12263,N_12098,N_12143);
xnor U12264 (N_12264,N_12030,N_12069);
nor U12265 (N_12265,N_12110,N_12044);
nor U12266 (N_12266,N_12122,N_12026);
nand U12267 (N_12267,N_12139,N_12050);
nor U12268 (N_12268,N_12029,N_12003);
and U12269 (N_12269,N_12078,N_12057);
xor U12270 (N_12270,N_12023,N_12139);
nand U12271 (N_12271,N_12122,N_12029);
nor U12272 (N_12272,N_12002,N_12098);
and U12273 (N_12273,N_12012,N_12130);
nor U12274 (N_12274,N_12077,N_12145);
or U12275 (N_12275,N_12133,N_12148);
or U12276 (N_12276,N_12079,N_12077);
or U12277 (N_12277,N_12146,N_12005);
nand U12278 (N_12278,N_12006,N_12019);
xor U12279 (N_12279,N_12086,N_12111);
xnor U12280 (N_12280,N_12057,N_12052);
and U12281 (N_12281,N_12091,N_12119);
xnor U12282 (N_12282,N_12103,N_12043);
and U12283 (N_12283,N_12079,N_12088);
or U12284 (N_12284,N_12112,N_12023);
and U12285 (N_12285,N_12091,N_12062);
and U12286 (N_12286,N_12098,N_12017);
nor U12287 (N_12287,N_12074,N_12020);
xor U12288 (N_12288,N_12116,N_12127);
xnor U12289 (N_12289,N_12060,N_12141);
nor U12290 (N_12290,N_12072,N_12133);
and U12291 (N_12291,N_12106,N_12104);
or U12292 (N_12292,N_12055,N_12042);
or U12293 (N_12293,N_12088,N_12045);
nand U12294 (N_12294,N_12013,N_12073);
xnor U12295 (N_12295,N_12065,N_12074);
xnor U12296 (N_12296,N_12113,N_12083);
and U12297 (N_12297,N_12100,N_12135);
nor U12298 (N_12298,N_12094,N_12136);
nor U12299 (N_12299,N_12114,N_12112);
nand U12300 (N_12300,N_12174,N_12235);
or U12301 (N_12301,N_12204,N_12270);
or U12302 (N_12302,N_12228,N_12186);
or U12303 (N_12303,N_12259,N_12209);
xnor U12304 (N_12304,N_12285,N_12221);
or U12305 (N_12305,N_12179,N_12287);
or U12306 (N_12306,N_12260,N_12189);
and U12307 (N_12307,N_12153,N_12266);
and U12308 (N_12308,N_12190,N_12195);
nand U12309 (N_12309,N_12162,N_12196);
xor U12310 (N_12310,N_12288,N_12211);
nor U12311 (N_12311,N_12250,N_12242);
nor U12312 (N_12312,N_12281,N_12200);
nand U12313 (N_12313,N_12150,N_12166);
xnor U12314 (N_12314,N_12165,N_12220);
nand U12315 (N_12315,N_12293,N_12216);
and U12316 (N_12316,N_12255,N_12158);
xor U12317 (N_12317,N_12219,N_12208);
or U12318 (N_12318,N_12203,N_12292);
nor U12319 (N_12319,N_12249,N_12183);
and U12320 (N_12320,N_12257,N_12198);
nand U12321 (N_12321,N_12241,N_12201);
or U12322 (N_12322,N_12264,N_12262);
xor U12323 (N_12323,N_12295,N_12194);
or U12324 (N_12324,N_12230,N_12181);
nand U12325 (N_12325,N_12251,N_12298);
and U12326 (N_12326,N_12226,N_12247);
xnor U12327 (N_12327,N_12283,N_12252);
or U12328 (N_12328,N_12212,N_12157);
or U12329 (N_12329,N_12271,N_12156);
nand U12330 (N_12330,N_12289,N_12178);
or U12331 (N_12331,N_12282,N_12197);
nor U12332 (N_12332,N_12224,N_12152);
nor U12333 (N_12333,N_12294,N_12154);
xnor U12334 (N_12334,N_12248,N_12233);
nand U12335 (N_12335,N_12170,N_12199);
and U12336 (N_12336,N_12180,N_12191);
and U12337 (N_12337,N_12163,N_12243);
nor U12338 (N_12338,N_12175,N_12263);
nor U12339 (N_12339,N_12276,N_12232);
nand U12340 (N_12340,N_12164,N_12160);
and U12341 (N_12341,N_12168,N_12290);
xnor U12342 (N_12342,N_12188,N_12206);
xnor U12343 (N_12343,N_12269,N_12291);
nand U12344 (N_12344,N_12286,N_12268);
xor U12345 (N_12345,N_12278,N_12225);
or U12346 (N_12346,N_12229,N_12171);
nand U12347 (N_12347,N_12261,N_12234);
nor U12348 (N_12348,N_12237,N_12254);
nor U12349 (N_12349,N_12256,N_12185);
nor U12350 (N_12350,N_12217,N_12246);
xnor U12351 (N_12351,N_12215,N_12244);
or U12352 (N_12352,N_12245,N_12167);
xnor U12353 (N_12353,N_12159,N_12238);
xor U12354 (N_12354,N_12182,N_12192);
xnor U12355 (N_12355,N_12155,N_12231);
and U12356 (N_12356,N_12299,N_12184);
nand U12357 (N_12357,N_12239,N_12172);
or U12358 (N_12358,N_12267,N_12265);
xor U12359 (N_12359,N_12280,N_12258);
or U12360 (N_12360,N_12227,N_12213);
nand U12361 (N_12361,N_12218,N_12161);
xnor U12362 (N_12362,N_12205,N_12214);
or U12363 (N_12363,N_12273,N_12193);
nor U12364 (N_12364,N_12275,N_12176);
xnor U12365 (N_12365,N_12240,N_12202);
and U12366 (N_12366,N_12207,N_12169);
and U12367 (N_12367,N_12210,N_12279);
nor U12368 (N_12368,N_12296,N_12272);
nor U12369 (N_12369,N_12253,N_12222);
and U12370 (N_12370,N_12277,N_12177);
nor U12371 (N_12371,N_12284,N_12297);
and U12372 (N_12372,N_12151,N_12236);
or U12373 (N_12373,N_12173,N_12223);
nand U12374 (N_12374,N_12274,N_12187);
nand U12375 (N_12375,N_12190,N_12281);
and U12376 (N_12376,N_12274,N_12174);
nand U12377 (N_12377,N_12269,N_12278);
or U12378 (N_12378,N_12168,N_12240);
xor U12379 (N_12379,N_12265,N_12168);
xor U12380 (N_12380,N_12152,N_12212);
or U12381 (N_12381,N_12298,N_12230);
xnor U12382 (N_12382,N_12237,N_12153);
or U12383 (N_12383,N_12269,N_12159);
nor U12384 (N_12384,N_12297,N_12246);
nand U12385 (N_12385,N_12254,N_12198);
xnor U12386 (N_12386,N_12182,N_12154);
nor U12387 (N_12387,N_12152,N_12255);
nor U12388 (N_12388,N_12208,N_12249);
nor U12389 (N_12389,N_12264,N_12243);
nor U12390 (N_12390,N_12218,N_12176);
and U12391 (N_12391,N_12170,N_12298);
or U12392 (N_12392,N_12254,N_12289);
nand U12393 (N_12393,N_12243,N_12283);
nand U12394 (N_12394,N_12179,N_12296);
xnor U12395 (N_12395,N_12225,N_12204);
or U12396 (N_12396,N_12271,N_12252);
nor U12397 (N_12397,N_12161,N_12283);
and U12398 (N_12398,N_12187,N_12250);
nand U12399 (N_12399,N_12192,N_12159);
and U12400 (N_12400,N_12231,N_12259);
and U12401 (N_12401,N_12222,N_12261);
nor U12402 (N_12402,N_12155,N_12171);
or U12403 (N_12403,N_12190,N_12260);
nand U12404 (N_12404,N_12152,N_12175);
xnor U12405 (N_12405,N_12203,N_12218);
nand U12406 (N_12406,N_12189,N_12240);
nor U12407 (N_12407,N_12167,N_12199);
and U12408 (N_12408,N_12254,N_12207);
or U12409 (N_12409,N_12167,N_12239);
or U12410 (N_12410,N_12294,N_12266);
nor U12411 (N_12411,N_12195,N_12248);
or U12412 (N_12412,N_12157,N_12151);
nand U12413 (N_12413,N_12278,N_12193);
or U12414 (N_12414,N_12226,N_12222);
nor U12415 (N_12415,N_12298,N_12292);
nor U12416 (N_12416,N_12162,N_12150);
nor U12417 (N_12417,N_12254,N_12279);
nand U12418 (N_12418,N_12199,N_12276);
xor U12419 (N_12419,N_12183,N_12150);
nand U12420 (N_12420,N_12248,N_12200);
or U12421 (N_12421,N_12178,N_12271);
nor U12422 (N_12422,N_12232,N_12182);
nor U12423 (N_12423,N_12207,N_12271);
nor U12424 (N_12424,N_12227,N_12289);
nor U12425 (N_12425,N_12193,N_12259);
xnor U12426 (N_12426,N_12166,N_12181);
xor U12427 (N_12427,N_12161,N_12261);
nand U12428 (N_12428,N_12190,N_12271);
or U12429 (N_12429,N_12188,N_12225);
nand U12430 (N_12430,N_12217,N_12281);
nand U12431 (N_12431,N_12248,N_12159);
and U12432 (N_12432,N_12189,N_12193);
and U12433 (N_12433,N_12297,N_12275);
nor U12434 (N_12434,N_12228,N_12276);
or U12435 (N_12435,N_12284,N_12172);
nand U12436 (N_12436,N_12196,N_12293);
or U12437 (N_12437,N_12206,N_12248);
xnor U12438 (N_12438,N_12162,N_12295);
nand U12439 (N_12439,N_12178,N_12210);
or U12440 (N_12440,N_12256,N_12277);
nand U12441 (N_12441,N_12279,N_12204);
and U12442 (N_12442,N_12289,N_12167);
nor U12443 (N_12443,N_12267,N_12223);
nor U12444 (N_12444,N_12276,N_12227);
or U12445 (N_12445,N_12261,N_12157);
nand U12446 (N_12446,N_12288,N_12270);
and U12447 (N_12447,N_12219,N_12200);
and U12448 (N_12448,N_12284,N_12279);
or U12449 (N_12449,N_12295,N_12219);
and U12450 (N_12450,N_12421,N_12364);
nor U12451 (N_12451,N_12425,N_12328);
nor U12452 (N_12452,N_12304,N_12308);
and U12453 (N_12453,N_12430,N_12447);
xor U12454 (N_12454,N_12433,N_12344);
and U12455 (N_12455,N_12393,N_12377);
nand U12456 (N_12456,N_12427,N_12443);
xnor U12457 (N_12457,N_12371,N_12336);
nor U12458 (N_12458,N_12332,N_12335);
nor U12459 (N_12459,N_12424,N_12396);
and U12460 (N_12460,N_12326,N_12360);
xnor U12461 (N_12461,N_12323,N_12439);
xor U12462 (N_12462,N_12312,N_12440);
xnor U12463 (N_12463,N_12448,N_12338);
nand U12464 (N_12464,N_12366,N_12318);
nand U12465 (N_12465,N_12346,N_12317);
and U12466 (N_12466,N_12357,N_12353);
and U12467 (N_12467,N_12419,N_12356);
or U12468 (N_12468,N_12354,N_12362);
nand U12469 (N_12469,N_12417,N_12376);
and U12470 (N_12470,N_12388,N_12436);
or U12471 (N_12471,N_12413,N_12374);
nand U12472 (N_12472,N_12409,N_12408);
nand U12473 (N_12473,N_12340,N_12302);
nor U12474 (N_12474,N_12445,N_12434);
or U12475 (N_12475,N_12416,N_12390);
nand U12476 (N_12476,N_12309,N_12333);
and U12477 (N_12477,N_12387,N_12342);
nand U12478 (N_12478,N_12331,N_12442);
or U12479 (N_12479,N_12418,N_12321);
or U12480 (N_12480,N_12441,N_12389);
and U12481 (N_12481,N_12349,N_12370);
nor U12482 (N_12482,N_12301,N_12379);
or U12483 (N_12483,N_12395,N_12392);
and U12484 (N_12484,N_12345,N_12378);
nor U12485 (N_12485,N_12310,N_12423);
and U12486 (N_12486,N_12375,N_12369);
xor U12487 (N_12487,N_12407,N_12361);
nor U12488 (N_12488,N_12352,N_12400);
xor U12489 (N_12489,N_12446,N_12401);
nor U12490 (N_12490,N_12348,N_12320);
nor U12491 (N_12491,N_12324,N_12337);
or U12492 (N_12492,N_12315,N_12343);
nand U12493 (N_12493,N_12359,N_12382);
and U12494 (N_12494,N_12351,N_12411);
or U12495 (N_12495,N_12426,N_12404);
xor U12496 (N_12496,N_12319,N_12399);
xor U12497 (N_12497,N_12405,N_12347);
and U12498 (N_12498,N_12435,N_12316);
nand U12499 (N_12499,N_12412,N_12437);
nand U12500 (N_12500,N_12313,N_12420);
or U12501 (N_12501,N_12385,N_12431);
xnor U12502 (N_12502,N_12311,N_12428);
or U12503 (N_12503,N_12422,N_12329);
and U12504 (N_12504,N_12438,N_12414);
or U12505 (N_12505,N_12373,N_12384);
or U12506 (N_12506,N_12350,N_12334);
xor U12507 (N_12507,N_12363,N_12358);
xnor U12508 (N_12508,N_12383,N_12305);
xor U12509 (N_12509,N_12330,N_12386);
nand U12510 (N_12510,N_12397,N_12368);
nor U12511 (N_12511,N_12402,N_12325);
or U12512 (N_12512,N_12398,N_12432);
xnor U12513 (N_12513,N_12403,N_12365);
and U12514 (N_12514,N_12406,N_12381);
xor U12515 (N_12515,N_12300,N_12341);
nor U12516 (N_12516,N_12415,N_12372);
nor U12517 (N_12517,N_12367,N_12307);
and U12518 (N_12518,N_12314,N_12429);
and U12519 (N_12519,N_12444,N_12355);
xnor U12520 (N_12520,N_12394,N_12391);
and U12521 (N_12521,N_12449,N_12306);
nor U12522 (N_12522,N_12303,N_12410);
or U12523 (N_12523,N_12327,N_12380);
nor U12524 (N_12524,N_12339,N_12322);
nand U12525 (N_12525,N_12407,N_12324);
and U12526 (N_12526,N_12442,N_12314);
xnor U12527 (N_12527,N_12316,N_12322);
xor U12528 (N_12528,N_12393,N_12402);
xor U12529 (N_12529,N_12343,N_12429);
and U12530 (N_12530,N_12390,N_12373);
xor U12531 (N_12531,N_12337,N_12311);
or U12532 (N_12532,N_12363,N_12374);
xor U12533 (N_12533,N_12419,N_12303);
nor U12534 (N_12534,N_12430,N_12414);
nand U12535 (N_12535,N_12300,N_12303);
nand U12536 (N_12536,N_12383,N_12421);
nand U12537 (N_12537,N_12367,N_12393);
and U12538 (N_12538,N_12338,N_12331);
nand U12539 (N_12539,N_12339,N_12396);
xor U12540 (N_12540,N_12386,N_12418);
or U12541 (N_12541,N_12350,N_12344);
and U12542 (N_12542,N_12303,N_12316);
and U12543 (N_12543,N_12305,N_12327);
xor U12544 (N_12544,N_12311,N_12336);
nand U12545 (N_12545,N_12405,N_12349);
xor U12546 (N_12546,N_12305,N_12332);
xor U12547 (N_12547,N_12320,N_12400);
and U12548 (N_12548,N_12409,N_12324);
or U12549 (N_12549,N_12378,N_12360);
nor U12550 (N_12550,N_12334,N_12439);
nand U12551 (N_12551,N_12438,N_12339);
nand U12552 (N_12552,N_12335,N_12359);
xor U12553 (N_12553,N_12421,N_12351);
and U12554 (N_12554,N_12389,N_12366);
nor U12555 (N_12555,N_12425,N_12435);
nand U12556 (N_12556,N_12421,N_12347);
nand U12557 (N_12557,N_12437,N_12321);
xor U12558 (N_12558,N_12420,N_12359);
nor U12559 (N_12559,N_12320,N_12406);
nor U12560 (N_12560,N_12374,N_12384);
nand U12561 (N_12561,N_12356,N_12318);
xor U12562 (N_12562,N_12393,N_12333);
nor U12563 (N_12563,N_12422,N_12395);
xor U12564 (N_12564,N_12363,N_12425);
or U12565 (N_12565,N_12352,N_12427);
nor U12566 (N_12566,N_12349,N_12317);
nor U12567 (N_12567,N_12327,N_12396);
or U12568 (N_12568,N_12415,N_12357);
xnor U12569 (N_12569,N_12358,N_12366);
nand U12570 (N_12570,N_12369,N_12358);
nand U12571 (N_12571,N_12308,N_12359);
xor U12572 (N_12572,N_12363,N_12377);
or U12573 (N_12573,N_12316,N_12324);
xnor U12574 (N_12574,N_12304,N_12413);
nor U12575 (N_12575,N_12435,N_12332);
and U12576 (N_12576,N_12310,N_12312);
nand U12577 (N_12577,N_12355,N_12428);
or U12578 (N_12578,N_12387,N_12343);
nor U12579 (N_12579,N_12301,N_12338);
nand U12580 (N_12580,N_12317,N_12314);
nor U12581 (N_12581,N_12341,N_12346);
xnor U12582 (N_12582,N_12402,N_12438);
and U12583 (N_12583,N_12446,N_12347);
or U12584 (N_12584,N_12353,N_12310);
nand U12585 (N_12585,N_12348,N_12387);
xor U12586 (N_12586,N_12353,N_12396);
nand U12587 (N_12587,N_12418,N_12416);
nand U12588 (N_12588,N_12419,N_12443);
nand U12589 (N_12589,N_12428,N_12327);
and U12590 (N_12590,N_12445,N_12439);
and U12591 (N_12591,N_12442,N_12443);
xor U12592 (N_12592,N_12318,N_12380);
nor U12593 (N_12593,N_12418,N_12364);
nand U12594 (N_12594,N_12426,N_12407);
xor U12595 (N_12595,N_12438,N_12343);
or U12596 (N_12596,N_12385,N_12317);
xnor U12597 (N_12597,N_12394,N_12390);
and U12598 (N_12598,N_12369,N_12331);
or U12599 (N_12599,N_12370,N_12312);
nand U12600 (N_12600,N_12501,N_12517);
or U12601 (N_12601,N_12473,N_12585);
xnor U12602 (N_12602,N_12499,N_12561);
nand U12603 (N_12603,N_12476,N_12488);
xor U12604 (N_12604,N_12510,N_12482);
nand U12605 (N_12605,N_12454,N_12522);
or U12606 (N_12606,N_12569,N_12566);
xor U12607 (N_12607,N_12538,N_12554);
nor U12608 (N_12608,N_12458,N_12500);
xnor U12609 (N_12609,N_12514,N_12478);
xor U12610 (N_12610,N_12565,N_12583);
nand U12611 (N_12611,N_12556,N_12493);
and U12612 (N_12612,N_12559,N_12536);
nand U12613 (N_12613,N_12504,N_12481);
nand U12614 (N_12614,N_12576,N_12584);
and U12615 (N_12615,N_12581,N_12465);
xor U12616 (N_12616,N_12484,N_12487);
xor U12617 (N_12617,N_12579,N_12460);
or U12618 (N_12618,N_12523,N_12582);
nor U12619 (N_12619,N_12524,N_12477);
xnor U12620 (N_12620,N_12496,N_12527);
and U12621 (N_12621,N_12532,N_12558);
xor U12622 (N_12622,N_12570,N_12557);
nor U12623 (N_12623,N_12457,N_12474);
nor U12624 (N_12624,N_12545,N_12567);
xnor U12625 (N_12625,N_12498,N_12533);
or U12626 (N_12626,N_12525,N_12505);
nand U12627 (N_12627,N_12518,N_12492);
and U12628 (N_12628,N_12596,N_12589);
nand U12629 (N_12629,N_12489,N_12503);
nand U12630 (N_12630,N_12564,N_12571);
and U12631 (N_12631,N_12521,N_12469);
xnor U12632 (N_12632,N_12529,N_12586);
and U12633 (N_12633,N_12531,N_12450);
nor U12634 (N_12634,N_12575,N_12590);
and U12635 (N_12635,N_12459,N_12591);
nor U12636 (N_12636,N_12475,N_12549);
or U12637 (N_12637,N_12593,N_12592);
nor U12638 (N_12638,N_12555,N_12516);
xnor U12639 (N_12639,N_12451,N_12515);
or U12640 (N_12640,N_12599,N_12452);
or U12641 (N_12641,N_12463,N_12467);
and U12642 (N_12642,N_12468,N_12541);
or U12643 (N_12643,N_12461,N_12494);
and U12644 (N_12644,N_12466,N_12563);
nand U12645 (N_12645,N_12534,N_12480);
nor U12646 (N_12646,N_12572,N_12509);
and U12647 (N_12647,N_12588,N_12577);
nor U12648 (N_12648,N_12508,N_12464);
xor U12649 (N_12649,N_12456,N_12542);
or U12650 (N_12650,N_12544,N_12483);
and U12651 (N_12651,N_12540,N_12550);
nor U12652 (N_12652,N_12495,N_12519);
xor U12653 (N_12653,N_12486,N_12485);
nand U12654 (N_12654,N_12562,N_12455);
nor U12655 (N_12655,N_12462,N_12568);
nor U12656 (N_12656,N_12453,N_12546);
nor U12657 (N_12657,N_12553,N_12537);
nor U12658 (N_12658,N_12597,N_12490);
and U12659 (N_12659,N_12551,N_12502);
and U12660 (N_12660,N_12594,N_12470);
or U12661 (N_12661,N_12472,N_12595);
or U12662 (N_12662,N_12497,N_12539);
and U12663 (N_12663,N_12548,N_12530);
nor U12664 (N_12664,N_12578,N_12560);
nor U12665 (N_12665,N_12535,N_12513);
nor U12666 (N_12666,N_12511,N_12479);
xnor U12667 (N_12667,N_12598,N_12520);
nor U12668 (N_12668,N_12587,N_12491);
and U12669 (N_12669,N_12507,N_12573);
and U12670 (N_12670,N_12547,N_12506);
nand U12671 (N_12671,N_12526,N_12528);
nor U12672 (N_12672,N_12512,N_12552);
nor U12673 (N_12673,N_12543,N_12574);
nor U12674 (N_12674,N_12471,N_12580);
xor U12675 (N_12675,N_12599,N_12540);
and U12676 (N_12676,N_12583,N_12467);
or U12677 (N_12677,N_12578,N_12529);
or U12678 (N_12678,N_12555,N_12507);
nor U12679 (N_12679,N_12493,N_12547);
nand U12680 (N_12680,N_12562,N_12465);
or U12681 (N_12681,N_12513,N_12511);
xnor U12682 (N_12682,N_12588,N_12509);
nand U12683 (N_12683,N_12488,N_12543);
or U12684 (N_12684,N_12526,N_12454);
nor U12685 (N_12685,N_12583,N_12514);
xor U12686 (N_12686,N_12561,N_12551);
and U12687 (N_12687,N_12485,N_12567);
nor U12688 (N_12688,N_12576,N_12569);
nor U12689 (N_12689,N_12476,N_12503);
nand U12690 (N_12690,N_12484,N_12562);
nand U12691 (N_12691,N_12475,N_12454);
nor U12692 (N_12692,N_12570,N_12529);
xnor U12693 (N_12693,N_12550,N_12538);
or U12694 (N_12694,N_12499,N_12507);
nor U12695 (N_12695,N_12526,N_12505);
and U12696 (N_12696,N_12580,N_12479);
nand U12697 (N_12697,N_12563,N_12579);
xnor U12698 (N_12698,N_12537,N_12500);
nand U12699 (N_12699,N_12519,N_12590);
and U12700 (N_12700,N_12487,N_12455);
or U12701 (N_12701,N_12509,N_12539);
nor U12702 (N_12702,N_12583,N_12556);
or U12703 (N_12703,N_12516,N_12499);
nor U12704 (N_12704,N_12508,N_12546);
xor U12705 (N_12705,N_12559,N_12583);
and U12706 (N_12706,N_12552,N_12497);
and U12707 (N_12707,N_12469,N_12559);
xor U12708 (N_12708,N_12569,N_12504);
nand U12709 (N_12709,N_12568,N_12487);
or U12710 (N_12710,N_12494,N_12464);
xor U12711 (N_12711,N_12513,N_12451);
nor U12712 (N_12712,N_12554,N_12459);
nand U12713 (N_12713,N_12494,N_12475);
xnor U12714 (N_12714,N_12534,N_12498);
or U12715 (N_12715,N_12559,N_12460);
and U12716 (N_12716,N_12471,N_12584);
and U12717 (N_12717,N_12563,N_12519);
nand U12718 (N_12718,N_12595,N_12545);
and U12719 (N_12719,N_12516,N_12569);
or U12720 (N_12720,N_12583,N_12494);
and U12721 (N_12721,N_12528,N_12531);
nand U12722 (N_12722,N_12515,N_12547);
nor U12723 (N_12723,N_12513,N_12563);
and U12724 (N_12724,N_12454,N_12470);
and U12725 (N_12725,N_12460,N_12578);
nand U12726 (N_12726,N_12542,N_12590);
or U12727 (N_12727,N_12456,N_12524);
and U12728 (N_12728,N_12574,N_12538);
nand U12729 (N_12729,N_12574,N_12521);
or U12730 (N_12730,N_12539,N_12506);
or U12731 (N_12731,N_12558,N_12476);
or U12732 (N_12732,N_12580,N_12492);
or U12733 (N_12733,N_12538,N_12586);
and U12734 (N_12734,N_12581,N_12535);
or U12735 (N_12735,N_12513,N_12598);
or U12736 (N_12736,N_12499,N_12529);
nand U12737 (N_12737,N_12495,N_12587);
xor U12738 (N_12738,N_12588,N_12475);
xnor U12739 (N_12739,N_12499,N_12465);
and U12740 (N_12740,N_12471,N_12516);
xor U12741 (N_12741,N_12595,N_12511);
xor U12742 (N_12742,N_12471,N_12547);
xnor U12743 (N_12743,N_12487,N_12472);
nand U12744 (N_12744,N_12500,N_12552);
xor U12745 (N_12745,N_12595,N_12577);
nor U12746 (N_12746,N_12518,N_12587);
nor U12747 (N_12747,N_12458,N_12583);
and U12748 (N_12748,N_12566,N_12565);
and U12749 (N_12749,N_12532,N_12591);
and U12750 (N_12750,N_12673,N_12706);
and U12751 (N_12751,N_12738,N_12740);
xnor U12752 (N_12752,N_12705,N_12626);
nand U12753 (N_12753,N_12663,N_12745);
and U12754 (N_12754,N_12698,N_12631);
nor U12755 (N_12755,N_12610,N_12700);
and U12756 (N_12756,N_12617,N_12612);
xnor U12757 (N_12757,N_12647,N_12624);
and U12758 (N_12758,N_12627,N_12741);
and U12759 (N_12759,N_12608,N_12620);
nand U12760 (N_12760,N_12713,N_12629);
and U12761 (N_12761,N_12748,N_12644);
or U12762 (N_12762,N_12732,N_12600);
or U12763 (N_12763,N_12659,N_12699);
or U12764 (N_12764,N_12642,N_12630);
or U12765 (N_12765,N_12684,N_12743);
nand U12766 (N_12766,N_12625,N_12669);
nor U12767 (N_12767,N_12671,N_12731);
nor U12768 (N_12768,N_12662,N_12670);
nor U12769 (N_12769,N_12653,N_12747);
nand U12770 (N_12770,N_12672,N_12697);
xor U12771 (N_12771,N_12666,N_12694);
nand U12772 (N_12772,N_12723,N_12667);
or U12773 (N_12773,N_12695,N_12712);
xnor U12774 (N_12774,N_12635,N_12616);
and U12775 (N_12775,N_12657,N_12707);
nor U12776 (N_12776,N_12729,N_12602);
xor U12777 (N_12777,N_12744,N_12674);
nor U12778 (N_12778,N_12676,N_12702);
xnor U12779 (N_12779,N_12643,N_12640);
and U12780 (N_12780,N_12716,N_12689);
nor U12781 (N_12781,N_12655,N_12749);
or U12782 (N_12782,N_12677,N_12680);
and U12783 (N_12783,N_12734,N_12633);
xnor U12784 (N_12784,N_12742,N_12604);
and U12785 (N_12785,N_12726,N_12687);
or U12786 (N_12786,N_12603,N_12660);
nor U12787 (N_12787,N_12727,N_12609);
and U12788 (N_12788,N_12658,N_12639);
nor U12789 (N_12789,N_12668,N_12691);
and U12790 (N_12790,N_12715,N_12721);
xor U12791 (N_12791,N_12621,N_12696);
or U12792 (N_12792,N_12637,N_12645);
or U12793 (N_12793,N_12692,N_12638);
or U12794 (N_12794,N_12704,N_12628);
or U12795 (N_12795,N_12720,N_12652);
nand U12796 (N_12796,N_12736,N_12724);
nor U12797 (N_12797,N_12675,N_12618);
nor U12798 (N_12798,N_12606,N_12685);
or U12799 (N_12799,N_12656,N_12661);
xnor U12800 (N_12800,N_12681,N_12701);
and U12801 (N_12801,N_12722,N_12665);
nand U12802 (N_12802,N_12739,N_12623);
and U12803 (N_12803,N_12651,N_12619);
nand U12804 (N_12804,N_12654,N_12708);
or U12805 (N_12805,N_12714,N_12634);
or U12806 (N_12806,N_12730,N_12613);
or U12807 (N_12807,N_12688,N_12601);
or U12808 (N_12808,N_12641,N_12615);
and U12809 (N_12809,N_12683,N_12711);
xor U12810 (N_12810,N_12632,N_12717);
xnor U12811 (N_12811,N_12686,N_12605);
and U12812 (N_12812,N_12622,N_12728);
nand U12813 (N_12813,N_12646,N_12725);
nor U12814 (N_12814,N_12710,N_12614);
and U12815 (N_12815,N_12678,N_12733);
or U12816 (N_12816,N_12648,N_12611);
xor U12817 (N_12817,N_12703,N_12679);
nand U12818 (N_12818,N_12690,N_12636);
nand U12819 (N_12819,N_12650,N_12607);
or U12820 (N_12820,N_12746,N_12719);
and U12821 (N_12821,N_12718,N_12737);
or U12822 (N_12822,N_12693,N_12709);
nand U12823 (N_12823,N_12664,N_12649);
nand U12824 (N_12824,N_12682,N_12735);
or U12825 (N_12825,N_12670,N_12686);
nand U12826 (N_12826,N_12639,N_12609);
nand U12827 (N_12827,N_12623,N_12686);
and U12828 (N_12828,N_12723,N_12668);
xnor U12829 (N_12829,N_12653,N_12738);
nor U12830 (N_12830,N_12719,N_12622);
xnor U12831 (N_12831,N_12645,N_12675);
xor U12832 (N_12832,N_12602,N_12605);
or U12833 (N_12833,N_12639,N_12608);
xor U12834 (N_12834,N_12611,N_12607);
nand U12835 (N_12835,N_12712,N_12679);
xor U12836 (N_12836,N_12649,N_12679);
nor U12837 (N_12837,N_12635,N_12662);
nor U12838 (N_12838,N_12654,N_12689);
nand U12839 (N_12839,N_12740,N_12606);
or U12840 (N_12840,N_12740,N_12663);
nor U12841 (N_12841,N_12705,N_12651);
and U12842 (N_12842,N_12613,N_12741);
nor U12843 (N_12843,N_12713,N_12648);
xnor U12844 (N_12844,N_12685,N_12705);
nor U12845 (N_12845,N_12694,N_12688);
xor U12846 (N_12846,N_12746,N_12643);
xnor U12847 (N_12847,N_12601,N_12605);
nand U12848 (N_12848,N_12705,N_12637);
nor U12849 (N_12849,N_12646,N_12735);
nor U12850 (N_12850,N_12619,N_12602);
or U12851 (N_12851,N_12748,N_12685);
and U12852 (N_12852,N_12690,N_12695);
xnor U12853 (N_12853,N_12679,N_12718);
nand U12854 (N_12854,N_12694,N_12629);
nand U12855 (N_12855,N_12690,N_12628);
and U12856 (N_12856,N_12680,N_12651);
or U12857 (N_12857,N_12657,N_12618);
xnor U12858 (N_12858,N_12749,N_12628);
nand U12859 (N_12859,N_12716,N_12744);
and U12860 (N_12860,N_12697,N_12692);
xor U12861 (N_12861,N_12709,N_12673);
or U12862 (N_12862,N_12693,N_12670);
or U12863 (N_12863,N_12649,N_12728);
or U12864 (N_12864,N_12738,N_12707);
nor U12865 (N_12865,N_12735,N_12611);
and U12866 (N_12866,N_12747,N_12733);
and U12867 (N_12867,N_12648,N_12666);
or U12868 (N_12868,N_12634,N_12603);
nor U12869 (N_12869,N_12704,N_12692);
or U12870 (N_12870,N_12721,N_12651);
nor U12871 (N_12871,N_12616,N_12651);
or U12872 (N_12872,N_12631,N_12628);
or U12873 (N_12873,N_12643,N_12625);
or U12874 (N_12874,N_12661,N_12718);
and U12875 (N_12875,N_12732,N_12711);
and U12876 (N_12876,N_12624,N_12606);
nand U12877 (N_12877,N_12624,N_12617);
nor U12878 (N_12878,N_12647,N_12638);
nand U12879 (N_12879,N_12657,N_12667);
nor U12880 (N_12880,N_12612,N_12642);
or U12881 (N_12881,N_12736,N_12692);
xnor U12882 (N_12882,N_12656,N_12621);
nor U12883 (N_12883,N_12660,N_12655);
nand U12884 (N_12884,N_12650,N_12710);
or U12885 (N_12885,N_12617,N_12727);
nand U12886 (N_12886,N_12632,N_12747);
nand U12887 (N_12887,N_12716,N_12608);
and U12888 (N_12888,N_12640,N_12746);
or U12889 (N_12889,N_12625,N_12675);
and U12890 (N_12890,N_12682,N_12646);
xor U12891 (N_12891,N_12744,N_12664);
nand U12892 (N_12892,N_12729,N_12692);
xor U12893 (N_12893,N_12711,N_12637);
nand U12894 (N_12894,N_12744,N_12654);
and U12895 (N_12895,N_12623,N_12720);
nand U12896 (N_12896,N_12718,N_12638);
nor U12897 (N_12897,N_12748,N_12681);
and U12898 (N_12898,N_12676,N_12717);
nand U12899 (N_12899,N_12632,N_12707);
nand U12900 (N_12900,N_12827,N_12849);
and U12901 (N_12901,N_12810,N_12868);
nand U12902 (N_12902,N_12751,N_12760);
xor U12903 (N_12903,N_12767,N_12845);
xor U12904 (N_12904,N_12848,N_12863);
nand U12905 (N_12905,N_12778,N_12887);
nand U12906 (N_12906,N_12784,N_12765);
xor U12907 (N_12907,N_12779,N_12753);
xnor U12908 (N_12908,N_12890,N_12832);
or U12909 (N_12909,N_12752,N_12831);
nand U12910 (N_12910,N_12830,N_12835);
nor U12911 (N_12911,N_12799,N_12841);
or U12912 (N_12912,N_12815,N_12822);
nor U12913 (N_12913,N_12823,N_12802);
or U12914 (N_12914,N_12793,N_12854);
xor U12915 (N_12915,N_12794,N_12857);
or U12916 (N_12916,N_12861,N_12895);
xor U12917 (N_12917,N_12804,N_12801);
xnor U12918 (N_12918,N_12782,N_12812);
nand U12919 (N_12919,N_12783,N_12791);
nor U12920 (N_12920,N_12888,N_12786);
or U12921 (N_12921,N_12780,N_12893);
and U12922 (N_12922,N_12851,N_12787);
or U12923 (N_12923,N_12843,N_12803);
or U12924 (N_12924,N_12766,N_12870);
nand U12925 (N_12925,N_12864,N_12816);
xor U12926 (N_12926,N_12761,N_12800);
nor U12927 (N_12927,N_12859,N_12825);
or U12928 (N_12928,N_12880,N_12875);
xnor U12929 (N_12929,N_12789,N_12770);
or U12930 (N_12930,N_12807,N_12750);
nor U12931 (N_12931,N_12762,N_12818);
and U12932 (N_12932,N_12883,N_12808);
nor U12933 (N_12933,N_12775,N_12867);
nor U12934 (N_12934,N_12834,N_12814);
nand U12935 (N_12935,N_12858,N_12809);
nor U12936 (N_12936,N_12840,N_12886);
nand U12937 (N_12937,N_12754,N_12855);
nand U12938 (N_12938,N_12769,N_12837);
nor U12939 (N_12939,N_12836,N_12891);
xnor U12940 (N_12940,N_12838,N_12853);
and U12941 (N_12941,N_12811,N_12869);
xor U12942 (N_12942,N_12758,N_12862);
and U12943 (N_12943,N_12860,N_12873);
and U12944 (N_12944,N_12877,N_12764);
nor U12945 (N_12945,N_12897,N_12846);
or U12946 (N_12946,N_12852,N_12768);
xnor U12947 (N_12947,N_12756,N_12833);
nor U12948 (N_12948,N_12774,N_12805);
nand U12949 (N_12949,N_12874,N_12757);
or U12950 (N_12950,N_12885,N_12844);
and U12951 (N_12951,N_12790,N_12892);
xor U12952 (N_12952,N_12881,N_12829);
or U12953 (N_12953,N_12824,N_12828);
nand U12954 (N_12954,N_12788,N_12896);
nor U12955 (N_12955,N_12781,N_12776);
nand U12956 (N_12956,N_12797,N_12894);
and U12957 (N_12957,N_12889,N_12777);
xor U12958 (N_12958,N_12878,N_12847);
or U12959 (N_12959,N_12821,N_12872);
nand U12960 (N_12960,N_12856,N_12806);
or U12961 (N_12961,N_12785,N_12839);
nor U12962 (N_12962,N_12795,N_12796);
or U12963 (N_12963,N_12865,N_12813);
xor U12964 (N_12964,N_12866,N_12759);
or U12965 (N_12965,N_12842,N_12773);
nor U12966 (N_12966,N_12819,N_12879);
nor U12967 (N_12967,N_12850,N_12899);
or U12968 (N_12968,N_12763,N_12755);
xor U12969 (N_12969,N_12798,N_12820);
nand U12970 (N_12970,N_12876,N_12871);
or U12971 (N_12971,N_12898,N_12817);
or U12972 (N_12972,N_12771,N_12772);
and U12973 (N_12973,N_12882,N_12884);
and U12974 (N_12974,N_12826,N_12792);
nand U12975 (N_12975,N_12829,N_12811);
nand U12976 (N_12976,N_12809,N_12814);
and U12977 (N_12977,N_12821,N_12849);
xor U12978 (N_12978,N_12815,N_12840);
nand U12979 (N_12979,N_12865,N_12832);
and U12980 (N_12980,N_12860,N_12859);
and U12981 (N_12981,N_12893,N_12880);
nand U12982 (N_12982,N_12808,N_12788);
xor U12983 (N_12983,N_12837,N_12774);
nor U12984 (N_12984,N_12841,N_12769);
or U12985 (N_12985,N_12890,N_12881);
nand U12986 (N_12986,N_12838,N_12841);
nor U12987 (N_12987,N_12795,N_12846);
or U12988 (N_12988,N_12883,N_12875);
xnor U12989 (N_12989,N_12772,N_12816);
and U12990 (N_12990,N_12825,N_12805);
or U12991 (N_12991,N_12766,N_12830);
and U12992 (N_12992,N_12867,N_12830);
nor U12993 (N_12993,N_12878,N_12766);
and U12994 (N_12994,N_12865,N_12896);
xnor U12995 (N_12995,N_12791,N_12882);
nand U12996 (N_12996,N_12870,N_12791);
or U12997 (N_12997,N_12851,N_12793);
xnor U12998 (N_12998,N_12773,N_12859);
nand U12999 (N_12999,N_12773,N_12763);
or U13000 (N_13000,N_12762,N_12855);
and U13001 (N_13001,N_12756,N_12866);
nand U13002 (N_13002,N_12755,N_12866);
nand U13003 (N_13003,N_12755,N_12830);
or U13004 (N_13004,N_12785,N_12770);
and U13005 (N_13005,N_12872,N_12848);
nor U13006 (N_13006,N_12889,N_12771);
xor U13007 (N_13007,N_12840,N_12827);
nor U13008 (N_13008,N_12785,N_12891);
and U13009 (N_13009,N_12883,N_12889);
or U13010 (N_13010,N_12785,N_12871);
nand U13011 (N_13011,N_12885,N_12787);
xor U13012 (N_13012,N_12822,N_12777);
and U13013 (N_13013,N_12829,N_12890);
nor U13014 (N_13014,N_12756,N_12864);
or U13015 (N_13015,N_12783,N_12771);
nand U13016 (N_13016,N_12859,N_12769);
and U13017 (N_13017,N_12787,N_12757);
xor U13018 (N_13018,N_12844,N_12889);
nor U13019 (N_13019,N_12881,N_12758);
or U13020 (N_13020,N_12851,N_12861);
xnor U13021 (N_13021,N_12787,N_12794);
nand U13022 (N_13022,N_12877,N_12782);
nand U13023 (N_13023,N_12808,N_12774);
xnor U13024 (N_13024,N_12799,N_12884);
nor U13025 (N_13025,N_12896,N_12801);
or U13026 (N_13026,N_12818,N_12896);
xor U13027 (N_13027,N_12882,N_12763);
xnor U13028 (N_13028,N_12867,N_12750);
and U13029 (N_13029,N_12753,N_12865);
nor U13030 (N_13030,N_12807,N_12894);
or U13031 (N_13031,N_12831,N_12866);
nand U13032 (N_13032,N_12841,N_12820);
or U13033 (N_13033,N_12813,N_12882);
nor U13034 (N_13034,N_12851,N_12829);
nand U13035 (N_13035,N_12874,N_12837);
nand U13036 (N_13036,N_12794,N_12771);
and U13037 (N_13037,N_12872,N_12781);
nor U13038 (N_13038,N_12810,N_12849);
or U13039 (N_13039,N_12895,N_12770);
and U13040 (N_13040,N_12894,N_12808);
nand U13041 (N_13041,N_12762,N_12768);
nor U13042 (N_13042,N_12802,N_12856);
nor U13043 (N_13043,N_12833,N_12868);
or U13044 (N_13044,N_12840,N_12813);
nor U13045 (N_13045,N_12811,N_12825);
and U13046 (N_13046,N_12767,N_12876);
nor U13047 (N_13047,N_12874,N_12879);
nor U13048 (N_13048,N_12758,N_12885);
nor U13049 (N_13049,N_12884,N_12851);
or U13050 (N_13050,N_12910,N_13000);
and U13051 (N_13051,N_13018,N_13024);
nand U13052 (N_13052,N_13012,N_12947);
xnor U13053 (N_13053,N_12914,N_13048);
and U13054 (N_13054,N_13037,N_12976);
xor U13055 (N_13055,N_13004,N_13027);
xor U13056 (N_13056,N_12937,N_12955);
nand U13057 (N_13057,N_13044,N_12906);
nand U13058 (N_13058,N_12965,N_12926);
nand U13059 (N_13059,N_12983,N_12970);
and U13060 (N_13060,N_12908,N_13042);
nand U13061 (N_13061,N_12980,N_13015);
and U13062 (N_13062,N_12988,N_12928);
and U13063 (N_13063,N_12918,N_12944);
and U13064 (N_13064,N_13029,N_12956);
xnor U13065 (N_13065,N_12999,N_12938);
or U13066 (N_13066,N_12951,N_12979);
nor U13067 (N_13067,N_13014,N_13028);
xor U13068 (N_13068,N_12936,N_12907);
xor U13069 (N_13069,N_12911,N_12978);
nor U13070 (N_13070,N_13036,N_13045);
nor U13071 (N_13071,N_12982,N_12996);
xor U13072 (N_13072,N_12927,N_12957);
and U13073 (N_13073,N_12919,N_12950);
and U13074 (N_13074,N_13047,N_12923);
nand U13075 (N_13075,N_13034,N_12990);
nand U13076 (N_13076,N_12973,N_13041);
or U13077 (N_13077,N_12925,N_12963);
nand U13078 (N_13078,N_12933,N_12959);
nand U13079 (N_13079,N_12989,N_12909);
or U13080 (N_13080,N_12968,N_12945);
xor U13081 (N_13081,N_13022,N_12939);
nand U13082 (N_13082,N_12913,N_12969);
nor U13083 (N_13083,N_12952,N_13021);
xnor U13084 (N_13084,N_12958,N_12940);
nor U13085 (N_13085,N_12992,N_12949);
nand U13086 (N_13086,N_12917,N_13011);
nand U13087 (N_13087,N_13040,N_12901);
nor U13088 (N_13088,N_13001,N_12929);
nor U13089 (N_13089,N_12942,N_12900);
nor U13090 (N_13090,N_12986,N_12946);
nor U13091 (N_13091,N_12998,N_12977);
xor U13092 (N_13092,N_12995,N_12922);
or U13093 (N_13093,N_12994,N_12924);
or U13094 (N_13094,N_13046,N_12904);
nor U13095 (N_13095,N_12915,N_13033);
nand U13096 (N_13096,N_13016,N_13035);
or U13097 (N_13097,N_12974,N_12997);
nand U13098 (N_13098,N_13002,N_12905);
and U13099 (N_13099,N_12941,N_13013);
xor U13100 (N_13100,N_13030,N_12967);
nand U13101 (N_13101,N_12934,N_13038);
and U13102 (N_13102,N_13005,N_13020);
or U13103 (N_13103,N_12931,N_12962);
and U13104 (N_13104,N_12984,N_12964);
and U13105 (N_13105,N_12960,N_12943);
or U13106 (N_13106,N_12975,N_12961);
nand U13107 (N_13107,N_13006,N_13049);
and U13108 (N_13108,N_12987,N_12903);
and U13109 (N_13109,N_12930,N_13003);
or U13110 (N_13110,N_12932,N_12971);
and U13111 (N_13111,N_13023,N_13043);
nand U13112 (N_13112,N_12954,N_12985);
nand U13113 (N_13113,N_12991,N_13025);
and U13114 (N_13114,N_12993,N_12920);
nand U13115 (N_13115,N_12912,N_13032);
nor U13116 (N_13116,N_12935,N_12916);
and U13117 (N_13117,N_13010,N_13019);
nand U13118 (N_13118,N_13039,N_13017);
xor U13119 (N_13119,N_12921,N_13026);
xnor U13120 (N_13120,N_12981,N_13008);
or U13121 (N_13121,N_13031,N_12972);
nor U13122 (N_13122,N_12902,N_12948);
nor U13123 (N_13123,N_13007,N_13009);
xnor U13124 (N_13124,N_12953,N_12966);
nand U13125 (N_13125,N_13023,N_12999);
xnor U13126 (N_13126,N_12913,N_13020);
and U13127 (N_13127,N_12956,N_12937);
and U13128 (N_13128,N_12916,N_12963);
nor U13129 (N_13129,N_12902,N_12970);
xnor U13130 (N_13130,N_13012,N_12943);
nor U13131 (N_13131,N_12913,N_12906);
nor U13132 (N_13132,N_13018,N_13001);
xor U13133 (N_13133,N_12914,N_13035);
xor U13134 (N_13134,N_12947,N_13025);
nor U13135 (N_13135,N_12940,N_13004);
and U13136 (N_13136,N_13022,N_12948);
or U13137 (N_13137,N_12933,N_12921);
nand U13138 (N_13138,N_12906,N_12974);
nor U13139 (N_13139,N_12984,N_12919);
nand U13140 (N_13140,N_12966,N_12936);
or U13141 (N_13141,N_13032,N_13016);
nand U13142 (N_13142,N_12955,N_13028);
xnor U13143 (N_13143,N_12987,N_13048);
xor U13144 (N_13144,N_13033,N_12955);
or U13145 (N_13145,N_12957,N_12991);
and U13146 (N_13146,N_12953,N_12973);
xor U13147 (N_13147,N_12989,N_12999);
nand U13148 (N_13148,N_12901,N_12921);
nor U13149 (N_13149,N_12916,N_12949);
nand U13150 (N_13150,N_13019,N_12989);
nor U13151 (N_13151,N_13044,N_12978);
xnor U13152 (N_13152,N_12942,N_12997);
nor U13153 (N_13153,N_12939,N_13013);
xor U13154 (N_13154,N_12938,N_13030);
xnor U13155 (N_13155,N_12914,N_13005);
and U13156 (N_13156,N_13033,N_13002);
xnor U13157 (N_13157,N_12977,N_12999);
nor U13158 (N_13158,N_12901,N_12925);
xor U13159 (N_13159,N_13037,N_13007);
nor U13160 (N_13160,N_12984,N_12942);
xor U13161 (N_13161,N_12944,N_13024);
xor U13162 (N_13162,N_13041,N_13014);
nor U13163 (N_13163,N_12984,N_12936);
or U13164 (N_13164,N_13029,N_12982);
nor U13165 (N_13165,N_12931,N_12963);
or U13166 (N_13166,N_12913,N_12954);
and U13167 (N_13167,N_13000,N_12909);
nor U13168 (N_13168,N_13048,N_12957);
and U13169 (N_13169,N_13047,N_13049);
nor U13170 (N_13170,N_13025,N_12934);
nand U13171 (N_13171,N_13010,N_12998);
nand U13172 (N_13172,N_12931,N_12973);
or U13173 (N_13173,N_13028,N_13046);
and U13174 (N_13174,N_12920,N_12949);
nand U13175 (N_13175,N_12989,N_13026);
or U13176 (N_13176,N_12936,N_13019);
nor U13177 (N_13177,N_13016,N_12946);
or U13178 (N_13178,N_12966,N_13045);
xnor U13179 (N_13179,N_12989,N_12962);
and U13180 (N_13180,N_12985,N_12910);
or U13181 (N_13181,N_12963,N_13037);
xor U13182 (N_13182,N_13046,N_12926);
nand U13183 (N_13183,N_12970,N_12980);
nor U13184 (N_13184,N_13013,N_13029);
and U13185 (N_13185,N_13020,N_12962);
nor U13186 (N_13186,N_13048,N_12943);
nor U13187 (N_13187,N_12921,N_12910);
xor U13188 (N_13188,N_13037,N_13048);
or U13189 (N_13189,N_12939,N_12909);
or U13190 (N_13190,N_12993,N_13030);
or U13191 (N_13191,N_13030,N_13016);
nand U13192 (N_13192,N_12938,N_13021);
and U13193 (N_13193,N_12917,N_12985);
nand U13194 (N_13194,N_13023,N_12929);
or U13195 (N_13195,N_12947,N_13028);
or U13196 (N_13196,N_12954,N_12919);
xor U13197 (N_13197,N_12921,N_12935);
nand U13198 (N_13198,N_13004,N_12926);
nor U13199 (N_13199,N_12906,N_13006);
and U13200 (N_13200,N_13173,N_13181);
nand U13201 (N_13201,N_13146,N_13088);
xnor U13202 (N_13202,N_13135,N_13105);
and U13203 (N_13203,N_13157,N_13171);
nand U13204 (N_13204,N_13094,N_13182);
nor U13205 (N_13205,N_13198,N_13128);
or U13206 (N_13206,N_13185,N_13114);
nand U13207 (N_13207,N_13111,N_13194);
or U13208 (N_13208,N_13090,N_13070);
or U13209 (N_13209,N_13193,N_13163);
and U13210 (N_13210,N_13058,N_13110);
or U13211 (N_13211,N_13151,N_13116);
and U13212 (N_13212,N_13099,N_13167);
nor U13213 (N_13213,N_13176,N_13124);
xor U13214 (N_13214,N_13068,N_13100);
or U13215 (N_13215,N_13140,N_13168);
xor U13216 (N_13216,N_13106,N_13084);
and U13217 (N_13217,N_13131,N_13109);
nor U13218 (N_13218,N_13187,N_13149);
nand U13219 (N_13219,N_13190,N_13152);
nand U13220 (N_13220,N_13175,N_13098);
xnor U13221 (N_13221,N_13166,N_13091);
and U13222 (N_13222,N_13067,N_13199);
and U13223 (N_13223,N_13071,N_13092);
nand U13224 (N_13224,N_13062,N_13112);
or U13225 (N_13225,N_13178,N_13072);
nand U13226 (N_13226,N_13069,N_13192);
or U13227 (N_13227,N_13055,N_13136);
nor U13228 (N_13228,N_13159,N_13082);
nand U13229 (N_13229,N_13086,N_13189);
and U13230 (N_13230,N_13059,N_13188);
xor U13231 (N_13231,N_13161,N_13119);
and U13232 (N_13232,N_13080,N_13093);
xor U13233 (N_13233,N_13153,N_13150);
nand U13234 (N_13234,N_13061,N_13134);
and U13235 (N_13235,N_13078,N_13197);
or U13236 (N_13236,N_13170,N_13083);
or U13237 (N_13237,N_13180,N_13147);
or U13238 (N_13238,N_13121,N_13052);
and U13239 (N_13239,N_13117,N_13191);
nor U13240 (N_13240,N_13133,N_13075);
or U13241 (N_13241,N_13057,N_13169);
and U13242 (N_13242,N_13063,N_13139);
nor U13243 (N_13243,N_13183,N_13115);
and U13244 (N_13244,N_13126,N_13060);
or U13245 (N_13245,N_13148,N_13195);
or U13246 (N_13246,N_13054,N_13053);
and U13247 (N_13247,N_13144,N_13127);
xnor U13248 (N_13248,N_13165,N_13184);
xnor U13249 (N_13249,N_13196,N_13142);
and U13250 (N_13250,N_13079,N_13143);
nor U13251 (N_13251,N_13095,N_13097);
nor U13252 (N_13252,N_13051,N_13123);
and U13253 (N_13253,N_13122,N_13066);
or U13254 (N_13254,N_13172,N_13096);
nor U13255 (N_13255,N_13174,N_13141);
or U13256 (N_13256,N_13103,N_13156);
nand U13257 (N_13257,N_13056,N_13104);
or U13258 (N_13258,N_13107,N_13138);
nand U13259 (N_13259,N_13137,N_13155);
and U13260 (N_13260,N_13125,N_13085);
or U13261 (N_13261,N_13087,N_13064);
and U13262 (N_13262,N_13081,N_13118);
or U13263 (N_13263,N_13154,N_13076);
or U13264 (N_13264,N_13089,N_13179);
and U13265 (N_13265,N_13162,N_13077);
or U13266 (N_13266,N_13108,N_13130);
xnor U13267 (N_13267,N_13101,N_13160);
nor U13268 (N_13268,N_13129,N_13113);
nand U13269 (N_13269,N_13102,N_13132);
xnor U13270 (N_13270,N_13050,N_13120);
nand U13271 (N_13271,N_13073,N_13186);
xnor U13272 (N_13272,N_13074,N_13164);
xnor U13273 (N_13273,N_13065,N_13145);
nor U13274 (N_13274,N_13158,N_13177);
nor U13275 (N_13275,N_13137,N_13090);
xor U13276 (N_13276,N_13079,N_13064);
xnor U13277 (N_13277,N_13132,N_13178);
and U13278 (N_13278,N_13143,N_13070);
and U13279 (N_13279,N_13139,N_13099);
nor U13280 (N_13280,N_13135,N_13066);
or U13281 (N_13281,N_13121,N_13123);
xnor U13282 (N_13282,N_13171,N_13059);
nor U13283 (N_13283,N_13150,N_13090);
nor U13284 (N_13284,N_13096,N_13146);
xnor U13285 (N_13285,N_13178,N_13051);
or U13286 (N_13286,N_13146,N_13050);
nand U13287 (N_13287,N_13147,N_13171);
xor U13288 (N_13288,N_13160,N_13093);
xor U13289 (N_13289,N_13064,N_13186);
nor U13290 (N_13290,N_13111,N_13138);
and U13291 (N_13291,N_13110,N_13093);
xor U13292 (N_13292,N_13198,N_13124);
or U13293 (N_13293,N_13137,N_13140);
nor U13294 (N_13294,N_13061,N_13193);
or U13295 (N_13295,N_13179,N_13057);
nor U13296 (N_13296,N_13165,N_13189);
or U13297 (N_13297,N_13090,N_13179);
or U13298 (N_13298,N_13076,N_13056);
xnor U13299 (N_13299,N_13156,N_13198);
nand U13300 (N_13300,N_13101,N_13184);
and U13301 (N_13301,N_13186,N_13156);
and U13302 (N_13302,N_13199,N_13135);
nor U13303 (N_13303,N_13141,N_13053);
and U13304 (N_13304,N_13080,N_13129);
nand U13305 (N_13305,N_13154,N_13089);
xnor U13306 (N_13306,N_13114,N_13159);
and U13307 (N_13307,N_13141,N_13080);
nand U13308 (N_13308,N_13087,N_13111);
xnor U13309 (N_13309,N_13135,N_13188);
xor U13310 (N_13310,N_13159,N_13149);
xnor U13311 (N_13311,N_13178,N_13152);
and U13312 (N_13312,N_13199,N_13102);
nor U13313 (N_13313,N_13067,N_13084);
or U13314 (N_13314,N_13132,N_13075);
nor U13315 (N_13315,N_13096,N_13163);
and U13316 (N_13316,N_13109,N_13118);
xnor U13317 (N_13317,N_13127,N_13186);
nor U13318 (N_13318,N_13053,N_13166);
nor U13319 (N_13319,N_13154,N_13186);
and U13320 (N_13320,N_13111,N_13092);
or U13321 (N_13321,N_13188,N_13061);
nand U13322 (N_13322,N_13198,N_13168);
or U13323 (N_13323,N_13106,N_13126);
or U13324 (N_13324,N_13083,N_13177);
nand U13325 (N_13325,N_13179,N_13131);
nor U13326 (N_13326,N_13186,N_13175);
nor U13327 (N_13327,N_13071,N_13097);
nand U13328 (N_13328,N_13149,N_13095);
nand U13329 (N_13329,N_13112,N_13130);
or U13330 (N_13330,N_13111,N_13085);
and U13331 (N_13331,N_13119,N_13110);
or U13332 (N_13332,N_13114,N_13157);
nand U13333 (N_13333,N_13161,N_13166);
nor U13334 (N_13334,N_13157,N_13146);
nand U13335 (N_13335,N_13152,N_13066);
nand U13336 (N_13336,N_13189,N_13143);
nor U13337 (N_13337,N_13101,N_13052);
nor U13338 (N_13338,N_13110,N_13072);
nor U13339 (N_13339,N_13181,N_13196);
xor U13340 (N_13340,N_13090,N_13076);
xnor U13341 (N_13341,N_13194,N_13132);
nand U13342 (N_13342,N_13081,N_13186);
xor U13343 (N_13343,N_13192,N_13143);
nand U13344 (N_13344,N_13150,N_13175);
nand U13345 (N_13345,N_13144,N_13095);
xnor U13346 (N_13346,N_13052,N_13057);
nor U13347 (N_13347,N_13160,N_13094);
xor U13348 (N_13348,N_13069,N_13135);
or U13349 (N_13349,N_13178,N_13199);
xnor U13350 (N_13350,N_13228,N_13329);
xor U13351 (N_13351,N_13263,N_13281);
or U13352 (N_13352,N_13303,N_13200);
and U13353 (N_13353,N_13206,N_13262);
nand U13354 (N_13354,N_13276,N_13256);
nand U13355 (N_13355,N_13333,N_13264);
and U13356 (N_13356,N_13250,N_13280);
xnor U13357 (N_13357,N_13305,N_13313);
nor U13358 (N_13358,N_13239,N_13201);
nor U13359 (N_13359,N_13267,N_13340);
and U13360 (N_13360,N_13240,N_13279);
nand U13361 (N_13361,N_13237,N_13326);
nand U13362 (N_13362,N_13271,N_13300);
and U13363 (N_13363,N_13310,N_13323);
or U13364 (N_13364,N_13234,N_13316);
and U13365 (N_13365,N_13223,N_13222);
nand U13366 (N_13366,N_13244,N_13347);
nand U13367 (N_13367,N_13324,N_13221);
nand U13368 (N_13368,N_13336,N_13252);
nor U13369 (N_13369,N_13295,N_13242);
or U13370 (N_13370,N_13290,N_13211);
and U13371 (N_13371,N_13273,N_13284);
or U13372 (N_13372,N_13259,N_13288);
nor U13373 (N_13373,N_13301,N_13229);
or U13374 (N_13374,N_13246,N_13226);
xnor U13375 (N_13375,N_13224,N_13249);
or U13376 (N_13376,N_13275,N_13298);
xnor U13377 (N_13377,N_13322,N_13328);
nor U13378 (N_13378,N_13317,N_13248);
or U13379 (N_13379,N_13230,N_13245);
and U13380 (N_13380,N_13217,N_13208);
nand U13381 (N_13381,N_13210,N_13269);
nor U13382 (N_13382,N_13287,N_13241);
nor U13383 (N_13383,N_13346,N_13325);
xnor U13384 (N_13384,N_13297,N_13342);
or U13385 (N_13385,N_13247,N_13257);
nor U13386 (N_13386,N_13205,N_13341);
xor U13387 (N_13387,N_13207,N_13219);
or U13388 (N_13388,N_13233,N_13349);
and U13389 (N_13389,N_13312,N_13282);
or U13390 (N_13390,N_13214,N_13302);
or U13391 (N_13391,N_13338,N_13320);
or U13392 (N_13392,N_13265,N_13260);
xnor U13393 (N_13393,N_13339,N_13261);
nor U13394 (N_13394,N_13231,N_13327);
and U13395 (N_13395,N_13243,N_13292);
nor U13396 (N_13396,N_13232,N_13348);
or U13397 (N_13397,N_13345,N_13319);
and U13398 (N_13398,N_13318,N_13212);
nand U13399 (N_13399,N_13291,N_13274);
and U13400 (N_13400,N_13215,N_13321);
or U13401 (N_13401,N_13253,N_13343);
and U13402 (N_13402,N_13289,N_13307);
or U13403 (N_13403,N_13220,N_13334);
xnor U13404 (N_13404,N_13225,N_13283);
and U13405 (N_13405,N_13227,N_13308);
nor U13406 (N_13406,N_13286,N_13335);
nand U13407 (N_13407,N_13331,N_13218);
and U13408 (N_13408,N_13266,N_13255);
or U13409 (N_13409,N_13311,N_13213);
or U13410 (N_13410,N_13306,N_13203);
xnor U13411 (N_13411,N_13332,N_13268);
nor U13412 (N_13412,N_13258,N_13202);
or U13413 (N_13413,N_13236,N_13294);
or U13414 (N_13414,N_13330,N_13277);
or U13415 (N_13415,N_13272,N_13209);
or U13416 (N_13416,N_13270,N_13204);
nand U13417 (N_13417,N_13235,N_13216);
nor U13418 (N_13418,N_13251,N_13309);
or U13419 (N_13419,N_13285,N_13344);
xnor U13420 (N_13420,N_13254,N_13238);
nand U13421 (N_13421,N_13337,N_13296);
nand U13422 (N_13422,N_13315,N_13278);
xor U13423 (N_13423,N_13299,N_13293);
nor U13424 (N_13424,N_13304,N_13314);
xor U13425 (N_13425,N_13263,N_13286);
or U13426 (N_13426,N_13236,N_13291);
xnor U13427 (N_13427,N_13219,N_13233);
and U13428 (N_13428,N_13256,N_13272);
nor U13429 (N_13429,N_13243,N_13258);
and U13430 (N_13430,N_13278,N_13295);
or U13431 (N_13431,N_13254,N_13342);
nand U13432 (N_13432,N_13273,N_13228);
or U13433 (N_13433,N_13250,N_13343);
or U13434 (N_13434,N_13290,N_13265);
nor U13435 (N_13435,N_13277,N_13333);
or U13436 (N_13436,N_13332,N_13239);
and U13437 (N_13437,N_13295,N_13258);
and U13438 (N_13438,N_13328,N_13298);
xor U13439 (N_13439,N_13298,N_13259);
nand U13440 (N_13440,N_13296,N_13270);
and U13441 (N_13441,N_13279,N_13268);
xnor U13442 (N_13442,N_13313,N_13232);
nand U13443 (N_13443,N_13253,N_13224);
and U13444 (N_13444,N_13304,N_13261);
xnor U13445 (N_13445,N_13244,N_13331);
nor U13446 (N_13446,N_13235,N_13229);
or U13447 (N_13447,N_13201,N_13251);
and U13448 (N_13448,N_13338,N_13325);
or U13449 (N_13449,N_13291,N_13335);
nor U13450 (N_13450,N_13211,N_13304);
nand U13451 (N_13451,N_13275,N_13303);
xor U13452 (N_13452,N_13342,N_13282);
nor U13453 (N_13453,N_13296,N_13271);
xnor U13454 (N_13454,N_13227,N_13244);
and U13455 (N_13455,N_13344,N_13282);
nor U13456 (N_13456,N_13243,N_13344);
nor U13457 (N_13457,N_13323,N_13308);
nor U13458 (N_13458,N_13212,N_13279);
nand U13459 (N_13459,N_13209,N_13242);
or U13460 (N_13460,N_13262,N_13226);
nand U13461 (N_13461,N_13283,N_13265);
nand U13462 (N_13462,N_13339,N_13312);
nor U13463 (N_13463,N_13241,N_13259);
nand U13464 (N_13464,N_13331,N_13208);
xnor U13465 (N_13465,N_13312,N_13316);
and U13466 (N_13466,N_13341,N_13274);
nand U13467 (N_13467,N_13257,N_13283);
nand U13468 (N_13468,N_13345,N_13324);
or U13469 (N_13469,N_13247,N_13220);
nor U13470 (N_13470,N_13304,N_13290);
xnor U13471 (N_13471,N_13277,N_13241);
nor U13472 (N_13472,N_13229,N_13219);
or U13473 (N_13473,N_13288,N_13308);
and U13474 (N_13474,N_13223,N_13333);
nand U13475 (N_13475,N_13280,N_13200);
or U13476 (N_13476,N_13278,N_13325);
xor U13477 (N_13477,N_13277,N_13310);
nand U13478 (N_13478,N_13337,N_13341);
or U13479 (N_13479,N_13224,N_13234);
nor U13480 (N_13480,N_13326,N_13212);
or U13481 (N_13481,N_13309,N_13218);
xnor U13482 (N_13482,N_13339,N_13299);
nand U13483 (N_13483,N_13269,N_13311);
or U13484 (N_13484,N_13213,N_13277);
nand U13485 (N_13485,N_13329,N_13248);
and U13486 (N_13486,N_13206,N_13300);
and U13487 (N_13487,N_13323,N_13276);
xor U13488 (N_13488,N_13228,N_13337);
and U13489 (N_13489,N_13308,N_13324);
nand U13490 (N_13490,N_13240,N_13313);
or U13491 (N_13491,N_13244,N_13305);
xor U13492 (N_13492,N_13317,N_13307);
xnor U13493 (N_13493,N_13349,N_13314);
nor U13494 (N_13494,N_13201,N_13298);
or U13495 (N_13495,N_13203,N_13340);
nor U13496 (N_13496,N_13264,N_13273);
and U13497 (N_13497,N_13278,N_13263);
nand U13498 (N_13498,N_13272,N_13270);
nand U13499 (N_13499,N_13202,N_13240);
nor U13500 (N_13500,N_13378,N_13479);
and U13501 (N_13501,N_13470,N_13476);
and U13502 (N_13502,N_13401,N_13362);
nor U13503 (N_13503,N_13386,N_13391);
xnor U13504 (N_13504,N_13357,N_13413);
nand U13505 (N_13505,N_13404,N_13383);
xnor U13506 (N_13506,N_13465,N_13380);
xor U13507 (N_13507,N_13405,N_13367);
and U13508 (N_13508,N_13381,N_13353);
nor U13509 (N_13509,N_13359,N_13395);
nor U13510 (N_13510,N_13435,N_13365);
and U13511 (N_13511,N_13437,N_13369);
nor U13512 (N_13512,N_13416,N_13373);
nand U13513 (N_13513,N_13471,N_13429);
or U13514 (N_13514,N_13419,N_13450);
or U13515 (N_13515,N_13432,N_13461);
or U13516 (N_13516,N_13485,N_13393);
nor U13517 (N_13517,N_13441,N_13451);
nor U13518 (N_13518,N_13350,N_13411);
or U13519 (N_13519,N_13444,N_13370);
or U13520 (N_13520,N_13418,N_13371);
or U13521 (N_13521,N_13354,N_13430);
or U13522 (N_13522,N_13448,N_13403);
and U13523 (N_13523,N_13466,N_13488);
xnor U13524 (N_13524,N_13460,N_13385);
nor U13525 (N_13525,N_13421,N_13355);
and U13526 (N_13526,N_13374,N_13422);
or U13527 (N_13527,N_13425,N_13377);
nor U13528 (N_13528,N_13462,N_13472);
nand U13529 (N_13529,N_13474,N_13475);
or U13530 (N_13530,N_13487,N_13478);
nor U13531 (N_13531,N_13351,N_13452);
xor U13532 (N_13532,N_13449,N_13490);
nor U13533 (N_13533,N_13440,N_13439);
or U13534 (N_13534,N_13483,N_13356);
nor U13535 (N_13535,N_13360,N_13469);
nand U13536 (N_13536,N_13406,N_13398);
nand U13537 (N_13537,N_13396,N_13494);
xnor U13538 (N_13538,N_13443,N_13455);
nor U13539 (N_13539,N_13489,N_13394);
and U13540 (N_13540,N_13493,N_13454);
or U13541 (N_13541,N_13467,N_13453);
or U13542 (N_13542,N_13361,N_13482);
xnor U13543 (N_13543,N_13447,N_13400);
or U13544 (N_13544,N_13410,N_13388);
or U13545 (N_13545,N_13468,N_13375);
and U13546 (N_13546,N_13473,N_13408);
and U13547 (N_13547,N_13442,N_13481);
nand U13548 (N_13548,N_13382,N_13423);
xnor U13549 (N_13549,N_13428,N_13415);
or U13550 (N_13550,N_13499,N_13376);
xnor U13551 (N_13551,N_13379,N_13392);
nor U13552 (N_13552,N_13399,N_13497);
and U13553 (N_13553,N_13389,N_13420);
and U13554 (N_13554,N_13434,N_13484);
xor U13555 (N_13555,N_13456,N_13464);
and U13556 (N_13556,N_13352,N_13463);
and U13557 (N_13557,N_13477,N_13417);
nor U13558 (N_13558,N_13364,N_13431);
or U13559 (N_13559,N_13433,N_13445);
or U13560 (N_13560,N_13491,N_13409);
nand U13561 (N_13561,N_13402,N_13366);
or U13562 (N_13562,N_13480,N_13372);
nand U13563 (N_13563,N_13436,N_13384);
nor U13564 (N_13564,N_13426,N_13486);
xor U13565 (N_13565,N_13390,N_13358);
and U13566 (N_13566,N_13446,N_13438);
xnor U13567 (N_13567,N_13492,N_13496);
or U13568 (N_13568,N_13363,N_13414);
nor U13569 (N_13569,N_13495,N_13368);
or U13570 (N_13570,N_13412,N_13387);
or U13571 (N_13571,N_13427,N_13407);
or U13572 (N_13572,N_13397,N_13459);
nand U13573 (N_13573,N_13458,N_13457);
or U13574 (N_13574,N_13424,N_13498);
nor U13575 (N_13575,N_13463,N_13454);
nand U13576 (N_13576,N_13390,N_13480);
or U13577 (N_13577,N_13364,N_13357);
or U13578 (N_13578,N_13417,N_13445);
xnor U13579 (N_13579,N_13407,N_13484);
and U13580 (N_13580,N_13403,N_13447);
nand U13581 (N_13581,N_13441,N_13432);
nand U13582 (N_13582,N_13457,N_13405);
and U13583 (N_13583,N_13482,N_13490);
or U13584 (N_13584,N_13449,N_13381);
or U13585 (N_13585,N_13418,N_13445);
and U13586 (N_13586,N_13469,N_13373);
xnor U13587 (N_13587,N_13497,N_13429);
or U13588 (N_13588,N_13414,N_13397);
xor U13589 (N_13589,N_13490,N_13498);
nor U13590 (N_13590,N_13490,N_13389);
nor U13591 (N_13591,N_13466,N_13438);
nand U13592 (N_13592,N_13450,N_13487);
nor U13593 (N_13593,N_13457,N_13436);
or U13594 (N_13594,N_13464,N_13373);
or U13595 (N_13595,N_13441,N_13490);
xor U13596 (N_13596,N_13473,N_13369);
xnor U13597 (N_13597,N_13392,N_13439);
xnor U13598 (N_13598,N_13366,N_13446);
nor U13599 (N_13599,N_13377,N_13363);
nand U13600 (N_13600,N_13397,N_13418);
xnor U13601 (N_13601,N_13389,N_13427);
xnor U13602 (N_13602,N_13478,N_13463);
or U13603 (N_13603,N_13486,N_13450);
or U13604 (N_13604,N_13438,N_13490);
and U13605 (N_13605,N_13477,N_13375);
and U13606 (N_13606,N_13382,N_13353);
nand U13607 (N_13607,N_13417,N_13455);
and U13608 (N_13608,N_13403,N_13365);
and U13609 (N_13609,N_13481,N_13425);
and U13610 (N_13610,N_13429,N_13374);
and U13611 (N_13611,N_13397,N_13352);
and U13612 (N_13612,N_13375,N_13459);
nand U13613 (N_13613,N_13478,N_13362);
nor U13614 (N_13614,N_13356,N_13373);
and U13615 (N_13615,N_13405,N_13425);
xnor U13616 (N_13616,N_13486,N_13476);
nand U13617 (N_13617,N_13467,N_13353);
and U13618 (N_13618,N_13496,N_13455);
nor U13619 (N_13619,N_13365,N_13448);
nor U13620 (N_13620,N_13359,N_13389);
xor U13621 (N_13621,N_13468,N_13485);
and U13622 (N_13622,N_13409,N_13443);
xor U13623 (N_13623,N_13470,N_13496);
nand U13624 (N_13624,N_13499,N_13440);
nor U13625 (N_13625,N_13498,N_13473);
nor U13626 (N_13626,N_13487,N_13394);
or U13627 (N_13627,N_13453,N_13395);
or U13628 (N_13628,N_13431,N_13471);
nor U13629 (N_13629,N_13423,N_13493);
xnor U13630 (N_13630,N_13437,N_13353);
nand U13631 (N_13631,N_13487,N_13369);
nor U13632 (N_13632,N_13480,N_13436);
xor U13633 (N_13633,N_13424,N_13364);
nand U13634 (N_13634,N_13390,N_13471);
xor U13635 (N_13635,N_13378,N_13352);
xor U13636 (N_13636,N_13375,N_13361);
or U13637 (N_13637,N_13469,N_13441);
xnor U13638 (N_13638,N_13389,N_13426);
or U13639 (N_13639,N_13351,N_13353);
nor U13640 (N_13640,N_13396,N_13497);
nor U13641 (N_13641,N_13456,N_13484);
and U13642 (N_13642,N_13425,N_13482);
nor U13643 (N_13643,N_13395,N_13445);
xnor U13644 (N_13644,N_13497,N_13473);
xnor U13645 (N_13645,N_13479,N_13386);
and U13646 (N_13646,N_13478,N_13442);
or U13647 (N_13647,N_13479,N_13499);
nand U13648 (N_13648,N_13474,N_13403);
nand U13649 (N_13649,N_13362,N_13353);
nand U13650 (N_13650,N_13606,N_13555);
xor U13651 (N_13651,N_13538,N_13544);
xor U13652 (N_13652,N_13515,N_13605);
nor U13653 (N_13653,N_13579,N_13576);
or U13654 (N_13654,N_13560,N_13573);
and U13655 (N_13655,N_13589,N_13626);
and U13656 (N_13656,N_13604,N_13612);
nand U13657 (N_13657,N_13595,N_13556);
nand U13658 (N_13658,N_13549,N_13533);
and U13659 (N_13659,N_13565,N_13582);
xnor U13660 (N_13660,N_13586,N_13599);
or U13661 (N_13661,N_13639,N_13646);
nor U13662 (N_13662,N_13553,N_13510);
xor U13663 (N_13663,N_13640,N_13545);
and U13664 (N_13664,N_13516,N_13504);
nor U13665 (N_13665,N_13506,N_13524);
xnor U13666 (N_13666,N_13642,N_13601);
or U13667 (N_13667,N_13641,N_13630);
nor U13668 (N_13668,N_13539,N_13645);
xnor U13669 (N_13669,N_13534,N_13648);
nor U13670 (N_13670,N_13591,N_13634);
xor U13671 (N_13671,N_13611,N_13578);
and U13672 (N_13672,N_13546,N_13531);
nor U13673 (N_13673,N_13637,N_13632);
or U13674 (N_13674,N_13629,N_13529);
xor U13675 (N_13675,N_13572,N_13503);
or U13676 (N_13676,N_13532,N_13603);
nand U13677 (N_13677,N_13547,N_13541);
nand U13678 (N_13678,N_13635,N_13600);
and U13679 (N_13679,N_13557,N_13624);
nor U13680 (N_13680,N_13574,N_13644);
xor U13681 (N_13681,N_13633,N_13602);
nor U13682 (N_13682,N_13625,N_13583);
nor U13683 (N_13683,N_13563,N_13518);
and U13684 (N_13684,N_13543,N_13527);
or U13685 (N_13685,N_13567,N_13592);
nor U13686 (N_13686,N_13550,N_13571);
nand U13687 (N_13687,N_13614,N_13566);
nor U13688 (N_13688,N_13535,N_13581);
or U13689 (N_13689,N_13525,N_13522);
and U13690 (N_13690,N_13521,N_13569);
nand U13691 (N_13691,N_13559,N_13638);
nand U13692 (N_13692,N_13508,N_13613);
and U13693 (N_13693,N_13537,N_13500);
or U13694 (N_13694,N_13540,N_13584);
nand U13695 (N_13695,N_13501,N_13615);
nor U13696 (N_13696,N_13607,N_13643);
nand U13697 (N_13697,N_13519,N_13616);
or U13698 (N_13698,N_13621,N_13505);
xnor U13699 (N_13699,N_13608,N_13530);
xnor U13700 (N_13700,N_13552,N_13507);
and U13701 (N_13701,N_13561,N_13517);
nand U13702 (N_13702,N_13588,N_13628);
nand U13703 (N_13703,N_13587,N_13511);
nand U13704 (N_13704,N_13514,N_13528);
and U13705 (N_13705,N_13627,N_13593);
xor U13706 (N_13706,N_13523,N_13623);
xnor U13707 (N_13707,N_13568,N_13597);
and U13708 (N_13708,N_13619,N_13610);
xnor U13709 (N_13709,N_13649,N_13647);
xnor U13710 (N_13710,N_13548,N_13596);
or U13711 (N_13711,N_13622,N_13585);
nand U13712 (N_13712,N_13575,N_13620);
xor U13713 (N_13713,N_13520,N_13509);
and U13714 (N_13714,N_13636,N_13558);
nand U13715 (N_13715,N_13570,N_13513);
or U13716 (N_13716,N_13631,N_13554);
and U13717 (N_13717,N_13526,N_13617);
xnor U13718 (N_13718,N_13609,N_13562);
or U13719 (N_13719,N_13502,N_13564);
xnor U13720 (N_13720,N_13577,N_13551);
nor U13721 (N_13721,N_13594,N_13536);
nand U13722 (N_13722,N_13580,N_13512);
or U13723 (N_13723,N_13590,N_13618);
or U13724 (N_13724,N_13542,N_13598);
and U13725 (N_13725,N_13567,N_13636);
xor U13726 (N_13726,N_13540,N_13646);
nor U13727 (N_13727,N_13614,N_13537);
nand U13728 (N_13728,N_13568,N_13592);
and U13729 (N_13729,N_13616,N_13543);
nor U13730 (N_13730,N_13647,N_13623);
nand U13731 (N_13731,N_13527,N_13627);
nor U13732 (N_13732,N_13546,N_13551);
nand U13733 (N_13733,N_13516,N_13557);
or U13734 (N_13734,N_13649,N_13506);
nand U13735 (N_13735,N_13605,N_13517);
nand U13736 (N_13736,N_13636,N_13549);
or U13737 (N_13737,N_13641,N_13636);
or U13738 (N_13738,N_13625,N_13621);
nand U13739 (N_13739,N_13523,N_13590);
or U13740 (N_13740,N_13597,N_13585);
or U13741 (N_13741,N_13539,N_13569);
nor U13742 (N_13742,N_13585,N_13642);
nand U13743 (N_13743,N_13516,N_13509);
nand U13744 (N_13744,N_13572,N_13511);
xnor U13745 (N_13745,N_13626,N_13523);
xor U13746 (N_13746,N_13639,N_13574);
or U13747 (N_13747,N_13519,N_13592);
nor U13748 (N_13748,N_13569,N_13555);
xor U13749 (N_13749,N_13631,N_13550);
and U13750 (N_13750,N_13555,N_13644);
or U13751 (N_13751,N_13584,N_13647);
and U13752 (N_13752,N_13552,N_13530);
or U13753 (N_13753,N_13597,N_13594);
and U13754 (N_13754,N_13541,N_13556);
and U13755 (N_13755,N_13570,N_13506);
nor U13756 (N_13756,N_13622,N_13506);
nand U13757 (N_13757,N_13565,N_13638);
or U13758 (N_13758,N_13534,N_13642);
or U13759 (N_13759,N_13549,N_13542);
nand U13760 (N_13760,N_13541,N_13643);
or U13761 (N_13761,N_13608,N_13561);
nand U13762 (N_13762,N_13506,N_13518);
or U13763 (N_13763,N_13637,N_13628);
or U13764 (N_13764,N_13522,N_13649);
nor U13765 (N_13765,N_13589,N_13554);
nor U13766 (N_13766,N_13635,N_13505);
nand U13767 (N_13767,N_13596,N_13589);
or U13768 (N_13768,N_13510,N_13591);
and U13769 (N_13769,N_13506,N_13521);
nor U13770 (N_13770,N_13574,N_13576);
and U13771 (N_13771,N_13516,N_13639);
xor U13772 (N_13772,N_13503,N_13580);
xnor U13773 (N_13773,N_13548,N_13606);
and U13774 (N_13774,N_13562,N_13510);
or U13775 (N_13775,N_13504,N_13579);
or U13776 (N_13776,N_13573,N_13509);
or U13777 (N_13777,N_13602,N_13611);
nand U13778 (N_13778,N_13542,N_13604);
and U13779 (N_13779,N_13532,N_13535);
xor U13780 (N_13780,N_13523,N_13521);
or U13781 (N_13781,N_13585,N_13502);
xnor U13782 (N_13782,N_13634,N_13513);
nand U13783 (N_13783,N_13545,N_13556);
or U13784 (N_13784,N_13633,N_13533);
and U13785 (N_13785,N_13508,N_13563);
xor U13786 (N_13786,N_13515,N_13607);
and U13787 (N_13787,N_13514,N_13619);
nor U13788 (N_13788,N_13622,N_13594);
nor U13789 (N_13789,N_13615,N_13541);
xnor U13790 (N_13790,N_13623,N_13637);
xnor U13791 (N_13791,N_13504,N_13559);
nor U13792 (N_13792,N_13552,N_13532);
or U13793 (N_13793,N_13562,N_13502);
nand U13794 (N_13794,N_13614,N_13519);
nor U13795 (N_13795,N_13545,N_13536);
and U13796 (N_13796,N_13594,N_13554);
xor U13797 (N_13797,N_13525,N_13605);
nand U13798 (N_13798,N_13630,N_13566);
xnor U13799 (N_13799,N_13648,N_13640);
xor U13800 (N_13800,N_13741,N_13751);
nand U13801 (N_13801,N_13670,N_13681);
xor U13802 (N_13802,N_13686,N_13688);
or U13803 (N_13803,N_13661,N_13668);
or U13804 (N_13804,N_13746,N_13710);
and U13805 (N_13805,N_13750,N_13764);
nand U13806 (N_13806,N_13684,N_13709);
or U13807 (N_13807,N_13669,N_13716);
nand U13808 (N_13808,N_13776,N_13725);
xor U13809 (N_13809,N_13728,N_13656);
nand U13810 (N_13810,N_13791,N_13671);
and U13811 (N_13811,N_13753,N_13678);
xnor U13812 (N_13812,N_13650,N_13660);
xnor U13813 (N_13813,N_13754,N_13722);
xnor U13814 (N_13814,N_13667,N_13677);
nor U13815 (N_13815,N_13798,N_13740);
and U13816 (N_13816,N_13729,N_13745);
xor U13817 (N_13817,N_13666,N_13659);
xnor U13818 (N_13818,N_13773,N_13760);
and U13819 (N_13819,N_13654,N_13711);
or U13820 (N_13820,N_13782,N_13763);
nand U13821 (N_13821,N_13736,N_13733);
nand U13822 (N_13822,N_13738,N_13663);
xnor U13823 (N_13823,N_13685,N_13653);
nor U13824 (N_13824,N_13689,N_13757);
nor U13825 (N_13825,N_13680,N_13726);
xnor U13826 (N_13826,N_13713,N_13690);
or U13827 (N_13827,N_13698,N_13702);
nand U13828 (N_13828,N_13752,N_13775);
nor U13829 (N_13829,N_13693,N_13789);
or U13830 (N_13830,N_13735,N_13767);
or U13831 (N_13831,N_13774,N_13703);
or U13832 (N_13832,N_13694,N_13714);
nor U13833 (N_13833,N_13664,N_13687);
or U13834 (N_13834,N_13717,N_13796);
and U13835 (N_13835,N_13720,N_13744);
or U13836 (N_13836,N_13692,N_13781);
xnor U13837 (N_13837,N_13742,N_13759);
or U13838 (N_13838,N_13734,N_13718);
or U13839 (N_13839,N_13665,N_13793);
and U13840 (N_13840,N_13657,N_13758);
or U13841 (N_13841,N_13780,N_13795);
nand U13842 (N_13842,N_13769,N_13790);
xnor U13843 (N_13843,N_13679,N_13676);
nand U13844 (N_13844,N_13785,N_13699);
xnor U13845 (N_13845,N_13797,N_13705);
and U13846 (N_13846,N_13674,N_13675);
nor U13847 (N_13847,N_13731,N_13655);
nand U13848 (N_13848,N_13771,N_13682);
or U13849 (N_13849,N_13697,N_13770);
and U13850 (N_13850,N_13786,N_13787);
and U13851 (N_13851,N_13691,N_13652);
nand U13852 (N_13852,N_13730,N_13712);
nor U13853 (N_13853,N_13700,N_13778);
and U13854 (N_13854,N_13799,N_13755);
xnor U13855 (N_13855,N_13766,N_13715);
xnor U13856 (N_13856,N_13761,N_13777);
or U13857 (N_13857,N_13662,N_13792);
xnor U13858 (N_13858,N_13743,N_13707);
nand U13859 (N_13859,N_13708,N_13784);
nand U13860 (N_13860,N_13772,N_13695);
or U13861 (N_13861,N_13658,N_13756);
nor U13862 (N_13862,N_13721,N_13794);
and U13863 (N_13863,N_13724,N_13747);
nor U13864 (N_13864,N_13749,N_13783);
or U13865 (N_13865,N_13739,N_13706);
nand U13866 (N_13866,N_13701,N_13768);
and U13867 (N_13867,N_13696,N_13737);
xor U13868 (N_13868,N_13683,N_13719);
nor U13869 (N_13869,N_13673,N_13672);
nor U13870 (N_13870,N_13651,N_13779);
nand U13871 (N_13871,N_13765,N_13723);
nand U13872 (N_13872,N_13704,N_13732);
nor U13873 (N_13873,N_13748,N_13788);
nand U13874 (N_13874,N_13727,N_13762);
and U13875 (N_13875,N_13690,N_13663);
nand U13876 (N_13876,N_13767,N_13667);
or U13877 (N_13877,N_13739,N_13662);
nor U13878 (N_13878,N_13742,N_13693);
or U13879 (N_13879,N_13687,N_13700);
nor U13880 (N_13880,N_13655,N_13760);
xnor U13881 (N_13881,N_13689,N_13739);
nand U13882 (N_13882,N_13695,N_13756);
xor U13883 (N_13883,N_13760,N_13736);
or U13884 (N_13884,N_13774,N_13791);
xnor U13885 (N_13885,N_13688,N_13716);
xnor U13886 (N_13886,N_13710,N_13742);
nand U13887 (N_13887,N_13745,N_13669);
nand U13888 (N_13888,N_13699,N_13704);
and U13889 (N_13889,N_13759,N_13767);
nand U13890 (N_13890,N_13759,N_13666);
xnor U13891 (N_13891,N_13653,N_13748);
and U13892 (N_13892,N_13782,N_13732);
or U13893 (N_13893,N_13719,N_13755);
nand U13894 (N_13894,N_13739,N_13763);
and U13895 (N_13895,N_13788,N_13711);
nand U13896 (N_13896,N_13658,N_13695);
xor U13897 (N_13897,N_13772,N_13782);
nor U13898 (N_13898,N_13737,N_13709);
xnor U13899 (N_13899,N_13745,N_13785);
nand U13900 (N_13900,N_13718,N_13714);
nand U13901 (N_13901,N_13778,N_13794);
nor U13902 (N_13902,N_13687,N_13791);
nor U13903 (N_13903,N_13795,N_13723);
nand U13904 (N_13904,N_13793,N_13766);
or U13905 (N_13905,N_13755,N_13690);
xnor U13906 (N_13906,N_13692,N_13752);
xor U13907 (N_13907,N_13784,N_13693);
and U13908 (N_13908,N_13765,N_13683);
or U13909 (N_13909,N_13667,N_13775);
nand U13910 (N_13910,N_13650,N_13746);
or U13911 (N_13911,N_13731,N_13709);
and U13912 (N_13912,N_13690,N_13772);
or U13913 (N_13913,N_13708,N_13683);
or U13914 (N_13914,N_13694,N_13661);
xnor U13915 (N_13915,N_13680,N_13690);
or U13916 (N_13916,N_13781,N_13765);
nor U13917 (N_13917,N_13681,N_13778);
nor U13918 (N_13918,N_13789,N_13746);
xnor U13919 (N_13919,N_13757,N_13658);
or U13920 (N_13920,N_13767,N_13778);
xnor U13921 (N_13921,N_13711,N_13748);
nand U13922 (N_13922,N_13738,N_13789);
and U13923 (N_13923,N_13680,N_13783);
xor U13924 (N_13924,N_13711,N_13652);
and U13925 (N_13925,N_13782,N_13771);
nor U13926 (N_13926,N_13688,N_13770);
and U13927 (N_13927,N_13665,N_13743);
or U13928 (N_13928,N_13700,N_13675);
nor U13929 (N_13929,N_13775,N_13710);
nor U13930 (N_13930,N_13666,N_13744);
nor U13931 (N_13931,N_13769,N_13719);
nand U13932 (N_13932,N_13791,N_13739);
and U13933 (N_13933,N_13795,N_13776);
nand U13934 (N_13934,N_13703,N_13657);
and U13935 (N_13935,N_13676,N_13695);
nand U13936 (N_13936,N_13695,N_13797);
and U13937 (N_13937,N_13747,N_13707);
xnor U13938 (N_13938,N_13672,N_13793);
xnor U13939 (N_13939,N_13736,N_13798);
or U13940 (N_13940,N_13726,N_13655);
or U13941 (N_13941,N_13751,N_13760);
nor U13942 (N_13942,N_13766,N_13713);
and U13943 (N_13943,N_13664,N_13792);
nor U13944 (N_13944,N_13797,N_13716);
xor U13945 (N_13945,N_13703,N_13744);
xor U13946 (N_13946,N_13733,N_13731);
nor U13947 (N_13947,N_13795,N_13697);
and U13948 (N_13948,N_13663,N_13654);
and U13949 (N_13949,N_13654,N_13668);
and U13950 (N_13950,N_13826,N_13885);
xnor U13951 (N_13951,N_13869,N_13859);
xnor U13952 (N_13952,N_13866,N_13831);
and U13953 (N_13953,N_13895,N_13824);
nor U13954 (N_13954,N_13883,N_13843);
nand U13955 (N_13955,N_13941,N_13891);
xnor U13956 (N_13956,N_13870,N_13809);
xnor U13957 (N_13957,N_13898,N_13886);
xnor U13958 (N_13958,N_13838,N_13821);
xor U13959 (N_13959,N_13915,N_13935);
and U13960 (N_13960,N_13832,N_13827);
nand U13961 (N_13961,N_13939,N_13911);
nor U13962 (N_13962,N_13892,N_13855);
nand U13963 (N_13963,N_13852,N_13874);
xor U13964 (N_13964,N_13848,N_13919);
or U13965 (N_13965,N_13924,N_13921);
and U13966 (N_13966,N_13867,N_13890);
nor U13967 (N_13967,N_13850,N_13808);
nor U13968 (N_13968,N_13815,N_13948);
or U13969 (N_13969,N_13925,N_13835);
or U13970 (N_13970,N_13912,N_13871);
nor U13971 (N_13971,N_13825,N_13909);
xor U13972 (N_13972,N_13899,N_13929);
or U13973 (N_13973,N_13856,N_13907);
and U13974 (N_13974,N_13932,N_13837);
or U13975 (N_13975,N_13936,N_13849);
nor U13976 (N_13976,N_13940,N_13946);
nand U13977 (N_13977,N_13851,N_13902);
and U13978 (N_13978,N_13931,N_13914);
nor U13979 (N_13979,N_13860,N_13893);
nor U13980 (N_13980,N_13853,N_13820);
nand U13981 (N_13981,N_13830,N_13880);
nor U13982 (N_13982,N_13805,N_13842);
and U13983 (N_13983,N_13845,N_13943);
nor U13984 (N_13984,N_13888,N_13889);
xor U13985 (N_13985,N_13814,N_13872);
and U13986 (N_13986,N_13829,N_13844);
nor U13987 (N_13987,N_13882,N_13894);
and U13988 (N_13988,N_13910,N_13807);
nor U13989 (N_13989,N_13938,N_13896);
xnor U13990 (N_13990,N_13822,N_13873);
nand U13991 (N_13991,N_13933,N_13944);
xor U13992 (N_13992,N_13916,N_13813);
xnor U13993 (N_13993,N_13828,N_13801);
or U13994 (N_13994,N_13854,N_13857);
nor U13995 (N_13995,N_13811,N_13803);
or U13996 (N_13996,N_13865,N_13881);
or U13997 (N_13997,N_13934,N_13875);
and U13998 (N_13998,N_13818,N_13858);
nand U13999 (N_13999,N_13800,N_13841);
and U14000 (N_14000,N_13804,N_13864);
and U14001 (N_14001,N_13908,N_13819);
or U14002 (N_14002,N_13922,N_13812);
xnor U14003 (N_14003,N_13897,N_13868);
nor U14004 (N_14004,N_13802,N_13817);
nand U14005 (N_14005,N_13879,N_13913);
nor U14006 (N_14006,N_13836,N_13945);
or U14007 (N_14007,N_13903,N_13878);
xnor U14008 (N_14008,N_13917,N_13937);
or U14009 (N_14009,N_13863,N_13923);
nor U14010 (N_14010,N_13920,N_13806);
and U14011 (N_14011,N_13877,N_13833);
nand U14012 (N_14012,N_13846,N_13839);
or U14013 (N_14013,N_13949,N_13900);
nand U14014 (N_14014,N_13876,N_13810);
or U14015 (N_14015,N_13904,N_13942);
and U14016 (N_14016,N_13847,N_13884);
xor U14017 (N_14017,N_13928,N_13823);
nor U14018 (N_14018,N_13887,N_13926);
and U14019 (N_14019,N_13906,N_13901);
nor U14020 (N_14020,N_13918,N_13861);
xor U14021 (N_14021,N_13816,N_13862);
or U14022 (N_14022,N_13930,N_13834);
nor U14023 (N_14023,N_13905,N_13840);
nand U14024 (N_14024,N_13947,N_13927);
nor U14025 (N_14025,N_13837,N_13824);
nor U14026 (N_14026,N_13889,N_13864);
nor U14027 (N_14027,N_13925,N_13905);
or U14028 (N_14028,N_13830,N_13823);
xor U14029 (N_14029,N_13832,N_13917);
and U14030 (N_14030,N_13932,N_13854);
xor U14031 (N_14031,N_13862,N_13945);
nor U14032 (N_14032,N_13911,N_13892);
and U14033 (N_14033,N_13863,N_13838);
or U14034 (N_14034,N_13924,N_13930);
and U14035 (N_14035,N_13934,N_13836);
xnor U14036 (N_14036,N_13884,N_13880);
or U14037 (N_14037,N_13861,N_13919);
and U14038 (N_14038,N_13871,N_13816);
nor U14039 (N_14039,N_13865,N_13931);
nand U14040 (N_14040,N_13937,N_13912);
or U14041 (N_14041,N_13879,N_13878);
or U14042 (N_14042,N_13874,N_13902);
or U14043 (N_14043,N_13817,N_13922);
nand U14044 (N_14044,N_13854,N_13871);
or U14045 (N_14045,N_13871,N_13801);
nor U14046 (N_14046,N_13892,N_13877);
xor U14047 (N_14047,N_13837,N_13848);
and U14048 (N_14048,N_13891,N_13920);
and U14049 (N_14049,N_13836,N_13844);
xor U14050 (N_14050,N_13801,N_13884);
nand U14051 (N_14051,N_13830,N_13910);
xor U14052 (N_14052,N_13928,N_13803);
nor U14053 (N_14053,N_13886,N_13868);
and U14054 (N_14054,N_13843,N_13865);
nand U14055 (N_14055,N_13815,N_13843);
nor U14056 (N_14056,N_13891,N_13837);
and U14057 (N_14057,N_13800,N_13942);
xnor U14058 (N_14058,N_13931,N_13909);
nand U14059 (N_14059,N_13895,N_13861);
nand U14060 (N_14060,N_13856,N_13823);
xnor U14061 (N_14061,N_13936,N_13831);
and U14062 (N_14062,N_13818,N_13804);
or U14063 (N_14063,N_13901,N_13880);
or U14064 (N_14064,N_13854,N_13900);
and U14065 (N_14065,N_13917,N_13814);
xnor U14066 (N_14066,N_13929,N_13866);
nor U14067 (N_14067,N_13813,N_13898);
xor U14068 (N_14068,N_13912,N_13898);
or U14069 (N_14069,N_13937,N_13802);
or U14070 (N_14070,N_13911,N_13830);
or U14071 (N_14071,N_13861,N_13920);
nor U14072 (N_14072,N_13850,N_13805);
nand U14073 (N_14073,N_13916,N_13841);
and U14074 (N_14074,N_13856,N_13810);
and U14075 (N_14075,N_13847,N_13920);
or U14076 (N_14076,N_13870,N_13894);
nand U14077 (N_14077,N_13858,N_13910);
xnor U14078 (N_14078,N_13877,N_13862);
and U14079 (N_14079,N_13869,N_13858);
or U14080 (N_14080,N_13902,N_13822);
and U14081 (N_14081,N_13815,N_13848);
and U14082 (N_14082,N_13868,N_13902);
or U14083 (N_14083,N_13876,N_13880);
and U14084 (N_14084,N_13818,N_13820);
and U14085 (N_14085,N_13827,N_13852);
and U14086 (N_14086,N_13945,N_13848);
nand U14087 (N_14087,N_13930,N_13936);
and U14088 (N_14088,N_13865,N_13882);
nand U14089 (N_14089,N_13847,N_13891);
or U14090 (N_14090,N_13903,N_13816);
xnor U14091 (N_14091,N_13866,N_13949);
nand U14092 (N_14092,N_13823,N_13864);
and U14093 (N_14093,N_13827,N_13851);
or U14094 (N_14094,N_13937,N_13800);
nor U14095 (N_14095,N_13802,N_13801);
nand U14096 (N_14096,N_13944,N_13830);
or U14097 (N_14097,N_13931,N_13925);
nor U14098 (N_14098,N_13832,N_13830);
xnor U14099 (N_14099,N_13809,N_13886);
nand U14100 (N_14100,N_13961,N_14013);
and U14101 (N_14101,N_14052,N_13992);
and U14102 (N_14102,N_14086,N_14009);
nor U14103 (N_14103,N_14068,N_14006);
nor U14104 (N_14104,N_13991,N_13954);
nand U14105 (N_14105,N_14048,N_13990);
and U14106 (N_14106,N_14043,N_14044);
nor U14107 (N_14107,N_13964,N_14029);
nor U14108 (N_14108,N_14017,N_14089);
and U14109 (N_14109,N_14018,N_14032);
nand U14110 (N_14110,N_14078,N_13950);
xor U14111 (N_14111,N_14038,N_13985);
and U14112 (N_14112,N_13976,N_14080);
nand U14113 (N_14113,N_13957,N_14001);
and U14114 (N_14114,N_14058,N_14045);
or U14115 (N_14115,N_14099,N_13959);
xnor U14116 (N_14116,N_14010,N_14066);
xnor U14117 (N_14117,N_14035,N_14059);
nand U14118 (N_14118,N_14085,N_14008);
nor U14119 (N_14119,N_14019,N_14034);
or U14120 (N_14120,N_13958,N_14060);
or U14121 (N_14121,N_13970,N_13960);
nand U14122 (N_14122,N_14098,N_13993);
or U14123 (N_14123,N_13968,N_14051);
nor U14124 (N_14124,N_13971,N_14088);
or U14125 (N_14125,N_13978,N_13966);
or U14126 (N_14126,N_14083,N_14016);
and U14127 (N_14127,N_14037,N_14096);
nor U14128 (N_14128,N_14055,N_13967);
or U14129 (N_14129,N_14065,N_13986);
nand U14130 (N_14130,N_14030,N_14011);
or U14131 (N_14131,N_14069,N_13955);
and U14132 (N_14132,N_13994,N_13953);
nand U14133 (N_14133,N_14040,N_14095);
and U14134 (N_14134,N_13987,N_14061);
nand U14135 (N_14135,N_14076,N_14075);
xnor U14136 (N_14136,N_14046,N_14004);
nand U14137 (N_14137,N_14092,N_14015);
nand U14138 (N_14138,N_14014,N_13962);
or U14139 (N_14139,N_13983,N_14027);
nand U14140 (N_14140,N_14097,N_14062);
nand U14141 (N_14141,N_13988,N_13963);
xnor U14142 (N_14142,N_14023,N_14071);
xnor U14143 (N_14143,N_14000,N_13979);
and U14144 (N_14144,N_14082,N_14002);
or U14145 (N_14145,N_14081,N_14057);
xor U14146 (N_14146,N_14026,N_13975);
nor U14147 (N_14147,N_14064,N_14087);
or U14148 (N_14148,N_13999,N_13965);
or U14149 (N_14149,N_14028,N_14073);
nor U14150 (N_14150,N_14022,N_13989);
or U14151 (N_14151,N_14039,N_14041);
xnor U14152 (N_14152,N_13956,N_13973);
nand U14153 (N_14153,N_13972,N_13974);
or U14154 (N_14154,N_13998,N_14094);
nand U14155 (N_14155,N_14007,N_13969);
nand U14156 (N_14156,N_13996,N_14090);
nand U14157 (N_14157,N_13977,N_14024);
nor U14158 (N_14158,N_13980,N_13952);
nand U14159 (N_14159,N_14084,N_13997);
nand U14160 (N_14160,N_13951,N_14033);
or U14161 (N_14161,N_14020,N_14093);
xor U14162 (N_14162,N_14005,N_14070);
and U14163 (N_14163,N_14025,N_14053);
nor U14164 (N_14164,N_14079,N_14012);
or U14165 (N_14165,N_14056,N_14031);
nand U14166 (N_14166,N_14021,N_14047);
and U14167 (N_14167,N_14072,N_14036);
or U14168 (N_14168,N_14042,N_14063);
xnor U14169 (N_14169,N_14049,N_14067);
or U14170 (N_14170,N_13982,N_13981);
xnor U14171 (N_14171,N_14091,N_14050);
nor U14172 (N_14172,N_14074,N_13984);
and U14173 (N_14173,N_14003,N_13995);
and U14174 (N_14174,N_14054,N_14077);
nor U14175 (N_14175,N_14064,N_13987);
nand U14176 (N_14176,N_14014,N_13964);
xor U14177 (N_14177,N_13968,N_14070);
nand U14178 (N_14178,N_14036,N_13989);
and U14179 (N_14179,N_14052,N_14089);
nand U14180 (N_14180,N_14057,N_13974);
or U14181 (N_14181,N_13965,N_13975);
xnor U14182 (N_14182,N_13976,N_14086);
nand U14183 (N_14183,N_14086,N_13974);
xnor U14184 (N_14184,N_14044,N_14046);
and U14185 (N_14185,N_14034,N_14060);
nand U14186 (N_14186,N_14083,N_14048);
xor U14187 (N_14187,N_13951,N_14002);
and U14188 (N_14188,N_14020,N_13955);
nor U14189 (N_14189,N_13998,N_14023);
nor U14190 (N_14190,N_14062,N_13958);
nand U14191 (N_14191,N_14019,N_13959);
nand U14192 (N_14192,N_13963,N_13966);
nand U14193 (N_14193,N_14096,N_14086);
and U14194 (N_14194,N_14079,N_14092);
or U14195 (N_14195,N_14062,N_14038);
xor U14196 (N_14196,N_13989,N_14042);
or U14197 (N_14197,N_14008,N_14011);
nor U14198 (N_14198,N_13964,N_13968);
or U14199 (N_14199,N_14059,N_14072);
xor U14200 (N_14200,N_13971,N_14024);
or U14201 (N_14201,N_14041,N_14051);
xnor U14202 (N_14202,N_14085,N_14020);
or U14203 (N_14203,N_14009,N_13974);
nor U14204 (N_14204,N_14046,N_14036);
or U14205 (N_14205,N_14050,N_14083);
nor U14206 (N_14206,N_14000,N_13970);
xor U14207 (N_14207,N_13963,N_14052);
nand U14208 (N_14208,N_13979,N_13995);
xor U14209 (N_14209,N_13971,N_13992);
nor U14210 (N_14210,N_14014,N_13981);
nor U14211 (N_14211,N_13975,N_14025);
nand U14212 (N_14212,N_14078,N_14020);
or U14213 (N_14213,N_13957,N_14008);
nand U14214 (N_14214,N_14024,N_14097);
xnor U14215 (N_14215,N_14029,N_14073);
nor U14216 (N_14216,N_14095,N_14078);
xor U14217 (N_14217,N_14097,N_14064);
xor U14218 (N_14218,N_14036,N_13984);
and U14219 (N_14219,N_14017,N_13965);
nor U14220 (N_14220,N_14006,N_14046);
xnor U14221 (N_14221,N_14093,N_14076);
nand U14222 (N_14222,N_13965,N_14092);
nor U14223 (N_14223,N_13986,N_13970);
or U14224 (N_14224,N_13950,N_14025);
nor U14225 (N_14225,N_14026,N_14069);
xor U14226 (N_14226,N_14015,N_13987);
or U14227 (N_14227,N_14019,N_13982);
nor U14228 (N_14228,N_14020,N_14033);
nor U14229 (N_14229,N_14072,N_14062);
or U14230 (N_14230,N_14094,N_14086);
or U14231 (N_14231,N_14003,N_14026);
xor U14232 (N_14232,N_13977,N_14004);
and U14233 (N_14233,N_14037,N_13997);
xnor U14234 (N_14234,N_14047,N_13954);
xor U14235 (N_14235,N_13968,N_14030);
nor U14236 (N_14236,N_14068,N_14052);
nand U14237 (N_14237,N_14056,N_13990);
or U14238 (N_14238,N_13993,N_14085);
nor U14239 (N_14239,N_14068,N_13982);
and U14240 (N_14240,N_13955,N_13967);
nor U14241 (N_14241,N_14088,N_14057);
nor U14242 (N_14242,N_14096,N_14080);
nor U14243 (N_14243,N_14012,N_14001);
or U14244 (N_14244,N_14056,N_13992);
nor U14245 (N_14245,N_14023,N_14048);
or U14246 (N_14246,N_14065,N_13981);
xnor U14247 (N_14247,N_14085,N_14098);
nand U14248 (N_14248,N_13987,N_13996);
or U14249 (N_14249,N_14061,N_13989);
or U14250 (N_14250,N_14107,N_14105);
and U14251 (N_14251,N_14116,N_14104);
nor U14252 (N_14252,N_14192,N_14204);
and U14253 (N_14253,N_14194,N_14179);
or U14254 (N_14254,N_14103,N_14231);
or U14255 (N_14255,N_14111,N_14189);
nand U14256 (N_14256,N_14165,N_14223);
xnor U14257 (N_14257,N_14178,N_14222);
nand U14258 (N_14258,N_14201,N_14237);
and U14259 (N_14259,N_14124,N_14235);
and U14260 (N_14260,N_14206,N_14118);
or U14261 (N_14261,N_14173,N_14160);
xor U14262 (N_14262,N_14213,N_14159);
xor U14263 (N_14263,N_14123,N_14143);
nand U14264 (N_14264,N_14161,N_14154);
and U14265 (N_14265,N_14149,N_14207);
xnor U14266 (N_14266,N_14113,N_14114);
nand U14267 (N_14267,N_14140,N_14101);
xor U14268 (N_14268,N_14243,N_14247);
xnor U14269 (N_14269,N_14198,N_14153);
nand U14270 (N_14270,N_14164,N_14227);
or U14271 (N_14271,N_14144,N_14163);
nand U14272 (N_14272,N_14244,N_14112);
or U14273 (N_14273,N_14126,N_14193);
xnor U14274 (N_14274,N_14125,N_14249);
xor U14275 (N_14275,N_14229,N_14106);
nor U14276 (N_14276,N_14135,N_14129);
nand U14277 (N_14277,N_14128,N_14230);
and U14278 (N_14278,N_14172,N_14134);
or U14279 (N_14279,N_14174,N_14168);
nor U14280 (N_14280,N_14233,N_14148);
and U14281 (N_14281,N_14145,N_14182);
nor U14282 (N_14282,N_14132,N_14171);
and U14283 (N_14283,N_14209,N_14158);
nand U14284 (N_14284,N_14130,N_14219);
nor U14285 (N_14285,N_14208,N_14191);
nand U14286 (N_14286,N_14188,N_14131);
nor U14287 (N_14287,N_14226,N_14150);
nor U14288 (N_14288,N_14210,N_14175);
nand U14289 (N_14289,N_14157,N_14186);
nand U14290 (N_14290,N_14122,N_14166);
nor U14291 (N_14291,N_14248,N_14183);
xnor U14292 (N_14292,N_14127,N_14133);
nor U14293 (N_14293,N_14100,N_14121);
or U14294 (N_14294,N_14214,N_14176);
nand U14295 (N_14295,N_14202,N_14185);
and U14296 (N_14296,N_14180,N_14200);
and U14297 (N_14297,N_14108,N_14203);
nand U14298 (N_14298,N_14141,N_14246);
xnor U14299 (N_14299,N_14162,N_14218);
and U14300 (N_14300,N_14241,N_14199);
and U14301 (N_14301,N_14195,N_14196);
nor U14302 (N_14302,N_14102,N_14228);
xor U14303 (N_14303,N_14216,N_14137);
nor U14304 (N_14304,N_14110,N_14109);
or U14305 (N_14305,N_14138,N_14215);
and U14306 (N_14306,N_14245,N_14169);
nand U14307 (N_14307,N_14181,N_14119);
and U14308 (N_14308,N_14197,N_14221);
nand U14309 (N_14309,N_14238,N_14184);
xor U14310 (N_14310,N_14155,N_14220);
nand U14311 (N_14311,N_14146,N_14217);
and U14312 (N_14312,N_14170,N_14152);
nor U14313 (N_14313,N_14136,N_14236);
and U14314 (N_14314,N_14239,N_14115);
nand U14315 (N_14315,N_14147,N_14117);
and U14316 (N_14316,N_14212,N_14190);
xnor U14317 (N_14317,N_14225,N_14139);
or U14318 (N_14318,N_14156,N_14151);
or U14319 (N_14319,N_14120,N_14234);
or U14320 (N_14320,N_14167,N_14242);
and U14321 (N_14321,N_14232,N_14211);
nor U14322 (N_14322,N_14187,N_14205);
nand U14323 (N_14323,N_14224,N_14177);
nor U14324 (N_14324,N_14142,N_14240);
and U14325 (N_14325,N_14242,N_14221);
nand U14326 (N_14326,N_14229,N_14186);
xnor U14327 (N_14327,N_14134,N_14202);
xor U14328 (N_14328,N_14165,N_14242);
nor U14329 (N_14329,N_14112,N_14187);
nor U14330 (N_14330,N_14246,N_14145);
and U14331 (N_14331,N_14167,N_14113);
xnor U14332 (N_14332,N_14163,N_14175);
nor U14333 (N_14333,N_14203,N_14229);
and U14334 (N_14334,N_14127,N_14145);
or U14335 (N_14335,N_14170,N_14234);
nand U14336 (N_14336,N_14247,N_14192);
xor U14337 (N_14337,N_14185,N_14104);
or U14338 (N_14338,N_14241,N_14157);
nor U14339 (N_14339,N_14199,N_14202);
nand U14340 (N_14340,N_14110,N_14192);
and U14341 (N_14341,N_14240,N_14246);
nor U14342 (N_14342,N_14153,N_14139);
nor U14343 (N_14343,N_14247,N_14241);
xnor U14344 (N_14344,N_14108,N_14240);
xor U14345 (N_14345,N_14201,N_14133);
and U14346 (N_14346,N_14196,N_14182);
and U14347 (N_14347,N_14215,N_14134);
xnor U14348 (N_14348,N_14197,N_14234);
nand U14349 (N_14349,N_14159,N_14161);
or U14350 (N_14350,N_14212,N_14108);
xnor U14351 (N_14351,N_14242,N_14195);
xnor U14352 (N_14352,N_14184,N_14221);
nand U14353 (N_14353,N_14106,N_14215);
or U14354 (N_14354,N_14144,N_14236);
xnor U14355 (N_14355,N_14140,N_14238);
or U14356 (N_14356,N_14190,N_14118);
nor U14357 (N_14357,N_14144,N_14235);
or U14358 (N_14358,N_14116,N_14240);
nor U14359 (N_14359,N_14239,N_14220);
nand U14360 (N_14360,N_14226,N_14196);
xnor U14361 (N_14361,N_14213,N_14191);
xnor U14362 (N_14362,N_14186,N_14127);
nand U14363 (N_14363,N_14245,N_14109);
nand U14364 (N_14364,N_14104,N_14190);
xor U14365 (N_14365,N_14116,N_14162);
nor U14366 (N_14366,N_14223,N_14106);
and U14367 (N_14367,N_14149,N_14242);
nand U14368 (N_14368,N_14174,N_14143);
or U14369 (N_14369,N_14132,N_14120);
and U14370 (N_14370,N_14222,N_14155);
and U14371 (N_14371,N_14187,N_14108);
nor U14372 (N_14372,N_14102,N_14191);
nand U14373 (N_14373,N_14232,N_14130);
xor U14374 (N_14374,N_14229,N_14175);
and U14375 (N_14375,N_14244,N_14100);
xnor U14376 (N_14376,N_14103,N_14167);
nand U14377 (N_14377,N_14202,N_14180);
or U14378 (N_14378,N_14113,N_14245);
or U14379 (N_14379,N_14169,N_14231);
and U14380 (N_14380,N_14199,N_14148);
nand U14381 (N_14381,N_14176,N_14230);
and U14382 (N_14382,N_14120,N_14154);
and U14383 (N_14383,N_14168,N_14203);
or U14384 (N_14384,N_14163,N_14109);
or U14385 (N_14385,N_14203,N_14224);
nand U14386 (N_14386,N_14226,N_14167);
or U14387 (N_14387,N_14194,N_14136);
nand U14388 (N_14388,N_14226,N_14117);
nor U14389 (N_14389,N_14210,N_14132);
nand U14390 (N_14390,N_14198,N_14140);
nor U14391 (N_14391,N_14223,N_14111);
nand U14392 (N_14392,N_14143,N_14200);
and U14393 (N_14393,N_14197,N_14106);
or U14394 (N_14394,N_14211,N_14220);
nand U14395 (N_14395,N_14101,N_14190);
and U14396 (N_14396,N_14156,N_14141);
or U14397 (N_14397,N_14202,N_14172);
xnor U14398 (N_14398,N_14229,N_14135);
and U14399 (N_14399,N_14195,N_14227);
nor U14400 (N_14400,N_14318,N_14339);
xnor U14401 (N_14401,N_14277,N_14316);
or U14402 (N_14402,N_14335,N_14293);
nand U14403 (N_14403,N_14331,N_14366);
nor U14404 (N_14404,N_14269,N_14398);
nor U14405 (N_14405,N_14304,N_14354);
nor U14406 (N_14406,N_14343,N_14349);
xnor U14407 (N_14407,N_14399,N_14369);
nand U14408 (N_14408,N_14251,N_14279);
nor U14409 (N_14409,N_14393,N_14348);
xnor U14410 (N_14410,N_14288,N_14261);
nor U14411 (N_14411,N_14295,N_14376);
or U14412 (N_14412,N_14291,N_14365);
nand U14413 (N_14413,N_14262,N_14266);
nand U14414 (N_14414,N_14363,N_14297);
nor U14415 (N_14415,N_14308,N_14352);
xnor U14416 (N_14416,N_14258,N_14347);
and U14417 (N_14417,N_14270,N_14392);
or U14418 (N_14418,N_14358,N_14283);
nand U14419 (N_14419,N_14296,N_14282);
nand U14420 (N_14420,N_14368,N_14382);
and U14421 (N_14421,N_14355,N_14264);
and U14422 (N_14422,N_14325,N_14390);
nor U14423 (N_14423,N_14272,N_14311);
and U14424 (N_14424,N_14329,N_14298);
nand U14425 (N_14425,N_14252,N_14386);
xor U14426 (N_14426,N_14327,N_14273);
nand U14427 (N_14427,N_14315,N_14367);
xor U14428 (N_14428,N_14271,N_14359);
nand U14429 (N_14429,N_14377,N_14381);
or U14430 (N_14430,N_14306,N_14330);
nand U14431 (N_14431,N_14360,N_14340);
and U14432 (N_14432,N_14250,N_14286);
nand U14433 (N_14433,N_14259,N_14319);
xor U14434 (N_14434,N_14391,N_14371);
nor U14435 (N_14435,N_14389,N_14253);
nand U14436 (N_14436,N_14396,N_14289);
or U14437 (N_14437,N_14345,N_14361);
xnor U14438 (N_14438,N_14268,N_14254);
nand U14439 (N_14439,N_14388,N_14346);
nor U14440 (N_14440,N_14362,N_14353);
and U14441 (N_14441,N_14278,N_14385);
nand U14442 (N_14442,N_14350,N_14285);
nand U14443 (N_14443,N_14374,N_14314);
or U14444 (N_14444,N_14342,N_14256);
nand U14445 (N_14445,N_14263,N_14395);
or U14446 (N_14446,N_14265,N_14370);
xnor U14447 (N_14447,N_14372,N_14310);
nor U14448 (N_14448,N_14344,N_14292);
and U14449 (N_14449,N_14302,N_14380);
xnor U14450 (N_14450,N_14305,N_14307);
nand U14451 (N_14451,N_14300,N_14337);
and U14452 (N_14452,N_14280,N_14338);
xor U14453 (N_14453,N_14303,N_14284);
or U14454 (N_14454,N_14334,N_14317);
nand U14455 (N_14455,N_14379,N_14260);
nor U14456 (N_14456,N_14276,N_14373);
nand U14457 (N_14457,N_14320,N_14321);
nand U14458 (N_14458,N_14313,N_14332);
nor U14459 (N_14459,N_14322,N_14294);
nor U14460 (N_14460,N_14336,N_14274);
or U14461 (N_14461,N_14257,N_14255);
nor U14462 (N_14462,N_14312,N_14287);
nand U14463 (N_14463,N_14394,N_14387);
and U14464 (N_14464,N_14383,N_14323);
and U14465 (N_14465,N_14328,N_14299);
and U14466 (N_14466,N_14357,N_14378);
nor U14467 (N_14467,N_14384,N_14397);
nand U14468 (N_14468,N_14356,N_14309);
nor U14469 (N_14469,N_14364,N_14324);
nand U14470 (N_14470,N_14333,N_14281);
or U14471 (N_14471,N_14375,N_14326);
xnor U14472 (N_14472,N_14341,N_14275);
xnor U14473 (N_14473,N_14301,N_14267);
nor U14474 (N_14474,N_14290,N_14351);
or U14475 (N_14475,N_14361,N_14295);
and U14476 (N_14476,N_14313,N_14312);
nor U14477 (N_14477,N_14312,N_14382);
nor U14478 (N_14478,N_14346,N_14324);
nand U14479 (N_14479,N_14294,N_14395);
xnor U14480 (N_14480,N_14320,N_14344);
or U14481 (N_14481,N_14326,N_14302);
and U14482 (N_14482,N_14308,N_14270);
or U14483 (N_14483,N_14297,N_14379);
xnor U14484 (N_14484,N_14324,N_14258);
nor U14485 (N_14485,N_14298,N_14282);
nor U14486 (N_14486,N_14290,N_14295);
and U14487 (N_14487,N_14260,N_14316);
nor U14488 (N_14488,N_14312,N_14338);
and U14489 (N_14489,N_14392,N_14326);
nor U14490 (N_14490,N_14319,N_14372);
nor U14491 (N_14491,N_14267,N_14332);
nor U14492 (N_14492,N_14289,N_14306);
and U14493 (N_14493,N_14303,N_14263);
nor U14494 (N_14494,N_14345,N_14277);
xnor U14495 (N_14495,N_14254,N_14272);
and U14496 (N_14496,N_14340,N_14258);
nor U14497 (N_14497,N_14340,N_14316);
nor U14498 (N_14498,N_14280,N_14288);
nor U14499 (N_14499,N_14300,N_14281);
nor U14500 (N_14500,N_14307,N_14312);
or U14501 (N_14501,N_14370,N_14341);
xnor U14502 (N_14502,N_14342,N_14251);
nor U14503 (N_14503,N_14380,N_14317);
or U14504 (N_14504,N_14261,N_14302);
and U14505 (N_14505,N_14264,N_14289);
nor U14506 (N_14506,N_14363,N_14359);
xor U14507 (N_14507,N_14316,N_14305);
xnor U14508 (N_14508,N_14252,N_14316);
and U14509 (N_14509,N_14353,N_14332);
or U14510 (N_14510,N_14379,N_14323);
nand U14511 (N_14511,N_14391,N_14285);
or U14512 (N_14512,N_14390,N_14278);
nand U14513 (N_14513,N_14387,N_14318);
nand U14514 (N_14514,N_14335,N_14379);
and U14515 (N_14515,N_14348,N_14279);
nand U14516 (N_14516,N_14285,N_14293);
xor U14517 (N_14517,N_14283,N_14278);
nor U14518 (N_14518,N_14269,N_14356);
nor U14519 (N_14519,N_14306,N_14263);
and U14520 (N_14520,N_14364,N_14308);
xnor U14521 (N_14521,N_14260,N_14323);
nor U14522 (N_14522,N_14390,N_14351);
nor U14523 (N_14523,N_14352,N_14267);
and U14524 (N_14524,N_14356,N_14259);
nand U14525 (N_14525,N_14322,N_14360);
nor U14526 (N_14526,N_14250,N_14371);
or U14527 (N_14527,N_14373,N_14258);
and U14528 (N_14528,N_14352,N_14317);
and U14529 (N_14529,N_14349,N_14271);
nand U14530 (N_14530,N_14356,N_14335);
nor U14531 (N_14531,N_14349,N_14342);
nor U14532 (N_14532,N_14266,N_14376);
nor U14533 (N_14533,N_14368,N_14299);
nor U14534 (N_14534,N_14312,N_14347);
xor U14535 (N_14535,N_14382,N_14292);
nand U14536 (N_14536,N_14373,N_14333);
nand U14537 (N_14537,N_14283,N_14378);
or U14538 (N_14538,N_14380,N_14275);
and U14539 (N_14539,N_14282,N_14399);
nand U14540 (N_14540,N_14325,N_14286);
nand U14541 (N_14541,N_14378,N_14372);
xor U14542 (N_14542,N_14307,N_14376);
and U14543 (N_14543,N_14283,N_14319);
nor U14544 (N_14544,N_14252,N_14261);
nor U14545 (N_14545,N_14357,N_14345);
and U14546 (N_14546,N_14277,N_14342);
xor U14547 (N_14547,N_14339,N_14291);
xnor U14548 (N_14548,N_14391,N_14361);
or U14549 (N_14549,N_14303,N_14278);
and U14550 (N_14550,N_14527,N_14464);
nand U14551 (N_14551,N_14423,N_14543);
nand U14552 (N_14552,N_14403,N_14407);
nand U14553 (N_14553,N_14532,N_14467);
and U14554 (N_14554,N_14498,N_14444);
and U14555 (N_14555,N_14458,N_14411);
and U14556 (N_14556,N_14420,N_14495);
xor U14557 (N_14557,N_14529,N_14402);
nand U14558 (N_14558,N_14470,N_14507);
nor U14559 (N_14559,N_14435,N_14419);
and U14560 (N_14560,N_14413,N_14461);
and U14561 (N_14561,N_14491,N_14503);
or U14562 (N_14562,N_14446,N_14525);
and U14563 (N_14563,N_14449,N_14521);
nand U14564 (N_14564,N_14499,N_14434);
nand U14565 (N_14565,N_14482,N_14522);
and U14566 (N_14566,N_14416,N_14520);
nand U14567 (N_14567,N_14451,N_14511);
xor U14568 (N_14568,N_14481,N_14547);
or U14569 (N_14569,N_14439,N_14542);
nand U14570 (N_14570,N_14422,N_14426);
nor U14571 (N_14571,N_14436,N_14414);
or U14572 (N_14572,N_14489,N_14534);
and U14573 (N_14573,N_14438,N_14406);
nor U14574 (N_14574,N_14526,N_14490);
xor U14575 (N_14575,N_14493,N_14424);
or U14576 (N_14576,N_14538,N_14468);
and U14577 (N_14577,N_14508,N_14428);
nand U14578 (N_14578,N_14517,N_14408);
nor U14579 (N_14579,N_14431,N_14484);
xor U14580 (N_14580,N_14433,N_14533);
nand U14581 (N_14581,N_14471,N_14440);
nand U14582 (N_14582,N_14465,N_14475);
nand U14583 (N_14583,N_14514,N_14535);
xor U14584 (N_14584,N_14497,N_14457);
or U14585 (N_14585,N_14421,N_14501);
and U14586 (N_14586,N_14404,N_14415);
or U14587 (N_14587,N_14445,N_14405);
nand U14588 (N_14588,N_14456,N_14513);
and U14589 (N_14589,N_14429,N_14518);
nor U14590 (N_14590,N_14450,N_14430);
nor U14591 (N_14591,N_14479,N_14510);
or U14592 (N_14592,N_14473,N_14410);
nor U14593 (N_14593,N_14441,N_14487);
and U14594 (N_14594,N_14412,N_14537);
nor U14595 (N_14595,N_14469,N_14447);
xnor U14596 (N_14596,N_14541,N_14530);
or U14597 (N_14597,N_14540,N_14474);
xnor U14598 (N_14598,N_14528,N_14425);
and U14599 (N_14599,N_14427,N_14488);
nor U14600 (N_14600,N_14459,N_14486);
and U14601 (N_14601,N_14506,N_14515);
nand U14602 (N_14602,N_14509,N_14417);
nor U14603 (N_14603,N_14492,N_14442);
nand U14604 (N_14604,N_14483,N_14494);
nand U14605 (N_14605,N_14545,N_14505);
and U14606 (N_14606,N_14476,N_14460);
or U14607 (N_14607,N_14448,N_14466);
nand U14608 (N_14608,N_14549,N_14432);
xnor U14609 (N_14609,N_14546,N_14500);
or U14610 (N_14610,N_14531,N_14502);
and U14611 (N_14611,N_14400,N_14409);
and U14612 (N_14612,N_14480,N_14452);
and U14613 (N_14613,N_14443,N_14519);
nand U14614 (N_14614,N_14454,N_14496);
and U14615 (N_14615,N_14453,N_14544);
xor U14616 (N_14616,N_14504,N_14536);
and U14617 (N_14617,N_14524,N_14437);
nand U14618 (N_14618,N_14478,N_14523);
and U14619 (N_14619,N_14539,N_14516);
nor U14620 (N_14620,N_14463,N_14472);
or U14621 (N_14621,N_14477,N_14512);
and U14622 (N_14622,N_14548,N_14462);
nor U14623 (N_14623,N_14401,N_14455);
and U14624 (N_14624,N_14485,N_14418);
xnor U14625 (N_14625,N_14510,N_14419);
and U14626 (N_14626,N_14449,N_14422);
nand U14627 (N_14627,N_14460,N_14418);
nor U14628 (N_14628,N_14411,N_14532);
and U14629 (N_14629,N_14514,N_14479);
nor U14630 (N_14630,N_14419,N_14523);
and U14631 (N_14631,N_14498,N_14405);
or U14632 (N_14632,N_14492,N_14401);
nor U14633 (N_14633,N_14410,N_14511);
xnor U14634 (N_14634,N_14470,N_14441);
nor U14635 (N_14635,N_14466,N_14412);
xnor U14636 (N_14636,N_14424,N_14528);
nand U14637 (N_14637,N_14519,N_14522);
and U14638 (N_14638,N_14527,N_14524);
or U14639 (N_14639,N_14484,N_14442);
or U14640 (N_14640,N_14419,N_14471);
xor U14641 (N_14641,N_14490,N_14518);
or U14642 (N_14642,N_14427,N_14523);
nand U14643 (N_14643,N_14407,N_14415);
or U14644 (N_14644,N_14478,N_14426);
xor U14645 (N_14645,N_14543,N_14492);
or U14646 (N_14646,N_14479,N_14531);
xor U14647 (N_14647,N_14500,N_14474);
nor U14648 (N_14648,N_14426,N_14439);
and U14649 (N_14649,N_14444,N_14477);
and U14650 (N_14650,N_14431,N_14437);
nor U14651 (N_14651,N_14539,N_14444);
or U14652 (N_14652,N_14513,N_14408);
nand U14653 (N_14653,N_14481,N_14433);
nor U14654 (N_14654,N_14541,N_14400);
xnor U14655 (N_14655,N_14428,N_14501);
xnor U14656 (N_14656,N_14496,N_14462);
xor U14657 (N_14657,N_14473,N_14414);
xnor U14658 (N_14658,N_14443,N_14476);
xor U14659 (N_14659,N_14510,N_14436);
nand U14660 (N_14660,N_14519,N_14503);
nand U14661 (N_14661,N_14457,N_14483);
xor U14662 (N_14662,N_14461,N_14426);
and U14663 (N_14663,N_14515,N_14513);
and U14664 (N_14664,N_14517,N_14498);
and U14665 (N_14665,N_14510,N_14542);
and U14666 (N_14666,N_14440,N_14464);
nand U14667 (N_14667,N_14516,N_14493);
nand U14668 (N_14668,N_14478,N_14511);
xor U14669 (N_14669,N_14536,N_14547);
and U14670 (N_14670,N_14531,N_14525);
nand U14671 (N_14671,N_14459,N_14487);
nor U14672 (N_14672,N_14534,N_14434);
and U14673 (N_14673,N_14532,N_14524);
or U14674 (N_14674,N_14450,N_14407);
nor U14675 (N_14675,N_14525,N_14487);
nand U14676 (N_14676,N_14465,N_14488);
or U14677 (N_14677,N_14516,N_14416);
and U14678 (N_14678,N_14510,N_14408);
nand U14679 (N_14679,N_14416,N_14405);
or U14680 (N_14680,N_14532,N_14545);
nor U14681 (N_14681,N_14515,N_14457);
or U14682 (N_14682,N_14423,N_14417);
and U14683 (N_14683,N_14470,N_14460);
nor U14684 (N_14684,N_14408,N_14467);
or U14685 (N_14685,N_14468,N_14518);
xnor U14686 (N_14686,N_14478,N_14504);
nor U14687 (N_14687,N_14443,N_14459);
nand U14688 (N_14688,N_14510,N_14484);
nor U14689 (N_14689,N_14522,N_14520);
nor U14690 (N_14690,N_14542,N_14434);
nor U14691 (N_14691,N_14444,N_14443);
or U14692 (N_14692,N_14475,N_14493);
and U14693 (N_14693,N_14430,N_14463);
and U14694 (N_14694,N_14532,N_14517);
nor U14695 (N_14695,N_14527,N_14435);
nand U14696 (N_14696,N_14453,N_14435);
nor U14697 (N_14697,N_14406,N_14516);
nor U14698 (N_14698,N_14419,N_14423);
and U14699 (N_14699,N_14527,N_14417);
xor U14700 (N_14700,N_14692,N_14636);
xnor U14701 (N_14701,N_14656,N_14563);
or U14702 (N_14702,N_14651,N_14606);
nor U14703 (N_14703,N_14630,N_14689);
xor U14704 (N_14704,N_14690,N_14647);
nor U14705 (N_14705,N_14620,N_14586);
or U14706 (N_14706,N_14675,N_14592);
or U14707 (N_14707,N_14614,N_14595);
nor U14708 (N_14708,N_14652,N_14635);
nor U14709 (N_14709,N_14590,N_14684);
nor U14710 (N_14710,N_14555,N_14599);
nand U14711 (N_14711,N_14655,N_14583);
nor U14712 (N_14712,N_14609,N_14696);
or U14713 (N_14713,N_14639,N_14564);
nor U14714 (N_14714,N_14676,N_14648);
and U14715 (N_14715,N_14669,N_14560);
or U14716 (N_14716,N_14670,N_14685);
or U14717 (N_14717,N_14673,N_14566);
xor U14718 (N_14718,N_14662,N_14587);
xor U14719 (N_14719,N_14626,N_14672);
nor U14720 (N_14720,N_14633,N_14578);
or U14721 (N_14721,N_14604,N_14551);
nor U14722 (N_14722,N_14621,N_14624);
or U14723 (N_14723,N_14550,N_14686);
xnor U14724 (N_14724,N_14661,N_14631);
or U14725 (N_14725,N_14569,N_14645);
nor U14726 (N_14726,N_14638,N_14580);
or U14727 (N_14727,N_14622,N_14605);
or U14728 (N_14728,N_14571,N_14602);
or U14729 (N_14729,N_14699,N_14570);
nor U14730 (N_14730,N_14657,N_14559);
and U14731 (N_14731,N_14557,N_14629);
nand U14732 (N_14732,N_14634,N_14577);
or U14733 (N_14733,N_14597,N_14610);
xnor U14734 (N_14734,N_14591,N_14553);
or U14735 (N_14735,N_14565,N_14572);
and U14736 (N_14736,N_14653,N_14691);
xor U14737 (N_14737,N_14646,N_14666);
nor U14738 (N_14738,N_14660,N_14593);
nand U14739 (N_14739,N_14693,N_14596);
nand U14740 (N_14740,N_14678,N_14619);
nor U14741 (N_14741,N_14695,N_14556);
nor U14742 (N_14742,N_14637,N_14658);
nand U14743 (N_14743,N_14698,N_14640);
nand U14744 (N_14744,N_14679,N_14567);
nand U14745 (N_14745,N_14663,N_14674);
or U14746 (N_14746,N_14584,N_14601);
nand U14747 (N_14747,N_14642,N_14554);
nand U14748 (N_14748,N_14562,N_14576);
nand U14749 (N_14749,N_14668,N_14568);
or U14750 (N_14750,N_14628,N_14574);
nand U14751 (N_14751,N_14649,N_14575);
or U14752 (N_14752,N_14598,N_14694);
nor U14753 (N_14753,N_14594,N_14659);
nor U14754 (N_14754,N_14615,N_14600);
nor U14755 (N_14755,N_14680,N_14664);
nand U14756 (N_14756,N_14603,N_14681);
xnor U14757 (N_14757,N_14650,N_14611);
nor U14758 (N_14758,N_14618,N_14697);
and U14759 (N_14759,N_14608,N_14607);
and U14760 (N_14760,N_14589,N_14613);
or U14761 (N_14761,N_14644,N_14561);
nand U14762 (N_14762,N_14641,N_14582);
nand U14763 (N_14763,N_14558,N_14617);
and U14764 (N_14764,N_14677,N_14667);
or U14765 (N_14765,N_14573,N_14627);
nor U14766 (N_14766,N_14688,N_14552);
and U14767 (N_14767,N_14654,N_14625);
nand U14768 (N_14768,N_14612,N_14623);
nand U14769 (N_14769,N_14687,N_14588);
or U14770 (N_14770,N_14581,N_14632);
or U14771 (N_14771,N_14616,N_14682);
nand U14772 (N_14772,N_14665,N_14579);
or U14773 (N_14773,N_14671,N_14683);
or U14774 (N_14774,N_14585,N_14643);
and U14775 (N_14775,N_14590,N_14668);
nor U14776 (N_14776,N_14657,N_14651);
nand U14777 (N_14777,N_14685,N_14671);
or U14778 (N_14778,N_14628,N_14681);
nand U14779 (N_14779,N_14621,N_14668);
or U14780 (N_14780,N_14586,N_14654);
and U14781 (N_14781,N_14677,N_14568);
and U14782 (N_14782,N_14592,N_14582);
nor U14783 (N_14783,N_14626,N_14656);
and U14784 (N_14784,N_14611,N_14581);
xnor U14785 (N_14785,N_14621,N_14647);
nand U14786 (N_14786,N_14617,N_14614);
and U14787 (N_14787,N_14622,N_14563);
or U14788 (N_14788,N_14676,N_14678);
and U14789 (N_14789,N_14634,N_14586);
or U14790 (N_14790,N_14566,N_14602);
xnor U14791 (N_14791,N_14598,N_14585);
nand U14792 (N_14792,N_14689,N_14569);
xnor U14793 (N_14793,N_14579,N_14610);
nand U14794 (N_14794,N_14673,N_14650);
nand U14795 (N_14795,N_14683,N_14607);
and U14796 (N_14796,N_14652,N_14677);
or U14797 (N_14797,N_14623,N_14698);
nor U14798 (N_14798,N_14675,N_14679);
nand U14799 (N_14799,N_14591,N_14613);
and U14800 (N_14800,N_14611,N_14653);
xor U14801 (N_14801,N_14566,N_14563);
xnor U14802 (N_14802,N_14642,N_14690);
nand U14803 (N_14803,N_14595,N_14641);
nor U14804 (N_14804,N_14650,N_14612);
nand U14805 (N_14805,N_14611,N_14555);
xor U14806 (N_14806,N_14610,N_14584);
nand U14807 (N_14807,N_14664,N_14563);
or U14808 (N_14808,N_14675,N_14677);
or U14809 (N_14809,N_14607,N_14670);
and U14810 (N_14810,N_14608,N_14582);
and U14811 (N_14811,N_14568,N_14690);
and U14812 (N_14812,N_14553,N_14697);
xnor U14813 (N_14813,N_14698,N_14625);
and U14814 (N_14814,N_14605,N_14632);
or U14815 (N_14815,N_14667,N_14600);
nand U14816 (N_14816,N_14680,N_14585);
nand U14817 (N_14817,N_14583,N_14612);
nand U14818 (N_14818,N_14658,N_14639);
and U14819 (N_14819,N_14666,N_14571);
nor U14820 (N_14820,N_14622,N_14618);
nor U14821 (N_14821,N_14655,N_14584);
or U14822 (N_14822,N_14610,N_14573);
nor U14823 (N_14823,N_14631,N_14636);
nor U14824 (N_14824,N_14669,N_14642);
or U14825 (N_14825,N_14601,N_14565);
nor U14826 (N_14826,N_14602,N_14697);
nand U14827 (N_14827,N_14673,N_14631);
xor U14828 (N_14828,N_14668,N_14644);
nand U14829 (N_14829,N_14649,N_14592);
and U14830 (N_14830,N_14688,N_14682);
nor U14831 (N_14831,N_14607,N_14669);
nand U14832 (N_14832,N_14666,N_14628);
or U14833 (N_14833,N_14565,N_14608);
or U14834 (N_14834,N_14694,N_14660);
nor U14835 (N_14835,N_14606,N_14621);
nor U14836 (N_14836,N_14581,N_14692);
nor U14837 (N_14837,N_14676,N_14617);
nor U14838 (N_14838,N_14663,N_14672);
nor U14839 (N_14839,N_14691,N_14619);
or U14840 (N_14840,N_14591,N_14569);
and U14841 (N_14841,N_14624,N_14686);
nor U14842 (N_14842,N_14639,N_14699);
or U14843 (N_14843,N_14619,N_14611);
or U14844 (N_14844,N_14677,N_14607);
xor U14845 (N_14845,N_14565,N_14590);
nand U14846 (N_14846,N_14582,N_14568);
and U14847 (N_14847,N_14584,N_14676);
xnor U14848 (N_14848,N_14564,N_14698);
or U14849 (N_14849,N_14583,N_14673);
and U14850 (N_14850,N_14778,N_14818);
nor U14851 (N_14851,N_14805,N_14765);
or U14852 (N_14852,N_14844,N_14722);
xnor U14853 (N_14853,N_14766,N_14812);
nor U14854 (N_14854,N_14709,N_14758);
nor U14855 (N_14855,N_14828,N_14751);
or U14856 (N_14856,N_14799,N_14845);
and U14857 (N_14857,N_14727,N_14721);
or U14858 (N_14858,N_14729,N_14769);
and U14859 (N_14859,N_14759,N_14777);
nand U14860 (N_14860,N_14724,N_14717);
nor U14861 (N_14861,N_14723,N_14795);
nor U14862 (N_14862,N_14782,N_14757);
xnor U14863 (N_14863,N_14787,N_14710);
nand U14864 (N_14864,N_14746,N_14817);
and U14865 (N_14865,N_14848,N_14772);
nand U14866 (N_14866,N_14798,N_14832);
nand U14867 (N_14867,N_14701,N_14781);
nor U14868 (N_14868,N_14792,N_14733);
or U14869 (N_14869,N_14768,N_14770);
or U14870 (N_14870,N_14815,N_14809);
xor U14871 (N_14871,N_14725,N_14750);
or U14872 (N_14872,N_14707,N_14700);
or U14873 (N_14873,N_14788,N_14703);
xor U14874 (N_14874,N_14748,N_14706);
xnor U14875 (N_14875,N_14806,N_14827);
and U14876 (N_14876,N_14735,N_14771);
or U14877 (N_14877,N_14780,N_14764);
or U14878 (N_14878,N_14839,N_14720);
nor U14879 (N_14879,N_14824,N_14836);
and U14880 (N_14880,N_14820,N_14800);
nand U14881 (N_14881,N_14785,N_14761);
or U14882 (N_14882,N_14776,N_14767);
or U14883 (N_14883,N_14745,N_14754);
or U14884 (N_14884,N_14741,N_14756);
or U14885 (N_14885,N_14846,N_14714);
or U14886 (N_14886,N_14779,N_14813);
xor U14887 (N_14887,N_14775,N_14712);
nor U14888 (N_14888,N_14796,N_14837);
nand U14889 (N_14889,N_14830,N_14802);
and U14890 (N_14890,N_14705,N_14713);
and U14891 (N_14891,N_14840,N_14842);
and U14892 (N_14892,N_14719,N_14791);
nor U14893 (N_14893,N_14834,N_14801);
xor U14894 (N_14894,N_14718,N_14816);
xor U14895 (N_14895,N_14739,N_14755);
nand U14896 (N_14896,N_14743,N_14753);
nand U14897 (N_14897,N_14808,N_14794);
nand U14898 (N_14898,N_14797,N_14737);
or U14899 (N_14899,N_14742,N_14807);
nor U14900 (N_14900,N_14752,N_14841);
nor U14901 (N_14901,N_14822,N_14826);
nor U14902 (N_14902,N_14784,N_14793);
or U14903 (N_14903,N_14702,N_14789);
nand U14904 (N_14904,N_14773,N_14716);
nand U14905 (N_14905,N_14740,N_14849);
xor U14906 (N_14906,N_14762,N_14715);
xnor U14907 (N_14907,N_14749,N_14708);
and U14908 (N_14908,N_14704,N_14732);
or U14909 (N_14909,N_14760,N_14843);
or U14910 (N_14910,N_14783,N_14811);
and U14911 (N_14911,N_14825,N_14790);
nand U14912 (N_14912,N_14711,N_14747);
or U14913 (N_14913,N_14786,N_14814);
and U14914 (N_14914,N_14831,N_14738);
nor U14915 (N_14915,N_14847,N_14821);
and U14916 (N_14916,N_14731,N_14819);
nand U14917 (N_14917,N_14726,N_14810);
nor U14918 (N_14918,N_14736,N_14803);
or U14919 (N_14919,N_14763,N_14804);
nand U14920 (N_14920,N_14829,N_14734);
xnor U14921 (N_14921,N_14835,N_14728);
xor U14922 (N_14922,N_14730,N_14744);
nor U14923 (N_14923,N_14833,N_14838);
and U14924 (N_14924,N_14823,N_14774);
nor U14925 (N_14925,N_14801,N_14798);
and U14926 (N_14926,N_14741,N_14766);
nor U14927 (N_14927,N_14833,N_14706);
nor U14928 (N_14928,N_14737,N_14785);
nand U14929 (N_14929,N_14736,N_14818);
nor U14930 (N_14930,N_14820,N_14798);
nand U14931 (N_14931,N_14849,N_14832);
and U14932 (N_14932,N_14744,N_14716);
and U14933 (N_14933,N_14702,N_14710);
xor U14934 (N_14934,N_14823,N_14772);
nor U14935 (N_14935,N_14801,N_14780);
nand U14936 (N_14936,N_14806,N_14740);
and U14937 (N_14937,N_14791,N_14805);
xor U14938 (N_14938,N_14824,N_14718);
or U14939 (N_14939,N_14796,N_14700);
or U14940 (N_14940,N_14782,N_14833);
and U14941 (N_14941,N_14724,N_14825);
nand U14942 (N_14942,N_14750,N_14783);
nor U14943 (N_14943,N_14791,N_14796);
xor U14944 (N_14944,N_14743,N_14817);
and U14945 (N_14945,N_14797,N_14744);
nor U14946 (N_14946,N_14771,N_14772);
nor U14947 (N_14947,N_14827,N_14812);
or U14948 (N_14948,N_14833,N_14725);
or U14949 (N_14949,N_14818,N_14806);
nor U14950 (N_14950,N_14720,N_14803);
and U14951 (N_14951,N_14761,N_14843);
or U14952 (N_14952,N_14770,N_14796);
and U14953 (N_14953,N_14819,N_14765);
nand U14954 (N_14954,N_14795,N_14799);
xnor U14955 (N_14955,N_14761,N_14717);
xnor U14956 (N_14956,N_14758,N_14777);
xor U14957 (N_14957,N_14775,N_14737);
or U14958 (N_14958,N_14742,N_14810);
nand U14959 (N_14959,N_14833,N_14827);
xnor U14960 (N_14960,N_14818,N_14823);
and U14961 (N_14961,N_14769,N_14814);
or U14962 (N_14962,N_14799,N_14826);
nand U14963 (N_14963,N_14707,N_14825);
and U14964 (N_14964,N_14733,N_14757);
xor U14965 (N_14965,N_14778,N_14807);
nor U14966 (N_14966,N_14736,N_14801);
or U14967 (N_14967,N_14750,N_14702);
nor U14968 (N_14968,N_14757,N_14822);
nor U14969 (N_14969,N_14831,N_14796);
nor U14970 (N_14970,N_14739,N_14710);
xnor U14971 (N_14971,N_14725,N_14708);
or U14972 (N_14972,N_14774,N_14713);
nand U14973 (N_14973,N_14706,N_14767);
xnor U14974 (N_14974,N_14712,N_14818);
nor U14975 (N_14975,N_14759,N_14752);
and U14976 (N_14976,N_14818,N_14700);
xnor U14977 (N_14977,N_14844,N_14813);
or U14978 (N_14978,N_14763,N_14806);
nand U14979 (N_14979,N_14827,N_14746);
nor U14980 (N_14980,N_14713,N_14814);
xor U14981 (N_14981,N_14742,N_14736);
or U14982 (N_14982,N_14841,N_14825);
nand U14983 (N_14983,N_14722,N_14834);
xnor U14984 (N_14984,N_14786,N_14822);
xnor U14985 (N_14985,N_14810,N_14750);
nand U14986 (N_14986,N_14748,N_14725);
nand U14987 (N_14987,N_14810,N_14712);
or U14988 (N_14988,N_14744,N_14833);
nand U14989 (N_14989,N_14701,N_14831);
or U14990 (N_14990,N_14741,N_14733);
or U14991 (N_14991,N_14795,N_14801);
and U14992 (N_14992,N_14714,N_14820);
or U14993 (N_14993,N_14755,N_14808);
nor U14994 (N_14994,N_14718,N_14828);
xnor U14995 (N_14995,N_14782,N_14718);
xnor U14996 (N_14996,N_14786,N_14741);
nor U14997 (N_14997,N_14799,N_14779);
nor U14998 (N_14998,N_14702,N_14833);
nand U14999 (N_14999,N_14791,N_14708);
nand UO_0 (O_0,N_14887,N_14918);
nor UO_1 (O_1,N_14881,N_14922);
and UO_2 (O_2,N_14997,N_14920);
or UO_3 (O_3,N_14977,N_14921);
or UO_4 (O_4,N_14933,N_14851);
and UO_5 (O_5,N_14855,N_14987);
nor UO_6 (O_6,N_14992,N_14939);
nor UO_7 (O_7,N_14882,N_14972);
xnor UO_8 (O_8,N_14923,N_14935);
and UO_9 (O_9,N_14989,N_14946);
and UO_10 (O_10,N_14995,N_14870);
nor UO_11 (O_11,N_14911,N_14890);
xnor UO_12 (O_12,N_14862,N_14913);
xnor UO_13 (O_13,N_14871,N_14938);
nor UO_14 (O_14,N_14856,N_14970);
nand UO_15 (O_15,N_14934,N_14858);
and UO_16 (O_16,N_14969,N_14941);
nor UO_17 (O_17,N_14879,N_14967);
nand UO_18 (O_18,N_14964,N_14877);
and UO_19 (O_19,N_14876,N_14948);
and UO_20 (O_20,N_14963,N_14954);
xor UO_21 (O_21,N_14873,N_14901);
nand UO_22 (O_22,N_14960,N_14884);
and UO_23 (O_23,N_14945,N_14949);
nand UO_24 (O_24,N_14915,N_14943);
nand UO_25 (O_25,N_14864,N_14908);
xnor UO_26 (O_26,N_14958,N_14947);
and UO_27 (O_27,N_14962,N_14898);
nor UO_28 (O_28,N_14975,N_14981);
nand UO_29 (O_29,N_14937,N_14905);
or UO_30 (O_30,N_14883,N_14936);
nor UO_31 (O_31,N_14988,N_14929);
nor UO_32 (O_32,N_14925,N_14978);
and UO_33 (O_33,N_14854,N_14968);
nand UO_34 (O_34,N_14897,N_14903);
nor UO_35 (O_35,N_14872,N_14880);
xnor UO_36 (O_36,N_14912,N_14896);
xor UO_37 (O_37,N_14961,N_14924);
nor UO_38 (O_38,N_14886,N_14926);
xnor UO_39 (O_39,N_14953,N_14983);
and UO_40 (O_40,N_14867,N_14956);
and UO_41 (O_41,N_14917,N_14971);
xnor UO_42 (O_42,N_14850,N_14966);
nand UO_43 (O_43,N_14885,N_14861);
nand UO_44 (O_44,N_14865,N_14944);
nor UO_45 (O_45,N_14916,N_14927);
xor UO_46 (O_46,N_14931,N_14952);
nor UO_47 (O_47,N_14857,N_14999);
and UO_48 (O_48,N_14930,N_14899);
or UO_49 (O_49,N_14904,N_14998);
xnor UO_50 (O_50,N_14979,N_14852);
xnor UO_51 (O_51,N_14888,N_14902);
or UO_52 (O_52,N_14914,N_14973);
xnor UO_53 (O_53,N_14928,N_14900);
nand UO_54 (O_54,N_14996,N_14940);
and UO_55 (O_55,N_14906,N_14957);
or UO_56 (O_56,N_14932,N_14907);
and UO_57 (O_57,N_14869,N_14909);
nor UO_58 (O_58,N_14891,N_14874);
nor UO_59 (O_59,N_14853,N_14984);
or UO_60 (O_60,N_14919,N_14955);
nand UO_61 (O_61,N_14878,N_14974);
or UO_62 (O_62,N_14950,N_14863);
or UO_63 (O_63,N_14895,N_14951);
nor UO_64 (O_64,N_14976,N_14875);
xor UO_65 (O_65,N_14982,N_14866);
nor UO_66 (O_66,N_14859,N_14892);
nand UO_67 (O_67,N_14910,N_14985);
xor UO_68 (O_68,N_14894,N_14994);
nor UO_69 (O_69,N_14991,N_14990);
and UO_70 (O_70,N_14860,N_14893);
or UO_71 (O_71,N_14986,N_14965);
xor UO_72 (O_72,N_14868,N_14980);
xor UO_73 (O_73,N_14959,N_14942);
or UO_74 (O_74,N_14993,N_14889);
nand UO_75 (O_75,N_14962,N_14881);
nor UO_76 (O_76,N_14914,N_14923);
nand UO_77 (O_77,N_14995,N_14898);
and UO_78 (O_78,N_14969,N_14982);
xnor UO_79 (O_79,N_14888,N_14862);
nor UO_80 (O_80,N_14952,N_14883);
nand UO_81 (O_81,N_14899,N_14994);
nand UO_82 (O_82,N_14944,N_14973);
and UO_83 (O_83,N_14856,N_14967);
and UO_84 (O_84,N_14863,N_14962);
xnor UO_85 (O_85,N_14994,N_14949);
nand UO_86 (O_86,N_14903,N_14871);
xor UO_87 (O_87,N_14864,N_14888);
xnor UO_88 (O_88,N_14918,N_14892);
nor UO_89 (O_89,N_14947,N_14975);
nand UO_90 (O_90,N_14927,N_14982);
xor UO_91 (O_91,N_14889,N_14979);
and UO_92 (O_92,N_14887,N_14976);
nand UO_93 (O_93,N_14927,N_14943);
or UO_94 (O_94,N_14891,N_14865);
nand UO_95 (O_95,N_14859,N_14912);
xor UO_96 (O_96,N_14916,N_14992);
nand UO_97 (O_97,N_14956,N_14894);
or UO_98 (O_98,N_14927,N_14999);
xor UO_99 (O_99,N_14940,N_14947);
or UO_100 (O_100,N_14984,N_14874);
nand UO_101 (O_101,N_14954,N_14865);
nand UO_102 (O_102,N_14855,N_14942);
xor UO_103 (O_103,N_14938,N_14939);
and UO_104 (O_104,N_14908,N_14981);
nand UO_105 (O_105,N_14919,N_14903);
xnor UO_106 (O_106,N_14981,N_14921);
nor UO_107 (O_107,N_14949,N_14893);
xor UO_108 (O_108,N_14898,N_14940);
nand UO_109 (O_109,N_14961,N_14962);
xor UO_110 (O_110,N_14938,N_14964);
nor UO_111 (O_111,N_14935,N_14928);
xnor UO_112 (O_112,N_14916,N_14974);
xor UO_113 (O_113,N_14931,N_14875);
and UO_114 (O_114,N_14867,N_14904);
or UO_115 (O_115,N_14860,N_14901);
and UO_116 (O_116,N_14858,N_14885);
or UO_117 (O_117,N_14897,N_14951);
or UO_118 (O_118,N_14983,N_14907);
or UO_119 (O_119,N_14936,N_14929);
or UO_120 (O_120,N_14975,N_14872);
xnor UO_121 (O_121,N_14949,N_14886);
or UO_122 (O_122,N_14967,N_14890);
nand UO_123 (O_123,N_14864,N_14925);
or UO_124 (O_124,N_14995,N_14864);
and UO_125 (O_125,N_14902,N_14885);
and UO_126 (O_126,N_14933,N_14913);
nor UO_127 (O_127,N_14916,N_14874);
xnor UO_128 (O_128,N_14888,N_14996);
and UO_129 (O_129,N_14866,N_14908);
nand UO_130 (O_130,N_14961,N_14950);
xor UO_131 (O_131,N_14877,N_14875);
or UO_132 (O_132,N_14856,N_14966);
and UO_133 (O_133,N_14927,N_14884);
or UO_134 (O_134,N_14992,N_14921);
nor UO_135 (O_135,N_14893,N_14885);
and UO_136 (O_136,N_14999,N_14856);
and UO_137 (O_137,N_14941,N_14869);
or UO_138 (O_138,N_14880,N_14960);
and UO_139 (O_139,N_14856,N_14881);
and UO_140 (O_140,N_14945,N_14980);
xor UO_141 (O_141,N_14887,N_14952);
and UO_142 (O_142,N_14963,N_14855);
nor UO_143 (O_143,N_14970,N_14925);
nand UO_144 (O_144,N_14872,N_14963);
or UO_145 (O_145,N_14998,N_14975);
and UO_146 (O_146,N_14881,N_14958);
nor UO_147 (O_147,N_14868,N_14969);
nand UO_148 (O_148,N_14940,N_14914);
nand UO_149 (O_149,N_14989,N_14964);
nor UO_150 (O_150,N_14910,N_14880);
xnor UO_151 (O_151,N_14886,N_14923);
or UO_152 (O_152,N_14939,N_14909);
nor UO_153 (O_153,N_14948,N_14886);
and UO_154 (O_154,N_14869,N_14961);
xor UO_155 (O_155,N_14980,N_14906);
nor UO_156 (O_156,N_14879,N_14870);
nand UO_157 (O_157,N_14983,N_14873);
xnor UO_158 (O_158,N_14898,N_14996);
xor UO_159 (O_159,N_14921,N_14938);
and UO_160 (O_160,N_14879,N_14928);
or UO_161 (O_161,N_14922,N_14953);
nand UO_162 (O_162,N_14893,N_14912);
nand UO_163 (O_163,N_14946,N_14952);
xor UO_164 (O_164,N_14864,N_14865);
and UO_165 (O_165,N_14972,N_14949);
and UO_166 (O_166,N_14860,N_14858);
or UO_167 (O_167,N_14872,N_14939);
nor UO_168 (O_168,N_14881,N_14985);
or UO_169 (O_169,N_14901,N_14992);
xor UO_170 (O_170,N_14967,N_14870);
nor UO_171 (O_171,N_14860,N_14934);
nor UO_172 (O_172,N_14928,N_14961);
and UO_173 (O_173,N_14984,N_14878);
nor UO_174 (O_174,N_14970,N_14966);
xor UO_175 (O_175,N_14879,N_14980);
or UO_176 (O_176,N_14875,N_14885);
xor UO_177 (O_177,N_14929,N_14966);
and UO_178 (O_178,N_14981,N_14888);
or UO_179 (O_179,N_14946,N_14975);
xor UO_180 (O_180,N_14896,N_14857);
xnor UO_181 (O_181,N_14953,N_14867);
or UO_182 (O_182,N_14868,N_14924);
nor UO_183 (O_183,N_14904,N_14978);
xor UO_184 (O_184,N_14972,N_14915);
xor UO_185 (O_185,N_14919,N_14884);
nand UO_186 (O_186,N_14925,N_14984);
nand UO_187 (O_187,N_14910,N_14867);
or UO_188 (O_188,N_14909,N_14882);
nor UO_189 (O_189,N_14941,N_14989);
and UO_190 (O_190,N_14907,N_14959);
nand UO_191 (O_191,N_14976,N_14940);
and UO_192 (O_192,N_14924,N_14864);
nor UO_193 (O_193,N_14871,N_14875);
and UO_194 (O_194,N_14889,N_14963);
nand UO_195 (O_195,N_14873,N_14874);
nor UO_196 (O_196,N_14891,N_14901);
nand UO_197 (O_197,N_14878,N_14967);
or UO_198 (O_198,N_14933,N_14914);
or UO_199 (O_199,N_14958,N_14898);
nor UO_200 (O_200,N_14907,N_14955);
nand UO_201 (O_201,N_14970,N_14999);
and UO_202 (O_202,N_14863,N_14956);
xnor UO_203 (O_203,N_14884,N_14877);
xor UO_204 (O_204,N_14899,N_14912);
and UO_205 (O_205,N_14919,N_14926);
and UO_206 (O_206,N_14883,N_14953);
nand UO_207 (O_207,N_14993,N_14955);
or UO_208 (O_208,N_14994,N_14920);
or UO_209 (O_209,N_14967,N_14895);
nand UO_210 (O_210,N_14919,N_14895);
or UO_211 (O_211,N_14907,N_14938);
and UO_212 (O_212,N_14961,N_14876);
nor UO_213 (O_213,N_14998,N_14881);
or UO_214 (O_214,N_14934,N_14878);
nand UO_215 (O_215,N_14988,N_14935);
and UO_216 (O_216,N_14989,N_14982);
xor UO_217 (O_217,N_14897,N_14954);
xor UO_218 (O_218,N_14882,N_14991);
nor UO_219 (O_219,N_14960,N_14990);
nor UO_220 (O_220,N_14882,N_14956);
nor UO_221 (O_221,N_14989,N_14882);
and UO_222 (O_222,N_14971,N_14865);
xor UO_223 (O_223,N_14944,N_14956);
nor UO_224 (O_224,N_14936,N_14873);
nand UO_225 (O_225,N_14956,N_14959);
nor UO_226 (O_226,N_14983,N_14918);
or UO_227 (O_227,N_14939,N_14994);
nand UO_228 (O_228,N_14895,N_14924);
nor UO_229 (O_229,N_14928,N_14922);
nor UO_230 (O_230,N_14931,N_14941);
xnor UO_231 (O_231,N_14903,N_14937);
nor UO_232 (O_232,N_14868,N_14855);
and UO_233 (O_233,N_14954,N_14982);
or UO_234 (O_234,N_14866,N_14974);
nand UO_235 (O_235,N_14895,N_14891);
nor UO_236 (O_236,N_14917,N_14897);
nand UO_237 (O_237,N_14940,N_14939);
or UO_238 (O_238,N_14944,N_14891);
and UO_239 (O_239,N_14904,N_14875);
nor UO_240 (O_240,N_14983,N_14904);
nor UO_241 (O_241,N_14981,N_14852);
nor UO_242 (O_242,N_14854,N_14919);
nand UO_243 (O_243,N_14881,N_14863);
and UO_244 (O_244,N_14864,N_14980);
nand UO_245 (O_245,N_14901,N_14881);
nor UO_246 (O_246,N_14974,N_14990);
nor UO_247 (O_247,N_14981,N_14879);
xnor UO_248 (O_248,N_14916,N_14884);
or UO_249 (O_249,N_14854,N_14965);
nand UO_250 (O_250,N_14960,N_14996);
and UO_251 (O_251,N_14948,N_14951);
or UO_252 (O_252,N_14928,N_14987);
or UO_253 (O_253,N_14958,N_14922);
or UO_254 (O_254,N_14937,N_14971);
or UO_255 (O_255,N_14984,N_14913);
xor UO_256 (O_256,N_14872,N_14991);
or UO_257 (O_257,N_14948,N_14980);
xnor UO_258 (O_258,N_14934,N_14871);
nand UO_259 (O_259,N_14911,N_14874);
or UO_260 (O_260,N_14942,N_14990);
or UO_261 (O_261,N_14930,N_14933);
nand UO_262 (O_262,N_14924,N_14876);
nand UO_263 (O_263,N_14901,N_14954);
nand UO_264 (O_264,N_14933,N_14890);
and UO_265 (O_265,N_14903,N_14970);
and UO_266 (O_266,N_14904,N_14873);
nor UO_267 (O_267,N_14914,N_14970);
xnor UO_268 (O_268,N_14924,N_14877);
and UO_269 (O_269,N_14882,N_14858);
and UO_270 (O_270,N_14934,N_14954);
nand UO_271 (O_271,N_14932,N_14997);
nand UO_272 (O_272,N_14901,N_14914);
nand UO_273 (O_273,N_14985,N_14957);
and UO_274 (O_274,N_14996,N_14961);
xnor UO_275 (O_275,N_14877,N_14894);
nor UO_276 (O_276,N_14964,N_14997);
nand UO_277 (O_277,N_14970,N_14992);
and UO_278 (O_278,N_14856,N_14909);
xnor UO_279 (O_279,N_14996,N_14976);
nor UO_280 (O_280,N_14876,N_14960);
xor UO_281 (O_281,N_14992,N_14954);
xor UO_282 (O_282,N_14870,N_14983);
nor UO_283 (O_283,N_14937,N_14922);
xnor UO_284 (O_284,N_14935,N_14974);
nor UO_285 (O_285,N_14874,N_14986);
nor UO_286 (O_286,N_14912,N_14906);
nor UO_287 (O_287,N_14998,N_14860);
nor UO_288 (O_288,N_14962,N_14868);
or UO_289 (O_289,N_14963,N_14875);
nor UO_290 (O_290,N_14929,N_14851);
nor UO_291 (O_291,N_14865,N_14884);
nor UO_292 (O_292,N_14973,N_14903);
xnor UO_293 (O_293,N_14998,N_14944);
or UO_294 (O_294,N_14980,N_14923);
nor UO_295 (O_295,N_14937,N_14921);
xor UO_296 (O_296,N_14889,N_14953);
nor UO_297 (O_297,N_14876,N_14908);
and UO_298 (O_298,N_14947,N_14955);
and UO_299 (O_299,N_14956,N_14910);
and UO_300 (O_300,N_14859,N_14862);
and UO_301 (O_301,N_14926,N_14897);
nand UO_302 (O_302,N_14964,N_14980);
or UO_303 (O_303,N_14891,N_14993);
or UO_304 (O_304,N_14978,N_14932);
nor UO_305 (O_305,N_14876,N_14885);
xnor UO_306 (O_306,N_14868,N_14871);
or UO_307 (O_307,N_14902,N_14944);
nand UO_308 (O_308,N_14916,N_14870);
and UO_309 (O_309,N_14865,N_14873);
nand UO_310 (O_310,N_14999,N_14933);
nand UO_311 (O_311,N_14973,N_14984);
xor UO_312 (O_312,N_14853,N_14938);
and UO_313 (O_313,N_14877,N_14958);
nor UO_314 (O_314,N_14918,N_14958);
xor UO_315 (O_315,N_14940,N_14994);
nor UO_316 (O_316,N_14924,N_14972);
xor UO_317 (O_317,N_14968,N_14919);
and UO_318 (O_318,N_14908,N_14942);
or UO_319 (O_319,N_14907,N_14953);
nand UO_320 (O_320,N_14961,N_14972);
xor UO_321 (O_321,N_14957,N_14967);
and UO_322 (O_322,N_14912,N_14853);
and UO_323 (O_323,N_14898,N_14997);
nor UO_324 (O_324,N_14953,N_14862);
nand UO_325 (O_325,N_14993,N_14971);
nand UO_326 (O_326,N_14915,N_14927);
and UO_327 (O_327,N_14936,N_14890);
or UO_328 (O_328,N_14861,N_14991);
nand UO_329 (O_329,N_14936,N_14927);
nand UO_330 (O_330,N_14855,N_14918);
nand UO_331 (O_331,N_14857,N_14870);
xnor UO_332 (O_332,N_14908,N_14899);
nand UO_333 (O_333,N_14856,N_14875);
nor UO_334 (O_334,N_14943,N_14850);
xor UO_335 (O_335,N_14937,N_14958);
nand UO_336 (O_336,N_14852,N_14905);
nor UO_337 (O_337,N_14984,N_14988);
and UO_338 (O_338,N_14917,N_14852);
and UO_339 (O_339,N_14910,N_14936);
nand UO_340 (O_340,N_14978,N_14984);
nand UO_341 (O_341,N_14877,N_14979);
nand UO_342 (O_342,N_14980,N_14888);
nor UO_343 (O_343,N_14932,N_14985);
nor UO_344 (O_344,N_14982,N_14896);
nor UO_345 (O_345,N_14891,N_14980);
xnor UO_346 (O_346,N_14866,N_14906);
nor UO_347 (O_347,N_14888,N_14857);
nor UO_348 (O_348,N_14886,N_14952);
nor UO_349 (O_349,N_14895,N_14876);
nand UO_350 (O_350,N_14858,N_14959);
and UO_351 (O_351,N_14970,N_14926);
xnor UO_352 (O_352,N_14914,N_14988);
and UO_353 (O_353,N_14870,N_14999);
nor UO_354 (O_354,N_14963,N_14907);
xor UO_355 (O_355,N_14862,N_14852);
nand UO_356 (O_356,N_14960,N_14955);
nor UO_357 (O_357,N_14987,N_14983);
or UO_358 (O_358,N_14862,N_14998);
xnor UO_359 (O_359,N_14896,N_14948);
and UO_360 (O_360,N_14983,N_14924);
nand UO_361 (O_361,N_14967,N_14924);
nor UO_362 (O_362,N_14873,N_14863);
and UO_363 (O_363,N_14949,N_14992);
xor UO_364 (O_364,N_14893,N_14897);
nand UO_365 (O_365,N_14897,N_14891);
or UO_366 (O_366,N_14965,N_14921);
nor UO_367 (O_367,N_14875,N_14880);
xnor UO_368 (O_368,N_14860,N_14851);
nand UO_369 (O_369,N_14903,N_14987);
nor UO_370 (O_370,N_14852,N_14978);
and UO_371 (O_371,N_14892,N_14946);
nand UO_372 (O_372,N_14902,N_14946);
nor UO_373 (O_373,N_14978,N_14991);
xor UO_374 (O_374,N_14885,N_14972);
and UO_375 (O_375,N_14958,N_14936);
nor UO_376 (O_376,N_14918,N_14920);
and UO_377 (O_377,N_14930,N_14891);
nor UO_378 (O_378,N_14986,N_14933);
and UO_379 (O_379,N_14866,N_14993);
or UO_380 (O_380,N_14947,N_14977);
or UO_381 (O_381,N_14944,N_14990);
nor UO_382 (O_382,N_14854,N_14858);
and UO_383 (O_383,N_14973,N_14908);
and UO_384 (O_384,N_14899,N_14980);
or UO_385 (O_385,N_14937,N_14973);
nand UO_386 (O_386,N_14969,N_14948);
nand UO_387 (O_387,N_14941,N_14955);
or UO_388 (O_388,N_14869,N_14991);
and UO_389 (O_389,N_14967,N_14888);
nor UO_390 (O_390,N_14961,N_14925);
and UO_391 (O_391,N_14850,N_14857);
xnor UO_392 (O_392,N_14879,N_14934);
nand UO_393 (O_393,N_14867,N_14964);
nor UO_394 (O_394,N_14870,N_14934);
nand UO_395 (O_395,N_14978,N_14935);
or UO_396 (O_396,N_14968,N_14922);
and UO_397 (O_397,N_14929,N_14877);
nand UO_398 (O_398,N_14902,N_14916);
or UO_399 (O_399,N_14957,N_14893);
xor UO_400 (O_400,N_14853,N_14923);
or UO_401 (O_401,N_14978,N_14958);
nor UO_402 (O_402,N_14852,N_14885);
nand UO_403 (O_403,N_14850,N_14957);
nor UO_404 (O_404,N_14971,N_14907);
or UO_405 (O_405,N_14852,N_14929);
nand UO_406 (O_406,N_14915,N_14861);
or UO_407 (O_407,N_14945,N_14887);
nand UO_408 (O_408,N_14983,N_14850);
nor UO_409 (O_409,N_14963,N_14910);
nand UO_410 (O_410,N_14988,N_14949);
or UO_411 (O_411,N_14942,N_14963);
or UO_412 (O_412,N_14943,N_14896);
nor UO_413 (O_413,N_14897,N_14875);
nand UO_414 (O_414,N_14958,N_14870);
nand UO_415 (O_415,N_14980,N_14981);
xor UO_416 (O_416,N_14908,N_14980);
or UO_417 (O_417,N_14944,N_14955);
nand UO_418 (O_418,N_14921,N_14959);
nand UO_419 (O_419,N_14873,N_14914);
nand UO_420 (O_420,N_14926,N_14965);
nor UO_421 (O_421,N_14890,N_14958);
nand UO_422 (O_422,N_14972,N_14916);
and UO_423 (O_423,N_14900,N_14990);
or UO_424 (O_424,N_14939,N_14987);
xnor UO_425 (O_425,N_14908,N_14880);
or UO_426 (O_426,N_14863,N_14943);
nand UO_427 (O_427,N_14871,N_14987);
or UO_428 (O_428,N_14922,N_14891);
nor UO_429 (O_429,N_14851,N_14964);
or UO_430 (O_430,N_14947,N_14918);
xnor UO_431 (O_431,N_14918,N_14981);
xnor UO_432 (O_432,N_14945,N_14957);
nor UO_433 (O_433,N_14908,N_14871);
or UO_434 (O_434,N_14937,N_14981);
or UO_435 (O_435,N_14966,N_14872);
xnor UO_436 (O_436,N_14887,N_14866);
and UO_437 (O_437,N_14854,N_14880);
nor UO_438 (O_438,N_14915,N_14936);
or UO_439 (O_439,N_14906,N_14972);
or UO_440 (O_440,N_14989,N_14911);
xor UO_441 (O_441,N_14997,N_14880);
xnor UO_442 (O_442,N_14924,N_14899);
nand UO_443 (O_443,N_14990,N_14924);
nand UO_444 (O_444,N_14921,N_14863);
and UO_445 (O_445,N_14976,N_14851);
nor UO_446 (O_446,N_14899,N_14931);
nand UO_447 (O_447,N_14965,N_14874);
nor UO_448 (O_448,N_14905,N_14922);
nand UO_449 (O_449,N_14872,N_14851);
nor UO_450 (O_450,N_14961,N_14966);
and UO_451 (O_451,N_14922,N_14960);
and UO_452 (O_452,N_14883,N_14961);
and UO_453 (O_453,N_14871,N_14929);
and UO_454 (O_454,N_14977,N_14991);
xor UO_455 (O_455,N_14898,N_14985);
and UO_456 (O_456,N_14936,N_14906);
xor UO_457 (O_457,N_14899,N_14891);
nor UO_458 (O_458,N_14970,N_14851);
xnor UO_459 (O_459,N_14894,N_14871);
or UO_460 (O_460,N_14881,N_14997);
or UO_461 (O_461,N_14987,N_14865);
nor UO_462 (O_462,N_14960,N_14855);
nand UO_463 (O_463,N_14964,N_14855);
xor UO_464 (O_464,N_14896,N_14936);
and UO_465 (O_465,N_14884,N_14998);
xor UO_466 (O_466,N_14967,N_14889);
nor UO_467 (O_467,N_14984,N_14938);
nand UO_468 (O_468,N_14997,N_14991);
xnor UO_469 (O_469,N_14915,N_14973);
nand UO_470 (O_470,N_14897,N_14994);
and UO_471 (O_471,N_14957,N_14936);
xnor UO_472 (O_472,N_14963,N_14857);
xor UO_473 (O_473,N_14941,N_14904);
or UO_474 (O_474,N_14987,N_14943);
or UO_475 (O_475,N_14854,N_14981);
or UO_476 (O_476,N_14900,N_14913);
and UO_477 (O_477,N_14980,N_14877);
and UO_478 (O_478,N_14908,N_14958);
nand UO_479 (O_479,N_14883,N_14925);
nor UO_480 (O_480,N_14999,N_14892);
and UO_481 (O_481,N_14998,N_14899);
nand UO_482 (O_482,N_14855,N_14992);
or UO_483 (O_483,N_14978,N_14959);
and UO_484 (O_484,N_14857,N_14960);
nor UO_485 (O_485,N_14913,N_14938);
nor UO_486 (O_486,N_14943,N_14895);
and UO_487 (O_487,N_14889,N_14997);
or UO_488 (O_488,N_14958,N_14911);
and UO_489 (O_489,N_14945,N_14960);
and UO_490 (O_490,N_14928,N_14948);
and UO_491 (O_491,N_14885,N_14897);
xnor UO_492 (O_492,N_14979,N_14892);
nor UO_493 (O_493,N_14899,N_14961);
and UO_494 (O_494,N_14931,N_14951);
nand UO_495 (O_495,N_14926,N_14987);
nor UO_496 (O_496,N_14892,N_14853);
and UO_497 (O_497,N_14885,N_14930);
xor UO_498 (O_498,N_14875,N_14957);
nor UO_499 (O_499,N_14935,N_14899);
or UO_500 (O_500,N_14909,N_14976);
or UO_501 (O_501,N_14988,N_14882);
or UO_502 (O_502,N_14873,N_14884);
or UO_503 (O_503,N_14860,N_14974);
xnor UO_504 (O_504,N_14922,N_14857);
or UO_505 (O_505,N_14970,N_14983);
xnor UO_506 (O_506,N_14863,N_14904);
nor UO_507 (O_507,N_14884,N_14956);
or UO_508 (O_508,N_14912,N_14969);
and UO_509 (O_509,N_14854,N_14874);
nand UO_510 (O_510,N_14895,N_14883);
nor UO_511 (O_511,N_14904,N_14991);
nand UO_512 (O_512,N_14851,N_14856);
and UO_513 (O_513,N_14897,N_14982);
nand UO_514 (O_514,N_14860,N_14855);
nand UO_515 (O_515,N_14997,N_14863);
and UO_516 (O_516,N_14921,N_14961);
nor UO_517 (O_517,N_14884,N_14933);
or UO_518 (O_518,N_14979,N_14881);
nor UO_519 (O_519,N_14980,N_14875);
nor UO_520 (O_520,N_14884,N_14852);
and UO_521 (O_521,N_14898,N_14979);
xor UO_522 (O_522,N_14937,N_14957);
and UO_523 (O_523,N_14987,N_14898);
nor UO_524 (O_524,N_14850,N_14861);
nor UO_525 (O_525,N_14989,N_14915);
or UO_526 (O_526,N_14910,N_14904);
nand UO_527 (O_527,N_14947,N_14889);
nand UO_528 (O_528,N_14952,N_14948);
xor UO_529 (O_529,N_14894,N_14973);
or UO_530 (O_530,N_14943,N_14946);
nand UO_531 (O_531,N_14919,N_14911);
nor UO_532 (O_532,N_14889,N_14908);
nor UO_533 (O_533,N_14910,N_14996);
nor UO_534 (O_534,N_14877,N_14914);
or UO_535 (O_535,N_14926,N_14903);
or UO_536 (O_536,N_14861,N_14960);
and UO_537 (O_537,N_14985,N_14893);
xor UO_538 (O_538,N_14936,N_14981);
nor UO_539 (O_539,N_14870,N_14937);
xor UO_540 (O_540,N_14884,N_14893);
or UO_541 (O_541,N_14907,N_14880);
nor UO_542 (O_542,N_14883,N_14872);
nand UO_543 (O_543,N_14949,N_14930);
and UO_544 (O_544,N_14979,N_14969);
nand UO_545 (O_545,N_14928,N_14999);
or UO_546 (O_546,N_14966,N_14894);
nor UO_547 (O_547,N_14873,N_14932);
nor UO_548 (O_548,N_14875,N_14858);
nand UO_549 (O_549,N_14864,N_14998);
xnor UO_550 (O_550,N_14871,N_14873);
nor UO_551 (O_551,N_14990,N_14962);
nand UO_552 (O_552,N_14873,N_14998);
nor UO_553 (O_553,N_14931,N_14857);
nor UO_554 (O_554,N_14897,N_14928);
nand UO_555 (O_555,N_14856,N_14878);
and UO_556 (O_556,N_14884,N_14991);
xor UO_557 (O_557,N_14886,N_14944);
xnor UO_558 (O_558,N_14974,N_14964);
nand UO_559 (O_559,N_14913,N_14999);
nand UO_560 (O_560,N_14897,N_14955);
and UO_561 (O_561,N_14976,N_14920);
xnor UO_562 (O_562,N_14983,N_14993);
or UO_563 (O_563,N_14942,N_14852);
xnor UO_564 (O_564,N_14932,N_14904);
nand UO_565 (O_565,N_14938,N_14910);
nor UO_566 (O_566,N_14900,N_14968);
and UO_567 (O_567,N_14858,N_14943);
and UO_568 (O_568,N_14983,N_14949);
nand UO_569 (O_569,N_14899,N_14934);
nor UO_570 (O_570,N_14993,N_14896);
and UO_571 (O_571,N_14904,N_14957);
nand UO_572 (O_572,N_14924,N_14969);
nor UO_573 (O_573,N_14970,N_14861);
or UO_574 (O_574,N_14949,N_14852);
xor UO_575 (O_575,N_14874,N_14914);
nor UO_576 (O_576,N_14853,N_14902);
nand UO_577 (O_577,N_14914,N_14860);
nand UO_578 (O_578,N_14898,N_14960);
and UO_579 (O_579,N_14851,N_14903);
nor UO_580 (O_580,N_14887,N_14936);
nor UO_581 (O_581,N_14985,N_14897);
xnor UO_582 (O_582,N_14991,N_14994);
xnor UO_583 (O_583,N_14873,N_14976);
or UO_584 (O_584,N_14920,N_14975);
xor UO_585 (O_585,N_14956,N_14859);
nor UO_586 (O_586,N_14870,N_14994);
nor UO_587 (O_587,N_14918,N_14907);
xor UO_588 (O_588,N_14996,N_14963);
xnor UO_589 (O_589,N_14999,N_14997);
and UO_590 (O_590,N_14943,N_14966);
nor UO_591 (O_591,N_14935,N_14873);
xor UO_592 (O_592,N_14955,N_14940);
xor UO_593 (O_593,N_14851,N_14869);
nor UO_594 (O_594,N_14905,N_14902);
nor UO_595 (O_595,N_14912,N_14939);
and UO_596 (O_596,N_14896,N_14893);
nor UO_597 (O_597,N_14940,N_14965);
nor UO_598 (O_598,N_14879,N_14881);
nand UO_599 (O_599,N_14923,N_14979);
and UO_600 (O_600,N_14883,N_14864);
xor UO_601 (O_601,N_14901,N_14988);
nand UO_602 (O_602,N_14977,N_14976);
nand UO_603 (O_603,N_14872,N_14874);
and UO_604 (O_604,N_14956,N_14949);
and UO_605 (O_605,N_14902,N_14922);
and UO_606 (O_606,N_14969,N_14926);
nand UO_607 (O_607,N_14928,N_14944);
xnor UO_608 (O_608,N_14866,N_14938);
or UO_609 (O_609,N_14971,N_14906);
and UO_610 (O_610,N_14948,N_14999);
nand UO_611 (O_611,N_14994,N_14929);
and UO_612 (O_612,N_14862,N_14981);
and UO_613 (O_613,N_14882,N_14898);
and UO_614 (O_614,N_14932,N_14912);
nor UO_615 (O_615,N_14861,N_14990);
xor UO_616 (O_616,N_14893,N_14904);
xor UO_617 (O_617,N_14934,N_14983);
nand UO_618 (O_618,N_14918,N_14950);
nand UO_619 (O_619,N_14931,N_14876);
xor UO_620 (O_620,N_14933,N_14882);
and UO_621 (O_621,N_14850,N_14980);
or UO_622 (O_622,N_14934,N_14855);
and UO_623 (O_623,N_14903,N_14863);
and UO_624 (O_624,N_14950,N_14983);
or UO_625 (O_625,N_14880,N_14866);
xor UO_626 (O_626,N_14926,N_14948);
nor UO_627 (O_627,N_14987,N_14949);
or UO_628 (O_628,N_14876,N_14882);
or UO_629 (O_629,N_14858,N_14923);
and UO_630 (O_630,N_14866,N_14875);
and UO_631 (O_631,N_14990,N_14948);
and UO_632 (O_632,N_14896,N_14966);
xor UO_633 (O_633,N_14897,N_14869);
nand UO_634 (O_634,N_14879,N_14989);
nor UO_635 (O_635,N_14892,N_14869);
nor UO_636 (O_636,N_14874,N_14868);
nand UO_637 (O_637,N_14989,N_14896);
xnor UO_638 (O_638,N_14868,N_14904);
or UO_639 (O_639,N_14866,N_14885);
and UO_640 (O_640,N_14922,N_14942);
nand UO_641 (O_641,N_14914,N_14964);
and UO_642 (O_642,N_14932,N_14925);
nor UO_643 (O_643,N_14912,N_14984);
or UO_644 (O_644,N_14868,N_14908);
nand UO_645 (O_645,N_14899,N_14950);
and UO_646 (O_646,N_14915,N_14920);
nor UO_647 (O_647,N_14880,N_14973);
xor UO_648 (O_648,N_14850,N_14974);
and UO_649 (O_649,N_14914,N_14987);
xnor UO_650 (O_650,N_14969,N_14925);
and UO_651 (O_651,N_14860,N_14884);
and UO_652 (O_652,N_14920,N_14985);
nor UO_653 (O_653,N_14879,N_14912);
nor UO_654 (O_654,N_14881,N_14905);
xnor UO_655 (O_655,N_14851,N_14971);
and UO_656 (O_656,N_14998,N_14953);
and UO_657 (O_657,N_14902,N_14990);
nor UO_658 (O_658,N_14902,N_14980);
nand UO_659 (O_659,N_14859,N_14987);
or UO_660 (O_660,N_14977,N_14873);
nand UO_661 (O_661,N_14902,N_14958);
or UO_662 (O_662,N_14896,N_14886);
nor UO_663 (O_663,N_14900,N_14893);
xnor UO_664 (O_664,N_14920,N_14941);
or UO_665 (O_665,N_14993,N_14895);
xor UO_666 (O_666,N_14981,N_14868);
and UO_667 (O_667,N_14983,N_14913);
and UO_668 (O_668,N_14950,N_14938);
xnor UO_669 (O_669,N_14986,N_14871);
nor UO_670 (O_670,N_14863,N_14866);
nor UO_671 (O_671,N_14971,N_14943);
nand UO_672 (O_672,N_14875,N_14965);
and UO_673 (O_673,N_14891,N_14936);
nand UO_674 (O_674,N_14930,N_14981);
and UO_675 (O_675,N_14934,N_14982);
or UO_676 (O_676,N_14977,N_14995);
and UO_677 (O_677,N_14923,N_14938);
xnor UO_678 (O_678,N_14935,N_14854);
or UO_679 (O_679,N_14935,N_14857);
and UO_680 (O_680,N_14957,N_14984);
xnor UO_681 (O_681,N_14870,N_14941);
or UO_682 (O_682,N_14869,N_14932);
and UO_683 (O_683,N_14968,N_14918);
nand UO_684 (O_684,N_14894,N_14921);
and UO_685 (O_685,N_14978,N_14887);
nor UO_686 (O_686,N_14862,N_14945);
xnor UO_687 (O_687,N_14921,N_14944);
or UO_688 (O_688,N_14894,N_14852);
and UO_689 (O_689,N_14999,N_14956);
nor UO_690 (O_690,N_14955,N_14908);
or UO_691 (O_691,N_14926,N_14916);
xnor UO_692 (O_692,N_14960,N_14907);
nor UO_693 (O_693,N_14920,N_14936);
nand UO_694 (O_694,N_14964,N_14900);
or UO_695 (O_695,N_14886,N_14862);
and UO_696 (O_696,N_14935,N_14976);
xor UO_697 (O_697,N_14935,N_14909);
nor UO_698 (O_698,N_14906,N_14874);
and UO_699 (O_699,N_14930,N_14861);
or UO_700 (O_700,N_14957,N_14920);
or UO_701 (O_701,N_14961,N_14857);
nor UO_702 (O_702,N_14875,N_14986);
xnor UO_703 (O_703,N_14963,N_14966);
and UO_704 (O_704,N_14971,N_14879);
xor UO_705 (O_705,N_14876,N_14962);
xor UO_706 (O_706,N_14949,N_14913);
and UO_707 (O_707,N_14905,N_14913);
and UO_708 (O_708,N_14996,N_14895);
nand UO_709 (O_709,N_14980,N_14897);
nor UO_710 (O_710,N_14980,N_14890);
and UO_711 (O_711,N_14937,N_14967);
xor UO_712 (O_712,N_14865,N_14900);
nand UO_713 (O_713,N_14867,N_14923);
or UO_714 (O_714,N_14906,N_14934);
or UO_715 (O_715,N_14870,N_14891);
and UO_716 (O_716,N_14934,N_14986);
nand UO_717 (O_717,N_14873,N_14981);
nor UO_718 (O_718,N_14879,N_14902);
xnor UO_719 (O_719,N_14917,N_14880);
and UO_720 (O_720,N_14872,N_14989);
nor UO_721 (O_721,N_14884,N_14951);
nand UO_722 (O_722,N_14907,N_14942);
nand UO_723 (O_723,N_14974,N_14857);
nand UO_724 (O_724,N_14926,N_14946);
nand UO_725 (O_725,N_14988,N_14986);
xor UO_726 (O_726,N_14948,N_14972);
nor UO_727 (O_727,N_14998,N_14911);
nor UO_728 (O_728,N_14949,N_14946);
nand UO_729 (O_729,N_14984,N_14923);
and UO_730 (O_730,N_14932,N_14964);
nor UO_731 (O_731,N_14967,N_14958);
and UO_732 (O_732,N_14865,N_14860);
nand UO_733 (O_733,N_14904,N_14980);
or UO_734 (O_734,N_14986,N_14902);
nand UO_735 (O_735,N_14893,N_14876);
xor UO_736 (O_736,N_14895,N_14985);
xnor UO_737 (O_737,N_14870,N_14886);
or UO_738 (O_738,N_14937,N_14900);
xnor UO_739 (O_739,N_14946,N_14887);
nand UO_740 (O_740,N_14894,N_14858);
nor UO_741 (O_741,N_14909,N_14891);
and UO_742 (O_742,N_14973,N_14938);
or UO_743 (O_743,N_14998,N_14946);
nand UO_744 (O_744,N_14994,N_14892);
xnor UO_745 (O_745,N_14937,N_14929);
nand UO_746 (O_746,N_14942,N_14885);
xnor UO_747 (O_747,N_14888,N_14852);
or UO_748 (O_748,N_14870,N_14864);
or UO_749 (O_749,N_14986,N_14938);
xnor UO_750 (O_750,N_14880,N_14925);
or UO_751 (O_751,N_14956,N_14856);
or UO_752 (O_752,N_14858,N_14896);
nor UO_753 (O_753,N_14921,N_14987);
nor UO_754 (O_754,N_14933,N_14998);
or UO_755 (O_755,N_14866,N_14989);
or UO_756 (O_756,N_14862,N_14895);
and UO_757 (O_757,N_14877,N_14996);
xor UO_758 (O_758,N_14904,N_14908);
or UO_759 (O_759,N_14959,N_14970);
or UO_760 (O_760,N_14873,N_14893);
or UO_761 (O_761,N_14911,N_14987);
nand UO_762 (O_762,N_14909,N_14921);
or UO_763 (O_763,N_14911,N_14879);
or UO_764 (O_764,N_14990,N_14886);
nor UO_765 (O_765,N_14873,N_14941);
nor UO_766 (O_766,N_14910,N_14862);
and UO_767 (O_767,N_14918,N_14990);
or UO_768 (O_768,N_14888,N_14882);
nor UO_769 (O_769,N_14945,N_14998);
and UO_770 (O_770,N_14983,N_14976);
or UO_771 (O_771,N_14867,N_14894);
nand UO_772 (O_772,N_14863,N_14874);
and UO_773 (O_773,N_14946,N_14853);
xnor UO_774 (O_774,N_14971,N_14933);
and UO_775 (O_775,N_14930,N_14982);
nor UO_776 (O_776,N_14865,N_14872);
or UO_777 (O_777,N_14983,N_14947);
nor UO_778 (O_778,N_14985,N_14875);
xnor UO_779 (O_779,N_14988,N_14930);
nor UO_780 (O_780,N_14887,N_14919);
and UO_781 (O_781,N_14954,N_14855);
nand UO_782 (O_782,N_14951,N_14926);
or UO_783 (O_783,N_14996,N_14896);
xor UO_784 (O_784,N_14850,N_14929);
xor UO_785 (O_785,N_14978,N_14909);
nand UO_786 (O_786,N_14928,N_14857);
xor UO_787 (O_787,N_14879,N_14909);
nand UO_788 (O_788,N_14911,N_14907);
or UO_789 (O_789,N_14994,N_14891);
nor UO_790 (O_790,N_14915,N_14962);
nor UO_791 (O_791,N_14998,N_14901);
xnor UO_792 (O_792,N_14896,N_14883);
nand UO_793 (O_793,N_14857,N_14955);
xor UO_794 (O_794,N_14895,N_14968);
nor UO_795 (O_795,N_14879,N_14882);
or UO_796 (O_796,N_14906,N_14859);
nand UO_797 (O_797,N_14949,N_14964);
nand UO_798 (O_798,N_14874,N_14983);
xor UO_799 (O_799,N_14878,N_14911);
nor UO_800 (O_800,N_14963,N_14887);
nand UO_801 (O_801,N_14912,N_14908);
and UO_802 (O_802,N_14871,N_14858);
xnor UO_803 (O_803,N_14869,N_14914);
nor UO_804 (O_804,N_14916,N_14853);
or UO_805 (O_805,N_14903,N_14859);
nand UO_806 (O_806,N_14867,N_14932);
or UO_807 (O_807,N_14872,N_14854);
xor UO_808 (O_808,N_14864,N_14918);
nand UO_809 (O_809,N_14861,N_14962);
or UO_810 (O_810,N_14954,N_14851);
nand UO_811 (O_811,N_14932,N_14940);
nand UO_812 (O_812,N_14864,N_14954);
xnor UO_813 (O_813,N_14895,N_14945);
or UO_814 (O_814,N_14932,N_14898);
xor UO_815 (O_815,N_14982,N_14958);
nand UO_816 (O_816,N_14928,N_14959);
or UO_817 (O_817,N_14880,N_14897);
and UO_818 (O_818,N_14927,N_14968);
or UO_819 (O_819,N_14886,N_14910);
nor UO_820 (O_820,N_14990,N_14907);
or UO_821 (O_821,N_14864,N_14956);
nand UO_822 (O_822,N_14872,N_14879);
and UO_823 (O_823,N_14963,N_14921);
and UO_824 (O_824,N_14955,N_14901);
nor UO_825 (O_825,N_14983,N_14997);
or UO_826 (O_826,N_14858,N_14856);
nand UO_827 (O_827,N_14945,N_14918);
xnor UO_828 (O_828,N_14850,N_14944);
nor UO_829 (O_829,N_14859,N_14865);
and UO_830 (O_830,N_14898,N_14890);
nand UO_831 (O_831,N_14873,N_14909);
nand UO_832 (O_832,N_14852,N_14909);
xnor UO_833 (O_833,N_14904,N_14888);
xnor UO_834 (O_834,N_14958,N_14854);
nor UO_835 (O_835,N_14876,N_14992);
and UO_836 (O_836,N_14891,N_14992);
xor UO_837 (O_837,N_14927,N_14988);
xor UO_838 (O_838,N_14954,N_14957);
and UO_839 (O_839,N_14974,N_14897);
nand UO_840 (O_840,N_14851,N_14996);
or UO_841 (O_841,N_14896,N_14882);
or UO_842 (O_842,N_14870,N_14913);
xnor UO_843 (O_843,N_14883,N_14940);
nor UO_844 (O_844,N_14900,N_14853);
nor UO_845 (O_845,N_14876,N_14956);
or UO_846 (O_846,N_14975,N_14982);
and UO_847 (O_847,N_14863,N_14861);
nand UO_848 (O_848,N_14867,N_14892);
or UO_849 (O_849,N_14967,N_14873);
and UO_850 (O_850,N_14893,N_14865);
xnor UO_851 (O_851,N_14933,N_14898);
or UO_852 (O_852,N_14896,N_14971);
nor UO_853 (O_853,N_14871,N_14950);
xor UO_854 (O_854,N_14989,N_14951);
nand UO_855 (O_855,N_14896,N_14926);
xor UO_856 (O_856,N_14936,N_14893);
nor UO_857 (O_857,N_14935,N_14929);
or UO_858 (O_858,N_14917,N_14954);
nor UO_859 (O_859,N_14914,N_14894);
or UO_860 (O_860,N_14969,N_14986);
xnor UO_861 (O_861,N_14978,N_14979);
and UO_862 (O_862,N_14866,N_14977);
nand UO_863 (O_863,N_14948,N_14941);
or UO_864 (O_864,N_14927,N_14864);
xor UO_865 (O_865,N_14901,N_14867);
nand UO_866 (O_866,N_14999,N_14862);
xnor UO_867 (O_867,N_14953,N_14951);
or UO_868 (O_868,N_14936,N_14956);
or UO_869 (O_869,N_14856,N_14987);
nor UO_870 (O_870,N_14906,N_14887);
or UO_871 (O_871,N_14901,N_14999);
nor UO_872 (O_872,N_14943,N_14870);
nand UO_873 (O_873,N_14912,N_14894);
or UO_874 (O_874,N_14915,N_14862);
xnor UO_875 (O_875,N_14981,N_14997);
and UO_876 (O_876,N_14949,N_14877);
or UO_877 (O_877,N_14975,N_14869);
nor UO_878 (O_878,N_14865,N_14857);
or UO_879 (O_879,N_14935,N_14958);
or UO_880 (O_880,N_14876,N_14878);
nand UO_881 (O_881,N_14870,N_14900);
and UO_882 (O_882,N_14944,N_14984);
nor UO_883 (O_883,N_14987,N_14970);
xor UO_884 (O_884,N_14966,N_14900);
or UO_885 (O_885,N_14996,N_14893);
or UO_886 (O_886,N_14857,N_14964);
or UO_887 (O_887,N_14908,N_14922);
nor UO_888 (O_888,N_14899,N_14873);
xor UO_889 (O_889,N_14975,N_14925);
xnor UO_890 (O_890,N_14929,N_14908);
xnor UO_891 (O_891,N_14963,N_14903);
or UO_892 (O_892,N_14993,N_14919);
or UO_893 (O_893,N_14854,N_14983);
nor UO_894 (O_894,N_14947,N_14927);
and UO_895 (O_895,N_14961,N_14971);
nor UO_896 (O_896,N_14885,N_14868);
nand UO_897 (O_897,N_14917,N_14898);
xor UO_898 (O_898,N_14986,N_14947);
and UO_899 (O_899,N_14998,N_14893);
xnor UO_900 (O_900,N_14990,N_14981);
nor UO_901 (O_901,N_14955,N_14917);
nor UO_902 (O_902,N_14975,N_14865);
xnor UO_903 (O_903,N_14850,N_14995);
nor UO_904 (O_904,N_14984,N_14994);
nand UO_905 (O_905,N_14972,N_14969);
or UO_906 (O_906,N_14869,N_14887);
or UO_907 (O_907,N_14976,N_14993);
and UO_908 (O_908,N_14885,N_14993);
nor UO_909 (O_909,N_14946,N_14987);
nand UO_910 (O_910,N_14964,N_14881);
nor UO_911 (O_911,N_14985,N_14999);
or UO_912 (O_912,N_14923,N_14972);
and UO_913 (O_913,N_14924,N_14960);
xnor UO_914 (O_914,N_14894,N_14886);
or UO_915 (O_915,N_14992,N_14996);
xnor UO_916 (O_916,N_14930,N_14971);
or UO_917 (O_917,N_14861,N_14978);
nand UO_918 (O_918,N_14941,N_14939);
or UO_919 (O_919,N_14968,N_14886);
xnor UO_920 (O_920,N_14907,N_14902);
nor UO_921 (O_921,N_14862,N_14952);
nor UO_922 (O_922,N_14900,N_14954);
nand UO_923 (O_923,N_14970,N_14893);
or UO_924 (O_924,N_14989,N_14944);
xor UO_925 (O_925,N_14940,N_14938);
or UO_926 (O_926,N_14877,N_14933);
and UO_927 (O_927,N_14920,N_14929);
nand UO_928 (O_928,N_14879,N_14973);
nor UO_929 (O_929,N_14921,N_14861);
and UO_930 (O_930,N_14941,N_14963);
nor UO_931 (O_931,N_14899,N_14897);
xnor UO_932 (O_932,N_14888,N_14889);
or UO_933 (O_933,N_14858,N_14851);
and UO_934 (O_934,N_14915,N_14921);
and UO_935 (O_935,N_14873,N_14885);
xnor UO_936 (O_936,N_14990,N_14925);
and UO_937 (O_937,N_14986,N_14857);
xnor UO_938 (O_938,N_14989,N_14883);
or UO_939 (O_939,N_14872,N_14875);
and UO_940 (O_940,N_14898,N_14903);
nand UO_941 (O_941,N_14883,N_14975);
nand UO_942 (O_942,N_14963,N_14946);
and UO_943 (O_943,N_14972,N_14974);
nand UO_944 (O_944,N_14974,N_14958);
or UO_945 (O_945,N_14996,N_14881);
and UO_946 (O_946,N_14920,N_14988);
or UO_947 (O_947,N_14989,N_14990);
or UO_948 (O_948,N_14949,N_14965);
nor UO_949 (O_949,N_14854,N_14868);
nand UO_950 (O_950,N_14895,N_14896);
nor UO_951 (O_951,N_14916,N_14864);
and UO_952 (O_952,N_14972,N_14889);
and UO_953 (O_953,N_14949,N_14929);
xor UO_954 (O_954,N_14972,N_14918);
xor UO_955 (O_955,N_14932,N_14998);
xor UO_956 (O_956,N_14902,N_14859);
nor UO_957 (O_957,N_14892,N_14877);
xnor UO_958 (O_958,N_14865,N_14977);
nor UO_959 (O_959,N_14965,N_14878);
xor UO_960 (O_960,N_14921,N_14878);
or UO_961 (O_961,N_14880,N_14942);
and UO_962 (O_962,N_14883,N_14991);
and UO_963 (O_963,N_14875,N_14907);
nand UO_964 (O_964,N_14921,N_14974);
and UO_965 (O_965,N_14988,N_14987);
nand UO_966 (O_966,N_14875,N_14890);
nand UO_967 (O_967,N_14872,N_14934);
xor UO_968 (O_968,N_14855,N_14922);
nor UO_969 (O_969,N_14930,N_14961);
nand UO_970 (O_970,N_14933,N_14881);
nor UO_971 (O_971,N_14990,N_14973);
nand UO_972 (O_972,N_14979,N_14897);
nand UO_973 (O_973,N_14893,N_14992);
and UO_974 (O_974,N_14922,N_14956);
xor UO_975 (O_975,N_14893,N_14888);
nand UO_976 (O_976,N_14864,N_14881);
xnor UO_977 (O_977,N_14996,N_14933);
xor UO_978 (O_978,N_14975,N_14997);
xor UO_979 (O_979,N_14914,N_14866);
xnor UO_980 (O_980,N_14876,N_14989);
xor UO_981 (O_981,N_14975,N_14944);
or UO_982 (O_982,N_14903,N_14850);
or UO_983 (O_983,N_14977,N_14879);
xor UO_984 (O_984,N_14868,N_14925);
xor UO_985 (O_985,N_14982,N_14940);
nand UO_986 (O_986,N_14888,N_14868);
and UO_987 (O_987,N_14884,N_14937);
and UO_988 (O_988,N_14913,N_14978);
nand UO_989 (O_989,N_14853,N_14930);
xnor UO_990 (O_990,N_14888,N_14922);
nand UO_991 (O_991,N_14869,N_14927);
and UO_992 (O_992,N_14852,N_14956);
xor UO_993 (O_993,N_14978,N_14900);
or UO_994 (O_994,N_14852,N_14940);
or UO_995 (O_995,N_14997,N_14872);
xnor UO_996 (O_996,N_14897,N_14941);
and UO_997 (O_997,N_14910,N_14926);
and UO_998 (O_998,N_14923,N_14927);
nor UO_999 (O_999,N_14856,N_14993);
nand UO_1000 (O_1000,N_14878,N_14957);
nand UO_1001 (O_1001,N_14876,N_14970);
and UO_1002 (O_1002,N_14912,N_14852);
nor UO_1003 (O_1003,N_14893,N_14890);
or UO_1004 (O_1004,N_14989,N_14906);
nor UO_1005 (O_1005,N_14957,N_14944);
nand UO_1006 (O_1006,N_14965,N_14905);
nor UO_1007 (O_1007,N_14873,N_14860);
or UO_1008 (O_1008,N_14884,N_14875);
and UO_1009 (O_1009,N_14894,N_14889);
xor UO_1010 (O_1010,N_14960,N_14853);
and UO_1011 (O_1011,N_14977,N_14943);
and UO_1012 (O_1012,N_14865,N_14911);
xor UO_1013 (O_1013,N_14948,N_14923);
nor UO_1014 (O_1014,N_14949,N_14853);
xnor UO_1015 (O_1015,N_14987,N_14900);
xor UO_1016 (O_1016,N_14923,N_14997);
nor UO_1017 (O_1017,N_14915,N_14888);
xor UO_1018 (O_1018,N_14923,N_14956);
xor UO_1019 (O_1019,N_14947,N_14872);
nand UO_1020 (O_1020,N_14967,N_14925);
nand UO_1021 (O_1021,N_14864,N_14932);
nand UO_1022 (O_1022,N_14989,N_14878);
or UO_1023 (O_1023,N_14905,N_14850);
xnor UO_1024 (O_1024,N_14946,N_14888);
nor UO_1025 (O_1025,N_14988,N_14874);
nor UO_1026 (O_1026,N_14990,N_14856);
nand UO_1027 (O_1027,N_14946,N_14939);
and UO_1028 (O_1028,N_14862,N_14959);
nand UO_1029 (O_1029,N_14983,N_14852);
nor UO_1030 (O_1030,N_14947,N_14997);
and UO_1031 (O_1031,N_14900,N_14953);
nor UO_1032 (O_1032,N_14882,N_14919);
and UO_1033 (O_1033,N_14960,N_14854);
or UO_1034 (O_1034,N_14995,N_14912);
and UO_1035 (O_1035,N_14852,N_14928);
xor UO_1036 (O_1036,N_14939,N_14864);
and UO_1037 (O_1037,N_14875,N_14970);
nand UO_1038 (O_1038,N_14905,N_14997);
xnor UO_1039 (O_1039,N_14851,N_14912);
and UO_1040 (O_1040,N_14989,N_14930);
xor UO_1041 (O_1041,N_14913,N_14867);
xnor UO_1042 (O_1042,N_14948,N_14907);
nor UO_1043 (O_1043,N_14853,N_14905);
and UO_1044 (O_1044,N_14908,N_14851);
nor UO_1045 (O_1045,N_14854,N_14945);
nand UO_1046 (O_1046,N_14947,N_14957);
and UO_1047 (O_1047,N_14902,N_14952);
or UO_1048 (O_1048,N_14858,N_14969);
or UO_1049 (O_1049,N_14956,N_14978);
nor UO_1050 (O_1050,N_14950,N_14975);
or UO_1051 (O_1051,N_14918,N_14883);
nor UO_1052 (O_1052,N_14928,N_14916);
and UO_1053 (O_1053,N_14867,N_14914);
xor UO_1054 (O_1054,N_14973,N_14993);
or UO_1055 (O_1055,N_14881,N_14910);
nand UO_1056 (O_1056,N_14997,N_14936);
nand UO_1057 (O_1057,N_14968,N_14996);
nand UO_1058 (O_1058,N_14942,N_14884);
xor UO_1059 (O_1059,N_14878,N_14997);
nand UO_1060 (O_1060,N_14932,N_14975);
nand UO_1061 (O_1061,N_14956,N_14901);
nor UO_1062 (O_1062,N_14975,N_14957);
or UO_1063 (O_1063,N_14976,N_14933);
xnor UO_1064 (O_1064,N_14945,N_14954);
xnor UO_1065 (O_1065,N_14852,N_14948);
and UO_1066 (O_1066,N_14891,N_14910);
nand UO_1067 (O_1067,N_14920,N_14874);
xor UO_1068 (O_1068,N_14929,N_14853);
nand UO_1069 (O_1069,N_14857,N_14973);
and UO_1070 (O_1070,N_14902,N_14850);
nor UO_1071 (O_1071,N_14924,N_14982);
or UO_1072 (O_1072,N_14877,N_14934);
and UO_1073 (O_1073,N_14985,N_14980);
nor UO_1074 (O_1074,N_14852,N_14866);
nand UO_1075 (O_1075,N_14869,N_14923);
or UO_1076 (O_1076,N_14942,N_14920);
nand UO_1077 (O_1077,N_14997,N_14993);
xnor UO_1078 (O_1078,N_14999,N_14949);
nand UO_1079 (O_1079,N_14995,N_14886);
or UO_1080 (O_1080,N_14872,N_14969);
nor UO_1081 (O_1081,N_14897,N_14850);
or UO_1082 (O_1082,N_14974,N_14892);
and UO_1083 (O_1083,N_14852,N_14927);
xor UO_1084 (O_1084,N_14917,N_14928);
xnor UO_1085 (O_1085,N_14974,N_14912);
xnor UO_1086 (O_1086,N_14912,N_14876);
xor UO_1087 (O_1087,N_14923,N_14879);
nand UO_1088 (O_1088,N_14913,N_14930);
and UO_1089 (O_1089,N_14942,N_14900);
xnor UO_1090 (O_1090,N_14863,N_14981);
and UO_1091 (O_1091,N_14923,N_14911);
nand UO_1092 (O_1092,N_14888,N_14883);
and UO_1093 (O_1093,N_14869,N_14879);
or UO_1094 (O_1094,N_14889,N_14981);
or UO_1095 (O_1095,N_14904,N_14853);
nor UO_1096 (O_1096,N_14925,N_14972);
nand UO_1097 (O_1097,N_14949,N_14980);
nor UO_1098 (O_1098,N_14976,N_14903);
and UO_1099 (O_1099,N_14962,N_14874);
xnor UO_1100 (O_1100,N_14961,N_14957);
nand UO_1101 (O_1101,N_14990,N_14928);
or UO_1102 (O_1102,N_14906,N_14888);
or UO_1103 (O_1103,N_14961,N_14953);
nand UO_1104 (O_1104,N_14938,N_14879);
or UO_1105 (O_1105,N_14853,N_14925);
nand UO_1106 (O_1106,N_14856,N_14958);
or UO_1107 (O_1107,N_14921,N_14870);
or UO_1108 (O_1108,N_14978,N_14876);
xor UO_1109 (O_1109,N_14988,N_14969);
and UO_1110 (O_1110,N_14988,N_14963);
xor UO_1111 (O_1111,N_14975,N_14968);
and UO_1112 (O_1112,N_14912,N_14895);
xnor UO_1113 (O_1113,N_14924,N_14918);
and UO_1114 (O_1114,N_14939,N_14871);
nand UO_1115 (O_1115,N_14944,N_14997);
or UO_1116 (O_1116,N_14934,N_14975);
nor UO_1117 (O_1117,N_14886,N_14958);
or UO_1118 (O_1118,N_14900,N_14896);
and UO_1119 (O_1119,N_14928,N_14908);
nor UO_1120 (O_1120,N_14915,N_14935);
nand UO_1121 (O_1121,N_14851,N_14917);
and UO_1122 (O_1122,N_14895,N_14941);
and UO_1123 (O_1123,N_14970,N_14952);
nor UO_1124 (O_1124,N_14854,N_14877);
xor UO_1125 (O_1125,N_14893,N_14880);
and UO_1126 (O_1126,N_14953,N_14916);
or UO_1127 (O_1127,N_14986,N_14959);
nand UO_1128 (O_1128,N_14859,N_14914);
nand UO_1129 (O_1129,N_14967,N_14935);
nand UO_1130 (O_1130,N_14958,N_14995);
or UO_1131 (O_1131,N_14989,N_14855);
and UO_1132 (O_1132,N_14996,N_14875);
nand UO_1133 (O_1133,N_14905,N_14956);
nand UO_1134 (O_1134,N_14971,N_14953);
nor UO_1135 (O_1135,N_14943,N_14956);
xor UO_1136 (O_1136,N_14913,N_14887);
xor UO_1137 (O_1137,N_14867,N_14893);
xnor UO_1138 (O_1138,N_14921,N_14991);
nand UO_1139 (O_1139,N_14867,N_14882);
and UO_1140 (O_1140,N_14870,N_14855);
or UO_1141 (O_1141,N_14912,N_14913);
xnor UO_1142 (O_1142,N_14854,N_14995);
nand UO_1143 (O_1143,N_14907,N_14864);
nand UO_1144 (O_1144,N_14962,N_14859);
nor UO_1145 (O_1145,N_14979,N_14975);
nor UO_1146 (O_1146,N_14975,N_14894);
xnor UO_1147 (O_1147,N_14934,N_14859);
and UO_1148 (O_1148,N_14959,N_14859);
and UO_1149 (O_1149,N_14970,N_14873);
xnor UO_1150 (O_1150,N_14858,N_14997);
nor UO_1151 (O_1151,N_14909,N_14874);
and UO_1152 (O_1152,N_14871,N_14911);
or UO_1153 (O_1153,N_14979,N_14988);
and UO_1154 (O_1154,N_14984,N_14981);
and UO_1155 (O_1155,N_14890,N_14895);
nor UO_1156 (O_1156,N_14996,N_14962);
nand UO_1157 (O_1157,N_14987,N_14915);
nor UO_1158 (O_1158,N_14932,N_14914);
or UO_1159 (O_1159,N_14933,N_14934);
nand UO_1160 (O_1160,N_14926,N_14862);
nor UO_1161 (O_1161,N_14929,N_14999);
xnor UO_1162 (O_1162,N_14856,N_14965);
or UO_1163 (O_1163,N_14966,N_14926);
and UO_1164 (O_1164,N_14886,N_14997);
xor UO_1165 (O_1165,N_14933,N_14940);
nor UO_1166 (O_1166,N_14888,N_14986);
nor UO_1167 (O_1167,N_14862,N_14958);
or UO_1168 (O_1168,N_14942,N_14977);
and UO_1169 (O_1169,N_14895,N_14944);
xor UO_1170 (O_1170,N_14851,N_14914);
xnor UO_1171 (O_1171,N_14897,N_14973);
and UO_1172 (O_1172,N_14850,N_14955);
or UO_1173 (O_1173,N_14954,N_14946);
and UO_1174 (O_1174,N_14880,N_14946);
nand UO_1175 (O_1175,N_14997,N_14995);
or UO_1176 (O_1176,N_14960,N_14871);
and UO_1177 (O_1177,N_14976,N_14904);
or UO_1178 (O_1178,N_14935,N_14913);
and UO_1179 (O_1179,N_14969,N_14930);
nand UO_1180 (O_1180,N_14945,N_14910);
nand UO_1181 (O_1181,N_14926,N_14958);
xor UO_1182 (O_1182,N_14868,N_14955);
nand UO_1183 (O_1183,N_14892,N_14930);
or UO_1184 (O_1184,N_14907,N_14946);
or UO_1185 (O_1185,N_14942,N_14991);
xnor UO_1186 (O_1186,N_14891,N_14863);
xor UO_1187 (O_1187,N_14866,N_14997);
and UO_1188 (O_1188,N_14911,N_14933);
or UO_1189 (O_1189,N_14853,N_14964);
nor UO_1190 (O_1190,N_14906,N_14894);
xor UO_1191 (O_1191,N_14861,N_14890);
xor UO_1192 (O_1192,N_14958,N_14899);
nor UO_1193 (O_1193,N_14882,N_14960);
xnor UO_1194 (O_1194,N_14873,N_14891);
xor UO_1195 (O_1195,N_14970,N_14912);
or UO_1196 (O_1196,N_14912,N_14890);
xnor UO_1197 (O_1197,N_14994,N_14921);
nand UO_1198 (O_1198,N_14901,N_14975);
nand UO_1199 (O_1199,N_14855,N_14852);
nor UO_1200 (O_1200,N_14970,N_14880);
nand UO_1201 (O_1201,N_14850,N_14867);
and UO_1202 (O_1202,N_14967,N_14916);
and UO_1203 (O_1203,N_14983,N_14862);
or UO_1204 (O_1204,N_14927,N_14946);
and UO_1205 (O_1205,N_14909,N_14924);
or UO_1206 (O_1206,N_14959,N_14977);
xnor UO_1207 (O_1207,N_14920,N_14952);
xor UO_1208 (O_1208,N_14857,N_14880);
or UO_1209 (O_1209,N_14851,N_14928);
nor UO_1210 (O_1210,N_14969,N_14935);
nor UO_1211 (O_1211,N_14909,N_14910);
or UO_1212 (O_1212,N_14960,N_14972);
nor UO_1213 (O_1213,N_14914,N_14888);
or UO_1214 (O_1214,N_14945,N_14881);
nor UO_1215 (O_1215,N_14870,N_14978);
or UO_1216 (O_1216,N_14937,N_14994);
nand UO_1217 (O_1217,N_14860,N_14972);
xor UO_1218 (O_1218,N_14907,N_14855);
or UO_1219 (O_1219,N_14903,N_14979);
or UO_1220 (O_1220,N_14908,N_14999);
nand UO_1221 (O_1221,N_14992,N_14887);
and UO_1222 (O_1222,N_14990,N_14938);
or UO_1223 (O_1223,N_14855,N_14950);
or UO_1224 (O_1224,N_14856,N_14864);
nand UO_1225 (O_1225,N_14913,N_14892);
and UO_1226 (O_1226,N_14987,N_14936);
xnor UO_1227 (O_1227,N_14975,N_14939);
xor UO_1228 (O_1228,N_14946,N_14885);
xor UO_1229 (O_1229,N_14913,N_14921);
nand UO_1230 (O_1230,N_14863,N_14934);
nand UO_1231 (O_1231,N_14937,N_14955);
xor UO_1232 (O_1232,N_14880,N_14981);
xor UO_1233 (O_1233,N_14985,N_14969);
xnor UO_1234 (O_1234,N_14943,N_14950);
nand UO_1235 (O_1235,N_14902,N_14966);
xnor UO_1236 (O_1236,N_14910,N_14998);
xnor UO_1237 (O_1237,N_14862,N_14923);
nand UO_1238 (O_1238,N_14871,N_14930);
nor UO_1239 (O_1239,N_14936,N_14952);
nor UO_1240 (O_1240,N_14901,N_14887);
xnor UO_1241 (O_1241,N_14929,N_14875);
or UO_1242 (O_1242,N_14871,N_14928);
nand UO_1243 (O_1243,N_14895,N_14947);
or UO_1244 (O_1244,N_14936,N_14851);
nor UO_1245 (O_1245,N_14898,N_14957);
nand UO_1246 (O_1246,N_14968,N_14951);
nand UO_1247 (O_1247,N_14957,N_14958);
nor UO_1248 (O_1248,N_14988,N_14916);
nand UO_1249 (O_1249,N_14969,N_14980);
nand UO_1250 (O_1250,N_14876,N_14863);
or UO_1251 (O_1251,N_14869,N_14974);
nor UO_1252 (O_1252,N_14942,N_14909);
and UO_1253 (O_1253,N_14851,N_14866);
xnor UO_1254 (O_1254,N_14944,N_14996);
nand UO_1255 (O_1255,N_14973,N_14966);
xor UO_1256 (O_1256,N_14976,N_14855);
nor UO_1257 (O_1257,N_14957,N_14891);
and UO_1258 (O_1258,N_14905,N_14875);
and UO_1259 (O_1259,N_14904,N_14927);
nor UO_1260 (O_1260,N_14993,N_14959);
nor UO_1261 (O_1261,N_14916,N_14930);
nor UO_1262 (O_1262,N_14932,N_14973);
or UO_1263 (O_1263,N_14937,N_14910);
xnor UO_1264 (O_1264,N_14918,N_14869);
and UO_1265 (O_1265,N_14945,N_14859);
nand UO_1266 (O_1266,N_14861,N_14955);
nand UO_1267 (O_1267,N_14991,N_14951);
nor UO_1268 (O_1268,N_14873,N_14888);
nor UO_1269 (O_1269,N_14887,N_14944);
nand UO_1270 (O_1270,N_14991,N_14949);
and UO_1271 (O_1271,N_14889,N_14944);
and UO_1272 (O_1272,N_14888,N_14875);
nor UO_1273 (O_1273,N_14958,N_14999);
or UO_1274 (O_1274,N_14871,N_14879);
and UO_1275 (O_1275,N_14917,N_14919);
nand UO_1276 (O_1276,N_14851,N_14870);
nor UO_1277 (O_1277,N_14959,N_14935);
and UO_1278 (O_1278,N_14851,N_14983);
and UO_1279 (O_1279,N_14919,N_14981);
nor UO_1280 (O_1280,N_14903,N_14883);
or UO_1281 (O_1281,N_14977,N_14878);
and UO_1282 (O_1282,N_14915,N_14954);
and UO_1283 (O_1283,N_14950,N_14991);
xor UO_1284 (O_1284,N_14872,N_14995);
nor UO_1285 (O_1285,N_14958,N_14977);
xnor UO_1286 (O_1286,N_14889,N_14865);
and UO_1287 (O_1287,N_14940,N_14935);
nor UO_1288 (O_1288,N_14922,N_14927);
or UO_1289 (O_1289,N_14918,N_14853);
or UO_1290 (O_1290,N_14853,N_14881);
xnor UO_1291 (O_1291,N_14936,N_14970);
and UO_1292 (O_1292,N_14853,N_14976);
or UO_1293 (O_1293,N_14863,N_14959);
nor UO_1294 (O_1294,N_14957,N_14919);
nor UO_1295 (O_1295,N_14919,N_14937);
or UO_1296 (O_1296,N_14959,N_14913);
or UO_1297 (O_1297,N_14944,N_14918);
nor UO_1298 (O_1298,N_14918,N_14977);
xnor UO_1299 (O_1299,N_14914,N_14995);
or UO_1300 (O_1300,N_14937,N_14873);
or UO_1301 (O_1301,N_14957,N_14977);
and UO_1302 (O_1302,N_14874,N_14975);
nand UO_1303 (O_1303,N_14988,N_14918);
nor UO_1304 (O_1304,N_14872,N_14912);
or UO_1305 (O_1305,N_14874,N_14875);
nand UO_1306 (O_1306,N_14888,N_14988);
or UO_1307 (O_1307,N_14900,N_14963);
or UO_1308 (O_1308,N_14881,N_14897);
and UO_1309 (O_1309,N_14896,N_14939);
or UO_1310 (O_1310,N_14917,N_14970);
xor UO_1311 (O_1311,N_14969,N_14864);
nand UO_1312 (O_1312,N_14986,N_14863);
xnor UO_1313 (O_1313,N_14906,N_14910);
xor UO_1314 (O_1314,N_14971,N_14970);
and UO_1315 (O_1315,N_14872,N_14998);
xnor UO_1316 (O_1316,N_14867,N_14998);
nor UO_1317 (O_1317,N_14978,N_14854);
xor UO_1318 (O_1318,N_14907,N_14950);
nand UO_1319 (O_1319,N_14923,N_14976);
nor UO_1320 (O_1320,N_14867,N_14986);
and UO_1321 (O_1321,N_14975,N_14871);
nand UO_1322 (O_1322,N_14912,N_14934);
xnor UO_1323 (O_1323,N_14983,N_14955);
or UO_1324 (O_1324,N_14933,N_14861);
xor UO_1325 (O_1325,N_14851,N_14958);
nand UO_1326 (O_1326,N_14916,N_14860);
and UO_1327 (O_1327,N_14905,N_14966);
nor UO_1328 (O_1328,N_14983,N_14980);
nand UO_1329 (O_1329,N_14866,N_14962);
nor UO_1330 (O_1330,N_14993,N_14904);
and UO_1331 (O_1331,N_14925,N_14929);
nor UO_1332 (O_1332,N_14893,N_14978);
or UO_1333 (O_1333,N_14891,N_14898);
and UO_1334 (O_1334,N_14881,N_14961);
nand UO_1335 (O_1335,N_14990,N_14972);
and UO_1336 (O_1336,N_14881,N_14900);
and UO_1337 (O_1337,N_14865,N_14868);
nand UO_1338 (O_1338,N_14955,N_14999);
and UO_1339 (O_1339,N_14875,N_14961);
xor UO_1340 (O_1340,N_14932,N_14915);
or UO_1341 (O_1341,N_14988,N_14950);
nor UO_1342 (O_1342,N_14907,N_14898);
and UO_1343 (O_1343,N_14968,N_14877);
xor UO_1344 (O_1344,N_14991,N_14984);
nor UO_1345 (O_1345,N_14872,N_14857);
xor UO_1346 (O_1346,N_14927,N_14935);
and UO_1347 (O_1347,N_14962,N_14946);
nand UO_1348 (O_1348,N_14992,N_14930);
or UO_1349 (O_1349,N_14910,N_14871);
nand UO_1350 (O_1350,N_14915,N_14922);
xnor UO_1351 (O_1351,N_14905,N_14863);
nand UO_1352 (O_1352,N_14894,N_14965);
nor UO_1353 (O_1353,N_14897,N_14939);
and UO_1354 (O_1354,N_14996,N_14858);
or UO_1355 (O_1355,N_14997,N_14996);
or UO_1356 (O_1356,N_14922,N_14904);
nor UO_1357 (O_1357,N_14872,N_14974);
and UO_1358 (O_1358,N_14934,N_14936);
xor UO_1359 (O_1359,N_14921,N_14876);
nand UO_1360 (O_1360,N_14850,N_14933);
nor UO_1361 (O_1361,N_14897,N_14865);
nand UO_1362 (O_1362,N_14874,N_14885);
and UO_1363 (O_1363,N_14918,N_14870);
and UO_1364 (O_1364,N_14894,N_14936);
or UO_1365 (O_1365,N_14900,N_14899);
and UO_1366 (O_1366,N_14960,N_14902);
or UO_1367 (O_1367,N_14981,N_14875);
nor UO_1368 (O_1368,N_14924,N_14865);
nor UO_1369 (O_1369,N_14873,N_14956);
or UO_1370 (O_1370,N_14954,N_14873);
nand UO_1371 (O_1371,N_14930,N_14889);
or UO_1372 (O_1372,N_14929,N_14972);
xnor UO_1373 (O_1373,N_14884,N_14866);
nand UO_1374 (O_1374,N_14951,N_14870);
or UO_1375 (O_1375,N_14919,N_14907);
and UO_1376 (O_1376,N_14916,N_14959);
and UO_1377 (O_1377,N_14856,N_14880);
xor UO_1378 (O_1378,N_14896,N_14944);
xnor UO_1379 (O_1379,N_14905,N_14931);
nand UO_1380 (O_1380,N_14959,N_14856);
or UO_1381 (O_1381,N_14978,N_14885);
and UO_1382 (O_1382,N_14980,N_14920);
nand UO_1383 (O_1383,N_14906,N_14983);
xnor UO_1384 (O_1384,N_14954,N_14998);
nand UO_1385 (O_1385,N_14919,N_14877);
xnor UO_1386 (O_1386,N_14958,N_14909);
nand UO_1387 (O_1387,N_14968,N_14899);
xor UO_1388 (O_1388,N_14868,N_14965);
or UO_1389 (O_1389,N_14964,N_14907);
nand UO_1390 (O_1390,N_14981,N_14985);
nand UO_1391 (O_1391,N_14891,N_14864);
or UO_1392 (O_1392,N_14950,N_14925);
xnor UO_1393 (O_1393,N_14889,N_14901);
and UO_1394 (O_1394,N_14914,N_14966);
nand UO_1395 (O_1395,N_14912,N_14885);
nand UO_1396 (O_1396,N_14970,N_14919);
xor UO_1397 (O_1397,N_14887,N_14867);
nor UO_1398 (O_1398,N_14873,N_14902);
nand UO_1399 (O_1399,N_14970,N_14909);
nand UO_1400 (O_1400,N_14973,N_14919);
nand UO_1401 (O_1401,N_14968,N_14894);
nor UO_1402 (O_1402,N_14929,N_14901);
and UO_1403 (O_1403,N_14924,N_14995);
nor UO_1404 (O_1404,N_14953,N_14935);
xnor UO_1405 (O_1405,N_14916,N_14907);
nor UO_1406 (O_1406,N_14973,N_14867);
or UO_1407 (O_1407,N_14994,N_14914);
nor UO_1408 (O_1408,N_14886,N_14950);
nand UO_1409 (O_1409,N_14947,N_14888);
nor UO_1410 (O_1410,N_14944,N_14985);
xor UO_1411 (O_1411,N_14990,N_14956);
or UO_1412 (O_1412,N_14866,N_14984);
and UO_1413 (O_1413,N_14982,N_14889);
or UO_1414 (O_1414,N_14898,N_14943);
or UO_1415 (O_1415,N_14890,N_14926);
xor UO_1416 (O_1416,N_14980,N_14915);
nor UO_1417 (O_1417,N_14854,N_14933);
and UO_1418 (O_1418,N_14932,N_14955);
and UO_1419 (O_1419,N_14881,N_14906);
and UO_1420 (O_1420,N_14851,N_14916);
and UO_1421 (O_1421,N_14968,N_14901);
or UO_1422 (O_1422,N_14947,N_14887);
xor UO_1423 (O_1423,N_14992,N_14856);
nand UO_1424 (O_1424,N_14929,N_14857);
and UO_1425 (O_1425,N_14855,N_14889);
nand UO_1426 (O_1426,N_14903,N_14924);
xor UO_1427 (O_1427,N_14861,N_14888);
or UO_1428 (O_1428,N_14996,N_14860);
or UO_1429 (O_1429,N_14966,N_14955);
and UO_1430 (O_1430,N_14901,N_14978);
xnor UO_1431 (O_1431,N_14939,N_14958);
nor UO_1432 (O_1432,N_14904,N_14880);
and UO_1433 (O_1433,N_14989,N_14890);
or UO_1434 (O_1434,N_14887,N_14961);
and UO_1435 (O_1435,N_14958,N_14882);
nand UO_1436 (O_1436,N_14914,N_14965);
or UO_1437 (O_1437,N_14901,N_14851);
nand UO_1438 (O_1438,N_14903,N_14964);
or UO_1439 (O_1439,N_14885,N_14899);
nor UO_1440 (O_1440,N_14966,N_14892);
or UO_1441 (O_1441,N_14980,N_14944);
or UO_1442 (O_1442,N_14901,N_14931);
nand UO_1443 (O_1443,N_14945,N_14946);
nand UO_1444 (O_1444,N_14947,N_14963);
or UO_1445 (O_1445,N_14895,N_14980);
nor UO_1446 (O_1446,N_14927,N_14920);
and UO_1447 (O_1447,N_14868,N_14910);
nand UO_1448 (O_1448,N_14990,N_14993);
xnor UO_1449 (O_1449,N_14908,N_14857);
and UO_1450 (O_1450,N_14914,N_14880);
or UO_1451 (O_1451,N_14942,N_14903);
nand UO_1452 (O_1452,N_14931,N_14895);
and UO_1453 (O_1453,N_14873,N_14878);
nor UO_1454 (O_1454,N_14890,N_14993);
and UO_1455 (O_1455,N_14862,N_14922);
xnor UO_1456 (O_1456,N_14979,N_14983);
xnor UO_1457 (O_1457,N_14916,N_14960);
nor UO_1458 (O_1458,N_14903,N_14867);
nand UO_1459 (O_1459,N_14910,N_14969);
nor UO_1460 (O_1460,N_14922,N_14959);
nand UO_1461 (O_1461,N_14951,N_14863);
xnor UO_1462 (O_1462,N_14887,N_14917);
nand UO_1463 (O_1463,N_14905,N_14933);
or UO_1464 (O_1464,N_14981,N_14935);
or UO_1465 (O_1465,N_14972,N_14861);
and UO_1466 (O_1466,N_14902,N_14875);
xnor UO_1467 (O_1467,N_14868,N_14994);
and UO_1468 (O_1468,N_14854,N_14870);
xor UO_1469 (O_1469,N_14883,N_14852);
nor UO_1470 (O_1470,N_14884,N_14982);
nor UO_1471 (O_1471,N_14963,N_14920);
and UO_1472 (O_1472,N_14887,N_14870);
nor UO_1473 (O_1473,N_14931,N_14929);
nor UO_1474 (O_1474,N_14877,N_14944);
xnor UO_1475 (O_1475,N_14951,N_14924);
or UO_1476 (O_1476,N_14906,N_14950);
xnor UO_1477 (O_1477,N_14959,N_14931);
or UO_1478 (O_1478,N_14861,N_14947);
xor UO_1479 (O_1479,N_14871,N_14968);
nor UO_1480 (O_1480,N_14908,N_14854);
xor UO_1481 (O_1481,N_14961,N_14937);
nand UO_1482 (O_1482,N_14858,N_14870);
nor UO_1483 (O_1483,N_14884,N_14941);
xor UO_1484 (O_1484,N_14908,N_14863);
xnor UO_1485 (O_1485,N_14921,N_14998);
nand UO_1486 (O_1486,N_14895,N_14933);
nand UO_1487 (O_1487,N_14915,N_14982);
xnor UO_1488 (O_1488,N_14913,N_14922);
or UO_1489 (O_1489,N_14913,N_14981);
and UO_1490 (O_1490,N_14975,N_14954);
nand UO_1491 (O_1491,N_14961,N_14945);
nand UO_1492 (O_1492,N_14881,N_14943);
xnor UO_1493 (O_1493,N_14948,N_14970);
nor UO_1494 (O_1494,N_14944,N_14855);
nor UO_1495 (O_1495,N_14915,N_14956);
nor UO_1496 (O_1496,N_14952,N_14935);
nor UO_1497 (O_1497,N_14882,N_14913);
nand UO_1498 (O_1498,N_14963,N_14909);
nor UO_1499 (O_1499,N_14859,N_14923);
nor UO_1500 (O_1500,N_14987,N_14857);
or UO_1501 (O_1501,N_14888,N_14960);
or UO_1502 (O_1502,N_14915,N_14967);
nand UO_1503 (O_1503,N_14924,N_14940);
xnor UO_1504 (O_1504,N_14950,N_14940);
xnor UO_1505 (O_1505,N_14876,N_14965);
and UO_1506 (O_1506,N_14851,N_14982);
nor UO_1507 (O_1507,N_14954,N_14898);
or UO_1508 (O_1508,N_14876,N_14855);
xor UO_1509 (O_1509,N_14930,N_14963);
or UO_1510 (O_1510,N_14969,N_14869);
xnor UO_1511 (O_1511,N_14934,N_14890);
nand UO_1512 (O_1512,N_14855,N_14972);
or UO_1513 (O_1513,N_14953,N_14853);
nor UO_1514 (O_1514,N_14923,N_14881);
nand UO_1515 (O_1515,N_14907,N_14979);
nand UO_1516 (O_1516,N_14997,N_14909);
nand UO_1517 (O_1517,N_14991,N_14929);
or UO_1518 (O_1518,N_14887,N_14858);
nand UO_1519 (O_1519,N_14952,N_14929);
and UO_1520 (O_1520,N_14915,N_14887);
nor UO_1521 (O_1521,N_14921,N_14866);
nand UO_1522 (O_1522,N_14939,N_14959);
or UO_1523 (O_1523,N_14966,N_14909);
or UO_1524 (O_1524,N_14971,N_14870);
and UO_1525 (O_1525,N_14980,N_14953);
nor UO_1526 (O_1526,N_14934,N_14918);
xnor UO_1527 (O_1527,N_14872,N_14881);
or UO_1528 (O_1528,N_14924,N_14911);
nand UO_1529 (O_1529,N_14898,N_14860);
or UO_1530 (O_1530,N_14982,N_14904);
nand UO_1531 (O_1531,N_14998,N_14919);
and UO_1532 (O_1532,N_14911,N_14957);
nor UO_1533 (O_1533,N_14923,N_14852);
xor UO_1534 (O_1534,N_14958,N_14951);
or UO_1535 (O_1535,N_14995,N_14917);
or UO_1536 (O_1536,N_14894,N_14974);
nor UO_1537 (O_1537,N_14884,N_14947);
xor UO_1538 (O_1538,N_14917,N_14974);
or UO_1539 (O_1539,N_14920,N_14937);
nor UO_1540 (O_1540,N_14886,N_14854);
nand UO_1541 (O_1541,N_14968,N_14973);
nor UO_1542 (O_1542,N_14901,N_14981);
xnor UO_1543 (O_1543,N_14867,N_14862);
xor UO_1544 (O_1544,N_14951,N_14986);
nor UO_1545 (O_1545,N_14979,N_14888);
xor UO_1546 (O_1546,N_14960,N_14889);
nor UO_1547 (O_1547,N_14880,N_14971);
and UO_1548 (O_1548,N_14923,N_14882);
and UO_1549 (O_1549,N_14912,N_14883);
nor UO_1550 (O_1550,N_14962,N_14867);
nand UO_1551 (O_1551,N_14965,N_14987);
nor UO_1552 (O_1552,N_14947,N_14960);
xnor UO_1553 (O_1553,N_14863,N_14968);
or UO_1554 (O_1554,N_14868,N_14911);
and UO_1555 (O_1555,N_14857,N_14984);
and UO_1556 (O_1556,N_14955,N_14970);
xnor UO_1557 (O_1557,N_14931,N_14996);
and UO_1558 (O_1558,N_14930,N_14890);
xnor UO_1559 (O_1559,N_14870,N_14890);
and UO_1560 (O_1560,N_14978,N_14993);
or UO_1561 (O_1561,N_14852,N_14964);
and UO_1562 (O_1562,N_14867,N_14875);
nand UO_1563 (O_1563,N_14857,N_14894);
xnor UO_1564 (O_1564,N_14941,N_14856);
xor UO_1565 (O_1565,N_14860,N_14930);
and UO_1566 (O_1566,N_14998,N_14937);
or UO_1567 (O_1567,N_14980,N_14918);
or UO_1568 (O_1568,N_14885,N_14915);
and UO_1569 (O_1569,N_14901,N_14882);
or UO_1570 (O_1570,N_14851,N_14879);
and UO_1571 (O_1571,N_14909,N_14883);
xnor UO_1572 (O_1572,N_14924,N_14882);
or UO_1573 (O_1573,N_14962,N_14966);
or UO_1574 (O_1574,N_14851,N_14906);
xor UO_1575 (O_1575,N_14988,N_14858);
nor UO_1576 (O_1576,N_14871,N_14856);
and UO_1577 (O_1577,N_14922,N_14996);
xor UO_1578 (O_1578,N_14872,N_14961);
xor UO_1579 (O_1579,N_14939,N_14862);
nor UO_1580 (O_1580,N_14924,N_14997);
or UO_1581 (O_1581,N_14947,N_14879);
and UO_1582 (O_1582,N_14963,N_14858);
or UO_1583 (O_1583,N_14988,N_14889);
or UO_1584 (O_1584,N_14854,N_14939);
nand UO_1585 (O_1585,N_14916,N_14993);
and UO_1586 (O_1586,N_14938,N_14900);
or UO_1587 (O_1587,N_14910,N_14900);
nor UO_1588 (O_1588,N_14943,N_14868);
and UO_1589 (O_1589,N_14960,N_14872);
xor UO_1590 (O_1590,N_14871,N_14914);
nand UO_1591 (O_1591,N_14922,N_14951);
xnor UO_1592 (O_1592,N_14970,N_14935);
and UO_1593 (O_1593,N_14853,N_14872);
and UO_1594 (O_1594,N_14861,N_14870);
nor UO_1595 (O_1595,N_14984,N_14861);
nand UO_1596 (O_1596,N_14950,N_14857);
xor UO_1597 (O_1597,N_14912,N_14948);
xnor UO_1598 (O_1598,N_14883,N_14879);
or UO_1599 (O_1599,N_14947,N_14915);
nand UO_1600 (O_1600,N_14991,N_14952);
nand UO_1601 (O_1601,N_14991,N_14955);
or UO_1602 (O_1602,N_14975,N_14873);
and UO_1603 (O_1603,N_14855,N_14979);
or UO_1604 (O_1604,N_14909,N_14893);
nand UO_1605 (O_1605,N_14968,N_14954);
nand UO_1606 (O_1606,N_14971,N_14877);
nor UO_1607 (O_1607,N_14958,N_14989);
or UO_1608 (O_1608,N_14888,N_14936);
or UO_1609 (O_1609,N_14867,N_14889);
nand UO_1610 (O_1610,N_14876,N_14918);
xor UO_1611 (O_1611,N_14943,N_14993);
nand UO_1612 (O_1612,N_14891,N_14884);
nand UO_1613 (O_1613,N_14956,N_14976);
nor UO_1614 (O_1614,N_14883,N_14875);
nand UO_1615 (O_1615,N_14937,N_14898);
nand UO_1616 (O_1616,N_14912,N_14871);
or UO_1617 (O_1617,N_14853,N_14866);
or UO_1618 (O_1618,N_14958,N_14891);
nor UO_1619 (O_1619,N_14920,N_14854);
xor UO_1620 (O_1620,N_14883,N_14942);
xnor UO_1621 (O_1621,N_14966,N_14977);
xor UO_1622 (O_1622,N_14995,N_14925);
and UO_1623 (O_1623,N_14954,N_14911);
nor UO_1624 (O_1624,N_14926,N_14864);
or UO_1625 (O_1625,N_14851,N_14952);
nor UO_1626 (O_1626,N_14999,N_14934);
or UO_1627 (O_1627,N_14884,N_14994);
and UO_1628 (O_1628,N_14892,N_14921);
xnor UO_1629 (O_1629,N_14997,N_14962);
xor UO_1630 (O_1630,N_14972,N_14950);
and UO_1631 (O_1631,N_14919,N_14879);
xor UO_1632 (O_1632,N_14880,N_14870);
or UO_1633 (O_1633,N_14973,N_14888);
or UO_1634 (O_1634,N_14965,N_14908);
or UO_1635 (O_1635,N_14867,N_14865);
or UO_1636 (O_1636,N_14920,N_14998);
nand UO_1637 (O_1637,N_14925,N_14977);
or UO_1638 (O_1638,N_14946,N_14886);
nand UO_1639 (O_1639,N_14953,N_14963);
xor UO_1640 (O_1640,N_14957,N_14976);
and UO_1641 (O_1641,N_14896,N_14918);
nand UO_1642 (O_1642,N_14851,N_14909);
nand UO_1643 (O_1643,N_14877,N_14886);
and UO_1644 (O_1644,N_14952,N_14953);
or UO_1645 (O_1645,N_14878,N_14963);
nand UO_1646 (O_1646,N_14988,N_14885);
and UO_1647 (O_1647,N_14875,N_14901);
nor UO_1648 (O_1648,N_14993,N_14911);
nand UO_1649 (O_1649,N_14911,N_14945);
nand UO_1650 (O_1650,N_14851,N_14993);
nor UO_1651 (O_1651,N_14918,N_14874);
nand UO_1652 (O_1652,N_14875,N_14927);
xor UO_1653 (O_1653,N_14942,N_14962);
nor UO_1654 (O_1654,N_14969,N_14933);
nand UO_1655 (O_1655,N_14970,N_14982);
and UO_1656 (O_1656,N_14895,N_14989);
nand UO_1657 (O_1657,N_14974,N_14931);
or UO_1658 (O_1658,N_14873,N_14919);
nor UO_1659 (O_1659,N_14889,N_14965);
nor UO_1660 (O_1660,N_14875,N_14958);
and UO_1661 (O_1661,N_14920,N_14999);
and UO_1662 (O_1662,N_14991,N_14853);
and UO_1663 (O_1663,N_14924,N_14968);
nor UO_1664 (O_1664,N_14903,N_14856);
and UO_1665 (O_1665,N_14965,N_14861);
nor UO_1666 (O_1666,N_14926,N_14882);
nand UO_1667 (O_1667,N_14893,N_14950);
nor UO_1668 (O_1668,N_14927,N_14995);
or UO_1669 (O_1669,N_14906,N_14979);
xnor UO_1670 (O_1670,N_14945,N_14968);
or UO_1671 (O_1671,N_14902,N_14981);
or UO_1672 (O_1672,N_14917,N_14981);
xnor UO_1673 (O_1673,N_14852,N_14853);
or UO_1674 (O_1674,N_14858,N_14859);
nor UO_1675 (O_1675,N_14872,N_14911);
or UO_1676 (O_1676,N_14895,N_14940);
nand UO_1677 (O_1677,N_14977,N_14997);
or UO_1678 (O_1678,N_14998,N_14930);
or UO_1679 (O_1679,N_14945,N_14864);
or UO_1680 (O_1680,N_14922,N_14874);
nand UO_1681 (O_1681,N_14940,N_14884);
xnor UO_1682 (O_1682,N_14860,N_14977);
and UO_1683 (O_1683,N_14977,N_14874);
and UO_1684 (O_1684,N_14954,N_14999);
nand UO_1685 (O_1685,N_14944,N_14967);
xnor UO_1686 (O_1686,N_14950,N_14926);
and UO_1687 (O_1687,N_14998,N_14936);
nor UO_1688 (O_1688,N_14983,N_14985);
or UO_1689 (O_1689,N_14880,N_14891);
xor UO_1690 (O_1690,N_14935,N_14888);
nor UO_1691 (O_1691,N_14945,N_14896);
and UO_1692 (O_1692,N_14999,N_14937);
and UO_1693 (O_1693,N_14857,N_14900);
nor UO_1694 (O_1694,N_14926,N_14967);
nor UO_1695 (O_1695,N_14992,N_14918);
and UO_1696 (O_1696,N_14851,N_14854);
nand UO_1697 (O_1697,N_14895,N_14952);
or UO_1698 (O_1698,N_14864,N_14959);
nor UO_1699 (O_1699,N_14858,N_14992);
xnor UO_1700 (O_1700,N_14912,N_14966);
or UO_1701 (O_1701,N_14951,N_14967);
nand UO_1702 (O_1702,N_14913,N_14945);
nor UO_1703 (O_1703,N_14883,N_14937);
nor UO_1704 (O_1704,N_14996,N_14927);
xnor UO_1705 (O_1705,N_14885,N_14862);
xor UO_1706 (O_1706,N_14974,N_14928);
and UO_1707 (O_1707,N_14923,N_14905);
nor UO_1708 (O_1708,N_14865,N_14950);
and UO_1709 (O_1709,N_14933,N_14915);
nor UO_1710 (O_1710,N_14903,N_14874);
nor UO_1711 (O_1711,N_14898,N_14861);
nor UO_1712 (O_1712,N_14986,N_14910);
nand UO_1713 (O_1713,N_14858,N_14914);
nand UO_1714 (O_1714,N_14888,N_14886);
or UO_1715 (O_1715,N_14990,N_14866);
and UO_1716 (O_1716,N_14933,N_14867);
xnor UO_1717 (O_1717,N_14963,N_14977);
nor UO_1718 (O_1718,N_14951,N_14893);
xor UO_1719 (O_1719,N_14942,N_14866);
and UO_1720 (O_1720,N_14949,N_14996);
nor UO_1721 (O_1721,N_14850,N_14976);
nor UO_1722 (O_1722,N_14907,N_14936);
or UO_1723 (O_1723,N_14994,N_14923);
and UO_1724 (O_1724,N_14965,N_14925);
xor UO_1725 (O_1725,N_14979,N_14900);
nor UO_1726 (O_1726,N_14924,N_14906);
nor UO_1727 (O_1727,N_14861,N_14913);
nand UO_1728 (O_1728,N_14920,N_14964);
nor UO_1729 (O_1729,N_14894,N_14927);
or UO_1730 (O_1730,N_14997,N_14859);
xnor UO_1731 (O_1731,N_14984,N_14989);
nor UO_1732 (O_1732,N_14889,N_14946);
xor UO_1733 (O_1733,N_14926,N_14954);
xor UO_1734 (O_1734,N_14919,N_14972);
xnor UO_1735 (O_1735,N_14909,N_14930);
xor UO_1736 (O_1736,N_14927,N_14879);
xnor UO_1737 (O_1737,N_14937,N_14939);
and UO_1738 (O_1738,N_14854,N_14860);
nand UO_1739 (O_1739,N_14967,N_14884);
and UO_1740 (O_1740,N_14903,N_14935);
nand UO_1741 (O_1741,N_14956,N_14917);
nand UO_1742 (O_1742,N_14917,N_14862);
and UO_1743 (O_1743,N_14931,N_14900);
or UO_1744 (O_1744,N_14872,N_14906);
or UO_1745 (O_1745,N_14879,N_14908);
and UO_1746 (O_1746,N_14952,N_14939);
xnor UO_1747 (O_1747,N_14883,N_14910);
and UO_1748 (O_1748,N_14971,N_14974);
or UO_1749 (O_1749,N_14913,N_14958);
and UO_1750 (O_1750,N_14997,N_14945);
nand UO_1751 (O_1751,N_14932,N_14926);
or UO_1752 (O_1752,N_14893,N_14857);
nand UO_1753 (O_1753,N_14971,N_14889);
nor UO_1754 (O_1754,N_14993,N_14940);
or UO_1755 (O_1755,N_14925,N_14992);
or UO_1756 (O_1756,N_14922,N_14999);
and UO_1757 (O_1757,N_14921,N_14880);
nand UO_1758 (O_1758,N_14924,N_14964);
or UO_1759 (O_1759,N_14852,N_14891);
or UO_1760 (O_1760,N_14899,N_14895);
or UO_1761 (O_1761,N_14871,N_14895);
xor UO_1762 (O_1762,N_14895,N_14894);
and UO_1763 (O_1763,N_14864,N_14964);
nor UO_1764 (O_1764,N_14912,N_14973);
or UO_1765 (O_1765,N_14935,N_14892);
or UO_1766 (O_1766,N_14931,N_14994);
or UO_1767 (O_1767,N_14913,N_14878);
or UO_1768 (O_1768,N_14926,N_14852);
xnor UO_1769 (O_1769,N_14886,N_14865);
nor UO_1770 (O_1770,N_14949,N_14947);
xnor UO_1771 (O_1771,N_14998,N_14960);
or UO_1772 (O_1772,N_14949,N_14924);
nor UO_1773 (O_1773,N_14950,N_14942);
nand UO_1774 (O_1774,N_14903,N_14977);
or UO_1775 (O_1775,N_14924,N_14915);
nand UO_1776 (O_1776,N_14934,N_14969);
nor UO_1777 (O_1777,N_14901,N_14871);
xor UO_1778 (O_1778,N_14973,N_14901);
nor UO_1779 (O_1779,N_14891,N_14862);
or UO_1780 (O_1780,N_14884,N_14905);
xnor UO_1781 (O_1781,N_14923,N_14951);
and UO_1782 (O_1782,N_14956,N_14889);
xor UO_1783 (O_1783,N_14991,N_14903);
nand UO_1784 (O_1784,N_14963,N_14890);
and UO_1785 (O_1785,N_14883,N_14911);
and UO_1786 (O_1786,N_14895,N_14898);
xor UO_1787 (O_1787,N_14999,N_14872);
nand UO_1788 (O_1788,N_14941,N_14927);
nor UO_1789 (O_1789,N_14878,N_14922);
nor UO_1790 (O_1790,N_14963,N_14982);
and UO_1791 (O_1791,N_14987,N_14866);
xnor UO_1792 (O_1792,N_14896,N_14923);
xor UO_1793 (O_1793,N_14940,N_14889);
nand UO_1794 (O_1794,N_14957,N_14980);
nor UO_1795 (O_1795,N_14972,N_14921);
xor UO_1796 (O_1796,N_14866,N_14878);
nor UO_1797 (O_1797,N_14947,N_14973);
or UO_1798 (O_1798,N_14938,N_14924);
or UO_1799 (O_1799,N_14967,N_14881);
nand UO_1800 (O_1800,N_14865,N_14942);
or UO_1801 (O_1801,N_14882,N_14900);
xnor UO_1802 (O_1802,N_14886,N_14951);
xnor UO_1803 (O_1803,N_14920,N_14974);
nor UO_1804 (O_1804,N_14894,N_14919);
xnor UO_1805 (O_1805,N_14881,N_14959);
nor UO_1806 (O_1806,N_14887,N_14970);
xor UO_1807 (O_1807,N_14994,N_14907);
and UO_1808 (O_1808,N_14995,N_14938);
or UO_1809 (O_1809,N_14954,N_14970);
nand UO_1810 (O_1810,N_14886,N_14928);
xnor UO_1811 (O_1811,N_14963,N_14935);
nor UO_1812 (O_1812,N_14890,N_14941);
and UO_1813 (O_1813,N_14987,N_14954);
and UO_1814 (O_1814,N_14972,N_14868);
nor UO_1815 (O_1815,N_14963,N_14949);
nor UO_1816 (O_1816,N_14941,N_14947);
xor UO_1817 (O_1817,N_14851,N_14975);
and UO_1818 (O_1818,N_14912,N_14930);
xor UO_1819 (O_1819,N_14886,N_14975);
nor UO_1820 (O_1820,N_14984,N_14922);
nand UO_1821 (O_1821,N_14956,N_14886);
or UO_1822 (O_1822,N_14925,N_14854);
xor UO_1823 (O_1823,N_14951,N_14854);
nor UO_1824 (O_1824,N_14858,N_14880);
nor UO_1825 (O_1825,N_14959,N_14995);
nand UO_1826 (O_1826,N_14873,N_14951);
or UO_1827 (O_1827,N_14862,N_14877);
nor UO_1828 (O_1828,N_14911,N_14885);
xnor UO_1829 (O_1829,N_14885,N_14910);
nor UO_1830 (O_1830,N_14973,N_14965);
xnor UO_1831 (O_1831,N_14907,N_14920);
or UO_1832 (O_1832,N_14971,N_14882);
and UO_1833 (O_1833,N_14921,N_14917);
xor UO_1834 (O_1834,N_14916,N_14980);
nand UO_1835 (O_1835,N_14993,N_14867);
nor UO_1836 (O_1836,N_14869,N_14912);
or UO_1837 (O_1837,N_14981,N_14904);
xnor UO_1838 (O_1838,N_14992,N_14851);
nor UO_1839 (O_1839,N_14923,N_14947);
or UO_1840 (O_1840,N_14966,N_14986);
nand UO_1841 (O_1841,N_14990,N_14855);
or UO_1842 (O_1842,N_14996,N_14979);
nor UO_1843 (O_1843,N_14857,N_14874);
and UO_1844 (O_1844,N_14962,N_14905);
xnor UO_1845 (O_1845,N_14869,N_14954);
or UO_1846 (O_1846,N_14945,N_14866);
or UO_1847 (O_1847,N_14998,N_14939);
xnor UO_1848 (O_1848,N_14974,N_14881);
nor UO_1849 (O_1849,N_14856,N_14926);
and UO_1850 (O_1850,N_14959,N_14944);
or UO_1851 (O_1851,N_14903,N_14855);
nor UO_1852 (O_1852,N_14989,N_14894);
or UO_1853 (O_1853,N_14915,N_14958);
nand UO_1854 (O_1854,N_14890,N_14876);
or UO_1855 (O_1855,N_14950,N_14948);
and UO_1856 (O_1856,N_14963,N_14922);
and UO_1857 (O_1857,N_14888,N_14912);
xnor UO_1858 (O_1858,N_14921,N_14951);
nor UO_1859 (O_1859,N_14943,N_14941);
and UO_1860 (O_1860,N_14990,N_14894);
and UO_1861 (O_1861,N_14883,N_14962);
nand UO_1862 (O_1862,N_14952,N_14968);
and UO_1863 (O_1863,N_14907,N_14951);
and UO_1864 (O_1864,N_14873,N_14950);
nand UO_1865 (O_1865,N_14974,N_14909);
nor UO_1866 (O_1866,N_14990,N_14881);
nor UO_1867 (O_1867,N_14913,N_14947);
nand UO_1868 (O_1868,N_14895,N_14986);
or UO_1869 (O_1869,N_14935,N_14934);
nand UO_1870 (O_1870,N_14935,N_14855);
and UO_1871 (O_1871,N_14890,N_14882);
nand UO_1872 (O_1872,N_14960,N_14968);
nor UO_1873 (O_1873,N_14923,N_14974);
nand UO_1874 (O_1874,N_14996,N_14879);
nor UO_1875 (O_1875,N_14982,N_14888);
xor UO_1876 (O_1876,N_14934,N_14984);
nand UO_1877 (O_1877,N_14909,N_14886);
xor UO_1878 (O_1878,N_14911,N_14852);
xor UO_1879 (O_1879,N_14992,N_14861);
nand UO_1880 (O_1880,N_14901,N_14951);
nand UO_1881 (O_1881,N_14903,N_14996);
and UO_1882 (O_1882,N_14945,N_14952);
nand UO_1883 (O_1883,N_14971,N_14990);
or UO_1884 (O_1884,N_14874,N_14924);
nor UO_1885 (O_1885,N_14920,N_14871);
nand UO_1886 (O_1886,N_14945,N_14853);
and UO_1887 (O_1887,N_14911,N_14915);
nand UO_1888 (O_1888,N_14996,N_14953);
and UO_1889 (O_1889,N_14876,N_14917);
xor UO_1890 (O_1890,N_14862,N_14902);
or UO_1891 (O_1891,N_14973,N_14929);
and UO_1892 (O_1892,N_14890,N_14959);
and UO_1893 (O_1893,N_14968,N_14862);
and UO_1894 (O_1894,N_14892,N_14889);
or UO_1895 (O_1895,N_14983,N_14883);
xnor UO_1896 (O_1896,N_14948,N_14954);
xnor UO_1897 (O_1897,N_14921,N_14883);
nor UO_1898 (O_1898,N_14852,N_14871);
or UO_1899 (O_1899,N_14896,N_14913);
or UO_1900 (O_1900,N_14979,N_14876);
nand UO_1901 (O_1901,N_14892,N_14863);
nand UO_1902 (O_1902,N_14994,N_14945);
xnor UO_1903 (O_1903,N_14919,N_14945);
xnor UO_1904 (O_1904,N_14931,N_14987);
and UO_1905 (O_1905,N_14964,N_14957);
nor UO_1906 (O_1906,N_14873,N_14997);
or UO_1907 (O_1907,N_14966,N_14868);
nor UO_1908 (O_1908,N_14938,N_14891);
xor UO_1909 (O_1909,N_14992,N_14988);
xor UO_1910 (O_1910,N_14988,N_14972);
xor UO_1911 (O_1911,N_14854,N_14859);
xor UO_1912 (O_1912,N_14982,N_14867);
or UO_1913 (O_1913,N_14914,N_14929);
or UO_1914 (O_1914,N_14909,N_14961);
or UO_1915 (O_1915,N_14994,N_14855);
or UO_1916 (O_1916,N_14910,N_14965);
or UO_1917 (O_1917,N_14995,N_14861);
nand UO_1918 (O_1918,N_14865,N_14861);
nand UO_1919 (O_1919,N_14933,N_14946);
nor UO_1920 (O_1920,N_14909,N_14906);
nand UO_1921 (O_1921,N_14920,N_14931);
and UO_1922 (O_1922,N_14940,N_14874);
nand UO_1923 (O_1923,N_14978,N_14879);
and UO_1924 (O_1924,N_14874,N_14982);
nand UO_1925 (O_1925,N_14944,N_14987);
and UO_1926 (O_1926,N_14992,N_14942);
and UO_1927 (O_1927,N_14869,N_14925);
xor UO_1928 (O_1928,N_14950,N_14980);
or UO_1929 (O_1929,N_14921,N_14947);
and UO_1930 (O_1930,N_14934,N_14941);
and UO_1931 (O_1931,N_14876,N_14925);
nand UO_1932 (O_1932,N_14994,N_14905);
nor UO_1933 (O_1933,N_14944,N_14971);
nor UO_1934 (O_1934,N_14993,N_14989);
nor UO_1935 (O_1935,N_14956,N_14953);
xor UO_1936 (O_1936,N_14934,N_14916);
nor UO_1937 (O_1937,N_14940,N_14910);
nand UO_1938 (O_1938,N_14891,N_14903);
nand UO_1939 (O_1939,N_14973,N_14859);
and UO_1940 (O_1940,N_14859,N_14946);
and UO_1941 (O_1941,N_14934,N_14958);
nand UO_1942 (O_1942,N_14862,N_14919);
xor UO_1943 (O_1943,N_14907,N_14906);
xnor UO_1944 (O_1944,N_14992,N_14874);
nand UO_1945 (O_1945,N_14931,N_14947);
xnor UO_1946 (O_1946,N_14864,N_14941);
nor UO_1947 (O_1947,N_14955,N_14998);
and UO_1948 (O_1948,N_14899,N_14896);
nand UO_1949 (O_1949,N_14921,N_14927);
nor UO_1950 (O_1950,N_14979,N_14936);
nor UO_1951 (O_1951,N_14971,N_14858);
and UO_1952 (O_1952,N_14858,N_14999);
or UO_1953 (O_1953,N_14943,N_14894);
nor UO_1954 (O_1954,N_14917,N_14932);
nand UO_1955 (O_1955,N_14945,N_14885);
and UO_1956 (O_1956,N_14907,N_14980);
xnor UO_1957 (O_1957,N_14884,N_14910);
nand UO_1958 (O_1958,N_14876,N_14873);
or UO_1959 (O_1959,N_14888,N_14918);
nand UO_1960 (O_1960,N_14989,N_14921);
nand UO_1961 (O_1961,N_14964,N_14975);
and UO_1962 (O_1962,N_14907,N_14892);
nor UO_1963 (O_1963,N_14952,N_14993);
xor UO_1964 (O_1964,N_14866,N_14930);
nand UO_1965 (O_1965,N_14996,N_14861);
xor UO_1966 (O_1966,N_14908,N_14874);
nand UO_1967 (O_1967,N_14986,N_14942);
xnor UO_1968 (O_1968,N_14924,N_14921);
and UO_1969 (O_1969,N_14969,N_14966);
or UO_1970 (O_1970,N_14910,N_14916);
xnor UO_1971 (O_1971,N_14876,N_14957);
and UO_1972 (O_1972,N_14908,N_14998);
and UO_1973 (O_1973,N_14871,N_14887);
nand UO_1974 (O_1974,N_14979,N_14939);
and UO_1975 (O_1975,N_14988,N_14970);
xnor UO_1976 (O_1976,N_14982,N_14879);
and UO_1977 (O_1977,N_14976,N_14961);
nor UO_1978 (O_1978,N_14864,N_14937);
and UO_1979 (O_1979,N_14943,N_14942);
nand UO_1980 (O_1980,N_14935,N_14921);
nand UO_1981 (O_1981,N_14890,N_14984);
and UO_1982 (O_1982,N_14863,N_14919);
or UO_1983 (O_1983,N_14880,N_14935);
or UO_1984 (O_1984,N_14857,N_14873);
nor UO_1985 (O_1985,N_14928,N_14894);
and UO_1986 (O_1986,N_14981,N_14906);
nor UO_1987 (O_1987,N_14904,N_14964);
nand UO_1988 (O_1988,N_14915,N_14879);
and UO_1989 (O_1989,N_14915,N_14912);
nor UO_1990 (O_1990,N_14910,N_14863);
and UO_1991 (O_1991,N_14929,N_14897);
or UO_1992 (O_1992,N_14902,N_14921);
and UO_1993 (O_1993,N_14978,N_14889);
nand UO_1994 (O_1994,N_14884,N_14988);
or UO_1995 (O_1995,N_14995,N_14863);
xor UO_1996 (O_1996,N_14985,N_14908);
xnor UO_1997 (O_1997,N_14931,N_14860);
xor UO_1998 (O_1998,N_14977,N_14981);
and UO_1999 (O_1999,N_14941,N_14874);
endmodule