module basic_2000_20000_2500_20_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_413,In_580);
nand U1 (N_1,In_1936,In_145);
nor U2 (N_2,In_1281,In_943);
xnor U3 (N_3,In_1795,In_1084);
or U4 (N_4,In_82,In_45);
xor U5 (N_5,In_284,In_233);
xor U6 (N_6,In_271,In_887);
and U7 (N_7,In_1643,In_208);
or U8 (N_8,In_1240,In_1639);
and U9 (N_9,In_1482,In_1834);
or U10 (N_10,In_388,In_1431);
nand U11 (N_11,In_1940,In_1667);
nor U12 (N_12,In_1284,In_391);
nor U13 (N_13,In_1656,In_1621);
nand U14 (N_14,In_390,In_1833);
nand U15 (N_15,In_1011,In_1215);
xnor U16 (N_16,In_1417,In_544);
nor U17 (N_17,In_1471,In_44);
and U18 (N_18,In_541,In_482);
nand U19 (N_19,In_218,In_1190);
xnor U20 (N_20,In_748,In_1577);
nor U21 (N_21,In_1949,In_1370);
nand U22 (N_22,In_891,In_1919);
xor U23 (N_23,In_1758,In_1119);
nand U24 (N_24,In_1021,In_1477);
and U25 (N_25,In_1756,In_1313);
nor U26 (N_26,In_1699,In_1306);
nand U27 (N_27,In_357,In_1800);
xor U28 (N_28,In_1245,In_817);
nor U29 (N_29,In_1268,In_837);
nand U30 (N_30,In_20,In_1506);
or U31 (N_31,In_553,In_1596);
xor U32 (N_32,In_1874,In_1077);
or U33 (N_33,In_1124,In_1752);
xnor U34 (N_34,In_1972,In_1252);
nand U35 (N_35,In_1439,In_1899);
and U36 (N_36,In_59,In_1408);
or U37 (N_37,In_246,In_1052);
xnor U38 (N_38,In_40,In_66);
xnor U39 (N_39,In_1060,In_1200);
xor U40 (N_40,In_708,In_1869);
nand U41 (N_41,In_1279,In_336);
and U42 (N_42,In_221,In_285);
nor U43 (N_43,In_1427,In_344);
nand U44 (N_44,In_1681,In_124);
nor U45 (N_45,In_1135,In_899);
nor U46 (N_46,In_399,In_621);
nand U47 (N_47,In_1932,In_993);
nor U48 (N_48,In_113,In_1700);
or U49 (N_49,In_1340,In_868);
or U50 (N_50,In_1532,In_535);
nand U51 (N_51,In_1794,In_1314);
xor U52 (N_52,In_1958,In_1541);
or U53 (N_53,In_1520,In_610);
nand U54 (N_54,In_272,In_971);
nand U55 (N_55,In_1988,In_1887);
and U56 (N_56,In_1209,In_1322);
or U57 (N_57,In_1309,In_1548);
nor U58 (N_58,In_1538,In_1232);
nor U59 (N_59,In_297,In_230);
and U60 (N_60,In_649,In_1774);
and U61 (N_61,In_849,In_77);
nand U62 (N_62,In_873,In_633);
nor U63 (N_63,In_161,In_1065);
and U64 (N_64,In_127,In_1813);
and U65 (N_65,In_515,In_1104);
nor U66 (N_66,In_416,In_625);
or U67 (N_67,In_611,In_1922);
or U68 (N_68,In_779,In_1790);
nor U69 (N_69,In_1654,In_770);
or U70 (N_70,In_958,In_472);
or U71 (N_71,In_61,In_1285);
xnor U72 (N_72,In_1625,In_1273);
nand U73 (N_73,In_1838,In_1634);
or U74 (N_74,In_139,In_371);
xor U75 (N_75,In_1895,In_1177);
nor U76 (N_76,In_1264,In_63);
nand U77 (N_77,In_148,In_250);
or U78 (N_78,In_1057,In_1100);
and U79 (N_79,In_765,In_1705);
nor U80 (N_80,In_1751,In_1396);
or U81 (N_81,In_116,In_1341);
or U82 (N_82,In_893,In_119);
nand U83 (N_83,In_491,In_475);
or U84 (N_84,In_980,In_76);
nor U85 (N_85,In_790,In_33);
and U86 (N_86,In_653,In_1943);
nor U87 (N_87,In_108,In_128);
and U88 (N_88,In_30,In_1853);
or U89 (N_89,In_191,In_920);
nand U90 (N_90,In_353,In_1063);
xor U91 (N_91,In_955,In_16);
and U92 (N_92,In_402,In_478);
or U93 (N_93,In_500,In_841);
or U94 (N_94,In_165,In_314);
or U95 (N_95,In_1999,In_976);
or U96 (N_96,In_492,In_1201);
xor U97 (N_97,In_1875,In_1425);
and U98 (N_98,In_1684,In_1069);
nand U99 (N_99,In_1557,In_1331);
nand U100 (N_100,In_827,In_1113);
nand U101 (N_101,In_1632,In_859);
or U102 (N_102,In_700,In_1324);
nand U103 (N_103,In_1300,In_769);
nor U104 (N_104,In_115,In_641);
and U105 (N_105,In_1320,In_586);
and U106 (N_106,In_104,In_1615);
or U107 (N_107,In_38,In_1034);
or U108 (N_108,In_1402,In_1508);
nand U109 (N_109,In_100,In_1574);
nor U110 (N_110,In_407,In_1501);
or U111 (N_111,In_152,In_932);
nor U112 (N_112,In_1059,In_319);
nand U113 (N_113,In_957,In_617);
and U114 (N_114,In_1670,In_1918);
xnor U115 (N_115,In_28,In_4);
nor U116 (N_116,In_916,In_95);
xnor U117 (N_117,In_1224,In_669);
or U118 (N_118,In_1585,In_1525);
and U119 (N_119,In_741,In_941);
or U120 (N_120,In_660,In_1116);
nand U121 (N_121,In_311,In_522);
nand U122 (N_122,In_1765,In_1474);
nor U123 (N_123,In_898,In_1682);
or U124 (N_124,In_1792,In_676);
nor U125 (N_125,In_270,In_1952);
or U126 (N_126,In_711,In_895);
or U127 (N_127,In_1844,In_1469);
and U128 (N_128,In_1801,In_1005);
or U129 (N_129,In_1053,In_366);
nand U130 (N_130,In_1823,In_204);
and U131 (N_131,In_992,In_1769);
or U132 (N_132,In_141,In_1329);
nor U133 (N_133,In_620,In_810);
or U134 (N_134,In_1561,In_1154);
and U135 (N_135,In_731,In_456);
nand U136 (N_136,In_1207,In_1914);
or U137 (N_137,In_539,In_1444);
nor U138 (N_138,In_1981,In_1270);
xnor U139 (N_139,In_1205,In_1079);
xor U140 (N_140,In_1961,In_1421);
and U141 (N_141,In_1357,In_651);
nand U142 (N_142,In_1206,In_394);
nand U143 (N_143,In_650,In_1767);
or U144 (N_144,In_24,In_1848);
nor U145 (N_145,In_158,In_1360);
or U146 (N_146,In_328,In_195);
or U147 (N_147,In_334,In_292);
or U148 (N_148,In_1509,In_251);
and U149 (N_149,In_1570,In_93);
nor U150 (N_150,In_1,In_1301);
and U151 (N_151,In_836,In_933);
nor U152 (N_152,In_310,In_367);
nor U153 (N_153,In_1407,In_1707);
xor U154 (N_154,In_1088,In_1489);
and U155 (N_155,In_1435,In_961);
nand U156 (N_156,In_690,In_1158);
and U157 (N_157,In_231,In_1709);
nand U158 (N_158,In_1722,In_1911);
or U159 (N_159,In_1576,In_1990);
nand U160 (N_160,In_35,In_1120);
nor U161 (N_161,In_1250,In_1286);
or U162 (N_162,In_533,In_1092);
or U163 (N_163,In_1122,In_707);
and U164 (N_164,In_760,In_333);
nand U165 (N_165,In_1708,In_369);
nor U166 (N_166,In_1162,In_316);
nand U167 (N_167,In_1624,In_1455);
nand U168 (N_168,In_1980,In_126);
nor U169 (N_169,In_1864,In_1995);
and U170 (N_170,In_142,In_561);
nand U171 (N_171,In_1235,In_280);
nand U172 (N_172,In_1406,In_639);
and U173 (N_173,In_1371,In_1846);
and U174 (N_174,In_793,In_1013);
or U175 (N_175,In_928,In_1738);
and U176 (N_176,In_1609,In_1725);
or U177 (N_177,In_229,In_188);
and U178 (N_178,In_1544,In_480);
or U179 (N_179,In_1002,In_1663);
and U180 (N_180,In_1275,In_332);
nand U181 (N_181,In_1437,In_791);
xor U182 (N_182,In_10,In_466);
and U183 (N_183,In_1590,In_1677);
nor U184 (N_184,In_91,In_757);
nor U185 (N_185,In_1037,In_838);
and U186 (N_186,In_546,In_138);
and U187 (N_187,In_430,In_906);
or U188 (N_188,In_1377,In_697);
and U189 (N_189,In_1890,In_1132);
xor U190 (N_190,In_1825,In_293);
nand U191 (N_191,In_29,In_1636);
or U192 (N_192,In_1759,In_1802);
nor U193 (N_193,In_36,In_1165);
or U194 (N_194,In_1103,In_1083);
nor U195 (N_195,In_1989,In_684);
or U196 (N_196,In_1903,In_249);
and U197 (N_197,In_423,In_1698);
or U198 (N_198,In_1137,In_1645);
nand U199 (N_199,In_1798,In_245);
nand U200 (N_200,In_243,In_175);
nor U201 (N_201,In_418,In_308);
or U202 (N_202,In_1204,In_834);
or U203 (N_203,In_1770,In_947);
nor U204 (N_204,In_1464,In_1696);
or U205 (N_205,In_112,In_1829);
and U206 (N_206,In_1603,In_1236);
nand U207 (N_207,In_25,In_1522);
nand U208 (N_208,In_585,In_860);
and U209 (N_209,In_428,In_805);
and U210 (N_210,In_970,In_979);
nand U211 (N_211,In_798,In_1781);
or U212 (N_212,In_1893,In_737);
or U213 (N_213,In_260,In_234);
xor U214 (N_214,In_819,In_1025);
nand U215 (N_215,In_504,In_1026);
and U216 (N_216,In_443,In_1099);
and U217 (N_217,In_694,In_1977);
nor U218 (N_218,In_1287,In_1278);
or U219 (N_219,In_1657,In_733);
and U220 (N_220,In_1163,In_1046);
or U221 (N_221,In_612,In_1262);
nor U222 (N_222,In_839,In_1228);
nand U223 (N_223,In_160,In_1121);
nand U224 (N_224,In_454,In_1673);
nand U225 (N_225,In_1463,In_643);
and U226 (N_226,In_704,In_1889);
xnor U227 (N_227,In_1894,In_1367);
nand U228 (N_228,In_341,In_203);
and U229 (N_229,In_1014,In_393);
nor U230 (N_230,In_170,In_1880);
or U231 (N_231,In_1998,In_940);
or U232 (N_232,In_1420,In_845);
nand U233 (N_233,In_52,In_1736);
nor U234 (N_234,In_616,In_634);
nor U235 (N_235,In_1897,In_442);
and U236 (N_236,In_706,In_1164);
and U237 (N_237,In_742,In_21);
nand U238 (N_238,In_703,In_1928);
or U239 (N_239,In_1174,In_12);
nand U240 (N_240,In_349,In_862);
or U241 (N_241,In_754,In_1571);
nand U242 (N_242,In_125,In_1554);
nor U243 (N_243,In_1959,In_109);
and U244 (N_244,In_959,In_408);
nor U245 (N_245,In_1832,In_1676);
or U246 (N_246,In_1076,In_944);
or U247 (N_247,In_909,In_851);
or U248 (N_248,In_241,In_678);
nor U249 (N_249,In_1246,In_1983);
nand U250 (N_250,In_1533,In_1335);
and U251 (N_251,In_1024,In_1058);
nor U252 (N_252,In_702,In_362);
nand U253 (N_253,In_542,In_655);
nand U254 (N_254,In_1850,In_1465);
or U255 (N_255,In_821,In_1569);
or U256 (N_256,In_631,In_1938);
and U257 (N_257,In_441,In_1272);
nand U258 (N_258,In_1022,In_1985);
and U259 (N_259,In_1424,In_347);
nor U260 (N_260,In_1726,In_1716);
nand U261 (N_261,In_1824,In_1619);
nor U262 (N_262,In_784,In_1534);
and U263 (N_263,In_97,In_1841);
nand U264 (N_264,In_1159,In_1865);
nand U265 (N_265,In_823,In_276);
and U266 (N_266,In_459,In_1884);
and U267 (N_267,In_1480,In_521);
or U268 (N_268,In_1234,In_1746);
or U269 (N_269,In_1267,In_457);
nor U270 (N_270,In_1450,In_1452);
nor U271 (N_271,In_435,In_745);
and U272 (N_272,In_1595,In_681);
or U273 (N_273,In_603,In_912);
or U274 (N_274,In_325,In_306);
or U275 (N_275,In_930,In_1835);
or U276 (N_276,In_88,In_1068);
or U277 (N_277,In_186,In_1883);
or U278 (N_278,In_1136,In_1493);
nand U279 (N_279,In_224,In_1566);
or U280 (N_280,In_6,In_1964);
nand U281 (N_281,In_1152,In_1404);
nand U282 (N_282,In_181,In_871);
nor U283 (N_283,In_747,In_1876);
nor U284 (N_284,In_1238,In_1908);
nand U285 (N_285,In_330,In_1161);
and U286 (N_286,In_1748,In_950);
nand U287 (N_287,In_1644,In_518);
nor U288 (N_288,In_1879,In_1967);
or U289 (N_289,In_80,In_1242);
nand U290 (N_290,In_1664,In_579);
nand U291 (N_291,In_1613,In_865);
nand U292 (N_292,In_831,In_667);
and U293 (N_293,In_1945,In_22);
xor U294 (N_294,In_1105,In_1671);
and U295 (N_295,In_286,In_1931);
nor U296 (N_296,In_1669,In_1757);
nand U297 (N_297,In_1602,In_1074);
and U298 (N_298,In_225,In_874);
or U299 (N_299,In_1735,In_963);
xnor U300 (N_300,In_1701,In_1788);
nor U301 (N_301,In_1502,In_190);
or U302 (N_302,In_571,In_1433);
and U303 (N_303,In_431,In_1653);
nand U304 (N_304,In_194,In_1146);
xor U305 (N_305,In_219,In_386);
nand U306 (N_306,In_753,In_695);
and U307 (N_307,In_1184,In_410);
nor U308 (N_308,In_1041,In_182);
nand U309 (N_309,In_1363,In_1712);
or U310 (N_310,In_575,In_532);
nor U311 (N_311,In_445,In_309);
or U312 (N_312,In_1148,In_1536);
nand U313 (N_313,In_763,In_304);
or U314 (N_314,In_278,In_451);
nor U315 (N_315,In_759,In_74);
nor U316 (N_316,In_1739,In_908);
or U317 (N_317,In_426,In_1710);
and U318 (N_318,In_58,In_395);
or U319 (N_319,In_589,In_904);
or U320 (N_320,In_490,In_1783);
nand U321 (N_321,In_1860,In_1365);
xnor U322 (N_322,In_1902,In_123);
nor U323 (N_323,In_1582,In_352);
and U324 (N_324,In_1690,In_1719);
nand U325 (N_325,In_1649,In_513);
nand U326 (N_326,In_1115,In_828);
nand U327 (N_327,In_853,In_1523);
or U328 (N_328,In_1706,In_848);
nor U329 (N_329,In_531,In_212);
and U330 (N_330,In_926,In_781);
or U331 (N_331,In_1727,In_1906);
or U332 (N_332,In_659,In_818);
nor U333 (N_333,In_987,In_274);
nand U334 (N_334,In_679,In_265);
nand U335 (N_335,In_121,In_381);
and U336 (N_336,In_137,In_417);
nand U337 (N_337,In_342,In_1044);
nor U338 (N_338,In_449,In_1171);
nand U339 (N_339,In_867,In_592);
nand U340 (N_340,In_1606,In_401);
xnor U341 (N_341,In_356,In_214);
nand U342 (N_342,In_645,In_830);
nor U343 (N_343,In_1003,In_155);
and U344 (N_344,In_1109,In_244);
xor U345 (N_345,In_1353,In_90);
nand U346 (N_346,In_1346,In_785);
nand U347 (N_347,In_1599,In_146);
nand U348 (N_348,In_96,In_105);
nor U349 (N_349,In_1219,In_279);
nand U350 (N_350,In_675,In_1456);
nor U351 (N_351,In_664,In_1097);
nor U352 (N_352,In_584,In_1498);
and U353 (N_353,In_795,In_0);
nor U354 (N_354,In_807,In_1933);
nand U355 (N_355,In_1255,In_483);
or U356 (N_356,In_615,In_370);
or U357 (N_357,In_1260,In_1458);
or U358 (N_358,In_481,In_1123);
nor U359 (N_359,In_134,In_1316);
nand U360 (N_360,In_597,In_1304);
nor U361 (N_361,In_802,In_630);
nor U362 (N_362,In_952,In_869);
and U363 (N_363,In_776,In_1188);
nor U364 (N_364,In_935,In_471);
and U365 (N_365,In_1168,In_1511);
and U366 (N_366,In_1648,In_1913);
nand U367 (N_367,In_1578,In_1855);
and U368 (N_368,In_213,In_680);
xnor U369 (N_369,In_1799,In_530);
and U370 (N_370,In_1356,In_861);
nand U371 (N_371,In_436,In_1486);
and U372 (N_372,In_782,In_1466);
nand U373 (N_373,In_1637,In_1185);
or U374 (N_374,In_1091,In_1552);
nand U375 (N_375,In_81,In_1358);
nor U376 (N_376,In_414,In_1755);
or U377 (N_377,In_850,In_588);
nor U378 (N_378,In_1409,In_622);
or U379 (N_379,In_397,In_1231);
and U380 (N_380,In_147,In_674);
or U381 (N_381,In_1310,In_574);
nor U382 (N_382,In_291,In_647);
or U383 (N_383,In_1968,In_902);
nand U384 (N_384,In_1912,In_582);
or U385 (N_385,In_355,In_51);
nand U386 (N_386,In_686,In_1873);
nand U387 (N_387,In_854,In_1539);
nand U388 (N_388,In_464,In_1973);
and U389 (N_389,In_1035,In_50);
and U390 (N_390,In_705,In_1540);
nor U391 (N_391,In_1020,In_211);
xnor U392 (N_392,In_199,In_360);
or U393 (N_393,In_1916,In_1061);
and U394 (N_394,In_1323,In_485);
xnor U395 (N_395,In_1378,In_296);
nand U396 (N_396,In_1797,In_1862);
or U397 (N_397,In_938,In_1110);
nand U398 (N_398,In_1473,In_1369);
nand U399 (N_399,In_406,In_1447);
nor U400 (N_400,In_783,In_1027);
and U401 (N_401,In_210,In_1047);
or U402 (N_402,In_894,In_1740);
nor U403 (N_403,In_1344,In_167);
and U404 (N_404,In_710,In_1479);
nand U405 (N_405,In_786,In_1332);
nand U406 (N_406,In_824,In_1429);
and U407 (N_407,In_1768,In_53);
nand U408 (N_408,In_1745,In_1975);
xor U409 (N_409,In_433,In_1957);
and U410 (N_410,In_1885,In_338);
nand U411 (N_411,In_1966,In_1001);
or U412 (N_412,In_1763,In_517);
xor U413 (N_413,In_354,In_984);
and U414 (N_414,In_1987,In_247);
nand U415 (N_415,In_1153,In_1512);
or U416 (N_416,In_140,In_1556);
nor U417 (N_417,In_1192,In_497);
and U418 (N_418,In_1400,In_877);
or U419 (N_419,In_1411,In_392);
or U420 (N_420,In_1297,In_1265);
nand U421 (N_421,In_1317,In_196);
nor U422 (N_422,In_41,In_714);
or U423 (N_423,In_1937,In_519);
nand U424 (N_424,In_596,In_600);
or U425 (N_425,In_1584,In_57);
and U426 (N_426,In_1956,In_1218);
or U427 (N_427,In_149,In_1229);
nor U428 (N_428,In_1826,In_71);
nand U429 (N_429,In_129,In_881);
or U430 (N_430,In_1514,In_486);
or U431 (N_431,In_1082,In_788);
xor U432 (N_432,In_1543,In_1662);
nand U433 (N_433,In_720,In_1274);
nor U434 (N_434,In_982,In_896);
xor U435 (N_435,In_1375,In_1986);
nand U436 (N_436,In_1457,In_1842);
nor U437 (N_437,In_238,In_1694);
nor U438 (N_438,In_5,In_729);
or U439 (N_439,In_1172,In_1315);
nor U440 (N_440,In_1808,In_1167);
nor U441 (N_441,In_1376,In_844);
nand U442 (N_442,In_1391,In_640);
and U443 (N_443,In_1470,In_346);
or U444 (N_444,In_1319,In_717);
or U445 (N_445,In_79,In_1073);
nand U446 (N_446,In_396,In_1398);
and U447 (N_447,In_1348,In_1840);
and U448 (N_448,In_351,In_317);
xnor U449 (N_449,In_1308,In_556);
nor U450 (N_450,In_1812,In_1666);
nand U451 (N_451,In_1863,In_1546);
and U452 (N_452,In_405,In_951);
and U453 (N_453,In_1927,In_842);
nand U454 (N_454,In_1261,In_666);
and U455 (N_455,In_882,In_1816);
nand U456 (N_456,In_1550,In_1950);
nand U457 (N_457,In_1620,In_174);
or U458 (N_458,In_668,In_1854);
nor U459 (N_459,In_1318,In_84);
nor U460 (N_460,In_1328,In_1955);
xnor U461 (N_461,In_150,In_606);
nor U462 (N_462,In_825,In_1296);
nor U463 (N_463,In_1772,In_969);
and U464 (N_464,In_361,In_1779);
or U465 (N_465,In_1312,In_448);
and U466 (N_466,In_1327,In_209);
xnor U467 (N_467,In_1909,In_520);
nand U468 (N_468,In_814,In_833);
and U469 (N_469,In_1762,In_1720);
nor U470 (N_470,In_1009,In_1647);
or U471 (N_471,In_1807,In_1761);
nand U472 (N_472,In_657,In_855);
nor U473 (N_473,In_685,In_1886);
or U474 (N_474,In_1686,In_1588);
nor U475 (N_475,In_1610,In_1067);
nor U476 (N_476,In_590,In_1194);
xnor U477 (N_477,In_1438,In_1269);
or U478 (N_478,In_463,In_327);
xor U479 (N_479,In_1107,In_1045);
or U480 (N_480,In_602,In_348);
nor U481 (N_481,In_1160,In_1542);
or U482 (N_482,In_1836,In_83);
nand U483 (N_483,In_568,In_326);
and U484 (N_484,In_281,In_1978);
nand U485 (N_485,In_473,In_1098);
nand U486 (N_486,In_1294,In_1593);
and U487 (N_487,In_1379,In_1211);
nor U488 (N_488,In_400,In_1691);
and U489 (N_489,In_323,In_587);
and U490 (N_490,In_1528,In_14);
nand U491 (N_491,In_777,In_421);
nor U492 (N_492,In_1049,In_768);
and U493 (N_493,In_133,In_1040);
nor U494 (N_494,In_1641,In_313);
or U495 (N_495,In_1085,In_545);
xnor U496 (N_496,In_1626,In_570);
nand U497 (N_497,In_766,In_890);
xor U498 (N_498,In_1481,In_455);
xor U499 (N_499,In_536,In_144);
or U500 (N_500,In_1773,In_1651);
nand U501 (N_501,In_499,In_1861);
nand U502 (N_502,In_1965,In_1338);
xnor U503 (N_503,In_1868,In_1586);
xor U504 (N_504,In_879,In_983);
or U505 (N_505,In_92,In_1389);
and U506 (N_506,In_778,In_168);
nand U507 (N_507,In_990,In_1693);
nor U508 (N_508,In_235,In_799);
nand U509 (N_509,In_1617,In_1640);
and U510 (N_510,In_673,In_797);
xnor U511 (N_511,In_446,In_1095);
nand U512 (N_512,In_508,In_350);
nor U513 (N_513,In_965,In_1926);
nor U514 (N_514,In_609,In_1605);
xnor U515 (N_515,In_173,In_812);
or U516 (N_516,In_1394,In_460);
nor U517 (N_517,In_60,In_1000);
and U518 (N_518,In_1924,In_1598);
nor U519 (N_519,In_253,In_258);
or U520 (N_520,In_1106,In_1659);
nor U521 (N_521,In_1239,In_815);
or U522 (N_522,In_331,In_1891);
nand U523 (N_523,In_502,In_1963);
nor U524 (N_524,In_1565,In_750);
nand U525 (N_525,In_206,In_886);
nand U526 (N_526,In_1233,In_294);
nor U527 (N_527,In_826,In_217);
or U528 (N_528,In_724,In_252);
xor U529 (N_529,In_507,In_1029);
and U530 (N_530,In_1403,In_1896);
and U531 (N_531,In_1422,In_1149);
or U532 (N_532,In_343,In_1917);
and U533 (N_533,In_1871,In_1345);
and U534 (N_534,In_936,In_691);
or U535 (N_535,In_1111,In_15);
xor U536 (N_536,In_1197,In_427);
and U537 (N_537,In_897,In_1991);
and U538 (N_538,In_1195,In_438);
xor U539 (N_539,In_1791,In_1495);
nand U540 (N_540,In_636,In_1054);
nor U541 (N_541,In_543,In_1361);
nor U542 (N_542,In_1081,In_1038);
nor U543 (N_543,In_1302,In_687);
nand U544 (N_544,In_223,In_883);
nand U545 (N_545,In_1970,In_1490);
nand U546 (N_546,In_1526,In_3);
xnor U547 (N_547,In_1695,In_70);
nor U548 (N_548,In_907,In_1721);
xnor U549 (N_549,In_1213,In_1764);
and U550 (N_550,In_1776,In_380);
or U551 (N_551,In_237,In_98);
and U552 (N_552,In_220,In_207);
nand U553 (N_553,In_422,In_1230);
nor U554 (N_554,In_1675,In_1108);
nand U555 (N_555,In_1128,In_450);
nor U556 (N_556,In_496,In_153);
and U557 (N_557,In_78,In_915);
or U558 (N_558,In_528,In_185);
xnor U559 (N_559,In_384,In_1388);
and U560 (N_560,In_232,In_7);
nor U561 (N_561,In_884,In_295);
and U562 (N_562,In_613,In_648);
nand U563 (N_563,In_1775,In_716);
or U564 (N_564,In_954,In_1954);
or U565 (N_565,In_359,In_1157);
xnor U566 (N_566,In_136,In_498);
nor U567 (N_567,In_1333,In_1156);
nand U568 (N_568,In_382,In_1446);
xnor U569 (N_569,In_1689,In_1380);
nor U570 (N_570,In_1687,In_1384);
nor U571 (N_571,In_1307,In_577);
nor U572 (N_572,In_322,In_569);
nor U573 (N_573,In_1374,In_111);
or U574 (N_574,In_1831,In_661);
nand U575 (N_575,In_1551,In_1142);
and U576 (N_576,In_1276,In_192);
or U577 (N_577,In_1786,In_488);
or U578 (N_578,In_267,In_179);
nor U579 (N_579,In_484,In_1150);
nand U580 (N_580,In_755,In_1646);
nor U581 (N_581,In_756,In_1553);
and U582 (N_582,In_1290,In_1661);
nand U583 (N_583,In_437,In_439);
and U584 (N_584,In_524,In_419);
or U585 (N_585,In_1485,In_701);
nor U586 (N_586,In_1780,In_1638);
nor U587 (N_587,In_166,In_434);
nand U588 (N_588,In_1507,In_1352);
nor U589 (N_589,In_719,In_156);
nor U590 (N_590,In_487,In_1930);
or U591 (N_591,In_1043,In_1382);
nor U592 (N_592,In_822,In_289);
nand U593 (N_593,In_1347,In_1907);
nor U594 (N_594,In_792,In_107);
nand U595 (N_595,In_1017,In_550);
and U596 (N_596,In_1849,In_725);
nor U597 (N_597,In_1530,In_672);
nand U598 (N_598,In_102,In_1289);
and U599 (N_599,In_1608,In_1901);
or U600 (N_600,In_72,In_1220);
and U601 (N_601,In_1244,In_1866);
xnor U602 (N_602,In_1387,In_9);
xor U603 (N_603,In_746,In_1453);
nor U604 (N_604,In_1852,In_607);
and U605 (N_605,In_1845,In_1257);
nand U606 (N_606,In_302,In_1086);
nand U607 (N_607,In_389,In_595);
nor U608 (N_608,In_1483,In_283);
or U609 (N_609,In_376,In_1817);
nor U610 (N_610,In_1616,In_1527);
or U611 (N_611,In_1697,In_409);
xnor U612 (N_612,In_1101,In_803);
nor U613 (N_613,In_1016,In_227);
and U614 (N_614,In_248,In_503);
nand U615 (N_615,In_1857,In_1881);
nor U616 (N_616,In_1343,In_476);
and U617 (N_617,In_1193,In_1545);
nand U618 (N_618,In_572,In_889);
or U619 (N_619,In_925,In_945);
and U620 (N_620,In_804,In_1847);
xnor U621 (N_621,In_1633,In_65);
nand U622 (N_622,In_429,In_1182);
nor U623 (N_623,In_1071,In_866);
nor U624 (N_624,In_1732,In_345);
or U625 (N_625,In_171,In_614);
or U626 (N_626,In_734,In_1935);
and U627 (N_627,In_924,In_1715);
and U628 (N_628,In_843,In_608);
nand U629 (N_629,In_1583,In_1870);
nor U630 (N_630,In_1743,In_671);
and U631 (N_631,In_892,In_566);
and U632 (N_632,In_560,In_373);
nor U633 (N_633,In_1976,In_698);
nand U634 (N_634,In_962,In_385);
and U635 (N_635,In_365,In_1173);
or U636 (N_636,In_432,In_1217);
and U637 (N_637,In_1248,In_1227);
nor U638 (N_638,In_1434,In_1519);
nor U639 (N_639,In_876,In_1292);
and U640 (N_640,In_1283,In_75);
nor U641 (N_641,In_23,In_727);
xnor U642 (N_642,In_1216,In_1898);
nand U643 (N_643,In_303,In_501);
or U644 (N_644,In_1713,In_1820);
nand U645 (N_645,In_162,In_1405);
and U646 (N_646,In_1920,In_49);
or U647 (N_647,In_151,In_1187);
and U648 (N_648,In_1851,In_120);
nand U649 (N_649,In_808,In_960);
nor U650 (N_650,In_1683,In_1189);
or U651 (N_651,In_1655,In_629);
or U652 (N_652,In_1782,In_1096);
nand U653 (N_653,In_934,In_1702);
and U654 (N_654,In_163,In_1126);
nor U655 (N_655,In_557,In_1336);
or U656 (N_656,In_1793,In_1023);
and U657 (N_657,In_1476,In_1672);
nand U658 (N_658,In_403,In_1630);
nor U659 (N_659,In_1397,In_806);
nor U660 (N_660,In_1703,In_601);
or U661 (N_661,In_477,In_1789);
and U662 (N_662,In_1665,In_37);
or U663 (N_663,In_1445,In_259);
nor U664 (N_664,In_1734,In_1467);
and U665 (N_665,In_1028,In_994);
nand U666 (N_666,In_548,In_1760);
and U667 (N_667,In_1856,In_494);
or U668 (N_668,In_1811,In_820);
xor U669 (N_669,In_635,In_525);
and U670 (N_670,In_1910,In_1947);
nand U671 (N_671,In_1724,In_878);
and U672 (N_672,In_46,In_329);
nand U673 (N_673,In_956,In_1915);
and U674 (N_674,In_379,In_578);
or U675 (N_675,In_1385,In_55);
nand U676 (N_676,In_619,In_277);
nand U677 (N_677,In_1141,In_19);
nand U678 (N_678,In_1254,In_1175);
nor U679 (N_679,In_654,In_479);
nand U680 (N_680,In_1923,In_775);
and U681 (N_681,In_1771,In_903);
xor U682 (N_682,In_1821,In_858);
nand U683 (N_683,In_424,In_1056);
nand U684 (N_684,In_114,In_64);
nand U685 (N_685,In_193,In_299);
nor U686 (N_686,In_1560,In_1125);
or U687 (N_687,In_670,In_665);
nand U688 (N_688,In_411,In_1948);
nor U689 (N_689,In_73,In_1518);
xnor U690 (N_690,In_1366,In_1678);
nand U691 (N_691,In_1859,In_318);
and U692 (N_692,In_1423,In_662);
and U693 (N_693,In_1858,In_658);
nand U694 (N_694,In_1785,In_470);
nand U695 (N_695,In_721,In_1839);
xnor U696 (N_696,In_864,In_103);
and U697 (N_697,In_728,In_996);
or U698 (N_698,In_1475,In_262);
nand U699 (N_699,In_1428,In_1888);
or U700 (N_700,In_1612,In_835);
and U701 (N_701,In_1741,In_1139);
xor U702 (N_702,In_68,In_1766);
and U703 (N_703,In_1253,In_39);
nor U704 (N_704,In_54,In_937);
nor U705 (N_705,In_89,In_444);
nand U706 (N_706,In_48,In_1183);
xor U707 (N_707,In_1680,In_1237);
xor U708 (N_708,In_978,In_69);
xnor U709 (N_709,In_1604,In_468);
nand U710 (N_710,In_1117,In_722);
and U711 (N_711,In_180,In_383);
nand U712 (N_712,In_169,In_1305);
nor U713 (N_713,In_176,In_1131);
nand U714 (N_714,In_154,In_1731);
or U715 (N_715,In_1145,In_398);
nor U716 (N_716,In_1652,In_642);
nand U717 (N_717,In_254,In_652);
or U718 (N_718,In_989,In_913);
nor U719 (N_719,In_1221,In_387);
and U720 (N_720,In_34,In_264);
nand U721 (N_721,In_931,In_692);
nand U722 (N_722,In_1390,In_723);
and U723 (N_723,In_1442,In_239);
and U724 (N_724,In_1144,In_1266);
nand U725 (N_725,In_130,In_1251);
and U726 (N_726,In_31,In_255);
or U727 (N_727,In_1941,In_863);
nor U728 (N_728,In_1837,In_1742);
and U729 (N_729,In_1062,In_1679);
nand U730 (N_730,In_1729,In_1436);
or U731 (N_731,In_1549,In_1225);
nand U732 (N_732,In_462,In_1969);
nor U733 (N_733,In_1355,In_320);
nand U734 (N_734,In_1472,In_626);
nor U735 (N_735,In_122,In_1496);
nand U736 (N_736,In_1787,In_273);
and U737 (N_737,In_440,In_269);
or U738 (N_738,In_1622,In_1151);
and U739 (N_739,In_364,In_975);
or U740 (N_740,In_1226,In_1454);
nand U741 (N_741,In_1494,In_739);
xnor U742 (N_742,In_540,In_452);
and U743 (N_743,In_1460,In_772);
and U744 (N_744,In_2,In_1572);
and U745 (N_745,In_1796,In_527);
nor U746 (N_746,In_87,In_946);
and U747 (N_747,In_1198,In_420);
or U748 (N_748,In_594,In_1547);
nor U749 (N_749,In_511,In_538);
xnor U750 (N_750,In_988,In_813);
nand U751 (N_751,In_581,In_1462);
nor U752 (N_752,In_559,In_27);
xor U753 (N_753,In_771,In_964);
nand U754 (N_754,In_1878,In_1996);
and U755 (N_755,In_1432,In_1033);
or U756 (N_756,In_1055,In_282);
nor U757 (N_757,In_949,In_1631);
xor U758 (N_758,In_800,In_1997);
and U759 (N_759,In_1129,In_1827);
nor U760 (N_760,In_198,In_628);
nand U761 (N_761,In_1298,In_1714);
and U762 (N_762,In_101,In_919);
xor U763 (N_763,In_1510,In_1618);
or U764 (N_764,In_461,In_1992);
xor U765 (N_765,In_1008,In_1203);
nand U766 (N_766,In_1562,In_335);
nor U767 (N_767,In_534,In_1170);
and U768 (N_768,In_1867,In_305);
nand U769 (N_769,In_1401,In_715);
nor U770 (N_770,In_1499,In_732);
and U771 (N_771,In_774,In_1243);
nor U772 (N_772,In_1668,In_1354);
nor U773 (N_773,In_261,In_1629);
or U774 (N_774,In_197,In_1191);
nor U775 (N_775,In_885,In_1822);
xor U776 (N_776,In_576,In_1249);
nor U777 (N_777,In_1478,In_489);
nor U778 (N_778,In_1090,In_1186);
nor U779 (N_779,In_573,In_1810);
xor U780 (N_780,In_1087,In_85);
nand U781 (N_781,In_870,In_973);
nor U782 (N_782,In_1030,In_1971);
nor U783 (N_783,In_1291,In_275);
and U784 (N_784,In_563,In_1373);
or U785 (N_785,In_1468,In_1042);
and U786 (N_786,In_604,In_1819);
or U787 (N_787,In_1537,In_743);
nor U788 (N_788,In_967,In_42);
or U789 (N_789,In_1416,In_1282);
and U790 (N_790,In_1247,In_1492);
nand U791 (N_791,In_736,In_1176);
or U792 (N_792,In_469,In_735);
xor U793 (N_793,In_1597,In_816);
or U794 (N_794,In_1951,In_1487);
or U795 (N_795,In_1223,In_202);
and U796 (N_796,In_922,In_1753);
nor U797 (N_797,In_857,In_143);
nand U798 (N_798,In_1449,In_598);
nand U799 (N_799,In_514,In_1386);
xnor U800 (N_800,In_1650,In_1750);
nand U801 (N_801,In_509,In_1214);
nand U802 (N_802,In_1368,In_118);
and U803 (N_803,In_929,In_8);
xnor U804 (N_804,In_605,In_1934);
nor U805 (N_805,In_1078,In_288);
xor U806 (N_806,In_927,In_591);
xor U807 (N_807,In_888,In_1515);
nand U808 (N_808,In_762,In_1381);
or U809 (N_809,In_942,In_709);
and U810 (N_810,In_1905,In_1364);
or U811 (N_811,In_751,In_1089);
nand U812 (N_812,In_178,In_242);
nand U813 (N_813,In_1155,In_738);
nand U814 (N_814,In_730,In_981);
nand U815 (N_815,In_1180,In_1395);
nor U816 (N_816,In_1127,In_1744);
and U817 (N_817,In_811,In_339);
nand U818 (N_818,In_953,In_17);
or U819 (N_819,In_718,In_1440);
nand U820 (N_820,In_632,In_266);
and U821 (N_821,In_1419,In_1169);
or U822 (N_822,In_94,In_1600);
nor U823 (N_823,In_1134,In_749);
nand U824 (N_824,In_1594,In_846);
or U825 (N_825,In_1051,In_752);
nand U826 (N_826,In_1426,In_1521);
and U827 (N_827,In_1007,In_425);
and U828 (N_828,In_999,In_1628);
nor U829 (N_829,In_555,In_627);
nor U830 (N_830,In_744,In_1564);
nand U831 (N_831,In_1418,In_447);
and U832 (N_832,In_1138,In_1383);
nand U833 (N_833,In_1828,In_11);
nand U834 (N_834,In_875,In_1448);
or U835 (N_835,In_921,In_1635);
nand U836 (N_836,In_1607,In_1580);
or U837 (N_837,In_847,In_740);
or U838 (N_838,In_1984,In_1342);
and U839 (N_839,In_1830,In_240);
nand U840 (N_840,In_1050,In_558);
and U841 (N_841,In_1258,In_1623);
xor U842 (N_842,In_47,In_1321);
nor U843 (N_843,In_1410,In_1777);
nor U844 (N_844,In_1730,In_159);
or U845 (N_845,In_26,In_222);
nor U846 (N_846,In_1491,In_337);
or U847 (N_847,In_187,In_1718);
and U848 (N_848,In_974,In_1524);
or U849 (N_849,In_1349,In_1939);
and U850 (N_850,In_966,In_1711);
nor U851 (N_851,In_985,In_1337);
xnor U852 (N_852,In_567,In_995);
nor U853 (N_853,In_1277,In_1212);
nor U854 (N_854,In_1179,In_801);
or U855 (N_855,In_1504,In_547);
and U856 (N_856,In_693,In_551);
xor U857 (N_857,In_1196,In_829);
and U858 (N_858,In_378,In_1946);
or U859 (N_859,In_1147,In_1392);
or U860 (N_860,In_1326,In_618);
and U861 (N_861,In_505,In_1372);
xor U862 (N_862,In_1114,In_86);
nor U863 (N_863,In_1809,In_713);
nor U864 (N_864,In_300,In_1627);
or U865 (N_865,In_968,In_307);
and U866 (N_866,In_372,In_1587);
nand U867 (N_867,In_1459,In_1032);
nand U868 (N_868,In_1093,In_1359);
and U869 (N_869,In_453,In_552);
nor U870 (N_870,In_1642,In_368);
or U871 (N_871,In_1778,In_1199);
and U872 (N_872,In_1688,In_1592);
nand U873 (N_873,In_157,In_901);
nor U874 (N_874,In_1685,In_268);
and U875 (N_875,In_1012,In_1872);
nor U876 (N_876,In_1075,In_1953);
and U877 (N_877,In_948,In_18);
nand U878 (N_878,In_1295,In_415);
and U879 (N_879,In_132,In_997);
or U880 (N_880,In_256,In_506);
or U881 (N_881,In_1299,In_1733);
xnor U882 (N_882,In_562,In_637);
xor U883 (N_883,In_787,In_832);
and U884 (N_884,In_1993,In_1133);
and U885 (N_885,In_493,In_911);
nand U886 (N_886,In_683,In_1555);
nor U887 (N_887,In_1960,In_510);
xnor U888 (N_888,In_1080,In_1843);
nor U889 (N_889,In_1658,In_1614);
nand U890 (N_890,In_215,In_1517);
and U891 (N_891,In_1601,In_13);
nor U892 (N_892,In_767,In_840);
nor U893 (N_893,In_1529,In_1102);
and U894 (N_894,In_236,In_1350);
and U895 (N_895,In_905,In_1263);
and U896 (N_896,In_1036,In_644);
or U897 (N_897,In_1516,In_1303);
xnor U898 (N_898,In_1503,In_1288);
and U899 (N_899,In_852,In_623);
nor U900 (N_900,In_56,In_656);
nand U901 (N_901,In_663,In_646);
or U902 (N_902,In_712,In_1723);
and U903 (N_903,In_117,In_1575);
nand U904 (N_904,In_43,In_1015);
nor U905 (N_905,In_1925,In_1330);
or U906 (N_906,In_638,In_758);
and U907 (N_907,In_106,In_512);
or U908 (N_908,In_404,In_780);
and U909 (N_909,In_1018,In_1535);
xor U910 (N_910,In_1441,In_1573);
or U911 (N_911,In_1451,In_1814);
nand U912 (N_912,In_1804,In_1399);
or U913 (N_913,In_564,In_1413);
nor U914 (N_914,In_1674,In_324);
nand U915 (N_915,In_593,In_374);
nand U916 (N_916,In_216,In_677);
and U917 (N_917,In_526,In_363);
nor U918 (N_918,In_1241,In_696);
nor U919 (N_919,In_910,In_1010);
or U920 (N_920,In_177,In_1567);
nand U921 (N_921,In_1325,In_1589);
or U922 (N_922,In_1339,In_1280);
nor U923 (N_923,In_1611,In_914);
nand U924 (N_924,In_172,In_1181);
nor U925 (N_925,In_1166,In_1944);
nor U926 (N_926,In_200,In_1351);
and U927 (N_927,In_298,In_1066);
nor U928 (N_928,In_1784,In_1031);
or U929 (N_929,In_1581,In_1143);
or U930 (N_930,In_1805,In_917);
xnor U931 (N_931,In_880,In_1311);
nor U932 (N_932,In_1362,In_1882);
nand U933 (N_933,In_773,In_1256);
nor U934 (N_934,In_465,In_183);
xor U935 (N_935,In_537,In_110);
or U936 (N_936,In_131,In_1982);
and U937 (N_937,In_529,In_1443);
nor U938 (N_938,In_583,In_699);
nor U939 (N_939,In_1900,In_32);
xnor U940 (N_940,In_1039,In_474);
nor U941 (N_941,In_315,In_972);
xor U942 (N_942,In_856,In_1004);
nor U943 (N_943,In_1563,In_761);
nand U944 (N_944,In_1660,In_872);
nor U945 (N_945,In_1334,In_1293);
or U946 (N_946,In_467,In_599);
nor U947 (N_947,In_135,In_164);
xor U948 (N_948,In_1815,In_1692);
xor U949 (N_949,In_1500,In_201);
nor U950 (N_950,In_1259,In_688);
or U951 (N_951,In_796,In_1497);
nor U952 (N_952,In_1064,In_991);
nor U953 (N_953,In_1559,In_1112);
nand U954 (N_954,In_62,In_1747);
nor U955 (N_955,In_1806,In_1072);
nand U956 (N_956,In_986,In_1222);
nor U957 (N_957,In_1414,In_377);
and U958 (N_958,In_794,In_358);
nor U959 (N_959,In_226,In_977);
nand U960 (N_960,In_458,In_1803);
nand U961 (N_961,In_1505,In_809);
nand U962 (N_962,In_1754,In_205);
nand U963 (N_963,In_554,In_1210);
nor U964 (N_964,In_1118,In_1140);
nor U965 (N_965,In_1393,In_682);
and U966 (N_966,In_1461,In_1488);
and U967 (N_967,In_918,In_257);
and U968 (N_968,In_1178,In_1048);
and U969 (N_969,In_1415,In_516);
and U970 (N_970,In_1704,In_228);
nand U971 (N_971,In_900,In_1749);
nor U972 (N_972,In_523,In_1892);
xnor U973 (N_973,In_1019,In_624);
xor U974 (N_974,In_1568,In_1717);
nor U975 (N_975,In_1962,In_495);
and U976 (N_976,In_263,In_764);
or U977 (N_977,In_1558,In_1430);
nor U978 (N_978,In_1929,In_1904);
nand U979 (N_979,In_923,In_1979);
nor U980 (N_980,In_1994,In_321);
nor U981 (N_981,In_375,In_67);
nor U982 (N_982,In_1737,In_1070);
or U983 (N_983,In_340,In_1579);
nor U984 (N_984,In_184,In_1412);
and U985 (N_985,In_287,In_99);
nand U986 (N_986,In_1877,In_1818);
nand U987 (N_987,In_412,In_1942);
nand U988 (N_988,In_789,In_189);
nand U989 (N_989,In_1271,In_312);
xnor U990 (N_990,In_1921,In_1006);
nor U991 (N_991,In_1130,In_1531);
xor U992 (N_992,In_1202,In_290);
nor U993 (N_993,In_939,In_689);
or U994 (N_994,In_1208,In_1513);
or U995 (N_995,In_1094,In_301);
or U996 (N_996,In_726,In_1591);
nand U997 (N_997,In_998,In_549);
or U998 (N_998,In_1974,In_1484);
nor U999 (N_999,In_1728,In_565);
nand U1000 (N_1000,N_842,N_598);
nor U1001 (N_1001,N_498,N_399);
or U1002 (N_1002,N_936,N_309);
xor U1003 (N_1003,N_561,N_84);
nor U1004 (N_1004,N_221,N_768);
or U1005 (N_1005,N_571,N_761);
nor U1006 (N_1006,N_892,N_750);
nand U1007 (N_1007,N_942,N_655);
nor U1008 (N_1008,N_943,N_459);
or U1009 (N_1009,N_981,N_957);
and U1010 (N_1010,N_658,N_595);
or U1011 (N_1011,N_521,N_965);
and U1012 (N_1012,N_850,N_127);
and U1013 (N_1013,N_139,N_111);
and U1014 (N_1014,N_582,N_752);
xnor U1015 (N_1015,N_114,N_134);
nor U1016 (N_1016,N_803,N_470);
and U1017 (N_1017,N_997,N_531);
or U1018 (N_1018,N_427,N_570);
nand U1019 (N_1019,N_450,N_695);
and U1020 (N_1020,N_988,N_108);
and U1021 (N_1021,N_339,N_419);
and U1022 (N_1022,N_808,N_387);
nand U1023 (N_1023,N_220,N_101);
nor U1024 (N_1024,N_744,N_184);
or U1025 (N_1025,N_441,N_182);
nor U1026 (N_1026,N_370,N_204);
nand U1027 (N_1027,N_237,N_157);
nand U1028 (N_1028,N_219,N_929);
or U1029 (N_1029,N_44,N_356);
or U1030 (N_1030,N_466,N_240);
nor U1031 (N_1031,N_626,N_416);
nand U1032 (N_1032,N_281,N_169);
nand U1033 (N_1033,N_980,N_522);
and U1034 (N_1034,N_104,N_707);
or U1035 (N_1035,N_479,N_94);
or U1036 (N_1036,N_946,N_654);
xor U1037 (N_1037,N_923,N_241);
or U1038 (N_1038,N_393,N_349);
nor U1039 (N_1039,N_178,N_420);
and U1040 (N_1040,N_123,N_162);
and U1041 (N_1041,N_351,N_916);
nor U1042 (N_1042,N_870,N_699);
and U1043 (N_1043,N_268,N_95);
and U1044 (N_1044,N_966,N_766);
nand U1045 (N_1045,N_39,N_407);
xor U1046 (N_1046,N_506,N_222);
nor U1047 (N_1047,N_200,N_830);
or U1048 (N_1048,N_238,N_501);
and U1049 (N_1049,N_481,N_728);
nand U1050 (N_1050,N_684,N_312);
and U1051 (N_1051,N_274,N_110);
xor U1052 (N_1052,N_945,N_906);
and U1053 (N_1053,N_218,N_831);
nand U1054 (N_1054,N_235,N_900);
or U1055 (N_1055,N_853,N_671);
nand U1056 (N_1056,N_395,N_856);
and U1057 (N_1057,N_857,N_810);
nand U1058 (N_1058,N_775,N_21);
and U1059 (N_1059,N_961,N_740);
nand U1060 (N_1060,N_635,N_207);
and U1061 (N_1061,N_871,N_10);
nor U1062 (N_1062,N_786,N_852);
nand U1063 (N_1063,N_913,N_990);
or U1064 (N_1064,N_128,N_27);
and U1065 (N_1065,N_85,N_7);
nand U1066 (N_1066,N_310,N_422);
nand U1067 (N_1067,N_998,N_230);
and U1068 (N_1068,N_777,N_637);
or U1069 (N_1069,N_860,N_720);
or U1070 (N_1070,N_26,N_565);
or U1071 (N_1071,N_130,N_978);
or U1072 (N_1072,N_181,N_597);
nor U1073 (N_1073,N_46,N_624);
or U1074 (N_1074,N_279,N_782);
and U1075 (N_1075,N_403,N_993);
xor U1076 (N_1076,N_697,N_974);
and U1077 (N_1077,N_953,N_524);
nand U1078 (N_1078,N_18,N_549);
and U1079 (N_1079,N_541,N_250);
nand U1080 (N_1080,N_909,N_784);
or U1081 (N_1081,N_553,N_348);
nor U1082 (N_1082,N_424,N_193);
nor U1083 (N_1083,N_618,N_4);
xnor U1084 (N_1084,N_319,N_359);
nand U1085 (N_1085,N_61,N_662);
nand U1086 (N_1086,N_35,N_791);
and U1087 (N_1087,N_849,N_176);
nor U1088 (N_1088,N_2,N_669);
or U1089 (N_1089,N_337,N_639);
nor U1090 (N_1090,N_989,N_733);
or U1091 (N_1091,N_800,N_578);
and U1092 (N_1092,N_537,N_632);
xor U1093 (N_1093,N_180,N_622);
nand U1094 (N_1094,N_834,N_560);
or U1095 (N_1095,N_600,N_71);
xor U1096 (N_1096,N_273,N_764);
and U1097 (N_1097,N_429,N_136);
nand U1098 (N_1098,N_225,N_443);
nor U1099 (N_1099,N_66,N_673);
nor U1100 (N_1100,N_794,N_760);
nand U1101 (N_1101,N_342,N_303);
or U1102 (N_1102,N_28,N_523);
nor U1103 (N_1103,N_43,N_864);
xor U1104 (N_1104,N_891,N_45);
and U1105 (N_1105,N_380,N_776);
or U1106 (N_1106,N_848,N_383);
or U1107 (N_1107,N_558,N_79);
or U1108 (N_1108,N_924,N_855);
or U1109 (N_1109,N_890,N_772);
or U1110 (N_1110,N_836,N_217);
and U1111 (N_1111,N_539,N_267);
and U1112 (N_1112,N_709,N_664);
nor U1113 (N_1113,N_227,N_869);
and U1114 (N_1114,N_233,N_31);
xnor U1115 (N_1115,N_64,N_68);
xnor U1116 (N_1116,N_0,N_982);
nand U1117 (N_1117,N_996,N_838);
or U1118 (N_1118,N_436,N_615);
and U1119 (N_1119,N_647,N_748);
xor U1120 (N_1120,N_390,N_398);
nor U1121 (N_1121,N_584,N_379);
and U1122 (N_1122,N_247,N_674);
or U1123 (N_1123,N_140,N_455);
and U1124 (N_1124,N_119,N_333);
nand U1125 (N_1125,N_724,N_629);
nor U1126 (N_1126,N_745,N_801);
nor U1127 (N_1127,N_513,N_69);
nor U1128 (N_1128,N_463,N_311);
nand U1129 (N_1129,N_691,N_528);
nand U1130 (N_1130,N_76,N_505);
or U1131 (N_1131,N_234,N_163);
nand U1132 (N_1132,N_425,N_291);
nor U1133 (N_1133,N_354,N_323);
xnor U1134 (N_1134,N_797,N_362);
or U1135 (N_1135,N_253,N_670);
nand U1136 (N_1136,N_195,N_880);
or U1137 (N_1137,N_576,N_353);
or U1138 (N_1138,N_484,N_895);
nor U1139 (N_1139,N_133,N_885);
and U1140 (N_1140,N_821,N_569);
and U1141 (N_1141,N_36,N_708);
or U1142 (N_1142,N_283,N_471);
or U1143 (N_1143,N_503,N_756);
or U1144 (N_1144,N_210,N_401);
or U1145 (N_1145,N_574,N_117);
or U1146 (N_1146,N_488,N_566);
nor U1147 (N_1147,N_179,N_91);
nor U1148 (N_1148,N_879,N_377);
nor U1149 (N_1149,N_154,N_34);
xor U1150 (N_1150,N_121,N_249);
nand U1151 (N_1151,N_366,N_438);
nand U1152 (N_1152,N_944,N_986);
nand U1153 (N_1153,N_738,N_712);
and U1154 (N_1154,N_586,N_82);
nand U1155 (N_1155,N_889,N_171);
nor U1156 (N_1156,N_282,N_256);
nand U1157 (N_1157,N_208,N_552);
nor U1158 (N_1158,N_486,N_858);
and U1159 (N_1159,N_700,N_115);
or U1160 (N_1160,N_440,N_819);
nand U1161 (N_1161,N_361,N_826);
nor U1162 (N_1162,N_107,N_129);
nor U1163 (N_1163,N_882,N_587);
and U1164 (N_1164,N_694,N_947);
and U1165 (N_1165,N_305,N_198);
or U1166 (N_1166,N_960,N_321);
or U1167 (N_1167,N_734,N_640);
nand U1168 (N_1168,N_285,N_196);
and U1169 (N_1169,N_649,N_809);
nand U1170 (N_1170,N_703,N_839);
nand U1171 (N_1171,N_109,N_706);
nand U1172 (N_1172,N_434,N_844);
nor U1173 (N_1173,N_596,N_341);
nand U1174 (N_1174,N_275,N_87);
or U1175 (N_1175,N_994,N_442);
nand U1176 (N_1176,N_952,N_770);
nand U1177 (N_1177,N_259,N_641);
or U1178 (N_1178,N_755,N_32);
nor U1179 (N_1179,N_502,N_446);
nor U1180 (N_1180,N_785,N_741);
and U1181 (N_1181,N_350,N_33);
nor U1182 (N_1182,N_465,N_435);
nor U1183 (N_1183,N_473,N_261);
or U1184 (N_1184,N_874,N_244);
nand U1185 (N_1185,N_286,N_53);
nor U1186 (N_1186,N_421,N_384);
nand U1187 (N_1187,N_665,N_388);
and U1188 (N_1188,N_332,N_818);
nand U1189 (N_1189,N_754,N_508);
and U1190 (N_1190,N_767,N_74);
nand U1191 (N_1191,N_517,N_676);
and U1192 (N_1192,N_611,N_185);
nand U1193 (N_1193,N_914,N_326);
nand U1194 (N_1194,N_845,N_369);
or U1195 (N_1195,N_49,N_40);
nor U1196 (N_1196,N_645,N_168);
and U1197 (N_1197,N_543,N_668);
nor U1198 (N_1198,N_749,N_663);
nand U1199 (N_1199,N_992,N_716);
or U1200 (N_1200,N_60,N_616);
xor U1201 (N_1201,N_589,N_677);
nor U1202 (N_1202,N_209,N_704);
or U1203 (N_1203,N_710,N_191);
nand U1204 (N_1204,N_451,N_229);
or U1205 (N_1205,N_432,N_80);
nand U1206 (N_1206,N_563,N_73);
and U1207 (N_1207,N_302,N_170);
nor U1208 (N_1208,N_940,N_941);
xor U1209 (N_1209,N_20,N_93);
and U1210 (N_1210,N_392,N_58);
nor U1211 (N_1211,N_16,N_12);
and U1212 (N_1212,N_964,N_788);
nand U1213 (N_1213,N_346,N_55);
or U1214 (N_1214,N_202,N_410);
nor U1215 (N_1215,N_813,N_462);
nand U1216 (N_1216,N_160,N_272);
nand U1217 (N_1217,N_447,N_445);
and U1218 (N_1218,N_771,N_973);
nor U1219 (N_1219,N_365,N_469);
nand U1220 (N_1220,N_89,N_555);
or U1221 (N_1221,N_683,N_491);
nand U1222 (N_1222,N_780,N_526);
and U1223 (N_1223,N_335,N_5);
nor U1224 (N_1224,N_304,N_186);
or U1225 (N_1225,N_148,N_367);
xor U1226 (N_1226,N_899,N_496);
nor U1227 (N_1227,N_859,N_623);
nand U1228 (N_1228,N_423,N_824);
or U1229 (N_1229,N_925,N_426);
nor U1230 (N_1230,N_29,N_461);
or U1231 (N_1231,N_9,N_317);
or U1232 (N_1232,N_939,N_666);
nor U1233 (N_1233,N_861,N_314);
xor U1234 (N_1234,N_783,N_591);
and U1235 (N_1235,N_894,N_535);
xor U1236 (N_1236,N_146,N_48);
nand U1237 (N_1237,N_15,N_13);
or U1238 (N_1238,N_886,N_854);
nor U1239 (N_1239,N_643,N_276);
nand U1240 (N_1240,N_843,N_612);
xor U1241 (N_1241,N_188,N_150);
and U1242 (N_1242,N_347,N_391);
nand U1243 (N_1243,N_721,N_500);
and U1244 (N_1244,N_903,N_456);
nor U1245 (N_1245,N_251,N_642);
and U1246 (N_1246,N_70,N_969);
and U1247 (N_1247,N_37,N_125);
or U1248 (N_1248,N_628,N_255);
and U1249 (N_1249,N_904,N_689);
nor U1250 (N_1250,N_922,N_102);
or U1251 (N_1251,N_65,N_343);
or U1252 (N_1252,N_897,N_141);
nand U1253 (N_1253,N_245,N_585);
nand U1254 (N_1254,N_564,N_829);
nand U1255 (N_1255,N_759,N_120);
or U1256 (N_1256,N_675,N_98);
or U1257 (N_1257,N_472,N_696);
nand U1258 (N_1258,N_527,N_294);
xor U1259 (N_1259,N_30,N_702);
nor U1260 (N_1260,N_873,N_201);
nand U1261 (N_1261,N_557,N_203);
or U1262 (N_1262,N_402,N_765);
or U1263 (N_1263,N_577,N_725);
or U1264 (N_1264,N_968,N_475);
nor U1265 (N_1265,N_409,N_580);
nand U1266 (N_1266,N_715,N_345);
and U1267 (N_1267,N_287,N_536);
xnor U1268 (N_1268,N_933,N_542);
and U1269 (N_1269,N_404,N_787);
xnor U1270 (N_1270,N_138,N_548);
or U1271 (N_1271,N_340,N_389);
nand U1272 (N_1272,N_495,N_534);
or U1273 (N_1273,N_510,N_687);
nor U1274 (N_1274,N_105,N_567);
or U1275 (N_1275,N_173,N_713);
nand U1276 (N_1276,N_652,N_727);
and U1277 (N_1277,N_667,N_551);
or U1278 (N_1278,N_215,N_520);
nand U1279 (N_1279,N_360,N_497);
nor U1280 (N_1280,N_88,N_877);
xor U1281 (N_1281,N_701,N_908);
nor U1282 (N_1282,N_375,N_547);
and U1283 (N_1283,N_962,N_56);
nand U1284 (N_1284,N_747,N_751);
nand U1285 (N_1285,N_688,N_866);
or U1286 (N_1286,N_711,N_289);
and U1287 (N_1287,N_896,N_405);
and U1288 (N_1288,N_984,N_621);
xor U1289 (N_1289,N_805,N_83);
or U1290 (N_1290,N_75,N_828);
xor U1291 (N_1291,N_544,N_183);
nand U1292 (N_1292,N_292,N_653);
and U1293 (N_1293,N_126,N_987);
or U1294 (N_1294,N_802,N_814);
nand U1295 (N_1295,N_735,N_514);
nand U1296 (N_1296,N_532,N_812);
and U1297 (N_1297,N_164,N_116);
and U1298 (N_1298,N_930,N_609);
nand U1299 (N_1299,N_512,N_189);
and U1300 (N_1300,N_919,N_530);
and U1301 (N_1301,N_297,N_951);
nor U1302 (N_1302,N_722,N_729);
or U1303 (N_1303,N_257,N_166);
nor U1304 (N_1304,N_817,N_149);
or U1305 (N_1305,N_627,N_62);
or U1306 (N_1306,N_328,N_482);
and U1307 (N_1307,N_122,N_153);
nor U1308 (N_1308,N_263,N_301);
nand U1309 (N_1309,N_991,N_418);
and U1310 (N_1310,N_242,N_827);
or U1311 (N_1311,N_373,N_862);
nor U1312 (N_1312,N_971,N_67);
or U1313 (N_1313,N_660,N_630);
xor U1314 (N_1314,N_672,N_307);
nand U1315 (N_1315,N_846,N_790);
or U1316 (N_1316,N_572,N_413);
or U1317 (N_1317,N_757,N_415);
nand U1318 (N_1318,N_868,N_685);
nand U1319 (N_1319,N_232,N_816);
and U1320 (N_1320,N_357,N_468);
nor U1321 (N_1321,N_118,N_588);
or U1322 (N_1322,N_206,N_478);
and U1323 (N_1323,N_318,N_264);
nand U1324 (N_1324,N_476,N_698);
nor U1325 (N_1325,N_374,N_975);
and U1326 (N_1326,N_773,N_902);
or U1327 (N_1327,N_950,N_231);
or U1328 (N_1328,N_932,N_499);
and U1329 (N_1329,N_604,N_739);
and U1330 (N_1330,N_51,N_847);
nor U1331 (N_1331,N_278,N_519);
and U1332 (N_1332,N_270,N_22);
nor U1333 (N_1333,N_147,N_863);
nor U1334 (N_1334,N_99,N_876);
nor U1335 (N_1335,N_533,N_631);
nor U1336 (N_1336,N_921,N_57);
and U1337 (N_1337,N_265,N_559);
and U1338 (N_1338,N_17,N_156);
and U1339 (N_1339,N_280,N_90);
nand U1340 (N_1340,N_714,N_78);
and U1341 (N_1341,N_865,N_602);
and U1342 (N_1342,N_358,N_888);
nor U1343 (N_1343,N_97,N_884);
nor U1344 (N_1344,N_492,N_400);
nand U1345 (N_1345,N_983,N_197);
or U1346 (N_1346,N_690,N_959);
nand U1347 (N_1347,N_485,N_833);
or U1348 (N_1348,N_334,N_737);
nand U1349 (N_1349,N_19,N_100);
or U1350 (N_1350,N_594,N_406);
nand U1351 (N_1351,N_659,N_228);
nand U1352 (N_1352,N_718,N_324);
nor U1353 (N_1353,N_758,N_474);
nand U1354 (N_1354,N_288,N_54);
nor U1355 (N_1355,N_252,N_158);
or U1356 (N_1356,N_550,N_601);
nor U1357 (N_1357,N_832,N_917);
nand U1358 (N_1358,N_507,N_736);
or U1359 (N_1359,N_656,N_454);
and U1360 (N_1360,N_433,N_518);
or U1361 (N_1361,N_792,N_545);
or U1362 (N_1362,N_368,N_226);
nor U1363 (N_1363,N_554,N_236);
and U1364 (N_1364,N_408,N_382);
or U1365 (N_1365,N_41,N_778);
or U1366 (N_1366,N_42,N_575);
and U1367 (N_1367,N_266,N_789);
nor U1368 (N_1368,N_428,N_515);
nand U1369 (N_1369,N_967,N_841);
nor U1370 (N_1370,N_956,N_633);
xor U1371 (N_1371,N_298,N_344);
or U1372 (N_1372,N_732,N_137);
nor U1373 (N_1373,N_719,N_460);
nand U1374 (N_1374,N_14,N_371);
or U1375 (N_1375,N_92,N_692);
or U1376 (N_1376,N_636,N_277);
or U1377 (N_1377,N_135,N_928);
and U1378 (N_1378,N_490,N_320);
nor U1379 (N_1379,N_386,N_439);
or U1380 (N_1380,N_705,N_124);
nor U1381 (N_1381,N_151,N_905);
nand U1382 (N_1382,N_680,N_417);
or U1383 (N_1383,N_806,N_187);
nand U1384 (N_1384,N_644,N_835);
or U1385 (N_1385,N_431,N_605);
and U1386 (N_1386,N_603,N_540);
and U1387 (N_1387,N_72,N_437);
nor U1388 (N_1388,N_926,N_887);
or U1389 (N_1389,N_972,N_867);
nand U1390 (N_1390,N_258,N_931);
and U1391 (N_1391,N_910,N_161);
nor U1392 (N_1392,N_59,N_175);
nor U1393 (N_1393,N_325,N_650);
and U1394 (N_1394,N_23,N_920);
and U1395 (N_1395,N_38,N_316);
and U1396 (N_1396,N_493,N_330);
nand U1397 (N_1397,N_338,N_397);
nand U1398 (N_1398,N_753,N_412);
or U1399 (N_1399,N_875,N_47);
and U1400 (N_1400,N_103,N_948);
and U1401 (N_1401,N_284,N_504);
nand U1402 (N_1402,N_331,N_50);
xnor U1403 (N_1403,N_372,N_619);
and U1404 (N_1404,N_295,N_131);
and U1405 (N_1405,N_840,N_246);
or U1406 (N_1406,N_781,N_614);
nand U1407 (N_1407,N_793,N_799);
or U1408 (N_1408,N_63,N_746);
or U1409 (N_1409,N_556,N_144);
nand U1410 (N_1410,N_396,N_610);
and U1411 (N_1411,N_911,N_606);
nor U1412 (N_1412,N_977,N_113);
nor U1413 (N_1413,N_260,N_24);
xnor U1414 (N_1414,N_779,N_872);
and U1415 (N_1415,N_958,N_807);
or U1416 (N_1416,N_617,N_581);
xor U1417 (N_1417,N_949,N_205);
nand U1418 (N_1418,N_213,N_452);
nand U1419 (N_1419,N_661,N_152);
xnor U1420 (N_1420,N_448,N_613);
and U1421 (N_1421,N_937,N_648);
and U1422 (N_1422,N_106,N_516);
nand U1423 (N_1423,N_112,N_3);
and U1424 (N_1424,N_385,N_199);
nor U1425 (N_1425,N_254,N_329);
nor U1426 (N_1426,N_458,N_243);
or U1427 (N_1427,N_322,N_308);
nor U1428 (N_1428,N_86,N_955);
nor U1429 (N_1429,N_820,N_8);
nand U1430 (N_1430,N_239,N_1);
or U1431 (N_1431,N_592,N_825);
nand U1432 (N_1432,N_174,N_376);
and U1433 (N_1433,N_907,N_464);
or U1434 (N_1434,N_480,N_769);
nand U1435 (N_1435,N_798,N_795);
or U1436 (N_1436,N_963,N_511);
and U1437 (N_1437,N_625,N_901);
and U1438 (N_1438,N_763,N_726);
nand U1439 (N_1439,N_599,N_883);
and U1440 (N_1440,N_444,N_743);
nand U1441 (N_1441,N_262,N_77);
or U1442 (N_1442,N_411,N_651);
or U1443 (N_1443,N_934,N_300);
or U1444 (N_1444,N_525,N_248);
nand U1445 (N_1445,N_25,N_6);
nor U1446 (N_1446,N_995,N_211);
and U1447 (N_1447,N_562,N_893);
nor U1448 (N_1448,N_878,N_327);
nand U1449 (N_1449,N_620,N_823);
and U1450 (N_1450,N_693,N_573);
nand U1451 (N_1451,N_796,N_731);
nand U1452 (N_1452,N_11,N_837);
or U1453 (N_1453,N_212,N_985);
nand U1454 (N_1454,N_190,N_414);
and U1455 (N_1455,N_290,N_679);
nor U1456 (N_1456,N_142,N_593);
or U1457 (N_1457,N_296,N_143);
nand U1458 (N_1458,N_315,N_159);
xor U1459 (N_1459,N_352,N_538);
nor U1460 (N_1460,N_590,N_935);
nand U1461 (N_1461,N_52,N_96);
nand U1462 (N_1462,N_430,N_177);
nor U1463 (N_1463,N_483,N_172);
nand U1464 (N_1464,N_381,N_918);
and U1465 (N_1465,N_313,N_494);
or U1466 (N_1466,N_912,N_132);
or U1467 (N_1467,N_579,N_194);
xnor U1468 (N_1468,N_938,N_898);
nand U1469 (N_1469,N_634,N_364);
nand U1470 (N_1470,N_489,N_638);
or U1471 (N_1471,N_607,N_970);
or U1472 (N_1472,N_509,N_804);
and U1473 (N_1473,N_686,N_954);
nor U1474 (N_1474,N_681,N_224);
nor U1475 (N_1475,N_851,N_394);
xnor U1476 (N_1476,N_192,N_378);
or U1477 (N_1477,N_487,N_646);
nor U1478 (N_1478,N_723,N_811);
nand U1479 (N_1479,N_269,N_822);
or U1480 (N_1480,N_467,N_81);
and U1481 (N_1481,N_165,N_155);
nor U1482 (N_1482,N_216,N_657);
or U1483 (N_1483,N_453,N_762);
or U1484 (N_1484,N_999,N_214);
nand U1485 (N_1485,N_881,N_336);
nor U1486 (N_1486,N_271,N_717);
and U1487 (N_1487,N_682,N_299);
or U1488 (N_1488,N_976,N_306);
nand U1489 (N_1489,N_678,N_167);
and U1490 (N_1490,N_927,N_529);
nor U1491 (N_1491,N_583,N_730);
nand U1492 (N_1492,N_546,N_774);
nand U1493 (N_1493,N_568,N_355);
or U1494 (N_1494,N_608,N_457);
and U1495 (N_1495,N_742,N_363);
or U1496 (N_1496,N_223,N_979);
and U1497 (N_1497,N_145,N_477);
nand U1498 (N_1498,N_915,N_449);
and U1499 (N_1499,N_815,N_293);
nand U1500 (N_1500,N_498,N_884);
and U1501 (N_1501,N_925,N_919);
nor U1502 (N_1502,N_302,N_301);
nor U1503 (N_1503,N_40,N_919);
nand U1504 (N_1504,N_190,N_895);
nand U1505 (N_1505,N_525,N_637);
nor U1506 (N_1506,N_412,N_662);
and U1507 (N_1507,N_698,N_867);
and U1508 (N_1508,N_332,N_545);
xor U1509 (N_1509,N_28,N_362);
nand U1510 (N_1510,N_585,N_769);
nand U1511 (N_1511,N_940,N_430);
and U1512 (N_1512,N_105,N_658);
and U1513 (N_1513,N_499,N_677);
and U1514 (N_1514,N_592,N_636);
and U1515 (N_1515,N_88,N_759);
or U1516 (N_1516,N_484,N_725);
nand U1517 (N_1517,N_647,N_26);
or U1518 (N_1518,N_879,N_748);
or U1519 (N_1519,N_319,N_298);
and U1520 (N_1520,N_765,N_296);
nor U1521 (N_1521,N_126,N_58);
and U1522 (N_1522,N_933,N_879);
nand U1523 (N_1523,N_514,N_358);
and U1524 (N_1524,N_229,N_84);
nor U1525 (N_1525,N_26,N_673);
nand U1526 (N_1526,N_916,N_9);
or U1527 (N_1527,N_470,N_578);
and U1528 (N_1528,N_494,N_475);
nand U1529 (N_1529,N_378,N_702);
or U1530 (N_1530,N_634,N_36);
nor U1531 (N_1531,N_873,N_649);
or U1532 (N_1532,N_108,N_417);
and U1533 (N_1533,N_848,N_612);
or U1534 (N_1534,N_407,N_551);
nor U1535 (N_1535,N_812,N_111);
xnor U1536 (N_1536,N_132,N_633);
and U1537 (N_1537,N_997,N_378);
and U1538 (N_1538,N_296,N_723);
nor U1539 (N_1539,N_6,N_507);
nand U1540 (N_1540,N_367,N_984);
or U1541 (N_1541,N_814,N_552);
xor U1542 (N_1542,N_637,N_628);
and U1543 (N_1543,N_612,N_695);
and U1544 (N_1544,N_558,N_180);
nand U1545 (N_1545,N_705,N_877);
and U1546 (N_1546,N_600,N_929);
and U1547 (N_1547,N_468,N_524);
nor U1548 (N_1548,N_105,N_334);
xor U1549 (N_1549,N_104,N_425);
and U1550 (N_1550,N_314,N_678);
nor U1551 (N_1551,N_971,N_208);
xor U1552 (N_1552,N_663,N_832);
nor U1553 (N_1553,N_583,N_208);
and U1554 (N_1554,N_460,N_938);
and U1555 (N_1555,N_181,N_83);
nor U1556 (N_1556,N_657,N_939);
and U1557 (N_1557,N_536,N_228);
and U1558 (N_1558,N_925,N_104);
or U1559 (N_1559,N_422,N_242);
nor U1560 (N_1560,N_490,N_910);
nor U1561 (N_1561,N_962,N_489);
or U1562 (N_1562,N_709,N_490);
and U1563 (N_1563,N_981,N_328);
or U1564 (N_1564,N_342,N_373);
and U1565 (N_1565,N_587,N_161);
or U1566 (N_1566,N_674,N_309);
and U1567 (N_1567,N_116,N_999);
and U1568 (N_1568,N_882,N_697);
xnor U1569 (N_1569,N_183,N_151);
and U1570 (N_1570,N_750,N_483);
nand U1571 (N_1571,N_674,N_57);
and U1572 (N_1572,N_602,N_213);
or U1573 (N_1573,N_942,N_491);
and U1574 (N_1574,N_60,N_460);
and U1575 (N_1575,N_255,N_856);
and U1576 (N_1576,N_227,N_150);
or U1577 (N_1577,N_215,N_970);
and U1578 (N_1578,N_615,N_544);
nand U1579 (N_1579,N_602,N_682);
and U1580 (N_1580,N_679,N_120);
or U1581 (N_1581,N_760,N_433);
nor U1582 (N_1582,N_75,N_738);
or U1583 (N_1583,N_551,N_581);
or U1584 (N_1584,N_378,N_970);
and U1585 (N_1585,N_631,N_702);
and U1586 (N_1586,N_39,N_207);
and U1587 (N_1587,N_2,N_747);
or U1588 (N_1588,N_387,N_457);
and U1589 (N_1589,N_233,N_980);
and U1590 (N_1590,N_102,N_61);
or U1591 (N_1591,N_347,N_92);
and U1592 (N_1592,N_229,N_598);
xnor U1593 (N_1593,N_25,N_640);
nand U1594 (N_1594,N_952,N_601);
or U1595 (N_1595,N_927,N_909);
nand U1596 (N_1596,N_24,N_232);
nand U1597 (N_1597,N_975,N_248);
nor U1598 (N_1598,N_352,N_829);
xor U1599 (N_1599,N_442,N_820);
or U1600 (N_1600,N_556,N_242);
nand U1601 (N_1601,N_12,N_950);
and U1602 (N_1602,N_40,N_718);
nor U1603 (N_1603,N_399,N_848);
nand U1604 (N_1604,N_44,N_894);
and U1605 (N_1605,N_595,N_742);
and U1606 (N_1606,N_611,N_911);
or U1607 (N_1607,N_815,N_205);
nand U1608 (N_1608,N_962,N_185);
or U1609 (N_1609,N_139,N_796);
or U1610 (N_1610,N_69,N_527);
nand U1611 (N_1611,N_957,N_802);
nor U1612 (N_1612,N_210,N_988);
nand U1613 (N_1613,N_156,N_40);
nand U1614 (N_1614,N_164,N_646);
nand U1615 (N_1615,N_186,N_67);
nor U1616 (N_1616,N_365,N_747);
or U1617 (N_1617,N_906,N_775);
xor U1618 (N_1618,N_802,N_412);
and U1619 (N_1619,N_399,N_486);
nand U1620 (N_1620,N_752,N_985);
nand U1621 (N_1621,N_631,N_85);
nor U1622 (N_1622,N_92,N_752);
and U1623 (N_1623,N_927,N_630);
and U1624 (N_1624,N_453,N_888);
or U1625 (N_1625,N_455,N_605);
nand U1626 (N_1626,N_733,N_90);
and U1627 (N_1627,N_395,N_323);
or U1628 (N_1628,N_198,N_297);
and U1629 (N_1629,N_475,N_446);
nor U1630 (N_1630,N_832,N_980);
xnor U1631 (N_1631,N_967,N_523);
and U1632 (N_1632,N_20,N_721);
nand U1633 (N_1633,N_365,N_506);
nand U1634 (N_1634,N_392,N_338);
and U1635 (N_1635,N_103,N_75);
and U1636 (N_1636,N_192,N_603);
nor U1637 (N_1637,N_709,N_254);
and U1638 (N_1638,N_526,N_992);
xnor U1639 (N_1639,N_94,N_862);
xor U1640 (N_1640,N_312,N_951);
or U1641 (N_1641,N_149,N_16);
and U1642 (N_1642,N_165,N_112);
or U1643 (N_1643,N_624,N_767);
or U1644 (N_1644,N_876,N_466);
xor U1645 (N_1645,N_919,N_386);
nor U1646 (N_1646,N_346,N_515);
or U1647 (N_1647,N_64,N_932);
and U1648 (N_1648,N_26,N_959);
nand U1649 (N_1649,N_433,N_79);
or U1650 (N_1650,N_240,N_571);
or U1651 (N_1651,N_458,N_207);
and U1652 (N_1652,N_878,N_834);
and U1653 (N_1653,N_412,N_770);
nor U1654 (N_1654,N_899,N_311);
nand U1655 (N_1655,N_783,N_76);
nand U1656 (N_1656,N_497,N_912);
or U1657 (N_1657,N_584,N_867);
and U1658 (N_1658,N_25,N_270);
or U1659 (N_1659,N_646,N_633);
nor U1660 (N_1660,N_27,N_796);
nand U1661 (N_1661,N_789,N_651);
xor U1662 (N_1662,N_469,N_688);
or U1663 (N_1663,N_445,N_274);
and U1664 (N_1664,N_395,N_789);
or U1665 (N_1665,N_830,N_826);
nand U1666 (N_1666,N_328,N_301);
nor U1667 (N_1667,N_272,N_90);
and U1668 (N_1668,N_966,N_548);
or U1669 (N_1669,N_801,N_599);
nand U1670 (N_1670,N_265,N_616);
or U1671 (N_1671,N_88,N_768);
nand U1672 (N_1672,N_915,N_178);
nor U1673 (N_1673,N_538,N_84);
and U1674 (N_1674,N_480,N_328);
nand U1675 (N_1675,N_699,N_794);
nor U1676 (N_1676,N_911,N_641);
nand U1677 (N_1677,N_354,N_836);
nand U1678 (N_1678,N_27,N_718);
or U1679 (N_1679,N_949,N_310);
nand U1680 (N_1680,N_45,N_611);
and U1681 (N_1681,N_832,N_996);
xor U1682 (N_1682,N_716,N_136);
or U1683 (N_1683,N_336,N_642);
nor U1684 (N_1684,N_949,N_430);
or U1685 (N_1685,N_358,N_7);
nor U1686 (N_1686,N_572,N_347);
or U1687 (N_1687,N_785,N_377);
and U1688 (N_1688,N_40,N_311);
nand U1689 (N_1689,N_75,N_709);
nand U1690 (N_1690,N_547,N_945);
or U1691 (N_1691,N_100,N_86);
or U1692 (N_1692,N_251,N_840);
and U1693 (N_1693,N_820,N_859);
nand U1694 (N_1694,N_676,N_131);
and U1695 (N_1695,N_815,N_472);
nor U1696 (N_1696,N_21,N_562);
nor U1697 (N_1697,N_116,N_165);
nand U1698 (N_1698,N_98,N_954);
or U1699 (N_1699,N_447,N_575);
nand U1700 (N_1700,N_60,N_914);
nor U1701 (N_1701,N_1,N_435);
nor U1702 (N_1702,N_661,N_985);
and U1703 (N_1703,N_8,N_673);
nor U1704 (N_1704,N_696,N_978);
or U1705 (N_1705,N_105,N_737);
nand U1706 (N_1706,N_386,N_495);
nand U1707 (N_1707,N_891,N_336);
nand U1708 (N_1708,N_108,N_921);
and U1709 (N_1709,N_703,N_408);
nand U1710 (N_1710,N_608,N_160);
and U1711 (N_1711,N_2,N_309);
nand U1712 (N_1712,N_151,N_456);
and U1713 (N_1713,N_581,N_727);
and U1714 (N_1714,N_82,N_375);
nor U1715 (N_1715,N_196,N_391);
and U1716 (N_1716,N_4,N_968);
or U1717 (N_1717,N_648,N_82);
nand U1718 (N_1718,N_823,N_228);
or U1719 (N_1719,N_738,N_817);
nand U1720 (N_1720,N_924,N_868);
xor U1721 (N_1721,N_569,N_554);
xor U1722 (N_1722,N_767,N_586);
and U1723 (N_1723,N_73,N_448);
nand U1724 (N_1724,N_441,N_631);
nor U1725 (N_1725,N_955,N_671);
or U1726 (N_1726,N_875,N_34);
or U1727 (N_1727,N_63,N_739);
nor U1728 (N_1728,N_513,N_356);
nor U1729 (N_1729,N_779,N_414);
xor U1730 (N_1730,N_640,N_914);
nand U1731 (N_1731,N_420,N_699);
nand U1732 (N_1732,N_249,N_357);
nor U1733 (N_1733,N_75,N_701);
nand U1734 (N_1734,N_9,N_562);
nand U1735 (N_1735,N_62,N_687);
nand U1736 (N_1736,N_405,N_879);
nor U1737 (N_1737,N_912,N_70);
or U1738 (N_1738,N_151,N_788);
nand U1739 (N_1739,N_696,N_993);
or U1740 (N_1740,N_127,N_790);
nand U1741 (N_1741,N_64,N_250);
and U1742 (N_1742,N_119,N_378);
or U1743 (N_1743,N_861,N_989);
nor U1744 (N_1744,N_925,N_472);
or U1745 (N_1745,N_178,N_685);
or U1746 (N_1746,N_263,N_739);
nor U1747 (N_1747,N_484,N_326);
nor U1748 (N_1748,N_321,N_696);
nand U1749 (N_1749,N_931,N_455);
and U1750 (N_1750,N_305,N_470);
xnor U1751 (N_1751,N_251,N_495);
or U1752 (N_1752,N_538,N_271);
or U1753 (N_1753,N_591,N_676);
xnor U1754 (N_1754,N_317,N_231);
and U1755 (N_1755,N_940,N_40);
and U1756 (N_1756,N_850,N_926);
and U1757 (N_1757,N_117,N_689);
xnor U1758 (N_1758,N_496,N_167);
nor U1759 (N_1759,N_935,N_446);
nor U1760 (N_1760,N_494,N_42);
xnor U1761 (N_1761,N_66,N_51);
and U1762 (N_1762,N_254,N_455);
nor U1763 (N_1763,N_829,N_397);
nor U1764 (N_1764,N_253,N_974);
xnor U1765 (N_1765,N_573,N_575);
nand U1766 (N_1766,N_454,N_14);
or U1767 (N_1767,N_893,N_523);
nor U1768 (N_1768,N_504,N_650);
nor U1769 (N_1769,N_373,N_830);
nand U1770 (N_1770,N_828,N_11);
nand U1771 (N_1771,N_917,N_511);
nor U1772 (N_1772,N_706,N_24);
or U1773 (N_1773,N_688,N_134);
nor U1774 (N_1774,N_693,N_170);
or U1775 (N_1775,N_505,N_877);
nor U1776 (N_1776,N_584,N_536);
or U1777 (N_1777,N_453,N_615);
nand U1778 (N_1778,N_67,N_861);
nand U1779 (N_1779,N_887,N_747);
or U1780 (N_1780,N_73,N_878);
nor U1781 (N_1781,N_801,N_311);
and U1782 (N_1782,N_941,N_401);
and U1783 (N_1783,N_192,N_607);
nand U1784 (N_1784,N_234,N_774);
and U1785 (N_1785,N_624,N_736);
and U1786 (N_1786,N_403,N_443);
nor U1787 (N_1787,N_432,N_883);
or U1788 (N_1788,N_955,N_885);
or U1789 (N_1789,N_256,N_311);
or U1790 (N_1790,N_974,N_84);
nor U1791 (N_1791,N_65,N_135);
nand U1792 (N_1792,N_647,N_696);
or U1793 (N_1793,N_758,N_281);
and U1794 (N_1794,N_525,N_178);
and U1795 (N_1795,N_117,N_108);
or U1796 (N_1796,N_652,N_289);
nand U1797 (N_1797,N_878,N_3);
and U1798 (N_1798,N_82,N_37);
and U1799 (N_1799,N_7,N_353);
and U1800 (N_1800,N_199,N_81);
or U1801 (N_1801,N_198,N_489);
nand U1802 (N_1802,N_204,N_624);
nand U1803 (N_1803,N_970,N_833);
nor U1804 (N_1804,N_115,N_490);
nor U1805 (N_1805,N_134,N_708);
nand U1806 (N_1806,N_518,N_578);
nand U1807 (N_1807,N_963,N_162);
nor U1808 (N_1808,N_86,N_567);
and U1809 (N_1809,N_785,N_777);
nand U1810 (N_1810,N_652,N_648);
or U1811 (N_1811,N_921,N_231);
or U1812 (N_1812,N_169,N_251);
or U1813 (N_1813,N_540,N_58);
or U1814 (N_1814,N_959,N_461);
or U1815 (N_1815,N_502,N_557);
nor U1816 (N_1816,N_155,N_350);
nand U1817 (N_1817,N_317,N_849);
nand U1818 (N_1818,N_137,N_782);
nor U1819 (N_1819,N_819,N_838);
nand U1820 (N_1820,N_711,N_78);
nand U1821 (N_1821,N_799,N_881);
nand U1822 (N_1822,N_268,N_158);
xnor U1823 (N_1823,N_137,N_853);
or U1824 (N_1824,N_227,N_21);
xnor U1825 (N_1825,N_405,N_185);
or U1826 (N_1826,N_7,N_343);
nand U1827 (N_1827,N_741,N_146);
or U1828 (N_1828,N_724,N_752);
or U1829 (N_1829,N_164,N_239);
or U1830 (N_1830,N_89,N_37);
nand U1831 (N_1831,N_821,N_35);
nand U1832 (N_1832,N_374,N_487);
nand U1833 (N_1833,N_478,N_443);
nor U1834 (N_1834,N_106,N_730);
and U1835 (N_1835,N_450,N_315);
or U1836 (N_1836,N_141,N_913);
xnor U1837 (N_1837,N_987,N_298);
nand U1838 (N_1838,N_416,N_778);
nand U1839 (N_1839,N_552,N_642);
and U1840 (N_1840,N_845,N_687);
and U1841 (N_1841,N_632,N_617);
and U1842 (N_1842,N_865,N_508);
nand U1843 (N_1843,N_844,N_224);
nand U1844 (N_1844,N_582,N_937);
and U1845 (N_1845,N_826,N_978);
xor U1846 (N_1846,N_771,N_89);
xnor U1847 (N_1847,N_83,N_806);
xnor U1848 (N_1848,N_332,N_813);
or U1849 (N_1849,N_339,N_68);
and U1850 (N_1850,N_556,N_714);
or U1851 (N_1851,N_285,N_845);
nor U1852 (N_1852,N_140,N_194);
and U1853 (N_1853,N_97,N_54);
or U1854 (N_1854,N_321,N_492);
xnor U1855 (N_1855,N_24,N_28);
or U1856 (N_1856,N_113,N_769);
and U1857 (N_1857,N_648,N_670);
nor U1858 (N_1858,N_800,N_351);
nand U1859 (N_1859,N_46,N_420);
and U1860 (N_1860,N_504,N_362);
xnor U1861 (N_1861,N_726,N_935);
and U1862 (N_1862,N_726,N_66);
nor U1863 (N_1863,N_594,N_614);
and U1864 (N_1864,N_735,N_167);
xnor U1865 (N_1865,N_772,N_118);
nand U1866 (N_1866,N_555,N_501);
nor U1867 (N_1867,N_974,N_247);
nand U1868 (N_1868,N_621,N_837);
or U1869 (N_1869,N_872,N_279);
nand U1870 (N_1870,N_636,N_942);
and U1871 (N_1871,N_213,N_425);
xor U1872 (N_1872,N_926,N_70);
and U1873 (N_1873,N_629,N_83);
or U1874 (N_1874,N_23,N_615);
nor U1875 (N_1875,N_634,N_644);
nand U1876 (N_1876,N_589,N_575);
nand U1877 (N_1877,N_603,N_751);
nor U1878 (N_1878,N_481,N_923);
nor U1879 (N_1879,N_587,N_107);
nor U1880 (N_1880,N_529,N_267);
or U1881 (N_1881,N_859,N_714);
xor U1882 (N_1882,N_633,N_913);
nand U1883 (N_1883,N_29,N_556);
nor U1884 (N_1884,N_911,N_462);
nand U1885 (N_1885,N_316,N_634);
and U1886 (N_1886,N_578,N_58);
nor U1887 (N_1887,N_980,N_22);
nor U1888 (N_1888,N_157,N_590);
nand U1889 (N_1889,N_598,N_142);
nand U1890 (N_1890,N_826,N_981);
xor U1891 (N_1891,N_721,N_101);
nand U1892 (N_1892,N_887,N_111);
nand U1893 (N_1893,N_419,N_263);
or U1894 (N_1894,N_820,N_761);
nor U1895 (N_1895,N_275,N_349);
nor U1896 (N_1896,N_764,N_243);
nor U1897 (N_1897,N_787,N_706);
or U1898 (N_1898,N_69,N_317);
or U1899 (N_1899,N_776,N_37);
nor U1900 (N_1900,N_59,N_532);
nand U1901 (N_1901,N_415,N_70);
nand U1902 (N_1902,N_626,N_826);
nor U1903 (N_1903,N_330,N_508);
and U1904 (N_1904,N_34,N_568);
and U1905 (N_1905,N_841,N_468);
nand U1906 (N_1906,N_531,N_635);
and U1907 (N_1907,N_975,N_221);
nand U1908 (N_1908,N_942,N_861);
nor U1909 (N_1909,N_433,N_51);
nor U1910 (N_1910,N_551,N_805);
or U1911 (N_1911,N_399,N_378);
nor U1912 (N_1912,N_39,N_767);
nor U1913 (N_1913,N_471,N_265);
xnor U1914 (N_1914,N_423,N_194);
nand U1915 (N_1915,N_597,N_961);
nor U1916 (N_1916,N_797,N_192);
or U1917 (N_1917,N_711,N_91);
and U1918 (N_1918,N_909,N_590);
nor U1919 (N_1919,N_963,N_461);
nor U1920 (N_1920,N_191,N_284);
nor U1921 (N_1921,N_335,N_895);
and U1922 (N_1922,N_913,N_423);
nand U1923 (N_1923,N_872,N_733);
or U1924 (N_1924,N_1,N_620);
nor U1925 (N_1925,N_575,N_810);
nand U1926 (N_1926,N_105,N_872);
or U1927 (N_1927,N_807,N_534);
nand U1928 (N_1928,N_850,N_516);
and U1929 (N_1929,N_761,N_834);
nand U1930 (N_1930,N_461,N_669);
or U1931 (N_1931,N_65,N_741);
nor U1932 (N_1932,N_280,N_963);
nand U1933 (N_1933,N_793,N_539);
xnor U1934 (N_1934,N_97,N_902);
nor U1935 (N_1935,N_531,N_154);
nand U1936 (N_1936,N_689,N_253);
and U1937 (N_1937,N_298,N_271);
xnor U1938 (N_1938,N_351,N_719);
and U1939 (N_1939,N_561,N_722);
and U1940 (N_1940,N_874,N_204);
and U1941 (N_1941,N_986,N_136);
xor U1942 (N_1942,N_653,N_506);
and U1943 (N_1943,N_352,N_395);
nor U1944 (N_1944,N_691,N_910);
nand U1945 (N_1945,N_798,N_773);
and U1946 (N_1946,N_645,N_556);
nor U1947 (N_1947,N_836,N_210);
nand U1948 (N_1948,N_932,N_972);
nor U1949 (N_1949,N_772,N_918);
nor U1950 (N_1950,N_864,N_428);
nand U1951 (N_1951,N_118,N_310);
xnor U1952 (N_1952,N_216,N_718);
and U1953 (N_1953,N_653,N_843);
and U1954 (N_1954,N_309,N_868);
nor U1955 (N_1955,N_94,N_786);
and U1956 (N_1956,N_373,N_646);
nand U1957 (N_1957,N_134,N_946);
or U1958 (N_1958,N_137,N_408);
or U1959 (N_1959,N_650,N_837);
nor U1960 (N_1960,N_649,N_549);
nor U1961 (N_1961,N_833,N_297);
and U1962 (N_1962,N_653,N_463);
or U1963 (N_1963,N_720,N_639);
nor U1964 (N_1964,N_582,N_602);
or U1965 (N_1965,N_634,N_817);
nand U1966 (N_1966,N_723,N_487);
nor U1967 (N_1967,N_301,N_942);
nor U1968 (N_1968,N_747,N_954);
nor U1969 (N_1969,N_5,N_298);
xor U1970 (N_1970,N_458,N_858);
and U1971 (N_1971,N_138,N_451);
nand U1972 (N_1972,N_887,N_602);
nor U1973 (N_1973,N_565,N_263);
nand U1974 (N_1974,N_840,N_592);
nand U1975 (N_1975,N_44,N_887);
nor U1976 (N_1976,N_248,N_68);
and U1977 (N_1977,N_34,N_950);
nand U1978 (N_1978,N_361,N_514);
nor U1979 (N_1979,N_151,N_445);
and U1980 (N_1980,N_663,N_977);
and U1981 (N_1981,N_278,N_88);
and U1982 (N_1982,N_132,N_579);
nand U1983 (N_1983,N_89,N_661);
xor U1984 (N_1984,N_734,N_122);
nand U1985 (N_1985,N_215,N_68);
nand U1986 (N_1986,N_5,N_519);
and U1987 (N_1987,N_859,N_239);
and U1988 (N_1988,N_657,N_529);
nand U1989 (N_1989,N_27,N_730);
xor U1990 (N_1990,N_556,N_53);
nor U1991 (N_1991,N_720,N_581);
nor U1992 (N_1992,N_538,N_228);
and U1993 (N_1993,N_32,N_618);
and U1994 (N_1994,N_201,N_521);
or U1995 (N_1995,N_226,N_280);
xor U1996 (N_1996,N_497,N_15);
and U1997 (N_1997,N_472,N_714);
nor U1998 (N_1998,N_788,N_94);
nand U1999 (N_1999,N_585,N_641);
or U2000 (N_2000,N_1510,N_1378);
and U2001 (N_2001,N_1201,N_1120);
nor U2002 (N_2002,N_1054,N_1333);
and U2003 (N_2003,N_1039,N_1462);
nand U2004 (N_2004,N_1211,N_1920);
nand U2005 (N_2005,N_1259,N_1401);
and U2006 (N_2006,N_1800,N_1826);
nor U2007 (N_2007,N_1816,N_1564);
or U2008 (N_2008,N_1310,N_1690);
and U2009 (N_2009,N_1587,N_1523);
or U2010 (N_2010,N_1829,N_1136);
and U2011 (N_2011,N_1827,N_1192);
or U2012 (N_2012,N_1285,N_1659);
and U2013 (N_2013,N_1427,N_1700);
xor U2014 (N_2014,N_1075,N_1250);
nand U2015 (N_2015,N_1731,N_1871);
and U2016 (N_2016,N_1802,N_1282);
nand U2017 (N_2017,N_1594,N_1189);
or U2018 (N_2018,N_1193,N_1864);
and U2019 (N_2019,N_1957,N_1517);
nor U2020 (N_2020,N_1290,N_1820);
nor U2021 (N_2021,N_1768,N_1244);
nor U2022 (N_2022,N_1420,N_1933);
and U2023 (N_2023,N_1653,N_1545);
nor U2024 (N_2024,N_1955,N_1058);
nand U2025 (N_2025,N_1279,N_1844);
nand U2026 (N_2026,N_1969,N_1086);
or U2027 (N_2027,N_1603,N_1437);
nor U2028 (N_2028,N_1887,N_1410);
and U2029 (N_2029,N_1724,N_1038);
nor U2030 (N_2030,N_1552,N_1286);
and U2031 (N_2031,N_1614,N_1831);
and U2032 (N_2032,N_1861,N_1952);
nand U2033 (N_2033,N_1267,N_1576);
or U2034 (N_2034,N_1238,N_1801);
or U2035 (N_2035,N_1509,N_1111);
or U2036 (N_2036,N_1818,N_1892);
nand U2037 (N_2037,N_1063,N_1563);
or U2038 (N_2038,N_1315,N_1258);
or U2039 (N_2039,N_1956,N_1155);
and U2040 (N_2040,N_1916,N_1703);
and U2041 (N_2041,N_1930,N_1766);
nand U2042 (N_2042,N_1464,N_1328);
and U2043 (N_2043,N_1675,N_1484);
nand U2044 (N_2044,N_1668,N_1584);
or U2045 (N_2045,N_1135,N_1036);
or U2046 (N_2046,N_1592,N_1886);
xnor U2047 (N_2047,N_1651,N_1536);
and U2048 (N_2048,N_1216,N_1405);
or U2049 (N_2049,N_1415,N_1301);
nor U2050 (N_2050,N_1667,N_1003);
nor U2051 (N_2051,N_1123,N_1775);
nand U2052 (N_2052,N_1072,N_1316);
nand U2053 (N_2053,N_1602,N_1317);
or U2054 (N_2054,N_1746,N_1689);
or U2055 (N_2055,N_1747,N_1237);
xnor U2056 (N_2056,N_1117,N_1839);
nor U2057 (N_2057,N_1591,N_1953);
nor U2058 (N_2058,N_1765,N_1336);
and U2059 (N_2059,N_1056,N_1247);
or U2060 (N_2060,N_1698,N_1254);
nand U2061 (N_2061,N_1434,N_1806);
nor U2062 (N_2062,N_1781,N_1882);
and U2063 (N_2063,N_1736,N_1388);
or U2064 (N_2064,N_1044,N_1593);
and U2065 (N_2065,N_1113,N_1265);
nor U2066 (N_2066,N_1283,N_1202);
nor U2067 (N_2067,N_1455,N_1977);
xnor U2068 (N_2068,N_1028,N_1187);
and U2069 (N_2069,N_1959,N_1449);
and U2070 (N_2070,N_1496,N_1419);
nand U2071 (N_2071,N_1218,N_1494);
xor U2072 (N_2072,N_1233,N_1371);
and U2073 (N_2073,N_1191,N_1574);
xnor U2074 (N_2074,N_1146,N_1467);
and U2075 (N_2075,N_1092,N_1624);
or U2076 (N_2076,N_1425,N_1495);
xor U2077 (N_2077,N_1701,N_1376);
nand U2078 (N_2078,N_1795,N_1853);
nand U2079 (N_2079,N_1209,N_1207);
nand U2080 (N_2080,N_1666,N_1981);
or U2081 (N_2081,N_1224,N_1068);
nor U2082 (N_2082,N_1059,N_1687);
nand U2083 (N_2083,N_1786,N_1069);
xnor U2084 (N_2084,N_1791,N_1688);
or U2085 (N_2085,N_1253,N_1715);
or U2086 (N_2086,N_1983,N_1100);
or U2087 (N_2087,N_1012,N_1513);
nor U2088 (N_2088,N_1526,N_1463);
nand U2089 (N_2089,N_1106,N_1011);
nand U2090 (N_2090,N_1714,N_1656);
nor U2091 (N_2091,N_1243,N_1280);
nor U2092 (N_2092,N_1423,N_1119);
nand U2093 (N_2093,N_1738,N_1447);
nand U2094 (N_2094,N_1035,N_1629);
nor U2095 (N_2095,N_1379,N_1020);
or U2096 (N_2096,N_1612,N_1256);
or U2097 (N_2097,N_1384,N_1077);
and U2098 (N_2098,N_1176,N_1348);
nor U2099 (N_2099,N_1809,N_1091);
nand U2100 (N_2100,N_1524,N_1677);
or U2101 (N_2101,N_1099,N_1712);
nand U2102 (N_2102,N_1108,N_1852);
or U2103 (N_2103,N_1654,N_1836);
nand U2104 (N_2104,N_1445,N_1974);
and U2105 (N_2105,N_1421,N_1922);
nor U2106 (N_2106,N_1570,N_1598);
and U2107 (N_2107,N_1787,N_1352);
nand U2108 (N_2108,N_1580,N_1025);
nor U2109 (N_2109,N_1021,N_1184);
or U2110 (N_2110,N_1723,N_1777);
and U2111 (N_2111,N_1792,N_1895);
nor U2112 (N_2112,N_1506,N_1159);
nand U2113 (N_2113,N_1263,N_1620);
or U2114 (N_2114,N_1302,N_1917);
and U2115 (N_2115,N_1569,N_1399);
nand U2116 (N_2116,N_1571,N_1982);
or U2117 (N_2117,N_1160,N_1018);
xor U2118 (N_2118,N_1753,N_1082);
xnor U2119 (N_2119,N_1344,N_1461);
nand U2120 (N_2120,N_1067,N_1903);
nand U2121 (N_2121,N_1085,N_1287);
and U2122 (N_2122,N_1845,N_1126);
nor U2123 (N_2123,N_1626,N_1133);
and U2124 (N_2124,N_1261,N_1305);
nand U2125 (N_2125,N_1230,N_1469);
or U2126 (N_2126,N_1572,N_1488);
nor U2127 (N_2127,N_1601,N_1772);
or U2128 (N_2128,N_1973,N_1718);
or U2129 (N_2129,N_1986,N_1755);
nor U2130 (N_2130,N_1595,N_1497);
xnor U2131 (N_2131,N_1522,N_1562);
and U2132 (N_2132,N_1949,N_1748);
nand U2133 (N_2133,N_1533,N_1181);
nand U2134 (N_2134,N_1431,N_1527);
or U2135 (N_2135,N_1931,N_1220);
nor U2136 (N_2136,N_1678,N_1101);
or U2137 (N_2137,N_1157,N_1749);
or U2138 (N_2138,N_1239,N_1942);
and U2139 (N_2139,N_1568,N_1112);
xor U2140 (N_2140,N_1650,N_1289);
or U2141 (N_2141,N_1671,N_1512);
nand U2142 (N_2142,N_1634,N_1177);
or U2143 (N_2143,N_1711,N_1630);
and U2144 (N_2144,N_1778,N_1492);
or U2145 (N_2145,N_1231,N_1550);
or U2146 (N_2146,N_1759,N_1362);
or U2147 (N_2147,N_1293,N_1727);
or U2148 (N_2148,N_1304,N_1166);
xnor U2149 (N_2149,N_1124,N_1297);
xor U2150 (N_2150,N_1888,N_1402);
and U2151 (N_2151,N_1869,N_1270);
and U2152 (N_2152,N_1409,N_1087);
or U2153 (N_2153,N_1234,N_1197);
or U2154 (N_2154,N_1334,N_1851);
and U2155 (N_2155,N_1141,N_1182);
or U2156 (N_2156,N_1742,N_1740);
nor U2157 (N_2157,N_1008,N_1648);
nand U2158 (N_2158,N_1432,N_1222);
nand U2159 (N_2159,N_1165,N_1782);
nor U2160 (N_2160,N_1394,N_1860);
nor U2161 (N_2161,N_1055,N_1451);
or U2162 (N_2162,N_1876,N_1936);
nand U2163 (N_2163,N_1185,N_1683);
nand U2164 (N_2164,N_1913,N_1862);
or U2165 (N_2165,N_1377,N_1456);
xnor U2166 (N_2166,N_1963,N_1728);
and U2167 (N_2167,N_1206,N_1422);
or U2168 (N_2168,N_1354,N_1453);
and U2169 (N_2169,N_1652,N_1565);
nor U2170 (N_2170,N_1383,N_1271);
nor U2171 (N_2171,N_1066,N_1487);
nand U2172 (N_2172,N_1313,N_1296);
and U2173 (N_2173,N_1590,N_1537);
nand U2174 (N_2174,N_1103,N_1705);
or U2175 (N_2175,N_1228,N_1483);
and U2176 (N_2176,N_1040,N_1979);
nand U2177 (N_2177,N_1118,N_1978);
nand U2178 (N_2178,N_1465,N_1625);
or U2179 (N_2179,N_1776,N_1885);
nand U2180 (N_2180,N_1902,N_1719);
or U2181 (N_2181,N_1906,N_1470);
and U2182 (N_2182,N_1618,N_1240);
or U2183 (N_2183,N_1442,N_1139);
nor U2184 (N_2184,N_1094,N_1713);
nor U2185 (N_2185,N_1874,N_1554);
or U2186 (N_2186,N_1636,N_1518);
or U2187 (N_2187,N_1414,N_1971);
and U2188 (N_2188,N_1169,N_1924);
nor U2189 (N_2189,N_1127,N_1985);
or U2190 (N_2190,N_1016,N_1918);
nand U2191 (N_2191,N_1529,N_1693);
or U2192 (N_2192,N_1345,N_1032);
or U2193 (N_2193,N_1142,N_1140);
and U2194 (N_2194,N_1551,N_1622);
or U2195 (N_2195,N_1941,N_1761);
or U2196 (N_2196,N_1684,N_1382);
or U2197 (N_2197,N_1796,N_1632);
and U2198 (N_2198,N_1850,N_1227);
nand U2199 (N_2199,N_1125,N_1443);
nand U2200 (N_2200,N_1349,N_1459);
and U2201 (N_2201,N_1122,N_1048);
or U2202 (N_2202,N_1084,N_1863);
and U2203 (N_2203,N_1751,N_1663);
nor U2204 (N_2204,N_1821,N_1739);
or U2205 (N_2205,N_1367,N_1951);
nor U2206 (N_2206,N_1799,N_1436);
nand U2207 (N_2207,N_1219,N_1696);
or U2208 (N_2208,N_1655,N_1406);
and U2209 (N_2209,N_1010,N_1001);
nand U2210 (N_2210,N_1346,N_1501);
nand U2211 (N_2211,N_1204,N_1961);
or U2212 (N_2212,N_1789,N_1466);
nor U2213 (N_2213,N_1438,N_1002);
or U2214 (N_2214,N_1249,N_1074);
nor U2215 (N_2215,N_1104,N_1407);
nor U2216 (N_2216,N_1843,N_1531);
xnor U2217 (N_2217,N_1132,N_1880);
nor U2218 (N_2218,N_1109,N_1288);
xnor U2219 (N_2219,N_1964,N_1060);
and U2220 (N_2220,N_1340,N_1832);
and U2221 (N_2221,N_1877,N_1045);
nand U2222 (N_2222,N_1278,N_1528);
nor U2223 (N_2223,N_1604,N_1901);
xnor U2224 (N_2224,N_1621,N_1923);
nand U2225 (N_2225,N_1446,N_1312);
nor U2226 (N_2226,N_1131,N_1398);
nand U2227 (N_2227,N_1392,N_1549);
nand U2228 (N_2228,N_1994,N_1566);
nor U2229 (N_2229,N_1031,N_1268);
xnor U2230 (N_2230,N_1426,N_1743);
xnor U2231 (N_2231,N_1514,N_1276);
nand U2232 (N_2232,N_1245,N_1217);
and U2233 (N_2233,N_1842,N_1006);
and U2234 (N_2234,N_1252,N_1695);
or U2235 (N_2235,N_1940,N_1321);
or U2236 (N_2236,N_1374,N_1670);
nand U2237 (N_2237,N_1645,N_1583);
or U2238 (N_2238,N_1788,N_1635);
and U2239 (N_2239,N_1559,N_1476);
nand U2240 (N_2240,N_1617,N_1685);
or U2241 (N_2241,N_1186,N_1548);
xor U2242 (N_2242,N_1105,N_1458);
and U2243 (N_2243,N_1539,N_1485);
or U2244 (N_2244,N_1733,N_1319);
and U2245 (N_2245,N_1337,N_1558);
nand U2246 (N_2246,N_1277,N_1229);
and U2247 (N_2247,N_1585,N_1413);
nor U2248 (N_2248,N_1642,N_1707);
nor U2249 (N_2249,N_1729,N_1946);
nand U2250 (N_2250,N_1049,N_1722);
or U2251 (N_2251,N_1052,N_1757);
xor U2252 (N_2252,N_1195,N_1291);
or U2253 (N_2253,N_1479,N_1295);
and U2254 (N_2254,N_1647,N_1534);
nor U2255 (N_2255,N_1014,N_1760);
nor U2256 (N_2256,N_1516,N_1359);
and U2257 (N_2257,N_1990,N_1855);
nand U2258 (N_2258,N_1669,N_1368);
and U2259 (N_2259,N_1573,N_1335);
nor U2260 (N_2260,N_1856,N_1215);
or U2261 (N_2261,N_1107,N_1174);
or U2262 (N_2262,N_1987,N_1318);
xor U2263 (N_2263,N_1947,N_1921);
nor U2264 (N_2264,N_1812,N_1454);
or U2265 (N_2265,N_1934,N_1780);
nor U2266 (N_2266,N_1898,N_1500);
nor U2267 (N_2267,N_1452,N_1486);
nor U2268 (N_2268,N_1331,N_1370);
nand U2269 (N_2269,N_1619,N_1638);
and U2270 (N_2270,N_1556,N_1793);
nor U2271 (N_2271,N_1322,N_1661);
nand U2272 (N_2272,N_1158,N_1081);
xor U2273 (N_2273,N_1730,N_1163);
nor U2274 (N_2274,N_1389,N_1199);
and U2275 (N_2275,N_1726,N_1457);
or U2276 (N_2276,N_1424,N_1530);
nand U2277 (N_2277,N_1395,N_1633);
and U2278 (N_2278,N_1897,N_1521);
nor U2279 (N_2279,N_1854,N_1950);
nor U2280 (N_2280,N_1332,N_1241);
or U2281 (N_2281,N_1435,N_1608);
xor U2282 (N_2282,N_1150,N_1676);
or U2283 (N_2283,N_1657,N_1721);
and U2284 (N_2284,N_1893,N_1269);
and U2285 (N_2285,N_1910,N_1073);
and U2286 (N_2286,N_1762,N_1752);
and U2287 (N_2287,N_1995,N_1363);
nor U2288 (N_2288,N_1369,N_1024);
and U2289 (N_2289,N_1027,N_1386);
or U2290 (N_2290,N_1543,N_1764);
nand U2291 (N_2291,N_1519,N_1779);
and U2292 (N_2292,N_1997,N_1507);
or U2293 (N_2293,N_1912,N_1212);
nand U2294 (N_2294,N_1699,N_1847);
nand U2295 (N_2295,N_1255,N_1029);
or U2296 (N_2296,N_1408,N_1682);
nor U2297 (N_2297,N_1720,N_1996);
or U2298 (N_2298,N_1857,N_1046);
nor U2299 (N_2299,N_1828,N_1393);
nand U2300 (N_2300,N_1062,N_1037);
nand U2301 (N_2301,N_1355,N_1605);
nor U2302 (N_2302,N_1970,N_1175);
and U2303 (N_2303,N_1915,N_1837);
xor U2304 (N_2304,N_1965,N_1623);
or U2305 (N_2305,N_1868,N_1147);
or U2306 (N_2306,N_1637,N_1129);
xnor U2307 (N_2307,N_1375,N_1783);
nand U2308 (N_2308,N_1292,N_1341);
and U2309 (N_2309,N_1889,N_1324);
xnor U2310 (N_2310,N_1498,N_1347);
nor U2311 (N_2311,N_1674,N_1515);
nor U2312 (N_2312,N_1520,N_1939);
nor U2313 (N_2313,N_1841,N_1050);
or U2314 (N_2314,N_1004,N_1342);
and U2315 (N_2315,N_1579,N_1803);
or U2316 (N_2316,N_1954,N_1351);
nor U2317 (N_2317,N_1366,N_1178);
nand U2318 (N_2318,N_1482,N_1905);
nor U2319 (N_2319,N_1875,N_1785);
or U2320 (N_2320,N_1859,N_1145);
nand U2321 (N_2321,N_1737,N_1691);
or U2322 (N_2322,N_1489,N_1274);
or U2323 (N_2323,N_1541,N_1967);
or U2324 (N_2324,N_1927,N_1872);
nor U2325 (N_2325,N_1089,N_1825);
or U2326 (N_2326,N_1908,N_1894);
nor U2327 (N_2327,N_1899,N_1242);
nand U2328 (N_2328,N_1441,N_1702);
nand U2329 (N_2329,N_1544,N_1833);
or U2330 (N_2330,N_1708,N_1444);
xor U2331 (N_2331,N_1555,N_1834);
nand U2332 (N_2332,N_1180,N_1148);
or U2333 (N_2333,N_1866,N_1391);
nand U2334 (N_2334,N_1450,N_1968);
nand U2335 (N_2335,N_1980,N_1013);
and U2336 (N_2336,N_1097,N_1798);
xor U2337 (N_2337,N_1744,N_1272);
and U2338 (N_2338,N_1628,N_1750);
or U2339 (N_2339,N_1116,N_1033);
or U2340 (N_2340,N_1311,N_1717);
nand U2341 (N_2341,N_1214,N_1611);
xnor U2342 (N_2342,N_1273,N_1194);
or U2343 (N_2343,N_1102,N_1814);
nor U2344 (N_2344,N_1472,N_1339);
xnor U2345 (N_2345,N_1198,N_1840);
or U2346 (N_2346,N_1115,N_1121);
nand U2347 (N_2347,N_1929,N_1606);
nor U2348 (N_2348,N_1473,N_1914);
nor U2349 (N_2349,N_1017,N_1298);
nand U2350 (N_2350,N_1599,N_1412);
xnor U2351 (N_2351,N_1043,N_1704);
or U2352 (N_2352,N_1538,N_1773);
and U2353 (N_2353,N_1071,N_1535);
and U2354 (N_2354,N_1835,N_1813);
or U2355 (N_2355,N_1439,N_1303);
nand U2356 (N_2356,N_1998,N_1525);
or U2357 (N_2357,N_1741,N_1480);
and U2358 (N_2358,N_1007,N_1962);
nand U2359 (N_2359,N_1716,N_1686);
or U2360 (N_2360,N_1190,N_1758);
and U2361 (N_2361,N_1428,N_1095);
or U2362 (N_2362,N_1532,N_1203);
nor U2363 (N_2363,N_1284,N_1658);
and U2364 (N_2364,N_1266,N_1810);
nor U2365 (N_2365,N_1468,N_1137);
nor U2366 (N_2366,N_1356,N_1323);
or U2367 (N_2367,N_1546,N_1096);
and U2368 (N_2368,N_1065,N_1560);
nand U2369 (N_2369,N_1053,N_1015);
nand U2370 (N_2370,N_1794,N_1478);
and U2371 (N_2371,N_1830,N_1080);
or U2372 (N_2372,N_1884,N_1665);
and U2373 (N_2373,N_1154,N_1948);
nor U2374 (N_2374,N_1338,N_1294);
and U2375 (N_2375,N_1372,N_1364);
nand U2376 (N_2376,N_1320,N_1070);
nor U2377 (N_2377,N_1999,N_1911);
and U2378 (N_2378,N_1090,N_1188);
nor U2379 (N_2379,N_1732,N_1083);
nor U2380 (N_2380,N_1078,N_1143);
or U2381 (N_2381,N_1815,N_1246);
and U2382 (N_2382,N_1925,N_1196);
xor U2383 (N_2383,N_1168,N_1361);
xnor U2384 (N_2384,N_1183,N_1225);
or U2385 (N_2385,N_1009,N_1330);
xor U2386 (N_2386,N_1314,N_1578);
nor U2387 (N_2387,N_1430,N_1173);
nor U2388 (N_2388,N_1022,N_1387);
nand U2389 (N_2389,N_1575,N_1975);
and U2390 (N_2390,N_1577,N_1325);
xnor U2391 (N_2391,N_1822,N_1047);
nor U2392 (N_2392,N_1681,N_1477);
nand U2393 (N_2393,N_1607,N_1891);
nor U2394 (N_2394,N_1380,N_1232);
or U2395 (N_2395,N_1542,N_1588);
or U2396 (N_2396,N_1172,N_1989);
nor U2397 (N_2397,N_1474,N_1680);
nor U2398 (N_2398,N_1460,N_1327);
nor U2399 (N_2399,N_1491,N_1260);
nand U2400 (N_2400,N_1631,N_1616);
nor U2401 (N_2401,N_1448,N_1756);
or U2402 (N_2402,N_1151,N_1932);
nand U2403 (N_2403,N_1030,N_1649);
and U2404 (N_2404,N_1672,N_1061);
or U2405 (N_2405,N_1000,N_1205);
or U2406 (N_2406,N_1943,N_1805);
and U2407 (N_2407,N_1471,N_1019);
and U2408 (N_2408,N_1213,N_1609);
or U2409 (N_2409,N_1023,N_1938);
or U2410 (N_2410,N_1926,N_1026);
or U2411 (N_2411,N_1493,N_1307);
nor U2412 (N_2412,N_1170,N_1846);
nor U2413 (N_2413,N_1919,N_1540);
and U2414 (N_2414,N_1397,N_1597);
or U2415 (N_2415,N_1396,N_1365);
nand U2416 (N_2416,N_1064,N_1694);
nand U2417 (N_2417,N_1966,N_1771);
xnor U2418 (N_2418,N_1144,N_1644);
and U2419 (N_2419,N_1403,N_1499);
nand U2420 (N_2420,N_1257,N_1804);
and U2421 (N_2421,N_1589,N_1329);
nand U2422 (N_2422,N_1041,N_1051);
or U2423 (N_2423,N_1679,N_1646);
or U2424 (N_2424,N_1504,N_1360);
or U2425 (N_2425,N_1935,N_1208);
or U2426 (N_2426,N_1418,N_1928);
or U2427 (N_2427,N_1808,N_1664);
nor U2428 (N_2428,N_1110,N_1817);
nor U2429 (N_2429,N_1156,N_1561);
nand U2430 (N_2430,N_1390,N_1904);
nand U2431 (N_2431,N_1896,N_1610);
nand U2432 (N_2432,N_1867,N_1130);
xnor U2433 (N_2433,N_1152,N_1660);
nor U2434 (N_2434,N_1508,N_1088);
nand U2435 (N_2435,N_1210,N_1076);
nor U2436 (N_2436,N_1138,N_1811);
nor U2437 (N_2437,N_1823,N_1153);
and U2438 (N_2438,N_1502,N_1945);
or U2439 (N_2439,N_1057,N_1824);
or U2440 (N_2440,N_1236,N_1343);
xnor U2441 (N_2441,N_1404,N_1162);
and U2442 (N_2442,N_1308,N_1769);
nand U2443 (N_2443,N_1221,N_1627);
and U2444 (N_2444,N_1640,N_1385);
nand U2445 (N_2445,N_1567,N_1890);
nand U2446 (N_2446,N_1878,N_1306);
nand U2447 (N_2447,N_1641,N_1264);
and U2448 (N_2448,N_1164,N_1400);
nor U2449 (N_2449,N_1582,N_1433);
nor U2450 (N_2450,N_1440,N_1774);
or U2451 (N_2451,N_1991,N_1960);
nand U2452 (N_2452,N_1300,N_1784);
or U2453 (N_2453,N_1958,N_1417);
nand U2454 (N_2454,N_1281,N_1819);
nor U2455 (N_2455,N_1235,N_1873);
and U2456 (N_2456,N_1993,N_1557);
and U2457 (N_2457,N_1511,N_1042);
and U2458 (N_2458,N_1770,N_1870);
nand U2459 (N_2459,N_1429,N_1639);
nor U2460 (N_2460,N_1988,N_1251);
and U2461 (N_2461,N_1161,N_1149);
or U2462 (N_2462,N_1128,N_1505);
nand U2463 (N_2463,N_1849,N_1807);
and U2464 (N_2464,N_1381,N_1790);
or U2465 (N_2465,N_1763,N_1248);
nand U2466 (N_2466,N_1879,N_1357);
nand U2467 (N_2467,N_1937,N_1179);
and U2468 (N_2468,N_1673,N_1503);
nand U2469 (N_2469,N_1171,N_1754);
nand U2470 (N_2470,N_1262,N_1838);
nor U2471 (N_2471,N_1547,N_1093);
nor U2472 (N_2472,N_1353,N_1299);
or U2473 (N_2473,N_1475,N_1883);
nor U2474 (N_2474,N_1992,N_1600);
and U2475 (N_2475,N_1697,N_1223);
and U2476 (N_2476,N_1907,N_1098);
xnor U2477 (N_2477,N_1167,N_1881);
nor U2478 (N_2478,N_1034,N_1596);
nor U2479 (N_2479,N_1858,N_1944);
nor U2480 (N_2480,N_1553,N_1767);
or U2481 (N_2481,N_1581,N_1358);
nand U2482 (N_2482,N_1350,N_1411);
nand U2483 (N_2483,N_1114,N_1745);
xnor U2484 (N_2484,N_1326,N_1734);
and U2485 (N_2485,N_1662,N_1226);
xor U2486 (N_2486,N_1643,N_1275);
nor U2487 (N_2487,N_1613,N_1865);
nand U2488 (N_2488,N_1725,N_1373);
nand U2489 (N_2489,N_1200,N_1976);
xor U2490 (N_2490,N_1490,N_1735);
nand U2491 (N_2491,N_1797,N_1909);
xnor U2492 (N_2492,N_1984,N_1710);
nand U2493 (N_2493,N_1615,N_1692);
and U2494 (N_2494,N_1706,N_1134);
nand U2495 (N_2495,N_1900,N_1848);
or U2496 (N_2496,N_1416,N_1481);
or U2497 (N_2497,N_1972,N_1709);
or U2498 (N_2498,N_1309,N_1079);
xnor U2499 (N_2499,N_1586,N_1005);
xnor U2500 (N_2500,N_1072,N_1123);
or U2501 (N_2501,N_1511,N_1306);
or U2502 (N_2502,N_1283,N_1929);
nor U2503 (N_2503,N_1394,N_1666);
or U2504 (N_2504,N_1922,N_1295);
and U2505 (N_2505,N_1345,N_1128);
or U2506 (N_2506,N_1966,N_1991);
nand U2507 (N_2507,N_1466,N_1101);
and U2508 (N_2508,N_1280,N_1156);
and U2509 (N_2509,N_1187,N_1049);
nor U2510 (N_2510,N_1542,N_1396);
or U2511 (N_2511,N_1316,N_1877);
nor U2512 (N_2512,N_1719,N_1573);
or U2513 (N_2513,N_1408,N_1226);
and U2514 (N_2514,N_1004,N_1862);
nor U2515 (N_2515,N_1178,N_1336);
nor U2516 (N_2516,N_1719,N_1011);
nand U2517 (N_2517,N_1215,N_1581);
and U2518 (N_2518,N_1049,N_1048);
and U2519 (N_2519,N_1410,N_1863);
and U2520 (N_2520,N_1975,N_1566);
and U2521 (N_2521,N_1176,N_1491);
nor U2522 (N_2522,N_1933,N_1594);
and U2523 (N_2523,N_1906,N_1450);
or U2524 (N_2524,N_1664,N_1073);
or U2525 (N_2525,N_1660,N_1944);
nand U2526 (N_2526,N_1854,N_1624);
or U2527 (N_2527,N_1452,N_1186);
and U2528 (N_2528,N_1944,N_1430);
nand U2529 (N_2529,N_1888,N_1310);
nand U2530 (N_2530,N_1935,N_1402);
and U2531 (N_2531,N_1783,N_1423);
nor U2532 (N_2532,N_1893,N_1988);
or U2533 (N_2533,N_1149,N_1067);
and U2534 (N_2534,N_1088,N_1875);
or U2535 (N_2535,N_1565,N_1542);
nor U2536 (N_2536,N_1181,N_1132);
or U2537 (N_2537,N_1442,N_1620);
or U2538 (N_2538,N_1388,N_1791);
nand U2539 (N_2539,N_1743,N_1564);
nor U2540 (N_2540,N_1732,N_1805);
nand U2541 (N_2541,N_1618,N_1266);
nor U2542 (N_2542,N_1977,N_1167);
xnor U2543 (N_2543,N_1600,N_1255);
nand U2544 (N_2544,N_1122,N_1400);
and U2545 (N_2545,N_1536,N_1425);
nand U2546 (N_2546,N_1601,N_1842);
nor U2547 (N_2547,N_1603,N_1151);
xor U2548 (N_2548,N_1123,N_1639);
or U2549 (N_2549,N_1109,N_1117);
nor U2550 (N_2550,N_1514,N_1712);
and U2551 (N_2551,N_1814,N_1074);
and U2552 (N_2552,N_1828,N_1231);
nor U2553 (N_2553,N_1614,N_1544);
and U2554 (N_2554,N_1082,N_1030);
or U2555 (N_2555,N_1165,N_1321);
nor U2556 (N_2556,N_1972,N_1017);
or U2557 (N_2557,N_1255,N_1421);
nor U2558 (N_2558,N_1237,N_1221);
nand U2559 (N_2559,N_1208,N_1673);
nand U2560 (N_2560,N_1874,N_1781);
and U2561 (N_2561,N_1203,N_1501);
and U2562 (N_2562,N_1078,N_1919);
nor U2563 (N_2563,N_1451,N_1955);
nor U2564 (N_2564,N_1548,N_1961);
and U2565 (N_2565,N_1818,N_1281);
nor U2566 (N_2566,N_1162,N_1785);
or U2567 (N_2567,N_1780,N_1878);
nand U2568 (N_2568,N_1370,N_1845);
or U2569 (N_2569,N_1369,N_1724);
nor U2570 (N_2570,N_1453,N_1673);
and U2571 (N_2571,N_1019,N_1942);
nor U2572 (N_2572,N_1093,N_1632);
nand U2573 (N_2573,N_1416,N_1975);
or U2574 (N_2574,N_1561,N_1134);
nor U2575 (N_2575,N_1681,N_1934);
or U2576 (N_2576,N_1290,N_1305);
and U2577 (N_2577,N_1645,N_1596);
and U2578 (N_2578,N_1102,N_1940);
and U2579 (N_2579,N_1361,N_1139);
and U2580 (N_2580,N_1525,N_1927);
nor U2581 (N_2581,N_1192,N_1392);
and U2582 (N_2582,N_1419,N_1067);
and U2583 (N_2583,N_1999,N_1623);
nor U2584 (N_2584,N_1056,N_1665);
or U2585 (N_2585,N_1103,N_1997);
and U2586 (N_2586,N_1775,N_1891);
or U2587 (N_2587,N_1289,N_1340);
and U2588 (N_2588,N_1423,N_1724);
and U2589 (N_2589,N_1172,N_1500);
and U2590 (N_2590,N_1113,N_1383);
and U2591 (N_2591,N_1906,N_1771);
or U2592 (N_2592,N_1775,N_1607);
nand U2593 (N_2593,N_1371,N_1954);
or U2594 (N_2594,N_1553,N_1030);
xnor U2595 (N_2595,N_1334,N_1804);
and U2596 (N_2596,N_1617,N_1757);
or U2597 (N_2597,N_1129,N_1424);
nor U2598 (N_2598,N_1849,N_1023);
nor U2599 (N_2599,N_1705,N_1613);
and U2600 (N_2600,N_1540,N_1652);
and U2601 (N_2601,N_1278,N_1142);
nand U2602 (N_2602,N_1589,N_1048);
or U2603 (N_2603,N_1805,N_1877);
or U2604 (N_2604,N_1509,N_1728);
or U2605 (N_2605,N_1633,N_1203);
and U2606 (N_2606,N_1762,N_1828);
nand U2607 (N_2607,N_1672,N_1697);
nor U2608 (N_2608,N_1302,N_1466);
and U2609 (N_2609,N_1433,N_1072);
or U2610 (N_2610,N_1272,N_1523);
nor U2611 (N_2611,N_1955,N_1170);
nor U2612 (N_2612,N_1591,N_1499);
xor U2613 (N_2613,N_1079,N_1579);
nor U2614 (N_2614,N_1174,N_1547);
or U2615 (N_2615,N_1865,N_1612);
or U2616 (N_2616,N_1630,N_1794);
nand U2617 (N_2617,N_1244,N_1246);
and U2618 (N_2618,N_1994,N_1537);
or U2619 (N_2619,N_1103,N_1473);
nor U2620 (N_2620,N_1580,N_1643);
and U2621 (N_2621,N_1201,N_1941);
or U2622 (N_2622,N_1832,N_1483);
nand U2623 (N_2623,N_1265,N_1253);
and U2624 (N_2624,N_1321,N_1935);
nor U2625 (N_2625,N_1296,N_1981);
nor U2626 (N_2626,N_1047,N_1169);
or U2627 (N_2627,N_1892,N_1495);
and U2628 (N_2628,N_1640,N_1787);
or U2629 (N_2629,N_1035,N_1789);
and U2630 (N_2630,N_1991,N_1615);
nand U2631 (N_2631,N_1021,N_1871);
or U2632 (N_2632,N_1355,N_1961);
and U2633 (N_2633,N_1525,N_1846);
xnor U2634 (N_2634,N_1964,N_1466);
nand U2635 (N_2635,N_1728,N_1733);
or U2636 (N_2636,N_1620,N_1380);
nor U2637 (N_2637,N_1463,N_1393);
and U2638 (N_2638,N_1919,N_1090);
nor U2639 (N_2639,N_1956,N_1111);
xor U2640 (N_2640,N_1410,N_1620);
nor U2641 (N_2641,N_1393,N_1715);
or U2642 (N_2642,N_1034,N_1682);
or U2643 (N_2643,N_1356,N_1621);
and U2644 (N_2644,N_1783,N_1425);
xnor U2645 (N_2645,N_1693,N_1178);
and U2646 (N_2646,N_1533,N_1622);
and U2647 (N_2647,N_1669,N_1865);
nor U2648 (N_2648,N_1341,N_1027);
or U2649 (N_2649,N_1470,N_1501);
xor U2650 (N_2650,N_1978,N_1695);
or U2651 (N_2651,N_1114,N_1521);
or U2652 (N_2652,N_1030,N_1443);
and U2653 (N_2653,N_1868,N_1755);
nand U2654 (N_2654,N_1861,N_1352);
and U2655 (N_2655,N_1872,N_1871);
nand U2656 (N_2656,N_1672,N_1656);
or U2657 (N_2657,N_1033,N_1058);
or U2658 (N_2658,N_1208,N_1995);
nor U2659 (N_2659,N_1005,N_1617);
and U2660 (N_2660,N_1807,N_1440);
nand U2661 (N_2661,N_1126,N_1435);
nor U2662 (N_2662,N_1830,N_1885);
nand U2663 (N_2663,N_1965,N_1098);
nand U2664 (N_2664,N_1380,N_1348);
and U2665 (N_2665,N_1538,N_1195);
nor U2666 (N_2666,N_1891,N_1522);
and U2667 (N_2667,N_1641,N_1281);
and U2668 (N_2668,N_1787,N_1203);
xnor U2669 (N_2669,N_1894,N_1303);
and U2670 (N_2670,N_1253,N_1156);
nor U2671 (N_2671,N_1016,N_1652);
nor U2672 (N_2672,N_1125,N_1894);
nand U2673 (N_2673,N_1965,N_1477);
or U2674 (N_2674,N_1934,N_1747);
nand U2675 (N_2675,N_1269,N_1539);
and U2676 (N_2676,N_1387,N_1996);
and U2677 (N_2677,N_1723,N_1973);
and U2678 (N_2678,N_1861,N_1225);
nor U2679 (N_2679,N_1100,N_1744);
and U2680 (N_2680,N_1259,N_1046);
nand U2681 (N_2681,N_1405,N_1687);
nand U2682 (N_2682,N_1064,N_1202);
nor U2683 (N_2683,N_1482,N_1388);
and U2684 (N_2684,N_1468,N_1221);
nor U2685 (N_2685,N_1044,N_1478);
xor U2686 (N_2686,N_1376,N_1918);
or U2687 (N_2687,N_1702,N_1118);
nor U2688 (N_2688,N_1289,N_1179);
xnor U2689 (N_2689,N_1722,N_1652);
nor U2690 (N_2690,N_1965,N_1185);
nor U2691 (N_2691,N_1658,N_1676);
or U2692 (N_2692,N_1868,N_1328);
or U2693 (N_2693,N_1950,N_1762);
nand U2694 (N_2694,N_1466,N_1000);
nand U2695 (N_2695,N_1470,N_1529);
nor U2696 (N_2696,N_1930,N_1877);
xor U2697 (N_2697,N_1813,N_1997);
or U2698 (N_2698,N_1432,N_1269);
nand U2699 (N_2699,N_1741,N_1514);
nor U2700 (N_2700,N_1374,N_1109);
nor U2701 (N_2701,N_1168,N_1578);
nand U2702 (N_2702,N_1062,N_1600);
or U2703 (N_2703,N_1262,N_1702);
and U2704 (N_2704,N_1463,N_1450);
nor U2705 (N_2705,N_1753,N_1187);
and U2706 (N_2706,N_1994,N_1247);
nand U2707 (N_2707,N_1653,N_1549);
and U2708 (N_2708,N_1323,N_1992);
nand U2709 (N_2709,N_1134,N_1615);
nand U2710 (N_2710,N_1083,N_1349);
nand U2711 (N_2711,N_1896,N_1617);
or U2712 (N_2712,N_1525,N_1035);
xor U2713 (N_2713,N_1578,N_1824);
or U2714 (N_2714,N_1892,N_1141);
and U2715 (N_2715,N_1711,N_1627);
or U2716 (N_2716,N_1716,N_1123);
nand U2717 (N_2717,N_1676,N_1815);
or U2718 (N_2718,N_1983,N_1102);
and U2719 (N_2719,N_1679,N_1522);
nor U2720 (N_2720,N_1418,N_1384);
or U2721 (N_2721,N_1629,N_1838);
or U2722 (N_2722,N_1402,N_1730);
nor U2723 (N_2723,N_1315,N_1709);
nor U2724 (N_2724,N_1135,N_1255);
nor U2725 (N_2725,N_1410,N_1963);
or U2726 (N_2726,N_1226,N_1689);
xor U2727 (N_2727,N_1696,N_1276);
or U2728 (N_2728,N_1320,N_1590);
or U2729 (N_2729,N_1710,N_1982);
xor U2730 (N_2730,N_1210,N_1849);
xor U2731 (N_2731,N_1371,N_1094);
nor U2732 (N_2732,N_1014,N_1985);
and U2733 (N_2733,N_1031,N_1764);
or U2734 (N_2734,N_1446,N_1384);
nor U2735 (N_2735,N_1005,N_1852);
nor U2736 (N_2736,N_1142,N_1510);
nand U2737 (N_2737,N_1792,N_1744);
or U2738 (N_2738,N_1264,N_1951);
nor U2739 (N_2739,N_1156,N_1482);
or U2740 (N_2740,N_1501,N_1504);
and U2741 (N_2741,N_1602,N_1065);
nand U2742 (N_2742,N_1587,N_1548);
nand U2743 (N_2743,N_1392,N_1945);
nand U2744 (N_2744,N_1615,N_1347);
nand U2745 (N_2745,N_1645,N_1507);
or U2746 (N_2746,N_1249,N_1285);
nor U2747 (N_2747,N_1913,N_1363);
xor U2748 (N_2748,N_1848,N_1672);
and U2749 (N_2749,N_1666,N_1959);
and U2750 (N_2750,N_1223,N_1118);
or U2751 (N_2751,N_1607,N_1126);
and U2752 (N_2752,N_1797,N_1396);
or U2753 (N_2753,N_1247,N_1921);
xor U2754 (N_2754,N_1183,N_1541);
nor U2755 (N_2755,N_1023,N_1298);
and U2756 (N_2756,N_1464,N_1523);
nor U2757 (N_2757,N_1047,N_1944);
and U2758 (N_2758,N_1505,N_1011);
nand U2759 (N_2759,N_1189,N_1757);
and U2760 (N_2760,N_1757,N_1412);
and U2761 (N_2761,N_1995,N_1008);
xnor U2762 (N_2762,N_1791,N_1580);
nand U2763 (N_2763,N_1824,N_1989);
nand U2764 (N_2764,N_1189,N_1067);
nand U2765 (N_2765,N_1358,N_1281);
nand U2766 (N_2766,N_1831,N_1205);
or U2767 (N_2767,N_1296,N_1938);
nand U2768 (N_2768,N_1272,N_1914);
xor U2769 (N_2769,N_1863,N_1090);
nor U2770 (N_2770,N_1143,N_1475);
and U2771 (N_2771,N_1806,N_1792);
and U2772 (N_2772,N_1290,N_1420);
nand U2773 (N_2773,N_1689,N_1554);
or U2774 (N_2774,N_1245,N_1632);
nor U2775 (N_2775,N_1878,N_1402);
nand U2776 (N_2776,N_1865,N_1916);
or U2777 (N_2777,N_1438,N_1745);
and U2778 (N_2778,N_1173,N_1116);
nand U2779 (N_2779,N_1465,N_1851);
nor U2780 (N_2780,N_1759,N_1476);
or U2781 (N_2781,N_1035,N_1111);
or U2782 (N_2782,N_1910,N_1133);
or U2783 (N_2783,N_1164,N_1535);
and U2784 (N_2784,N_1044,N_1253);
xnor U2785 (N_2785,N_1464,N_1888);
or U2786 (N_2786,N_1451,N_1244);
or U2787 (N_2787,N_1553,N_1055);
xnor U2788 (N_2788,N_1372,N_1260);
nand U2789 (N_2789,N_1706,N_1463);
or U2790 (N_2790,N_1783,N_1033);
xor U2791 (N_2791,N_1204,N_1172);
nand U2792 (N_2792,N_1926,N_1148);
nand U2793 (N_2793,N_1895,N_1131);
or U2794 (N_2794,N_1107,N_1287);
or U2795 (N_2795,N_1865,N_1971);
and U2796 (N_2796,N_1633,N_1169);
nand U2797 (N_2797,N_1834,N_1359);
nand U2798 (N_2798,N_1615,N_1403);
and U2799 (N_2799,N_1674,N_1810);
nor U2800 (N_2800,N_1917,N_1707);
xnor U2801 (N_2801,N_1203,N_1596);
and U2802 (N_2802,N_1165,N_1817);
xor U2803 (N_2803,N_1515,N_1063);
nor U2804 (N_2804,N_1955,N_1417);
nand U2805 (N_2805,N_1097,N_1391);
or U2806 (N_2806,N_1242,N_1137);
nor U2807 (N_2807,N_1722,N_1025);
nand U2808 (N_2808,N_1062,N_1671);
nand U2809 (N_2809,N_1874,N_1516);
nand U2810 (N_2810,N_1497,N_1589);
and U2811 (N_2811,N_1570,N_1110);
nor U2812 (N_2812,N_1272,N_1271);
nand U2813 (N_2813,N_1117,N_1783);
xnor U2814 (N_2814,N_1069,N_1607);
nand U2815 (N_2815,N_1523,N_1493);
nor U2816 (N_2816,N_1624,N_1058);
and U2817 (N_2817,N_1334,N_1125);
and U2818 (N_2818,N_1331,N_1911);
and U2819 (N_2819,N_1394,N_1705);
and U2820 (N_2820,N_1145,N_1354);
nor U2821 (N_2821,N_1281,N_1750);
nand U2822 (N_2822,N_1098,N_1900);
xor U2823 (N_2823,N_1743,N_1276);
or U2824 (N_2824,N_1516,N_1015);
or U2825 (N_2825,N_1530,N_1284);
and U2826 (N_2826,N_1665,N_1287);
or U2827 (N_2827,N_1104,N_1139);
nand U2828 (N_2828,N_1738,N_1270);
nand U2829 (N_2829,N_1837,N_1415);
nand U2830 (N_2830,N_1277,N_1033);
or U2831 (N_2831,N_1428,N_1272);
and U2832 (N_2832,N_1813,N_1345);
nor U2833 (N_2833,N_1721,N_1431);
xnor U2834 (N_2834,N_1999,N_1358);
or U2835 (N_2835,N_1794,N_1241);
or U2836 (N_2836,N_1251,N_1831);
nand U2837 (N_2837,N_1292,N_1872);
nand U2838 (N_2838,N_1385,N_1118);
or U2839 (N_2839,N_1564,N_1125);
nor U2840 (N_2840,N_1482,N_1572);
nand U2841 (N_2841,N_1845,N_1047);
and U2842 (N_2842,N_1049,N_1655);
and U2843 (N_2843,N_1629,N_1862);
nor U2844 (N_2844,N_1952,N_1025);
nand U2845 (N_2845,N_1137,N_1527);
and U2846 (N_2846,N_1242,N_1377);
nor U2847 (N_2847,N_1949,N_1365);
or U2848 (N_2848,N_1219,N_1128);
nor U2849 (N_2849,N_1991,N_1861);
and U2850 (N_2850,N_1135,N_1780);
and U2851 (N_2851,N_1163,N_1662);
nand U2852 (N_2852,N_1158,N_1177);
nor U2853 (N_2853,N_1624,N_1129);
xor U2854 (N_2854,N_1520,N_1698);
and U2855 (N_2855,N_1259,N_1101);
xor U2856 (N_2856,N_1076,N_1705);
and U2857 (N_2857,N_1858,N_1723);
nand U2858 (N_2858,N_1898,N_1014);
and U2859 (N_2859,N_1500,N_1480);
nand U2860 (N_2860,N_1022,N_1911);
xnor U2861 (N_2861,N_1080,N_1319);
nand U2862 (N_2862,N_1603,N_1914);
and U2863 (N_2863,N_1183,N_1548);
or U2864 (N_2864,N_1856,N_1481);
nand U2865 (N_2865,N_1271,N_1728);
nand U2866 (N_2866,N_1769,N_1000);
or U2867 (N_2867,N_1789,N_1992);
or U2868 (N_2868,N_1393,N_1531);
or U2869 (N_2869,N_1906,N_1496);
nor U2870 (N_2870,N_1327,N_1651);
nor U2871 (N_2871,N_1194,N_1258);
and U2872 (N_2872,N_1348,N_1638);
xnor U2873 (N_2873,N_1074,N_1085);
and U2874 (N_2874,N_1962,N_1891);
and U2875 (N_2875,N_1000,N_1091);
nand U2876 (N_2876,N_1390,N_1477);
nand U2877 (N_2877,N_1570,N_1423);
nand U2878 (N_2878,N_1511,N_1138);
nand U2879 (N_2879,N_1813,N_1017);
and U2880 (N_2880,N_1787,N_1704);
nand U2881 (N_2881,N_1440,N_1342);
and U2882 (N_2882,N_1732,N_1203);
nand U2883 (N_2883,N_1395,N_1644);
and U2884 (N_2884,N_1310,N_1771);
nor U2885 (N_2885,N_1409,N_1229);
xor U2886 (N_2886,N_1852,N_1256);
nor U2887 (N_2887,N_1968,N_1073);
xor U2888 (N_2888,N_1449,N_1680);
nor U2889 (N_2889,N_1409,N_1960);
and U2890 (N_2890,N_1228,N_1317);
nand U2891 (N_2891,N_1041,N_1815);
or U2892 (N_2892,N_1716,N_1662);
and U2893 (N_2893,N_1711,N_1693);
or U2894 (N_2894,N_1198,N_1471);
nor U2895 (N_2895,N_1218,N_1598);
nor U2896 (N_2896,N_1236,N_1795);
nor U2897 (N_2897,N_1840,N_1395);
nor U2898 (N_2898,N_1510,N_1069);
or U2899 (N_2899,N_1023,N_1376);
and U2900 (N_2900,N_1977,N_1079);
or U2901 (N_2901,N_1195,N_1391);
or U2902 (N_2902,N_1601,N_1419);
or U2903 (N_2903,N_1139,N_1313);
nand U2904 (N_2904,N_1193,N_1359);
nand U2905 (N_2905,N_1430,N_1155);
nand U2906 (N_2906,N_1734,N_1220);
or U2907 (N_2907,N_1580,N_1723);
or U2908 (N_2908,N_1638,N_1697);
and U2909 (N_2909,N_1686,N_1581);
or U2910 (N_2910,N_1422,N_1380);
and U2911 (N_2911,N_1739,N_1404);
or U2912 (N_2912,N_1579,N_1450);
nand U2913 (N_2913,N_1323,N_1577);
or U2914 (N_2914,N_1185,N_1340);
and U2915 (N_2915,N_1450,N_1926);
nand U2916 (N_2916,N_1997,N_1793);
xnor U2917 (N_2917,N_1746,N_1767);
nor U2918 (N_2918,N_1618,N_1505);
nor U2919 (N_2919,N_1164,N_1051);
and U2920 (N_2920,N_1437,N_1200);
xor U2921 (N_2921,N_1575,N_1011);
or U2922 (N_2922,N_1064,N_1357);
nand U2923 (N_2923,N_1955,N_1184);
nor U2924 (N_2924,N_1143,N_1949);
and U2925 (N_2925,N_1129,N_1368);
or U2926 (N_2926,N_1493,N_1492);
or U2927 (N_2927,N_1753,N_1381);
and U2928 (N_2928,N_1682,N_1788);
or U2929 (N_2929,N_1224,N_1477);
and U2930 (N_2930,N_1820,N_1088);
or U2931 (N_2931,N_1373,N_1857);
and U2932 (N_2932,N_1235,N_1788);
and U2933 (N_2933,N_1135,N_1228);
nand U2934 (N_2934,N_1321,N_1009);
and U2935 (N_2935,N_1096,N_1515);
nor U2936 (N_2936,N_1822,N_1623);
or U2937 (N_2937,N_1950,N_1408);
or U2938 (N_2938,N_1269,N_1458);
xor U2939 (N_2939,N_1020,N_1960);
or U2940 (N_2940,N_1921,N_1269);
and U2941 (N_2941,N_1399,N_1435);
and U2942 (N_2942,N_1188,N_1454);
and U2943 (N_2943,N_1517,N_1537);
and U2944 (N_2944,N_1707,N_1839);
or U2945 (N_2945,N_1352,N_1018);
and U2946 (N_2946,N_1657,N_1989);
nor U2947 (N_2947,N_1578,N_1388);
xnor U2948 (N_2948,N_1493,N_1762);
and U2949 (N_2949,N_1345,N_1398);
nand U2950 (N_2950,N_1344,N_1762);
nand U2951 (N_2951,N_1047,N_1093);
nand U2952 (N_2952,N_1975,N_1195);
or U2953 (N_2953,N_1675,N_1228);
xor U2954 (N_2954,N_1203,N_1522);
and U2955 (N_2955,N_1126,N_1874);
or U2956 (N_2956,N_1474,N_1231);
and U2957 (N_2957,N_1952,N_1355);
nand U2958 (N_2958,N_1427,N_1944);
nand U2959 (N_2959,N_1911,N_1044);
nor U2960 (N_2960,N_1979,N_1253);
and U2961 (N_2961,N_1989,N_1028);
nor U2962 (N_2962,N_1534,N_1204);
or U2963 (N_2963,N_1690,N_1994);
nand U2964 (N_2964,N_1577,N_1544);
and U2965 (N_2965,N_1080,N_1591);
nand U2966 (N_2966,N_1301,N_1609);
xnor U2967 (N_2967,N_1012,N_1586);
nand U2968 (N_2968,N_1657,N_1793);
or U2969 (N_2969,N_1408,N_1067);
nor U2970 (N_2970,N_1831,N_1461);
nor U2971 (N_2971,N_1302,N_1796);
and U2972 (N_2972,N_1843,N_1911);
and U2973 (N_2973,N_1164,N_1089);
and U2974 (N_2974,N_1407,N_1100);
or U2975 (N_2975,N_1418,N_1365);
or U2976 (N_2976,N_1777,N_1740);
xnor U2977 (N_2977,N_1843,N_1255);
nor U2978 (N_2978,N_1226,N_1918);
nand U2979 (N_2979,N_1863,N_1907);
nor U2980 (N_2980,N_1995,N_1809);
xor U2981 (N_2981,N_1921,N_1380);
or U2982 (N_2982,N_1073,N_1368);
and U2983 (N_2983,N_1083,N_1126);
nand U2984 (N_2984,N_1716,N_1057);
nand U2985 (N_2985,N_1706,N_1135);
or U2986 (N_2986,N_1697,N_1242);
xor U2987 (N_2987,N_1922,N_1660);
nor U2988 (N_2988,N_1100,N_1422);
nor U2989 (N_2989,N_1680,N_1423);
xnor U2990 (N_2990,N_1663,N_1143);
nor U2991 (N_2991,N_1348,N_1403);
nand U2992 (N_2992,N_1094,N_1145);
xor U2993 (N_2993,N_1172,N_1206);
and U2994 (N_2994,N_1569,N_1021);
nand U2995 (N_2995,N_1534,N_1835);
nor U2996 (N_2996,N_1505,N_1327);
and U2997 (N_2997,N_1343,N_1533);
or U2998 (N_2998,N_1613,N_1739);
and U2999 (N_2999,N_1830,N_1112);
nor U3000 (N_3000,N_2502,N_2771);
or U3001 (N_3001,N_2872,N_2442);
and U3002 (N_3002,N_2334,N_2251);
nor U3003 (N_3003,N_2765,N_2075);
or U3004 (N_3004,N_2932,N_2778);
nand U3005 (N_3005,N_2793,N_2563);
and U3006 (N_3006,N_2378,N_2947);
and U3007 (N_3007,N_2377,N_2272);
nor U3008 (N_3008,N_2191,N_2840);
and U3009 (N_3009,N_2481,N_2930);
nor U3010 (N_3010,N_2753,N_2216);
nor U3011 (N_3011,N_2529,N_2000);
nand U3012 (N_3012,N_2819,N_2827);
xor U3013 (N_3013,N_2496,N_2069);
nand U3014 (N_3014,N_2803,N_2598);
nand U3015 (N_3015,N_2472,N_2056);
or U3016 (N_3016,N_2209,N_2305);
or U3017 (N_3017,N_2583,N_2749);
nor U3018 (N_3018,N_2610,N_2572);
nand U3019 (N_3019,N_2477,N_2602);
nand U3020 (N_3020,N_2278,N_2915);
nand U3021 (N_3021,N_2141,N_2814);
nand U3022 (N_3022,N_2329,N_2314);
and U3023 (N_3023,N_2663,N_2355);
nand U3024 (N_3024,N_2419,N_2726);
nand U3025 (N_3025,N_2405,N_2370);
or U3026 (N_3026,N_2674,N_2298);
and U3027 (N_3027,N_2256,N_2794);
and U3028 (N_3028,N_2660,N_2969);
nor U3029 (N_3029,N_2341,N_2899);
and U3030 (N_3030,N_2345,N_2004);
or U3031 (N_3031,N_2231,N_2770);
nand U3032 (N_3032,N_2903,N_2198);
nand U3033 (N_3033,N_2489,N_2908);
or U3034 (N_3034,N_2934,N_2754);
and U3035 (N_3035,N_2107,N_2296);
xnor U3036 (N_3036,N_2444,N_2025);
and U3037 (N_3037,N_2071,N_2239);
nand U3038 (N_3038,N_2177,N_2768);
nor U3039 (N_3039,N_2459,N_2796);
and U3040 (N_3040,N_2175,N_2153);
xnor U3041 (N_3041,N_2702,N_2810);
or U3042 (N_3042,N_2625,N_2517);
xor U3043 (N_3043,N_2923,N_2109);
and U3044 (N_3044,N_2902,N_2401);
nor U3045 (N_3045,N_2766,N_2804);
and U3046 (N_3046,N_2010,N_2577);
nand U3047 (N_3047,N_2330,N_2809);
nor U3048 (N_3048,N_2890,N_2190);
nand U3049 (N_3049,N_2556,N_2781);
or U3050 (N_3050,N_2669,N_2125);
nor U3051 (N_3051,N_2639,N_2710);
nor U3052 (N_3052,N_2288,N_2657);
and U3053 (N_3053,N_2463,N_2085);
nor U3054 (N_3054,N_2396,N_2937);
nor U3055 (N_3055,N_2093,N_2831);
nand U3056 (N_3056,N_2596,N_2964);
and U3057 (N_3057,N_2178,N_2959);
xor U3058 (N_3058,N_2418,N_2061);
and U3059 (N_3059,N_2464,N_2080);
or U3060 (N_3060,N_2568,N_2211);
xnor U3061 (N_3061,N_2253,N_2842);
and U3062 (N_3062,N_2850,N_2654);
nor U3063 (N_3063,N_2676,N_2587);
and U3064 (N_3064,N_2976,N_2133);
or U3065 (N_3065,N_2407,N_2828);
nand U3066 (N_3066,N_2817,N_2035);
or U3067 (N_3067,N_2928,N_2303);
nand U3068 (N_3068,N_2764,N_2539);
or U3069 (N_3069,N_2650,N_2551);
or U3070 (N_3070,N_2974,N_2328);
or U3071 (N_3071,N_2524,N_2203);
nor U3072 (N_3072,N_2126,N_2946);
xor U3073 (N_3073,N_2611,N_2561);
or U3074 (N_3074,N_2730,N_2222);
nand U3075 (N_3075,N_2255,N_2108);
and U3076 (N_3076,N_2187,N_2698);
nand U3077 (N_3077,N_2549,N_2628);
nor U3078 (N_3078,N_2200,N_2530);
nor U3079 (N_3079,N_2767,N_2362);
nor U3080 (N_3080,N_2824,N_2163);
and U3081 (N_3081,N_2634,N_2901);
and U3082 (N_3082,N_2315,N_2402);
or U3083 (N_3083,N_2366,N_2014);
nor U3084 (N_3084,N_2475,N_2036);
and U3085 (N_3085,N_2875,N_2065);
xnor U3086 (N_3086,N_2413,N_2927);
or U3087 (N_3087,N_2135,N_2834);
and U3088 (N_3088,N_2918,N_2961);
and U3089 (N_3089,N_2049,N_2759);
nand U3090 (N_3090,N_2990,N_2520);
and U3091 (N_3091,N_2054,N_2878);
nand U3092 (N_3092,N_2999,N_2668);
nor U3093 (N_3093,N_2039,N_2981);
nor U3094 (N_3094,N_2467,N_2436);
and U3095 (N_3095,N_2994,N_2034);
or U3096 (N_3096,N_2893,N_2072);
and U3097 (N_3097,N_2632,N_2262);
and U3098 (N_3098,N_2121,N_2829);
and U3099 (N_3099,N_2742,N_2258);
and U3100 (N_3100,N_2204,N_2601);
and U3101 (N_3101,N_2170,N_2326);
nand U3102 (N_3102,N_2704,N_2292);
xnor U3103 (N_3103,N_2168,N_2790);
nor U3104 (N_3104,N_2900,N_2331);
nand U3105 (N_3105,N_2041,N_2214);
nor U3106 (N_3106,N_2060,N_2174);
nand U3107 (N_3107,N_2707,N_2230);
nor U3108 (N_3108,N_2929,N_2183);
or U3109 (N_3109,N_2213,N_2869);
xnor U3110 (N_3110,N_2217,N_2042);
nor U3111 (N_3111,N_2666,N_2095);
or U3112 (N_3112,N_2486,N_2811);
nand U3113 (N_3113,N_2017,N_2207);
nand U3114 (N_3114,N_2219,N_2560);
and U3115 (N_3115,N_2115,N_2942);
nor U3116 (N_3116,N_2692,N_2302);
nand U3117 (N_3117,N_2623,N_2352);
or U3118 (N_3118,N_2067,N_2167);
nand U3119 (N_3119,N_2433,N_2184);
nor U3120 (N_3120,N_2374,N_2734);
nor U3121 (N_3121,N_2452,N_2414);
and U3122 (N_3122,N_2652,N_2408);
nand U3123 (N_3123,N_2088,N_2747);
nand U3124 (N_3124,N_2784,N_2166);
nand U3125 (N_3125,N_2680,N_2671);
nand U3126 (N_3126,N_2388,N_2430);
and U3127 (N_3127,N_2755,N_2252);
nor U3128 (N_3128,N_2830,N_2460);
nor U3129 (N_3129,N_2638,N_2565);
or U3130 (N_3130,N_2741,N_2679);
or U3131 (N_3131,N_2123,N_2287);
nand U3132 (N_3132,N_2357,N_2138);
and U3133 (N_3133,N_2238,N_2157);
or U3134 (N_3134,N_2554,N_2333);
and U3135 (N_3135,N_2971,N_2566);
nand U3136 (N_3136,N_2320,N_2892);
nor U3137 (N_3137,N_2289,N_2818);
or U3138 (N_3138,N_2826,N_2234);
xnor U3139 (N_3139,N_2979,N_2709);
or U3140 (N_3140,N_2488,N_2164);
or U3141 (N_3141,N_2547,N_2143);
or U3142 (N_3142,N_2505,N_2189);
nor U3143 (N_3143,N_2852,N_2494);
nor U3144 (N_3144,N_2142,N_2047);
or U3145 (N_3145,N_2607,N_2694);
xor U3146 (N_3146,N_2672,N_2241);
nor U3147 (N_3147,N_2462,N_2074);
and U3148 (N_3148,N_2291,N_2327);
or U3149 (N_3149,N_2787,N_2227);
nand U3150 (N_3150,N_2756,N_2931);
nor U3151 (N_3151,N_2373,N_2118);
nor U3152 (N_3152,N_2715,N_2732);
or U3153 (N_3153,N_2192,N_2954);
xor U3154 (N_3154,N_2386,N_2906);
or U3155 (N_3155,N_2853,N_2018);
or U3156 (N_3156,N_2030,N_2015);
or U3157 (N_3157,N_2678,N_2380);
xnor U3158 (N_3158,N_2914,N_2473);
or U3159 (N_3159,N_2874,N_2752);
nor U3160 (N_3160,N_2099,N_2703);
nor U3161 (N_3161,N_2132,N_2885);
nand U3162 (N_3162,N_2519,N_2283);
xor U3163 (N_3163,N_2604,N_2526);
and U3164 (N_3164,N_2548,N_2382);
nand U3165 (N_3165,N_2428,N_2960);
nand U3166 (N_3166,N_2581,N_2779);
nor U3167 (N_3167,N_2737,N_2063);
or U3168 (N_3168,N_2655,N_2465);
nor U3169 (N_3169,N_2336,N_2281);
nand U3170 (N_3170,N_2046,N_2735);
or U3171 (N_3171,N_2399,N_2497);
and U3172 (N_3172,N_2245,N_2265);
nand U3173 (N_3173,N_2195,N_2500);
and U3174 (N_3174,N_2171,N_2090);
nor U3175 (N_3175,N_2919,N_2510);
nor U3176 (N_3176,N_2555,N_2338);
or U3177 (N_3177,N_2359,N_2443);
or U3178 (N_3178,N_2651,N_2078);
and U3179 (N_3179,N_2422,N_2471);
and U3180 (N_3180,N_2996,N_2697);
nor U3181 (N_3181,N_2991,N_2938);
or U3182 (N_3182,N_2040,N_2627);
and U3183 (N_3183,N_2120,N_2727);
or U3184 (N_3184,N_2708,N_2441);
and U3185 (N_3185,N_2595,N_2570);
xnor U3186 (N_3186,N_2648,N_2096);
nor U3187 (N_3187,N_2432,N_2884);
or U3188 (N_3188,N_2867,N_2387);
or U3189 (N_3189,N_2206,N_2435);
or U3190 (N_3190,N_2220,N_2434);
nand U3191 (N_3191,N_2368,N_2713);
nand U3192 (N_3192,N_2487,N_2182);
nor U3193 (N_3193,N_2613,N_2316);
nor U3194 (N_3194,N_2169,N_2579);
or U3195 (N_3195,N_2677,N_2102);
or U3196 (N_3196,N_2273,N_2127);
nand U3197 (N_3197,N_2269,N_2323);
nand U3198 (N_3198,N_2662,N_2003);
nor U3199 (N_3199,N_2571,N_2275);
nor U3200 (N_3200,N_2147,N_2146);
and U3201 (N_3201,N_2600,N_2675);
and U3202 (N_3202,N_2729,N_2277);
and U3203 (N_3203,N_2240,N_2215);
nor U3204 (N_3204,N_2640,N_2263);
nor U3205 (N_3205,N_2744,N_2397);
or U3206 (N_3206,N_2006,N_2683);
and U3207 (N_3207,N_2887,N_2509);
and U3208 (N_3208,N_2823,N_2552);
or U3209 (N_3209,N_2599,N_2094);
nor U3210 (N_3210,N_2733,N_2635);
nand U3211 (N_3211,N_2910,N_2031);
nor U3212 (N_3212,N_2606,N_2385);
nor U3213 (N_3213,N_2087,N_2001);
nor U3214 (N_3214,N_2801,N_2986);
and U3215 (N_3215,N_2997,N_2681);
nand U3216 (N_3216,N_2210,N_2957);
nand U3217 (N_3217,N_2700,N_2024);
or U3218 (N_3218,N_2546,N_2337);
and U3219 (N_3219,N_2989,N_2920);
nor U3220 (N_3220,N_2369,N_2822);
and U3221 (N_3221,N_2670,N_2578);
or U3222 (N_3222,N_2409,N_2084);
nand U3223 (N_3223,N_2225,N_2347);
or U3224 (N_3224,N_2848,N_2151);
nand U3225 (N_3225,N_2798,N_2533);
nor U3226 (N_3226,N_2309,N_2975);
xnor U3227 (N_3227,N_2400,N_2592);
and U3228 (N_3228,N_2757,N_2866);
or U3229 (N_3229,N_2792,N_2614);
nand U3230 (N_3230,N_2939,N_2776);
or U3231 (N_3231,N_2699,N_2038);
nand U3232 (N_3232,N_2511,N_2145);
nand U3233 (N_3233,N_2130,N_2479);
nand U3234 (N_3234,N_2545,N_2013);
or U3235 (N_3235,N_2838,N_2806);
and U3236 (N_3236,N_2644,N_2447);
xor U3237 (N_3237,N_2706,N_2558);
nor U3238 (N_3238,N_2835,N_2398);
nand U3239 (N_3239,N_2395,N_2354);
and U3240 (N_3240,N_2940,N_2856);
xnor U3241 (N_3241,N_2955,N_2244);
or U3242 (N_3242,N_2005,N_2112);
and U3243 (N_3243,N_2912,N_2391);
and U3244 (N_3244,N_2980,N_2631);
and U3245 (N_3245,N_2507,N_2188);
and U3246 (N_3246,N_2807,N_2665);
nor U3247 (N_3247,N_2064,N_2228);
xnor U3248 (N_3248,N_2936,N_2185);
or U3249 (N_3249,N_2559,N_2103);
and U3250 (N_3250,N_2772,N_2506);
nand U3251 (N_3251,N_2091,N_2528);
nor U3252 (N_3252,N_2154,N_2297);
and U3253 (N_3253,N_2394,N_2935);
and U3254 (N_3254,N_2081,N_2636);
and U3255 (N_3255,N_2740,N_2023);
nor U3256 (N_3256,N_2448,N_2158);
or U3257 (N_3257,N_2594,N_2712);
and U3258 (N_3258,N_2274,N_2883);
or U3259 (N_3259,N_2523,N_2295);
or U3260 (N_3260,N_2027,N_2349);
nand U3261 (N_3261,N_2172,N_2689);
or U3262 (N_3262,N_2083,N_2128);
or U3263 (N_3263,N_2789,N_2290);
or U3264 (N_3264,N_2008,N_2421);
and U3265 (N_3265,N_2582,N_2514);
nor U3266 (N_3266,N_2492,N_2816);
and U3267 (N_3267,N_2136,N_2243);
nor U3268 (N_3268,N_2716,N_2978);
nand U3269 (N_3269,N_2201,N_2527);
or U3270 (N_3270,N_2116,N_2495);
nand U3271 (N_3271,N_2633,N_2012);
nor U3272 (N_3272,N_2724,N_2160);
nand U3273 (N_3273,N_2403,N_2339);
nand U3274 (N_3274,N_2237,N_2748);
nor U3275 (N_3275,N_2490,N_2114);
nor U3276 (N_3276,N_2846,N_2375);
nand U3277 (N_3277,N_2695,N_2854);
and U3278 (N_3278,N_2659,N_2567);
nand U3279 (N_3279,N_2445,N_2454);
nor U3280 (N_3280,N_2775,N_2294);
and U3281 (N_3281,N_2800,N_2322);
nand U3282 (N_3282,N_2493,N_2865);
nand U3283 (N_3283,N_2420,N_2149);
nand U3284 (N_3284,N_2233,N_2491);
or U3285 (N_3285,N_2905,N_2871);
and U3286 (N_3286,N_2925,N_2832);
xnor U3287 (N_3287,N_2522,N_2100);
or U3288 (N_3288,N_2621,N_2863);
nand U3289 (N_3289,N_2304,N_2310);
nor U3290 (N_3290,N_2332,N_2518);
nand U3291 (N_3291,N_2985,N_2907);
or U3292 (N_3292,N_2022,N_2647);
or U3293 (N_3293,N_2916,N_2603);
nor U3294 (N_3294,N_2426,N_2285);
or U3295 (N_3295,N_2247,N_2293);
xor U3296 (N_3296,N_2485,N_2881);
nand U3297 (N_3297,N_2714,N_2270);
and U3298 (N_3298,N_2193,N_2468);
xor U3299 (N_3299,N_2615,N_2845);
and U3300 (N_3300,N_2470,N_2371);
nor U3301 (N_3301,N_2970,N_2236);
and U3302 (N_3302,N_2791,N_2344);
nor U3303 (N_3303,N_2584,N_2951);
and U3304 (N_3304,N_2007,N_2267);
nand U3305 (N_3305,N_2643,N_2687);
or U3306 (N_3306,N_2739,N_2150);
and U3307 (N_3307,N_2324,N_2098);
nand U3308 (N_3308,N_2622,N_2858);
and U3309 (N_3309,N_2609,N_2686);
and U3310 (N_3310,N_2531,N_2879);
nor U3311 (N_3311,N_2542,N_2097);
or U3312 (N_3312,N_2284,N_2254);
nor U3313 (N_3313,N_2591,N_2082);
or U3314 (N_3314,N_2363,N_2966);
or U3315 (N_3315,N_2086,N_2246);
nor U3316 (N_3316,N_2537,N_2543);
and U3317 (N_3317,N_2588,N_2358);
or U3318 (N_3318,N_2690,N_2286);
or U3319 (N_3319,N_2498,N_2541);
xor U3320 (N_3320,N_2580,N_2043);
xnor U3321 (N_3321,N_2044,N_2788);
and U3322 (N_3322,N_2642,N_2629);
nand U3323 (N_3323,N_2381,N_2540);
nor U3324 (N_3324,N_2573,N_2995);
nand U3325 (N_3325,N_2673,N_2089);
or U3326 (N_3326,N_2924,N_2933);
nand U3327 (N_3327,N_2691,N_2474);
and U3328 (N_3328,N_2410,N_2943);
nand U3329 (N_3329,N_2282,N_2593);
and U3330 (N_3330,N_2965,N_2983);
or U3331 (N_3331,N_2799,N_2992);
and U3332 (N_3332,N_2656,N_2068);
nand U3333 (N_3333,N_2423,N_2346);
or U3334 (N_3334,N_2728,N_2221);
or U3335 (N_3335,N_2194,N_2825);
and U3336 (N_3336,N_2993,N_2562);
nor U3337 (N_3337,N_2684,N_2836);
nand U3338 (N_3338,N_2982,N_2877);
and U3339 (N_3339,N_2364,N_2637);
or U3340 (N_3340,N_2057,N_2967);
xnor U3341 (N_3341,N_2458,N_2750);
nor U3342 (N_3342,N_2389,N_2052);
nand U3343 (N_3343,N_2973,N_2199);
or U3344 (N_3344,N_2351,N_2406);
nor U3345 (N_3345,N_2279,N_2059);
nand U3346 (N_3346,N_2886,N_2751);
or U3347 (N_3347,N_2508,N_2722);
xnor U3348 (N_3348,N_2392,N_2372);
or U3349 (N_3349,N_2079,N_2913);
nand U3350 (N_3350,N_2544,N_2131);
and U3351 (N_3351,N_2589,N_2909);
nand U3352 (N_3352,N_2048,N_2503);
nor U3353 (N_3353,N_2101,N_2760);
and U3354 (N_3354,N_2844,N_2009);
nand U3355 (N_3355,N_2449,N_2894);
or U3356 (N_3356,N_2301,N_2257);
nor U3357 (N_3357,N_2029,N_2813);
xnor U3358 (N_3358,N_2319,N_2944);
nand U3359 (N_3359,N_2889,N_2646);
nand U3360 (N_3360,N_2110,N_2880);
or U3361 (N_3361,N_2941,N_2425);
or U3362 (N_3362,N_2956,N_2605);
nor U3363 (N_3363,N_2019,N_2888);
xnor U3364 (N_3364,N_2271,N_2597);
xnor U3365 (N_3365,N_2053,N_2513);
nand U3366 (N_3366,N_2176,N_2165);
or U3367 (N_3367,N_2313,N_2417);
or U3368 (N_3368,N_2427,N_2111);
and U3369 (N_3369,N_2725,N_2032);
and U3370 (N_3370,N_2312,N_2117);
and U3371 (N_3371,N_2620,N_2782);
nor U3372 (N_3372,N_2062,N_2862);
nand U3373 (N_3373,N_2129,N_2317);
nand U3374 (N_3374,N_2619,N_2917);
and U3375 (N_3375,N_2898,N_2325);
xnor U3376 (N_3376,N_2261,N_2950);
and U3377 (N_3377,N_2224,N_2761);
and U3378 (N_3378,N_2534,N_2229);
nor U3379 (N_3379,N_2055,N_2843);
and U3380 (N_3380,N_2576,N_2876);
or U3381 (N_3381,N_2365,N_2896);
nand U3382 (N_3382,N_2649,N_2104);
or U3383 (N_3383,N_2208,N_2461);
and U3384 (N_3384,N_2259,N_2984);
nor U3385 (N_3385,N_2682,N_2590);
nand U3386 (N_3386,N_2797,N_2066);
nor U3387 (N_3387,N_2242,N_2450);
nor U3388 (N_3388,N_2958,N_2155);
nor U3389 (N_3389,N_2311,N_2482);
nand U3390 (N_3390,N_2466,N_2617);
and U3391 (N_3391,N_2026,N_2348);
or U3392 (N_3392,N_2438,N_2033);
or U3393 (N_3393,N_2945,N_2837);
and U3394 (N_3394,N_2731,N_2028);
nor U3395 (N_3395,N_2140,N_2280);
nand U3396 (N_3396,N_2342,N_2773);
and U3397 (N_3397,N_2181,N_2179);
or U3398 (N_3398,N_2780,N_2411);
nor U3399 (N_3399,N_2306,N_2248);
nor U3400 (N_3400,N_2260,N_2717);
nand U3401 (N_3401,N_2456,N_2499);
or U3402 (N_3402,N_2963,N_2718);
or U3403 (N_3403,N_2353,N_2532);
xnor U3404 (N_3404,N_2076,N_2106);
nor U3405 (N_3405,N_2564,N_2557);
nor U3406 (N_3406,N_2521,N_2777);
nor U3407 (N_3407,N_2383,N_2839);
or U3408 (N_3408,N_2641,N_2988);
nor U3409 (N_3409,N_2808,N_2350);
nor U3410 (N_3410,N_2011,N_2525);
or U3411 (N_3411,N_2439,N_2073);
or U3412 (N_3412,N_2948,N_2833);
nor U3413 (N_3413,N_2020,N_2162);
or U3414 (N_3414,N_2361,N_2569);
nand U3415 (N_3415,N_2685,N_2343);
or U3416 (N_3416,N_2515,N_2002);
or U3417 (N_3417,N_2820,N_2849);
xnor U3418 (N_3418,N_2197,N_2202);
nand U3419 (N_3419,N_2720,N_2148);
nand U3420 (N_3420,N_2021,N_2119);
nand U3421 (N_3421,N_2616,N_2821);
nand U3422 (N_3422,N_2212,N_2701);
and U3423 (N_3423,N_2250,N_2977);
nand U3424 (N_3424,N_2667,N_2962);
or U3425 (N_3425,N_2437,N_2585);
nor U3426 (N_3426,N_2037,N_2318);
nor U3427 (N_3427,N_2746,N_2113);
nor U3428 (N_3428,N_2661,N_2376);
and U3429 (N_3429,N_2904,N_2868);
xnor U3430 (N_3430,N_2390,N_2618);
and U3431 (N_3431,N_2161,N_2841);
nor U3432 (N_3432,N_2105,N_2762);
or U3433 (N_3433,N_2805,N_2736);
or U3434 (N_3434,N_2952,N_2504);
nand U3435 (N_3435,N_2774,N_2308);
or U3436 (N_3436,N_2300,N_2516);
nand U3437 (N_3437,N_2815,N_2612);
or U3438 (N_3438,N_2745,N_2705);
nor U3439 (N_3439,N_2897,N_2608);
or U3440 (N_3440,N_2480,N_2264);
nor U3441 (N_3441,N_2550,N_2658);
nand U3442 (N_3442,N_2186,N_2512);
nor U3443 (N_3443,N_2144,N_2122);
nor U3444 (N_3444,N_2882,N_2645);
nand U3445 (N_3445,N_2783,N_2786);
nor U3446 (N_3446,N_2586,N_2738);
nor U3447 (N_3447,N_2453,N_2972);
and U3448 (N_3448,N_2223,N_2911);
and U3449 (N_3449,N_2152,N_2949);
or U3450 (N_3450,N_2196,N_2077);
or U3451 (N_3451,N_2360,N_2476);
nor U3452 (N_3452,N_2218,N_2501);
or U3453 (N_3453,N_2891,N_2469);
nand U3454 (N_3454,N_2926,N_2873);
nand U3455 (N_3455,N_2384,N_2268);
and U3456 (N_3456,N_2812,N_2173);
and U3457 (N_3457,N_2321,N_2451);
nor U3458 (N_3458,N_2860,N_2058);
nor U3459 (N_3459,N_2536,N_2299);
and U3460 (N_3460,N_2232,N_2226);
or U3461 (N_3461,N_2016,N_2457);
nand U3462 (N_3462,N_2847,N_2484);
xnor U3463 (N_3463,N_2429,N_2688);
nor U3464 (N_3464,N_2859,N_2235);
and U3465 (N_3465,N_2431,N_2743);
nand U3466 (N_3466,N_2412,N_2416);
xor U3467 (N_3467,N_2693,N_2180);
nand U3468 (N_3468,N_2404,N_2723);
nand U3469 (N_3469,N_2156,N_2953);
or U3470 (N_3470,N_2050,N_2092);
or U3471 (N_3471,N_2249,N_2266);
nand U3472 (N_3472,N_2851,N_2205);
nor U3473 (N_3473,N_2630,N_2575);
nand U3474 (N_3474,N_2478,N_2758);
nor U3475 (N_3475,N_2624,N_2998);
xor U3476 (N_3476,N_2070,N_2139);
and U3477 (N_3477,N_2802,N_2137);
nor U3478 (N_3478,N_2857,N_2711);
and U3479 (N_3479,N_2696,N_2626);
nand U3480 (N_3480,N_2455,N_2335);
or U3481 (N_3481,N_2719,N_2446);
or U3482 (N_3482,N_2861,N_2785);
nand U3483 (N_3483,N_2276,N_2968);
nor U3484 (N_3484,N_2367,N_2921);
nor U3485 (N_3485,N_2424,N_2483);
or U3486 (N_3486,N_2415,N_2922);
nand U3487 (N_3487,N_2340,N_2870);
nor U3488 (N_3488,N_2795,N_2987);
and U3489 (N_3489,N_2721,N_2051);
nand U3490 (N_3490,N_2440,N_2356);
or U3491 (N_3491,N_2763,N_2307);
nand U3492 (N_3492,N_2159,N_2538);
nor U3493 (N_3493,N_2393,N_2124);
or U3494 (N_3494,N_2855,N_2134);
and U3495 (N_3495,N_2574,N_2045);
or U3496 (N_3496,N_2769,N_2379);
and U3497 (N_3497,N_2653,N_2895);
or U3498 (N_3498,N_2864,N_2535);
nor U3499 (N_3499,N_2553,N_2664);
xor U3500 (N_3500,N_2083,N_2577);
and U3501 (N_3501,N_2832,N_2428);
or U3502 (N_3502,N_2521,N_2860);
nor U3503 (N_3503,N_2224,N_2949);
nor U3504 (N_3504,N_2270,N_2487);
and U3505 (N_3505,N_2818,N_2232);
nor U3506 (N_3506,N_2425,N_2421);
and U3507 (N_3507,N_2519,N_2831);
or U3508 (N_3508,N_2703,N_2297);
or U3509 (N_3509,N_2744,N_2898);
or U3510 (N_3510,N_2435,N_2770);
nor U3511 (N_3511,N_2744,N_2845);
nor U3512 (N_3512,N_2525,N_2351);
and U3513 (N_3513,N_2952,N_2790);
and U3514 (N_3514,N_2138,N_2590);
and U3515 (N_3515,N_2001,N_2086);
nand U3516 (N_3516,N_2692,N_2935);
nor U3517 (N_3517,N_2559,N_2220);
xnor U3518 (N_3518,N_2519,N_2540);
and U3519 (N_3519,N_2552,N_2471);
or U3520 (N_3520,N_2431,N_2342);
xor U3521 (N_3521,N_2186,N_2440);
nand U3522 (N_3522,N_2875,N_2930);
nand U3523 (N_3523,N_2539,N_2824);
and U3524 (N_3524,N_2427,N_2240);
nand U3525 (N_3525,N_2554,N_2858);
and U3526 (N_3526,N_2709,N_2864);
nor U3527 (N_3527,N_2297,N_2900);
nand U3528 (N_3528,N_2526,N_2987);
nor U3529 (N_3529,N_2211,N_2584);
or U3530 (N_3530,N_2168,N_2305);
nand U3531 (N_3531,N_2761,N_2112);
nor U3532 (N_3532,N_2854,N_2416);
nand U3533 (N_3533,N_2561,N_2316);
and U3534 (N_3534,N_2176,N_2315);
or U3535 (N_3535,N_2408,N_2057);
and U3536 (N_3536,N_2941,N_2569);
nor U3537 (N_3537,N_2317,N_2206);
and U3538 (N_3538,N_2382,N_2386);
or U3539 (N_3539,N_2583,N_2790);
nor U3540 (N_3540,N_2418,N_2092);
xor U3541 (N_3541,N_2863,N_2243);
nor U3542 (N_3542,N_2731,N_2737);
xor U3543 (N_3543,N_2739,N_2217);
nor U3544 (N_3544,N_2612,N_2748);
xor U3545 (N_3545,N_2445,N_2524);
nor U3546 (N_3546,N_2559,N_2335);
xor U3547 (N_3547,N_2938,N_2913);
and U3548 (N_3548,N_2814,N_2090);
nand U3549 (N_3549,N_2488,N_2197);
or U3550 (N_3550,N_2508,N_2556);
and U3551 (N_3551,N_2028,N_2446);
nand U3552 (N_3552,N_2272,N_2006);
nand U3553 (N_3553,N_2225,N_2399);
or U3554 (N_3554,N_2365,N_2911);
or U3555 (N_3555,N_2019,N_2244);
and U3556 (N_3556,N_2746,N_2415);
nand U3557 (N_3557,N_2678,N_2114);
or U3558 (N_3558,N_2432,N_2440);
and U3559 (N_3559,N_2194,N_2282);
or U3560 (N_3560,N_2790,N_2493);
nand U3561 (N_3561,N_2515,N_2510);
and U3562 (N_3562,N_2819,N_2947);
xor U3563 (N_3563,N_2175,N_2184);
nor U3564 (N_3564,N_2878,N_2525);
nand U3565 (N_3565,N_2961,N_2602);
nor U3566 (N_3566,N_2718,N_2427);
xor U3567 (N_3567,N_2558,N_2267);
nand U3568 (N_3568,N_2988,N_2535);
or U3569 (N_3569,N_2543,N_2328);
nor U3570 (N_3570,N_2013,N_2656);
nor U3571 (N_3571,N_2353,N_2158);
or U3572 (N_3572,N_2014,N_2050);
nor U3573 (N_3573,N_2496,N_2678);
or U3574 (N_3574,N_2821,N_2859);
or U3575 (N_3575,N_2574,N_2066);
nor U3576 (N_3576,N_2376,N_2701);
or U3577 (N_3577,N_2837,N_2465);
and U3578 (N_3578,N_2758,N_2955);
nand U3579 (N_3579,N_2773,N_2144);
and U3580 (N_3580,N_2774,N_2013);
xor U3581 (N_3581,N_2242,N_2848);
xor U3582 (N_3582,N_2712,N_2097);
and U3583 (N_3583,N_2860,N_2270);
xnor U3584 (N_3584,N_2117,N_2617);
and U3585 (N_3585,N_2864,N_2404);
and U3586 (N_3586,N_2839,N_2586);
nor U3587 (N_3587,N_2417,N_2307);
or U3588 (N_3588,N_2633,N_2507);
or U3589 (N_3589,N_2325,N_2021);
or U3590 (N_3590,N_2035,N_2020);
and U3591 (N_3591,N_2738,N_2864);
xor U3592 (N_3592,N_2175,N_2955);
and U3593 (N_3593,N_2199,N_2266);
nand U3594 (N_3594,N_2292,N_2230);
xor U3595 (N_3595,N_2423,N_2719);
or U3596 (N_3596,N_2410,N_2105);
nor U3597 (N_3597,N_2639,N_2915);
and U3598 (N_3598,N_2677,N_2950);
and U3599 (N_3599,N_2081,N_2473);
and U3600 (N_3600,N_2314,N_2301);
and U3601 (N_3601,N_2482,N_2276);
nand U3602 (N_3602,N_2431,N_2467);
xor U3603 (N_3603,N_2033,N_2371);
nand U3604 (N_3604,N_2356,N_2927);
or U3605 (N_3605,N_2283,N_2234);
nor U3606 (N_3606,N_2467,N_2029);
or U3607 (N_3607,N_2460,N_2740);
and U3608 (N_3608,N_2524,N_2519);
and U3609 (N_3609,N_2982,N_2351);
and U3610 (N_3610,N_2014,N_2949);
or U3611 (N_3611,N_2978,N_2739);
nand U3612 (N_3612,N_2609,N_2617);
or U3613 (N_3613,N_2642,N_2830);
and U3614 (N_3614,N_2258,N_2468);
nand U3615 (N_3615,N_2949,N_2340);
or U3616 (N_3616,N_2472,N_2359);
nand U3617 (N_3617,N_2935,N_2711);
nand U3618 (N_3618,N_2420,N_2213);
or U3619 (N_3619,N_2346,N_2721);
or U3620 (N_3620,N_2642,N_2884);
nor U3621 (N_3621,N_2056,N_2780);
nor U3622 (N_3622,N_2140,N_2901);
or U3623 (N_3623,N_2445,N_2851);
or U3624 (N_3624,N_2886,N_2020);
xor U3625 (N_3625,N_2049,N_2521);
nor U3626 (N_3626,N_2125,N_2373);
nand U3627 (N_3627,N_2538,N_2613);
or U3628 (N_3628,N_2327,N_2637);
and U3629 (N_3629,N_2725,N_2752);
nor U3630 (N_3630,N_2890,N_2775);
nor U3631 (N_3631,N_2103,N_2283);
or U3632 (N_3632,N_2059,N_2780);
and U3633 (N_3633,N_2957,N_2709);
or U3634 (N_3634,N_2985,N_2300);
nor U3635 (N_3635,N_2996,N_2393);
nor U3636 (N_3636,N_2366,N_2234);
nand U3637 (N_3637,N_2536,N_2649);
xnor U3638 (N_3638,N_2656,N_2435);
xor U3639 (N_3639,N_2265,N_2759);
nand U3640 (N_3640,N_2624,N_2691);
nor U3641 (N_3641,N_2134,N_2199);
and U3642 (N_3642,N_2355,N_2213);
or U3643 (N_3643,N_2698,N_2941);
and U3644 (N_3644,N_2343,N_2185);
xnor U3645 (N_3645,N_2879,N_2487);
or U3646 (N_3646,N_2918,N_2842);
nor U3647 (N_3647,N_2156,N_2741);
and U3648 (N_3648,N_2682,N_2400);
or U3649 (N_3649,N_2699,N_2712);
or U3650 (N_3650,N_2099,N_2121);
nand U3651 (N_3651,N_2504,N_2136);
nand U3652 (N_3652,N_2839,N_2294);
or U3653 (N_3653,N_2344,N_2524);
and U3654 (N_3654,N_2024,N_2976);
and U3655 (N_3655,N_2837,N_2487);
and U3656 (N_3656,N_2968,N_2847);
nand U3657 (N_3657,N_2295,N_2268);
and U3658 (N_3658,N_2413,N_2209);
or U3659 (N_3659,N_2290,N_2589);
and U3660 (N_3660,N_2901,N_2489);
nand U3661 (N_3661,N_2618,N_2945);
nand U3662 (N_3662,N_2787,N_2934);
and U3663 (N_3663,N_2545,N_2941);
or U3664 (N_3664,N_2290,N_2214);
nor U3665 (N_3665,N_2473,N_2957);
nor U3666 (N_3666,N_2643,N_2321);
xor U3667 (N_3667,N_2926,N_2024);
or U3668 (N_3668,N_2809,N_2061);
or U3669 (N_3669,N_2996,N_2030);
xor U3670 (N_3670,N_2634,N_2703);
and U3671 (N_3671,N_2030,N_2572);
and U3672 (N_3672,N_2353,N_2521);
and U3673 (N_3673,N_2063,N_2013);
nor U3674 (N_3674,N_2248,N_2789);
or U3675 (N_3675,N_2681,N_2353);
and U3676 (N_3676,N_2196,N_2161);
or U3677 (N_3677,N_2309,N_2476);
nor U3678 (N_3678,N_2604,N_2140);
nand U3679 (N_3679,N_2392,N_2627);
and U3680 (N_3680,N_2640,N_2477);
nand U3681 (N_3681,N_2822,N_2530);
and U3682 (N_3682,N_2202,N_2941);
and U3683 (N_3683,N_2848,N_2050);
nand U3684 (N_3684,N_2466,N_2519);
xor U3685 (N_3685,N_2607,N_2144);
nand U3686 (N_3686,N_2114,N_2272);
nand U3687 (N_3687,N_2073,N_2111);
xor U3688 (N_3688,N_2912,N_2144);
nand U3689 (N_3689,N_2824,N_2745);
xor U3690 (N_3690,N_2280,N_2007);
nand U3691 (N_3691,N_2553,N_2460);
or U3692 (N_3692,N_2623,N_2290);
and U3693 (N_3693,N_2325,N_2396);
and U3694 (N_3694,N_2120,N_2597);
or U3695 (N_3695,N_2423,N_2122);
and U3696 (N_3696,N_2312,N_2233);
and U3697 (N_3697,N_2142,N_2538);
nand U3698 (N_3698,N_2048,N_2852);
nor U3699 (N_3699,N_2863,N_2964);
nand U3700 (N_3700,N_2364,N_2046);
nor U3701 (N_3701,N_2056,N_2202);
nor U3702 (N_3702,N_2373,N_2121);
nand U3703 (N_3703,N_2668,N_2517);
or U3704 (N_3704,N_2556,N_2672);
or U3705 (N_3705,N_2787,N_2026);
nor U3706 (N_3706,N_2252,N_2775);
or U3707 (N_3707,N_2793,N_2037);
xnor U3708 (N_3708,N_2314,N_2707);
nor U3709 (N_3709,N_2320,N_2116);
nor U3710 (N_3710,N_2193,N_2361);
and U3711 (N_3711,N_2892,N_2769);
nor U3712 (N_3712,N_2088,N_2594);
or U3713 (N_3713,N_2053,N_2322);
or U3714 (N_3714,N_2017,N_2427);
nand U3715 (N_3715,N_2129,N_2770);
or U3716 (N_3716,N_2688,N_2264);
nand U3717 (N_3717,N_2686,N_2383);
xor U3718 (N_3718,N_2743,N_2645);
and U3719 (N_3719,N_2920,N_2380);
or U3720 (N_3720,N_2023,N_2955);
or U3721 (N_3721,N_2377,N_2743);
nand U3722 (N_3722,N_2796,N_2096);
and U3723 (N_3723,N_2121,N_2042);
xor U3724 (N_3724,N_2455,N_2860);
nand U3725 (N_3725,N_2637,N_2257);
nor U3726 (N_3726,N_2541,N_2301);
nor U3727 (N_3727,N_2385,N_2820);
and U3728 (N_3728,N_2169,N_2810);
nand U3729 (N_3729,N_2866,N_2244);
and U3730 (N_3730,N_2965,N_2005);
nor U3731 (N_3731,N_2150,N_2522);
nand U3732 (N_3732,N_2037,N_2946);
nand U3733 (N_3733,N_2422,N_2900);
or U3734 (N_3734,N_2381,N_2224);
nand U3735 (N_3735,N_2097,N_2638);
nand U3736 (N_3736,N_2665,N_2049);
nor U3737 (N_3737,N_2334,N_2327);
nor U3738 (N_3738,N_2780,N_2130);
and U3739 (N_3739,N_2948,N_2194);
nand U3740 (N_3740,N_2627,N_2331);
nand U3741 (N_3741,N_2594,N_2470);
or U3742 (N_3742,N_2063,N_2806);
nor U3743 (N_3743,N_2827,N_2977);
nand U3744 (N_3744,N_2427,N_2433);
nand U3745 (N_3745,N_2276,N_2229);
or U3746 (N_3746,N_2838,N_2361);
nor U3747 (N_3747,N_2051,N_2071);
and U3748 (N_3748,N_2875,N_2255);
nand U3749 (N_3749,N_2499,N_2251);
or U3750 (N_3750,N_2516,N_2801);
nor U3751 (N_3751,N_2920,N_2909);
nand U3752 (N_3752,N_2938,N_2648);
nand U3753 (N_3753,N_2676,N_2483);
and U3754 (N_3754,N_2396,N_2371);
nor U3755 (N_3755,N_2409,N_2103);
or U3756 (N_3756,N_2304,N_2214);
or U3757 (N_3757,N_2469,N_2988);
nand U3758 (N_3758,N_2183,N_2559);
or U3759 (N_3759,N_2208,N_2893);
or U3760 (N_3760,N_2700,N_2582);
nor U3761 (N_3761,N_2204,N_2983);
or U3762 (N_3762,N_2035,N_2894);
nor U3763 (N_3763,N_2713,N_2060);
nand U3764 (N_3764,N_2788,N_2471);
nand U3765 (N_3765,N_2881,N_2617);
nor U3766 (N_3766,N_2792,N_2118);
nand U3767 (N_3767,N_2949,N_2593);
or U3768 (N_3768,N_2392,N_2279);
and U3769 (N_3769,N_2256,N_2537);
nand U3770 (N_3770,N_2821,N_2688);
nor U3771 (N_3771,N_2907,N_2259);
nand U3772 (N_3772,N_2503,N_2713);
nor U3773 (N_3773,N_2134,N_2007);
or U3774 (N_3774,N_2418,N_2017);
and U3775 (N_3775,N_2131,N_2640);
and U3776 (N_3776,N_2020,N_2328);
nor U3777 (N_3777,N_2980,N_2261);
nand U3778 (N_3778,N_2569,N_2592);
or U3779 (N_3779,N_2169,N_2414);
or U3780 (N_3780,N_2444,N_2046);
nor U3781 (N_3781,N_2109,N_2512);
nor U3782 (N_3782,N_2966,N_2970);
and U3783 (N_3783,N_2712,N_2602);
or U3784 (N_3784,N_2672,N_2435);
xor U3785 (N_3785,N_2145,N_2220);
or U3786 (N_3786,N_2928,N_2675);
nor U3787 (N_3787,N_2790,N_2002);
and U3788 (N_3788,N_2498,N_2332);
nand U3789 (N_3789,N_2001,N_2529);
or U3790 (N_3790,N_2534,N_2073);
nand U3791 (N_3791,N_2151,N_2731);
nand U3792 (N_3792,N_2182,N_2459);
xor U3793 (N_3793,N_2031,N_2673);
xor U3794 (N_3794,N_2080,N_2114);
xnor U3795 (N_3795,N_2141,N_2591);
nor U3796 (N_3796,N_2440,N_2674);
nor U3797 (N_3797,N_2847,N_2975);
and U3798 (N_3798,N_2437,N_2921);
xor U3799 (N_3799,N_2674,N_2150);
and U3800 (N_3800,N_2576,N_2681);
nand U3801 (N_3801,N_2721,N_2840);
or U3802 (N_3802,N_2761,N_2318);
xor U3803 (N_3803,N_2946,N_2123);
nor U3804 (N_3804,N_2842,N_2609);
or U3805 (N_3805,N_2120,N_2355);
or U3806 (N_3806,N_2939,N_2086);
nand U3807 (N_3807,N_2560,N_2688);
nand U3808 (N_3808,N_2722,N_2368);
and U3809 (N_3809,N_2071,N_2404);
nand U3810 (N_3810,N_2835,N_2159);
xor U3811 (N_3811,N_2631,N_2927);
nand U3812 (N_3812,N_2690,N_2932);
nor U3813 (N_3813,N_2974,N_2644);
nand U3814 (N_3814,N_2046,N_2412);
or U3815 (N_3815,N_2106,N_2775);
nand U3816 (N_3816,N_2822,N_2771);
or U3817 (N_3817,N_2502,N_2895);
xnor U3818 (N_3818,N_2728,N_2928);
nand U3819 (N_3819,N_2033,N_2568);
nand U3820 (N_3820,N_2505,N_2403);
and U3821 (N_3821,N_2750,N_2606);
nand U3822 (N_3822,N_2940,N_2725);
nand U3823 (N_3823,N_2251,N_2453);
nor U3824 (N_3824,N_2722,N_2976);
and U3825 (N_3825,N_2113,N_2450);
or U3826 (N_3826,N_2971,N_2747);
nor U3827 (N_3827,N_2117,N_2556);
and U3828 (N_3828,N_2596,N_2366);
xnor U3829 (N_3829,N_2999,N_2747);
and U3830 (N_3830,N_2253,N_2114);
nand U3831 (N_3831,N_2987,N_2010);
nand U3832 (N_3832,N_2463,N_2500);
and U3833 (N_3833,N_2516,N_2946);
and U3834 (N_3834,N_2642,N_2783);
nand U3835 (N_3835,N_2796,N_2493);
nand U3836 (N_3836,N_2977,N_2226);
nand U3837 (N_3837,N_2020,N_2897);
and U3838 (N_3838,N_2298,N_2194);
nand U3839 (N_3839,N_2111,N_2563);
nand U3840 (N_3840,N_2492,N_2295);
xnor U3841 (N_3841,N_2653,N_2677);
nor U3842 (N_3842,N_2307,N_2699);
nor U3843 (N_3843,N_2496,N_2271);
xnor U3844 (N_3844,N_2849,N_2634);
or U3845 (N_3845,N_2761,N_2740);
or U3846 (N_3846,N_2471,N_2815);
and U3847 (N_3847,N_2496,N_2650);
and U3848 (N_3848,N_2155,N_2144);
nand U3849 (N_3849,N_2067,N_2358);
xnor U3850 (N_3850,N_2092,N_2822);
or U3851 (N_3851,N_2075,N_2452);
or U3852 (N_3852,N_2348,N_2914);
or U3853 (N_3853,N_2899,N_2279);
or U3854 (N_3854,N_2561,N_2764);
and U3855 (N_3855,N_2486,N_2397);
nand U3856 (N_3856,N_2348,N_2511);
nor U3857 (N_3857,N_2166,N_2972);
xnor U3858 (N_3858,N_2136,N_2803);
nand U3859 (N_3859,N_2534,N_2474);
nand U3860 (N_3860,N_2876,N_2012);
and U3861 (N_3861,N_2858,N_2507);
or U3862 (N_3862,N_2367,N_2049);
nor U3863 (N_3863,N_2122,N_2748);
or U3864 (N_3864,N_2841,N_2641);
or U3865 (N_3865,N_2571,N_2071);
or U3866 (N_3866,N_2517,N_2847);
nand U3867 (N_3867,N_2691,N_2412);
nor U3868 (N_3868,N_2088,N_2742);
nor U3869 (N_3869,N_2668,N_2131);
or U3870 (N_3870,N_2794,N_2588);
and U3871 (N_3871,N_2610,N_2248);
or U3872 (N_3872,N_2592,N_2660);
nor U3873 (N_3873,N_2967,N_2804);
and U3874 (N_3874,N_2376,N_2578);
xor U3875 (N_3875,N_2617,N_2296);
nor U3876 (N_3876,N_2744,N_2958);
or U3877 (N_3877,N_2761,N_2517);
xor U3878 (N_3878,N_2961,N_2356);
nor U3879 (N_3879,N_2166,N_2745);
or U3880 (N_3880,N_2086,N_2030);
and U3881 (N_3881,N_2667,N_2779);
nor U3882 (N_3882,N_2012,N_2052);
or U3883 (N_3883,N_2579,N_2844);
or U3884 (N_3884,N_2178,N_2003);
nor U3885 (N_3885,N_2927,N_2573);
nand U3886 (N_3886,N_2293,N_2900);
nand U3887 (N_3887,N_2041,N_2614);
or U3888 (N_3888,N_2833,N_2315);
and U3889 (N_3889,N_2152,N_2530);
nor U3890 (N_3890,N_2307,N_2695);
nand U3891 (N_3891,N_2114,N_2510);
nor U3892 (N_3892,N_2367,N_2968);
nor U3893 (N_3893,N_2601,N_2786);
xnor U3894 (N_3894,N_2407,N_2404);
nor U3895 (N_3895,N_2229,N_2816);
xnor U3896 (N_3896,N_2537,N_2051);
xor U3897 (N_3897,N_2566,N_2288);
or U3898 (N_3898,N_2543,N_2428);
or U3899 (N_3899,N_2312,N_2849);
or U3900 (N_3900,N_2097,N_2395);
nor U3901 (N_3901,N_2524,N_2735);
nor U3902 (N_3902,N_2104,N_2245);
or U3903 (N_3903,N_2627,N_2991);
and U3904 (N_3904,N_2807,N_2632);
and U3905 (N_3905,N_2262,N_2272);
or U3906 (N_3906,N_2851,N_2932);
xnor U3907 (N_3907,N_2633,N_2795);
and U3908 (N_3908,N_2453,N_2078);
nor U3909 (N_3909,N_2731,N_2383);
or U3910 (N_3910,N_2743,N_2980);
nand U3911 (N_3911,N_2191,N_2904);
or U3912 (N_3912,N_2831,N_2784);
or U3913 (N_3913,N_2276,N_2628);
nor U3914 (N_3914,N_2629,N_2592);
nand U3915 (N_3915,N_2225,N_2901);
or U3916 (N_3916,N_2909,N_2327);
xnor U3917 (N_3917,N_2289,N_2865);
nand U3918 (N_3918,N_2450,N_2709);
nor U3919 (N_3919,N_2953,N_2490);
or U3920 (N_3920,N_2301,N_2618);
nand U3921 (N_3921,N_2364,N_2835);
nand U3922 (N_3922,N_2945,N_2925);
nand U3923 (N_3923,N_2100,N_2226);
xor U3924 (N_3924,N_2836,N_2301);
and U3925 (N_3925,N_2982,N_2794);
nor U3926 (N_3926,N_2311,N_2879);
nor U3927 (N_3927,N_2386,N_2652);
and U3928 (N_3928,N_2876,N_2292);
nand U3929 (N_3929,N_2723,N_2468);
and U3930 (N_3930,N_2364,N_2315);
or U3931 (N_3931,N_2954,N_2217);
and U3932 (N_3932,N_2971,N_2878);
nand U3933 (N_3933,N_2111,N_2609);
and U3934 (N_3934,N_2532,N_2869);
xnor U3935 (N_3935,N_2343,N_2219);
nand U3936 (N_3936,N_2134,N_2786);
nor U3937 (N_3937,N_2113,N_2216);
or U3938 (N_3938,N_2003,N_2791);
nor U3939 (N_3939,N_2075,N_2644);
or U3940 (N_3940,N_2024,N_2705);
nor U3941 (N_3941,N_2704,N_2177);
nand U3942 (N_3942,N_2116,N_2828);
nor U3943 (N_3943,N_2730,N_2215);
nand U3944 (N_3944,N_2170,N_2499);
and U3945 (N_3945,N_2344,N_2620);
nand U3946 (N_3946,N_2310,N_2997);
and U3947 (N_3947,N_2483,N_2191);
nor U3948 (N_3948,N_2078,N_2950);
or U3949 (N_3949,N_2899,N_2978);
nand U3950 (N_3950,N_2306,N_2404);
xor U3951 (N_3951,N_2531,N_2456);
nor U3952 (N_3952,N_2174,N_2742);
or U3953 (N_3953,N_2544,N_2726);
nand U3954 (N_3954,N_2765,N_2383);
and U3955 (N_3955,N_2018,N_2214);
nand U3956 (N_3956,N_2357,N_2812);
nor U3957 (N_3957,N_2519,N_2038);
and U3958 (N_3958,N_2307,N_2984);
nand U3959 (N_3959,N_2782,N_2276);
or U3960 (N_3960,N_2906,N_2787);
or U3961 (N_3961,N_2052,N_2816);
nand U3962 (N_3962,N_2608,N_2814);
nand U3963 (N_3963,N_2398,N_2797);
nand U3964 (N_3964,N_2624,N_2144);
nand U3965 (N_3965,N_2991,N_2871);
nand U3966 (N_3966,N_2195,N_2389);
xnor U3967 (N_3967,N_2494,N_2133);
nor U3968 (N_3968,N_2740,N_2415);
nor U3969 (N_3969,N_2768,N_2319);
xnor U3970 (N_3970,N_2544,N_2123);
nor U3971 (N_3971,N_2861,N_2322);
nor U3972 (N_3972,N_2533,N_2032);
nand U3973 (N_3973,N_2649,N_2396);
or U3974 (N_3974,N_2318,N_2381);
or U3975 (N_3975,N_2609,N_2025);
xnor U3976 (N_3976,N_2781,N_2960);
nor U3977 (N_3977,N_2578,N_2149);
and U3978 (N_3978,N_2699,N_2286);
xnor U3979 (N_3979,N_2021,N_2314);
and U3980 (N_3980,N_2119,N_2763);
or U3981 (N_3981,N_2079,N_2290);
and U3982 (N_3982,N_2773,N_2108);
and U3983 (N_3983,N_2231,N_2990);
or U3984 (N_3984,N_2059,N_2050);
nand U3985 (N_3985,N_2161,N_2513);
xnor U3986 (N_3986,N_2533,N_2212);
or U3987 (N_3987,N_2601,N_2450);
nor U3988 (N_3988,N_2569,N_2909);
nor U3989 (N_3989,N_2063,N_2169);
nand U3990 (N_3990,N_2919,N_2731);
or U3991 (N_3991,N_2985,N_2084);
nor U3992 (N_3992,N_2829,N_2975);
nor U3993 (N_3993,N_2685,N_2194);
or U3994 (N_3994,N_2700,N_2435);
and U3995 (N_3995,N_2356,N_2286);
and U3996 (N_3996,N_2420,N_2939);
or U3997 (N_3997,N_2727,N_2870);
or U3998 (N_3998,N_2019,N_2202);
nand U3999 (N_3999,N_2669,N_2872);
or U4000 (N_4000,N_3595,N_3141);
or U4001 (N_4001,N_3713,N_3812);
nor U4002 (N_4002,N_3465,N_3246);
and U4003 (N_4003,N_3195,N_3518);
nor U4004 (N_4004,N_3034,N_3940);
xnor U4005 (N_4005,N_3950,N_3997);
nand U4006 (N_4006,N_3572,N_3004);
or U4007 (N_4007,N_3459,N_3776);
nand U4008 (N_4008,N_3882,N_3641);
nor U4009 (N_4009,N_3382,N_3039);
and U4010 (N_4010,N_3969,N_3495);
nor U4011 (N_4011,N_3892,N_3718);
nor U4012 (N_4012,N_3282,N_3388);
nand U4013 (N_4013,N_3489,N_3687);
or U4014 (N_4014,N_3847,N_3856);
or U4015 (N_4015,N_3561,N_3667);
nand U4016 (N_4016,N_3234,N_3135);
or U4017 (N_4017,N_3634,N_3203);
nor U4018 (N_4018,N_3524,N_3149);
and U4019 (N_4019,N_3418,N_3414);
nor U4020 (N_4020,N_3439,N_3804);
or U4021 (N_4021,N_3939,N_3673);
and U4022 (N_4022,N_3824,N_3497);
or U4023 (N_4023,N_3065,N_3769);
xnor U4024 (N_4024,N_3823,N_3333);
xor U4025 (N_4025,N_3581,N_3469);
nand U4026 (N_4026,N_3486,N_3512);
xor U4027 (N_4027,N_3881,N_3636);
or U4028 (N_4028,N_3573,N_3755);
or U4029 (N_4029,N_3154,N_3575);
and U4030 (N_4030,N_3364,N_3980);
nor U4031 (N_4031,N_3528,N_3691);
nand U4032 (N_4032,N_3244,N_3833);
nand U4033 (N_4033,N_3785,N_3952);
and U4034 (N_4034,N_3837,N_3089);
and U4035 (N_4035,N_3336,N_3690);
and U4036 (N_4036,N_3668,N_3194);
and U4037 (N_4037,N_3557,N_3620);
nand U4038 (N_4038,N_3555,N_3240);
and U4039 (N_4039,N_3009,N_3630);
nand U4040 (N_4040,N_3883,N_3844);
or U4041 (N_4041,N_3629,N_3296);
xor U4042 (N_4042,N_3948,N_3097);
and U4043 (N_4043,N_3462,N_3770);
nor U4044 (N_4044,N_3488,N_3662);
nand U4045 (N_4045,N_3242,N_3323);
xor U4046 (N_4046,N_3126,N_3276);
nand U4047 (N_4047,N_3106,N_3519);
nand U4048 (N_4048,N_3565,N_3248);
nand U4049 (N_4049,N_3127,N_3068);
or U4050 (N_4050,N_3332,N_3777);
and U4051 (N_4051,N_3096,N_3016);
xor U4052 (N_4052,N_3263,N_3547);
nand U4053 (N_4053,N_3818,N_3256);
and U4054 (N_4054,N_3029,N_3008);
nor U4055 (N_4055,N_3604,N_3843);
nor U4056 (N_4056,N_3095,N_3836);
or U4057 (N_4057,N_3819,N_3801);
and U4058 (N_4058,N_3476,N_3995);
nand U4059 (N_4059,N_3903,N_3888);
and U4060 (N_4060,N_3485,N_3326);
or U4061 (N_4061,N_3594,N_3808);
and U4062 (N_4062,N_3609,N_3378);
and U4063 (N_4063,N_3092,N_3328);
xor U4064 (N_4064,N_3583,N_3644);
xnor U4065 (N_4065,N_3907,N_3304);
nor U4066 (N_4066,N_3729,N_3120);
nand U4067 (N_4067,N_3803,N_3807);
nand U4068 (N_4068,N_3404,N_3480);
xnor U4069 (N_4069,N_3551,N_3853);
or U4070 (N_4070,N_3360,N_3990);
nor U4071 (N_4071,N_3350,N_3230);
or U4072 (N_4072,N_3612,N_3788);
xnor U4073 (N_4073,N_3945,N_3744);
xnor U4074 (N_4074,N_3470,N_3906);
and U4075 (N_4075,N_3702,N_3928);
xor U4076 (N_4076,N_3429,N_3103);
and U4077 (N_4077,N_3317,N_3078);
xor U4078 (N_4078,N_3767,N_3455);
or U4079 (N_4079,N_3395,N_3757);
nor U4080 (N_4080,N_3142,N_3739);
nor U4081 (N_4081,N_3057,N_3002);
or U4082 (N_4082,N_3381,N_3814);
nand U4083 (N_4083,N_3834,N_3683);
nor U4084 (N_4084,N_3505,N_3558);
nand U4085 (N_4085,N_3471,N_3580);
or U4086 (N_4086,N_3874,N_3637);
and U4087 (N_4087,N_3265,N_3123);
and U4088 (N_4088,N_3199,N_3708);
nor U4089 (N_4089,N_3156,N_3701);
xor U4090 (N_4090,N_3049,N_3973);
nand U4091 (N_4091,N_3845,N_3370);
and U4092 (N_4092,N_3345,N_3977);
nand U4093 (N_4093,N_3310,N_3553);
or U4094 (N_4094,N_3018,N_3921);
nor U4095 (N_4095,N_3198,N_3879);
and U4096 (N_4096,N_3515,N_3937);
xnor U4097 (N_4097,N_3288,N_3251);
xnor U4098 (N_4098,N_3926,N_3077);
nand U4099 (N_4099,N_3165,N_3066);
xor U4100 (N_4100,N_3675,N_3390);
nand U4101 (N_4101,N_3682,N_3746);
or U4102 (N_4102,N_3197,N_3954);
nor U4103 (N_4103,N_3993,N_3955);
or U4104 (N_4104,N_3867,N_3070);
nand U4105 (N_4105,N_3369,N_3262);
nand U4106 (N_4106,N_3301,N_3653);
or U4107 (N_4107,N_3446,N_3438);
nand U4108 (N_4108,N_3221,N_3664);
and U4109 (N_4109,N_3417,N_3764);
and U4110 (N_4110,N_3163,N_3060);
or U4111 (N_4111,N_3058,N_3999);
nor U4112 (N_4112,N_3712,N_3901);
nand U4113 (N_4113,N_3707,N_3130);
or U4114 (N_4114,N_3705,N_3706);
or U4115 (N_4115,N_3622,N_3148);
nand U4116 (N_4116,N_3371,N_3478);
nand U4117 (N_4117,N_3064,N_3405);
xor U4118 (N_4118,N_3972,N_3929);
nor U4119 (N_4119,N_3021,N_3494);
nor U4120 (N_4120,N_3121,N_3107);
or U4121 (N_4121,N_3848,N_3475);
or U4122 (N_4122,N_3711,N_3229);
xnor U4123 (N_4123,N_3855,N_3187);
nor U4124 (N_4124,N_3925,N_3268);
nand U4125 (N_4125,N_3966,N_3436);
nor U4126 (N_4126,N_3665,N_3367);
or U4127 (N_4127,N_3212,N_3179);
nand U4128 (N_4128,N_3780,N_3136);
or U4129 (N_4129,N_3311,N_3491);
xor U4130 (N_4130,N_3958,N_3260);
and U4131 (N_4131,N_3463,N_3700);
nor U4132 (N_4132,N_3696,N_3584);
nor U4133 (N_4133,N_3458,N_3965);
nand U4134 (N_4134,N_3915,N_3619);
nand U4135 (N_4135,N_3544,N_3261);
nor U4136 (N_4136,N_3678,N_3527);
nor U4137 (N_4137,N_3434,N_3694);
and U4138 (N_4138,N_3181,N_3628);
nor U4139 (N_4139,N_3590,N_3428);
nor U4140 (N_4140,N_3292,N_3959);
nor U4141 (N_4141,N_3166,N_3151);
nand U4142 (N_4142,N_3456,N_3468);
or U4143 (N_4143,N_3781,N_3932);
or U4144 (N_4144,N_3758,N_3174);
xor U4145 (N_4145,N_3771,N_3810);
nor U4146 (N_4146,N_3806,N_3258);
nor U4147 (N_4147,N_3075,N_3492);
or U4148 (N_4148,N_3962,N_3137);
nand U4149 (N_4149,N_3502,N_3517);
or U4150 (N_4150,N_3433,N_3738);
or U4151 (N_4151,N_3361,N_3253);
nor U4152 (N_4152,N_3050,N_3271);
or U4153 (N_4153,N_3635,N_3542);
xnor U4154 (N_4154,N_3900,N_3394);
nor U4155 (N_4155,N_3822,N_3787);
or U4156 (N_4156,N_3010,N_3875);
nor U4157 (N_4157,N_3944,N_3927);
or U4158 (N_4158,N_3646,N_3331);
nor U4159 (N_4159,N_3943,N_3209);
or U4160 (N_4160,N_3909,N_3530);
or U4161 (N_4161,N_3571,N_3162);
and U4162 (N_4162,N_3490,N_3207);
nor U4163 (N_4163,N_3805,N_3727);
nand U4164 (N_4164,N_3895,N_3603);
nand U4165 (N_4165,N_3061,N_3793);
nand U4166 (N_4166,N_3750,N_3045);
nor U4167 (N_4167,N_3979,N_3693);
nand U4168 (N_4168,N_3539,N_3125);
nand U4169 (N_4169,N_3540,N_3407);
and U4170 (N_4170,N_3393,N_3661);
and U4171 (N_4171,N_3028,N_3213);
nand U4172 (N_4172,N_3354,N_3192);
or U4173 (N_4173,N_3211,N_3543);
nand U4174 (N_4174,N_3859,N_3625);
or U4175 (N_4175,N_3953,N_3864);
nor U4176 (N_4176,N_3698,N_3252);
and U4177 (N_4177,N_3109,N_3272);
xnor U4178 (N_4178,N_3308,N_3373);
nand U4179 (N_4179,N_3532,N_3286);
xor U4180 (N_4180,N_3379,N_3315);
and U4181 (N_4181,N_3460,N_3257);
nor U4182 (N_4182,N_3986,N_3509);
nand U4183 (N_4183,N_3567,N_3295);
and U4184 (N_4184,N_3910,N_3273);
or U4185 (N_4185,N_3756,N_3440);
nor U4186 (N_4186,N_3223,N_3051);
and U4187 (N_4187,N_3851,N_3117);
nand U4188 (N_4188,N_3415,N_3576);
nor U4189 (N_4189,N_3503,N_3423);
or U4190 (N_4190,N_3356,N_3173);
and U4191 (N_4191,N_3854,N_3365);
nand U4192 (N_4192,N_3281,N_3773);
or U4193 (N_4193,N_3613,N_3143);
and U4194 (N_4194,N_3487,N_3568);
nand U4195 (N_4195,N_3642,N_3586);
nor U4196 (N_4196,N_3098,N_3452);
nand U4197 (N_4197,N_3118,N_3032);
nor U4198 (N_4198,N_3047,N_3305);
xnor U4199 (N_4199,N_3798,N_3374);
and U4200 (N_4200,N_3936,N_3716);
or U4201 (N_4201,N_3931,N_3506);
xor U4202 (N_4202,N_3821,N_3726);
or U4203 (N_4203,N_3104,N_3608);
and U4204 (N_4204,N_3208,N_3355);
and U4205 (N_4205,N_3884,N_3048);
or U4206 (N_4206,N_3412,N_3504);
nor U4207 (N_4207,N_3671,N_3041);
and U4208 (N_4208,N_3432,N_3852);
and U4209 (N_4209,N_3563,N_3782);
nand U4210 (N_4210,N_3796,N_3579);
and U4211 (N_4211,N_3616,N_3055);
nand U4212 (N_4212,N_3912,N_3652);
xnor U4213 (N_4213,N_3627,N_3978);
xnor U4214 (N_4214,N_3402,N_3182);
nor U4215 (N_4215,N_3588,N_3832);
and U4216 (N_4216,N_3160,N_3466);
nor U4217 (N_4217,N_3632,N_3006);
or U4218 (N_4218,N_3084,N_3885);
nand U4219 (N_4219,N_3184,N_3264);
nand U4220 (N_4220,N_3984,N_3383);
and U4221 (N_4221,N_3283,N_3850);
and U4222 (N_4222,N_3663,N_3933);
nand U4223 (N_4223,N_3316,N_3873);
nor U4224 (N_4224,N_3059,N_3728);
or U4225 (N_4225,N_3347,N_3115);
or U4226 (N_4226,N_3090,N_3655);
xnor U4227 (N_4227,N_3645,N_3218);
and U4228 (N_4228,N_3397,N_3387);
nand U4229 (N_4229,N_3964,N_3200);
xor U4230 (N_4230,N_3091,N_3043);
nor U4231 (N_4231,N_3274,N_3243);
or U4232 (N_4232,N_3860,N_3507);
and U4233 (N_4233,N_3435,N_3709);
or U4234 (N_4234,N_3348,N_3139);
or U4235 (N_4235,N_3660,N_3680);
xnor U4236 (N_4236,N_3116,N_3224);
nor U4237 (N_4237,N_3501,N_3259);
nor U4238 (N_4238,N_3871,N_3000);
nor U4239 (N_4239,N_3930,N_3073);
and U4240 (N_4240,N_3217,N_3730);
xor U4241 (N_4241,N_3419,N_3886);
and U4242 (N_4242,N_3145,N_3062);
nor U4243 (N_4243,N_3560,N_3510);
or U4244 (N_4244,N_3731,N_3020);
or U4245 (N_4245,N_3922,N_3119);
or U4246 (N_4246,N_3422,N_3052);
and U4247 (N_4247,N_3724,N_3686);
nand U4248 (N_4248,N_3227,N_3177);
nand U4249 (N_4249,N_3222,N_3880);
nand U4250 (N_4250,N_3826,N_3030);
nand U4251 (N_4251,N_3896,N_3974);
and U4252 (N_4252,N_3684,N_3183);
and U4253 (N_4253,N_3285,N_3745);
or U4254 (N_4254,N_3320,N_3548);
or U4255 (N_4255,N_3623,N_3719);
and U4256 (N_4256,N_3451,N_3552);
and U4257 (N_4257,N_3759,N_3101);
nand U4258 (N_4258,N_3204,N_3359);
or U4259 (N_4259,N_3157,N_3362);
nor U4260 (N_4260,N_3255,N_3180);
nor U4261 (N_4261,N_3094,N_3626);
nand U4262 (N_4262,N_3266,N_3751);
or U4263 (N_4263,N_3113,N_3666);
nand U4264 (N_4264,N_3508,N_3531);
nor U4265 (N_4265,N_3024,N_3067);
nor U4266 (N_4266,N_3914,N_3550);
nand U4267 (N_4267,N_3786,N_3829);
nand U4268 (N_4268,N_3521,N_3441);
nor U4269 (N_4269,N_3516,N_3085);
and U4270 (N_4270,N_3040,N_3774);
xnor U4271 (N_4271,N_3249,N_3161);
or U4272 (N_4272,N_3889,N_3589);
or U4273 (N_4273,N_3005,N_3159);
nand U4274 (N_4274,N_3017,N_3158);
or U4275 (N_4275,N_3453,N_3278);
or U4276 (N_4276,N_3138,N_3302);
and U4277 (N_4277,N_3357,N_3124);
nor U4278 (N_4278,N_3330,N_3300);
xor U4279 (N_4279,N_3564,N_3437);
nand U4280 (N_4280,N_3591,N_3841);
nor U4281 (N_4281,N_3368,N_3099);
or U4282 (N_4282,N_3284,N_3870);
or U4283 (N_4283,N_3175,N_3046);
or U4284 (N_4284,N_3688,N_3538);
nand U4285 (N_4285,N_3743,N_3617);
nor U4286 (N_4286,N_3754,N_3069);
nor U4287 (N_4287,N_3277,N_3386);
and U4288 (N_4288,N_3566,N_3985);
and U4289 (N_4289,N_3778,N_3775);
xnor U4290 (N_4290,N_3890,N_3454);
nor U4291 (N_4291,N_3765,N_3679);
or U4292 (N_4292,N_3014,N_3991);
nand U4293 (N_4293,N_3520,N_3290);
or U4294 (N_4294,N_3868,N_3789);
xor U4295 (N_4295,N_3946,N_3898);
nand U4296 (N_4296,N_3659,N_3114);
nand U4297 (N_4297,N_3722,N_3858);
and U4298 (N_4298,N_3987,N_3989);
or U4299 (N_4299,N_3872,N_3171);
nand U4300 (N_4300,N_3214,N_3839);
nand U4301 (N_4301,N_3658,N_3430);
nor U4302 (N_4302,N_3447,N_3862);
nor U4303 (N_4303,N_3596,N_3790);
nand U4304 (N_4304,N_3086,N_3299);
and U4305 (N_4305,N_3410,N_3267);
and U4306 (N_4306,N_3013,N_3523);
nand U4307 (N_4307,N_3610,N_3377);
xnor U4308 (N_4308,N_3499,N_3245);
and U4309 (N_4309,N_3924,N_3140);
and U4310 (N_4310,N_3335,N_3408);
and U4311 (N_4311,N_3406,N_3254);
or U4312 (N_4312,N_3947,N_3772);
nor U4313 (N_4313,N_3827,N_3353);
and U4314 (N_4314,N_3577,N_3389);
or U4315 (N_4315,N_3319,N_3734);
and U4316 (N_4316,N_3102,N_3384);
nand U4317 (N_4317,N_3768,N_3904);
nor U4318 (N_4318,N_3809,N_3582);
nor U4319 (N_4319,N_3391,N_3122);
nor U4320 (N_4320,N_3971,N_3306);
or U4321 (N_4321,N_3887,N_3297);
and U4322 (N_4322,N_3036,N_3012);
nor U4323 (N_4323,N_3695,N_3082);
and U4324 (N_4324,N_3467,N_3970);
and U4325 (N_4325,N_3830,N_3087);
and U4326 (N_4326,N_3019,N_3275);
and U4327 (N_4327,N_3424,N_3574);
nor U4328 (N_4328,N_3100,N_3797);
nor U4329 (N_4329,N_3654,N_3732);
nor U4330 (N_4330,N_3657,N_3170);
nor U4331 (N_4331,N_3697,N_3513);
nand U4332 (N_4332,N_3536,N_3385);
and U4333 (N_4333,N_3026,N_3189);
nand U4334 (N_4334,N_3598,N_3399);
nand U4335 (N_4335,N_3105,N_3650);
xor U4336 (N_4336,N_3535,N_3293);
or U4337 (N_4337,N_3529,N_3704);
and U4338 (N_4338,N_3537,N_3236);
nand U4339 (N_4339,N_3951,N_3185);
nor U4340 (N_4340,N_3413,N_3420);
nand U4341 (N_4341,N_3800,N_3007);
nor U4342 (N_4342,N_3753,N_3640);
and U4343 (N_4343,N_3380,N_3220);
nand U4344 (N_4344,N_3349,N_3396);
nor U4345 (N_4345,N_3562,N_3134);
and U4346 (N_4346,N_3720,N_3846);
nor U4347 (N_4347,N_3038,N_3983);
nor U4348 (N_4348,N_3742,N_3811);
and U4349 (N_4349,N_3996,N_3309);
nor U4350 (N_4350,N_3554,N_3201);
nor U4351 (N_4351,N_3559,N_3474);
nand U4352 (N_4352,N_3401,N_3093);
nor U4353 (N_4353,N_3919,N_3534);
and U4354 (N_4354,N_3941,N_3992);
and U4355 (N_4355,N_3916,N_3442);
and U4356 (N_4356,N_3079,N_3376);
nor U4357 (N_4357,N_3219,N_3699);
and U4358 (N_4358,N_3083,N_3011);
nand U4359 (N_4359,N_3760,N_3146);
or U4360 (N_4360,N_3816,N_3444);
xor U4361 (N_4361,N_3820,N_3541);
nor U4362 (N_4362,N_3715,N_3291);
or U4363 (N_4363,N_3398,N_3842);
nor U4364 (N_4364,N_3270,N_3615);
or U4365 (N_4365,N_3313,N_3597);
nand U4366 (N_4366,N_3164,N_3196);
nor U4367 (N_4367,N_3496,N_3112);
and U4368 (N_4368,N_3714,N_3339);
nand U4369 (N_4369,N_3908,N_3611);
nor U4370 (N_4370,N_3733,N_3215);
and U4371 (N_4371,N_3238,N_3232);
nand U4372 (N_4372,N_3131,N_3526);
and U4373 (N_4373,N_3913,N_3600);
or U4374 (N_4374,N_3585,N_3735);
or U4375 (N_4375,N_3749,N_3366);
or U4376 (N_4376,N_3152,N_3570);
nor U4377 (N_4377,N_3602,N_3674);
and U4378 (N_4378,N_3685,N_3792);
or U4379 (N_4379,N_3477,N_3840);
and U4380 (N_4380,N_3737,N_3403);
or U4381 (N_4381,N_3001,N_3071);
and U4382 (N_4382,N_3147,N_3457);
nand U4383 (N_4383,N_3035,N_3421);
nor U4384 (N_4384,N_3624,N_3168);
and U4385 (N_4385,N_3761,N_3228);
nor U4386 (N_4386,N_3400,N_3464);
xor U4387 (N_4387,N_3338,N_3917);
or U4388 (N_4388,N_3762,N_3279);
nor U4389 (N_4389,N_3322,N_3838);
nand U4390 (N_4390,N_3072,N_3416);
nand U4391 (N_4391,N_3473,N_3703);
and U4392 (N_4392,N_3618,N_3968);
or U4393 (N_4393,N_3934,N_3191);
nand U4394 (N_4394,N_3111,N_3639);
and U4395 (N_4395,N_3784,N_3828);
and U4396 (N_4396,N_3525,N_3053);
and U4397 (N_4397,N_3717,N_3643);
nand U4398 (N_4398,N_3500,N_3269);
and U4399 (N_4399,N_3692,N_3076);
nor U4400 (N_4400,N_3479,N_3003);
and U4401 (N_4401,N_3905,N_3815);
xnor U4402 (N_4402,N_3031,N_3153);
xor U4403 (N_4403,N_3923,N_3710);
nand U4404 (N_4404,N_3763,N_3247);
nor U4405 (N_4405,N_3144,N_3605);
and U4406 (N_4406,N_3150,N_3294);
and U4407 (N_4407,N_3647,N_3994);
and U4408 (N_4408,N_3949,N_3344);
nand U4409 (N_4409,N_3472,N_3894);
and U4410 (N_4410,N_3411,N_3795);
and U4411 (N_4411,N_3186,N_3817);
or U4412 (N_4412,N_3802,N_3607);
and U4413 (N_4413,N_3878,N_3237);
and U4414 (N_4414,N_3298,N_3649);
and U4415 (N_4415,N_3448,N_3172);
or U4416 (N_4416,N_3975,N_3963);
nand U4417 (N_4417,N_3129,N_3445);
or U4418 (N_4418,N_3250,N_3409);
xor U4419 (N_4419,N_3813,N_3280);
nor U4420 (N_4420,N_3741,N_3863);
xor U4421 (N_4421,N_3231,N_3676);
nor U4422 (N_4422,N_3748,N_3314);
or U4423 (N_4423,N_3461,N_3303);
nor U4424 (N_4424,N_3897,N_3648);
nor U4425 (N_4425,N_3877,N_3202);
xor U4426 (N_4426,N_3342,N_3015);
or U4427 (N_4427,N_3631,N_3791);
and U4428 (N_4428,N_3312,N_3606);
or U4429 (N_4429,N_3723,N_3857);
or U4430 (N_4430,N_3651,N_3037);
xnor U4431 (N_4431,N_3918,N_3482);
and U4432 (N_4432,N_3831,N_3375);
or U4433 (N_4433,N_3998,N_3210);
or U4434 (N_4434,N_3981,N_3329);
xor U4435 (N_4435,N_3023,N_3920);
and U4436 (N_4436,N_3167,N_3340);
xnor U4437 (N_4437,N_3235,N_3522);
nand U4438 (N_4438,N_3358,N_3307);
nor U4439 (N_4439,N_3556,N_3022);
xor U4440 (N_4440,N_3861,N_3783);
or U4441 (N_4441,N_3108,N_3902);
nand U4442 (N_4442,N_3155,N_3938);
nand U4443 (N_4443,N_3351,N_3074);
xnor U4444 (N_4444,N_3876,N_3601);
and U4445 (N_4445,N_3239,N_3587);
and U4446 (N_4446,N_3960,N_3677);
nor U4447 (N_4447,N_3614,N_3545);
nand U4448 (N_4448,N_3935,N_3206);
and U4449 (N_4449,N_3766,N_3431);
nor U4450 (N_4450,N_3893,N_3233);
or U4451 (N_4451,N_3216,N_3865);
or U4452 (N_4452,N_3670,N_3835);
or U4453 (N_4453,N_3325,N_3533);
nand U4454 (N_4454,N_3080,N_3942);
and U4455 (N_4455,N_3427,N_3961);
and U4456 (N_4456,N_3638,N_3132);
xnor U4457 (N_4457,N_3483,N_3721);
nand U4458 (N_4458,N_3511,N_3967);
nand U4459 (N_4459,N_3176,N_3569);
and U4460 (N_4460,N_3740,N_3443);
or U4461 (N_4461,N_3110,N_3226);
or U4462 (N_4462,N_3493,N_3169);
and U4463 (N_4463,N_3736,N_3341);
or U4464 (N_4464,N_3689,N_3794);
and U4465 (N_4465,N_3289,N_3205);
xor U4466 (N_4466,N_3321,N_3063);
xnor U4467 (N_4467,N_3337,N_3287);
nor U4468 (N_4468,N_3033,N_3514);
and U4469 (N_4469,N_3956,N_3866);
or U4470 (N_4470,N_3799,N_3363);
or U4471 (N_4471,N_3621,N_3825);
and U4472 (N_4472,N_3449,N_3752);
xor U4473 (N_4473,N_3779,N_3042);
xor U4474 (N_4474,N_3725,N_3225);
and U4475 (N_4475,N_3484,N_3188);
nor U4476 (N_4476,N_3128,N_3747);
nor U4477 (N_4477,N_3178,N_3426);
or U4478 (N_4478,N_3633,N_3988);
nand U4479 (N_4479,N_3027,N_3425);
nand U4480 (N_4480,N_3372,N_3044);
nand U4481 (N_4481,N_3982,N_3334);
or U4482 (N_4482,N_3672,N_3190);
and U4483 (N_4483,N_3592,N_3849);
nor U4484 (N_4484,N_3450,N_3241);
and U4485 (N_4485,N_3599,N_3498);
and U4486 (N_4486,N_3324,N_3899);
and U4487 (N_4487,N_3957,N_3352);
or U4488 (N_4488,N_3318,N_3343);
and U4489 (N_4489,N_3656,N_3546);
xnor U4490 (N_4490,N_3327,N_3025);
and U4491 (N_4491,N_3392,N_3193);
or U4492 (N_4492,N_3056,N_3081);
and U4493 (N_4493,N_3054,N_3578);
nand U4494 (N_4494,N_3681,N_3593);
xor U4495 (N_4495,N_3891,N_3669);
nor U4496 (N_4496,N_3976,N_3911);
and U4497 (N_4497,N_3549,N_3133);
and U4498 (N_4498,N_3346,N_3088);
and U4499 (N_4499,N_3481,N_3869);
and U4500 (N_4500,N_3342,N_3305);
nand U4501 (N_4501,N_3588,N_3006);
or U4502 (N_4502,N_3888,N_3029);
nor U4503 (N_4503,N_3278,N_3793);
and U4504 (N_4504,N_3259,N_3590);
or U4505 (N_4505,N_3612,N_3167);
and U4506 (N_4506,N_3239,N_3613);
nor U4507 (N_4507,N_3149,N_3532);
or U4508 (N_4508,N_3473,N_3730);
nor U4509 (N_4509,N_3616,N_3463);
xnor U4510 (N_4510,N_3468,N_3415);
or U4511 (N_4511,N_3073,N_3108);
or U4512 (N_4512,N_3413,N_3800);
or U4513 (N_4513,N_3316,N_3789);
or U4514 (N_4514,N_3002,N_3022);
nand U4515 (N_4515,N_3102,N_3911);
nor U4516 (N_4516,N_3446,N_3990);
nor U4517 (N_4517,N_3737,N_3749);
nor U4518 (N_4518,N_3309,N_3271);
and U4519 (N_4519,N_3602,N_3776);
or U4520 (N_4520,N_3149,N_3441);
nor U4521 (N_4521,N_3448,N_3619);
and U4522 (N_4522,N_3496,N_3588);
or U4523 (N_4523,N_3664,N_3744);
nor U4524 (N_4524,N_3895,N_3962);
nand U4525 (N_4525,N_3243,N_3500);
nor U4526 (N_4526,N_3142,N_3616);
nor U4527 (N_4527,N_3342,N_3185);
nor U4528 (N_4528,N_3349,N_3554);
or U4529 (N_4529,N_3214,N_3463);
or U4530 (N_4530,N_3839,N_3405);
xnor U4531 (N_4531,N_3101,N_3417);
or U4532 (N_4532,N_3936,N_3228);
xnor U4533 (N_4533,N_3297,N_3519);
nor U4534 (N_4534,N_3236,N_3539);
nand U4535 (N_4535,N_3514,N_3206);
nor U4536 (N_4536,N_3428,N_3543);
nor U4537 (N_4537,N_3273,N_3254);
or U4538 (N_4538,N_3180,N_3664);
and U4539 (N_4539,N_3088,N_3105);
xor U4540 (N_4540,N_3206,N_3198);
or U4541 (N_4541,N_3418,N_3801);
and U4542 (N_4542,N_3829,N_3400);
nor U4543 (N_4543,N_3296,N_3541);
xnor U4544 (N_4544,N_3042,N_3348);
nand U4545 (N_4545,N_3052,N_3466);
and U4546 (N_4546,N_3188,N_3228);
nor U4547 (N_4547,N_3046,N_3880);
and U4548 (N_4548,N_3571,N_3800);
nand U4549 (N_4549,N_3729,N_3692);
or U4550 (N_4550,N_3966,N_3241);
or U4551 (N_4551,N_3346,N_3429);
nand U4552 (N_4552,N_3035,N_3032);
and U4553 (N_4553,N_3179,N_3553);
nand U4554 (N_4554,N_3519,N_3146);
nand U4555 (N_4555,N_3728,N_3261);
nand U4556 (N_4556,N_3574,N_3981);
nor U4557 (N_4557,N_3754,N_3033);
or U4558 (N_4558,N_3545,N_3651);
nor U4559 (N_4559,N_3052,N_3853);
nor U4560 (N_4560,N_3251,N_3417);
nand U4561 (N_4561,N_3550,N_3370);
and U4562 (N_4562,N_3650,N_3100);
and U4563 (N_4563,N_3280,N_3574);
nand U4564 (N_4564,N_3024,N_3233);
nand U4565 (N_4565,N_3992,N_3874);
nand U4566 (N_4566,N_3742,N_3590);
xor U4567 (N_4567,N_3497,N_3802);
and U4568 (N_4568,N_3274,N_3724);
nor U4569 (N_4569,N_3585,N_3704);
nor U4570 (N_4570,N_3261,N_3659);
or U4571 (N_4571,N_3087,N_3624);
or U4572 (N_4572,N_3664,N_3688);
and U4573 (N_4573,N_3111,N_3284);
nor U4574 (N_4574,N_3511,N_3902);
and U4575 (N_4575,N_3833,N_3022);
nor U4576 (N_4576,N_3315,N_3117);
and U4577 (N_4577,N_3213,N_3109);
nand U4578 (N_4578,N_3812,N_3540);
nor U4579 (N_4579,N_3911,N_3559);
nand U4580 (N_4580,N_3623,N_3994);
and U4581 (N_4581,N_3627,N_3076);
and U4582 (N_4582,N_3897,N_3593);
and U4583 (N_4583,N_3871,N_3329);
nand U4584 (N_4584,N_3843,N_3463);
nor U4585 (N_4585,N_3476,N_3098);
nand U4586 (N_4586,N_3655,N_3399);
and U4587 (N_4587,N_3211,N_3979);
and U4588 (N_4588,N_3692,N_3377);
xnor U4589 (N_4589,N_3549,N_3788);
or U4590 (N_4590,N_3698,N_3703);
nand U4591 (N_4591,N_3627,N_3132);
or U4592 (N_4592,N_3227,N_3973);
nand U4593 (N_4593,N_3574,N_3688);
and U4594 (N_4594,N_3010,N_3009);
and U4595 (N_4595,N_3868,N_3165);
nor U4596 (N_4596,N_3368,N_3905);
and U4597 (N_4597,N_3325,N_3571);
or U4598 (N_4598,N_3780,N_3394);
or U4599 (N_4599,N_3397,N_3575);
and U4600 (N_4600,N_3218,N_3894);
or U4601 (N_4601,N_3765,N_3561);
nor U4602 (N_4602,N_3733,N_3540);
or U4603 (N_4603,N_3067,N_3313);
xnor U4604 (N_4604,N_3630,N_3319);
nor U4605 (N_4605,N_3712,N_3178);
nor U4606 (N_4606,N_3500,N_3827);
nand U4607 (N_4607,N_3394,N_3362);
xor U4608 (N_4608,N_3497,N_3059);
and U4609 (N_4609,N_3634,N_3108);
nor U4610 (N_4610,N_3119,N_3477);
or U4611 (N_4611,N_3933,N_3034);
or U4612 (N_4612,N_3019,N_3147);
or U4613 (N_4613,N_3053,N_3570);
or U4614 (N_4614,N_3060,N_3825);
nor U4615 (N_4615,N_3973,N_3170);
and U4616 (N_4616,N_3672,N_3346);
or U4617 (N_4617,N_3178,N_3484);
nand U4618 (N_4618,N_3620,N_3010);
nand U4619 (N_4619,N_3945,N_3576);
or U4620 (N_4620,N_3000,N_3185);
nor U4621 (N_4621,N_3507,N_3513);
nor U4622 (N_4622,N_3221,N_3441);
or U4623 (N_4623,N_3866,N_3254);
nand U4624 (N_4624,N_3920,N_3195);
nor U4625 (N_4625,N_3079,N_3868);
nor U4626 (N_4626,N_3954,N_3949);
nor U4627 (N_4627,N_3342,N_3817);
nand U4628 (N_4628,N_3802,N_3170);
or U4629 (N_4629,N_3788,N_3882);
xor U4630 (N_4630,N_3152,N_3129);
and U4631 (N_4631,N_3213,N_3166);
or U4632 (N_4632,N_3927,N_3933);
xnor U4633 (N_4633,N_3633,N_3872);
and U4634 (N_4634,N_3422,N_3894);
and U4635 (N_4635,N_3342,N_3875);
nor U4636 (N_4636,N_3387,N_3916);
and U4637 (N_4637,N_3766,N_3584);
or U4638 (N_4638,N_3813,N_3381);
and U4639 (N_4639,N_3051,N_3042);
and U4640 (N_4640,N_3236,N_3925);
nor U4641 (N_4641,N_3061,N_3825);
and U4642 (N_4642,N_3966,N_3984);
nor U4643 (N_4643,N_3188,N_3362);
or U4644 (N_4644,N_3056,N_3139);
and U4645 (N_4645,N_3757,N_3422);
or U4646 (N_4646,N_3804,N_3289);
xnor U4647 (N_4647,N_3277,N_3782);
nand U4648 (N_4648,N_3513,N_3622);
and U4649 (N_4649,N_3048,N_3171);
nor U4650 (N_4650,N_3395,N_3089);
and U4651 (N_4651,N_3387,N_3939);
or U4652 (N_4652,N_3708,N_3735);
or U4653 (N_4653,N_3363,N_3013);
nor U4654 (N_4654,N_3052,N_3425);
nand U4655 (N_4655,N_3252,N_3856);
nor U4656 (N_4656,N_3618,N_3021);
or U4657 (N_4657,N_3940,N_3219);
and U4658 (N_4658,N_3020,N_3733);
nand U4659 (N_4659,N_3944,N_3763);
xnor U4660 (N_4660,N_3936,N_3913);
nand U4661 (N_4661,N_3795,N_3781);
and U4662 (N_4662,N_3041,N_3903);
and U4663 (N_4663,N_3883,N_3231);
nor U4664 (N_4664,N_3446,N_3290);
nand U4665 (N_4665,N_3460,N_3124);
and U4666 (N_4666,N_3175,N_3762);
nand U4667 (N_4667,N_3230,N_3553);
nor U4668 (N_4668,N_3448,N_3864);
nor U4669 (N_4669,N_3553,N_3994);
and U4670 (N_4670,N_3517,N_3456);
and U4671 (N_4671,N_3906,N_3723);
or U4672 (N_4672,N_3248,N_3888);
and U4673 (N_4673,N_3189,N_3917);
xor U4674 (N_4674,N_3361,N_3061);
nand U4675 (N_4675,N_3706,N_3443);
nand U4676 (N_4676,N_3592,N_3660);
nor U4677 (N_4677,N_3271,N_3763);
and U4678 (N_4678,N_3577,N_3396);
nor U4679 (N_4679,N_3483,N_3064);
nand U4680 (N_4680,N_3232,N_3802);
nand U4681 (N_4681,N_3813,N_3260);
nand U4682 (N_4682,N_3017,N_3698);
nand U4683 (N_4683,N_3663,N_3253);
or U4684 (N_4684,N_3839,N_3211);
nand U4685 (N_4685,N_3377,N_3164);
nor U4686 (N_4686,N_3019,N_3309);
and U4687 (N_4687,N_3853,N_3771);
nor U4688 (N_4688,N_3529,N_3750);
xor U4689 (N_4689,N_3401,N_3398);
nor U4690 (N_4690,N_3929,N_3288);
or U4691 (N_4691,N_3431,N_3324);
nand U4692 (N_4692,N_3381,N_3799);
nand U4693 (N_4693,N_3477,N_3896);
nor U4694 (N_4694,N_3769,N_3074);
xor U4695 (N_4695,N_3291,N_3467);
or U4696 (N_4696,N_3694,N_3989);
nand U4697 (N_4697,N_3506,N_3828);
and U4698 (N_4698,N_3923,N_3980);
nor U4699 (N_4699,N_3666,N_3179);
xor U4700 (N_4700,N_3244,N_3967);
or U4701 (N_4701,N_3134,N_3190);
and U4702 (N_4702,N_3832,N_3024);
and U4703 (N_4703,N_3220,N_3189);
xnor U4704 (N_4704,N_3425,N_3949);
xnor U4705 (N_4705,N_3754,N_3174);
and U4706 (N_4706,N_3479,N_3298);
and U4707 (N_4707,N_3936,N_3331);
or U4708 (N_4708,N_3592,N_3791);
nand U4709 (N_4709,N_3612,N_3842);
nand U4710 (N_4710,N_3542,N_3247);
nor U4711 (N_4711,N_3997,N_3842);
or U4712 (N_4712,N_3007,N_3911);
nand U4713 (N_4713,N_3166,N_3944);
nand U4714 (N_4714,N_3723,N_3858);
and U4715 (N_4715,N_3757,N_3649);
or U4716 (N_4716,N_3255,N_3909);
or U4717 (N_4717,N_3999,N_3272);
nor U4718 (N_4718,N_3089,N_3379);
or U4719 (N_4719,N_3173,N_3336);
nand U4720 (N_4720,N_3847,N_3848);
and U4721 (N_4721,N_3063,N_3624);
or U4722 (N_4722,N_3407,N_3276);
nand U4723 (N_4723,N_3300,N_3431);
and U4724 (N_4724,N_3293,N_3696);
nand U4725 (N_4725,N_3373,N_3278);
or U4726 (N_4726,N_3891,N_3685);
nor U4727 (N_4727,N_3733,N_3492);
nor U4728 (N_4728,N_3226,N_3067);
and U4729 (N_4729,N_3339,N_3681);
and U4730 (N_4730,N_3333,N_3151);
and U4731 (N_4731,N_3103,N_3293);
and U4732 (N_4732,N_3537,N_3169);
nand U4733 (N_4733,N_3100,N_3986);
and U4734 (N_4734,N_3554,N_3242);
nand U4735 (N_4735,N_3309,N_3759);
nor U4736 (N_4736,N_3977,N_3219);
and U4737 (N_4737,N_3584,N_3479);
and U4738 (N_4738,N_3979,N_3933);
or U4739 (N_4739,N_3787,N_3065);
and U4740 (N_4740,N_3639,N_3649);
and U4741 (N_4741,N_3408,N_3967);
xor U4742 (N_4742,N_3109,N_3254);
or U4743 (N_4743,N_3838,N_3445);
nand U4744 (N_4744,N_3455,N_3062);
nand U4745 (N_4745,N_3072,N_3541);
or U4746 (N_4746,N_3502,N_3915);
nand U4747 (N_4747,N_3721,N_3459);
nor U4748 (N_4748,N_3832,N_3675);
or U4749 (N_4749,N_3234,N_3318);
and U4750 (N_4750,N_3494,N_3768);
nand U4751 (N_4751,N_3430,N_3055);
nor U4752 (N_4752,N_3931,N_3196);
or U4753 (N_4753,N_3984,N_3071);
or U4754 (N_4754,N_3167,N_3128);
and U4755 (N_4755,N_3909,N_3605);
nand U4756 (N_4756,N_3720,N_3508);
or U4757 (N_4757,N_3002,N_3604);
or U4758 (N_4758,N_3345,N_3839);
nor U4759 (N_4759,N_3402,N_3210);
nand U4760 (N_4760,N_3981,N_3697);
and U4761 (N_4761,N_3866,N_3616);
nor U4762 (N_4762,N_3605,N_3853);
nor U4763 (N_4763,N_3234,N_3078);
nor U4764 (N_4764,N_3669,N_3045);
nor U4765 (N_4765,N_3186,N_3874);
nor U4766 (N_4766,N_3742,N_3721);
xor U4767 (N_4767,N_3816,N_3027);
nor U4768 (N_4768,N_3160,N_3769);
nor U4769 (N_4769,N_3571,N_3565);
xnor U4770 (N_4770,N_3326,N_3772);
and U4771 (N_4771,N_3004,N_3445);
or U4772 (N_4772,N_3507,N_3282);
nor U4773 (N_4773,N_3853,N_3327);
nor U4774 (N_4774,N_3681,N_3031);
nand U4775 (N_4775,N_3449,N_3262);
nand U4776 (N_4776,N_3034,N_3178);
nor U4777 (N_4777,N_3303,N_3802);
or U4778 (N_4778,N_3629,N_3171);
and U4779 (N_4779,N_3903,N_3610);
nor U4780 (N_4780,N_3505,N_3479);
nand U4781 (N_4781,N_3088,N_3198);
and U4782 (N_4782,N_3899,N_3844);
or U4783 (N_4783,N_3904,N_3781);
nor U4784 (N_4784,N_3854,N_3146);
nand U4785 (N_4785,N_3392,N_3595);
nor U4786 (N_4786,N_3322,N_3062);
or U4787 (N_4787,N_3380,N_3402);
xnor U4788 (N_4788,N_3117,N_3774);
or U4789 (N_4789,N_3737,N_3550);
and U4790 (N_4790,N_3776,N_3992);
nor U4791 (N_4791,N_3138,N_3242);
nand U4792 (N_4792,N_3655,N_3674);
xnor U4793 (N_4793,N_3124,N_3854);
nor U4794 (N_4794,N_3464,N_3076);
and U4795 (N_4795,N_3862,N_3820);
and U4796 (N_4796,N_3694,N_3815);
nor U4797 (N_4797,N_3820,N_3342);
or U4798 (N_4798,N_3296,N_3559);
nor U4799 (N_4799,N_3454,N_3041);
or U4800 (N_4800,N_3219,N_3703);
nor U4801 (N_4801,N_3300,N_3461);
nand U4802 (N_4802,N_3180,N_3602);
nand U4803 (N_4803,N_3513,N_3746);
nand U4804 (N_4804,N_3394,N_3238);
nor U4805 (N_4805,N_3640,N_3341);
nand U4806 (N_4806,N_3773,N_3970);
nand U4807 (N_4807,N_3642,N_3428);
nor U4808 (N_4808,N_3394,N_3359);
or U4809 (N_4809,N_3812,N_3625);
or U4810 (N_4810,N_3455,N_3148);
or U4811 (N_4811,N_3327,N_3392);
and U4812 (N_4812,N_3532,N_3101);
or U4813 (N_4813,N_3273,N_3829);
and U4814 (N_4814,N_3703,N_3862);
xnor U4815 (N_4815,N_3793,N_3986);
nor U4816 (N_4816,N_3299,N_3593);
and U4817 (N_4817,N_3553,N_3406);
nor U4818 (N_4818,N_3687,N_3884);
or U4819 (N_4819,N_3166,N_3017);
or U4820 (N_4820,N_3104,N_3899);
nor U4821 (N_4821,N_3826,N_3679);
or U4822 (N_4822,N_3101,N_3328);
and U4823 (N_4823,N_3114,N_3376);
and U4824 (N_4824,N_3926,N_3326);
or U4825 (N_4825,N_3390,N_3224);
nand U4826 (N_4826,N_3933,N_3337);
or U4827 (N_4827,N_3219,N_3501);
or U4828 (N_4828,N_3191,N_3759);
and U4829 (N_4829,N_3259,N_3492);
or U4830 (N_4830,N_3161,N_3715);
and U4831 (N_4831,N_3053,N_3551);
or U4832 (N_4832,N_3197,N_3726);
or U4833 (N_4833,N_3302,N_3580);
nor U4834 (N_4834,N_3830,N_3177);
and U4835 (N_4835,N_3895,N_3528);
or U4836 (N_4836,N_3589,N_3965);
or U4837 (N_4837,N_3846,N_3666);
and U4838 (N_4838,N_3008,N_3139);
nand U4839 (N_4839,N_3879,N_3170);
nor U4840 (N_4840,N_3518,N_3713);
nor U4841 (N_4841,N_3963,N_3931);
or U4842 (N_4842,N_3968,N_3120);
nor U4843 (N_4843,N_3728,N_3627);
nand U4844 (N_4844,N_3181,N_3032);
or U4845 (N_4845,N_3045,N_3395);
and U4846 (N_4846,N_3592,N_3725);
nand U4847 (N_4847,N_3417,N_3013);
and U4848 (N_4848,N_3166,N_3487);
or U4849 (N_4849,N_3702,N_3457);
or U4850 (N_4850,N_3866,N_3292);
xnor U4851 (N_4851,N_3143,N_3862);
nand U4852 (N_4852,N_3042,N_3914);
and U4853 (N_4853,N_3277,N_3596);
or U4854 (N_4854,N_3172,N_3538);
xnor U4855 (N_4855,N_3039,N_3020);
and U4856 (N_4856,N_3771,N_3685);
xnor U4857 (N_4857,N_3706,N_3397);
nand U4858 (N_4858,N_3983,N_3096);
nand U4859 (N_4859,N_3798,N_3398);
xor U4860 (N_4860,N_3568,N_3042);
nand U4861 (N_4861,N_3752,N_3652);
xnor U4862 (N_4862,N_3381,N_3522);
xor U4863 (N_4863,N_3544,N_3540);
and U4864 (N_4864,N_3443,N_3500);
nand U4865 (N_4865,N_3048,N_3836);
nand U4866 (N_4866,N_3628,N_3389);
xor U4867 (N_4867,N_3904,N_3236);
and U4868 (N_4868,N_3056,N_3274);
and U4869 (N_4869,N_3321,N_3118);
nor U4870 (N_4870,N_3980,N_3529);
nand U4871 (N_4871,N_3422,N_3906);
or U4872 (N_4872,N_3495,N_3447);
nand U4873 (N_4873,N_3852,N_3717);
or U4874 (N_4874,N_3117,N_3514);
nor U4875 (N_4875,N_3898,N_3835);
nand U4876 (N_4876,N_3552,N_3954);
nand U4877 (N_4877,N_3971,N_3366);
nor U4878 (N_4878,N_3006,N_3497);
or U4879 (N_4879,N_3972,N_3476);
nor U4880 (N_4880,N_3803,N_3311);
nand U4881 (N_4881,N_3120,N_3505);
nand U4882 (N_4882,N_3507,N_3025);
nand U4883 (N_4883,N_3912,N_3193);
or U4884 (N_4884,N_3251,N_3133);
nand U4885 (N_4885,N_3238,N_3623);
xnor U4886 (N_4886,N_3613,N_3555);
nor U4887 (N_4887,N_3565,N_3846);
or U4888 (N_4888,N_3859,N_3039);
nand U4889 (N_4889,N_3374,N_3846);
and U4890 (N_4890,N_3211,N_3398);
nand U4891 (N_4891,N_3425,N_3731);
or U4892 (N_4892,N_3096,N_3857);
nand U4893 (N_4893,N_3412,N_3212);
nor U4894 (N_4894,N_3718,N_3954);
or U4895 (N_4895,N_3336,N_3777);
or U4896 (N_4896,N_3811,N_3979);
or U4897 (N_4897,N_3612,N_3182);
or U4898 (N_4898,N_3413,N_3281);
and U4899 (N_4899,N_3774,N_3416);
nand U4900 (N_4900,N_3597,N_3446);
or U4901 (N_4901,N_3617,N_3983);
nand U4902 (N_4902,N_3012,N_3521);
nand U4903 (N_4903,N_3709,N_3570);
nor U4904 (N_4904,N_3690,N_3433);
nor U4905 (N_4905,N_3132,N_3084);
and U4906 (N_4906,N_3533,N_3328);
and U4907 (N_4907,N_3002,N_3324);
nand U4908 (N_4908,N_3424,N_3546);
nor U4909 (N_4909,N_3534,N_3166);
nand U4910 (N_4910,N_3808,N_3708);
nor U4911 (N_4911,N_3508,N_3533);
and U4912 (N_4912,N_3871,N_3485);
or U4913 (N_4913,N_3099,N_3370);
or U4914 (N_4914,N_3432,N_3900);
and U4915 (N_4915,N_3791,N_3866);
nand U4916 (N_4916,N_3116,N_3304);
nor U4917 (N_4917,N_3291,N_3750);
and U4918 (N_4918,N_3827,N_3883);
or U4919 (N_4919,N_3945,N_3707);
nor U4920 (N_4920,N_3917,N_3637);
or U4921 (N_4921,N_3283,N_3052);
nand U4922 (N_4922,N_3090,N_3826);
nor U4923 (N_4923,N_3737,N_3619);
nor U4924 (N_4924,N_3811,N_3791);
nand U4925 (N_4925,N_3153,N_3118);
and U4926 (N_4926,N_3357,N_3796);
and U4927 (N_4927,N_3312,N_3179);
or U4928 (N_4928,N_3988,N_3024);
xnor U4929 (N_4929,N_3142,N_3021);
nor U4930 (N_4930,N_3989,N_3470);
nor U4931 (N_4931,N_3837,N_3999);
nand U4932 (N_4932,N_3159,N_3479);
nand U4933 (N_4933,N_3181,N_3576);
or U4934 (N_4934,N_3742,N_3731);
and U4935 (N_4935,N_3246,N_3631);
nand U4936 (N_4936,N_3520,N_3280);
and U4937 (N_4937,N_3626,N_3034);
and U4938 (N_4938,N_3304,N_3639);
and U4939 (N_4939,N_3335,N_3043);
nand U4940 (N_4940,N_3437,N_3542);
or U4941 (N_4941,N_3947,N_3966);
nand U4942 (N_4942,N_3934,N_3206);
xor U4943 (N_4943,N_3524,N_3992);
nand U4944 (N_4944,N_3014,N_3084);
or U4945 (N_4945,N_3589,N_3076);
nor U4946 (N_4946,N_3480,N_3789);
or U4947 (N_4947,N_3982,N_3294);
and U4948 (N_4948,N_3505,N_3239);
nand U4949 (N_4949,N_3468,N_3484);
or U4950 (N_4950,N_3936,N_3412);
nand U4951 (N_4951,N_3265,N_3475);
xor U4952 (N_4952,N_3085,N_3495);
nand U4953 (N_4953,N_3423,N_3858);
and U4954 (N_4954,N_3136,N_3222);
nand U4955 (N_4955,N_3191,N_3699);
or U4956 (N_4956,N_3541,N_3407);
or U4957 (N_4957,N_3935,N_3357);
and U4958 (N_4958,N_3644,N_3229);
nor U4959 (N_4959,N_3737,N_3508);
and U4960 (N_4960,N_3919,N_3866);
nor U4961 (N_4961,N_3235,N_3565);
nand U4962 (N_4962,N_3361,N_3044);
nand U4963 (N_4963,N_3543,N_3556);
nand U4964 (N_4964,N_3548,N_3008);
nor U4965 (N_4965,N_3660,N_3247);
nand U4966 (N_4966,N_3873,N_3403);
nor U4967 (N_4967,N_3368,N_3446);
and U4968 (N_4968,N_3308,N_3909);
and U4969 (N_4969,N_3988,N_3983);
nand U4970 (N_4970,N_3149,N_3602);
nor U4971 (N_4971,N_3981,N_3321);
or U4972 (N_4972,N_3588,N_3363);
nand U4973 (N_4973,N_3669,N_3878);
and U4974 (N_4974,N_3905,N_3330);
or U4975 (N_4975,N_3521,N_3544);
or U4976 (N_4976,N_3982,N_3215);
or U4977 (N_4977,N_3990,N_3364);
and U4978 (N_4978,N_3812,N_3565);
nand U4979 (N_4979,N_3743,N_3458);
nor U4980 (N_4980,N_3178,N_3701);
nor U4981 (N_4981,N_3297,N_3570);
and U4982 (N_4982,N_3622,N_3883);
and U4983 (N_4983,N_3097,N_3601);
or U4984 (N_4984,N_3448,N_3794);
xor U4985 (N_4985,N_3002,N_3757);
or U4986 (N_4986,N_3630,N_3890);
or U4987 (N_4987,N_3343,N_3644);
nand U4988 (N_4988,N_3164,N_3390);
or U4989 (N_4989,N_3440,N_3033);
xnor U4990 (N_4990,N_3969,N_3292);
and U4991 (N_4991,N_3475,N_3315);
and U4992 (N_4992,N_3673,N_3945);
xnor U4993 (N_4993,N_3230,N_3064);
nand U4994 (N_4994,N_3304,N_3144);
or U4995 (N_4995,N_3487,N_3754);
and U4996 (N_4996,N_3035,N_3960);
nand U4997 (N_4997,N_3932,N_3090);
nand U4998 (N_4998,N_3309,N_3249);
nor U4999 (N_4999,N_3896,N_3764);
and U5000 (N_5000,N_4778,N_4490);
xnor U5001 (N_5001,N_4426,N_4488);
or U5002 (N_5002,N_4540,N_4724);
or U5003 (N_5003,N_4626,N_4777);
nor U5004 (N_5004,N_4604,N_4562);
nand U5005 (N_5005,N_4081,N_4617);
nand U5006 (N_5006,N_4761,N_4551);
and U5007 (N_5007,N_4500,N_4634);
and U5008 (N_5008,N_4425,N_4489);
nor U5009 (N_5009,N_4319,N_4690);
nor U5010 (N_5010,N_4367,N_4094);
or U5011 (N_5011,N_4035,N_4810);
nand U5012 (N_5012,N_4941,N_4910);
nor U5013 (N_5013,N_4046,N_4205);
and U5014 (N_5014,N_4541,N_4660);
nor U5015 (N_5015,N_4057,N_4861);
or U5016 (N_5016,N_4815,N_4918);
and U5017 (N_5017,N_4914,N_4392);
nor U5018 (N_5018,N_4354,N_4148);
or U5019 (N_5019,N_4729,N_4681);
and U5020 (N_5020,N_4475,N_4436);
or U5021 (N_5021,N_4024,N_4257);
xor U5022 (N_5022,N_4213,N_4041);
and U5023 (N_5023,N_4280,N_4323);
nor U5024 (N_5024,N_4445,N_4637);
and U5025 (N_5025,N_4357,N_4930);
and U5026 (N_5026,N_4740,N_4264);
and U5027 (N_5027,N_4977,N_4877);
nor U5028 (N_5028,N_4468,N_4347);
or U5029 (N_5029,N_4448,N_4242);
or U5030 (N_5030,N_4391,N_4162);
and U5031 (N_5031,N_4886,N_4145);
nor U5032 (N_5032,N_4752,N_4123);
and U5033 (N_5033,N_4458,N_4322);
or U5034 (N_5034,N_4568,N_4892);
nand U5035 (N_5035,N_4952,N_4888);
and U5036 (N_5036,N_4964,N_4827);
xor U5037 (N_5037,N_4498,N_4510);
nand U5038 (N_5038,N_4627,N_4653);
nand U5039 (N_5039,N_4420,N_4375);
nand U5040 (N_5040,N_4991,N_4485);
and U5041 (N_5041,N_4153,N_4151);
and U5042 (N_5042,N_4198,N_4271);
nand U5043 (N_5043,N_4460,N_4848);
or U5044 (N_5044,N_4048,N_4544);
and U5045 (N_5045,N_4782,N_4915);
nand U5046 (N_5046,N_4343,N_4206);
and U5047 (N_5047,N_4968,N_4352);
nor U5048 (N_5048,N_4350,N_4819);
nand U5049 (N_5049,N_4384,N_4454);
or U5050 (N_5050,N_4239,N_4300);
nand U5051 (N_5051,N_4452,N_4699);
xnor U5052 (N_5052,N_4766,N_4254);
xnor U5053 (N_5053,N_4382,N_4061);
nor U5054 (N_5054,N_4100,N_4756);
or U5055 (N_5055,N_4997,N_4502);
nand U5056 (N_5056,N_4386,N_4641);
and U5057 (N_5057,N_4763,N_4135);
and U5058 (N_5058,N_4836,N_4157);
or U5059 (N_5059,N_4528,N_4771);
or U5060 (N_5060,N_4349,N_4718);
and U5061 (N_5061,N_4530,N_4829);
nor U5062 (N_5062,N_4379,N_4484);
and U5063 (N_5063,N_4230,N_4809);
and U5064 (N_5064,N_4787,N_4291);
nand U5065 (N_5065,N_4253,N_4134);
and U5066 (N_5066,N_4029,N_4516);
nand U5067 (N_5067,N_4673,N_4825);
or U5068 (N_5068,N_4062,N_4000);
nor U5069 (N_5069,N_4372,N_4674);
nor U5070 (N_5070,N_4654,N_4723);
or U5071 (N_5071,N_4474,N_4579);
and U5072 (N_5072,N_4456,N_4422);
or U5073 (N_5073,N_4494,N_4665);
nand U5074 (N_5074,N_4947,N_4394);
or U5075 (N_5075,N_4181,N_4129);
xnor U5076 (N_5076,N_4446,N_4864);
and U5077 (N_5077,N_4549,N_4642);
nand U5078 (N_5078,N_4896,N_4019);
nand U5079 (N_5079,N_4767,N_4596);
nand U5080 (N_5080,N_4104,N_4328);
and U5081 (N_5081,N_4719,N_4635);
and U5082 (N_5082,N_4908,N_4734);
nor U5083 (N_5083,N_4138,N_4356);
nor U5084 (N_5084,N_4478,N_4417);
or U5085 (N_5085,N_4077,N_4262);
nor U5086 (N_5086,N_4389,N_4758);
or U5087 (N_5087,N_4017,N_4267);
nand U5088 (N_5088,N_4090,N_4192);
nand U5089 (N_5089,N_4305,N_4951);
nand U5090 (N_5090,N_4030,N_4649);
nand U5091 (N_5091,N_4508,N_4683);
nor U5092 (N_5092,N_4373,N_4402);
nor U5093 (N_5093,N_4353,N_4703);
or U5094 (N_5094,N_4221,N_4313);
nor U5095 (N_5095,N_4507,N_4677);
nand U5096 (N_5096,N_4950,N_4107);
and U5097 (N_5097,N_4419,N_4822);
and U5098 (N_5098,N_4139,N_4693);
or U5099 (N_5099,N_4571,N_4832);
nor U5100 (N_5100,N_4808,N_4376);
nand U5101 (N_5101,N_4237,N_4880);
and U5102 (N_5102,N_4633,N_4021);
or U5103 (N_5103,N_4937,N_4733);
or U5104 (N_5104,N_4773,N_4942);
nand U5105 (N_5105,N_4555,N_4894);
nand U5106 (N_5106,N_4140,N_4331);
xnor U5107 (N_5107,N_4272,N_4501);
nor U5108 (N_5108,N_4576,N_4973);
nor U5109 (N_5109,N_4444,N_4043);
nor U5110 (N_5110,N_4934,N_4797);
xor U5111 (N_5111,N_4016,N_4362);
or U5112 (N_5112,N_4482,N_4255);
nand U5113 (N_5113,N_4661,N_4757);
nor U5114 (N_5114,N_4847,N_4584);
or U5115 (N_5115,N_4039,N_4988);
and U5116 (N_5116,N_4212,N_4518);
and U5117 (N_5117,N_4390,N_4998);
nor U5118 (N_5118,N_4128,N_4190);
and U5119 (N_5119,N_4493,N_4383);
and U5120 (N_5120,N_4269,N_4109);
xor U5121 (N_5121,N_4177,N_4623);
nand U5122 (N_5122,N_4953,N_4089);
or U5123 (N_5123,N_4891,N_4595);
xnor U5124 (N_5124,N_4605,N_4286);
xor U5125 (N_5125,N_4005,N_4807);
and U5126 (N_5126,N_4462,N_4866);
and U5127 (N_5127,N_4900,N_4841);
xnor U5128 (N_5128,N_4435,N_4275);
and U5129 (N_5129,N_4209,N_4119);
nor U5130 (N_5130,N_4152,N_4545);
and U5131 (N_5131,N_4279,N_4053);
nor U5132 (N_5132,N_4059,N_4481);
nand U5133 (N_5133,N_4006,N_4058);
nand U5134 (N_5134,N_4725,N_4092);
or U5135 (N_5135,N_4688,N_4745);
or U5136 (N_5136,N_4408,N_4806);
or U5137 (N_5137,N_4141,N_4907);
xor U5138 (N_5138,N_4296,N_4614);
nand U5139 (N_5139,N_4547,N_4312);
or U5140 (N_5140,N_4543,N_4967);
nor U5141 (N_5141,N_4233,N_4936);
xor U5142 (N_5142,N_4285,N_4274);
nor U5143 (N_5143,N_4070,N_4290);
nor U5144 (N_5144,N_4054,N_4857);
and U5145 (N_5145,N_4015,N_4027);
or U5146 (N_5146,N_4929,N_4933);
or U5147 (N_5147,N_4479,N_4995);
nand U5148 (N_5148,N_4248,N_4049);
nand U5149 (N_5149,N_4122,N_4260);
nor U5150 (N_5150,N_4457,N_4166);
and U5151 (N_5151,N_4976,N_4803);
or U5152 (N_5152,N_4585,N_4890);
xor U5153 (N_5153,N_4040,N_4374);
xnor U5154 (N_5154,N_4440,N_4284);
or U5155 (N_5155,N_4193,N_4859);
nor U5156 (N_5156,N_4788,N_4429);
nor U5157 (N_5157,N_4158,N_4831);
nor U5158 (N_5158,N_4522,N_4939);
nor U5159 (N_5159,N_4324,N_4700);
nand U5160 (N_5160,N_4366,N_4339);
nand U5161 (N_5161,N_4603,N_4638);
xor U5162 (N_5162,N_4093,N_4833);
nand U5163 (N_5163,N_4423,N_4011);
nor U5164 (N_5164,N_4065,N_4755);
or U5165 (N_5165,N_4765,N_4852);
and U5166 (N_5166,N_4743,N_4293);
nand U5167 (N_5167,N_4762,N_4514);
nor U5168 (N_5168,N_4467,N_4567);
or U5169 (N_5169,N_4582,N_4801);
nand U5170 (N_5170,N_4091,N_4424);
and U5171 (N_5171,N_4033,N_4970);
or U5172 (N_5172,N_4639,N_4316);
and U5173 (N_5173,N_4117,N_4326);
and U5174 (N_5174,N_4625,N_4909);
or U5175 (N_5175,N_4946,N_4003);
and U5176 (N_5176,N_4685,N_4302);
or U5177 (N_5177,N_4956,N_4195);
nand U5178 (N_5178,N_4238,N_4668);
or U5179 (N_5179,N_4008,N_4670);
and U5180 (N_5180,N_4870,N_4464);
nand U5181 (N_5181,N_4586,N_4118);
and U5182 (N_5182,N_4110,N_4154);
or U5183 (N_5183,N_4728,N_4538);
or U5184 (N_5184,N_4051,N_4597);
or U5185 (N_5185,N_4520,N_4395);
nor U5186 (N_5186,N_4666,N_4304);
and U5187 (N_5187,N_4526,N_4266);
nor U5188 (N_5188,N_4747,N_4416);
and U5189 (N_5189,N_4557,N_4542);
and U5190 (N_5190,N_4984,N_4628);
and U5191 (N_5191,N_4176,N_4565);
and U5192 (N_5192,N_4958,N_4342);
and U5193 (N_5193,N_4632,N_4702);
nor U5194 (N_5194,N_4075,N_4731);
or U5195 (N_5195,N_4611,N_4959);
nor U5196 (N_5196,N_4405,N_4377);
nor U5197 (N_5197,N_4088,N_4472);
or U5198 (N_5198,N_4598,N_4564);
nor U5199 (N_5199,N_4449,N_4592);
and U5200 (N_5200,N_4931,N_4308);
and U5201 (N_5201,N_4513,N_4712);
nand U5202 (N_5202,N_4364,N_4009);
or U5203 (N_5203,N_4483,N_4790);
nand U5204 (N_5204,N_4330,N_4736);
or U5205 (N_5205,N_4981,N_4018);
and U5206 (N_5206,N_4295,N_4273);
nor U5207 (N_5207,N_4459,N_4903);
and U5208 (N_5208,N_4210,N_4980);
nor U5209 (N_5209,N_4706,N_4171);
xor U5210 (N_5210,N_4994,N_4669);
and U5211 (N_5211,N_4063,N_4846);
nand U5212 (N_5212,N_4341,N_4155);
nand U5213 (N_5213,N_4161,N_4160);
or U5214 (N_5214,N_4966,N_4969);
nand U5215 (N_5215,N_4218,N_4028);
nand U5216 (N_5216,N_4067,N_4183);
or U5217 (N_5217,N_4989,N_4471);
or U5218 (N_5218,N_4224,N_4816);
or U5219 (N_5219,N_4759,N_4412);
nand U5220 (N_5220,N_4663,N_4651);
and U5221 (N_5221,N_4684,N_4769);
or U5222 (N_5222,N_4270,N_4511);
nor U5223 (N_5223,N_4505,N_4780);
nand U5224 (N_5224,N_4486,N_4878);
nor U5225 (N_5225,N_4144,N_4671);
or U5226 (N_5226,N_4215,N_4175);
and U5227 (N_5227,N_4657,N_4996);
xor U5228 (N_5228,N_4113,N_4406);
xor U5229 (N_5229,N_4987,N_4199);
nand U5230 (N_5230,N_4811,N_4813);
or U5231 (N_5231,N_4231,N_4359);
or U5232 (N_5232,N_4850,N_4358);
nand U5233 (N_5233,N_4744,N_4414);
xnor U5234 (N_5234,N_4022,N_4536);
nand U5235 (N_5235,N_4537,N_4556);
nor U5236 (N_5236,N_4963,N_4561);
nand U5237 (N_5237,N_4678,N_4923);
nor U5238 (N_5238,N_4217,N_4949);
and U5239 (N_5239,N_4164,N_4524);
nand U5240 (N_5240,N_4147,N_4716);
nor U5241 (N_5241,N_4919,N_4796);
and U5242 (N_5242,N_4875,N_4034);
nor U5243 (N_5243,N_4791,N_4785);
nor U5244 (N_5244,N_4086,N_4036);
or U5245 (N_5245,N_4149,N_4361);
or U5246 (N_5246,N_4334,N_4052);
xnor U5247 (N_5247,N_4050,N_4108);
nand U5248 (N_5248,N_4717,N_4369);
xnor U5249 (N_5249,N_4512,N_4682);
and U5250 (N_5250,N_4243,N_4074);
or U5251 (N_5251,N_4979,N_4655);
nand U5252 (N_5252,N_4687,N_4944);
and U5253 (N_5253,N_4309,N_4509);
and U5254 (N_5254,N_4664,N_4594);
nor U5255 (N_5255,N_4187,N_4553);
xor U5256 (N_5256,N_4137,N_4658);
nor U5257 (N_5257,N_4698,N_4411);
or U5258 (N_5258,N_4012,N_4779);
and U5259 (N_5259,N_4609,N_4529);
or U5260 (N_5260,N_4225,N_4647);
xnor U5261 (N_5261,N_4120,N_4845);
nor U5262 (N_5262,N_4985,N_4403);
and U5263 (N_5263,N_4197,N_4283);
nor U5264 (N_5264,N_4245,N_4473);
xor U5265 (N_5265,N_4525,N_4306);
nand U5266 (N_5266,N_4125,N_4360);
xor U5267 (N_5267,N_4573,N_4645);
or U5268 (N_5268,N_4523,N_4563);
or U5269 (N_5269,N_4975,N_4962);
or U5270 (N_5270,N_4754,N_4532);
or U5271 (N_5271,N_4317,N_4868);
nor U5272 (N_5272,N_4708,N_4150);
nor U5273 (N_5273,N_4821,N_4060);
and U5274 (N_5274,N_4867,N_4901);
nor U5275 (N_5275,N_4805,N_4615);
and U5276 (N_5276,N_4593,N_4643);
xnor U5277 (N_5277,N_4202,N_4143);
nand U5278 (N_5278,N_4329,N_4607);
or U5279 (N_5279,N_4707,N_4581);
or U5280 (N_5280,N_4739,N_4726);
nor U5281 (N_5281,N_4083,N_4837);
nor U5282 (N_5282,N_4496,N_4616);
nor U5283 (N_5283,N_4772,N_4315);
or U5284 (N_5284,N_4672,N_4775);
or U5285 (N_5285,N_4619,N_4249);
and U5286 (N_5286,N_4082,N_4170);
and U5287 (N_5287,N_4168,N_4885);
or U5288 (N_5288,N_4802,N_4881);
or U5289 (N_5289,N_4131,N_4887);
or U5290 (N_5290,N_4325,N_4229);
xnor U5291 (N_5291,N_4826,N_4071);
or U5292 (N_5292,N_4746,N_4069);
nor U5293 (N_5293,N_4659,N_4400);
nor U5294 (N_5294,N_4078,N_4453);
nor U5295 (N_5295,N_4817,N_4132);
and U5296 (N_5296,N_4694,N_4727);
nand U5297 (N_5297,N_4679,N_4013);
or U5298 (N_5298,N_4159,N_4751);
nand U5299 (N_5299,N_4920,N_4142);
or U5300 (N_5300,N_4163,N_4534);
and U5301 (N_5301,N_4961,N_4853);
or U5302 (N_5302,N_4993,N_4842);
nor U5303 (N_5303,N_4889,N_4792);
or U5304 (N_5304,N_4748,N_4786);
and U5305 (N_5305,N_4550,N_4818);
nand U5306 (N_5306,N_4430,N_4025);
and U5307 (N_5307,N_4080,N_4252);
nor U5308 (N_5308,N_4872,N_4044);
or U5309 (N_5309,N_4007,N_4105);
or U5310 (N_5310,N_4957,N_4630);
nand U5311 (N_5311,N_4204,N_4574);
or U5312 (N_5312,N_4156,N_4413);
nor U5313 (N_5313,N_4207,N_4855);
or U5314 (N_5314,N_4259,N_4795);
nand U5315 (N_5315,N_4646,N_4421);
nand U5316 (N_5316,N_4636,N_4548);
or U5317 (N_5317,N_4720,N_4097);
nand U5318 (N_5318,N_4932,N_4240);
and U5319 (N_5319,N_4580,N_4469);
or U5320 (N_5320,N_4730,N_4776);
nor U5321 (N_5321,N_4004,N_4906);
nand U5322 (N_5322,N_4463,N_4102);
nand U5323 (N_5323,N_4711,N_4527);
nand U5324 (N_5324,N_4583,N_4999);
nand U5325 (N_5325,N_4814,N_4073);
nor U5326 (N_5326,N_4263,N_4201);
nor U5327 (N_5327,N_4432,N_4320);
xnor U5328 (N_5328,N_4506,N_4223);
or U5329 (N_5329,N_4455,N_4447);
xnor U5330 (N_5330,N_4539,N_4297);
or U5331 (N_5331,N_4960,N_4227);
nand U5332 (N_5332,N_4954,N_4606);
or U5333 (N_5333,N_4799,N_4351);
and U5334 (N_5334,N_4774,N_4431);
nand U5335 (N_5335,N_4492,N_4644);
or U5336 (N_5336,N_4363,N_4345);
xnor U5337 (N_5337,N_4823,N_4656);
and U5338 (N_5338,N_4184,N_4121);
nor U5339 (N_5339,N_4883,N_4874);
or U5340 (N_5340,N_4926,N_4610);
or U5341 (N_5341,N_4335,N_4172);
xor U5342 (N_5342,N_4236,N_4869);
xor U5343 (N_5343,N_4076,N_4495);
or U5344 (N_5344,N_4401,N_4618);
xnor U5345 (N_5345,N_4631,N_4904);
or U5346 (N_5346,N_4470,N_4935);
and U5347 (N_5347,N_4333,N_4265);
or U5348 (N_5348,N_4045,N_4517);
nand U5349 (N_5349,N_4348,N_4114);
or U5350 (N_5350,N_4650,N_4126);
nand U5351 (N_5351,N_4124,N_4268);
nand U5352 (N_5352,N_4844,N_4955);
or U5353 (N_5353,N_4047,N_4340);
and U5354 (N_5354,N_4174,N_4294);
nand U5355 (N_5355,N_4697,N_4781);
and U5356 (N_5356,N_4222,N_4552);
and U5357 (N_5357,N_4972,N_4715);
or U5358 (N_5358,N_4566,N_4261);
and U5359 (N_5359,N_4096,N_4519);
nand U5360 (N_5360,N_4393,N_4146);
and U5361 (N_5361,N_4032,N_4188);
xor U5362 (N_5362,N_4476,N_4912);
xor U5363 (N_5363,N_4241,N_4741);
or U5364 (N_5364,N_4721,N_4691);
and U5365 (N_5365,N_4234,N_4895);
nor U5366 (N_5366,N_4570,N_4127);
or U5367 (N_5367,N_4365,N_4608);
xnor U5368 (N_5368,N_4680,N_4397);
and U5369 (N_5369,N_4838,N_4443);
nand U5370 (N_5370,N_4042,N_4208);
or U5371 (N_5371,N_4064,N_4577);
nand U5372 (N_5372,N_4794,N_4327);
nor U5373 (N_5373,N_4913,N_4368);
and U5374 (N_5374,N_4676,N_4292);
or U5375 (N_5375,N_4344,N_4336);
and U5376 (N_5376,N_4737,N_4800);
xor U5377 (N_5377,N_4925,N_4084);
and U5378 (N_5378,N_4020,N_4735);
or U5379 (N_5379,N_4111,N_4893);
xnor U5380 (N_5380,N_4856,N_4732);
nand U5381 (N_5381,N_4418,N_4865);
nand U5382 (N_5382,N_4281,N_4196);
and U5383 (N_5383,N_4399,N_4098);
or U5384 (N_5384,N_4318,N_4169);
or U5385 (N_5385,N_4983,N_4165);
nand U5386 (N_5386,N_4251,N_4115);
nand U5387 (N_5387,N_4338,N_4216);
and U5388 (N_5388,N_4879,N_4497);
or U5389 (N_5389,N_4228,N_4554);
xnor U5390 (N_5390,N_4648,N_4873);
nand U5391 (N_5391,N_4437,N_4037);
and U5392 (N_5392,N_4804,N_4332);
nand U5393 (N_5393,N_4928,N_4396);
or U5394 (N_5394,N_4640,N_4533);
or U5395 (N_5395,N_4346,N_4710);
nor U5396 (N_5396,N_4531,N_4371);
nand U5397 (N_5397,N_4590,N_4990);
and U5398 (N_5398,N_4897,N_4173);
nor U5399 (N_5399,N_4095,N_4535);
and U5400 (N_5400,N_4905,N_4789);
nand U5401 (N_5401,N_4311,N_4499);
or U5402 (N_5402,N_4834,N_4310);
nand U5403 (N_5403,N_4480,N_4974);
nand U5404 (N_5404,N_4770,N_4858);
nor U5405 (N_5405,N_4835,N_4922);
xnor U5406 (N_5406,N_4849,N_4085);
and U5407 (N_5407,N_4410,N_4917);
or U5408 (N_5408,N_4911,N_4103);
nor U5409 (N_5409,N_4938,N_4387);
or U5410 (N_5410,N_4546,N_4200);
nor U5411 (N_5411,N_4023,N_4258);
nor U5412 (N_5412,N_4578,N_4840);
nor U5413 (N_5413,N_4948,N_4136);
nand U5414 (N_5414,N_4830,N_4714);
xnor U5415 (N_5415,N_4812,N_4876);
or U5416 (N_5416,N_4713,N_4978);
nor U5417 (N_5417,N_4288,N_4378);
nor U5418 (N_5418,N_4589,N_4451);
nor U5419 (N_5419,N_4899,N_4971);
and U5420 (N_5420,N_4705,N_4385);
nor U5421 (N_5421,N_4066,N_4784);
nand U5422 (N_5422,N_4986,N_4398);
and U5423 (N_5423,N_4185,N_4575);
or U5424 (N_5424,N_4101,N_4246);
nor U5425 (N_5425,N_4001,N_4180);
or U5426 (N_5426,N_4178,N_4862);
nand U5427 (N_5427,N_4355,N_4982);
nor U5428 (N_5428,N_4600,N_4031);
nor U5429 (N_5429,N_4587,N_4220);
and U5430 (N_5430,N_4613,N_4612);
xnor U5431 (N_5431,N_4843,N_4675);
nor U5432 (N_5432,N_4450,N_4521);
and U5433 (N_5433,N_4232,N_4760);
or U5434 (N_5434,N_4871,N_4186);
or U5435 (N_5435,N_4388,N_4667);
nand U5436 (N_5436,N_4056,N_4409);
and U5437 (N_5437,N_4828,N_4704);
and U5438 (N_5438,N_4851,N_4839);
or U5439 (N_5439,N_4287,N_4277);
nand U5440 (N_5440,N_4884,N_4860);
and U5441 (N_5441,N_4010,N_4824);
nand U5442 (N_5442,N_4079,N_4407);
or U5443 (N_5443,N_4965,N_4442);
nor U5444 (N_5444,N_4695,N_4924);
nand U5445 (N_5445,N_4191,N_4301);
xnor U5446 (N_5446,N_4298,N_4491);
or U5447 (N_5447,N_4182,N_4380);
and U5448 (N_5448,N_4055,N_4307);
and U5449 (N_5449,N_4211,N_4686);
nor U5450 (N_5450,N_4572,N_4167);
and U5451 (N_5451,N_4465,N_4370);
and U5452 (N_5452,N_4854,N_4189);
and U5453 (N_5453,N_4662,N_4219);
and U5454 (N_5454,N_4038,N_4902);
and U5455 (N_5455,N_4601,N_4898);
nand U5456 (N_5456,N_4337,N_4087);
nand U5457 (N_5457,N_4943,N_4116);
or U5458 (N_5458,N_4433,N_4133);
nand U5459 (N_5459,N_4194,N_4130);
nor U5460 (N_5460,N_4753,N_4321);
or U5461 (N_5461,N_4783,N_4689);
nand U5462 (N_5462,N_4404,N_4768);
xnor U5463 (N_5463,N_4504,N_4303);
nand U5464 (N_5464,N_4461,N_4652);
nor U5465 (N_5465,N_4428,N_4014);
and U5466 (N_5466,N_4434,N_4798);
and U5467 (N_5467,N_4738,N_4558);
and U5468 (N_5468,N_4620,N_4621);
or U5469 (N_5469,N_4381,N_4278);
and U5470 (N_5470,N_4750,N_4927);
nand U5471 (N_5471,N_4560,N_4477);
nand U5472 (N_5472,N_4099,N_4599);
xor U5473 (N_5473,N_4438,N_4226);
and U5474 (N_5474,N_4515,N_4276);
or U5475 (N_5475,N_4820,N_4256);
or U5476 (N_5476,N_4622,N_4441);
and U5477 (N_5477,N_4214,N_4466);
and U5478 (N_5478,N_4921,N_4427);
and U5479 (N_5479,N_4764,N_4749);
nor U5480 (N_5480,N_4244,N_4569);
and U5481 (N_5481,N_4106,N_4945);
nand U5482 (N_5482,N_4701,N_4863);
or U5483 (N_5483,N_4026,N_4439);
nor U5484 (N_5484,N_4068,N_4503);
nor U5485 (N_5485,N_4415,N_4591);
or U5486 (N_5486,N_4247,N_4696);
nand U5487 (N_5487,N_4559,N_4112);
nand U5488 (N_5488,N_4916,N_4709);
nand U5489 (N_5489,N_4940,N_4882);
nand U5490 (N_5490,N_4742,N_4487);
nand U5491 (N_5491,N_4624,N_4289);
nor U5492 (N_5492,N_4299,N_4235);
nor U5493 (N_5493,N_4179,N_4203);
and U5494 (N_5494,N_4692,N_4602);
or U5495 (N_5495,N_4793,N_4072);
or U5496 (N_5496,N_4629,N_4588);
nand U5497 (N_5497,N_4992,N_4002);
nor U5498 (N_5498,N_4722,N_4282);
and U5499 (N_5499,N_4314,N_4250);
nand U5500 (N_5500,N_4515,N_4230);
nand U5501 (N_5501,N_4859,N_4922);
nand U5502 (N_5502,N_4890,N_4434);
nor U5503 (N_5503,N_4310,N_4743);
nor U5504 (N_5504,N_4410,N_4079);
and U5505 (N_5505,N_4268,N_4797);
nor U5506 (N_5506,N_4907,N_4304);
or U5507 (N_5507,N_4850,N_4774);
or U5508 (N_5508,N_4373,N_4600);
nand U5509 (N_5509,N_4088,N_4864);
nand U5510 (N_5510,N_4876,N_4544);
or U5511 (N_5511,N_4683,N_4254);
nor U5512 (N_5512,N_4636,N_4856);
nand U5513 (N_5513,N_4915,N_4602);
and U5514 (N_5514,N_4217,N_4359);
nor U5515 (N_5515,N_4451,N_4397);
and U5516 (N_5516,N_4787,N_4646);
nor U5517 (N_5517,N_4751,N_4310);
or U5518 (N_5518,N_4537,N_4718);
nor U5519 (N_5519,N_4821,N_4308);
nand U5520 (N_5520,N_4718,N_4860);
nor U5521 (N_5521,N_4994,N_4573);
nand U5522 (N_5522,N_4247,N_4222);
nor U5523 (N_5523,N_4746,N_4976);
nand U5524 (N_5524,N_4659,N_4198);
and U5525 (N_5525,N_4730,N_4609);
or U5526 (N_5526,N_4003,N_4951);
or U5527 (N_5527,N_4864,N_4121);
nor U5528 (N_5528,N_4987,N_4298);
nor U5529 (N_5529,N_4777,N_4058);
nor U5530 (N_5530,N_4118,N_4366);
or U5531 (N_5531,N_4490,N_4451);
or U5532 (N_5532,N_4863,N_4028);
or U5533 (N_5533,N_4112,N_4817);
or U5534 (N_5534,N_4519,N_4280);
or U5535 (N_5535,N_4142,N_4295);
nand U5536 (N_5536,N_4456,N_4860);
and U5537 (N_5537,N_4481,N_4121);
nand U5538 (N_5538,N_4022,N_4365);
and U5539 (N_5539,N_4223,N_4211);
or U5540 (N_5540,N_4541,N_4832);
or U5541 (N_5541,N_4435,N_4013);
or U5542 (N_5542,N_4043,N_4395);
and U5543 (N_5543,N_4453,N_4398);
nand U5544 (N_5544,N_4232,N_4632);
and U5545 (N_5545,N_4271,N_4154);
nor U5546 (N_5546,N_4353,N_4112);
xnor U5547 (N_5547,N_4293,N_4970);
xnor U5548 (N_5548,N_4477,N_4005);
and U5549 (N_5549,N_4566,N_4033);
nor U5550 (N_5550,N_4234,N_4883);
nand U5551 (N_5551,N_4485,N_4696);
and U5552 (N_5552,N_4302,N_4786);
nor U5553 (N_5553,N_4481,N_4334);
nand U5554 (N_5554,N_4248,N_4784);
or U5555 (N_5555,N_4292,N_4766);
xnor U5556 (N_5556,N_4161,N_4249);
nor U5557 (N_5557,N_4482,N_4981);
nand U5558 (N_5558,N_4300,N_4551);
or U5559 (N_5559,N_4563,N_4307);
or U5560 (N_5560,N_4747,N_4787);
and U5561 (N_5561,N_4265,N_4812);
xor U5562 (N_5562,N_4016,N_4506);
nand U5563 (N_5563,N_4602,N_4753);
and U5564 (N_5564,N_4997,N_4115);
and U5565 (N_5565,N_4009,N_4826);
and U5566 (N_5566,N_4515,N_4648);
nor U5567 (N_5567,N_4510,N_4631);
nor U5568 (N_5568,N_4351,N_4122);
or U5569 (N_5569,N_4855,N_4409);
or U5570 (N_5570,N_4207,N_4943);
nor U5571 (N_5571,N_4480,N_4444);
or U5572 (N_5572,N_4742,N_4270);
nand U5573 (N_5573,N_4030,N_4783);
xnor U5574 (N_5574,N_4002,N_4192);
nor U5575 (N_5575,N_4077,N_4110);
or U5576 (N_5576,N_4750,N_4374);
or U5577 (N_5577,N_4697,N_4174);
and U5578 (N_5578,N_4982,N_4528);
nand U5579 (N_5579,N_4038,N_4026);
nor U5580 (N_5580,N_4049,N_4983);
xnor U5581 (N_5581,N_4387,N_4996);
nand U5582 (N_5582,N_4013,N_4911);
nand U5583 (N_5583,N_4737,N_4994);
nand U5584 (N_5584,N_4486,N_4079);
or U5585 (N_5585,N_4324,N_4217);
or U5586 (N_5586,N_4656,N_4248);
or U5587 (N_5587,N_4576,N_4624);
xnor U5588 (N_5588,N_4805,N_4171);
or U5589 (N_5589,N_4836,N_4777);
xor U5590 (N_5590,N_4578,N_4964);
nor U5591 (N_5591,N_4387,N_4490);
or U5592 (N_5592,N_4824,N_4970);
or U5593 (N_5593,N_4637,N_4295);
or U5594 (N_5594,N_4347,N_4761);
or U5595 (N_5595,N_4501,N_4224);
nand U5596 (N_5596,N_4145,N_4934);
or U5597 (N_5597,N_4277,N_4071);
or U5598 (N_5598,N_4154,N_4601);
nor U5599 (N_5599,N_4518,N_4444);
nor U5600 (N_5600,N_4678,N_4854);
xor U5601 (N_5601,N_4697,N_4299);
or U5602 (N_5602,N_4944,N_4234);
nor U5603 (N_5603,N_4161,N_4239);
and U5604 (N_5604,N_4652,N_4842);
or U5605 (N_5605,N_4742,N_4496);
nand U5606 (N_5606,N_4754,N_4042);
nor U5607 (N_5607,N_4859,N_4703);
and U5608 (N_5608,N_4872,N_4485);
or U5609 (N_5609,N_4308,N_4512);
nor U5610 (N_5610,N_4771,N_4167);
and U5611 (N_5611,N_4649,N_4467);
nand U5612 (N_5612,N_4843,N_4124);
nor U5613 (N_5613,N_4137,N_4038);
or U5614 (N_5614,N_4072,N_4103);
and U5615 (N_5615,N_4765,N_4456);
nand U5616 (N_5616,N_4537,N_4452);
nand U5617 (N_5617,N_4779,N_4643);
nor U5618 (N_5618,N_4207,N_4382);
and U5619 (N_5619,N_4488,N_4388);
or U5620 (N_5620,N_4147,N_4877);
and U5621 (N_5621,N_4669,N_4085);
or U5622 (N_5622,N_4645,N_4295);
and U5623 (N_5623,N_4379,N_4296);
nand U5624 (N_5624,N_4168,N_4171);
nor U5625 (N_5625,N_4404,N_4876);
nand U5626 (N_5626,N_4328,N_4585);
or U5627 (N_5627,N_4244,N_4820);
and U5628 (N_5628,N_4514,N_4027);
or U5629 (N_5629,N_4217,N_4246);
nand U5630 (N_5630,N_4840,N_4178);
or U5631 (N_5631,N_4440,N_4066);
nor U5632 (N_5632,N_4491,N_4151);
and U5633 (N_5633,N_4773,N_4379);
or U5634 (N_5634,N_4685,N_4347);
xnor U5635 (N_5635,N_4527,N_4649);
nand U5636 (N_5636,N_4075,N_4063);
nand U5637 (N_5637,N_4479,N_4371);
nor U5638 (N_5638,N_4413,N_4279);
nor U5639 (N_5639,N_4061,N_4632);
nand U5640 (N_5640,N_4279,N_4072);
and U5641 (N_5641,N_4015,N_4716);
nor U5642 (N_5642,N_4576,N_4783);
or U5643 (N_5643,N_4488,N_4781);
and U5644 (N_5644,N_4654,N_4514);
or U5645 (N_5645,N_4399,N_4804);
nor U5646 (N_5646,N_4323,N_4185);
or U5647 (N_5647,N_4256,N_4057);
xnor U5648 (N_5648,N_4556,N_4646);
nand U5649 (N_5649,N_4171,N_4895);
or U5650 (N_5650,N_4522,N_4314);
xnor U5651 (N_5651,N_4434,N_4648);
nor U5652 (N_5652,N_4549,N_4350);
nand U5653 (N_5653,N_4124,N_4530);
nor U5654 (N_5654,N_4210,N_4365);
nor U5655 (N_5655,N_4039,N_4715);
or U5656 (N_5656,N_4287,N_4756);
and U5657 (N_5657,N_4591,N_4537);
and U5658 (N_5658,N_4277,N_4497);
nor U5659 (N_5659,N_4646,N_4893);
nor U5660 (N_5660,N_4312,N_4346);
xor U5661 (N_5661,N_4489,N_4471);
nand U5662 (N_5662,N_4502,N_4879);
and U5663 (N_5663,N_4543,N_4304);
nor U5664 (N_5664,N_4144,N_4095);
and U5665 (N_5665,N_4699,N_4657);
nand U5666 (N_5666,N_4520,N_4458);
nor U5667 (N_5667,N_4567,N_4766);
or U5668 (N_5668,N_4289,N_4385);
nand U5669 (N_5669,N_4861,N_4130);
nor U5670 (N_5670,N_4488,N_4430);
nand U5671 (N_5671,N_4579,N_4807);
or U5672 (N_5672,N_4205,N_4487);
nor U5673 (N_5673,N_4621,N_4865);
or U5674 (N_5674,N_4756,N_4945);
xor U5675 (N_5675,N_4776,N_4813);
nor U5676 (N_5676,N_4273,N_4057);
nor U5677 (N_5677,N_4330,N_4632);
nand U5678 (N_5678,N_4328,N_4919);
and U5679 (N_5679,N_4478,N_4751);
or U5680 (N_5680,N_4019,N_4298);
nor U5681 (N_5681,N_4242,N_4488);
xnor U5682 (N_5682,N_4272,N_4880);
xor U5683 (N_5683,N_4256,N_4060);
and U5684 (N_5684,N_4661,N_4886);
xor U5685 (N_5685,N_4187,N_4953);
nor U5686 (N_5686,N_4643,N_4609);
xnor U5687 (N_5687,N_4052,N_4516);
and U5688 (N_5688,N_4291,N_4391);
or U5689 (N_5689,N_4462,N_4080);
and U5690 (N_5690,N_4889,N_4882);
or U5691 (N_5691,N_4611,N_4341);
or U5692 (N_5692,N_4968,N_4481);
or U5693 (N_5693,N_4491,N_4260);
nor U5694 (N_5694,N_4531,N_4145);
xnor U5695 (N_5695,N_4895,N_4533);
xor U5696 (N_5696,N_4211,N_4975);
nor U5697 (N_5697,N_4730,N_4326);
nand U5698 (N_5698,N_4573,N_4476);
nor U5699 (N_5699,N_4379,N_4830);
nand U5700 (N_5700,N_4785,N_4506);
or U5701 (N_5701,N_4583,N_4211);
nor U5702 (N_5702,N_4318,N_4070);
and U5703 (N_5703,N_4018,N_4594);
and U5704 (N_5704,N_4583,N_4036);
nor U5705 (N_5705,N_4340,N_4847);
xor U5706 (N_5706,N_4150,N_4480);
nor U5707 (N_5707,N_4554,N_4112);
or U5708 (N_5708,N_4146,N_4770);
nand U5709 (N_5709,N_4883,N_4107);
nand U5710 (N_5710,N_4954,N_4958);
or U5711 (N_5711,N_4653,N_4696);
xnor U5712 (N_5712,N_4924,N_4469);
nand U5713 (N_5713,N_4513,N_4141);
nand U5714 (N_5714,N_4759,N_4196);
nand U5715 (N_5715,N_4685,N_4415);
nor U5716 (N_5716,N_4440,N_4074);
or U5717 (N_5717,N_4618,N_4599);
nor U5718 (N_5718,N_4888,N_4463);
and U5719 (N_5719,N_4304,N_4908);
nand U5720 (N_5720,N_4108,N_4915);
nand U5721 (N_5721,N_4014,N_4415);
nor U5722 (N_5722,N_4241,N_4726);
nand U5723 (N_5723,N_4577,N_4852);
nor U5724 (N_5724,N_4072,N_4308);
and U5725 (N_5725,N_4691,N_4270);
nor U5726 (N_5726,N_4912,N_4954);
nor U5727 (N_5727,N_4167,N_4071);
or U5728 (N_5728,N_4158,N_4601);
nand U5729 (N_5729,N_4033,N_4895);
or U5730 (N_5730,N_4259,N_4122);
or U5731 (N_5731,N_4909,N_4922);
and U5732 (N_5732,N_4018,N_4663);
or U5733 (N_5733,N_4510,N_4419);
and U5734 (N_5734,N_4180,N_4208);
nor U5735 (N_5735,N_4047,N_4011);
and U5736 (N_5736,N_4364,N_4321);
nor U5737 (N_5737,N_4038,N_4016);
xnor U5738 (N_5738,N_4706,N_4531);
nand U5739 (N_5739,N_4587,N_4710);
nand U5740 (N_5740,N_4303,N_4339);
nand U5741 (N_5741,N_4502,N_4742);
and U5742 (N_5742,N_4061,N_4401);
or U5743 (N_5743,N_4824,N_4335);
nand U5744 (N_5744,N_4146,N_4853);
xor U5745 (N_5745,N_4659,N_4920);
or U5746 (N_5746,N_4681,N_4694);
xor U5747 (N_5747,N_4273,N_4689);
nand U5748 (N_5748,N_4628,N_4798);
nor U5749 (N_5749,N_4419,N_4128);
nand U5750 (N_5750,N_4338,N_4559);
nor U5751 (N_5751,N_4853,N_4244);
nor U5752 (N_5752,N_4949,N_4931);
or U5753 (N_5753,N_4969,N_4249);
nor U5754 (N_5754,N_4686,N_4046);
nand U5755 (N_5755,N_4392,N_4780);
nand U5756 (N_5756,N_4796,N_4086);
or U5757 (N_5757,N_4821,N_4707);
or U5758 (N_5758,N_4175,N_4803);
or U5759 (N_5759,N_4398,N_4868);
or U5760 (N_5760,N_4670,N_4761);
nor U5761 (N_5761,N_4117,N_4321);
and U5762 (N_5762,N_4532,N_4579);
nor U5763 (N_5763,N_4572,N_4660);
nor U5764 (N_5764,N_4771,N_4704);
nor U5765 (N_5765,N_4398,N_4580);
xor U5766 (N_5766,N_4952,N_4050);
and U5767 (N_5767,N_4124,N_4468);
or U5768 (N_5768,N_4062,N_4024);
nand U5769 (N_5769,N_4304,N_4164);
or U5770 (N_5770,N_4670,N_4574);
nor U5771 (N_5771,N_4629,N_4549);
nand U5772 (N_5772,N_4773,N_4516);
nand U5773 (N_5773,N_4567,N_4027);
xor U5774 (N_5774,N_4696,N_4548);
and U5775 (N_5775,N_4591,N_4503);
and U5776 (N_5776,N_4079,N_4219);
nand U5777 (N_5777,N_4735,N_4488);
or U5778 (N_5778,N_4311,N_4664);
nor U5779 (N_5779,N_4122,N_4091);
and U5780 (N_5780,N_4896,N_4362);
and U5781 (N_5781,N_4567,N_4561);
nand U5782 (N_5782,N_4150,N_4449);
nand U5783 (N_5783,N_4923,N_4279);
nand U5784 (N_5784,N_4049,N_4763);
or U5785 (N_5785,N_4185,N_4828);
or U5786 (N_5786,N_4576,N_4842);
nand U5787 (N_5787,N_4788,N_4756);
nor U5788 (N_5788,N_4116,N_4810);
nor U5789 (N_5789,N_4758,N_4586);
nand U5790 (N_5790,N_4982,N_4004);
nor U5791 (N_5791,N_4236,N_4593);
or U5792 (N_5792,N_4475,N_4336);
nand U5793 (N_5793,N_4958,N_4411);
nand U5794 (N_5794,N_4581,N_4745);
or U5795 (N_5795,N_4349,N_4101);
nor U5796 (N_5796,N_4613,N_4751);
or U5797 (N_5797,N_4216,N_4782);
nand U5798 (N_5798,N_4419,N_4211);
nor U5799 (N_5799,N_4668,N_4750);
nand U5800 (N_5800,N_4665,N_4935);
or U5801 (N_5801,N_4938,N_4631);
nand U5802 (N_5802,N_4670,N_4623);
and U5803 (N_5803,N_4401,N_4045);
and U5804 (N_5804,N_4289,N_4295);
nand U5805 (N_5805,N_4207,N_4292);
nor U5806 (N_5806,N_4296,N_4500);
xnor U5807 (N_5807,N_4567,N_4476);
nor U5808 (N_5808,N_4813,N_4291);
and U5809 (N_5809,N_4570,N_4245);
nor U5810 (N_5810,N_4925,N_4394);
or U5811 (N_5811,N_4017,N_4282);
and U5812 (N_5812,N_4372,N_4696);
nor U5813 (N_5813,N_4183,N_4874);
or U5814 (N_5814,N_4468,N_4407);
xnor U5815 (N_5815,N_4844,N_4279);
and U5816 (N_5816,N_4336,N_4263);
and U5817 (N_5817,N_4581,N_4454);
or U5818 (N_5818,N_4716,N_4936);
and U5819 (N_5819,N_4570,N_4463);
and U5820 (N_5820,N_4309,N_4226);
or U5821 (N_5821,N_4008,N_4575);
and U5822 (N_5822,N_4732,N_4742);
or U5823 (N_5823,N_4828,N_4878);
or U5824 (N_5824,N_4473,N_4484);
nand U5825 (N_5825,N_4113,N_4498);
nand U5826 (N_5826,N_4918,N_4310);
nand U5827 (N_5827,N_4793,N_4170);
nor U5828 (N_5828,N_4062,N_4800);
and U5829 (N_5829,N_4074,N_4371);
nor U5830 (N_5830,N_4778,N_4566);
or U5831 (N_5831,N_4352,N_4299);
nor U5832 (N_5832,N_4468,N_4098);
nand U5833 (N_5833,N_4965,N_4945);
nor U5834 (N_5834,N_4818,N_4359);
nand U5835 (N_5835,N_4914,N_4345);
nand U5836 (N_5836,N_4446,N_4357);
and U5837 (N_5837,N_4248,N_4787);
and U5838 (N_5838,N_4566,N_4678);
or U5839 (N_5839,N_4478,N_4112);
nor U5840 (N_5840,N_4417,N_4223);
or U5841 (N_5841,N_4117,N_4992);
nand U5842 (N_5842,N_4033,N_4208);
or U5843 (N_5843,N_4678,N_4499);
nor U5844 (N_5844,N_4972,N_4273);
and U5845 (N_5845,N_4702,N_4914);
or U5846 (N_5846,N_4827,N_4414);
nor U5847 (N_5847,N_4827,N_4240);
nand U5848 (N_5848,N_4729,N_4085);
xor U5849 (N_5849,N_4545,N_4109);
nor U5850 (N_5850,N_4247,N_4173);
and U5851 (N_5851,N_4537,N_4894);
nor U5852 (N_5852,N_4543,N_4020);
or U5853 (N_5853,N_4774,N_4891);
and U5854 (N_5854,N_4876,N_4390);
or U5855 (N_5855,N_4978,N_4430);
and U5856 (N_5856,N_4419,N_4682);
or U5857 (N_5857,N_4740,N_4039);
nor U5858 (N_5858,N_4529,N_4901);
or U5859 (N_5859,N_4027,N_4804);
nand U5860 (N_5860,N_4495,N_4873);
and U5861 (N_5861,N_4762,N_4682);
nand U5862 (N_5862,N_4642,N_4161);
nor U5863 (N_5863,N_4372,N_4494);
xnor U5864 (N_5864,N_4355,N_4230);
and U5865 (N_5865,N_4867,N_4263);
nand U5866 (N_5866,N_4622,N_4090);
nor U5867 (N_5867,N_4932,N_4754);
or U5868 (N_5868,N_4878,N_4935);
nor U5869 (N_5869,N_4457,N_4263);
and U5870 (N_5870,N_4684,N_4353);
and U5871 (N_5871,N_4666,N_4675);
and U5872 (N_5872,N_4485,N_4296);
nand U5873 (N_5873,N_4700,N_4167);
and U5874 (N_5874,N_4576,N_4127);
or U5875 (N_5875,N_4912,N_4259);
nor U5876 (N_5876,N_4847,N_4199);
and U5877 (N_5877,N_4074,N_4730);
or U5878 (N_5878,N_4650,N_4545);
or U5879 (N_5879,N_4502,N_4775);
nand U5880 (N_5880,N_4192,N_4716);
and U5881 (N_5881,N_4631,N_4157);
nor U5882 (N_5882,N_4097,N_4939);
or U5883 (N_5883,N_4532,N_4935);
or U5884 (N_5884,N_4165,N_4910);
nor U5885 (N_5885,N_4382,N_4558);
xnor U5886 (N_5886,N_4132,N_4398);
nor U5887 (N_5887,N_4196,N_4216);
xor U5888 (N_5888,N_4000,N_4754);
and U5889 (N_5889,N_4913,N_4173);
and U5890 (N_5890,N_4804,N_4916);
and U5891 (N_5891,N_4377,N_4440);
or U5892 (N_5892,N_4328,N_4776);
or U5893 (N_5893,N_4270,N_4413);
nor U5894 (N_5894,N_4753,N_4229);
xor U5895 (N_5895,N_4803,N_4189);
or U5896 (N_5896,N_4284,N_4072);
nor U5897 (N_5897,N_4046,N_4245);
and U5898 (N_5898,N_4228,N_4971);
nand U5899 (N_5899,N_4036,N_4289);
or U5900 (N_5900,N_4309,N_4573);
xnor U5901 (N_5901,N_4530,N_4669);
nor U5902 (N_5902,N_4318,N_4231);
nand U5903 (N_5903,N_4093,N_4994);
or U5904 (N_5904,N_4417,N_4438);
and U5905 (N_5905,N_4704,N_4659);
nand U5906 (N_5906,N_4172,N_4117);
or U5907 (N_5907,N_4860,N_4553);
or U5908 (N_5908,N_4079,N_4635);
nor U5909 (N_5909,N_4250,N_4957);
or U5910 (N_5910,N_4389,N_4718);
or U5911 (N_5911,N_4650,N_4119);
and U5912 (N_5912,N_4304,N_4982);
nand U5913 (N_5913,N_4477,N_4693);
nor U5914 (N_5914,N_4664,N_4292);
xnor U5915 (N_5915,N_4249,N_4384);
nor U5916 (N_5916,N_4152,N_4007);
and U5917 (N_5917,N_4074,N_4332);
nand U5918 (N_5918,N_4399,N_4663);
or U5919 (N_5919,N_4824,N_4290);
nor U5920 (N_5920,N_4928,N_4652);
xnor U5921 (N_5921,N_4622,N_4123);
or U5922 (N_5922,N_4719,N_4055);
xnor U5923 (N_5923,N_4316,N_4127);
or U5924 (N_5924,N_4264,N_4589);
or U5925 (N_5925,N_4535,N_4892);
xor U5926 (N_5926,N_4176,N_4384);
or U5927 (N_5927,N_4685,N_4093);
nor U5928 (N_5928,N_4423,N_4667);
and U5929 (N_5929,N_4374,N_4623);
nand U5930 (N_5930,N_4997,N_4833);
nand U5931 (N_5931,N_4863,N_4886);
and U5932 (N_5932,N_4042,N_4511);
nor U5933 (N_5933,N_4422,N_4486);
nand U5934 (N_5934,N_4979,N_4958);
and U5935 (N_5935,N_4970,N_4088);
or U5936 (N_5936,N_4532,N_4247);
xor U5937 (N_5937,N_4111,N_4190);
nor U5938 (N_5938,N_4499,N_4078);
and U5939 (N_5939,N_4388,N_4381);
or U5940 (N_5940,N_4506,N_4397);
and U5941 (N_5941,N_4702,N_4813);
nand U5942 (N_5942,N_4892,N_4043);
and U5943 (N_5943,N_4576,N_4723);
nor U5944 (N_5944,N_4876,N_4207);
and U5945 (N_5945,N_4769,N_4115);
xor U5946 (N_5946,N_4062,N_4811);
and U5947 (N_5947,N_4244,N_4484);
nand U5948 (N_5948,N_4641,N_4266);
nor U5949 (N_5949,N_4577,N_4181);
or U5950 (N_5950,N_4759,N_4301);
nor U5951 (N_5951,N_4398,N_4973);
and U5952 (N_5952,N_4393,N_4331);
nor U5953 (N_5953,N_4164,N_4165);
nor U5954 (N_5954,N_4654,N_4589);
and U5955 (N_5955,N_4280,N_4007);
nand U5956 (N_5956,N_4256,N_4223);
nand U5957 (N_5957,N_4182,N_4771);
nand U5958 (N_5958,N_4558,N_4288);
or U5959 (N_5959,N_4215,N_4665);
nand U5960 (N_5960,N_4943,N_4440);
or U5961 (N_5961,N_4205,N_4740);
nor U5962 (N_5962,N_4194,N_4956);
nor U5963 (N_5963,N_4277,N_4840);
or U5964 (N_5964,N_4601,N_4909);
or U5965 (N_5965,N_4533,N_4718);
and U5966 (N_5966,N_4724,N_4648);
nand U5967 (N_5967,N_4284,N_4136);
nand U5968 (N_5968,N_4056,N_4960);
and U5969 (N_5969,N_4466,N_4008);
nand U5970 (N_5970,N_4558,N_4124);
nor U5971 (N_5971,N_4055,N_4005);
nor U5972 (N_5972,N_4441,N_4425);
nor U5973 (N_5973,N_4159,N_4964);
or U5974 (N_5974,N_4260,N_4346);
and U5975 (N_5975,N_4114,N_4919);
xor U5976 (N_5976,N_4645,N_4749);
nand U5977 (N_5977,N_4714,N_4682);
or U5978 (N_5978,N_4944,N_4446);
nor U5979 (N_5979,N_4952,N_4406);
nor U5980 (N_5980,N_4016,N_4094);
nor U5981 (N_5981,N_4689,N_4494);
or U5982 (N_5982,N_4444,N_4904);
nor U5983 (N_5983,N_4921,N_4602);
or U5984 (N_5984,N_4994,N_4520);
xnor U5985 (N_5985,N_4098,N_4011);
nor U5986 (N_5986,N_4802,N_4526);
xnor U5987 (N_5987,N_4256,N_4054);
xor U5988 (N_5988,N_4043,N_4427);
nand U5989 (N_5989,N_4474,N_4644);
and U5990 (N_5990,N_4652,N_4923);
or U5991 (N_5991,N_4061,N_4465);
xnor U5992 (N_5992,N_4937,N_4830);
nor U5993 (N_5993,N_4498,N_4508);
xnor U5994 (N_5994,N_4056,N_4177);
xnor U5995 (N_5995,N_4958,N_4651);
and U5996 (N_5996,N_4692,N_4040);
xor U5997 (N_5997,N_4047,N_4893);
nor U5998 (N_5998,N_4522,N_4167);
and U5999 (N_5999,N_4493,N_4388);
xnor U6000 (N_6000,N_5783,N_5487);
or U6001 (N_6001,N_5892,N_5836);
nand U6002 (N_6002,N_5765,N_5824);
and U6003 (N_6003,N_5705,N_5296);
or U6004 (N_6004,N_5440,N_5541);
nor U6005 (N_6005,N_5031,N_5166);
nor U6006 (N_6006,N_5211,N_5328);
nor U6007 (N_6007,N_5317,N_5297);
or U6008 (N_6008,N_5772,N_5723);
nand U6009 (N_6009,N_5147,N_5554);
nand U6010 (N_6010,N_5394,N_5999);
nor U6011 (N_6011,N_5965,N_5202);
and U6012 (N_6012,N_5600,N_5371);
nand U6013 (N_6013,N_5428,N_5033);
nor U6014 (N_6014,N_5351,N_5981);
xnor U6015 (N_6015,N_5054,N_5261);
nand U6016 (N_6016,N_5866,N_5458);
and U6017 (N_6017,N_5514,N_5167);
and U6018 (N_6018,N_5905,N_5753);
nor U6019 (N_6019,N_5254,N_5959);
nand U6020 (N_6020,N_5225,N_5642);
nor U6021 (N_6021,N_5365,N_5421);
nand U6022 (N_6022,N_5376,N_5862);
nand U6023 (N_6023,N_5855,N_5511);
or U6024 (N_6024,N_5145,N_5976);
nor U6025 (N_6025,N_5271,N_5689);
nor U6026 (N_6026,N_5092,N_5738);
and U6027 (N_6027,N_5633,N_5242);
xor U6028 (N_6028,N_5382,N_5764);
and U6029 (N_6029,N_5672,N_5653);
nor U6030 (N_6030,N_5333,N_5098);
nor U6031 (N_6031,N_5559,N_5178);
or U6032 (N_6032,N_5538,N_5477);
nor U6033 (N_6033,N_5832,N_5336);
and U6034 (N_6034,N_5160,N_5008);
nor U6035 (N_6035,N_5443,N_5692);
or U6036 (N_6036,N_5728,N_5006);
xnor U6037 (N_6037,N_5956,N_5679);
nor U6038 (N_6038,N_5597,N_5707);
and U6039 (N_6039,N_5932,N_5262);
and U6040 (N_6040,N_5907,N_5757);
and U6041 (N_6041,N_5940,N_5208);
nor U6042 (N_6042,N_5716,N_5185);
and U6043 (N_6043,N_5038,N_5220);
and U6044 (N_6044,N_5978,N_5209);
nand U6045 (N_6045,N_5341,N_5933);
nand U6046 (N_6046,N_5076,N_5936);
nand U6047 (N_6047,N_5485,N_5348);
nand U6048 (N_6048,N_5563,N_5044);
nor U6049 (N_6049,N_5164,N_5230);
and U6050 (N_6050,N_5708,N_5312);
nand U6051 (N_6051,N_5687,N_5389);
or U6052 (N_6052,N_5276,N_5378);
nand U6053 (N_6053,N_5015,N_5973);
nand U6054 (N_6054,N_5503,N_5318);
nand U6055 (N_6055,N_5391,N_5291);
or U6056 (N_6056,N_5839,N_5567);
and U6057 (N_6057,N_5626,N_5986);
and U6058 (N_6058,N_5950,N_5722);
nor U6059 (N_6059,N_5762,N_5255);
nand U6060 (N_6060,N_5499,N_5424);
nand U6061 (N_6061,N_5065,N_5850);
and U6062 (N_6062,N_5077,N_5073);
nand U6063 (N_6063,N_5158,N_5875);
or U6064 (N_6064,N_5683,N_5280);
or U6065 (N_6065,N_5685,N_5449);
nor U6066 (N_6066,N_5081,N_5340);
and U6067 (N_6067,N_5800,N_5446);
nor U6068 (N_6068,N_5970,N_5465);
nand U6069 (N_6069,N_5466,N_5364);
xor U6070 (N_6070,N_5086,N_5741);
nor U6071 (N_6071,N_5051,N_5068);
nor U6072 (N_6072,N_5174,N_5525);
nand U6073 (N_6073,N_5372,N_5612);
nor U6074 (N_6074,N_5769,N_5890);
nand U6075 (N_6075,N_5645,N_5197);
nor U6076 (N_6076,N_5238,N_5544);
or U6077 (N_6077,N_5183,N_5740);
or U6078 (N_6078,N_5789,N_5447);
nand U6079 (N_6079,N_5087,N_5593);
nand U6080 (N_6080,N_5797,N_5621);
nor U6081 (N_6081,N_5259,N_5265);
nor U6082 (N_6082,N_5019,N_5732);
and U6083 (N_6083,N_5515,N_5669);
or U6084 (N_6084,N_5561,N_5321);
and U6085 (N_6085,N_5270,N_5283);
nand U6086 (N_6086,N_5121,N_5591);
nor U6087 (N_6087,N_5982,N_5420);
nand U6088 (N_6088,N_5657,N_5100);
nor U6089 (N_6089,N_5846,N_5310);
or U6090 (N_6090,N_5269,N_5278);
and U6091 (N_6091,N_5405,N_5848);
nor U6092 (N_6092,N_5078,N_5432);
nor U6093 (N_6093,N_5744,N_5921);
or U6094 (N_6094,N_5709,N_5290);
nor U6095 (N_6095,N_5127,N_5878);
xnor U6096 (N_6096,N_5292,N_5095);
and U6097 (N_6097,N_5805,N_5287);
or U6098 (N_6098,N_5881,N_5506);
and U6099 (N_6099,N_5156,N_5461);
and U6100 (N_6100,N_5998,N_5129);
and U6101 (N_6101,N_5969,N_5879);
and U6102 (N_6102,N_5324,N_5688);
nor U6103 (N_6103,N_5693,N_5780);
nand U6104 (N_6104,N_5763,N_5471);
nor U6105 (N_6105,N_5751,N_5883);
nor U6106 (N_6106,N_5126,N_5216);
nor U6107 (N_6107,N_5553,N_5916);
nor U6108 (N_6108,N_5752,N_5516);
nor U6109 (N_6109,N_5545,N_5469);
nand U6110 (N_6110,N_5229,N_5074);
nor U6111 (N_6111,N_5686,N_5059);
nand U6112 (N_6112,N_5161,N_5429);
nor U6113 (N_6113,N_5279,N_5830);
or U6114 (N_6114,N_5346,N_5734);
nor U6115 (N_6115,N_5237,N_5355);
and U6116 (N_6116,N_5357,N_5188);
nor U6117 (N_6117,N_5856,N_5599);
xor U6118 (N_6118,N_5235,N_5628);
or U6119 (N_6119,N_5785,N_5569);
or U6120 (N_6120,N_5590,N_5402);
nor U6121 (N_6121,N_5968,N_5383);
nor U6122 (N_6122,N_5798,N_5560);
xor U6123 (N_6123,N_5223,N_5479);
and U6124 (N_6124,N_5681,N_5793);
or U6125 (N_6125,N_5721,N_5387);
and U6126 (N_6126,N_5849,N_5542);
and U6127 (N_6127,N_5775,N_5130);
nand U6128 (N_6128,N_5818,N_5462);
or U6129 (N_6129,N_5184,N_5580);
nor U6130 (N_6130,N_5181,N_5662);
and U6131 (N_6131,N_5467,N_5831);
and U6132 (N_6132,N_5901,N_5106);
nand U6133 (N_6133,N_5670,N_5408);
and U6134 (N_6134,N_5735,N_5637);
nor U6135 (N_6135,N_5241,N_5634);
xor U6136 (N_6136,N_5922,N_5674);
or U6137 (N_6137,N_5919,N_5007);
or U6138 (N_6138,N_5758,N_5551);
and U6139 (N_6139,N_5643,N_5110);
nand U6140 (N_6140,N_5997,N_5505);
or U6141 (N_6141,N_5954,N_5534);
nor U6142 (N_6142,N_5453,N_5690);
nand U6143 (N_6143,N_5894,N_5871);
or U6144 (N_6144,N_5934,N_5011);
nor U6145 (N_6145,N_5790,N_5718);
nor U6146 (N_6146,N_5345,N_5358);
nand U6147 (N_6147,N_5588,N_5049);
nand U6148 (N_6148,N_5491,N_5214);
or U6149 (N_6149,N_5926,N_5925);
and U6150 (N_6150,N_5729,N_5625);
nor U6151 (N_6151,N_5668,N_5808);
or U6152 (N_6152,N_5869,N_5966);
or U6153 (N_6153,N_5696,N_5444);
or U6154 (N_6154,N_5611,N_5946);
or U6155 (N_6155,N_5698,N_5598);
nand U6156 (N_6156,N_5566,N_5558);
and U6157 (N_6157,N_5097,N_5880);
nand U6158 (N_6158,N_5112,N_5826);
and U6159 (N_6159,N_5854,N_5517);
and U6160 (N_6160,N_5791,N_5114);
and U6161 (N_6161,N_5575,N_5811);
or U6162 (N_6162,N_5088,N_5961);
nor U6163 (N_6163,N_5974,N_5043);
xnor U6164 (N_6164,N_5638,N_5463);
or U6165 (N_6165,N_5017,N_5860);
and U6166 (N_6166,N_5799,N_5900);
and U6167 (N_6167,N_5963,N_5329);
xor U6168 (N_6168,N_5003,N_5748);
nand U6169 (N_6169,N_5437,N_5768);
and U6170 (N_6170,N_5400,N_5189);
nor U6171 (N_6171,N_5101,N_5293);
and U6172 (N_6172,N_5564,N_5439);
nor U6173 (N_6173,N_5971,N_5014);
and U6174 (N_6174,N_5330,N_5159);
nand U6175 (N_6175,N_5586,N_5825);
and U6176 (N_6176,N_5990,N_5834);
nor U6177 (N_6177,N_5964,N_5720);
nand U6178 (N_6178,N_5153,N_5710);
nand U6179 (N_6179,N_5574,N_5426);
and U6180 (N_6180,N_5838,N_5822);
nand U6181 (N_6181,N_5909,N_5029);
xor U6182 (N_6182,N_5996,N_5142);
or U6183 (N_6183,N_5360,N_5742);
nand U6184 (N_6184,N_5782,N_5908);
and U6185 (N_6185,N_5169,N_5170);
nand U6186 (N_6186,N_5256,N_5072);
or U6187 (N_6187,N_5131,N_5601);
and U6188 (N_6188,N_5647,N_5366);
or U6189 (N_6189,N_5770,N_5307);
and U6190 (N_6190,N_5585,N_5350);
and U6191 (N_6191,N_5109,N_5226);
nor U6192 (N_6192,N_5913,N_5141);
or U6193 (N_6193,N_5508,N_5306);
nor U6194 (N_6194,N_5117,N_5665);
nand U6195 (N_6195,N_5677,N_5386);
nor U6196 (N_6196,N_5781,N_5398);
nand U6197 (N_6197,N_5118,N_5565);
or U6198 (N_6198,N_5796,N_5263);
and U6199 (N_6199,N_5082,N_5935);
nor U6200 (N_6200,N_5396,N_5221);
or U6201 (N_6201,N_5438,N_5298);
nor U6202 (N_6202,N_5667,N_5388);
and U6203 (N_6203,N_5417,N_5552);
and U6204 (N_6204,N_5264,N_5979);
nor U6205 (N_6205,N_5102,N_5134);
nor U6206 (N_6206,N_5556,N_5246);
nand U6207 (N_6207,N_5149,N_5823);
or U6208 (N_6208,N_5039,N_5630);
nor U6209 (N_6209,N_5025,N_5171);
and U6210 (N_6210,N_5344,N_5532);
or U6211 (N_6211,N_5107,N_5509);
nand U6212 (N_6212,N_5460,N_5260);
xor U6213 (N_6213,N_5804,N_5457);
nand U6214 (N_6214,N_5172,N_5540);
and U6215 (N_6215,N_5309,N_5472);
or U6216 (N_6216,N_5018,N_5475);
nor U6217 (N_6217,N_5401,N_5481);
nor U6218 (N_6218,N_5085,N_5984);
and U6219 (N_6219,N_5062,N_5607);
xnor U6220 (N_6220,N_5887,N_5577);
or U6221 (N_6221,N_5198,N_5119);
nand U6222 (N_6222,N_5010,N_5652);
nand U6223 (N_6223,N_5803,N_5617);
and U6224 (N_6224,N_5434,N_5157);
nand U6225 (N_6225,N_5143,N_5406);
nor U6226 (N_6226,N_5442,N_5711);
nand U6227 (N_6227,N_5285,N_5841);
or U6228 (N_6228,N_5592,N_5493);
or U6229 (N_6229,N_5622,N_5247);
or U6230 (N_6230,N_5904,N_5616);
nor U6231 (N_6231,N_5245,N_5303);
nand U6232 (N_6232,N_5060,N_5064);
nor U6233 (N_6233,N_5058,N_5486);
nor U6234 (N_6234,N_5301,N_5089);
nand U6235 (N_6235,N_5299,N_5137);
nand U6236 (N_6236,N_5536,N_5635);
and U6237 (N_6237,N_5316,N_5222);
xor U6238 (N_6238,N_5882,N_5191);
or U6239 (N_6239,N_5473,N_5488);
nand U6240 (N_6240,N_5988,N_5323);
or U6241 (N_6241,N_5093,N_5132);
or U6242 (N_6242,N_5024,N_5608);
nor U6243 (N_6243,N_5951,N_5821);
nor U6244 (N_6244,N_5727,N_5650);
xnor U6245 (N_6245,N_5339,N_5148);
or U6246 (N_6246,N_5482,N_5792);
xnor U6247 (N_6247,N_5187,N_5067);
or U6248 (N_6248,N_5070,N_5726);
nand U6249 (N_6249,N_5828,N_5987);
nor U6250 (N_6250,N_5320,N_5352);
and U6251 (N_6251,N_5958,N_5957);
or U6252 (N_6252,N_5546,N_5801);
nand U6253 (N_6253,N_5991,N_5615);
nand U6254 (N_6254,N_5362,N_5123);
nand U6255 (N_6255,N_5243,N_5703);
nand U6256 (N_6256,N_5176,N_5928);
or U6257 (N_6257,N_5873,N_5817);
nor U6258 (N_6258,N_5195,N_5455);
or U6259 (N_6259,N_5224,N_5094);
and U6260 (N_6260,N_5527,N_5448);
and U6261 (N_6261,N_5530,N_5994);
xor U6262 (N_6262,N_5639,N_5390);
or U6263 (N_6263,N_5501,N_5807);
and U6264 (N_6264,N_5182,N_5993);
xnor U6265 (N_6265,N_5057,N_5080);
xor U6266 (N_6266,N_5613,N_5199);
and U6267 (N_6267,N_5368,N_5941);
nor U6268 (N_6268,N_5250,N_5234);
nor U6269 (N_6269,N_5138,N_5050);
or U6270 (N_6270,N_5699,N_5535);
nand U6271 (N_6271,N_5844,N_5743);
and U6272 (N_6272,N_5004,N_5655);
and U6273 (N_6273,N_5450,N_5203);
nand U6274 (N_6274,N_5146,N_5845);
or U6275 (N_6275,N_5717,N_5179);
nor U6276 (N_6276,N_5165,N_5498);
and U6277 (N_6277,N_5416,N_5659);
nor U6278 (N_6278,N_5194,N_5300);
nand U6279 (N_6279,N_5305,N_5929);
nand U6280 (N_6280,N_5370,N_5550);
nand U6281 (N_6281,N_5474,N_5651);
or U6282 (N_6282,N_5380,N_5190);
nor U6283 (N_6283,N_5528,N_5620);
xor U6284 (N_6284,N_5492,N_5512);
nand U6285 (N_6285,N_5927,N_5337);
or U6286 (N_6286,N_5867,N_5483);
nand U6287 (N_6287,N_5724,N_5034);
or U6288 (N_6288,N_5295,N_5713);
nand U6289 (N_6289,N_5331,N_5257);
and U6290 (N_6290,N_5543,N_5750);
nor U6291 (N_6291,N_5314,N_5009);
nand U6292 (N_6292,N_5409,N_5691);
or U6293 (N_6293,N_5374,N_5228);
nor U6294 (N_6294,N_5273,N_5572);
nand U6295 (N_6295,N_5335,N_5120);
nand U6296 (N_6296,N_5342,N_5864);
or U6297 (N_6297,N_5403,N_5837);
nand U6298 (N_6298,N_5454,N_5053);
nor U6299 (N_6299,N_5128,N_5500);
and U6300 (N_6300,N_5829,N_5624);
nor U6301 (N_6301,N_5938,N_5215);
and U6302 (N_6302,N_5016,N_5694);
nand U6303 (N_6303,N_5001,N_5452);
nand U6304 (N_6304,N_5524,N_5573);
and U6305 (N_6305,N_5952,N_5249);
or U6306 (N_6306,N_5464,N_5795);
nand U6307 (N_6307,N_5055,N_5893);
nor U6308 (N_6308,N_5985,N_5023);
nand U6309 (N_6309,N_5377,N_5806);
and U6310 (N_6310,N_5851,N_5902);
nand U6311 (N_6311,N_5857,N_5091);
or U6312 (N_6312,N_5910,N_5745);
nor U6313 (N_6313,N_5431,N_5213);
nand U6314 (N_6314,N_5407,N_5108);
and U6315 (N_6315,N_5605,N_5583);
nand U6316 (N_6316,N_5547,N_5771);
xnor U6317 (N_6317,N_5036,N_5787);
nor U6318 (N_6318,N_5139,N_5923);
xnor U6319 (N_6319,N_5361,N_5218);
or U6320 (N_6320,N_5529,N_5026);
nor U6321 (N_6321,N_5325,N_5338);
or U6322 (N_6322,N_5664,N_5210);
xnor U6323 (N_6323,N_5549,N_5570);
xor U6324 (N_6324,N_5392,N_5504);
nand U6325 (N_6325,N_5548,N_5779);
or U6326 (N_6326,N_5063,N_5332);
or U6327 (N_6327,N_5778,N_5356);
nand U6328 (N_6328,N_5267,N_5737);
and U6329 (N_6329,N_5497,N_5582);
or U6330 (N_6330,N_5914,N_5122);
nor U6331 (N_6331,N_5012,N_5168);
nor U6332 (N_6332,N_5843,N_5937);
and U6333 (N_6333,N_5980,N_5385);
or U6334 (N_6334,N_5173,N_5813);
or U6335 (N_6335,N_5676,N_5313);
nor U6336 (N_6336,N_5820,N_5510);
nor U6337 (N_6337,N_5456,N_5631);
or U6338 (N_6338,N_5819,N_5614);
and U6339 (N_6339,N_5111,N_5636);
nor U6340 (N_6340,N_5319,N_5103);
nand U6341 (N_6341,N_5842,N_5353);
nor U6342 (N_6342,N_5046,N_5595);
nand U6343 (N_6343,N_5289,N_5911);
nor U6344 (N_6344,N_5661,N_5606);
nand U6345 (N_6345,N_5571,N_5885);
or U6346 (N_6346,N_5193,N_5706);
and U6347 (N_6347,N_5150,N_5411);
or U6348 (N_6348,N_5872,N_5675);
or U6349 (N_6349,N_5253,N_5602);
or U6350 (N_6350,N_5468,N_5079);
nor U6351 (N_6351,N_5695,N_5373);
nand U6352 (N_6352,N_5747,N_5939);
or U6353 (N_6353,N_5186,N_5489);
nand U6354 (N_6354,N_5604,N_5136);
nor U6355 (N_6355,N_5140,N_5040);
nor U6356 (N_6356,N_5311,N_5833);
nor U6357 (N_6357,N_5632,N_5603);
or U6358 (N_6358,N_5920,N_5537);
or U6359 (N_6359,N_5495,N_5519);
nor U6360 (N_6360,N_5955,N_5056);
nand U6361 (N_6361,N_5702,N_5490);
or U6362 (N_6362,N_5644,N_5286);
and U6363 (N_6363,N_5144,N_5105);
or U6364 (N_6364,N_5863,N_5539);
or U6365 (N_6365,N_5725,N_5268);
and U6366 (N_6366,N_5349,N_5983);
nand U6367 (N_6367,N_5656,N_5281);
and U6368 (N_6368,N_5066,N_5113);
xor U6369 (N_6369,N_5619,N_5576);
xor U6370 (N_6370,N_5252,N_5413);
or U6371 (N_6371,N_5115,N_5163);
and U6372 (N_6372,N_5944,N_5354);
nor U6373 (N_6373,N_5714,N_5897);
and U6374 (N_6374,N_5419,N_5761);
xnor U6375 (N_6375,N_5589,N_5244);
and U6376 (N_6376,N_5212,N_5618);
and U6377 (N_6377,N_5096,N_5395);
and U6378 (N_6378,N_5272,N_5609);
and U6379 (N_6379,N_5898,N_5021);
and U6380 (N_6380,N_5304,N_5906);
nand U6381 (N_6381,N_5206,N_5410);
and U6382 (N_6382,N_5784,N_5042);
nand U6383 (N_6383,N_5816,N_5649);
nand U6384 (N_6384,N_5423,N_5531);
or U6385 (N_6385,N_5526,N_5302);
and U6386 (N_6386,N_5384,N_5562);
nor U6387 (N_6387,N_5673,N_5022);
or U6388 (N_6388,N_5217,N_5967);
or U6389 (N_6389,N_5629,N_5061);
nand U6390 (N_6390,N_5084,N_5731);
xnor U6391 (N_6391,N_5654,N_5903);
xnor U6392 (N_6392,N_5641,N_5523);
nor U6393 (N_6393,N_5658,N_5557);
and U6394 (N_6394,N_5786,N_5513);
nand U6395 (N_6395,N_5294,N_5041);
nor U6396 (N_6396,N_5322,N_5960);
xor U6397 (N_6397,N_5133,N_5759);
nor U6398 (N_6398,N_5404,N_5104);
nand U6399 (N_6399,N_5739,N_5258);
nand U6400 (N_6400,N_5874,N_5773);
nand U6401 (N_6401,N_5470,N_5663);
nor U6402 (N_6402,N_5367,N_5697);
nand U6403 (N_6403,N_5277,N_5135);
xnor U6404 (N_6404,N_5847,N_5840);
nand U6405 (N_6405,N_5918,N_5415);
nand U6406 (N_6406,N_5520,N_5436);
nor U6407 (N_6407,N_5746,N_5680);
and U6408 (N_6408,N_5766,N_5870);
nand U6409 (N_6409,N_5594,N_5877);
or U6410 (N_6410,N_5835,N_5712);
xnor U6411 (N_6411,N_5240,N_5930);
and U6412 (N_6412,N_5756,N_5155);
and U6413 (N_6413,N_5774,N_5427);
nor U6414 (N_6414,N_5949,N_5733);
nand U6415 (N_6415,N_5518,N_5414);
nand U6416 (N_6416,N_5977,N_5931);
or U6417 (N_6417,N_5700,N_5266);
nor U6418 (N_6418,N_5125,N_5480);
or U6419 (N_6419,N_5083,N_5578);
xor U6420 (N_6420,N_5975,N_5891);
nand U6421 (N_6421,N_5451,N_5852);
nand U6422 (N_6422,N_5175,N_5251);
and U6423 (N_6423,N_5484,N_5284);
xnor U6424 (N_6424,N_5719,N_5418);
nor U6425 (N_6425,N_5177,N_5204);
and U6426 (N_6426,N_5776,N_5942);
and U6427 (N_6427,N_5610,N_5522);
nand U6428 (N_6428,N_5777,N_5124);
nand U6429 (N_6429,N_5858,N_5200);
or U6430 (N_6430,N_5393,N_5555);
nand U6431 (N_6431,N_5648,N_5749);
nor U6432 (N_6432,N_5827,N_5888);
nor U6433 (N_6433,N_5627,N_5326);
nor U6434 (N_6434,N_5045,N_5399);
and U6435 (N_6435,N_5359,N_5381);
xor U6436 (N_6436,N_5682,N_5899);
nand U6437 (N_6437,N_5005,N_5507);
nand U6438 (N_6438,N_5227,N_5995);
xor U6439 (N_6439,N_5037,N_5496);
nand U6440 (N_6440,N_5945,N_5815);
or U6441 (N_6441,N_5116,N_5205);
or U6442 (N_6442,N_5917,N_5274);
and U6443 (N_6443,N_5347,N_5027);
and U6444 (N_6444,N_5861,N_5219);
nand U6445 (N_6445,N_5052,N_5275);
and U6446 (N_6446,N_5730,N_5886);
nor U6447 (N_6447,N_5868,N_5236);
nand U6448 (N_6448,N_5231,N_5099);
nor U6449 (N_6449,N_5239,N_5154);
nand U6450 (N_6450,N_5327,N_5048);
nor U6451 (N_6451,N_5736,N_5794);
xor U6452 (N_6452,N_5334,N_5075);
and U6453 (N_6453,N_5754,N_5912);
and U6454 (N_6454,N_5948,N_5678);
nor U6455 (N_6455,N_5884,N_5020);
or U6456 (N_6456,N_5315,N_5397);
or U6457 (N_6457,N_5028,N_5152);
nor U6458 (N_6458,N_5533,N_5032);
nand U6459 (N_6459,N_5915,N_5375);
or U6460 (N_6460,N_5412,N_5207);
or U6461 (N_6461,N_5000,N_5379);
and U6462 (N_6462,N_5002,N_5684);
and U6463 (N_6463,N_5895,N_5972);
nand U6464 (N_6464,N_5232,N_5445);
or U6465 (N_6465,N_5201,N_5701);
or U6466 (N_6466,N_5814,N_5853);
or U6467 (N_6467,N_5802,N_5308);
and U6468 (N_6468,N_5596,N_5992);
and U6469 (N_6469,N_5476,N_5671);
xor U6470 (N_6470,N_5579,N_5581);
nor U6471 (N_6471,N_5865,N_5013);
nand U6472 (N_6472,N_5760,N_5889);
nor U6473 (N_6473,N_5755,N_5069);
nand U6474 (N_6474,N_5896,N_5478);
nor U6475 (N_6475,N_5422,N_5876);
nor U6476 (N_6476,N_5030,N_5640);
xor U6477 (N_6477,N_5425,N_5282);
or U6478 (N_6478,N_5180,N_5071);
nand U6479 (N_6479,N_5584,N_5363);
nand U6480 (N_6480,N_5646,N_5192);
and U6481 (N_6481,N_5623,N_5810);
and U6482 (N_6482,N_5767,N_5568);
or U6483 (N_6483,N_5441,N_5704);
and U6484 (N_6484,N_5924,N_5859);
or U6485 (N_6485,N_5090,N_5288);
nor U6486 (N_6486,N_5162,N_5943);
nand U6487 (N_6487,N_5521,N_5494);
or U6488 (N_6488,N_5343,N_5947);
xnor U6489 (N_6489,N_5502,N_5435);
and U6490 (N_6490,N_5459,N_5788);
nand U6491 (N_6491,N_5233,N_5953);
nor U6492 (N_6492,N_5666,N_5812);
xnor U6493 (N_6493,N_5989,N_5962);
nand U6494 (N_6494,N_5715,N_5369);
and U6495 (N_6495,N_5809,N_5248);
or U6496 (N_6496,N_5433,N_5047);
and U6497 (N_6497,N_5587,N_5660);
nor U6498 (N_6498,N_5196,N_5151);
or U6499 (N_6499,N_5035,N_5430);
and U6500 (N_6500,N_5774,N_5448);
or U6501 (N_6501,N_5214,N_5807);
or U6502 (N_6502,N_5785,N_5692);
and U6503 (N_6503,N_5761,N_5681);
nor U6504 (N_6504,N_5790,N_5430);
nor U6505 (N_6505,N_5220,N_5474);
or U6506 (N_6506,N_5411,N_5164);
or U6507 (N_6507,N_5300,N_5038);
nand U6508 (N_6508,N_5983,N_5208);
and U6509 (N_6509,N_5378,N_5083);
nor U6510 (N_6510,N_5180,N_5749);
and U6511 (N_6511,N_5660,N_5058);
nor U6512 (N_6512,N_5853,N_5942);
nor U6513 (N_6513,N_5633,N_5332);
nand U6514 (N_6514,N_5524,N_5080);
nand U6515 (N_6515,N_5549,N_5305);
and U6516 (N_6516,N_5777,N_5430);
nor U6517 (N_6517,N_5391,N_5886);
nor U6518 (N_6518,N_5699,N_5568);
nor U6519 (N_6519,N_5215,N_5046);
nor U6520 (N_6520,N_5963,N_5974);
nor U6521 (N_6521,N_5804,N_5643);
or U6522 (N_6522,N_5249,N_5599);
nor U6523 (N_6523,N_5866,N_5709);
nand U6524 (N_6524,N_5773,N_5981);
and U6525 (N_6525,N_5154,N_5700);
or U6526 (N_6526,N_5071,N_5192);
xnor U6527 (N_6527,N_5950,N_5576);
and U6528 (N_6528,N_5562,N_5539);
or U6529 (N_6529,N_5842,N_5476);
nor U6530 (N_6530,N_5020,N_5707);
and U6531 (N_6531,N_5839,N_5111);
or U6532 (N_6532,N_5840,N_5541);
and U6533 (N_6533,N_5712,N_5546);
or U6534 (N_6534,N_5647,N_5031);
xor U6535 (N_6535,N_5721,N_5462);
nor U6536 (N_6536,N_5260,N_5645);
xnor U6537 (N_6537,N_5956,N_5308);
nor U6538 (N_6538,N_5951,N_5193);
nor U6539 (N_6539,N_5684,N_5154);
nor U6540 (N_6540,N_5837,N_5948);
xnor U6541 (N_6541,N_5613,N_5643);
nor U6542 (N_6542,N_5698,N_5300);
nand U6543 (N_6543,N_5475,N_5030);
and U6544 (N_6544,N_5392,N_5265);
or U6545 (N_6545,N_5103,N_5470);
nor U6546 (N_6546,N_5491,N_5965);
nor U6547 (N_6547,N_5785,N_5765);
xnor U6548 (N_6548,N_5762,N_5333);
xor U6549 (N_6549,N_5326,N_5135);
and U6550 (N_6550,N_5125,N_5907);
xnor U6551 (N_6551,N_5070,N_5290);
and U6552 (N_6552,N_5608,N_5027);
and U6553 (N_6553,N_5853,N_5277);
nor U6554 (N_6554,N_5574,N_5296);
and U6555 (N_6555,N_5141,N_5970);
and U6556 (N_6556,N_5803,N_5954);
nand U6557 (N_6557,N_5753,N_5222);
nor U6558 (N_6558,N_5857,N_5949);
or U6559 (N_6559,N_5954,N_5869);
and U6560 (N_6560,N_5588,N_5144);
and U6561 (N_6561,N_5466,N_5270);
or U6562 (N_6562,N_5667,N_5400);
or U6563 (N_6563,N_5013,N_5841);
xor U6564 (N_6564,N_5692,N_5847);
xor U6565 (N_6565,N_5617,N_5788);
or U6566 (N_6566,N_5785,N_5734);
nand U6567 (N_6567,N_5241,N_5557);
and U6568 (N_6568,N_5937,N_5329);
and U6569 (N_6569,N_5407,N_5652);
nand U6570 (N_6570,N_5994,N_5374);
nor U6571 (N_6571,N_5014,N_5729);
xnor U6572 (N_6572,N_5151,N_5955);
and U6573 (N_6573,N_5288,N_5392);
and U6574 (N_6574,N_5441,N_5336);
nor U6575 (N_6575,N_5296,N_5840);
and U6576 (N_6576,N_5415,N_5976);
nand U6577 (N_6577,N_5094,N_5336);
nand U6578 (N_6578,N_5018,N_5595);
and U6579 (N_6579,N_5922,N_5154);
and U6580 (N_6580,N_5147,N_5580);
and U6581 (N_6581,N_5366,N_5100);
nor U6582 (N_6582,N_5884,N_5840);
and U6583 (N_6583,N_5247,N_5575);
xnor U6584 (N_6584,N_5577,N_5769);
or U6585 (N_6585,N_5391,N_5926);
or U6586 (N_6586,N_5295,N_5947);
or U6587 (N_6587,N_5396,N_5008);
nand U6588 (N_6588,N_5384,N_5387);
and U6589 (N_6589,N_5110,N_5189);
or U6590 (N_6590,N_5297,N_5575);
and U6591 (N_6591,N_5830,N_5340);
nor U6592 (N_6592,N_5209,N_5256);
nor U6593 (N_6593,N_5825,N_5849);
nand U6594 (N_6594,N_5720,N_5693);
xor U6595 (N_6595,N_5833,N_5174);
xor U6596 (N_6596,N_5388,N_5319);
nor U6597 (N_6597,N_5314,N_5776);
xor U6598 (N_6598,N_5053,N_5211);
and U6599 (N_6599,N_5021,N_5884);
nor U6600 (N_6600,N_5823,N_5138);
or U6601 (N_6601,N_5700,N_5491);
nand U6602 (N_6602,N_5029,N_5027);
or U6603 (N_6603,N_5582,N_5584);
xnor U6604 (N_6604,N_5131,N_5037);
nor U6605 (N_6605,N_5204,N_5100);
and U6606 (N_6606,N_5047,N_5915);
or U6607 (N_6607,N_5778,N_5558);
nand U6608 (N_6608,N_5044,N_5832);
or U6609 (N_6609,N_5633,N_5637);
and U6610 (N_6610,N_5533,N_5661);
or U6611 (N_6611,N_5538,N_5239);
or U6612 (N_6612,N_5995,N_5887);
and U6613 (N_6613,N_5355,N_5763);
nand U6614 (N_6614,N_5650,N_5474);
and U6615 (N_6615,N_5422,N_5886);
or U6616 (N_6616,N_5200,N_5913);
and U6617 (N_6617,N_5182,N_5690);
nand U6618 (N_6618,N_5408,N_5853);
and U6619 (N_6619,N_5326,N_5874);
nand U6620 (N_6620,N_5108,N_5384);
or U6621 (N_6621,N_5304,N_5839);
xnor U6622 (N_6622,N_5044,N_5017);
nor U6623 (N_6623,N_5248,N_5715);
and U6624 (N_6624,N_5415,N_5807);
nor U6625 (N_6625,N_5888,N_5467);
xnor U6626 (N_6626,N_5174,N_5066);
nor U6627 (N_6627,N_5623,N_5196);
xor U6628 (N_6628,N_5535,N_5582);
nor U6629 (N_6629,N_5105,N_5267);
or U6630 (N_6630,N_5141,N_5874);
and U6631 (N_6631,N_5472,N_5816);
nor U6632 (N_6632,N_5426,N_5847);
and U6633 (N_6633,N_5105,N_5630);
or U6634 (N_6634,N_5571,N_5005);
and U6635 (N_6635,N_5663,N_5425);
and U6636 (N_6636,N_5336,N_5258);
and U6637 (N_6637,N_5364,N_5372);
nand U6638 (N_6638,N_5297,N_5630);
or U6639 (N_6639,N_5461,N_5051);
nor U6640 (N_6640,N_5594,N_5484);
or U6641 (N_6641,N_5817,N_5965);
and U6642 (N_6642,N_5990,N_5671);
and U6643 (N_6643,N_5982,N_5748);
nor U6644 (N_6644,N_5137,N_5007);
nor U6645 (N_6645,N_5448,N_5013);
nand U6646 (N_6646,N_5253,N_5557);
nand U6647 (N_6647,N_5266,N_5925);
nor U6648 (N_6648,N_5092,N_5614);
or U6649 (N_6649,N_5604,N_5416);
or U6650 (N_6650,N_5406,N_5250);
xor U6651 (N_6651,N_5863,N_5988);
or U6652 (N_6652,N_5137,N_5851);
or U6653 (N_6653,N_5885,N_5100);
and U6654 (N_6654,N_5660,N_5813);
xnor U6655 (N_6655,N_5576,N_5680);
nor U6656 (N_6656,N_5863,N_5509);
nor U6657 (N_6657,N_5957,N_5174);
and U6658 (N_6658,N_5794,N_5397);
nand U6659 (N_6659,N_5913,N_5841);
nor U6660 (N_6660,N_5358,N_5153);
and U6661 (N_6661,N_5950,N_5009);
nor U6662 (N_6662,N_5694,N_5247);
or U6663 (N_6663,N_5318,N_5841);
or U6664 (N_6664,N_5767,N_5231);
or U6665 (N_6665,N_5624,N_5155);
nand U6666 (N_6666,N_5786,N_5994);
xor U6667 (N_6667,N_5811,N_5979);
and U6668 (N_6668,N_5322,N_5613);
and U6669 (N_6669,N_5130,N_5075);
or U6670 (N_6670,N_5275,N_5605);
and U6671 (N_6671,N_5142,N_5213);
or U6672 (N_6672,N_5187,N_5295);
or U6673 (N_6673,N_5936,N_5825);
or U6674 (N_6674,N_5701,N_5238);
nor U6675 (N_6675,N_5670,N_5497);
or U6676 (N_6676,N_5740,N_5011);
and U6677 (N_6677,N_5587,N_5545);
and U6678 (N_6678,N_5441,N_5649);
nor U6679 (N_6679,N_5148,N_5587);
xor U6680 (N_6680,N_5143,N_5072);
nor U6681 (N_6681,N_5261,N_5617);
xnor U6682 (N_6682,N_5140,N_5467);
nand U6683 (N_6683,N_5397,N_5551);
nor U6684 (N_6684,N_5889,N_5383);
and U6685 (N_6685,N_5626,N_5343);
and U6686 (N_6686,N_5232,N_5842);
nor U6687 (N_6687,N_5011,N_5580);
or U6688 (N_6688,N_5738,N_5287);
or U6689 (N_6689,N_5814,N_5932);
nor U6690 (N_6690,N_5394,N_5283);
xnor U6691 (N_6691,N_5179,N_5033);
nor U6692 (N_6692,N_5468,N_5943);
xnor U6693 (N_6693,N_5931,N_5886);
or U6694 (N_6694,N_5448,N_5060);
or U6695 (N_6695,N_5127,N_5853);
nor U6696 (N_6696,N_5425,N_5631);
xor U6697 (N_6697,N_5328,N_5264);
nand U6698 (N_6698,N_5078,N_5365);
nor U6699 (N_6699,N_5107,N_5778);
nand U6700 (N_6700,N_5549,N_5147);
nor U6701 (N_6701,N_5443,N_5910);
and U6702 (N_6702,N_5091,N_5213);
nor U6703 (N_6703,N_5894,N_5928);
and U6704 (N_6704,N_5184,N_5713);
nand U6705 (N_6705,N_5678,N_5673);
nor U6706 (N_6706,N_5210,N_5901);
nand U6707 (N_6707,N_5191,N_5205);
and U6708 (N_6708,N_5511,N_5589);
and U6709 (N_6709,N_5202,N_5188);
nor U6710 (N_6710,N_5513,N_5943);
nand U6711 (N_6711,N_5652,N_5656);
and U6712 (N_6712,N_5687,N_5319);
xor U6713 (N_6713,N_5750,N_5097);
and U6714 (N_6714,N_5072,N_5849);
or U6715 (N_6715,N_5668,N_5814);
and U6716 (N_6716,N_5566,N_5936);
and U6717 (N_6717,N_5348,N_5133);
nand U6718 (N_6718,N_5793,N_5118);
and U6719 (N_6719,N_5792,N_5051);
nand U6720 (N_6720,N_5395,N_5649);
nand U6721 (N_6721,N_5647,N_5489);
or U6722 (N_6722,N_5089,N_5198);
xor U6723 (N_6723,N_5827,N_5632);
or U6724 (N_6724,N_5798,N_5073);
or U6725 (N_6725,N_5536,N_5265);
nor U6726 (N_6726,N_5407,N_5522);
nor U6727 (N_6727,N_5120,N_5545);
and U6728 (N_6728,N_5801,N_5051);
or U6729 (N_6729,N_5519,N_5328);
nor U6730 (N_6730,N_5879,N_5717);
nand U6731 (N_6731,N_5314,N_5455);
and U6732 (N_6732,N_5877,N_5048);
nand U6733 (N_6733,N_5226,N_5542);
and U6734 (N_6734,N_5955,N_5572);
or U6735 (N_6735,N_5906,N_5842);
and U6736 (N_6736,N_5552,N_5252);
xor U6737 (N_6737,N_5221,N_5952);
nand U6738 (N_6738,N_5719,N_5485);
nor U6739 (N_6739,N_5209,N_5327);
nor U6740 (N_6740,N_5559,N_5036);
and U6741 (N_6741,N_5918,N_5764);
and U6742 (N_6742,N_5234,N_5701);
or U6743 (N_6743,N_5234,N_5349);
or U6744 (N_6744,N_5526,N_5790);
and U6745 (N_6745,N_5368,N_5859);
nor U6746 (N_6746,N_5328,N_5799);
nand U6747 (N_6747,N_5321,N_5597);
or U6748 (N_6748,N_5521,N_5872);
xor U6749 (N_6749,N_5743,N_5258);
xor U6750 (N_6750,N_5059,N_5133);
nor U6751 (N_6751,N_5808,N_5937);
or U6752 (N_6752,N_5154,N_5575);
nor U6753 (N_6753,N_5337,N_5234);
or U6754 (N_6754,N_5214,N_5880);
or U6755 (N_6755,N_5555,N_5761);
nor U6756 (N_6756,N_5487,N_5164);
nor U6757 (N_6757,N_5183,N_5816);
and U6758 (N_6758,N_5497,N_5365);
or U6759 (N_6759,N_5800,N_5647);
xor U6760 (N_6760,N_5401,N_5318);
nor U6761 (N_6761,N_5321,N_5814);
xnor U6762 (N_6762,N_5999,N_5411);
nand U6763 (N_6763,N_5727,N_5130);
nor U6764 (N_6764,N_5704,N_5624);
nor U6765 (N_6765,N_5343,N_5752);
nand U6766 (N_6766,N_5875,N_5061);
or U6767 (N_6767,N_5909,N_5729);
nor U6768 (N_6768,N_5400,N_5402);
xor U6769 (N_6769,N_5157,N_5604);
nand U6770 (N_6770,N_5975,N_5777);
or U6771 (N_6771,N_5917,N_5190);
or U6772 (N_6772,N_5350,N_5704);
or U6773 (N_6773,N_5231,N_5539);
xor U6774 (N_6774,N_5449,N_5066);
nor U6775 (N_6775,N_5290,N_5711);
and U6776 (N_6776,N_5973,N_5980);
or U6777 (N_6777,N_5345,N_5986);
and U6778 (N_6778,N_5767,N_5055);
nand U6779 (N_6779,N_5881,N_5677);
nor U6780 (N_6780,N_5652,N_5985);
and U6781 (N_6781,N_5229,N_5286);
xor U6782 (N_6782,N_5353,N_5312);
xnor U6783 (N_6783,N_5071,N_5365);
or U6784 (N_6784,N_5712,N_5613);
and U6785 (N_6785,N_5628,N_5136);
nand U6786 (N_6786,N_5845,N_5140);
nand U6787 (N_6787,N_5038,N_5181);
and U6788 (N_6788,N_5453,N_5868);
nor U6789 (N_6789,N_5871,N_5414);
nand U6790 (N_6790,N_5994,N_5063);
xor U6791 (N_6791,N_5600,N_5577);
nor U6792 (N_6792,N_5246,N_5275);
nand U6793 (N_6793,N_5316,N_5848);
nand U6794 (N_6794,N_5034,N_5237);
or U6795 (N_6795,N_5142,N_5269);
or U6796 (N_6796,N_5226,N_5362);
nor U6797 (N_6797,N_5512,N_5729);
or U6798 (N_6798,N_5889,N_5040);
nand U6799 (N_6799,N_5256,N_5832);
or U6800 (N_6800,N_5217,N_5280);
nor U6801 (N_6801,N_5306,N_5104);
and U6802 (N_6802,N_5332,N_5471);
nand U6803 (N_6803,N_5502,N_5783);
nor U6804 (N_6804,N_5140,N_5211);
xor U6805 (N_6805,N_5915,N_5525);
nor U6806 (N_6806,N_5509,N_5190);
nor U6807 (N_6807,N_5181,N_5115);
xor U6808 (N_6808,N_5715,N_5737);
or U6809 (N_6809,N_5482,N_5691);
or U6810 (N_6810,N_5678,N_5953);
or U6811 (N_6811,N_5169,N_5318);
and U6812 (N_6812,N_5835,N_5968);
nand U6813 (N_6813,N_5587,N_5122);
and U6814 (N_6814,N_5178,N_5137);
nand U6815 (N_6815,N_5483,N_5511);
and U6816 (N_6816,N_5905,N_5446);
nor U6817 (N_6817,N_5898,N_5751);
nand U6818 (N_6818,N_5973,N_5302);
nand U6819 (N_6819,N_5952,N_5555);
nor U6820 (N_6820,N_5975,N_5259);
nor U6821 (N_6821,N_5333,N_5980);
or U6822 (N_6822,N_5481,N_5183);
nand U6823 (N_6823,N_5853,N_5664);
and U6824 (N_6824,N_5748,N_5474);
nand U6825 (N_6825,N_5484,N_5410);
and U6826 (N_6826,N_5985,N_5524);
nand U6827 (N_6827,N_5216,N_5875);
nand U6828 (N_6828,N_5881,N_5113);
nand U6829 (N_6829,N_5033,N_5354);
nand U6830 (N_6830,N_5021,N_5643);
nor U6831 (N_6831,N_5681,N_5463);
or U6832 (N_6832,N_5811,N_5475);
nor U6833 (N_6833,N_5079,N_5425);
or U6834 (N_6834,N_5873,N_5793);
nand U6835 (N_6835,N_5978,N_5787);
xor U6836 (N_6836,N_5109,N_5716);
nor U6837 (N_6837,N_5233,N_5468);
or U6838 (N_6838,N_5072,N_5865);
nand U6839 (N_6839,N_5920,N_5159);
nand U6840 (N_6840,N_5807,N_5383);
or U6841 (N_6841,N_5953,N_5934);
nor U6842 (N_6842,N_5529,N_5861);
and U6843 (N_6843,N_5941,N_5258);
nand U6844 (N_6844,N_5006,N_5911);
nor U6845 (N_6845,N_5872,N_5833);
and U6846 (N_6846,N_5038,N_5819);
xor U6847 (N_6847,N_5606,N_5663);
or U6848 (N_6848,N_5953,N_5335);
nand U6849 (N_6849,N_5585,N_5824);
or U6850 (N_6850,N_5849,N_5858);
xnor U6851 (N_6851,N_5669,N_5420);
or U6852 (N_6852,N_5090,N_5628);
or U6853 (N_6853,N_5497,N_5815);
or U6854 (N_6854,N_5345,N_5526);
xnor U6855 (N_6855,N_5542,N_5054);
nor U6856 (N_6856,N_5942,N_5732);
or U6857 (N_6857,N_5584,N_5094);
nand U6858 (N_6858,N_5267,N_5709);
or U6859 (N_6859,N_5057,N_5968);
nand U6860 (N_6860,N_5117,N_5715);
or U6861 (N_6861,N_5150,N_5443);
or U6862 (N_6862,N_5154,N_5784);
nand U6863 (N_6863,N_5199,N_5194);
nor U6864 (N_6864,N_5423,N_5455);
nor U6865 (N_6865,N_5381,N_5667);
nand U6866 (N_6866,N_5352,N_5259);
or U6867 (N_6867,N_5183,N_5725);
and U6868 (N_6868,N_5726,N_5834);
or U6869 (N_6869,N_5266,N_5773);
nand U6870 (N_6870,N_5363,N_5950);
nand U6871 (N_6871,N_5435,N_5708);
nand U6872 (N_6872,N_5639,N_5072);
nor U6873 (N_6873,N_5698,N_5071);
nand U6874 (N_6874,N_5777,N_5304);
and U6875 (N_6875,N_5248,N_5189);
and U6876 (N_6876,N_5508,N_5620);
and U6877 (N_6877,N_5290,N_5197);
nand U6878 (N_6878,N_5325,N_5802);
and U6879 (N_6879,N_5302,N_5630);
and U6880 (N_6880,N_5242,N_5880);
xor U6881 (N_6881,N_5603,N_5319);
nand U6882 (N_6882,N_5379,N_5104);
or U6883 (N_6883,N_5715,N_5886);
nand U6884 (N_6884,N_5815,N_5249);
xnor U6885 (N_6885,N_5848,N_5761);
nor U6886 (N_6886,N_5821,N_5107);
nand U6887 (N_6887,N_5660,N_5902);
or U6888 (N_6888,N_5630,N_5594);
nand U6889 (N_6889,N_5927,N_5932);
nor U6890 (N_6890,N_5732,N_5240);
and U6891 (N_6891,N_5073,N_5396);
nor U6892 (N_6892,N_5669,N_5294);
or U6893 (N_6893,N_5234,N_5352);
or U6894 (N_6894,N_5996,N_5179);
nand U6895 (N_6895,N_5950,N_5222);
xnor U6896 (N_6896,N_5507,N_5068);
xor U6897 (N_6897,N_5734,N_5050);
xnor U6898 (N_6898,N_5044,N_5966);
or U6899 (N_6899,N_5713,N_5695);
nand U6900 (N_6900,N_5303,N_5908);
nand U6901 (N_6901,N_5384,N_5770);
nand U6902 (N_6902,N_5026,N_5645);
nor U6903 (N_6903,N_5986,N_5991);
and U6904 (N_6904,N_5609,N_5324);
nor U6905 (N_6905,N_5076,N_5073);
nor U6906 (N_6906,N_5947,N_5323);
nand U6907 (N_6907,N_5385,N_5077);
nand U6908 (N_6908,N_5552,N_5433);
or U6909 (N_6909,N_5779,N_5510);
nand U6910 (N_6910,N_5545,N_5411);
nor U6911 (N_6911,N_5027,N_5245);
or U6912 (N_6912,N_5721,N_5184);
nand U6913 (N_6913,N_5617,N_5526);
or U6914 (N_6914,N_5269,N_5121);
or U6915 (N_6915,N_5680,N_5298);
or U6916 (N_6916,N_5682,N_5509);
and U6917 (N_6917,N_5504,N_5116);
nand U6918 (N_6918,N_5661,N_5879);
xor U6919 (N_6919,N_5874,N_5861);
nand U6920 (N_6920,N_5575,N_5475);
nand U6921 (N_6921,N_5532,N_5602);
or U6922 (N_6922,N_5512,N_5385);
or U6923 (N_6923,N_5087,N_5229);
nand U6924 (N_6924,N_5175,N_5951);
nand U6925 (N_6925,N_5617,N_5806);
nand U6926 (N_6926,N_5378,N_5009);
nand U6927 (N_6927,N_5401,N_5732);
nor U6928 (N_6928,N_5600,N_5620);
nor U6929 (N_6929,N_5022,N_5793);
nand U6930 (N_6930,N_5672,N_5534);
or U6931 (N_6931,N_5108,N_5966);
or U6932 (N_6932,N_5715,N_5629);
and U6933 (N_6933,N_5206,N_5055);
nor U6934 (N_6934,N_5114,N_5276);
or U6935 (N_6935,N_5528,N_5184);
and U6936 (N_6936,N_5474,N_5363);
and U6937 (N_6937,N_5898,N_5494);
or U6938 (N_6938,N_5896,N_5824);
and U6939 (N_6939,N_5845,N_5423);
or U6940 (N_6940,N_5944,N_5580);
nor U6941 (N_6941,N_5565,N_5317);
and U6942 (N_6942,N_5565,N_5734);
xnor U6943 (N_6943,N_5747,N_5086);
nand U6944 (N_6944,N_5260,N_5496);
xor U6945 (N_6945,N_5240,N_5203);
xor U6946 (N_6946,N_5470,N_5989);
and U6947 (N_6947,N_5247,N_5557);
nor U6948 (N_6948,N_5608,N_5913);
or U6949 (N_6949,N_5017,N_5939);
or U6950 (N_6950,N_5266,N_5361);
nand U6951 (N_6951,N_5869,N_5257);
and U6952 (N_6952,N_5849,N_5902);
nor U6953 (N_6953,N_5251,N_5384);
and U6954 (N_6954,N_5609,N_5128);
nand U6955 (N_6955,N_5988,N_5886);
nor U6956 (N_6956,N_5467,N_5084);
nand U6957 (N_6957,N_5652,N_5952);
or U6958 (N_6958,N_5063,N_5945);
and U6959 (N_6959,N_5779,N_5414);
and U6960 (N_6960,N_5084,N_5345);
or U6961 (N_6961,N_5769,N_5245);
and U6962 (N_6962,N_5782,N_5508);
nor U6963 (N_6963,N_5964,N_5258);
or U6964 (N_6964,N_5165,N_5545);
xnor U6965 (N_6965,N_5294,N_5986);
xnor U6966 (N_6966,N_5838,N_5855);
or U6967 (N_6967,N_5751,N_5735);
and U6968 (N_6968,N_5458,N_5716);
or U6969 (N_6969,N_5106,N_5580);
and U6970 (N_6970,N_5960,N_5833);
nand U6971 (N_6971,N_5436,N_5328);
and U6972 (N_6972,N_5623,N_5437);
and U6973 (N_6973,N_5176,N_5696);
nor U6974 (N_6974,N_5103,N_5979);
nor U6975 (N_6975,N_5914,N_5058);
nor U6976 (N_6976,N_5076,N_5333);
nand U6977 (N_6977,N_5363,N_5169);
and U6978 (N_6978,N_5750,N_5762);
nand U6979 (N_6979,N_5919,N_5523);
xnor U6980 (N_6980,N_5111,N_5632);
nand U6981 (N_6981,N_5938,N_5037);
nor U6982 (N_6982,N_5387,N_5987);
nand U6983 (N_6983,N_5307,N_5958);
nand U6984 (N_6984,N_5937,N_5799);
xnor U6985 (N_6985,N_5260,N_5741);
nor U6986 (N_6986,N_5099,N_5743);
nor U6987 (N_6987,N_5583,N_5997);
and U6988 (N_6988,N_5650,N_5540);
or U6989 (N_6989,N_5421,N_5036);
and U6990 (N_6990,N_5969,N_5014);
nand U6991 (N_6991,N_5695,N_5469);
xnor U6992 (N_6992,N_5926,N_5423);
and U6993 (N_6993,N_5514,N_5129);
nor U6994 (N_6994,N_5960,N_5245);
nand U6995 (N_6995,N_5152,N_5604);
or U6996 (N_6996,N_5221,N_5587);
nand U6997 (N_6997,N_5529,N_5825);
nand U6998 (N_6998,N_5477,N_5415);
nor U6999 (N_6999,N_5392,N_5841);
xnor U7000 (N_7000,N_6549,N_6386);
nor U7001 (N_7001,N_6175,N_6626);
and U7002 (N_7002,N_6470,N_6266);
or U7003 (N_7003,N_6436,N_6090);
or U7004 (N_7004,N_6025,N_6352);
or U7005 (N_7005,N_6716,N_6151);
and U7006 (N_7006,N_6561,N_6127);
and U7007 (N_7007,N_6592,N_6607);
nand U7008 (N_7008,N_6268,N_6524);
and U7009 (N_7009,N_6860,N_6174);
or U7010 (N_7010,N_6357,N_6778);
nor U7011 (N_7011,N_6141,N_6371);
xor U7012 (N_7012,N_6558,N_6795);
and U7013 (N_7013,N_6509,N_6548);
or U7014 (N_7014,N_6741,N_6279);
nand U7015 (N_7015,N_6440,N_6672);
and U7016 (N_7016,N_6269,N_6805);
nor U7017 (N_7017,N_6432,N_6425);
and U7018 (N_7018,N_6941,N_6932);
nand U7019 (N_7019,N_6999,N_6753);
or U7020 (N_7020,N_6583,N_6823);
or U7021 (N_7021,N_6924,N_6820);
or U7022 (N_7022,N_6661,N_6343);
or U7023 (N_7023,N_6565,N_6764);
and U7024 (N_7024,N_6671,N_6770);
nand U7025 (N_7025,N_6086,N_6728);
or U7026 (N_7026,N_6465,N_6946);
and U7027 (N_7027,N_6633,N_6152);
xnor U7028 (N_7028,N_6663,N_6226);
nand U7029 (N_7029,N_6400,N_6028);
and U7030 (N_7030,N_6111,N_6701);
xor U7031 (N_7031,N_6767,N_6403);
and U7032 (N_7032,N_6375,N_6115);
or U7033 (N_7033,N_6620,N_6445);
nand U7034 (N_7034,N_6071,N_6362);
and U7035 (N_7035,N_6281,N_6718);
nand U7036 (N_7036,N_6433,N_6793);
nor U7037 (N_7037,N_6893,N_6879);
xor U7038 (N_7038,N_6298,N_6504);
nor U7039 (N_7039,N_6133,N_6950);
xnor U7040 (N_7040,N_6032,N_6194);
and U7041 (N_7041,N_6595,N_6132);
or U7042 (N_7042,N_6316,N_6218);
nand U7043 (N_7043,N_6255,N_6596);
or U7044 (N_7044,N_6388,N_6724);
nand U7045 (N_7045,N_6027,N_6965);
nand U7046 (N_7046,N_6895,N_6689);
nor U7047 (N_7047,N_6271,N_6599);
xnor U7048 (N_7048,N_6700,N_6117);
or U7049 (N_7049,N_6286,N_6979);
and U7050 (N_7050,N_6840,N_6444);
or U7051 (N_7051,N_6878,N_6587);
and U7052 (N_7052,N_6710,N_6825);
or U7053 (N_7053,N_6926,N_6001);
and U7054 (N_7054,N_6870,N_6872);
nor U7055 (N_7055,N_6101,N_6802);
and U7056 (N_7056,N_6815,N_6069);
or U7057 (N_7057,N_6976,N_6240);
or U7058 (N_7058,N_6105,N_6227);
or U7059 (N_7059,N_6260,N_6065);
and U7060 (N_7060,N_6336,N_6295);
and U7061 (N_7061,N_6106,N_6201);
nor U7062 (N_7062,N_6231,N_6665);
nor U7063 (N_7063,N_6717,N_6224);
nor U7064 (N_7064,N_6833,N_6173);
or U7065 (N_7065,N_6679,N_6521);
or U7066 (N_7066,N_6576,N_6505);
or U7067 (N_7067,N_6278,N_6828);
or U7068 (N_7068,N_6922,N_6986);
or U7069 (N_7069,N_6858,N_6322);
or U7070 (N_7070,N_6978,N_6988);
nor U7071 (N_7071,N_6076,N_6088);
or U7072 (N_7072,N_6157,N_6422);
nor U7073 (N_7073,N_6514,N_6450);
nand U7074 (N_7074,N_6915,N_6329);
nor U7075 (N_7075,N_6604,N_6670);
and U7076 (N_7076,N_6799,N_6265);
nand U7077 (N_7077,N_6159,N_6874);
nor U7078 (N_7078,N_6708,N_6387);
nand U7079 (N_7079,N_6373,N_6654);
and U7080 (N_7080,N_6367,N_6768);
and U7081 (N_7081,N_6258,N_6696);
or U7082 (N_7082,N_6569,N_6546);
or U7083 (N_7083,N_6059,N_6109);
nand U7084 (N_7084,N_6300,N_6560);
or U7085 (N_7085,N_6486,N_6649);
or U7086 (N_7086,N_6966,N_6248);
nor U7087 (N_7087,N_6784,N_6692);
or U7088 (N_7088,N_6472,N_6423);
nor U7089 (N_7089,N_6952,N_6601);
nand U7090 (N_7090,N_6676,N_6681);
or U7091 (N_7091,N_6538,N_6098);
or U7092 (N_7092,N_6089,N_6222);
nor U7093 (N_7093,N_6605,N_6317);
nor U7094 (N_7094,N_6099,N_6721);
or U7095 (N_7095,N_6917,N_6745);
and U7096 (N_7096,N_6094,N_6324);
or U7097 (N_7097,N_6808,N_6064);
or U7098 (N_7098,N_6232,N_6835);
nor U7099 (N_7099,N_6185,N_6913);
nand U7100 (N_7100,N_6519,N_6624);
nor U7101 (N_7101,N_6429,N_6301);
nor U7102 (N_7102,N_6360,N_6983);
nor U7103 (N_7103,N_6156,N_6199);
nand U7104 (N_7104,N_6190,N_6817);
or U7105 (N_7105,N_6206,N_6339);
or U7106 (N_7106,N_6837,N_6454);
nand U7107 (N_7107,N_6209,N_6121);
nor U7108 (N_7108,N_6903,N_6853);
nand U7109 (N_7109,N_6398,N_6553);
or U7110 (N_7110,N_6280,N_6167);
or U7111 (N_7111,N_6822,N_6714);
or U7112 (N_7112,N_6818,N_6123);
or U7113 (N_7113,N_6245,N_6068);
nor U7114 (N_7114,N_6215,N_6697);
nand U7115 (N_7115,N_6467,N_6192);
nand U7116 (N_7116,N_6930,N_6685);
or U7117 (N_7117,N_6600,N_6434);
and U7118 (N_7118,N_6276,N_6451);
nand U7119 (N_7119,N_6294,N_6237);
xnor U7120 (N_7120,N_6660,N_6200);
and U7121 (N_7121,N_6586,N_6761);
and U7122 (N_7122,N_6752,N_6987);
nand U7123 (N_7123,N_6408,N_6892);
and U7124 (N_7124,N_6330,N_6350);
or U7125 (N_7125,N_6902,N_6923);
and U7126 (N_7126,N_6730,N_6072);
or U7127 (N_7127,N_6040,N_6179);
or U7128 (N_7128,N_6918,N_6694);
and U7129 (N_7129,N_6613,N_6341);
and U7130 (N_7130,N_6426,N_6827);
xnor U7131 (N_7131,N_6968,N_6325);
or U7132 (N_7132,N_6742,N_6899);
and U7133 (N_7133,N_6308,N_6116);
nand U7134 (N_7134,N_6385,N_6220);
nand U7135 (N_7135,N_6756,N_6442);
nor U7136 (N_7136,N_6533,N_6198);
nor U7137 (N_7137,N_6368,N_6452);
nand U7138 (N_7138,N_6614,N_6811);
and U7139 (N_7139,N_6079,N_6674);
and U7140 (N_7140,N_6120,N_6490);
xnor U7141 (N_7141,N_6551,N_6559);
or U7142 (N_7142,N_6698,N_6180);
and U7143 (N_7143,N_6137,N_6460);
nand U7144 (N_7144,N_6956,N_6499);
and U7145 (N_7145,N_6142,N_6766);
or U7146 (N_7146,N_6735,N_6464);
nor U7147 (N_7147,N_6901,N_6568);
and U7148 (N_7148,N_6187,N_6990);
and U7149 (N_7149,N_6774,N_6038);
or U7150 (N_7150,N_6898,N_6849);
and U7151 (N_7151,N_6830,N_6480);
or U7152 (N_7152,N_6230,N_6113);
nor U7153 (N_7153,N_6292,N_6949);
nor U7154 (N_7154,N_6847,N_6402);
xor U7155 (N_7155,N_6256,N_6522);
or U7156 (N_7156,N_6975,N_6481);
nor U7157 (N_7157,N_6036,N_6335);
nor U7158 (N_7158,N_6342,N_6338);
nor U7159 (N_7159,N_6695,N_6618);
nor U7160 (N_7160,N_6318,N_6951);
and U7161 (N_7161,N_6736,N_6684);
nor U7162 (N_7162,N_6852,N_6829);
nor U7163 (N_7163,N_6469,N_6729);
nand U7164 (N_7164,N_6877,N_6556);
or U7165 (N_7165,N_6969,N_6589);
nand U7166 (N_7166,N_6542,N_6639);
or U7167 (N_7167,N_6772,N_6683);
nand U7168 (N_7168,N_6435,N_6437);
or U7169 (N_7169,N_6785,N_6798);
or U7170 (N_7170,N_6520,N_6471);
nand U7171 (N_7171,N_6501,N_6290);
and U7172 (N_7172,N_6940,N_6331);
xnor U7173 (N_7173,N_6916,N_6967);
and U7174 (N_7174,N_6854,N_6372);
or U7175 (N_7175,N_6263,N_6821);
or U7176 (N_7176,N_6333,N_6616);
nor U7177 (N_7177,N_6500,N_6719);
nand U7178 (N_7178,N_6557,N_6925);
or U7179 (N_7179,N_6270,N_6351);
nor U7180 (N_7180,N_6751,N_6103);
or U7181 (N_7181,N_6091,N_6703);
or U7182 (N_7182,N_6783,N_6377);
xor U7183 (N_7183,N_6029,N_6886);
nand U7184 (N_7184,N_6163,N_6196);
nor U7185 (N_7185,N_6773,N_6045);
nand U7186 (N_7186,N_6732,N_6779);
xnor U7187 (N_7187,N_6138,N_6236);
or U7188 (N_7188,N_6702,N_6021);
or U7189 (N_7189,N_6075,N_6970);
xor U7190 (N_7190,N_6381,N_6347);
nor U7191 (N_7191,N_6754,N_6489);
or U7192 (N_7192,N_6758,N_6632);
and U7193 (N_7193,N_6836,N_6713);
nor U7194 (N_7194,N_6800,N_6527);
or U7195 (N_7195,N_6739,N_6356);
nand U7196 (N_7196,N_6482,N_6042);
and U7197 (N_7197,N_6037,N_6512);
and U7198 (N_7198,N_6535,N_6516);
xor U7199 (N_7199,N_6355,N_6876);
and U7200 (N_7200,N_6733,N_6114);
or U7201 (N_7201,N_6744,N_6246);
nand U7202 (N_7202,N_6740,N_6747);
nor U7203 (N_7203,N_6593,N_6792);
nand U7204 (N_7204,N_6746,N_6731);
nand U7205 (N_7205,N_6394,N_6439);
or U7206 (N_7206,N_6993,N_6931);
nor U7207 (N_7207,N_6484,N_6296);
xor U7208 (N_7208,N_6707,N_6315);
xor U7209 (N_7209,N_6030,N_6938);
and U7210 (N_7210,N_6962,N_6657);
nand U7211 (N_7211,N_6378,N_6291);
nand U7212 (N_7212,N_6653,N_6875);
and U7213 (N_7213,N_6645,N_6004);
or U7214 (N_7214,N_6264,N_6312);
xor U7215 (N_7215,N_6585,N_6345);
or U7216 (N_7216,N_6989,N_6711);
xor U7217 (N_7217,N_6927,N_6018);
or U7218 (N_7218,N_6659,N_6909);
nand U7219 (N_7219,N_6046,N_6310);
nand U7220 (N_7220,N_6992,N_6643);
xor U7221 (N_7221,N_6850,N_6225);
nand U7222 (N_7222,N_6478,N_6320);
and U7223 (N_7223,N_6349,N_6982);
nor U7224 (N_7224,N_6544,N_6885);
and U7225 (N_7225,N_6513,N_6788);
and U7226 (N_7226,N_6313,N_6189);
or U7227 (N_7227,N_6985,N_6051);
nand U7228 (N_7228,N_6508,N_6994);
nor U7229 (N_7229,N_6223,N_6666);
or U7230 (N_7230,N_6497,N_6762);
nor U7231 (N_7231,N_6384,N_6459);
nand U7232 (N_7232,N_6677,N_6699);
xnor U7233 (N_7233,N_6640,N_6831);
or U7234 (N_7234,N_6483,N_6182);
xnor U7235 (N_7235,N_6996,N_6297);
nor U7236 (N_7236,N_6498,N_6130);
or U7237 (N_7237,N_6203,N_6528);
nand U7238 (N_7238,N_6181,N_6407);
nand U7239 (N_7239,N_6619,N_6617);
nor U7240 (N_7240,N_6143,N_6705);
xor U7241 (N_7241,N_6477,N_6789);
and U7242 (N_7242,N_6539,N_6369);
xnor U7243 (N_7243,N_6963,N_6393);
or U7244 (N_7244,N_6244,N_6158);
nand U7245 (N_7245,N_6272,N_6406);
nand U7246 (N_7246,N_6379,N_6397);
and U7247 (N_7247,N_6552,N_6153);
nand U7248 (N_7248,N_6267,N_6326);
nor U7249 (N_7249,N_6005,N_6202);
nor U7250 (N_7250,N_6578,N_6933);
nor U7251 (N_7251,N_6612,N_6413);
nor U7252 (N_7252,N_6087,N_6590);
xor U7253 (N_7253,N_6610,N_6843);
and U7254 (N_7254,N_6636,N_6841);
xor U7255 (N_7255,N_6083,N_6547);
or U7256 (N_7256,N_6016,N_6419);
or U7257 (N_7257,N_6826,N_6488);
and U7258 (N_7258,N_6573,N_6449);
or U7259 (N_7259,N_6581,N_6247);
nor U7260 (N_7260,N_6166,N_6374);
xor U7261 (N_7261,N_6566,N_6957);
and U7262 (N_7262,N_6078,N_6842);
and U7263 (N_7263,N_6939,N_6791);
or U7264 (N_7264,N_6212,N_6077);
or U7265 (N_7265,N_6491,N_6602);
nand U7266 (N_7266,N_6074,N_6184);
nand U7267 (N_7267,N_6609,N_6461);
nand U7268 (N_7268,N_6009,N_6564);
and U7269 (N_7269,N_6466,N_6024);
and U7270 (N_7270,N_6582,N_6006);
xnor U7271 (N_7271,N_6107,N_6282);
xnor U7272 (N_7272,N_6288,N_6446);
and U7273 (N_7273,N_6060,N_6757);
nor U7274 (N_7274,N_6652,N_6502);
or U7275 (N_7275,N_6210,N_6096);
xor U7276 (N_7276,N_6093,N_6399);
or U7277 (N_7277,N_6543,N_6862);
nand U7278 (N_7278,N_6855,N_6139);
nor U7279 (N_7279,N_6346,N_6658);
xnor U7280 (N_7280,N_6363,N_6412);
or U7281 (N_7281,N_6848,N_6936);
xnor U7282 (N_7282,N_6554,N_6814);
or U7283 (N_7283,N_6887,N_6851);
nor U7284 (N_7284,N_6034,N_6252);
nand U7285 (N_7285,N_6813,N_6391);
nor U7286 (N_7286,N_6536,N_6673);
and U7287 (N_7287,N_6254,N_6550);
and U7288 (N_7288,N_6238,N_6463);
and U7289 (N_7289,N_6052,N_6311);
and U7290 (N_7290,N_6907,N_6353);
and U7291 (N_7291,N_6358,N_6305);
and U7292 (N_7292,N_6682,N_6906);
nand U7293 (N_7293,N_6631,N_6039);
xor U7294 (N_7294,N_6914,N_6606);
or U7295 (N_7295,N_6066,N_6904);
nor U7296 (N_7296,N_6404,N_6910);
nor U7297 (N_7297,N_6124,N_6284);
nand U7298 (N_7298,N_6621,N_6920);
nor U7299 (N_7299,N_6912,N_6627);
nor U7300 (N_7300,N_6421,N_6574);
or U7301 (N_7301,N_6947,N_6690);
or U7302 (N_7302,N_6380,N_6390);
and U7303 (N_7303,N_6468,N_6518);
nand U7304 (N_7304,N_6262,N_6834);
and U7305 (N_7305,N_6642,N_6438);
nand U7306 (N_7306,N_6867,N_6797);
and U7307 (N_7307,N_6871,N_6819);
and U7308 (N_7308,N_6641,N_6447);
nand U7309 (N_7309,N_6646,N_6479);
and U7310 (N_7310,N_6061,N_6759);
and U7311 (N_7311,N_6883,N_6948);
xnor U7312 (N_7312,N_6104,N_6344);
and U7313 (N_7313,N_6934,N_6882);
xnor U7314 (N_7314,N_6108,N_6134);
nor U7315 (N_7315,N_6242,N_6944);
nor U7316 (N_7316,N_6958,N_6168);
or U7317 (N_7317,N_6487,N_6002);
nor U7318 (N_7318,N_6884,N_6726);
or U7319 (N_7319,N_6801,N_6003);
nand U7320 (N_7320,N_6580,N_6525);
xnor U7321 (N_7321,N_6890,N_6796);
or U7322 (N_7322,N_6598,N_6303);
nor U7323 (N_7323,N_6998,N_6361);
and U7324 (N_7324,N_6176,N_6044);
nor U7325 (N_7325,N_6015,N_6678);
nand U7326 (N_7326,N_6687,N_6748);
and U7327 (N_7327,N_6251,N_6007);
nand U7328 (N_7328,N_6973,N_6769);
or U7329 (N_7329,N_6763,N_6188);
and U7330 (N_7330,N_6328,N_6457);
nand U7331 (N_7331,N_6473,N_6416);
and U7332 (N_7332,N_6359,N_6662);
nand U7333 (N_7333,N_6327,N_6804);
nand U7334 (N_7334,N_6935,N_6888);
nor U7335 (N_7335,N_6638,N_6129);
nand U7336 (N_7336,N_6891,N_6366);
or U7337 (N_7337,N_6495,N_6119);
and U7338 (N_7338,N_6810,N_6715);
nand U7339 (N_7339,N_6844,N_6462);
nor U7340 (N_7340,N_6110,N_6727);
or U7341 (N_7341,N_6147,N_6889);
nor U7342 (N_7342,N_6688,N_6896);
and U7343 (N_7343,N_6122,N_6628);
and U7344 (N_7344,N_6803,N_6567);
nor U7345 (N_7345,N_6974,N_6980);
or U7346 (N_7346,N_6146,N_6562);
nor U7347 (N_7347,N_6782,N_6971);
nand U7348 (N_7348,N_6775,N_6706);
nor U7349 (N_7349,N_6510,N_6577);
xor U7350 (N_7350,N_6790,N_6031);
nor U7351 (N_7351,N_6972,N_6228);
and U7352 (N_7352,N_6984,N_6997);
and U7353 (N_7353,N_6430,N_6507);
nand U7354 (N_7354,N_6165,N_6453);
xnor U7355 (N_7355,N_6208,N_6503);
and U7356 (N_7356,N_6160,N_6396);
nor U7357 (N_7357,N_6794,N_6526);
and U7358 (N_7358,N_6299,N_6597);
nand U7359 (N_7359,N_6523,N_6048);
and U7360 (N_7360,N_6364,N_6073);
and U7361 (N_7361,N_6304,N_6555);
xnor U7362 (N_7362,N_6017,N_6749);
nand U7363 (N_7363,N_6370,N_6722);
nor U7364 (N_7364,N_6410,N_6014);
xor U7365 (N_7365,N_6420,N_6136);
nor U7366 (N_7366,N_6448,N_6140);
nand U7367 (N_7367,N_6629,N_6149);
nor U7368 (N_7368,N_6217,N_6026);
nor U7369 (N_7369,N_6100,N_6171);
or U7370 (N_7370,N_6053,N_6771);
nand U7371 (N_7371,N_6492,N_6161);
nand U7372 (N_7372,N_6411,N_6234);
nand U7373 (N_7373,N_6824,N_6035);
or U7374 (N_7374,N_6275,N_6475);
nor U7375 (N_7375,N_6863,N_6084);
and U7376 (N_7376,N_6287,N_6183);
or U7377 (N_7377,N_6257,N_6953);
and U7378 (N_7378,N_6859,N_6214);
and U7379 (N_7379,N_6591,N_6022);
nand U7380 (N_7380,N_6418,N_6712);
nand U7381 (N_7381,N_6704,N_6650);
and U7382 (N_7382,N_6954,N_6424);
or U7383 (N_7383,N_6213,N_6162);
and U7384 (N_7384,N_6097,N_6013);
and U7385 (N_7385,N_6250,N_6443);
nand U7386 (N_7386,N_6723,N_6680);
nand U7387 (N_7387,N_6243,N_6937);
xnor U7388 (N_7388,N_6058,N_6102);
and U7389 (N_7389,N_6431,N_6047);
or U7390 (N_7390,N_6995,N_6177);
nand U7391 (N_7391,N_6839,N_6274);
xnor U7392 (N_7392,N_6807,N_6081);
and U7393 (N_7393,N_6376,N_6229);
nor U7394 (N_7394,N_6063,N_6169);
or U7395 (N_7395,N_6506,N_6570);
and U7396 (N_7396,N_6959,N_6321);
or U7397 (N_7397,N_6530,N_6865);
and U7398 (N_7398,N_6427,N_6382);
and U7399 (N_7399,N_6144,N_6571);
and U7400 (N_7400,N_6579,N_6055);
and U7401 (N_7401,N_6409,N_6456);
or U7402 (N_7402,N_6531,N_6128);
nand U7403 (N_7403,N_6720,N_6725);
nand U7404 (N_7404,N_6894,N_6118);
nor U7405 (N_7405,N_6955,N_6981);
nand U7406 (N_7406,N_6365,N_6928);
nor U7407 (N_7407,N_6233,N_6857);
xnor U7408 (N_7408,N_6337,N_6603);
nand U7409 (N_7409,N_6532,N_6383);
nand U7410 (N_7410,N_6145,N_6125);
or U7411 (N_7411,N_6277,N_6777);
nand U7412 (N_7412,N_6709,N_6669);
or U7413 (N_7413,N_6816,N_6611);
xor U7414 (N_7414,N_6511,N_6178);
nand U7415 (N_7415,N_6261,N_6354);
or U7416 (N_7416,N_6049,N_6838);
xor U7417 (N_7417,N_6881,N_6537);
xor U7418 (N_7418,N_6332,N_6991);
nand U7419 (N_7419,N_6070,N_6389);
nand U7420 (N_7420,N_6743,N_6170);
and U7421 (N_7421,N_6691,N_6575);
or U7422 (N_7422,N_6622,N_6219);
and U7423 (N_7423,N_6415,N_6942);
nor U7424 (N_7424,N_6655,N_6082);
nor U7425 (N_7425,N_6921,N_6786);
and U7426 (N_7426,N_6253,N_6832);
nand U7427 (N_7427,N_6873,N_6960);
nand U7428 (N_7428,N_6588,N_6405);
nor U7429 (N_7429,N_6781,N_6092);
xor U7430 (N_7430,N_6738,N_6126);
or U7431 (N_7431,N_6293,N_6594);
or U7432 (N_7432,N_6515,N_6540);
nand U7433 (N_7433,N_6647,N_6428);
nor U7434 (N_7434,N_6476,N_6235);
or U7435 (N_7435,N_6734,N_6534);
or U7436 (N_7436,N_6905,N_6529);
nor U7437 (N_7437,N_6010,N_6693);
and U7438 (N_7438,N_6191,N_6458);
xor U7439 (N_7439,N_6812,N_6307);
nand U7440 (N_7440,N_6545,N_6644);
and U7441 (N_7441,N_6765,N_6289);
nor U7442 (N_7442,N_6041,N_6776);
nand U7443 (N_7443,N_6911,N_6750);
nor U7444 (N_7444,N_6634,N_6760);
nor U7445 (N_7445,N_6787,N_6216);
and U7446 (N_7446,N_6067,N_6417);
and U7447 (N_7447,N_6155,N_6334);
or U7448 (N_7448,N_6000,N_6929);
nand U7449 (N_7449,N_6241,N_6302);
nor U7450 (N_7450,N_6668,N_6864);
nor U7451 (N_7451,N_6085,N_6011);
xnor U7452 (N_7452,N_6211,N_6135);
and U7453 (N_7453,N_6249,N_6056);
or U7454 (N_7454,N_6964,N_6977);
nor U7455 (N_7455,N_6474,N_6204);
nor U7456 (N_7456,N_6414,N_6637);
or U7457 (N_7457,N_6493,N_6205);
nand U7458 (N_7458,N_6861,N_6008);
nor U7459 (N_7459,N_6572,N_6664);
nor U7460 (N_7460,N_6148,N_6020);
nor U7461 (N_7461,N_6285,N_6755);
and U7462 (N_7462,N_6150,N_6667);
and U7463 (N_7463,N_6319,N_6283);
nor U7464 (N_7464,N_6080,N_6656);
nand U7465 (N_7465,N_6164,N_6455);
and U7466 (N_7466,N_6625,N_6172);
or U7467 (N_7467,N_6259,N_6441);
or U7468 (N_7468,N_6395,N_6623);
nor U7469 (N_7469,N_6239,N_6401);
and U7470 (N_7470,N_6323,N_6496);
nand U7471 (N_7471,N_6309,N_6880);
nor U7472 (N_7472,N_6054,N_6868);
or U7473 (N_7473,N_6207,N_6340);
nand U7474 (N_7474,N_6062,N_6651);
xnor U7475 (N_7475,N_6897,N_6186);
nand U7476 (N_7476,N_6945,N_6517);
nand U7477 (N_7477,N_6869,N_6635);
and U7478 (N_7478,N_6154,N_6648);
nor U7479 (N_7479,N_6193,N_6846);
or U7480 (N_7480,N_6541,N_6615);
nand U7481 (N_7481,N_6908,N_6112);
nor U7482 (N_7482,N_6392,N_6095);
and U7483 (N_7483,N_6608,N_6866);
and U7484 (N_7484,N_6900,N_6809);
nand U7485 (N_7485,N_6221,N_6012);
and U7486 (N_7486,N_6043,N_6057);
nor U7487 (N_7487,N_6584,N_6050);
or U7488 (N_7488,N_6919,N_6686);
or U7489 (N_7489,N_6314,N_6961);
nand U7490 (N_7490,N_6197,N_6023);
nand U7491 (N_7491,N_6675,N_6780);
and U7492 (N_7492,N_6348,N_6273);
nor U7493 (N_7493,N_6630,N_6806);
and U7494 (N_7494,N_6943,N_6195);
xor U7495 (N_7495,N_6737,N_6019);
or U7496 (N_7496,N_6856,N_6845);
and U7497 (N_7497,N_6494,N_6033);
nand U7498 (N_7498,N_6306,N_6563);
nor U7499 (N_7499,N_6131,N_6485);
nand U7500 (N_7500,N_6785,N_6541);
nor U7501 (N_7501,N_6197,N_6483);
xor U7502 (N_7502,N_6344,N_6476);
nor U7503 (N_7503,N_6192,N_6708);
nor U7504 (N_7504,N_6821,N_6946);
xor U7505 (N_7505,N_6217,N_6561);
or U7506 (N_7506,N_6188,N_6286);
or U7507 (N_7507,N_6189,N_6127);
or U7508 (N_7508,N_6733,N_6052);
nand U7509 (N_7509,N_6527,N_6692);
nor U7510 (N_7510,N_6088,N_6839);
and U7511 (N_7511,N_6874,N_6651);
nor U7512 (N_7512,N_6293,N_6526);
and U7513 (N_7513,N_6833,N_6465);
and U7514 (N_7514,N_6973,N_6803);
or U7515 (N_7515,N_6215,N_6368);
or U7516 (N_7516,N_6456,N_6692);
and U7517 (N_7517,N_6978,N_6334);
xor U7518 (N_7518,N_6554,N_6200);
nand U7519 (N_7519,N_6603,N_6953);
xnor U7520 (N_7520,N_6238,N_6680);
nand U7521 (N_7521,N_6039,N_6032);
and U7522 (N_7522,N_6796,N_6044);
and U7523 (N_7523,N_6696,N_6289);
and U7524 (N_7524,N_6825,N_6441);
nor U7525 (N_7525,N_6445,N_6951);
xor U7526 (N_7526,N_6711,N_6652);
or U7527 (N_7527,N_6827,N_6881);
nand U7528 (N_7528,N_6758,N_6795);
or U7529 (N_7529,N_6726,N_6179);
nand U7530 (N_7530,N_6551,N_6722);
nand U7531 (N_7531,N_6995,N_6491);
nor U7532 (N_7532,N_6138,N_6389);
nand U7533 (N_7533,N_6876,N_6490);
or U7534 (N_7534,N_6886,N_6055);
nor U7535 (N_7535,N_6679,N_6407);
nor U7536 (N_7536,N_6176,N_6278);
and U7537 (N_7537,N_6296,N_6083);
or U7538 (N_7538,N_6298,N_6906);
nand U7539 (N_7539,N_6744,N_6881);
or U7540 (N_7540,N_6116,N_6194);
nor U7541 (N_7541,N_6910,N_6879);
and U7542 (N_7542,N_6135,N_6614);
or U7543 (N_7543,N_6803,N_6870);
or U7544 (N_7544,N_6293,N_6776);
or U7545 (N_7545,N_6320,N_6743);
nand U7546 (N_7546,N_6601,N_6244);
nor U7547 (N_7547,N_6859,N_6617);
and U7548 (N_7548,N_6174,N_6020);
nand U7549 (N_7549,N_6452,N_6618);
or U7550 (N_7550,N_6611,N_6267);
and U7551 (N_7551,N_6829,N_6419);
or U7552 (N_7552,N_6676,N_6002);
nand U7553 (N_7553,N_6796,N_6864);
nor U7554 (N_7554,N_6671,N_6991);
and U7555 (N_7555,N_6256,N_6801);
or U7556 (N_7556,N_6173,N_6816);
nor U7557 (N_7557,N_6039,N_6170);
nand U7558 (N_7558,N_6136,N_6740);
nor U7559 (N_7559,N_6341,N_6570);
nand U7560 (N_7560,N_6681,N_6860);
or U7561 (N_7561,N_6856,N_6017);
nand U7562 (N_7562,N_6797,N_6816);
and U7563 (N_7563,N_6400,N_6752);
xor U7564 (N_7564,N_6981,N_6484);
and U7565 (N_7565,N_6158,N_6420);
xor U7566 (N_7566,N_6345,N_6646);
nand U7567 (N_7567,N_6580,N_6433);
nand U7568 (N_7568,N_6649,N_6571);
or U7569 (N_7569,N_6646,N_6749);
and U7570 (N_7570,N_6272,N_6329);
xnor U7571 (N_7571,N_6576,N_6957);
nor U7572 (N_7572,N_6054,N_6970);
or U7573 (N_7573,N_6071,N_6771);
and U7574 (N_7574,N_6890,N_6059);
and U7575 (N_7575,N_6966,N_6337);
and U7576 (N_7576,N_6648,N_6782);
nor U7577 (N_7577,N_6416,N_6386);
and U7578 (N_7578,N_6383,N_6705);
nand U7579 (N_7579,N_6388,N_6854);
nand U7580 (N_7580,N_6558,N_6480);
nand U7581 (N_7581,N_6350,N_6447);
and U7582 (N_7582,N_6095,N_6210);
and U7583 (N_7583,N_6926,N_6443);
nand U7584 (N_7584,N_6885,N_6658);
and U7585 (N_7585,N_6912,N_6496);
nand U7586 (N_7586,N_6201,N_6276);
nand U7587 (N_7587,N_6598,N_6825);
and U7588 (N_7588,N_6363,N_6703);
nand U7589 (N_7589,N_6924,N_6090);
nor U7590 (N_7590,N_6122,N_6892);
nor U7591 (N_7591,N_6662,N_6861);
and U7592 (N_7592,N_6516,N_6567);
and U7593 (N_7593,N_6996,N_6121);
or U7594 (N_7594,N_6125,N_6260);
nor U7595 (N_7595,N_6651,N_6885);
nand U7596 (N_7596,N_6153,N_6360);
or U7597 (N_7597,N_6712,N_6325);
and U7598 (N_7598,N_6253,N_6330);
or U7599 (N_7599,N_6317,N_6702);
or U7600 (N_7600,N_6724,N_6683);
and U7601 (N_7601,N_6848,N_6366);
or U7602 (N_7602,N_6739,N_6211);
or U7603 (N_7603,N_6228,N_6708);
or U7604 (N_7604,N_6288,N_6411);
or U7605 (N_7605,N_6055,N_6506);
and U7606 (N_7606,N_6776,N_6977);
or U7607 (N_7607,N_6132,N_6553);
or U7608 (N_7608,N_6299,N_6581);
or U7609 (N_7609,N_6914,N_6560);
nor U7610 (N_7610,N_6688,N_6173);
nand U7611 (N_7611,N_6834,N_6473);
nand U7612 (N_7612,N_6136,N_6156);
xor U7613 (N_7613,N_6777,N_6253);
xnor U7614 (N_7614,N_6054,N_6554);
and U7615 (N_7615,N_6989,N_6789);
or U7616 (N_7616,N_6925,N_6830);
xor U7617 (N_7617,N_6705,N_6881);
nor U7618 (N_7618,N_6375,N_6645);
and U7619 (N_7619,N_6843,N_6364);
or U7620 (N_7620,N_6265,N_6681);
nand U7621 (N_7621,N_6502,N_6097);
and U7622 (N_7622,N_6578,N_6863);
and U7623 (N_7623,N_6628,N_6102);
or U7624 (N_7624,N_6677,N_6555);
nand U7625 (N_7625,N_6367,N_6052);
or U7626 (N_7626,N_6446,N_6738);
nand U7627 (N_7627,N_6261,N_6144);
or U7628 (N_7628,N_6115,N_6567);
or U7629 (N_7629,N_6126,N_6225);
xnor U7630 (N_7630,N_6678,N_6895);
or U7631 (N_7631,N_6688,N_6648);
nor U7632 (N_7632,N_6895,N_6792);
nand U7633 (N_7633,N_6320,N_6234);
xnor U7634 (N_7634,N_6575,N_6971);
and U7635 (N_7635,N_6249,N_6267);
xor U7636 (N_7636,N_6213,N_6283);
xnor U7637 (N_7637,N_6207,N_6914);
or U7638 (N_7638,N_6130,N_6745);
nand U7639 (N_7639,N_6808,N_6020);
nor U7640 (N_7640,N_6828,N_6501);
nor U7641 (N_7641,N_6832,N_6995);
and U7642 (N_7642,N_6269,N_6534);
nand U7643 (N_7643,N_6927,N_6824);
or U7644 (N_7644,N_6656,N_6580);
nor U7645 (N_7645,N_6957,N_6727);
nor U7646 (N_7646,N_6366,N_6119);
or U7647 (N_7647,N_6381,N_6202);
nand U7648 (N_7648,N_6952,N_6967);
nand U7649 (N_7649,N_6694,N_6270);
xor U7650 (N_7650,N_6658,N_6165);
or U7651 (N_7651,N_6707,N_6531);
or U7652 (N_7652,N_6517,N_6923);
and U7653 (N_7653,N_6080,N_6472);
or U7654 (N_7654,N_6093,N_6244);
or U7655 (N_7655,N_6020,N_6033);
xor U7656 (N_7656,N_6798,N_6897);
and U7657 (N_7657,N_6242,N_6360);
nand U7658 (N_7658,N_6779,N_6026);
nand U7659 (N_7659,N_6062,N_6160);
and U7660 (N_7660,N_6667,N_6375);
xor U7661 (N_7661,N_6594,N_6087);
and U7662 (N_7662,N_6946,N_6966);
nor U7663 (N_7663,N_6252,N_6880);
xnor U7664 (N_7664,N_6117,N_6383);
nor U7665 (N_7665,N_6051,N_6232);
and U7666 (N_7666,N_6331,N_6009);
xor U7667 (N_7667,N_6775,N_6203);
xnor U7668 (N_7668,N_6082,N_6043);
and U7669 (N_7669,N_6216,N_6278);
nand U7670 (N_7670,N_6849,N_6214);
or U7671 (N_7671,N_6450,N_6778);
nor U7672 (N_7672,N_6544,N_6246);
or U7673 (N_7673,N_6535,N_6834);
and U7674 (N_7674,N_6613,N_6959);
and U7675 (N_7675,N_6392,N_6477);
nand U7676 (N_7676,N_6314,N_6196);
or U7677 (N_7677,N_6112,N_6022);
nor U7678 (N_7678,N_6388,N_6594);
and U7679 (N_7679,N_6944,N_6088);
or U7680 (N_7680,N_6742,N_6632);
nor U7681 (N_7681,N_6949,N_6226);
and U7682 (N_7682,N_6287,N_6299);
nor U7683 (N_7683,N_6809,N_6175);
nand U7684 (N_7684,N_6962,N_6391);
nor U7685 (N_7685,N_6177,N_6979);
or U7686 (N_7686,N_6002,N_6120);
or U7687 (N_7687,N_6225,N_6191);
nand U7688 (N_7688,N_6801,N_6282);
and U7689 (N_7689,N_6951,N_6783);
and U7690 (N_7690,N_6693,N_6737);
nand U7691 (N_7691,N_6425,N_6562);
and U7692 (N_7692,N_6758,N_6116);
and U7693 (N_7693,N_6841,N_6521);
xor U7694 (N_7694,N_6353,N_6348);
xnor U7695 (N_7695,N_6210,N_6075);
nor U7696 (N_7696,N_6407,N_6009);
nand U7697 (N_7697,N_6679,N_6329);
nand U7698 (N_7698,N_6925,N_6597);
nor U7699 (N_7699,N_6951,N_6145);
nand U7700 (N_7700,N_6565,N_6134);
and U7701 (N_7701,N_6144,N_6746);
and U7702 (N_7702,N_6296,N_6641);
nor U7703 (N_7703,N_6824,N_6578);
nand U7704 (N_7704,N_6358,N_6063);
or U7705 (N_7705,N_6702,N_6966);
nand U7706 (N_7706,N_6457,N_6326);
or U7707 (N_7707,N_6623,N_6068);
nand U7708 (N_7708,N_6024,N_6410);
and U7709 (N_7709,N_6053,N_6719);
and U7710 (N_7710,N_6856,N_6267);
nand U7711 (N_7711,N_6566,N_6577);
nor U7712 (N_7712,N_6834,N_6918);
and U7713 (N_7713,N_6910,N_6747);
xnor U7714 (N_7714,N_6279,N_6798);
or U7715 (N_7715,N_6181,N_6397);
nor U7716 (N_7716,N_6380,N_6637);
nor U7717 (N_7717,N_6360,N_6365);
xor U7718 (N_7718,N_6259,N_6761);
or U7719 (N_7719,N_6073,N_6042);
nor U7720 (N_7720,N_6634,N_6693);
or U7721 (N_7721,N_6891,N_6032);
nor U7722 (N_7722,N_6023,N_6578);
nor U7723 (N_7723,N_6704,N_6551);
and U7724 (N_7724,N_6452,N_6313);
nand U7725 (N_7725,N_6304,N_6073);
nand U7726 (N_7726,N_6907,N_6041);
xnor U7727 (N_7727,N_6912,N_6632);
and U7728 (N_7728,N_6827,N_6277);
nand U7729 (N_7729,N_6312,N_6704);
and U7730 (N_7730,N_6010,N_6564);
nand U7731 (N_7731,N_6958,N_6002);
nand U7732 (N_7732,N_6487,N_6773);
nor U7733 (N_7733,N_6741,N_6961);
nor U7734 (N_7734,N_6851,N_6073);
or U7735 (N_7735,N_6265,N_6955);
nand U7736 (N_7736,N_6737,N_6061);
xor U7737 (N_7737,N_6936,N_6817);
nand U7738 (N_7738,N_6970,N_6555);
nand U7739 (N_7739,N_6754,N_6192);
and U7740 (N_7740,N_6025,N_6133);
or U7741 (N_7741,N_6868,N_6247);
nor U7742 (N_7742,N_6244,N_6740);
nand U7743 (N_7743,N_6041,N_6952);
nor U7744 (N_7744,N_6547,N_6396);
nand U7745 (N_7745,N_6417,N_6108);
nor U7746 (N_7746,N_6139,N_6985);
nor U7747 (N_7747,N_6532,N_6111);
and U7748 (N_7748,N_6731,N_6435);
nand U7749 (N_7749,N_6837,N_6504);
nor U7750 (N_7750,N_6536,N_6905);
nor U7751 (N_7751,N_6804,N_6187);
or U7752 (N_7752,N_6056,N_6008);
xor U7753 (N_7753,N_6147,N_6214);
and U7754 (N_7754,N_6207,N_6740);
nand U7755 (N_7755,N_6568,N_6837);
and U7756 (N_7756,N_6262,N_6086);
and U7757 (N_7757,N_6571,N_6594);
and U7758 (N_7758,N_6895,N_6816);
nor U7759 (N_7759,N_6583,N_6800);
xnor U7760 (N_7760,N_6517,N_6844);
nand U7761 (N_7761,N_6284,N_6348);
and U7762 (N_7762,N_6680,N_6227);
xor U7763 (N_7763,N_6578,N_6138);
and U7764 (N_7764,N_6301,N_6534);
and U7765 (N_7765,N_6460,N_6458);
nand U7766 (N_7766,N_6485,N_6024);
nand U7767 (N_7767,N_6144,N_6697);
or U7768 (N_7768,N_6354,N_6554);
nand U7769 (N_7769,N_6090,N_6575);
nand U7770 (N_7770,N_6213,N_6201);
nand U7771 (N_7771,N_6057,N_6163);
and U7772 (N_7772,N_6514,N_6925);
nand U7773 (N_7773,N_6445,N_6779);
nand U7774 (N_7774,N_6983,N_6542);
nor U7775 (N_7775,N_6664,N_6039);
nor U7776 (N_7776,N_6214,N_6699);
nor U7777 (N_7777,N_6000,N_6546);
or U7778 (N_7778,N_6114,N_6391);
and U7779 (N_7779,N_6600,N_6321);
nor U7780 (N_7780,N_6319,N_6590);
nand U7781 (N_7781,N_6317,N_6668);
xor U7782 (N_7782,N_6814,N_6436);
nand U7783 (N_7783,N_6890,N_6640);
and U7784 (N_7784,N_6363,N_6023);
or U7785 (N_7785,N_6281,N_6152);
nor U7786 (N_7786,N_6891,N_6591);
nand U7787 (N_7787,N_6171,N_6700);
xnor U7788 (N_7788,N_6915,N_6754);
nor U7789 (N_7789,N_6991,N_6846);
nor U7790 (N_7790,N_6035,N_6172);
nor U7791 (N_7791,N_6226,N_6198);
or U7792 (N_7792,N_6306,N_6600);
nor U7793 (N_7793,N_6080,N_6096);
and U7794 (N_7794,N_6804,N_6565);
nor U7795 (N_7795,N_6255,N_6561);
nand U7796 (N_7796,N_6788,N_6442);
nand U7797 (N_7797,N_6122,N_6842);
or U7798 (N_7798,N_6293,N_6874);
or U7799 (N_7799,N_6381,N_6808);
xor U7800 (N_7800,N_6971,N_6476);
nor U7801 (N_7801,N_6682,N_6250);
xor U7802 (N_7802,N_6753,N_6252);
and U7803 (N_7803,N_6217,N_6190);
nor U7804 (N_7804,N_6962,N_6729);
nand U7805 (N_7805,N_6705,N_6484);
nand U7806 (N_7806,N_6103,N_6594);
nand U7807 (N_7807,N_6138,N_6988);
and U7808 (N_7808,N_6983,N_6487);
or U7809 (N_7809,N_6569,N_6908);
or U7810 (N_7810,N_6992,N_6254);
or U7811 (N_7811,N_6919,N_6509);
nand U7812 (N_7812,N_6899,N_6270);
or U7813 (N_7813,N_6487,N_6890);
nor U7814 (N_7814,N_6919,N_6362);
nor U7815 (N_7815,N_6233,N_6908);
and U7816 (N_7816,N_6448,N_6522);
or U7817 (N_7817,N_6907,N_6712);
or U7818 (N_7818,N_6080,N_6612);
and U7819 (N_7819,N_6917,N_6207);
or U7820 (N_7820,N_6952,N_6943);
nor U7821 (N_7821,N_6860,N_6619);
nor U7822 (N_7822,N_6240,N_6857);
xnor U7823 (N_7823,N_6889,N_6607);
nand U7824 (N_7824,N_6924,N_6994);
and U7825 (N_7825,N_6437,N_6813);
nand U7826 (N_7826,N_6497,N_6437);
or U7827 (N_7827,N_6716,N_6818);
or U7828 (N_7828,N_6413,N_6745);
and U7829 (N_7829,N_6549,N_6542);
nand U7830 (N_7830,N_6363,N_6737);
xor U7831 (N_7831,N_6476,N_6216);
and U7832 (N_7832,N_6828,N_6507);
xor U7833 (N_7833,N_6694,N_6984);
xnor U7834 (N_7834,N_6682,N_6781);
xor U7835 (N_7835,N_6672,N_6484);
and U7836 (N_7836,N_6559,N_6649);
or U7837 (N_7837,N_6484,N_6862);
and U7838 (N_7838,N_6815,N_6430);
and U7839 (N_7839,N_6021,N_6111);
nand U7840 (N_7840,N_6739,N_6281);
or U7841 (N_7841,N_6635,N_6056);
or U7842 (N_7842,N_6280,N_6841);
and U7843 (N_7843,N_6132,N_6339);
nand U7844 (N_7844,N_6418,N_6217);
nor U7845 (N_7845,N_6166,N_6047);
nand U7846 (N_7846,N_6231,N_6571);
or U7847 (N_7847,N_6595,N_6768);
or U7848 (N_7848,N_6619,N_6340);
nor U7849 (N_7849,N_6161,N_6690);
and U7850 (N_7850,N_6006,N_6207);
nor U7851 (N_7851,N_6880,N_6142);
or U7852 (N_7852,N_6692,N_6087);
or U7853 (N_7853,N_6586,N_6998);
nand U7854 (N_7854,N_6073,N_6315);
and U7855 (N_7855,N_6879,N_6250);
nand U7856 (N_7856,N_6457,N_6741);
nand U7857 (N_7857,N_6099,N_6408);
and U7858 (N_7858,N_6250,N_6195);
nor U7859 (N_7859,N_6683,N_6025);
nor U7860 (N_7860,N_6236,N_6754);
and U7861 (N_7861,N_6559,N_6396);
or U7862 (N_7862,N_6030,N_6221);
and U7863 (N_7863,N_6920,N_6010);
nor U7864 (N_7864,N_6060,N_6543);
and U7865 (N_7865,N_6195,N_6806);
and U7866 (N_7866,N_6707,N_6694);
nand U7867 (N_7867,N_6681,N_6313);
xnor U7868 (N_7868,N_6012,N_6393);
or U7869 (N_7869,N_6833,N_6215);
and U7870 (N_7870,N_6419,N_6376);
and U7871 (N_7871,N_6782,N_6841);
xor U7872 (N_7872,N_6082,N_6180);
xnor U7873 (N_7873,N_6122,N_6839);
xnor U7874 (N_7874,N_6287,N_6482);
nand U7875 (N_7875,N_6582,N_6091);
xnor U7876 (N_7876,N_6200,N_6208);
xnor U7877 (N_7877,N_6634,N_6813);
nand U7878 (N_7878,N_6081,N_6537);
and U7879 (N_7879,N_6419,N_6884);
nand U7880 (N_7880,N_6418,N_6716);
and U7881 (N_7881,N_6682,N_6403);
or U7882 (N_7882,N_6941,N_6570);
and U7883 (N_7883,N_6111,N_6699);
nand U7884 (N_7884,N_6470,N_6906);
xor U7885 (N_7885,N_6216,N_6957);
nor U7886 (N_7886,N_6011,N_6826);
and U7887 (N_7887,N_6300,N_6277);
nor U7888 (N_7888,N_6690,N_6700);
or U7889 (N_7889,N_6514,N_6983);
nand U7890 (N_7890,N_6598,N_6287);
and U7891 (N_7891,N_6788,N_6557);
nor U7892 (N_7892,N_6316,N_6830);
and U7893 (N_7893,N_6436,N_6523);
and U7894 (N_7894,N_6813,N_6929);
and U7895 (N_7895,N_6782,N_6364);
or U7896 (N_7896,N_6500,N_6055);
nand U7897 (N_7897,N_6036,N_6468);
and U7898 (N_7898,N_6937,N_6442);
nand U7899 (N_7899,N_6968,N_6851);
nand U7900 (N_7900,N_6000,N_6246);
or U7901 (N_7901,N_6460,N_6757);
nand U7902 (N_7902,N_6417,N_6564);
or U7903 (N_7903,N_6508,N_6979);
and U7904 (N_7904,N_6154,N_6634);
or U7905 (N_7905,N_6016,N_6638);
nand U7906 (N_7906,N_6828,N_6404);
nand U7907 (N_7907,N_6933,N_6664);
nand U7908 (N_7908,N_6035,N_6835);
or U7909 (N_7909,N_6112,N_6611);
nor U7910 (N_7910,N_6175,N_6513);
nand U7911 (N_7911,N_6759,N_6520);
nor U7912 (N_7912,N_6234,N_6354);
and U7913 (N_7913,N_6423,N_6242);
or U7914 (N_7914,N_6599,N_6999);
nor U7915 (N_7915,N_6398,N_6922);
nand U7916 (N_7916,N_6676,N_6985);
or U7917 (N_7917,N_6580,N_6922);
nor U7918 (N_7918,N_6213,N_6246);
nor U7919 (N_7919,N_6256,N_6561);
xor U7920 (N_7920,N_6526,N_6802);
or U7921 (N_7921,N_6593,N_6034);
nor U7922 (N_7922,N_6205,N_6130);
nor U7923 (N_7923,N_6441,N_6932);
or U7924 (N_7924,N_6187,N_6970);
nor U7925 (N_7925,N_6469,N_6357);
nand U7926 (N_7926,N_6156,N_6998);
nor U7927 (N_7927,N_6905,N_6057);
and U7928 (N_7928,N_6364,N_6132);
nor U7929 (N_7929,N_6093,N_6422);
nor U7930 (N_7930,N_6273,N_6895);
and U7931 (N_7931,N_6611,N_6851);
xnor U7932 (N_7932,N_6633,N_6770);
nand U7933 (N_7933,N_6722,N_6382);
nor U7934 (N_7934,N_6100,N_6494);
or U7935 (N_7935,N_6818,N_6608);
or U7936 (N_7936,N_6059,N_6580);
nor U7937 (N_7937,N_6018,N_6233);
nand U7938 (N_7938,N_6686,N_6499);
and U7939 (N_7939,N_6063,N_6198);
or U7940 (N_7940,N_6615,N_6362);
nand U7941 (N_7941,N_6120,N_6921);
nor U7942 (N_7942,N_6493,N_6644);
or U7943 (N_7943,N_6904,N_6742);
nand U7944 (N_7944,N_6145,N_6398);
or U7945 (N_7945,N_6755,N_6971);
nand U7946 (N_7946,N_6922,N_6524);
nor U7947 (N_7947,N_6437,N_6163);
nand U7948 (N_7948,N_6162,N_6329);
or U7949 (N_7949,N_6225,N_6148);
nand U7950 (N_7950,N_6554,N_6114);
nand U7951 (N_7951,N_6501,N_6534);
or U7952 (N_7952,N_6201,N_6059);
nand U7953 (N_7953,N_6974,N_6011);
nand U7954 (N_7954,N_6772,N_6358);
or U7955 (N_7955,N_6399,N_6654);
or U7956 (N_7956,N_6710,N_6682);
and U7957 (N_7957,N_6760,N_6413);
nor U7958 (N_7958,N_6867,N_6879);
nand U7959 (N_7959,N_6917,N_6458);
and U7960 (N_7960,N_6019,N_6102);
xor U7961 (N_7961,N_6661,N_6333);
or U7962 (N_7962,N_6367,N_6562);
nor U7963 (N_7963,N_6362,N_6009);
xor U7964 (N_7964,N_6528,N_6463);
and U7965 (N_7965,N_6986,N_6567);
and U7966 (N_7966,N_6762,N_6459);
and U7967 (N_7967,N_6274,N_6593);
xor U7968 (N_7968,N_6876,N_6296);
nor U7969 (N_7969,N_6047,N_6907);
nor U7970 (N_7970,N_6088,N_6542);
nor U7971 (N_7971,N_6731,N_6876);
xnor U7972 (N_7972,N_6945,N_6713);
nand U7973 (N_7973,N_6179,N_6779);
nand U7974 (N_7974,N_6814,N_6756);
xor U7975 (N_7975,N_6321,N_6246);
and U7976 (N_7976,N_6553,N_6341);
nand U7977 (N_7977,N_6506,N_6775);
or U7978 (N_7978,N_6648,N_6511);
or U7979 (N_7979,N_6507,N_6935);
and U7980 (N_7980,N_6805,N_6721);
nand U7981 (N_7981,N_6072,N_6436);
or U7982 (N_7982,N_6715,N_6319);
nor U7983 (N_7983,N_6134,N_6118);
nand U7984 (N_7984,N_6641,N_6779);
xor U7985 (N_7985,N_6759,N_6641);
nor U7986 (N_7986,N_6568,N_6790);
nor U7987 (N_7987,N_6633,N_6140);
xor U7988 (N_7988,N_6115,N_6449);
nor U7989 (N_7989,N_6370,N_6392);
and U7990 (N_7990,N_6207,N_6515);
nand U7991 (N_7991,N_6301,N_6069);
nand U7992 (N_7992,N_6236,N_6628);
or U7993 (N_7993,N_6044,N_6683);
or U7994 (N_7994,N_6822,N_6166);
and U7995 (N_7995,N_6750,N_6969);
or U7996 (N_7996,N_6949,N_6730);
nand U7997 (N_7997,N_6419,N_6805);
and U7998 (N_7998,N_6907,N_6461);
and U7999 (N_7999,N_6362,N_6608);
nand U8000 (N_8000,N_7292,N_7776);
xor U8001 (N_8001,N_7702,N_7359);
nand U8002 (N_8002,N_7074,N_7884);
nor U8003 (N_8003,N_7482,N_7503);
nand U8004 (N_8004,N_7034,N_7705);
and U8005 (N_8005,N_7000,N_7262);
and U8006 (N_8006,N_7852,N_7797);
and U8007 (N_8007,N_7231,N_7528);
nand U8008 (N_8008,N_7479,N_7440);
xor U8009 (N_8009,N_7144,N_7352);
xor U8010 (N_8010,N_7011,N_7239);
or U8011 (N_8011,N_7577,N_7882);
or U8012 (N_8012,N_7600,N_7115);
or U8013 (N_8013,N_7471,N_7271);
nand U8014 (N_8014,N_7757,N_7167);
nand U8015 (N_8015,N_7960,N_7159);
xor U8016 (N_8016,N_7826,N_7434);
nor U8017 (N_8017,N_7521,N_7507);
and U8018 (N_8018,N_7344,N_7936);
nand U8019 (N_8019,N_7018,N_7649);
nor U8020 (N_8020,N_7664,N_7931);
or U8021 (N_8021,N_7060,N_7963);
nand U8022 (N_8022,N_7904,N_7927);
or U8023 (N_8023,N_7297,N_7921);
nor U8024 (N_8024,N_7850,N_7300);
nor U8025 (N_8025,N_7427,N_7323);
nor U8026 (N_8026,N_7838,N_7501);
or U8027 (N_8027,N_7602,N_7943);
nor U8028 (N_8028,N_7338,N_7858);
and U8029 (N_8029,N_7619,N_7723);
and U8030 (N_8030,N_7730,N_7513);
nand U8031 (N_8031,N_7089,N_7994);
and U8032 (N_8032,N_7312,N_7306);
nand U8033 (N_8033,N_7182,N_7985);
or U8034 (N_8034,N_7714,N_7974);
nor U8035 (N_8035,N_7456,N_7106);
nand U8036 (N_8036,N_7532,N_7301);
nand U8037 (N_8037,N_7470,N_7047);
nand U8038 (N_8038,N_7367,N_7886);
nor U8039 (N_8039,N_7817,N_7995);
nor U8040 (N_8040,N_7895,N_7509);
or U8041 (N_8041,N_7918,N_7423);
nand U8042 (N_8042,N_7768,N_7123);
nand U8043 (N_8043,N_7962,N_7879);
nor U8044 (N_8044,N_7372,N_7582);
nand U8045 (N_8045,N_7021,N_7608);
nor U8046 (N_8046,N_7800,N_7540);
nor U8047 (N_8047,N_7706,N_7568);
and U8048 (N_8048,N_7908,N_7203);
nand U8049 (N_8049,N_7829,N_7105);
nand U8050 (N_8050,N_7117,N_7319);
nand U8051 (N_8051,N_7972,N_7808);
xnor U8052 (N_8052,N_7958,N_7631);
and U8053 (N_8053,N_7764,N_7846);
nand U8054 (N_8054,N_7790,N_7217);
and U8055 (N_8055,N_7779,N_7729);
nand U8056 (N_8056,N_7016,N_7265);
nand U8057 (N_8057,N_7576,N_7287);
nor U8058 (N_8058,N_7565,N_7221);
or U8059 (N_8059,N_7940,N_7032);
xor U8060 (N_8060,N_7594,N_7013);
and U8061 (N_8061,N_7303,N_7529);
or U8062 (N_8062,N_7067,N_7299);
xor U8063 (N_8063,N_7255,N_7014);
nor U8064 (N_8064,N_7928,N_7455);
or U8065 (N_8065,N_7320,N_7165);
and U8066 (N_8066,N_7481,N_7561);
or U8067 (N_8067,N_7238,N_7378);
nor U8068 (N_8068,N_7758,N_7857);
and U8069 (N_8069,N_7677,N_7487);
xnor U8070 (N_8070,N_7151,N_7726);
or U8071 (N_8071,N_7537,N_7530);
and U8072 (N_8072,N_7912,N_7294);
nor U8073 (N_8073,N_7461,N_7309);
or U8074 (N_8074,N_7674,N_7392);
or U8075 (N_8075,N_7272,N_7240);
and U8076 (N_8076,N_7101,N_7635);
or U8077 (N_8077,N_7458,N_7187);
or U8078 (N_8078,N_7062,N_7036);
nor U8079 (N_8079,N_7080,N_7172);
nor U8080 (N_8080,N_7515,N_7676);
and U8081 (N_8081,N_7870,N_7098);
nor U8082 (N_8082,N_7110,N_7787);
nor U8083 (N_8083,N_7666,N_7976);
nand U8084 (N_8084,N_7571,N_7542);
and U8085 (N_8085,N_7308,N_7526);
and U8086 (N_8086,N_7356,N_7129);
nand U8087 (N_8087,N_7999,N_7404);
or U8088 (N_8088,N_7346,N_7621);
xor U8089 (N_8089,N_7096,N_7745);
nand U8090 (N_8090,N_7951,N_7235);
nand U8091 (N_8091,N_7739,N_7026);
or U8092 (N_8092,N_7553,N_7006);
xnor U8093 (N_8093,N_7794,N_7788);
nor U8094 (N_8094,N_7875,N_7523);
nor U8095 (N_8095,N_7775,N_7317);
xor U8096 (N_8096,N_7865,N_7054);
nor U8097 (N_8097,N_7811,N_7896);
nor U8098 (N_8098,N_7448,N_7331);
or U8099 (N_8099,N_7048,N_7387);
nor U8100 (N_8100,N_7514,N_7212);
nor U8101 (N_8101,N_7930,N_7363);
and U8102 (N_8102,N_7848,N_7733);
and U8103 (N_8103,N_7942,N_7605);
xnor U8104 (N_8104,N_7206,N_7176);
and U8105 (N_8105,N_7349,N_7708);
or U8106 (N_8106,N_7008,N_7409);
and U8107 (N_8107,N_7329,N_7090);
or U8108 (N_8108,N_7925,N_7778);
nor U8109 (N_8109,N_7433,N_7044);
and U8110 (N_8110,N_7830,N_7717);
nor U8111 (N_8111,N_7780,N_7200);
or U8112 (N_8112,N_7593,N_7385);
nand U8113 (N_8113,N_7386,N_7075);
xor U8114 (N_8114,N_7570,N_7230);
nand U8115 (N_8115,N_7506,N_7658);
nand U8116 (N_8116,N_7397,N_7411);
or U8117 (N_8117,N_7375,N_7854);
xnor U8118 (N_8118,N_7480,N_7701);
nand U8119 (N_8119,N_7412,N_7224);
and U8120 (N_8120,N_7132,N_7087);
nand U8121 (N_8121,N_7724,N_7641);
nor U8122 (N_8122,N_7076,N_7831);
nand U8123 (N_8123,N_7073,N_7045);
or U8124 (N_8124,N_7406,N_7964);
or U8125 (N_8125,N_7396,N_7244);
nand U8126 (N_8126,N_7274,N_7228);
and U8127 (N_8127,N_7683,N_7276);
nor U8128 (N_8128,N_7148,N_7660);
or U8129 (N_8129,N_7825,N_7314);
and U8130 (N_8130,N_7969,N_7316);
nand U8131 (N_8131,N_7939,N_7141);
nor U8132 (N_8132,N_7107,N_7335);
nor U8133 (N_8133,N_7010,N_7465);
xor U8134 (N_8134,N_7145,N_7755);
nand U8135 (N_8135,N_7158,N_7219);
nor U8136 (N_8136,N_7613,N_7188);
and U8137 (N_8137,N_7178,N_7252);
or U8138 (N_8138,N_7659,N_7259);
nor U8139 (N_8139,N_7476,N_7686);
and U8140 (N_8140,N_7586,N_7562);
nor U8141 (N_8141,N_7247,N_7849);
nand U8142 (N_8142,N_7160,N_7707);
nand U8143 (N_8143,N_7863,N_7260);
and U8144 (N_8144,N_7256,N_7782);
and U8145 (N_8145,N_7688,N_7722);
nand U8146 (N_8146,N_7190,N_7606);
nor U8147 (N_8147,N_7245,N_7795);
or U8148 (N_8148,N_7332,N_7401);
or U8149 (N_8149,N_7901,N_7307);
and U8150 (N_8150,N_7747,N_7508);
xor U8151 (N_8151,N_7078,N_7358);
and U8152 (N_8152,N_7803,N_7590);
and U8153 (N_8153,N_7667,N_7700);
nand U8154 (N_8154,N_7202,N_7418);
or U8155 (N_8155,N_7833,N_7281);
xnor U8156 (N_8156,N_7862,N_7064);
nand U8157 (N_8157,N_7622,N_7947);
and U8158 (N_8158,N_7012,N_7545);
nand U8159 (N_8159,N_7236,N_7491);
nor U8160 (N_8160,N_7607,N_7398);
or U8161 (N_8161,N_7986,N_7524);
and U8162 (N_8162,N_7431,N_7368);
nor U8163 (N_8163,N_7258,N_7834);
or U8164 (N_8164,N_7836,N_7612);
and U8165 (N_8165,N_7337,N_7474);
nor U8166 (N_8166,N_7632,N_7469);
or U8167 (N_8167,N_7112,N_7761);
or U8168 (N_8168,N_7381,N_7327);
xnor U8169 (N_8169,N_7061,N_7818);
nand U8170 (N_8170,N_7801,N_7156);
or U8171 (N_8171,N_7166,N_7467);
nor U8172 (N_8172,N_7170,N_7139);
nand U8173 (N_8173,N_7365,N_7626);
and U8174 (N_8174,N_7192,N_7719);
and U8175 (N_8175,N_7634,N_7888);
nor U8176 (N_8176,N_7120,N_7116);
or U8177 (N_8177,N_7445,N_7580);
nand U8178 (N_8178,N_7710,N_7907);
nand U8179 (N_8179,N_7189,N_7791);
nand U8180 (N_8180,N_7598,N_7184);
and U8181 (N_8181,N_7589,N_7227);
and U8182 (N_8182,N_7222,N_7750);
or U8183 (N_8183,N_7655,N_7906);
xor U8184 (N_8184,N_7871,N_7620);
nor U8185 (N_8185,N_7454,N_7450);
and U8186 (N_8186,N_7922,N_7422);
and U8187 (N_8187,N_7806,N_7771);
nand U8188 (N_8188,N_7257,N_7390);
xor U8189 (N_8189,N_7715,N_7017);
nand U8190 (N_8190,N_7629,N_7304);
nor U8191 (N_8191,N_7822,N_7197);
or U8192 (N_8192,N_7040,N_7143);
and U8193 (N_8193,N_7547,N_7122);
nor U8194 (N_8194,N_7393,N_7127);
or U8195 (N_8195,N_7534,N_7627);
nand U8196 (N_8196,N_7805,N_7993);
or U8197 (N_8197,N_7214,N_7815);
and U8198 (N_8198,N_7373,N_7675);
nand U8199 (N_8199,N_7573,N_7201);
and U8200 (N_8200,N_7379,N_7874);
nand U8201 (N_8201,N_7002,N_7405);
or U8202 (N_8202,N_7867,N_7554);
nor U8203 (N_8203,N_7037,N_7732);
xnor U8204 (N_8204,N_7486,N_7114);
nand U8205 (N_8205,N_7001,N_7920);
xor U8206 (N_8206,N_7648,N_7211);
or U8207 (N_8207,N_7654,N_7519);
nor U8208 (N_8208,N_7687,N_7909);
nand U8209 (N_8209,N_7384,N_7760);
nand U8210 (N_8210,N_7694,N_7408);
or U8211 (N_8211,N_7934,N_7223);
or U8212 (N_8212,N_7269,N_7578);
nor U8213 (N_8213,N_7926,N_7389);
nand U8214 (N_8214,N_7816,N_7983);
nor U8215 (N_8215,N_7083,N_7793);
or U8216 (N_8216,N_7555,N_7483);
and U8217 (N_8217,N_7881,N_7682);
or U8218 (N_8218,N_7610,N_7426);
and U8219 (N_8219,N_7376,N_7885);
nor U8220 (N_8220,N_7277,N_7441);
nor U8221 (N_8221,N_7652,N_7585);
and U8222 (N_8222,N_7897,N_7414);
and U8223 (N_8223,N_7827,N_7351);
nand U8224 (N_8224,N_7341,N_7614);
and U8225 (N_8225,N_7168,N_7992);
nor U8226 (N_8226,N_7894,N_7961);
xor U8227 (N_8227,N_7699,N_7539);
nor U8228 (N_8228,N_7919,N_7334);
and U8229 (N_8229,N_7574,N_7394);
nand U8230 (N_8230,N_7743,N_7935);
and U8231 (N_8231,N_7740,N_7137);
or U8232 (N_8232,N_7058,N_7289);
nor U8233 (N_8233,N_7738,N_7859);
nand U8234 (N_8234,N_7004,N_7978);
and U8235 (N_8235,N_7847,N_7678);
nand U8236 (N_8236,N_7656,N_7302);
nand U8237 (N_8237,N_7280,N_7751);
and U8238 (N_8238,N_7877,N_7218);
xnor U8239 (N_8239,N_7956,N_7057);
or U8240 (N_8240,N_7009,N_7777);
nand U8241 (N_8241,N_7752,N_7169);
nand U8242 (N_8242,N_7024,N_7878);
nor U8243 (N_8243,N_7288,N_7633);
nor U8244 (N_8244,N_7042,N_7759);
nand U8245 (N_8245,N_7400,N_7371);
nand U8246 (N_8246,N_7975,N_7840);
nand U8247 (N_8247,N_7609,N_7429);
and U8248 (N_8248,N_7572,N_7510);
nor U8249 (N_8249,N_7873,N_7275);
nor U8250 (N_8250,N_7020,N_7611);
and U8251 (N_8251,N_7193,N_7679);
or U8252 (N_8252,N_7564,N_7603);
or U8253 (N_8253,N_7071,N_7027);
nor U8254 (N_8254,N_7196,N_7282);
nand U8255 (N_8255,N_7938,N_7949);
xor U8256 (N_8256,N_7597,N_7923);
and U8257 (N_8257,N_7615,N_7637);
nand U8258 (N_8258,N_7749,N_7842);
nand U8259 (N_8259,N_7003,N_7407);
nand U8260 (N_8260,N_7792,N_7097);
nand U8261 (N_8261,N_7070,N_7536);
and U8262 (N_8262,N_7866,N_7968);
nand U8263 (N_8263,N_7225,N_7543);
xor U8264 (N_8264,N_7796,N_7933);
nand U8265 (N_8265,N_7579,N_7742);
or U8266 (N_8266,N_7703,N_7518);
xnor U8267 (N_8267,N_7913,N_7581);
and U8268 (N_8268,N_7232,N_7033);
or U8269 (N_8269,N_7860,N_7059);
and U8270 (N_8270,N_7204,N_7250);
nand U8271 (N_8271,N_7497,N_7081);
or U8272 (N_8272,N_7601,N_7929);
and U8273 (N_8273,N_7814,N_7183);
nor U8274 (N_8274,N_7134,N_7869);
nand U8275 (N_8275,N_7522,N_7068);
xor U8276 (N_8276,N_7763,N_7459);
nor U8277 (N_8277,N_7551,N_7171);
xor U8278 (N_8278,N_7639,N_7485);
nor U8279 (N_8279,N_7488,N_7439);
nand U8280 (N_8280,N_7587,N_7413);
or U8281 (N_8281,N_7864,N_7462);
and U8282 (N_8282,N_7417,N_7944);
or U8283 (N_8283,N_7124,N_7069);
xor U8284 (N_8284,N_7911,N_7902);
nor U8285 (N_8285,N_7556,N_7741);
xnor U8286 (N_8286,N_7432,N_7802);
nand U8287 (N_8287,N_7030,N_7665);
nor U8288 (N_8288,N_7727,N_7436);
and U8289 (N_8289,N_7451,N_7950);
and U8290 (N_8290,N_7765,N_7689);
xor U8291 (N_8291,N_7584,N_7125);
nor U8292 (N_8292,N_7038,N_7162);
or U8293 (N_8293,N_7711,N_7546);
nand U8294 (N_8294,N_7208,N_7981);
and U8295 (N_8295,N_7511,N_7493);
xor U8296 (N_8296,N_7267,N_7893);
nand U8297 (N_8297,N_7948,N_7136);
or U8298 (N_8298,N_7813,N_7286);
nand U8299 (N_8299,N_7043,N_7149);
xnor U8300 (N_8300,N_7924,N_7642);
and U8301 (N_8301,N_7229,N_7498);
nand U8302 (N_8302,N_7118,N_7015);
and U8303 (N_8303,N_7173,N_7628);
nor U8304 (N_8304,N_7754,N_7851);
and U8305 (N_8305,N_7022,N_7100);
and U8306 (N_8306,N_7746,N_7653);
nand U8307 (N_8307,N_7916,N_7736);
or U8308 (N_8308,N_7366,N_7261);
xor U8309 (N_8309,N_7266,N_7824);
and U8310 (N_8310,N_7370,N_7504);
nand U8311 (N_8311,N_7861,N_7194);
and U8312 (N_8312,N_7377,N_7531);
nor U8313 (N_8313,N_7186,N_7636);
and U8314 (N_8314,N_7273,N_7987);
and U8315 (N_8315,N_7041,N_7290);
nor U8316 (N_8316,N_7399,N_7086);
or U8317 (N_8317,N_7326,N_7065);
and U8318 (N_8318,N_7638,N_7991);
nor U8319 (N_8319,N_7887,N_7880);
nor U8320 (N_8320,N_7889,N_7050);
nand U8321 (N_8321,N_7430,N_7246);
and U8322 (N_8322,N_7311,N_7077);
xor U8323 (N_8323,N_7416,N_7525);
nor U8324 (N_8324,N_7696,N_7322);
or U8325 (N_8325,N_7293,N_7369);
or U8326 (N_8326,N_7647,N_7671);
or U8327 (N_8327,N_7296,N_7820);
nor U8328 (N_8328,N_7391,N_7910);
nand U8329 (N_8329,N_7102,N_7126);
and U8330 (N_8330,N_7342,N_7198);
or U8331 (N_8331,N_7029,N_7180);
nor U8332 (N_8332,N_7163,N_7079);
or U8333 (N_8333,N_7548,N_7268);
nand U8334 (N_8334,N_7575,N_7155);
nand U8335 (N_8335,N_7899,N_7891);
nor U8336 (N_8336,N_7415,N_7446);
nor U8337 (N_8337,N_7199,N_7005);
and U8338 (N_8338,N_7807,N_7028);
or U8339 (N_8339,N_7959,N_7072);
xnor U8340 (N_8340,N_7599,N_7990);
and U8341 (N_8341,N_7977,N_7205);
or U8342 (N_8342,N_7443,N_7588);
or U8343 (N_8343,N_7955,N_7447);
or U8344 (N_8344,N_7063,N_7680);
nand U8345 (N_8345,N_7350,N_7616);
or U8346 (N_8346,N_7130,N_7147);
xnor U8347 (N_8347,N_7592,N_7552);
and U8348 (N_8348,N_7997,N_7785);
xor U8349 (N_8349,N_7684,N_7364);
xnor U8350 (N_8350,N_7868,N_7496);
nor U8351 (N_8351,N_7789,N_7357);
or U8352 (N_8352,N_7318,N_7313);
nor U8353 (N_8353,N_7783,N_7645);
nand U8354 (N_8354,N_7099,N_7725);
and U8355 (N_8355,N_7890,N_7971);
nand U8356 (N_8356,N_7770,N_7133);
and U8357 (N_8357,N_7544,N_7640);
nand U8358 (N_8358,N_7569,N_7291);
nand U8359 (N_8359,N_7898,N_7388);
or U8360 (N_8360,N_7786,N_7031);
and U8361 (N_8361,N_7767,N_7953);
and U8362 (N_8362,N_7263,N_7839);
or U8363 (N_8363,N_7812,N_7973);
nor U8364 (N_8364,N_7856,N_7354);
nand U8365 (N_8365,N_7735,N_7663);
and U8366 (N_8366,N_7175,N_7049);
xnor U8367 (N_8367,N_7685,N_7954);
nor U8368 (N_8368,N_7023,N_7734);
or U8369 (N_8369,N_7595,N_7035);
and U8370 (N_8370,N_7932,N_7821);
nor U8371 (N_8371,N_7138,N_7131);
and U8372 (N_8372,N_7512,N_7728);
and U8373 (N_8373,N_7494,N_7055);
nand U8374 (N_8374,N_7567,N_7108);
or U8375 (N_8375,N_7965,N_7563);
and U8376 (N_8376,N_7774,N_7091);
and U8377 (N_8377,N_7468,N_7650);
nor U8378 (N_8378,N_7784,N_7744);
nor U8379 (N_8379,N_7185,N_7917);
nor U8380 (N_8380,N_7718,N_7892);
and U8381 (N_8381,N_7695,N_7984);
nor U8382 (N_8382,N_7154,N_7477);
and U8383 (N_8383,N_7088,N_7243);
xnor U8384 (N_8384,N_7835,N_7690);
nor U8385 (N_8385,N_7713,N_7618);
and U8386 (N_8386,N_7502,N_7533);
or U8387 (N_8387,N_7437,N_7419);
nor U8388 (N_8388,N_7980,N_7111);
or U8389 (N_8389,N_7772,N_7104);
nor U8390 (N_8390,N_7355,N_7855);
or U8391 (N_8391,N_7668,N_7095);
and U8392 (N_8392,N_7270,N_7520);
or U8393 (N_8393,N_7428,N_7464);
xnor U8394 (N_8394,N_7492,N_7453);
nor U8395 (N_8395,N_7082,N_7698);
nand U8396 (N_8396,N_7844,N_7558);
and U8397 (N_8397,N_7146,N_7490);
or U8398 (N_8398,N_7946,N_7457);
or U8399 (N_8399,N_7460,N_7425);
nand U8400 (N_8400,N_7500,N_7720);
or U8401 (N_8401,N_7541,N_7538);
nor U8402 (N_8402,N_7403,N_7254);
or U8403 (N_8403,N_7053,N_7140);
nor U8404 (N_8404,N_7798,N_7809);
and U8405 (N_8405,N_7495,N_7085);
or U8406 (N_8406,N_7121,N_7216);
and U8407 (N_8407,N_7237,N_7672);
and U8408 (N_8408,N_7253,N_7161);
nand U8409 (N_8409,N_7915,N_7191);
nand U8410 (N_8410,N_7596,N_7452);
and U8411 (N_8411,N_7823,N_7819);
nor U8412 (N_8412,N_7348,N_7279);
or U8413 (N_8413,N_7285,N_7712);
nand U8414 (N_8414,N_7340,N_7941);
or U8415 (N_8415,N_7142,N_7937);
nor U8416 (N_8416,N_7952,N_7410);
and U8417 (N_8417,N_7421,N_7527);
or U8418 (N_8418,N_7233,N_7242);
or U8419 (N_8419,N_7853,N_7505);
xor U8420 (N_8420,N_7762,N_7651);
and U8421 (N_8421,N_7152,N_7177);
nor U8422 (N_8422,N_7310,N_7164);
nor U8423 (N_8423,N_7150,N_7623);
and U8424 (N_8424,N_7181,N_7845);
nor U8425 (N_8425,N_7153,N_7905);
xnor U8426 (N_8426,N_7025,N_7900);
and U8427 (N_8427,N_7345,N_7591);
nand U8428 (N_8428,N_7709,N_7324);
nand U8429 (N_8429,N_7996,N_7692);
or U8430 (N_8430,N_7438,N_7084);
nand U8431 (N_8431,N_7773,N_7325);
or U8432 (N_8432,N_7550,N_7007);
nor U8433 (N_8433,N_7264,N_7721);
or U8434 (N_8434,N_7673,N_7566);
nor U8435 (N_8435,N_7046,N_7693);
and U8436 (N_8436,N_7876,N_7226);
nor U8437 (N_8437,N_7420,N_7174);
nand U8438 (N_8438,N_7625,N_7799);
or U8439 (N_8439,N_7113,N_7957);
and U8440 (N_8440,N_7251,N_7557);
nand U8441 (N_8441,N_7516,N_7535);
nand U8442 (N_8442,N_7435,N_7872);
nor U8443 (N_8443,N_7119,N_7383);
and U8444 (N_8444,N_7837,N_7967);
xnor U8445 (N_8445,N_7103,N_7361);
nor U8446 (N_8446,N_7249,N_7475);
nor U8447 (N_8447,N_7328,N_7157);
nor U8448 (N_8448,N_7298,N_7662);
nand U8449 (N_8449,N_7748,N_7998);
or U8450 (N_8450,N_7449,N_7979);
nand U8451 (N_8451,N_7914,N_7731);
xnor U8452 (N_8452,N_7374,N_7330);
or U8453 (N_8453,N_7278,N_7644);
and U8454 (N_8454,N_7560,N_7333);
nor U8455 (N_8455,N_7362,N_7691);
xor U8456 (N_8456,N_7248,N_7210);
nor U8457 (N_8457,N_7988,N_7305);
nor U8458 (N_8458,N_7716,N_7234);
or U8459 (N_8459,N_7945,N_7472);
nand U8460 (N_8460,N_7617,N_7756);
and U8461 (N_8461,N_7810,N_7402);
nor U8462 (N_8462,N_7466,N_7339);
nor U8463 (N_8463,N_7473,N_7336);
or U8464 (N_8464,N_7681,N_7195);
or U8465 (N_8465,N_7583,N_7463);
and U8466 (N_8466,N_7737,N_7128);
and U8467 (N_8467,N_7360,N_7109);
or U8468 (N_8468,N_7670,N_7484);
nand U8469 (N_8469,N_7135,N_7559);
nor U8470 (N_8470,N_7321,N_7051);
nor U8471 (N_8471,N_7843,N_7630);
xnor U8472 (N_8472,N_7209,N_7424);
or U8473 (N_8473,N_7284,N_7444);
nor U8474 (N_8474,N_7382,N_7832);
and U8475 (N_8475,N_7295,N_7704);
or U8476 (N_8476,N_7643,N_7669);
xnor U8477 (N_8477,N_7395,N_7970);
and U8478 (N_8478,N_7781,N_7661);
nor U8479 (N_8479,N_7093,N_7315);
or U8480 (N_8480,N_7220,N_7207);
and U8481 (N_8481,N_7753,N_7841);
nand U8482 (N_8482,N_7213,N_7066);
nand U8483 (N_8483,N_7380,N_7353);
or U8484 (N_8484,N_7347,N_7517);
xnor U8485 (N_8485,N_7489,N_7241);
xor U8486 (N_8486,N_7094,N_7766);
and U8487 (N_8487,N_7804,N_7442);
nor U8488 (N_8488,N_7903,N_7039);
and U8489 (N_8489,N_7052,N_7982);
or U8490 (N_8490,N_7283,N_7657);
and U8491 (N_8491,N_7769,N_7478);
nor U8492 (N_8492,N_7499,N_7092);
and U8493 (N_8493,N_7828,N_7056);
and U8494 (N_8494,N_7989,N_7966);
nor U8495 (N_8495,N_7883,N_7697);
or U8496 (N_8496,N_7019,N_7215);
nor U8497 (N_8497,N_7624,N_7646);
xnor U8498 (N_8498,N_7179,N_7604);
nand U8499 (N_8499,N_7343,N_7549);
and U8500 (N_8500,N_7613,N_7817);
or U8501 (N_8501,N_7821,N_7352);
nand U8502 (N_8502,N_7308,N_7486);
xor U8503 (N_8503,N_7224,N_7676);
and U8504 (N_8504,N_7570,N_7847);
nor U8505 (N_8505,N_7388,N_7121);
and U8506 (N_8506,N_7905,N_7296);
nor U8507 (N_8507,N_7898,N_7972);
nor U8508 (N_8508,N_7177,N_7107);
and U8509 (N_8509,N_7708,N_7151);
and U8510 (N_8510,N_7162,N_7614);
or U8511 (N_8511,N_7023,N_7300);
nand U8512 (N_8512,N_7531,N_7448);
nor U8513 (N_8513,N_7092,N_7896);
nor U8514 (N_8514,N_7180,N_7887);
or U8515 (N_8515,N_7311,N_7577);
xor U8516 (N_8516,N_7957,N_7480);
and U8517 (N_8517,N_7571,N_7648);
or U8518 (N_8518,N_7721,N_7715);
nand U8519 (N_8519,N_7286,N_7801);
xnor U8520 (N_8520,N_7167,N_7256);
xor U8521 (N_8521,N_7498,N_7515);
and U8522 (N_8522,N_7380,N_7175);
nor U8523 (N_8523,N_7105,N_7547);
nor U8524 (N_8524,N_7849,N_7288);
and U8525 (N_8525,N_7162,N_7505);
nand U8526 (N_8526,N_7012,N_7801);
nor U8527 (N_8527,N_7037,N_7970);
nor U8528 (N_8528,N_7422,N_7309);
nor U8529 (N_8529,N_7644,N_7305);
or U8530 (N_8530,N_7522,N_7313);
nand U8531 (N_8531,N_7081,N_7611);
and U8532 (N_8532,N_7584,N_7870);
or U8533 (N_8533,N_7716,N_7158);
nor U8534 (N_8534,N_7816,N_7161);
nand U8535 (N_8535,N_7887,N_7424);
nand U8536 (N_8536,N_7532,N_7920);
and U8537 (N_8537,N_7918,N_7460);
and U8538 (N_8538,N_7121,N_7832);
nand U8539 (N_8539,N_7476,N_7049);
nor U8540 (N_8540,N_7543,N_7189);
and U8541 (N_8541,N_7982,N_7189);
or U8542 (N_8542,N_7938,N_7575);
and U8543 (N_8543,N_7812,N_7179);
or U8544 (N_8544,N_7808,N_7119);
or U8545 (N_8545,N_7792,N_7495);
or U8546 (N_8546,N_7009,N_7573);
and U8547 (N_8547,N_7159,N_7393);
and U8548 (N_8548,N_7879,N_7409);
nor U8549 (N_8549,N_7388,N_7814);
or U8550 (N_8550,N_7263,N_7414);
and U8551 (N_8551,N_7309,N_7493);
nand U8552 (N_8552,N_7061,N_7398);
nand U8553 (N_8553,N_7717,N_7647);
and U8554 (N_8554,N_7272,N_7090);
nor U8555 (N_8555,N_7259,N_7755);
nor U8556 (N_8556,N_7861,N_7899);
nand U8557 (N_8557,N_7583,N_7600);
nor U8558 (N_8558,N_7575,N_7224);
or U8559 (N_8559,N_7846,N_7944);
nor U8560 (N_8560,N_7973,N_7878);
nand U8561 (N_8561,N_7295,N_7003);
and U8562 (N_8562,N_7019,N_7369);
xor U8563 (N_8563,N_7570,N_7211);
and U8564 (N_8564,N_7074,N_7857);
and U8565 (N_8565,N_7043,N_7097);
nand U8566 (N_8566,N_7985,N_7752);
or U8567 (N_8567,N_7815,N_7673);
nand U8568 (N_8568,N_7830,N_7361);
and U8569 (N_8569,N_7766,N_7258);
nor U8570 (N_8570,N_7791,N_7497);
or U8571 (N_8571,N_7875,N_7708);
nand U8572 (N_8572,N_7002,N_7178);
or U8573 (N_8573,N_7566,N_7715);
nor U8574 (N_8574,N_7581,N_7283);
and U8575 (N_8575,N_7930,N_7634);
or U8576 (N_8576,N_7398,N_7858);
and U8577 (N_8577,N_7626,N_7018);
and U8578 (N_8578,N_7988,N_7377);
or U8579 (N_8579,N_7907,N_7465);
nor U8580 (N_8580,N_7838,N_7403);
or U8581 (N_8581,N_7750,N_7335);
or U8582 (N_8582,N_7269,N_7516);
xnor U8583 (N_8583,N_7315,N_7007);
nand U8584 (N_8584,N_7048,N_7003);
nor U8585 (N_8585,N_7514,N_7762);
nand U8586 (N_8586,N_7617,N_7971);
or U8587 (N_8587,N_7881,N_7226);
xnor U8588 (N_8588,N_7444,N_7949);
and U8589 (N_8589,N_7553,N_7651);
or U8590 (N_8590,N_7974,N_7200);
nand U8591 (N_8591,N_7412,N_7005);
xor U8592 (N_8592,N_7759,N_7191);
nor U8593 (N_8593,N_7876,N_7452);
or U8594 (N_8594,N_7273,N_7319);
nand U8595 (N_8595,N_7333,N_7784);
or U8596 (N_8596,N_7951,N_7810);
nand U8597 (N_8597,N_7344,N_7956);
or U8598 (N_8598,N_7979,N_7652);
and U8599 (N_8599,N_7077,N_7432);
or U8600 (N_8600,N_7174,N_7871);
or U8601 (N_8601,N_7209,N_7860);
xnor U8602 (N_8602,N_7193,N_7446);
and U8603 (N_8603,N_7682,N_7784);
nand U8604 (N_8604,N_7504,N_7550);
nand U8605 (N_8605,N_7492,N_7350);
nand U8606 (N_8606,N_7909,N_7679);
and U8607 (N_8607,N_7391,N_7046);
and U8608 (N_8608,N_7938,N_7331);
nor U8609 (N_8609,N_7469,N_7378);
nand U8610 (N_8610,N_7809,N_7791);
nand U8611 (N_8611,N_7029,N_7428);
xor U8612 (N_8612,N_7874,N_7356);
nand U8613 (N_8613,N_7312,N_7935);
and U8614 (N_8614,N_7097,N_7563);
xnor U8615 (N_8615,N_7550,N_7636);
and U8616 (N_8616,N_7195,N_7718);
and U8617 (N_8617,N_7931,N_7760);
nand U8618 (N_8618,N_7998,N_7559);
nor U8619 (N_8619,N_7425,N_7738);
or U8620 (N_8620,N_7629,N_7365);
nor U8621 (N_8621,N_7287,N_7522);
nand U8622 (N_8622,N_7220,N_7737);
nand U8623 (N_8623,N_7545,N_7792);
xnor U8624 (N_8624,N_7359,N_7939);
xor U8625 (N_8625,N_7087,N_7623);
and U8626 (N_8626,N_7786,N_7907);
xnor U8627 (N_8627,N_7100,N_7224);
xnor U8628 (N_8628,N_7696,N_7553);
and U8629 (N_8629,N_7819,N_7746);
nand U8630 (N_8630,N_7371,N_7049);
nand U8631 (N_8631,N_7968,N_7723);
or U8632 (N_8632,N_7455,N_7842);
or U8633 (N_8633,N_7700,N_7351);
nor U8634 (N_8634,N_7162,N_7187);
nor U8635 (N_8635,N_7089,N_7216);
and U8636 (N_8636,N_7257,N_7481);
nor U8637 (N_8637,N_7700,N_7105);
or U8638 (N_8638,N_7481,N_7649);
xnor U8639 (N_8639,N_7808,N_7992);
nor U8640 (N_8640,N_7800,N_7185);
or U8641 (N_8641,N_7925,N_7727);
nand U8642 (N_8642,N_7487,N_7965);
nand U8643 (N_8643,N_7887,N_7655);
xnor U8644 (N_8644,N_7241,N_7041);
nand U8645 (N_8645,N_7266,N_7458);
nand U8646 (N_8646,N_7555,N_7640);
and U8647 (N_8647,N_7887,N_7176);
nand U8648 (N_8648,N_7448,N_7991);
or U8649 (N_8649,N_7124,N_7365);
nor U8650 (N_8650,N_7163,N_7220);
nand U8651 (N_8651,N_7687,N_7241);
nand U8652 (N_8652,N_7093,N_7455);
nand U8653 (N_8653,N_7227,N_7632);
xnor U8654 (N_8654,N_7226,N_7924);
or U8655 (N_8655,N_7866,N_7566);
nand U8656 (N_8656,N_7174,N_7897);
nand U8657 (N_8657,N_7979,N_7281);
and U8658 (N_8658,N_7038,N_7144);
and U8659 (N_8659,N_7484,N_7447);
nand U8660 (N_8660,N_7989,N_7447);
or U8661 (N_8661,N_7115,N_7009);
or U8662 (N_8662,N_7972,N_7351);
nor U8663 (N_8663,N_7852,N_7406);
and U8664 (N_8664,N_7406,N_7186);
xnor U8665 (N_8665,N_7011,N_7688);
and U8666 (N_8666,N_7243,N_7273);
and U8667 (N_8667,N_7397,N_7945);
xnor U8668 (N_8668,N_7345,N_7056);
or U8669 (N_8669,N_7899,N_7466);
nand U8670 (N_8670,N_7326,N_7355);
nor U8671 (N_8671,N_7500,N_7678);
or U8672 (N_8672,N_7091,N_7248);
and U8673 (N_8673,N_7778,N_7333);
nor U8674 (N_8674,N_7941,N_7918);
or U8675 (N_8675,N_7297,N_7337);
nor U8676 (N_8676,N_7998,N_7640);
nor U8677 (N_8677,N_7838,N_7600);
and U8678 (N_8678,N_7232,N_7570);
or U8679 (N_8679,N_7764,N_7823);
nor U8680 (N_8680,N_7119,N_7090);
and U8681 (N_8681,N_7221,N_7332);
or U8682 (N_8682,N_7539,N_7191);
nand U8683 (N_8683,N_7971,N_7934);
nor U8684 (N_8684,N_7248,N_7888);
nor U8685 (N_8685,N_7927,N_7466);
nand U8686 (N_8686,N_7265,N_7686);
or U8687 (N_8687,N_7307,N_7393);
nor U8688 (N_8688,N_7211,N_7010);
nor U8689 (N_8689,N_7970,N_7152);
or U8690 (N_8690,N_7195,N_7614);
and U8691 (N_8691,N_7938,N_7114);
and U8692 (N_8692,N_7643,N_7289);
and U8693 (N_8693,N_7738,N_7407);
nor U8694 (N_8694,N_7373,N_7501);
nor U8695 (N_8695,N_7039,N_7835);
nand U8696 (N_8696,N_7171,N_7319);
or U8697 (N_8697,N_7068,N_7489);
nand U8698 (N_8698,N_7480,N_7844);
nor U8699 (N_8699,N_7903,N_7100);
and U8700 (N_8700,N_7715,N_7813);
or U8701 (N_8701,N_7725,N_7381);
nor U8702 (N_8702,N_7856,N_7444);
or U8703 (N_8703,N_7817,N_7770);
xor U8704 (N_8704,N_7813,N_7928);
and U8705 (N_8705,N_7118,N_7735);
nor U8706 (N_8706,N_7958,N_7514);
nor U8707 (N_8707,N_7810,N_7342);
nand U8708 (N_8708,N_7126,N_7371);
or U8709 (N_8709,N_7767,N_7144);
nand U8710 (N_8710,N_7764,N_7700);
nand U8711 (N_8711,N_7211,N_7645);
nand U8712 (N_8712,N_7392,N_7668);
and U8713 (N_8713,N_7045,N_7429);
or U8714 (N_8714,N_7441,N_7166);
or U8715 (N_8715,N_7219,N_7967);
xor U8716 (N_8716,N_7648,N_7420);
nand U8717 (N_8717,N_7680,N_7272);
nor U8718 (N_8718,N_7546,N_7484);
nand U8719 (N_8719,N_7782,N_7613);
or U8720 (N_8720,N_7763,N_7104);
or U8721 (N_8721,N_7945,N_7663);
nor U8722 (N_8722,N_7101,N_7143);
and U8723 (N_8723,N_7668,N_7771);
nor U8724 (N_8724,N_7853,N_7072);
and U8725 (N_8725,N_7810,N_7333);
or U8726 (N_8726,N_7971,N_7798);
and U8727 (N_8727,N_7203,N_7769);
or U8728 (N_8728,N_7626,N_7056);
nor U8729 (N_8729,N_7631,N_7040);
or U8730 (N_8730,N_7141,N_7620);
and U8731 (N_8731,N_7469,N_7686);
xor U8732 (N_8732,N_7416,N_7917);
xnor U8733 (N_8733,N_7075,N_7976);
nor U8734 (N_8734,N_7531,N_7254);
and U8735 (N_8735,N_7722,N_7914);
or U8736 (N_8736,N_7352,N_7509);
and U8737 (N_8737,N_7506,N_7892);
nor U8738 (N_8738,N_7524,N_7551);
or U8739 (N_8739,N_7603,N_7477);
nor U8740 (N_8740,N_7090,N_7990);
or U8741 (N_8741,N_7698,N_7167);
or U8742 (N_8742,N_7099,N_7805);
nor U8743 (N_8743,N_7423,N_7855);
nand U8744 (N_8744,N_7201,N_7822);
nor U8745 (N_8745,N_7314,N_7529);
xor U8746 (N_8746,N_7513,N_7413);
nor U8747 (N_8747,N_7188,N_7139);
and U8748 (N_8748,N_7910,N_7342);
and U8749 (N_8749,N_7225,N_7798);
or U8750 (N_8750,N_7947,N_7844);
and U8751 (N_8751,N_7196,N_7936);
and U8752 (N_8752,N_7279,N_7329);
or U8753 (N_8753,N_7097,N_7113);
xor U8754 (N_8754,N_7865,N_7205);
xor U8755 (N_8755,N_7828,N_7191);
nand U8756 (N_8756,N_7409,N_7504);
nand U8757 (N_8757,N_7781,N_7651);
nand U8758 (N_8758,N_7451,N_7324);
or U8759 (N_8759,N_7369,N_7754);
or U8760 (N_8760,N_7725,N_7345);
xnor U8761 (N_8761,N_7928,N_7556);
and U8762 (N_8762,N_7012,N_7775);
nand U8763 (N_8763,N_7406,N_7433);
or U8764 (N_8764,N_7913,N_7911);
and U8765 (N_8765,N_7339,N_7488);
nand U8766 (N_8766,N_7138,N_7277);
and U8767 (N_8767,N_7225,N_7692);
nand U8768 (N_8768,N_7984,N_7950);
and U8769 (N_8769,N_7351,N_7283);
nand U8770 (N_8770,N_7172,N_7514);
or U8771 (N_8771,N_7272,N_7829);
and U8772 (N_8772,N_7370,N_7302);
nand U8773 (N_8773,N_7209,N_7876);
and U8774 (N_8774,N_7876,N_7472);
nor U8775 (N_8775,N_7921,N_7799);
nor U8776 (N_8776,N_7592,N_7838);
and U8777 (N_8777,N_7669,N_7165);
nor U8778 (N_8778,N_7430,N_7164);
nand U8779 (N_8779,N_7702,N_7815);
and U8780 (N_8780,N_7114,N_7845);
nor U8781 (N_8781,N_7466,N_7748);
or U8782 (N_8782,N_7766,N_7133);
nand U8783 (N_8783,N_7437,N_7922);
nand U8784 (N_8784,N_7588,N_7331);
or U8785 (N_8785,N_7499,N_7983);
and U8786 (N_8786,N_7186,N_7316);
nor U8787 (N_8787,N_7230,N_7190);
and U8788 (N_8788,N_7290,N_7105);
or U8789 (N_8789,N_7419,N_7413);
nor U8790 (N_8790,N_7405,N_7286);
nand U8791 (N_8791,N_7903,N_7774);
or U8792 (N_8792,N_7086,N_7550);
nor U8793 (N_8793,N_7469,N_7156);
nor U8794 (N_8794,N_7657,N_7610);
xor U8795 (N_8795,N_7143,N_7724);
or U8796 (N_8796,N_7333,N_7907);
nand U8797 (N_8797,N_7200,N_7645);
nor U8798 (N_8798,N_7163,N_7447);
and U8799 (N_8799,N_7578,N_7649);
xor U8800 (N_8800,N_7536,N_7199);
nand U8801 (N_8801,N_7438,N_7507);
xor U8802 (N_8802,N_7684,N_7970);
xnor U8803 (N_8803,N_7493,N_7295);
and U8804 (N_8804,N_7322,N_7449);
or U8805 (N_8805,N_7186,N_7664);
or U8806 (N_8806,N_7578,N_7081);
nor U8807 (N_8807,N_7445,N_7940);
or U8808 (N_8808,N_7673,N_7301);
nand U8809 (N_8809,N_7596,N_7411);
and U8810 (N_8810,N_7090,N_7940);
nand U8811 (N_8811,N_7121,N_7300);
nor U8812 (N_8812,N_7604,N_7101);
nor U8813 (N_8813,N_7126,N_7344);
nor U8814 (N_8814,N_7462,N_7355);
or U8815 (N_8815,N_7739,N_7995);
nor U8816 (N_8816,N_7666,N_7048);
or U8817 (N_8817,N_7763,N_7607);
nand U8818 (N_8818,N_7487,N_7674);
nor U8819 (N_8819,N_7247,N_7015);
and U8820 (N_8820,N_7011,N_7111);
and U8821 (N_8821,N_7088,N_7917);
and U8822 (N_8822,N_7316,N_7082);
and U8823 (N_8823,N_7810,N_7060);
or U8824 (N_8824,N_7163,N_7776);
or U8825 (N_8825,N_7441,N_7400);
or U8826 (N_8826,N_7316,N_7880);
and U8827 (N_8827,N_7321,N_7408);
and U8828 (N_8828,N_7210,N_7258);
xnor U8829 (N_8829,N_7374,N_7461);
and U8830 (N_8830,N_7062,N_7693);
nand U8831 (N_8831,N_7989,N_7141);
xnor U8832 (N_8832,N_7618,N_7178);
and U8833 (N_8833,N_7580,N_7300);
and U8834 (N_8834,N_7129,N_7287);
nand U8835 (N_8835,N_7264,N_7507);
or U8836 (N_8836,N_7778,N_7617);
nor U8837 (N_8837,N_7915,N_7039);
nor U8838 (N_8838,N_7080,N_7073);
nor U8839 (N_8839,N_7083,N_7088);
and U8840 (N_8840,N_7356,N_7605);
nor U8841 (N_8841,N_7367,N_7192);
and U8842 (N_8842,N_7548,N_7572);
xnor U8843 (N_8843,N_7116,N_7393);
or U8844 (N_8844,N_7555,N_7882);
nor U8845 (N_8845,N_7100,N_7927);
and U8846 (N_8846,N_7365,N_7094);
nor U8847 (N_8847,N_7275,N_7049);
nand U8848 (N_8848,N_7242,N_7078);
nor U8849 (N_8849,N_7431,N_7845);
and U8850 (N_8850,N_7014,N_7256);
nor U8851 (N_8851,N_7049,N_7240);
nand U8852 (N_8852,N_7692,N_7730);
nand U8853 (N_8853,N_7233,N_7109);
nand U8854 (N_8854,N_7628,N_7113);
or U8855 (N_8855,N_7179,N_7551);
nor U8856 (N_8856,N_7051,N_7953);
nor U8857 (N_8857,N_7331,N_7078);
and U8858 (N_8858,N_7761,N_7826);
nor U8859 (N_8859,N_7693,N_7929);
xnor U8860 (N_8860,N_7932,N_7964);
nand U8861 (N_8861,N_7808,N_7058);
and U8862 (N_8862,N_7259,N_7145);
or U8863 (N_8863,N_7705,N_7105);
xnor U8864 (N_8864,N_7206,N_7906);
nand U8865 (N_8865,N_7036,N_7275);
nor U8866 (N_8866,N_7364,N_7767);
or U8867 (N_8867,N_7976,N_7139);
nand U8868 (N_8868,N_7192,N_7844);
nor U8869 (N_8869,N_7663,N_7928);
or U8870 (N_8870,N_7137,N_7398);
and U8871 (N_8871,N_7600,N_7828);
or U8872 (N_8872,N_7759,N_7252);
or U8873 (N_8873,N_7943,N_7014);
xor U8874 (N_8874,N_7046,N_7566);
or U8875 (N_8875,N_7698,N_7233);
nor U8876 (N_8876,N_7442,N_7250);
or U8877 (N_8877,N_7359,N_7148);
nor U8878 (N_8878,N_7122,N_7757);
nand U8879 (N_8879,N_7776,N_7862);
or U8880 (N_8880,N_7904,N_7218);
nor U8881 (N_8881,N_7550,N_7545);
or U8882 (N_8882,N_7506,N_7309);
nand U8883 (N_8883,N_7827,N_7902);
or U8884 (N_8884,N_7516,N_7237);
xor U8885 (N_8885,N_7928,N_7896);
and U8886 (N_8886,N_7264,N_7272);
nor U8887 (N_8887,N_7902,N_7306);
nor U8888 (N_8888,N_7679,N_7815);
nor U8889 (N_8889,N_7705,N_7742);
or U8890 (N_8890,N_7400,N_7580);
or U8891 (N_8891,N_7076,N_7975);
xor U8892 (N_8892,N_7163,N_7687);
nand U8893 (N_8893,N_7829,N_7725);
nand U8894 (N_8894,N_7149,N_7696);
nor U8895 (N_8895,N_7950,N_7782);
and U8896 (N_8896,N_7206,N_7734);
and U8897 (N_8897,N_7908,N_7486);
or U8898 (N_8898,N_7706,N_7970);
or U8899 (N_8899,N_7846,N_7253);
nand U8900 (N_8900,N_7992,N_7266);
and U8901 (N_8901,N_7230,N_7883);
and U8902 (N_8902,N_7893,N_7261);
nand U8903 (N_8903,N_7175,N_7930);
and U8904 (N_8904,N_7720,N_7857);
or U8905 (N_8905,N_7793,N_7313);
and U8906 (N_8906,N_7694,N_7654);
or U8907 (N_8907,N_7681,N_7772);
and U8908 (N_8908,N_7058,N_7036);
xnor U8909 (N_8909,N_7536,N_7538);
nor U8910 (N_8910,N_7436,N_7432);
nor U8911 (N_8911,N_7561,N_7602);
nand U8912 (N_8912,N_7071,N_7369);
xnor U8913 (N_8913,N_7798,N_7695);
and U8914 (N_8914,N_7588,N_7801);
nor U8915 (N_8915,N_7846,N_7402);
or U8916 (N_8916,N_7845,N_7800);
nand U8917 (N_8917,N_7203,N_7254);
nand U8918 (N_8918,N_7418,N_7287);
nand U8919 (N_8919,N_7252,N_7773);
and U8920 (N_8920,N_7481,N_7437);
and U8921 (N_8921,N_7677,N_7760);
nand U8922 (N_8922,N_7980,N_7556);
nor U8923 (N_8923,N_7734,N_7442);
nor U8924 (N_8924,N_7565,N_7961);
xnor U8925 (N_8925,N_7362,N_7506);
nor U8926 (N_8926,N_7355,N_7077);
or U8927 (N_8927,N_7145,N_7967);
nor U8928 (N_8928,N_7399,N_7130);
and U8929 (N_8929,N_7577,N_7659);
nor U8930 (N_8930,N_7509,N_7768);
and U8931 (N_8931,N_7762,N_7441);
nor U8932 (N_8932,N_7396,N_7074);
nand U8933 (N_8933,N_7243,N_7202);
or U8934 (N_8934,N_7995,N_7570);
nor U8935 (N_8935,N_7675,N_7401);
and U8936 (N_8936,N_7285,N_7591);
xor U8937 (N_8937,N_7673,N_7228);
or U8938 (N_8938,N_7384,N_7578);
or U8939 (N_8939,N_7694,N_7210);
nor U8940 (N_8940,N_7409,N_7037);
nand U8941 (N_8941,N_7260,N_7037);
nand U8942 (N_8942,N_7111,N_7545);
nand U8943 (N_8943,N_7961,N_7440);
nand U8944 (N_8944,N_7715,N_7977);
nand U8945 (N_8945,N_7916,N_7377);
and U8946 (N_8946,N_7478,N_7064);
and U8947 (N_8947,N_7618,N_7277);
nor U8948 (N_8948,N_7791,N_7305);
nand U8949 (N_8949,N_7214,N_7359);
nand U8950 (N_8950,N_7137,N_7417);
or U8951 (N_8951,N_7564,N_7714);
xnor U8952 (N_8952,N_7812,N_7982);
xor U8953 (N_8953,N_7487,N_7795);
and U8954 (N_8954,N_7041,N_7826);
and U8955 (N_8955,N_7275,N_7163);
nand U8956 (N_8956,N_7919,N_7361);
or U8957 (N_8957,N_7637,N_7125);
nand U8958 (N_8958,N_7121,N_7744);
nand U8959 (N_8959,N_7221,N_7313);
and U8960 (N_8960,N_7419,N_7577);
nand U8961 (N_8961,N_7168,N_7546);
nor U8962 (N_8962,N_7797,N_7881);
nor U8963 (N_8963,N_7990,N_7681);
or U8964 (N_8964,N_7141,N_7673);
nor U8965 (N_8965,N_7589,N_7130);
xnor U8966 (N_8966,N_7079,N_7329);
nand U8967 (N_8967,N_7023,N_7134);
nor U8968 (N_8968,N_7038,N_7840);
xor U8969 (N_8969,N_7767,N_7049);
or U8970 (N_8970,N_7646,N_7053);
or U8971 (N_8971,N_7359,N_7893);
nand U8972 (N_8972,N_7836,N_7606);
xor U8973 (N_8973,N_7209,N_7403);
and U8974 (N_8974,N_7575,N_7758);
xor U8975 (N_8975,N_7078,N_7420);
nor U8976 (N_8976,N_7792,N_7278);
nor U8977 (N_8977,N_7780,N_7457);
xnor U8978 (N_8978,N_7621,N_7630);
nand U8979 (N_8979,N_7730,N_7752);
nor U8980 (N_8980,N_7898,N_7461);
nor U8981 (N_8981,N_7558,N_7757);
nor U8982 (N_8982,N_7933,N_7724);
and U8983 (N_8983,N_7640,N_7898);
nand U8984 (N_8984,N_7144,N_7507);
or U8985 (N_8985,N_7770,N_7527);
nand U8986 (N_8986,N_7918,N_7491);
nand U8987 (N_8987,N_7803,N_7505);
and U8988 (N_8988,N_7918,N_7608);
nand U8989 (N_8989,N_7369,N_7099);
nor U8990 (N_8990,N_7038,N_7291);
nand U8991 (N_8991,N_7956,N_7888);
or U8992 (N_8992,N_7407,N_7380);
nor U8993 (N_8993,N_7116,N_7910);
nand U8994 (N_8994,N_7248,N_7619);
or U8995 (N_8995,N_7902,N_7228);
nand U8996 (N_8996,N_7967,N_7959);
and U8997 (N_8997,N_7100,N_7864);
nand U8998 (N_8998,N_7701,N_7387);
and U8999 (N_8999,N_7625,N_7478);
or U9000 (N_9000,N_8081,N_8675);
nor U9001 (N_9001,N_8176,N_8602);
nor U9002 (N_9002,N_8358,N_8731);
xnor U9003 (N_9003,N_8007,N_8540);
and U9004 (N_9004,N_8877,N_8080);
nand U9005 (N_9005,N_8534,N_8630);
and U9006 (N_9006,N_8656,N_8252);
nand U9007 (N_9007,N_8728,N_8657);
or U9008 (N_9008,N_8891,N_8855);
and U9009 (N_9009,N_8191,N_8320);
and U9010 (N_9010,N_8830,N_8350);
nand U9011 (N_9011,N_8392,N_8142);
or U9012 (N_9012,N_8973,N_8061);
nand U9013 (N_9013,N_8233,N_8687);
nand U9014 (N_9014,N_8296,N_8634);
or U9015 (N_9015,N_8663,N_8902);
nor U9016 (N_9016,N_8418,N_8098);
or U9017 (N_9017,N_8453,N_8118);
and U9018 (N_9018,N_8648,N_8730);
or U9019 (N_9019,N_8138,N_8203);
xnor U9020 (N_9020,N_8765,N_8958);
nor U9021 (N_9021,N_8810,N_8809);
nand U9022 (N_9022,N_8658,N_8521);
or U9023 (N_9023,N_8890,N_8088);
or U9024 (N_9024,N_8063,N_8395);
and U9025 (N_9025,N_8366,N_8002);
and U9026 (N_9026,N_8977,N_8225);
and U9027 (N_9027,N_8404,N_8122);
and U9028 (N_9028,N_8747,N_8722);
nor U9029 (N_9029,N_8432,N_8825);
or U9030 (N_9030,N_8172,N_8889);
and U9031 (N_9031,N_8433,N_8427);
nor U9032 (N_9032,N_8368,N_8413);
and U9033 (N_9033,N_8489,N_8270);
nand U9034 (N_9034,N_8504,N_8393);
and U9035 (N_9035,N_8463,N_8802);
nand U9036 (N_9036,N_8471,N_8506);
nor U9037 (N_9037,N_8291,N_8502);
nand U9038 (N_9038,N_8562,N_8935);
nand U9039 (N_9039,N_8120,N_8982);
and U9040 (N_9040,N_8068,N_8171);
xor U9041 (N_9041,N_8072,N_8460);
or U9042 (N_9042,N_8922,N_8603);
nand U9043 (N_9043,N_8276,N_8208);
nor U9044 (N_9044,N_8607,N_8929);
xor U9045 (N_9045,N_8420,N_8700);
or U9046 (N_9046,N_8292,N_8328);
nor U9047 (N_9047,N_8157,N_8381);
or U9048 (N_9048,N_8783,N_8874);
nor U9049 (N_9049,N_8965,N_8859);
or U9050 (N_9050,N_8762,N_8447);
nand U9051 (N_9051,N_8019,N_8078);
and U9052 (N_9052,N_8455,N_8197);
nand U9053 (N_9053,N_8593,N_8375);
or U9054 (N_9054,N_8582,N_8136);
nor U9055 (N_9055,N_8569,N_8649);
nand U9056 (N_9056,N_8016,N_8341);
and U9057 (N_9057,N_8570,N_8234);
nand U9058 (N_9058,N_8175,N_8268);
xor U9059 (N_9059,N_8969,N_8846);
and U9060 (N_9060,N_8373,N_8446);
nor U9061 (N_9061,N_8949,N_8133);
nor U9062 (N_9062,N_8772,N_8986);
and U9063 (N_9063,N_8071,N_8355);
or U9064 (N_9064,N_8470,N_8134);
or U9065 (N_9065,N_8140,N_8469);
or U9066 (N_9066,N_8887,N_8000);
nand U9067 (N_9067,N_8548,N_8474);
or U9068 (N_9068,N_8815,N_8983);
and U9069 (N_9069,N_8131,N_8883);
or U9070 (N_9070,N_8106,N_8340);
nand U9071 (N_9071,N_8031,N_8238);
and U9072 (N_9072,N_8995,N_8386);
and U9073 (N_9073,N_8147,N_8263);
or U9074 (N_9074,N_8561,N_8259);
nand U9075 (N_9075,N_8465,N_8996);
or U9076 (N_9076,N_8636,N_8339);
or U9077 (N_9077,N_8376,N_8187);
nor U9078 (N_9078,N_8261,N_8725);
nor U9079 (N_9079,N_8060,N_8854);
nand U9080 (N_9080,N_8492,N_8679);
nor U9081 (N_9081,N_8242,N_8847);
nand U9082 (N_9082,N_8473,N_8479);
or U9083 (N_9083,N_8039,N_8050);
nor U9084 (N_9084,N_8613,N_8978);
nand U9085 (N_9085,N_8149,N_8091);
nor U9086 (N_9086,N_8827,N_8262);
nor U9087 (N_9087,N_8835,N_8006);
xor U9088 (N_9088,N_8584,N_8282);
nor U9089 (N_9089,N_8462,N_8312);
nand U9090 (N_9090,N_8024,N_8037);
or U9091 (N_9091,N_8638,N_8493);
nand U9092 (N_9092,N_8383,N_8975);
xor U9093 (N_9093,N_8867,N_8084);
nor U9094 (N_9094,N_8338,N_8755);
and U9095 (N_9095,N_8763,N_8070);
and U9096 (N_9096,N_8448,N_8673);
and U9097 (N_9097,N_8522,N_8415);
or U9098 (N_9098,N_8429,N_8936);
nor U9099 (N_9099,N_8216,N_8255);
xnor U9100 (N_9100,N_8573,N_8436);
xor U9101 (N_9101,N_8293,N_8269);
nor U9102 (N_9102,N_8974,N_8520);
xor U9103 (N_9103,N_8198,N_8403);
or U9104 (N_9104,N_8004,N_8507);
and U9105 (N_9105,N_8440,N_8124);
nand U9106 (N_9106,N_8742,N_8665);
and U9107 (N_9107,N_8464,N_8989);
nor U9108 (N_9108,N_8231,N_8287);
or U9109 (N_9109,N_8457,N_8653);
or U9110 (N_9110,N_8500,N_8150);
or U9111 (N_9111,N_8606,N_8530);
or U9112 (N_9112,N_8964,N_8499);
nor U9113 (N_9113,N_8524,N_8597);
nand U9114 (N_9114,N_8402,N_8536);
or U9115 (N_9115,N_8456,N_8369);
nand U9116 (N_9116,N_8842,N_8260);
nor U9117 (N_9117,N_8750,N_8025);
or U9118 (N_9118,N_8953,N_8832);
xor U9119 (N_9119,N_8820,N_8876);
and U9120 (N_9120,N_8034,N_8184);
nor U9121 (N_9121,N_8099,N_8289);
or U9122 (N_9122,N_8871,N_8181);
nor U9123 (N_9123,N_8711,N_8856);
nor U9124 (N_9124,N_8961,N_8498);
or U9125 (N_9125,N_8999,N_8738);
nor U9126 (N_9126,N_8545,N_8523);
and U9127 (N_9127,N_8159,N_8107);
or U9128 (N_9128,N_8012,N_8170);
nor U9129 (N_9129,N_8863,N_8645);
nor U9130 (N_9130,N_8659,N_8706);
nand U9131 (N_9131,N_8406,N_8343);
nor U9132 (N_9132,N_8752,N_8251);
nor U9133 (N_9133,N_8941,N_8860);
or U9134 (N_9134,N_8027,N_8219);
or U9135 (N_9135,N_8180,N_8516);
nor U9136 (N_9136,N_8167,N_8563);
nand U9137 (N_9137,N_8839,N_8614);
or U9138 (N_9138,N_8049,N_8821);
nor U9139 (N_9139,N_8608,N_8271);
or U9140 (N_9140,N_8724,N_8051);
nor U9141 (N_9141,N_8549,N_8074);
nor U9142 (N_9142,N_8277,N_8990);
and U9143 (N_9143,N_8962,N_8959);
nand U9144 (N_9144,N_8344,N_8151);
nand U9145 (N_9145,N_8193,N_8680);
nor U9146 (N_9146,N_8513,N_8212);
nor U9147 (N_9147,N_8957,N_8458);
nand U9148 (N_9148,N_8301,N_8577);
and U9149 (N_9149,N_8664,N_8230);
nor U9150 (N_9150,N_8115,N_8773);
or U9151 (N_9151,N_8558,N_8250);
nand U9152 (N_9152,N_8955,N_8623);
xnor U9153 (N_9153,N_8137,N_8713);
or U9154 (N_9154,N_8079,N_8154);
nand U9155 (N_9155,N_8574,N_8192);
nand U9156 (N_9156,N_8278,N_8698);
and U9157 (N_9157,N_8281,N_8111);
nor U9158 (N_9158,N_8880,N_8984);
and U9159 (N_9159,N_8315,N_8550);
and U9160 (N_9160,N_8073,N_8719);
nor U9161 (N_9161,N_8491,N_8472);
or U9162 (N_9162,N_8654,N_8266);
and U9163 (N_9163,N_8003,N_8946);
or U9164 (N_9164,N_8591,N_8518);
or U9165 (N_9165,N_8644,N_8800);
or U9166 (N_9166,N_8824,N_8786);
and U9167 (N_9167,N_8617,N_8696);
nor U9168 (N_9168,N_8162,N_8590);
nor U9169 (N_9169,N_8611,N_8861);
nand U9170 (N_9170,N_8533,N_8241);
and U9171 (N_9171,N_8991,N_8714);
nor U9172 (N_9172,N_8411,N_8298);
nand U9173 (N_9173,N_8560,N_8264);
nor U9174 (N_9174,N_8834,N_8442);
nand U9175 (N_9175,N_8914,N_8308);
and U9176 (N_9176,N_8405,N_8626);
or U9177 (N_9177,N_8886,N_8580);
or U9178 (N_9178,N_8741,N_8677);
or U9179 (N_9179,N_8330,N_8173);
and U9180 (N_9180,N_8352,N_8213);
xor U9181 (N_9181,N_8697,N_8791);
or U9182 (N_9182,N_8319,N_8110);
and U9183 (N_9183,N_8754,N_8923);
and U9184 (N_9184,N_8888,N_8588);
nand U9185 (N_9185,N_8417,N_8721);
nor U9186 (N_9186,N_8908,N_8655);
or U9187 (N_9187,N_8937,N_8477);
nor U9188 (N_9188,N_8112,N_8579);
xor U9189 (N_9189,N_8356,N_8015);
or U9190 (N_9190,N_8723,N_8158);
and U9191 (N_9191,N_8589,N_8954);
and U9192 (N_9192,N_8629,N_8042);
and U9193 (N_9193,N_8503,N_8426);
nand U9194 (N_9194,N_8089,N_8085);
nand U9195 (N_9195,N_8913,N_8650);
nand U9196 (N_9196,N_8703,N_8912);
xor U9197 (N_9197,N_8434,N_8734);
or U9198 (N_9198,N_8598,N_8535);
and U9199 (N_9199,N_8988,N_8904);
or U9200 (N_9200,N_8667,N_8612);
nand U9201 (N_9201,N_8214,N_8481);
nand U9202 (N_9202,N_8565,N_8852);
and U9203 (N_9203,N_8485,N_8808);
nor U9204 (N_9204,N_8926,N_8186);
or U9205 (N_9205,N_8285,N_8310);
or U9206 (N_9206,N_8148,N_8021);
nor U9207 (N_9207,N_8666,N_8218);
nor U9208 (N_9208,N_8040,N_8119);
and U9209 (N_9209,N_8512,N_8057);
nor U9210 (N_9210,N_8105,N_8280);
xor U9211 (N_9211,N_8254,N_8726);
and U9212 (N_9212,N_8985,N_8439);
nand U9213 (N_9213,N_8660,N_8622);
nor U9214 (N_9214,N_8304,N_8793);
or U9215 (N_9215,N_8971,N_8114);
nor U9216 (N_9216,N_8715,N_8998);
nand U9217 (N_9217,N_8733,N_8831);
nand U9218 (N_9218,N_8360,N_8921);
nand U9219 (N_9219,N_8807,N_8302);
and U9220 (N_9220,N_8695,N_8275);
xor U9221 (N_9221,N_8435,N_8782);
nand U9222 (N_9222,N_8497,N_8910);
and U9223 (N_9223,N_8768,N_8979);
and U9224 (N_9224,N_8235,N_8424);
xnor U9225 (N_9225,N_8062,N_8215);
or U9226 (N_9226,N_8684,N_8746);
or U9227 (N_9227,N_8717,N_8482);
xor U9228 (N_9228,N_8316,N_8348);
and U9229 (N_9229,N_8920,N_8314);
and U9230 (N_9230,N_8283,N_8380);
or U9231 (N_9231,N_8257,N_8325);
and U9232 (N_9232,N_8190,N_8948);
or U9233 (N_9233,N_8329,N_8211);
nand U9234 (N_9234,N_8097,N_8100);
nand U9235 (N_9235,N_8798,N_8519);
or U9236 (N_9236,N_8539,N_8378);
nor U9237 (N_9237,N_8844,N_8610);
nor U9238 (N_9238,N_8616,N_8770);
or U9239 (N_9239,N_8430,N_8224);
nand U9240 (N_9240,N_8661,N_8875);
or U9241 (N_9241,N_8682,N_8841);
nor U9242 (N_9242,N_8884,N_8940);
and U9243 (N_9243,N_8384,N_8592);
nand U9244 (N_9244,N_8299,N_8764);
or U9245 (N_9245,N_8868,N_8774);
and U9246 (N_9246,N_8103,N_8641);
nand U9247 (N_9247,N_8438,N_8357);
nor U9248 (N_9248,N_8001,N_8372);
or U9249 (N_9249,N_8748,N_8163);
and U9250 (N_9250,N_8639,N_8419);
nand U9251 (N_9251,N_8605,N_8478);
nor U9252 (N_9252,N_8531,N_8652);
nor U9253 (N_9253,N_8688,N_8576);
and U9254 (N_9254,N_8567,N_8305);
nand U9255 (N_9255,N_8056,N_8745);
xnor U9256 (N_9256,N_8146,N_8803);
or U9257 (N_9257,N_8496,N_8526);
or U9258 (N_9258,N_8422,N_8981);
or U9259 (N_9259,N_8394,N_8155);
nand U9260 (N_9260,N_8253,N_8421);
and U9261 (N_9261,N_8317,N_8609);
or U9262 (N_9262,N_8126,N_8952);
or U9263 (N_9263,N_8351,N_8692);
nor U9264 (N_9264,N_8327,N_8205);
nand U9265 (N_9265,N_8113,N_8178);
and U9266 (N_9266,N_8288,N_8409);
and U9267 (N_9267,N_8484,N_8399);
and U9268 (N_9268,N_8572,N_8704);
xor U9269 (N_9269,N_8020,N_8347);
and U9270 (N_9270,N_8541,N_8443);
nor U9271 (N_9271,N_8836,N_8221);
nand U9272 (N_9272,N_8515,N_8766);
nor U9273 (N_9273,N_8236,N_8220);
xor U9274 (N_9274,N_8934,N_8087);
nor U9275 (N_9275,N_8761,N_8365);
nand U9276 (N_9276,N_8248,N_8416);
nor U9277 (N_9277,N_8053,N_8525);
or U9278 (N_9278,N_8321,N_8812);
nor U9279 (N_9279,N_8200,N_8086);
and U9280 (N_9280,N_8297,N_8045);
nand U9281 (N_9281,N_8017,N_8177);
nor U9282 (N_9282,N_8968,N_8813);
nor U9283 (N_9283,N_8632,N_8223);
and U9284 (N_9284,N_8538,N_8950);
xnor U9285 (N_9285,N_8780,N_8740);
and U9286 (N_9286,N_8082,N_8547);
nor U9287 (N_9287,N_8795,N_8128);
xor U9288 (N_9288,N_8095,N_8945);
nand U9289 (N_9289,N_8685,N_8129);
nor U9290 (N_9290,N_8851,N_8705);
or U9291 (N_9291,N_8816,N_8486);
xor U9292 (N_9292,N_8127,N_8686);
nand U9293 (N_9293,N_8942,N_8054);
and U9294 (N_9294,N_8182,N_8787);
or U9295 (N_9295,N_8967,N_8651);
nor U9296 (N_9296,N_8454,N_8374);
and U9297 (N_9297,N_8267,N_8028);
nor U9298 (N_9298,N_8823,N_8806);
nand U9299 (N_9299,N_8640,N_8370);
or U9300 (N_9300,N_8274,N_8067);
xnor U9301 (N_9301,N_8425,N_8326);
nor U9302 (N_9302,N_8872,N_8094);
nand U9303 (N_9303,N_8345,N_8822);
and U9304 (N_9304,N_8771,N_8188);
nand U9305 (N_9305,N_8707,N_8928);
nor U9306 (N_9306,N_8501,N_8833);
xor U9307 (N_9307,N_8153,N_8508);
or U9308 (N_9308,N_8033,N_8487);
or U9309 (N_9309,N_8681,N_8244);
xnor U9310 (N_9310,N_8618,N_8619);
or U9311 (N_9311,N_8690,N_8898);
and U9312 (N_9312,N_8691,N_8792);
nor U9313 (N_9313,N_8749,N_8599);
nor U9314 (N_9314,N_8564,N_8776);
nor U9315 (N_9315,N_8866,N_8018);
nor U9316 (N_9316,N_8896,N_8398);
or U9317 (N_9317,N_8899,N_8010);
or U9318 (N_9318,N_8966,N_8169);
nor U9319 (N_9319,N_8699,N_8354);
nand U9320 (N_9320,N_8805,N_8595);
or U9321 (N_9321,N_8165,N_8843);
nand U9322 (N_9322,N_8537,N_8226);
or U9323 (N_9323,N_8869,N_8108);
nand U9324 (N_9324,N_8359,N_8583);
or U9325 (N_9325,N_8029,N_8207);
or U9326 (N_9326,N_8647,N_8475);
nand U9327 (N_9327,N_8444,N_8390);
nor U9328 (N_9328,N_8069,N_8014);
or U9329 (N_9329,N_8139,N_8272);
nand U9330 (N_9330,N_8911,N_8760);
nor U9331 (N_9331,N_8837,N_8038);
or U9332 (N_9332,N_8581,N_8865);
nand U9333 (N_9333,N_8044,N_8013);
nand U9334 (N_9334,N_8976,N_8382);
nand U9335 (N_9335,N_8311,N_8817);
or U9336 (N_9336,N_8052,N_8468);
and U9337 (N_9337,N_8735,N_8870);
or U9338 (N_9338,N_8412,N_8845);
or U9339 (N_9339,N_8552,N_8273);
and U9340 (N_9340,N_8461,N_8718);
nand U9341 (N_9341,N_8228,N_8585);
or U9342 (N_9342,N_8919,N_8757);
nor U9343 (N_9343,N_8960,N_8363);
nor U9344 (N_9344,N_8206,N_8970);
and U9345 (N_9345,N_8026,N_8195);
xor U9346 (N_9346,N_8410,N_8318);
and U9347 (N_9347,N_8727,N_8441);
xor U9348 (N_9348,N_8391,N_8232);
or U9349 (N_9349,N_8878,N_8769);
and U9350 (N_9350,N_8209,N_8668);
and U9351 (N_9351,N_8451,N_8756);
or U9352 (N_9352,N_8559,N_8011);
or U9353 (N_9353,N_8848,N_8729);
nor U9354 (N_9354,N_8488,N_8586);
nor U9355 (N_9355,N_8437,N_8575);
or U9356 (N_9356,N_8939,N_8125);
or U9357 (N_9357,N_8801,N_8938);
xnor U9358 (N_9358,N_8881,N_8838);
nand U9359 (N_9359,N_8222,N_8217);
and U9360 (N_9360,N_8005,N_8712);
nand U9361 (N_9361,N_8514,N_8237);
xor U9362 (N_9362,N_8396,N_8553);
nor U9363 (N_9363,N_8956,N_8494);
nand U9364 (N_9364,N_8643,N_8388);
nor U9365 (N_9365,N_8483,N_8947);
and U9366 (N_9366,N_8096,N_8882);
xnor U9367 (N_9367,N_8900,N_8543);
or U9368 (N_9368,N_8879,N_8450);
and U9369 (N_9369,N_8035,N_8055);
xor U9370 (N_9370,N_8849,N_8737);
nand U9371 (N_9371,N_8059,N_8145);
or U9372 (N_9372,N_8030,N_8240);
or U9373 (N_9373,N_8116,N_8322);
and U9374 (N_9374,N_8303,N_8306);
nand U9375 (N_9375,N_8710,N_8332);
or U9376 (N_9376,N_8646,N_8490);
and U9377 (N_9377,N_8279,N_8143);
nor U9378 (N_9378,N_8864,N_8290);
nor U9379 (N_9379,N_8987,N_8708);
nor U9380 (N_9380,N_8117,N_8371);
and U9381 (N_9381,N_8788,N_8972);
or U9382 (N_9382,N_8048,N_8930);
nand U9383 (N_9383,N_8229,N_8627);
nor U9384 (N_9384,N_8980,N_8334);
nand U9385 (N_9385,N_8065,N_8924);
and U9386 (N_9386,N_8933,N_8452);
nor U9387 (N_9387,N_8633,N_8850);
or U9388 (N_9388,N_8245,N_8092);
nand U9389 (N_9389,N_8596,N_8389);
nor U9390 (N_9390,N_8476,N_8909);
or U9391 (N_9391,N_8367,N_8046);
and U9392 (N_9392,N_8775,N_8022);
nand U9393 (N_9393,N_8336,N_8379);
nand U9394 (N_9394,N_8032,N_8739);
nor U9395 (N_9395,N_8799,N_8858);
nor U9396 (N_9396,N_8578,N_8510);
or U9397 (N_9397,N_8732,N_8152);
nand U9398 (N_9398,N_8642,N_8784);
xnor U9399 (N_9399,N_8313,N_8628);
and U9400 (N_9400,N_8509,N_8227);
and U9401 (N_9401,N_8683,N_8135);
and U9402 (N_9402,N_8265,N_8814);
and U9403 (N_9403,N_8790,N_8480);
nand U9404 (N_9404,N_8058,N_8556);
and U9405 (N_9405,N_8511,N_8323);
and U9406 (N_9406,N_8594,N_8551);
nor U9407 (N_9407,N_8785,N_8467);
nand U9408 (N_9408,N_8546,N_8885);
nor U9409 (N_9409,N_8294,N_8342);
nor U9410 (N_9410,N_8179,N_8566);
or U9411 (N_9411,N_8362,N_8353);
nor U9412 (N_9412,N_8604,N_8075);
xor U9413 (N_9413,N_8615,N_8571);
nor U9414 (N_9414,N_8963,N_8797);
and U9415 (N_9415,N_8166,N_8532);
nand U9416 (N_9416,N_8174,N_8401);
nor U9417 (N_9417,N_8694,N_8529);
and U9418 (N_9418,N_8066,N_8811);
and U9419 (N_9419,N_8943,N_8104);
nand U9420 (N_9420,N_8631,N_8853);
or U9421 (N_9421,N_8123,N_8702);
nand U9422 (N_9422,N_8121,N_8753);
nor U9423 (N_9423,N_8204,N_8720);
nand U9424 (N_9424,N_8333,N_8689);
or U9425 (N_9425,N_8466,N_8161);
and U9426 (N_9426,N_8408,N_8400);
and U9427 (N_9427,N_8777,N_8751);
nor U9428 (N_9428,N_8160,N_8758);
or U9429 (N_9429,N_8101,N_8701);
xor U9430 (N_9430,N_8047,N_8361);
or U9431 (N_9431,N_8894,N_8385);
xnor U9432 (N_9432,N_8246,N_8199);
xor U9433 (N_9433,N_8671,N_8672);
and U9434 (N_9434,N_8528,N_8132);
nand U9435 (N_9435,N_8625,N_8951);
nor U9436 (N_9436,N_8036,N_8678);
or U9437 (N_9437,N_8144,N_8693);
nand U9438 (N_9438,N_8109,N_8023);
xor U9439 (N_9439,N_8670,N_8944);
and U9440 (N_9440,N_8819,N_8256);
nor U9441 (N_9441,N_8992,N_8164);
nand U9442 (N_9442,N_8829,N_8637);
xnor U9443 (N_9443,N_8669,N_8239);
or U9444 (N_9444,N_8767,N_8445);
nand U9445 (N_9445,N_8295,N_8554);
xor U9446 (N_9446,N_8527,N_8892);
or U9447 (N_9447,N_8840,N_8620);
and U9448 (N_9448,N_8997,N_8423);
nor U9449 (N_9449,N_8041,N_8716);
nor U9450 (N_9450,N_8893,N_8709);
nor U9451 (N_9451,N_8505,N_8789);
nor U9452 (N_9452,N_8794,N_8781);
nand U9453 (N_9453,N_8243,N_8674);
or U9454 (N_9454,N_8857,N_8495);
nand U9455 (N_9455,N_8517,N_8736);
or U9456 (N_9456,N_8918,N_8778);
nor U9457 (N_9457,N_8544,N_8927);
nand U9458 (N_9458,N_8141,N_8587);
or U9459 (N_9459,N_8102,N_8459);
and U9460 (N_9460,N_8431,N_8258);
nor U9461 (N_9461,N_8090,N_8196);
nor U9462 (N_9462,N_8993,N_8093);
nor U9463 (N_9463,N_8168,N_8804);
or U9464 (N_9464,N_8568,N_8779);
or U9465 (N_9465,N_8915,N_8907);
nand U9466 (N_9466,N_8828,N_8300);
nor U9467 (N_9467,N_8183,N_8903);
or U9468 (N_9468,N_8635,N_8185);
or U9469 (N_9469,N_8895,N_8542);
xor U9470 (N_9470,N_8676,N_8008);
or U9471 (N_9471,N_8307,N_8917);
nor U9472 (N_9472,N_8194,N_8156);
nand U9473 (N_9473,N_8337,N_8009);
nor U9474 (N_9474,N_8906,N_8043);
or U9475 (N_9475,N_8083,N_8916);
and U9476 (N_9476,N_8796,N_8601);
and U9477 (N_9477,N_8324,N_8449);
or U9478 (N_9478,N_8897,N_8932);
nor U9479 (N_9479,N_8901,N_8130);
nor U9480 (N_9480,N_8284,N_8335);
nand U9481 (N_9481,N_8201,N_8077);
nor U9482 (N_9482,N_8202,N_8557);
and U9483 (N_9483,N_8309,N_8247);
xor U9484 (N_9484,N_8624,N_8210);
xnor U9485 (N_9485,N_8744,N_8349);
and U9486 (N_9486,N_8076,N_8621);
or U9487 (N_9487,N_8862,N_8743);
xnor U9488 (N_9488,N_8346,N_8397);
and U9489 (N_9489,N_8994,N_8925);
nor U9490 (N_9490,N_8377,N_8873);
or U9491 (N_9491,N_8826,N_8364);
nand U9492 (N_9492,N_8818,N_8286);
xor U9493 (N_9493,N_8414,N_8064);
nand U9494 (N_9494,N_8662,N_8387);
nor U9495 (N_9495,N_8905,N_8931);
and U9496 (N_9496,N_8249,N_8600);
and U9497 (N_9497,N_8759,N_8555);
nor U9498 (N_9498,N_8407,N_8331);
or U9499 (N_9499,N_8428,N_8189);
nand U9500 (N_9500,N_8911,N_8489);
and U9501 (N_9501,N_8624,N_8525);
nand U9502 (N_9502,N_8041,N_8959);
or U9503 (N_9503,N_8663,N_8717);
nand U9504 (N_9504,N_8447,N_8802);
and U9505 (N_9505,N_8596,N_8489);
or U9506 (N_9506,N_8949,N_8713);
xor U9507 (N_9507,N_8861,N_8653);
nor U9508 (N_9508,N_8524,N_8194);
nand U9509 (N_9509,N_8569,N_8111);
or U9510 (N_9510,N_8881,N_8266);
nor U9511 (N_9511,N_8236,N_8922);
and U9512 (N_9512,N_8507,N_8355);
or U9513 (N_9513,N_8146,N_8274);
nor U9514 (N_9514,N_8106,N_8430);
nor U9515 (N_9515,N_8761,N_8256);
nand U9516 (N_9516,N_8354,N_8967);
nor U9517 (N_9517,N_8592,N_8705);
nor U9518 (N_9518,N_8507,N_8638);
nand U9519 (N_9519,N_8100,N_8053);
nand U9520 (N_9520,N_8825,N_8177);
or U9521 (N_9521,N_8720,N_8635);
nor U9522 (N_9522,N_8977,N_8962);
and U9523 (N_9523,N_8615,N_8150);
nor U9524 (N_9524,N_8387,N_8728);
nand U9525 (N_9525,N_8945,N_8697);
nand U9526 (N_9526,N_8787,N_8468);
and U9527 (N_9527,N_8497,N_8179);
xnor U9528 (N_9528,N_8466,N_8944);
and U9529 (N_9529,N_8468,N_8859);
nor U9530 (N_9530,N_8746,N_8352);
or U9531 (N_9531,N_8511,N_8102);
nand U9532 (N_9532,N_8751,N_8613);
nor U9533 (N_9533,N_8498,N_8434);
or U9534 (N_9534,N_8716,N_8767);
and U9535 (N_9535,N_8921,N_8487);
nor U9536 (N_9536,N_8663,N_8328);
nand U9537 (N_9537,N_8315,N_8267);
and U9538 (N_9538,N_8110,N_8423);
nor U9539 (N_9539,N_8125,N_8667);
nor U9540 (N_9540,N_8156,N_8011);
nand U9541 (N_9541,N_8681,N_8615);
xnor U9542 (N_9542,N_8728,N_8827);
or U9543 (N_9543,N_8796,N_8923);
and U9544 (N_9544,N_8469,N_8104);
and U9545 (N_9545,N_8553,N_8299);
nand U9546 (N_9546,N_8550,N_8344);
nor U9547 (N_9547,N_8133,N_8623);
or U9548 (N_9548,N_8346,N_8960);
nor U9549 (N_9549,N_8444,N_8274);
and U9550 (N_9550,N_8300,N_8703);
and U9551 (N_9551,N_8298,N_8161);
nor U9552 (N_9552,N_8745,N_8197);
nor U9553 (N_9553,N_8755,N_8710);
nand U9554 (N_9554,N_8781,N_8472);
and U9555 (N_9555,N_8904,N_8209);
or U9556 (N_9556,N_8768,N_8798);
nor U9557 (N_9557,N_8831,N_8670);
nor U9558 (N_9558,N_8823,N_8507);
or U9559 (N_9559,N_8004,N_8540);
or U9560 (N_9560,N_8692,N_8378);
or U9561 (N_9561,N_8108,N_8943);
or U9562 (N_9562,N_8254,N_8529);
or U9563 (N_9563,N_8595,N_8817);
and U9564 (N_9564,N_8040,N_8030);
xnor U9565 (N_9565,N_8566,N_8433);
xor U9566 (N_9566,N_8141,N_8776);
nor U9567 (N_9567,N_8754,N_8264);
or U9568 (N_9568,N_8830,N_8998);
nand U9569 (N_9569,N_8813,N_8712);
nor U9570 (N_9570,N_8370,N_8341);
nand U9571 (N_9571,N_8538,N_8565);
and U9572 (N_9572,N_8867,N_8199);
nor U9573 (N_9573,N_8049,N_8688);
and U9574 (N_9574,N_8384,N_8368);
nor U9575 (N_9575,N_8331,N_8193);
or U9576 (N_9576,N_8835,N_8928);
nand U9577 (N_9577,N_8089,N_8280);
nor U9578 (N_9578,N_8041,N_8027);
nor U9579 (N_9579,N_8663,N_8155);
xor U9580 (N_9580,N_8552,N_8251);
nor U9581 (N_9581,N_8645,N_8916);
nand U9582 (N_9582,N_8614,N_8586);
or U9583 (N_9583,N_8426,N_8419);
nor U9584 (N_9584,N_8182,N_8342);
nand U9585 (N_9585,N_8774,N_8925);
xnor U9586 (N_9586,N_8044,N_8847);
nand U9587 (N_9587,N_8447,N_8047);
nor U9588 (N_9588,N_8035,N_8177);
nand U9589 (N_9589,N_8002,N_8020);
or U9590 (N_9590,N_8636,N_8330);
and U9591 (N_9591,N_8820,N_8904);
nor U9592 (N_9592,N_8242,N_8235);
xnor U9593 (N_9593,N_8104,N_8364);
nand U9594 (N_9594,N_8576,N_8061);
xnor U9595 (N_9595,N_8335,N_8959);
or U9596 (N_9596,N_8901,N_8058);
nor U9597 (N_9597,N_8474,N_8774);
and U9598 (N_9598,N_8534,N_8992);
xor U9599 (N_9599,N_8967,N_8353);
or U9600 (N_9600,N_8448,N_8627);
nand U9601 (N_9601,N_8074,N_8969);
or U9602 (N_9602,N_8607,N_8460);
or U9603 (N_9603,N_8395,N_8182);
nand U9604 (N_9604,N_8463,N_8828);
nor U9605 (N_9605,N_8658,N_8214);
and U9606 (N_9606,N_8822,N_8262);
and U9607 (N_9607,N_8035,N_8591);
or U9608 (N_9608,N_8523,N_8538);
and U9609 (N_9609,N_8075,N_8139);
nand U9610 (N_9610,N_8406,N_8139);
or U9611 (N_9611,N_8671,N_8378);
or U9612 (N_9612,N_8626,N_8779);
nor U9613 (N_9613,N_8945,N_8388);
or U9614 (N_9614,N_8343,N_8377);
and U9615 (N_9615,N_8640,N_8314);
nand U9616 (N_9616,N_8016,N_8682);
and U9617 (N_9617,N_8097,N_8083);
or U9618 (N_9618,N_8302,N_8642);
or U9619 (N_9619,N_8836,N_8008);
nand U9620 (N_9620,N_8261,N_8674);
nor U9621 (N_9621,N_8586,N_8721);
nor U9622 (N_9622,N_8549,N_8853);
or U9623 (N_9623,N_8414,N_8896);
nor U9624 (N_9624,N_8529,N_8557);
or U9625 (N_9625,N_8872,N_8758);
or U9626 (N_9626,N_8099,N_8647);
or U9627 (N_9627,N_8836,N_8865);
xor U9628 (N_9628,N_8847,N_8192);
and U9629 (N_9629,N_8462,N_8330);
nor U9630 (N_9630,N_8705,N_8825);
nand U9631 (N_9631,N_8252,N_8974);
nor U9632 (N_9632,N_8662,N_8055);
or U9633 (N_9633,N_8490,N_8934);
nor U9634 (N_9634,N_8008,N_8878);
nand U9635 (N_9635,N_8609,N_8683);
and U9636 (N_9636,N_8791,N_8556);
nand U9637 (N_9637,N_8920,N_8584);
and U9638 (N_9638,N_8262,N_8041);
xnor U9639 (N_9639,N_8409,N_8262);
nand U9640 (N_9640,N_8009,N_8587);
and U9641 (N_9641,N_8612,N_8075);
and U9642 (N_9642,N_8813,N_8768);
nor U9643 (N_9643,N_8789,N_8400);
and U9644 (N_9644,N_8263,N_8185);
nor U9645 (N_9645,N_8357,N_8389);
nor U9646 (N_9646,N_8898,N_8529);
nor U9647 (N_9647,N_8932,N_8950);
or U9648 (N_9648,N_8644,N_8792);
or U9649 (N_9649,N_8055,N_8749);
or U9650 (N_9650,N_8922,N_8554);
or U9651 (N_9651,N_8674,N_8885);
and U9652 (N_9652,N_8895,N_8207);
nor U9653 (N_9653,N_8965,N_8203);
xor U9654 (N_9654,N_8144,N_8783);
nand U9655 (N_9655,N_8729,N_8522);
nor U9656 (N_9656,N_8756,N_8944);
or U9657 (N_9657,N_8240,N_8459);
or U9658 (N_9658,N_8132,N_8870);
nand U9659 (N_9659,N_8922,N_8730);
nand U9660 (N_9660,N_8184,N_8486);
nand U9661 (N_9661,N_8596,N_8751);
nor U9662 (N_9662,N_8899,N_8702);
or U9663 (N_9663,N_8179,N_8372);
nor U9664 (N_9664,N_8539,N_8157);
or U9665 (N_9665,N_8811,N_8491);
nand U9666 (N_9666,N_8385,N_8211);
or U9667 (N_9667,N_8833,N_8450);
nand U9668 (N_9668,N_8870,N_8613);
nor U9669 (N_9669,N_8207,N_8220);
and U9670 (N_9670,N_8588,N_8786);
nand U9671 (N_9671,N_8969,N_8577);
or U9672 (N_9672,N_8369,N_8663);
nor U9673 (N_9673,N_8943,N_8131);
nor U9674 (N_9674,N_8226,N_8492);
and U9675 (N_9675,N_8116,N_8518);
nor U9676 (N_9676,N_8817,N_8887);
nand U9677 (N_9677,N_8049,N_8031);
or U9678 (N_9678,N_8970,N_8223);
nor U9679 (N_9679,N_8514,N_8177);
nand U9680 (N_9680,N_8600,N_8734);
xor U9681 (N_9681,N_8504,N_8965);
nor U9682 (N_9682,N_8698,N_8319);
and U9683 (N_9683,N_8208,N_8871);
and U9684 (N_9684,N_8790,N_8376);
and U9685 (N_9685,N_8130,N_8952);
nor U9686 (N_9686,N_8053,N_8499);
nand U9687 (N_9687,N_8459,N_8688);
and U9688 (N_9688,N_8349,N_8411);
nand U9689 (N_9689,N_8811,N_8101);
nand U9690 (N_9690,N_8391,N_8548);
or U9691 (N_9691,N_8463,N_8341);
or U9692 (N_9692,N_8903,N_8411);
or U9693 (N_9693,N_8876,N_8931);
nand U9694 (N_9694,N_8756,N_8879);
nor U9695 (N_9695,N_8785,N_8915);
nor U9696 (N_9696,N_8487,N_8089);
and U9697 (N_9697,N_8737,N_8165);
nand U9698 (N_9698,N_8298,N_8632);
and U9699 (N_9699,N_8097,N_8673);
nand U9700 (N_9700,N_8026,N_8753);
or U9701 (N_9701,N_8549,N_8004);
and U9702 (N_9702,N_8121,N_8612);
nand U9703 (N_9703,N_8603,N_8527);
or U9704 (N_9704,N_8007,N_8092);
nor U9705 (N_9705,N_8462,N_8294);
or U9706 (N_9706,N_8194,N_8164);
nand U9707 (N_9707,N_8191,N_8482);
or U9708 (N_9708,N_8318,N_8870);
or U9709 (N_9709,N_8311,N_8559);
nand U9710 (N_9710,N_8823,N_8398);
and U9711 (N_9711,N_8745,N_8160);
nand U9712 (N_9712,N_8498,N_8545);
nor U9713 (N_9713,N_8627,N_8344);
or U9714 (N_9714,N_8266,N_8075);
or U9715 (N_9715,N_8739,N_8805);
or U9716 (N_9716,N_8464,N_8896);
nor U9717 (N_9717,N_8083,N_8879);
nor U9718 (N_9718,N_8751,N_8459);
xnor U9719 (N_9719,N_8580,N_8598);
and U9720 (N_9720,N_8376,N_8822);
and U9721 (N_9721,N_8484,N_8511);
or U9722 (N_9722,N_8659,N_8928);
and U9723 (N_9723,N_8007,N_8577);
nor U9724 (N_9724,N_8091,N_8879);
or U9725 (N_9725,N_8926,N_8570);
nor U9726 (N_9726,N_8897,N_8695);
nor U9727 (N_9727,N_8480,N_8360);
nor U9728 (N_9728,N_8098,N_8188);
or U9729 (N_9729,N_8483,N_8951);
and U9730 (N_9730,N_8283,N_8124);
or U9731 (N_9731,N_8836,N_8302);
nand U9732 (N_9732,N_8169,N_8785);
nor U9733 (N_9733,N_8074,N_8315);
nand U9734 (N_9734,N_8730,N_8226);
nor U9735 (N_9735,N_8228,N_8000);
or U9736 (N_9736,N_8594,N_8584);
and U9737 (N_9737,N_8408,N_8829);
nor U9738 (N_9738,N_8007,N_8792);
or U9739 (N_9739,N_8884,N_8043);
nand U9740 (N_9740,N_8665,N_8784);
and U9741 (N_9741,N_8399,N_8573);
xnor U9742 (N_9742,N_8870,N_8346);
nor U9743 (N_9743,N_8549,N_8883);
and U9744 (N_9744,N_8457,N_8449);
nand U9745 (N_9745,N_8211,N_8292);
or U9746 (N_9746,N_8719,N_8481);
and U9747 (N_9747,N_8740,N_8239);
nand U9748 (N_9748,N_8286,N_8771);
nor U9749 (N_9749,N_8320,N_8034);
or U9750 (N_9750,N_8823,N_8265);
and U9751 (N_9751,N_8547,N_8314);
or U9752 (N_9752,N_8191,N_8272);
nand U9753 (N_9753,N_8251,N_8186);
or U9754 (N_9754,N_8944,N_8275);
or U9755 (N_9755,N_8605,N_8622);
xnor U9756 (N_9756,N_8964,N_8723);
and U9757 (N_9757,N_8399,N_8075);
or U9758 (N_9758,N_8180,N_8647);
and U9759 (N_9759,N_8113,N_8027);
xor U9760 (N_9760,N_8881,N_8844);
nand U9761 (N_9761,N_8154,N_8591);
and U9762 (N_9762,N_8840,N_8852);
nor U9763 (N_9763,N_8318,N_8730);
or U9764 (N_9764,N_8046,N_8151);
xnor U9765 (N_9765,N_8705,N_8074);
or U9766 (N_9766,N_8322,N_8915);
nor U9767 (N_9767,N_8851,N_8069);
nand U9768 (N_9768,N_8294,N_8205);
and U9769 (N_9769,N_8169,N_8303);
xnor U9770 (N_9770,N_8473,N_8119);
nand U9771 (N_9771,N_8857,N_8142);
nand U9772 (N_9772,N_8411,N_8871);
or U9773 (N_9773,N_8374,N_8493);
nor U9774 (N_9774,N_8237,N_8242);
or U9775 (N_9775,N_8947,N_8423);
nor U9776 (N_9776,N_8720,N_8860);
and U9777 (N_9777,N_8796,N_8103);
or U9778 (N_9778,N_8817,N_8187);
xnor U9779 (N_9779,N_8240,N_8519);
nor U9780 (N_9780,N_8031,N_8298);
nor U9781 (N_9781,N_8691,N_8115);
nor U9782 (N_9782,N_8015,N_8443);
nand U9783 (N_9783,N_8117,N_8905);
nor U9784 (N_9784,N_8392,N_8829);
or U9785 (N_9785,N_8851,N_8831);
or U9786 (N_9786,N_8668,N_8418);
and U9787 (N_9787,N_8961,N_8416);
nand U9788 (N_9788,N_8109,N_8393);
nor U9789 (N_9789,N_8805,N_8163);
nand U9790 (N_9790,N_8645,N_8939);
nand U9791 (N_9791,N_8692,N_8779);
or U9792 (N_9792,N_8194,N_8221);
or U9793 (N_9793,N_8802,N_8119);
nor U9794 (N_9794,N_8876,N_8149);
or U9795 (N_9795,N_8928,N_8967);
xor U9796 (N_9796,N_8392,N_8389);
nand U9797 (N_9797,N_8296,N_8945);
and U9798 (N_9798,N_8817,N_8323);
or U9799 (N_9799,N_8386,N_8585);
and U9800 (N_9800,N_8004,N_8712);
nand U9801 (N_9801,N_8371,N_8276);
nand U9802 (N_9802,N_8886,N_8361);
or U9803 (N_9803,N_8652,N_8483);
or U9804 (N_9804,N_8083,N_8740);
nand U9805 (N_9805,N_8725,N_8597);
xnor U9806 (N_9806,N_8745,N_8378);
and U9807 (N_9807,N_8511,N_8161);
nor U9808 (N_9808,N_8826,N_8096);
nor U9809 (N_9809,N_8922,N_8586);
xnor U9810 (N_9810,N_8632,N_8129);
nor U9811 (N_9811,N_8213,N_8835);
xnor U9812 (N_9812,N_8729,N_8368);
or U9813 (N_9813,N_8812,N_8771);
nor U9814 (N_9814,N_8663,N_8949);
or U9815 (N_9815,N_8958,N_8641);
nand U9816 (N_9816,N_8178,N_8860);
or U9817 (N_9817,N_8389,N_8457);
or U9818 (N_9818,N_8087,N_8094);
xnor U9819 (N_9819,N_8326,N_8603);
xor U9820 (N_9820,N_8870,N_8008);
and U9821 (N_9821,N_8033,N_8514);
or U9822 (N_9822,N_8127,N_8776);
nand U9823 (N_9823,N_8132,N_8728);
and U9824 (N_9824,N_8874,N_8340);
or U9825 (N_9825,N_8173,N_8127);
nand U9826 (N_9826,N_8017,N_8385);
or U9827 (N_9827,N_8072,N_8178);
nand U9828 (N_9828,N_8191,N_8006);
and U9829 (N_9829,N_8579,N_8509);
and U9830 (N_9830,N_8371,N_8352);
or U9831 (N_9831,N_8197,N_8362);
or U9832 (N_9832,N_8320,N_8148);
or U9833 (N_9833,N_8358,N_8732);
or U9834 (N_9834,N_8368,N_8165);
nand U9835 (N_9835,N_8490,N_8248);
xor U9836 (N_9836,N_8318,N_8692);
xor U9837 (N_9837,N_8834,N_8500);
or U9838 (N_9838,N_8541,N_8634);
or U9839 (N_9839,N_8436,N_8305);
nor U9840 (N_9840,N_8023,N_8329);
or U9841 (N_9841,N_8989,N_8063);
and U9842 (N_9842,N_8987,N_8271);
nor U9843 (N_9843,N_8466,N_8799);
nand U9844 (N_9844,N_8114,N_8210);
and U9845 (N_9845,N_8672,N_8877);
nor U9846 (N_9846,N_8160,N_8364);
or U9847 (N_9847,N_8181,N_8982);
or U9848 (N_9848,N_8307,N_8412);
and U9849 (N_9849,N_8142,N_8606);
and U9850 (N_9850,N_8653,N_8699);
or U9851 (N_9851,N_8518,N_8325);
and U9852 (N_9852,N_8095,N_8974);
nor U9853 (N_9853,N_8378,N_8762);
or U9854 (N_9854,N_8573,N_8366);
nor U9855 (N_9855,N_8481,N_8578);
nand U9856 (N_9856,N_8381,N_8908);
xor U9857 (N_9857,N_8671,N_8318);
nor U9858 (N_9858,N_8091,N_8247);
and U9859 (N_9859,N_8990,N_8411);
nor U9860 (N_9860,N_8021,N_8264);
or U9861 (N_9861,N_8516,N_8093);
nor U9862 (N_9862,N_8371,N_8188);
nand U9863 (N_9863,N_8464,N_8721);
nor U9864 (N_9864,N_8232,N_8502);
nand U9865 (N_9865,N_8333,N_8081);
nand U9866 (N_9866,N_8358,N_8160);
nor U9867 (N_9867,N_8711,N_8950);
or U9868 (N_9868,N_8149,N_8223);
nor U9869 (N_9869,N_8506,N_8097);
and U9870 (N_9870,N_8051,N_8649);
xnor U9871 (N_9871,N_8012,N_8928);
or U9872 (N_9872,N_8787,N_8061);
and U9873 (N_9873,N_8149,N_8553);
nand U9874 (N_9874,N_8677,N_8619);
nor U9875 (N_9875,N_8234,N_8577);
or U9876 (N_9876,N_8744,N_8009);
nand U9877 (N_9877,N_8292,N_8532);
nor U9878 (N_9878,N_8210,N_8220);
or U9879 (N_9879,N_8951,N_8330);
xor U9880 (N_9880,N_8515,N_8121);
nand U9881 (N_9881,N_8048,N_8905);
and U9882 (N_9882,N_8442,N_8534);
and U9883 (N_9883,N_8664,N_8592);
xnor U9884 (N_9884,N_8891,N_8859);
or U9885 (N_9885,N_8582,N_8831);
and U9886 (N_9886,N_8715,N_8585);
nand U9887 (N_9887,N_8462,N_8929);
nor U9888 (N_9888,N_8618,N_8529);
nor U9889 (N_9889,N_8019,N_8209);
nor U9890 (N_9890,N_8481,N_8071);
xnor U9891 (N_9891,N_8554,N_8507);
nand U9892 (N_9892,N_8612,N_8704);
or U9893 (N_9893,N_8074,N_8924);
nor U9894 (N_9894,N_8855,N_8536);
and U9895 (N_9895,N_8829,N_8757);
or U9896 (N_9896,N_8348,N_8908);
or U9897 (N_9897,N_8994,N_8712);
and U9898 (N_9898,N_8449,N_8679);
nand U9899 (N_9899,N_8797,N_8586);
or U9900 (N_9900,N_8992,N_8114);
nand U9901 (N_9901,N_8022,N_8816);
or U9902 (N_9902,N_8534,N_8719);
or U9903 (N_9903,N_8395,N_8278);
or U9904 (N_9904,N_8496,N_8046);
nor U9905 (N_9905,N_8548,N_8397);
nor U9906 (N_9906,N_8184,N_8197);
nor U9907 (N_9907,N_8901,N_8828);
nor U9908 (N_9908,N_8037,N_8438);
and U9909 (N_9909,N_8019,N_8392);
nor U9910 (N_9910,N_8748,N_8528);
xnor U9911 (N_9911,N_8610,N_8845);
nor U9912 (N_9912,N_8156,N_8042);
xor U9913 (N_9913,N_8179,N_8092);
nor U9914 (N_9914,N_8378,N_8934);
and U9915 (N_9915,N_8300,N_8412);
xnor U9916 (N_9916,N_8611,N_8102);
nand U9917 (N_9917,N_8623,N_8629);
nand U9918 (N_9918,N_8900,N_8793);
or U9919 (N_9919,N_8836,N_8988);
and U9920 (N_9920,N_8999,N_8572);
or U9921 (N_9921,N_8600,N_8708);
and U9922 (N_9922,N_8705,N_8580);
nand U9923 (N_9923,N_8116,N_8069);
or U9924 (N_9924,N_8832,N_8534);
nand U9925 (N_9925,N_8829,N_8456);
and U9926 (N_9926,N_8068,N_8337);
and U9927 (N_9927,N_8416,N_8397);
nand U9928 (N_9928,N_8764,N_8676);
and U9929 (N_9929,N_8285,N_8812);
nand U9930 (N_9930,N_8498,N_8027);
or U9931 (N_9931,N_8424,N_8958);
xnor U9932 (N_9932,N_8603,N_8399);
and U9933 (N_9933,N_8047,N_8645);
and U9934 (N_9934,N_8248,N_8498);
or U9935 (N_9935,N_8885,N_8498);
and U9936 (N_9936,N_8424,N_8640);
nor U9937 (N_9937,N_8905,N_8697);
nor U9938 (N_9938,N_8061,N_8915);
or U9939 (N_9939,N_8161,N_8287);
or U9940 (N_9940,N_8427,N_8514);
and U9941 (N_9941,N_8110,N_8201);
nand U9942 (N_9942,N_8026,N_8244);
nor U9943 (N_9943,N_8869,N_8767);
or U9944 (N_9944,N_8380,N_8177);
and U9945 (N_9945,N_8939,N_8199);
or U9946 (N_9946,N_8457,N_8134);
and U9947 (N_9947,N_8463,N_8952);
xor U9948 (N_9948,N_8822,N_8682);
nor U9949 (N_9949,N_8718,N_8228);
and U9950 (N_9950,N_8791,N_8935);
xor U9951 (N_9951,N_8859,N_8712);
nor U9952 (N_9952,N_8161,N_8376);
or U9953 (N_9953,N_8311,N_8630);
nor U9954 (N_9954,N_8772,N_8301);
nand U9955 (N_9955,N_8524,N_8908);
and U9956 (N_9956,N_8254,N_8877);
nor U9957 (N_9957,N_8930,N_8671);
nand U9958 (N_9958,N_8678,N_8081);
and U9959 (N_9959,N_8041,N_8048);
nor U9960 (N_9960,N_8013,N_8642);
nand U9961 (N_9961,N_8407,N_8401);
or U9962 (N_9962,N_8385,N_8492);
and U9963 (N_9963,N_8059,N_8355);
and U9964 (N_9964,N_8550,N_8628);
nand U9965 (N_9965,N_8739,N_8779);
nor U9966 (N_9966,N_8013,N_8197);
nand U9967 (N_9967,N_8200,N_8165);
nor U9968 (N_9968,N_8513,N_8401);
xnor U9969 (N_9969,N_8825,N_8888);
nor U9970 (N_9970,N_8832,N_8264);
nor U9971 (N_9971,N_8516,N_8351);
nor U9972 (N_9972,N_8395,N_8676);
nor U9973 (N_9973,N_8768,N_8225);
nand U9974 (N_9974,N_8586,N_8188);
and U9975 (N_9975,N_8933,N_8009);
and U9976 (N_9976,N_8750,N_8835);
xnor U9977 (N_9977,N_8297,N_8587);
nand U9978 (N_9978,N_8555,N_8706);
or U9979 (N_9979,N_8649,N_8658);
nand U9980 (N_9980,N_8350,N_8507);
or U9981 (N_9981,N_8311,N_8536);
nor U9982 (N_9982,N_8812,N_8448);
or U9983 (N_9983,N_8147,N_8559);
and U9984 (N_9984,N_8001,N_8403);
or U9985 (N_9985,N_8155,N_8620);
or U9986 (N_9986,N_8281,N_8816);
nor U9987 (N_9987,N_8058,N_8766);
nand U9988 (N_9988,N_8939,N_8925);
and U9989 (N_9989,N_8838,N_8453);
and U9990 (N_9990,N_8642,N_8808);
nor U9991 (N_9991,N_8796,N_8453);
and U9992 (N_9992,N_8228,N_8930);
nor U9993 (N_9993,N_8298,N_8547);
or U9994 (N_9994,N_8293,N_8862);
nor U9995 (N_9995,N_8686,N_8803);
nand U9996 (N_9996,N_8356,N_8043);
xnor U9997 (N_9997,N_8273,N_8597);
nand U9998 (N_9998,N_8955,N_8046);
nor U9999 (N_9999,N_8955,N_8610);
nor U10000 (N_10000,N_9768,N_9569);
nand U10001 (N_10001,N_9349,N_9374);
nand U10002 (N_10002,N_9910,N_9684);
nand U10003 (N_10003,N_9459,N_9399);
nor U10004 (N_10004,N_9798,N_9361);
or U10005 (N_10005,N_9249,N_9025);
and U10006 (N_10006,N_9587,N_9849);
or U10007 (N_10007,N_9516,N_9393);
and U10008 (N_10008,N_9014,N_9287);
or U10009 (N_10009,N_9811,N_9278);
nand U10010 (N_10010,N_9661,N_9006);
and U10011 (N_10011,N_9963,N_9335);
nand U10012 (N_10012,N_9908,N_9188);
nand U10013 (N_10013,N_9513,N_9751);
xnor U10014 (N_10014,N_9038,N_9022);
xor U10015 (N_10015,N_9814,N_9450);
xor U10016 (N_10016,N_9184,N_9434);
nor U10017 (N_10017,N_9870,N_9427);
nor U10018 (N_10018,N_9899,N_9789);
nor U10019 (N_10019,N_9271,N_9639);
nand U10020 (N_10020,N_9795,N_9250);
nand U10021 (N_10021,N_9699,N_9955);
or U10022 (N_10022,N_9939,N_9246);
or U10023 (N_10023,N_9402,N_9075);
or U10024 (N_10024,N_9562,N_9536);
nand U10025 (N_10025,N_9218,N_9827);
or U10026 (N_10026,N_9260,N_9162);
nand U10027 (N_10027,N_9511,N_9183);
or U10028 (N_10028,N_9378,N_9883);
nand U10029 (N_10029,N_9767,N_9632);
and U10030 (N_10030,N_9835,N_9956);
nand U10031 (N_10031,N_9706,N_9128);
and U10032 (N_10032,N_9042,N_9410);
nand U10033 (N_10033,N_9600,N_9698);
nand U10034 (N_10034,N_9400,N_9294);
nand U10035 (N_10035,N_9051,N_9680);
and U10036 (N_10036,N_9417,N_9660);
and U10037 (N_10037,N_9640,N_9930);
or U10038 (N_10038,N_9238,N_9651);
xnor U10039 (N_10039,N_9046,N_9938);
nor U10040 (N_10040,N_9122,N_9888);
nor U10041 (N_10041,N_9013,N_9714);
or U10042 (N_10042,N_9103,N_9211);
and U10043 (N_10043,N_9097,N_9901);
nand U10044 (N_10044,N_9535,N_9317);
nor U10045 (N_10045,N_9653,N_9201);
nor U10046 (N_10046,N_9381,N_9059);
nor U10047 (N_10047,N_9072,N_9288);
or U10048 (N_10048,N_9048,N_9305);
or U10049 (N_10049,N_9725,N_9364);
or U10050 (N_10050,N_9894,N_9664);
or U10051 (N_10051,N_9416,N_9248);
nand U10052 (N_10052,N_9177,N_9957);
or U10053 (N_10053,N_9005,N_9225);
or U10054 (N_10054,N_9263,N_9323);
or U10055 (N_10055,N_9770,N_9848);
nand U10056 (N_10056,N_9360,N_9089);
and U10057 (N_10057,N_9439,N_9721);
xor U10058 (N_10058,N_9466,N_9406);
nor U10059 (N_10059,N_9228,N_9255);
and U10060 (N_10060,N_9669,N_9129);
or U10061 (N_10061,N_9800,N_9160);
xor U10062 (N_10062,N_9920,N_9605);
xor U10063 (N_10063,N_9233,N_9948);
or U10064 (N_10064,N_9921,N_9531);
nand U10065 (N_10065,N_9952,N_9745);
nor U10066 (N_10066,N_9585,N_9864);
or U10067 (N_10067,N_9504,N_9276);
or U10068 (N_10068,N_9766,N_9762);
or U10069 (N_10069,N_9510,N_9477);
nand U10070 (N_10070,N_9635,N_9886);
or U10071 (N_10071,N_9214,N_9623);
nor U10072 (N_10072,N_9873,N_9926);
nand U10073 (N_10073,N_9682,N_9186);
nand U10074 (N_10074,N_9016,N_9475);
or U10075 (N_10075,N_9134,N_9889);
or U10076 (N_10076,N_9710,N_9777);
nor U10077 (N_10077,N_9481,N_9769);
nand U10078 (N_10078,N_9702,N_9931);
nor U10079 (N_10079,N_9980,N_9350);
and U10080 (N_10080,N_9392,N_9776);
and U10081 (N_10081,N_9729,N_9482);
and U10082 (N_10082,N_9999,N_9990);
or U10083 (N_10083,N_9251,N_9805);
xor U10084 (N_10084,N_9234,N_9711);
nand U10085 (N_10085,N_9469,N_9825);
or U10086 (N_10086,N_9989,N_9689);
nand U10087 (N_10087,N_9471,N_9953);
xnor U10088 (N_10088,N_9296,N_9053);
or U10089 (N_10089,N_9227,N_9217);
xnor U10090 (N_10090,N_9633,N_9212);
or U10091 (N_10091,N_9914,N_9590);
or U10092 (N_10092,N_9572,N_9861);
nor U10093 (N_10093,N_9954,N_9951);
nor U10094 (N_10094,N_9026,N_9902);
xnor U10095 (N_10095,N_9101,N_9433);
nand U10096 (N_10096,N_9226,N_9525);
or U10097 (N_10097,N_9982,N_9192);
nand U10098 (N_10098,N_9891,N_9194);
xor U10099 (N_10099,N_9306,N_9817);
nand U10100 (N_10100,N_9937,N_9787);
nand U10101 (N_10101,N_9489,N_9332);
nor U10102 (N_10102,N_9541,N_9197);
or U10103 (N_10103,N_9913,N_9152);
or U10104 (N_10104,N_9505,N_9720);
and U10105 (N_10105,N_9297,N_9231);
nand U10106 (N_10106,N_9001,N_9803);
and U10107 (N_10107,N_9120,N_9259);
nor U10108 (N_10108,N_9688,N_9449);
nor U10109 (N_10109,N_9422,N_9851);
or U10110 (N_10110,N_9300,N_9380);
nand U10111 (N_10111,N_9693,N_9718);
nand U10112 (N_10112,N_9067,N_9498);
nor U10113 (N_10113,N_9991,N_9221);
and U10114 (N_10114,N_9039,N_9815);
xnor U10115 (N_10115,N_9918,N_9232);
nor U10116 (N_10116,N_9838,N_9836);
and U10117 (N_10117,N_9934,N_9379);
nor U10118 (N_10118,N_9696,N_9925);
and U10119 (N_10119,N_9539,N_9237);
or U10120 (N_10120,N_9662,N_9788);
or U10121 (N_10121,N_9842,N_9117);
or U10122 (N_10122,N_9448,N_9759);
or U10123 (N_10123,N_9834,N_9163);
and U10124 (N_10124,N_9880,N_9972);
or U10125 (N_10125,N_9791,N_9858);
nand U10126 (N_10126,N_9673,N_9521);
and U10127 (N_10127,N_9176,N_9890);
and U10128 (N_10128,N_9373,N_9049);
nand U10129 (N_10129,N_9312,N_9343);
and U10130 (N_10130,N_9494,N_9421);
xor U10131 (N_10131,N_9011,N_9998);
and U10132 (N_10132,N_9885,N_9372);
and U10133 (N_10133,N_9322,N_9385);
nand U10134 (N_10134,N_9619,N_9155);
or U10135 (N_10135,N_9601,N_9534);
nor U10136 (N_10136,N_9984,N_9734);
and U10137 (N_10137,N_9874,N_9205);
nor U10138 (N_10138,N_9922,N_9801);
and U10139 (N_10139,N_9345,N_9266);
nor U10140 (N_10140,N_9784,N_9333);
or U10141 (N_10141,N_9658,N_9057);
or U10142 (N_10142,N_9359,N_9451);
nand U10143 (N_10143,N_9193,N_9239);
or U10144 (N_10144,N_9964,N_9293);
or U10145 (N_10145,N_9644,N_9470);
nor U10146 (N_10146,N_9149,N_9522);
nor U10147 (N_10147,N_9070,N_9054);
nor U10148 (N_10148,N_9463,N_9114);
xnor U10149 (N_10149,N_9301,N_9987);
and U10150 (N_10150,N_9445,N_9617);
and U10151 (N_10151,N_9657,N_9544);
nand U10152 (N_10152,N_9747,N_9310);
and U10153 (N_10153,N_9659,N_9992);
nor U10154 (N_10154,N_9283,N_9377);
or U10155 (N_10155,N_9295,N_9198);
or U10156 (N_10156,N_9116,N_9465);
nor U10157 (N_10157,N_9764,N_9010);
nand U10158 (N_10158,N_9137,N_9037);
nand U10159 (N_10159,N_9031,N_9665);
xor U10160 (N_10160,N_9023,N_9969);
nand U10161 (N_10161,N_9329,N_9435);
or U10162 (N_10162,N_9358,N_9429);
nor U10163 (N_10163,N_9738,N_9040);
nand U10164 (N_10164,N_9876,N_9898);
nor U10165 (N_10165,N_9147,N_9576);
or U10166 (N_10166,N_9102,N_9012);
nand U10167 (N_10167,N_9589,N_9737);
and U10168 (N_10168,N_9882,N_9388);
or U10169 (N_10169,N_9119,N_9638);
nand U10170 (N_10170,N_9456,N_9960);
or U10171 (N_10171,N_9196,N_9367);
nand U10172 (N_10172,N_9857,N_9806);
nor U10173 (N_10173,N_9540,N_9809);
and U10174 (N_10174,N_9052,N_9760);
and U10175 (N_10175,N_9356,N_9065);
and U10176 (N_10176,N_9674,N_9277);
xnor U10177 (N_10177,N_9597,N_9109);
and U10178 (N_10178,N_9733,N_9782);
or U10179 (N_10179,N_9642,N_9017);
or U10180 (N_10180,N_9376,N_9141);
nor U10181 (N_10181,N_9761,N_9631);
nand U10182 (N_10182,N_9823,N_9919);
nor U10183 (N_10183,N_9143,N_9321);
and U10184 (N_10184,N_9113,N_9190);
and U10185 (N_10185,N_9003,N_9424);
nor U10186 (N_10186,N_9941,N_9743);
and U10187 (N_10187,N_9961,N_9903);
and U10188 (N_10188,N_9598,N_9905);
and U10189 (N_10189,N_9503,N_9911);
or U10190 (N_10190,N_9484,N_9032);
nor U10191 (N_10191,N_9896,N_9303);
or U10192 (N_10192,N_9512,N_9215);
nand U10193 (N_10193,N_9187,N_9492);
xnor U10194 (N_10194,N_9588,N_9528);
nor U10195 (N_10195,N_9181,N_9455);
xor U10196 (N_10196,N_9839,N_9092);
nand U10197 (N_10197,N_9501,N_9348);
nor U10198 (N_10198,N_9140,N_9900);
or U10199 (N_10199,N_9443,N_9326);
or U10200 (N_10200,N_9897,N_9123);
or U10201 (N_10201,N_9386,N_9676);
xnor U10202 (N_10202,N_9959,N_9907);
and U10203 (N_10203,N_9495,N_9508);
or U10204 (N_10204,N_9428,N_9004);
nand U10205 (N_10205,N_9558,N_9357);
or U10206 (N_10206,N_9912,N_9744);
or U10207 (N_10207,N_9229,N_9968);
nor U10208 (N_10208,N_9172,N_9906);
and U10209 (N_10209,N_9663,N_9950);
xnor U10210 (N_10210,N_9563,N_9547);
nor U10211 (N_10211,N_9780,N_9174);
xor U10212 (N_10212,N_9274,N_9337);
nor U10213 (N_10213,N_9866,N_9586);
and U10214 (N_10214,N_9420,N_9182);
or U10215 (N_10215,N_9750,N_9395);
and U10216 (N_10216,N_9088,N_9518);
nand U10217 (N_10217,N_9064,N_9491);
nand U10218 (N_10218,N_9254,N_9979);
nor U10219 (N_10219,N_9893,N_9872);
nand U10220 (N_10220,N_9869,N_9749);
and U10221 (N_10221,N_9695,N_9189);
nand U10222 (N_10222,N_9146,N_9523);
xnor U10223 (N_10223,N_9892,N_9154);
nand U10224 (N_10224,N_9216,N_9009);
xnor U10225 (N_10225,N_9486,N_9625);
xnor U10226 (N_10226,N_9976,N_9408);
or U10227 (N_10227,N_9325,N_9502);
nand U10228 (N_10228,N_9490,N_9790);
or U10229 (N_10229,N_9773,N_9881);
xnor U10230 (N_10230,N_9204,N_9082);
nand U10231 (N_10231,N_9180,N_9785);
and U10232 (N_10232,N_9175,N_9258);
nand U10233 (N_10233,N_9629,N_9008);
and U10234 (N_10234,N_9062,N_9077);
xnor U10235 (N_10235,N_9079,N_9375);
xnor U10236 (N_10236,N_9136,N_9257);
nand U10237 (N_10237,N_9222,N_9041);
nor U10238 (N_10238,N_9654,N_9515);
and U10239 (N_10239,N_9855,N_9068);
nor U10240 (N_10240,N_9656,N_9715);
and U10241 (N_10241,N_9850,N_9599);
or U10242 (N_10242,N_9530,N_9178);
nand U10243 (N_10243,N_9262,N_9087);
and U10244 (N_10244,N_9833,N_9647);
nor U10245 (N_10245,N_9407,N_9253);
and U10246 (N_10246,N_9369,N_9207);
nand U10247 (N_10247,N_9320,N_9159);
and U10248 (N_10248,N_9454,N_9363);
nor U10249 (N_10249,N_9135,N_9703);
nand U10250 (N_10250,N_9436,N_9098);
or U10251 (N_10251,N_9115,N_9002);
xnor U10252 (N_10252,N_9624,N_9138);
nor U10253 (N_10253,N_9820,N_9324);
nand U10254 (N_10254,N_9813,N_9020);
or U10255 (N_10255,N_9928,N_9110);
nand U10256 (N_10256,N_9550,N_9552);
and U10257 (N_10257,N_9243,N_9804);
xnor U10258 (N_10258,N_9816,N_9945);
xor U10259 (N_10259,N_9575,N_9126);
nor U10260 (N_10260,N_9637,N_9018);
or U10261 (N_10261,N_9583,N_9168);
nor U10262 (N_10262,N_9462,N_9464);
nand U10263 (N_10263,N_9500,N_9650);
or U10264 (N_10264,N_9083,N_9728);
nand U10265 (N_10265,N_9628,N_9104);
or U10266 (N_10266,N_9467,N_9602);
or U10267 (N_10267,N_9045,N_9863);
or U10268 (N_10268,N_9697,N_9112);
or U10269 (N_10269,N_9548,N_9778);
and U10270 (N_10270,N_9423,N_9797);
and U10271 (N_10271,N_9279,N_9167);
xnor U10272 (N_10272,N_9822,N_9405);
nor U10273 (N_10273,N_9557,N_9050);
nor U10274 (N_10274,N_9591,N_9856);
or U10275 (N_10275,N_9812,N_9754);
or U10276 (N_10276,N_9304,N_9268);
nand U10277 (N_10277,N_9574,N_9206);
nor U10278 (N_10278,N_9442,N_9944);
and U10279 (N_10279,N_9578,N_9997);
or U10280 (N_10280,N_9107,N_9735);
and U10281 (N_10281,N_9105,N_9289);
nand U10282 (N_10282,N_9610,N_9156);
and U10283 (N_10283,N_9568,N_9242);
or U10284 (N_10284,N_9819,N_9485);
or U10285 (N_10285,N_9165,N_9592);
or U10286 (N_10286,N_9208,N_9347);
nand U10287 (N_10287,N_9125,N_9063);
nor U10288 (N_10288,N_9543,N_9593);
nor U10289 (N_10289,N_9694,N_9265);
nand U10290 (N_10290,N_9840,N_9401);
and U10291 (N_10291,N_9626,N_9044);
nor U10292 (N_10292,N_9185,N_9291);
xor U10293 (N_10293,N_9086,N_9331);
nand U10294 (N_10294,N_9108,N_9438);
xnor U10295 (N_10295,N_9847,N_9556);
xor U10296 (N_10296,N_9245,N_9841);
and U10297 (N_10297,N_9425,N_9313);
nand U10298 (N_10298,N_9244,N_9994);
nor U10299 (N_10299,N_9757,N_9796);
nand U10300 (N_10300,N_9564,N_9074);
xor U10301 (N_10301,N_9821,N_9546);
and U10302 (N_10302,N_9270,N_9191);
and U10303 (N_10303,N_9690,N_9679);
nor U10304 (N_10304,N_9646,N_9121);
nor U10305 (N_10305,N_9717,N_9775);
and U10306 (N_10306,N_9076,N_9582);
nor U10307 (N_10307,N_9877,N_9567);
and U10308 (N_10308,N_9832,N_9852);
xnor U10309 (N_10309,N_9043,N_9584);
nor U10310 (N_10310,N_9634,N_9479);
or U10311 (N_10311,N_9387,N_9727);
nor U10312 (N_10312,N_9978,N_9752);
or U10313 (N_10313,N_9554,N_9342);
nand U10314 (N_10314,N_9826,N_9620);
or U10315 (N_10315,N_9837,N_9034);
xnor U10316 (N_10316,N_9645,N_9452);
nand U10317 (N_10317,N_9173,N_9327);
nor U10318 (N_10318,N_9247,N_9929);
and U10319 (N_10319,N_9404,N_9415);
and U10320 (N_10320,N_9517,N_9281);
nor U10321 (N_10321,N_9096,N_9370);
nor U10322 (N_10322,N_9731,N_9958);
or U10323 (N_10323,N_9028,N_9383);
nor U10324 (N_10324,N_9616,N_9319);
and U10325 (N_10325,N_9476,N_9709);
or U10326 (N_10326,N_9437,N_9648);
and U10327 (N_10327,N_9845,N_9480);
nor U10328 (N_10328,N_9966,N_9118);
and U10329 (N_10329,N_9615,N_9085);
nand U10330 (N_10330,N_9412,N_9532);
and U10331 (N_10331,N_9933,N_9506);
nand U10332 (N_10332,N_9444,N_9403);
and U10333 (N_10333,N_9807,N_9298);
nor U10334 (N_10334,N_9862,N_9150);
and U10335 (N_10335,N_9542,N_9252);
or U10336 (N_10336,N_9967,N_9603);
nand U10337 (N_10337,N_9351,N_9195);
nand U10338 (N_10338,N_9655,N_9431);
and U10339 (N_10339,N_9707,N_9701);
xnor U10340 (N_10340,N_9675,N_9672);
or U10341 (N_10341,N_9742,N_9519);
xnor U10342 (N_10342,N_9030,N_9171);
nor U10343 (N_10343,N_9621,N_9884);
or U10344 (N_10344,N_9533,N_9529);
or U10345 (N_10345,N_9947,N_9566);
xnor U10346 (N_10346,N_9949,N_9818);
nor U10347 (N_10347,N_9241,N_9055);
and U10348 (N_10348,N_9256,N_9396);
nand U10349 (N_10349,N_9895,N_9802);
and U10350 (N_10350,N_9553,N_9507);
nor U10351 (N_10351,N_9447,N_9981);
and U10352 (N_10352,N_9091,N_9771);
and U10353 (N_10353,N_9686,N_9594);
and U10354 (N_10354,N_9740,N_9514);
nor U10355 (N_10355,N_9318,N_9681);
and U10356 (N_10356,N_9124,N_9432);
nand U10357 (N_10357,N_9200,N_9723);
nor U10358 (N_10358,N_9577,N_9334);
nand U10359 (N_10359,N_9153,N_9878);
or U10360 (N_10360,N_9166,N_9843);
nand U10361 (N_10361,N_9923,N_9753);
or U10362 (N_10362,N_9170,N_9524);
nor U10363 (N_10363,N_9794,N_9223);
xnor U10364 (N_10364,N_9867,N_9346);
and U10365 (N_10365,N_9169,N_9179);
nand U10366 (N_10366,N_9604,N_9722);
or U10367 (N_10367,N_9366,N_9144);
nor U10368 (N_10368,N_9986,N_9461);
xnor U10369 (N_10369,N_9061,N_9398);
nor U10370 (N_10370,N_9988,N_9829);
nor U10371 (N_10371,N_9844,N_9545);
nor U10372 (N_10372,N_9139,N_9158);
xor U10373 (N_10373,N_9607,N_9779);
nor U10374 (N_10374,N_9286,N_9499);
and U10375 (N_10375,N_9133,N_9235);
and U10376 (N_10376,N_9924,N_9995);
nand U10377 (N_10377,N_9157,N_9993);
and U10378 (N_10378,N_9704,N_9354);
nor U10379 (N_10379,N_9571,N_9219);
or U10380 (N_10380,N_9419,N_9854);
nor U10381 (N_10381,N_9774,N_9783);
or U10382 (N_10382,N_9965,N_9127);
nand U10383 (N_10383,N_9970,N_9142);
nand U10384 (N_10384,N_9641,N_9460);
nor U10385 (N_10385,N_9763,N_9330);
or U10386 (N_10386,N_9394,N_9338);
nor U10387 (N_10387,N_9210,N_9468);
nor U10388 (N_10388,N_9830,N_9643);
and U10389 (N_10389,N_9875,N_9935);
nor U10390 (N_10390,N_9786,N_9060);
or U10391 (N_10391,N_9758,N_9942);
and U10392 (N_10392,N_9493,N_9909);
or U10393 (N_10393,N_9446,N_9478);
nand U10394 (N_10394,N_9781,N_9936);
or U10395 (N_10395,N_9799,N_9340);
xor U10396 (N_10396,N_9538,N_9203);
and U10397 (N_10397,N_9756,N_9078);
xor U10398 (N_10398,N_9971,N_9904);
nand U10399 (N_10399,N_9716,N_9549);
nand U10400 (N_10400,N_9609,N_9015);
nor U10401 (N_10401,N_9362,N_9299);
or U10402 (N_10402,N_9453,N_9151);
or U10403 (N_10403,N_9474,N_9622);
nand U10404 (N_10404,N_9457,N_9496);
and U10405 (N_10405,N_9831,N_9736);
nand U10406 (N_10406,N_9035,N_9560);
nor U10407 (N_10407,N_9213,N_9099);
or U10408 (N_10408,N_9916,N_9000);
or U10409 (N_10409,N_9666,N_9871);
nand U10410 (N_10410,N_9090,N_9100);
nand U10411 (N_10411,N_9084,N_9161);
nand U10412 (N_10412,N_9527,N_9440);
and U10413 (N_10413,N_9328,N_9284);
or U10414 (N_10414,N_9677,N_9290);
nor U10415 (N_10415,N_9962,N_9081);
nor U10416 (N_10416,N_9414,N_9036);
or U10417 (N_10417,N_9683,N_9371);
nor U10418 (N_10418,N_9473,N_9095);
nand U10419 (N_10419,N_9353,N_9810);
nand U10420 (N_10420,N_9868,N_9224);
and U10421 (N_10421,N_9355,N_9093);
nor U10422 (N_10422,N_9730,N_9687);
nor U10423 (N_10423,N_9390,N_9382);
nand U10424 (N_10424,N_9860,N_9595);
nor U10425 (N_10425,N_9391,N_9033);
and U10426 (N_10426,N_9739,N_9397);
and U10427 (N_10427,N_9282,N_9565);
or U10428 (N_10428,N_9946,N_9573);
and U10429 (N_10429,N_9199,N_9652);
nor U10430 (N_10430,N_9824,N_9741);
and U10431 (N_10431,N_9581,N_9220);
or U10432 (N_10432,N_9853,N_9019);
nand U10433 (N_10433,N_9069,N_9384);
and U10434 (N_10434,N_9649,N_9365);
and U10435 (N_10435,N_9808,N_9940);
nand U10436 (N_10436,N_9765,N_9755);
nand U10437 (N_10437,N_9846,N_9272);
or U10438 (N_10438,N_9418,N_9915);
nor U10439 (N_10439,N_9047,N_9859);
nor U10440 (N_10440,N_9708,N_9555);
nand U10441 (N_10441,N_9671,N_9561);
nor U10442 (N_10442,N_9685,N_9024);
and U10443 (N_10443,N_9292,N_9341);
and U10444 (N_10444,N_9732,N_9887);
and U10445 (N_10445,N_9596,N_9021);
nor U10446 (N_10446,N_9667,N_9977);
nand U10447 (N_10447,N_9712,N_9700);
nor U10448 (N_10448,N_9267,N_9027);
and U10449 (N_10449,N_9975,N_9273);
nand U10450 (N_10450,N_9389,N_9236);
or U10451 (N_10451,N_9106,N_9148);
and U10452 (N_10452,N_9748,N_9409);
nand U10453 (N_10453,N_9309,N_9285);
and U10454 (N_10454,N_9497,N_9996);
or U10455 (N_10455,N_9264,N_9488);
nor U10456 (N_10456,N_9275,N_9007);
and U10457 (N_10457,N_9613,N_9202);
nor U10458 (N_10458,N_9307,N_9441);
or U10459 (N_10459,N_9792,N_9094);
xnor U10460 (N_10460,N_9131,N_9071);
or U10461 (N_10461,N_9308,N_9080);
and U10462 (N_10462,N_9280,N_9472);
or U10463 (N_10463,N_9368,N_9828);
nor U10464 (N_10464,N_9526,N_9551);
nor U10465 (N_10465,N_9691,N_9487);
and U10466 (N_10466,N_9627,N_9705);
or U10467 (N_10467,N_9943,N_9692);
and U10468 (N_10468,N_9746,N_9058);
nand U10469 (N_10469,N_9719,N_9426);
and U10470 (N_10470,N_9772,N_9559);
and U10471 (N_10471,N_9269,N_9974);
nor U10472 (N_10472,N_9314,N_9614);
nor U10473 (N_10473,N_9336,N_9678);
and U10474 (N_10474,N_9606,N_9520);
and U10475 (N_10475,N_9579,N_9932);
and U10476 (N_10476,N_9580,N_9130);
nor U10477 (N_10477,N_9927,N_9413);
and U10478 (N_10478,N_9066,N_9315);
nor U10479 (N_10479,N_9316,N_9793);
or U10480 (N_10480,N_9111,N_9164);
and U10481 (N_10481,N_9618,N_9458);
nand U10482 (N_10482,N_9973,N_9029);
nor U10483 (N_10483,N_9339,N_9509);
or U10484 (N_10484,N_9917,N_9240);
and U10485 (N_10485,N_9611,N_9570);
nand U10486 (N_10486,N_9145,N_9983);
or U10487 (N_10487,N_9411,N_9430);
and U10488 (N_10488,N_9724,N_9879);
or U10489 (N_10489,N_9302,N_9630);
nor U10490 (N_10490,N_9209,N_9668);
nand U10491 (N_10491,N_9352,N_9132);
xor U10492 (N_10492,N_9056,N_9483);
xnor U10493 (N_10493,N_9311,N_9612);
xnor U10494 (N_10494,N_9670,N_9726);
nand U10495 (N_10495,N_9230,N_9865);
nor U10496 (N_10496,N_9537,N_9636);
nor U10497 (N_10497,N_9261,N_9608);
or U10498 (N_10498,N_9985,N_9344);
nor U10499 (N_10499,N_9713,N_9073);
and U10500 (N_10500,N_9155,N_9021);
nor U10501 (N_10501,N_9845,N_9293);
and U10502 (N_10502,N_9053,N_9580);
xor U10503 (N_10503,N_9939,N_9182);
nor U10504 (N_10504,N_9420,N_9657);
or U10505 (N_10505,N_9701,N_9879);
nand U10506 (N_10506,N_9512,N_9071);
nor U10507 (N_10507,N_9108,N_9676);
nand U10508 (N_10508,N_9524,N_9603);
or U10509 (N_10509,N_9944,N_9758);
and U10510 (N_10510,N_9788,N_9014);
nor U10511 (N_10511,N_9302,N_9006);
nand U10512 (N_10512,N_9954,N_9598);
and U10513 (N_10513,N_9788,N_9624);
xnor U10514 (N_10514,N_9399,N_9927);
nand U10515 (N_10515,N_9427,N_9569);
and U10516 (N_10516,N_9938,N_9055);
nor U10517 (N_10517,N_9995,N_9192);
or U10518 (N_10518,N_9872,N_9823);
or U10519 (N_10519,N_9320,N_9076);
or U10520 (N_10520,N_9441,N_9242);
or U10521 (N_10521,N_9063,N_9647);
nor U10522 (N_10522,N_9090,N_9647);
and U10523 (N_10523,N_9080,N_9610);
and U10524 (N_10524,N_9839,N_9099);
or U10525 (N_10525,N_9751,N_9448);
or U10526 (N_10526,N_9588,N_9415);
or U10527 (N_10527,N_9046,N_9435);
or U10528 (N_10528,N_9261,N_9169);
and U10529 (N_10529,N_9832,N_9723);
nand U10530 (N_10530,N_9885,N_9473);
nand U10531 (N_10531,N_9926,N_9378);
nor U10532 (N_10532,N_9148,N_9395);
or U10533 (N_10533,N_9771,N_9588);
or U10534 (N_10534,N_9166,N_9380);
nor U10535 (N_10535,N_9597,N_9287);
and U10536 (N_10536,N_9366,N_9829);
or U10537 (N_10537,N_9832,N_9167);
or U10538 (N_10538,N_9738,N_9027);
and U10539 (N_10539,N_9272,N_9730);
or U10540 (N_10540,N_9074,N_9433);
nand U10541 (N_10541,N_9603,N_9704);
or U10542 (N_10542,N_9955,N_9472);
nor U10543 (N_10543,N_9571,N_9656);
or U10544 (N_10544,N_9520,N_9236);
nand U10545 (N_10545,N_9567,N_9113);
or U10546 (N_10546,N_9799,N_9814);
nor U10547 (N_10547,N_9610,N_9257);
or U10548 (N_10548,N_9034,N_9751);
xnor U10549 (N_10549,N_9683,N_9481);
or U10550 (N_10550,N_9138,N_9370);
and U10551 (N_10551,N_9872,N_9119);
xor U10552 (N_10552,N_9068,N_9908);
nor U10553 (N_10553,N_9086,N_9931);
xnor U10554 (N_10554,N_9174,N_9853);
or U10555 (N_10555,N_9855,N_9960);
or U10556 (N_10556,N_9263,N_9747);
nand U10557 (N_10557,N_9919,N_9770);
or U10558 (N_10558,N_9221,N_9767);
nor U10559 (N_10559,N_9782,N_9371);
or U10560 (N_10560,N_9368,N_9816);
and U10561 (N_10561,N_9016,N_9498);
nand U10562 (N_10562,N_9324,N_9183);
or U10563 (N_10563,N_9974,N_9426);
nand U10564 (N_10564,N_9405,N_9101);
or U10565 (N_10565,N_9932,N_9477);
nor U10566 (N_10566,N_9381,N_9840);
nor U10567 (N_10567,N_9201,N_9899);
nand U10568 (N_10568,N_9174,N_9257);
or U10569 (N_10569,N_9540,N_9390);
nand U10570 (N_10570,N_9496,N_9077);
and U10571 (N_10571,N_9164,N_9432);
and U10572 (N_10572,N_9499,N_9285);
nor U10573 (N_10573,N_9707,N_9716);
nand U10574 (N_10574,N_9513,N_9252);
and U10575 (N_10575,N_9881,N_9630);
and U10576 (N_10576,N_9961,N_9591);
and U10577 (N_10577,N_9267,N_9568);
or U10578 (N_10578,N_9316,N_9057);
and U10579 (N_10579,N_9343,N_9912);
and U10580 (N_10580,N_9655,N_9929);
or U10581 (N_10581,N_9420,N_9786);
xnor U10582 (N_10582,N_9517,N_9924);
and U10583 (N_10583,N_9627,N_9467);
nand U10584 (N_10584,N_9574,N_9607);
nor U10585 (N_10585,N_9578,N_9941);
nand U10586 (N_10586,N_9202,N_9281);
and U10587 (N_10587,N_9095,N_9584);
nand U10588 (N_10588,N_9910,N_9822);
xnor U10589 (N_10589,N_9882,N_9232);
nor U10590 (N_10590,N_9999,N_9121);
or U10591 (N_10591,N_9483,N_9511);
or U10592 (N_10592,N_9755,N_9244);
nand U10593 (N_10593,N_9288,N_9086);
and U10594 (N_10594,N_9746,N_9181);
and U10595 (N_10595,N_9568,N_9663);
nand U10596 (N_10596,N_9676,N_9745);
or U10597 (N_10597,N_9087,N_9056);
or U10598 (N_10598,N_9749,N_9690);
or U10599 (N_10599,N_9674,N_9011);
or U10600 (N_10600,N_9486,N_9130);
or U10601 (N_10601,N_9614,N_9534);
and U10602 (N_10602,N_9180,N_9870);
nand U10603 (N_10603,N_9260,N_9636);
or U10604 (N_10604,N_9230,N_9382);
nor U10605 (N_10605,N_9579,N_9582);
nor U10606 (N_10606,N_9265,N_9810);
and U10607 (N_10607,N_9764,N_9951);
xor U10608 (N_10608,N_9421,N_9353);
nand U10609 (N_10609,N_9812,N_9331);
xor U10610 (N_10610,N_9397,N_9446);
or U10611 (N_10611,N_9479,N_9394);
and U10612 (N_10612,N_9421,N_9680);
and U10613 (N_10613,N_9461,N_9590);
nand U10614 (N_10614,N_9379,N_9595);
nor U10615 (N_10615,N_9762,N_9325);
nand U10616 (N_10616,N_9366,N_9188);
or U10617 (N_10617,N_9073,N_9376);
nand U10618 (N_10618,N_9064,N_9530);
nor U10619 (N_10619,N_9480,N_9610);
and U10620 (N_10620,N_9122,N_9350);
or U10621 (N_10621,N_9609,N_9896);
and U10622 (N_10622,N_9779,N_9200);
and U10623 (N_10623,N_9369,N_9458);
nand U10624 (N_10624,N_9742,N_9787);
nand U10625 (N_10625,N_9784,N_9788);
nor U10626 (N_10626,N_9399,N_9890);
nor U10627 (N_10627,N_9124,N_9507);
nand U10628 (N_10628,N_9777,N_9594);
nand U10629 (N_10629,N_9062,N_9777);
nand U10630 (N_10630,N_9051,N_9049);
and U10631 (N_10631,N_9666,N_9244);
nand U10632 (N_10632,N_9482,N_9081);
nand U10633 (N_10633,N_9310,N_9389);
and U10634 (N_10634,N_9252,N_9588);
nor U10635 (N_10635,N_9640,N_9016);
nor U10636 (N_10636,N_9678,N_9364);
nor U10637 (N_10637,N_9738,N_9056);
nand U10638 (N_10638,N_9903,N_9294);
or U10639 (N_10639,N_9334,N_9792);
and U10640 (N_10640,N_9347,N_9325);
and U10641 (N_10641,N_9174,N_9497);
nand U10642 (N_10642,N_9181,N_9772);
nor U10643 (N_10643,N_9638,N_9134);
or U10644 (N_10644,N_9285,N_9526);
nor U10645 (N_10645,N_9564,N_9951);
and U10646 (N_10646,N_9205,N_9158);
nor U10647 (N_10647,N_9171,N_9367);
nor U10648 (N_10648,N_9701,N_9111);
or U10649 (N_10649,N_9839,N_9408);
and U10650 (N_10650,N_9402,N_9508);
and U10651 (N_10651,N_9366,N_9832);
and U10652 (N_10652,N_9301,N_9629);
nand U10653 (N_10653,N_9580,N_9924);
xnor U10654 (N_10654,N_9001,N_9343);
and U10655 (N_10655,N_9600,N_9423);
nor U10656 (N_10656,N_9012,N_9058);
or U10657 (N_10657,N_9077,N_9575);
xnor U10658 (N_10658,N_9065,N_9037);
or U10659 (N_10659,N_9161,N_9345);
or U10660 (N_10660,N_9977,N_9785);
xnor U10661 (N_10661,N_9545,N_9761);
nor U10662 (N_10662,N_9713,N_9413);
nor U10663 (N_10663,N_9645,N_9810);
and U10664 (N_10664,N_9995,N_9583);
nand U10665 (N_10665,N_9955,N_9183);
nor U10666 (N_10666,N_9115,N_9758);
or U10667 (N_10667,N_9175,N_9934);
or U10668 (N_10668,N_9090,N_9635);
and U10669 (N_10669,N_9305,N_9721);
or U10670 (N_10670,N_9939,N_9282);
nand U10671 (N_10671,N_9393,N_9912);
nand U10672 (N_10672,N_9186,N_9711);
and U10673 (N_10673,N_9269,N_9370);
xnor U10674 (N_10674,N_9522,N_9258);
nor U10675 (N_10675,N_9418,N_9037);
nand U10676 (N_10676,N_9880,N_9175);
and U10677 (N_10677,N_9294,N_9303);
or U10678 (N_10678,N_9832,N_9433);
or U10679 (N_10679,N_9829,N_9811);
xnor U10680 (N_10680,N_9163,N_9972);
or U10681 (N_10681,N_9007,N_9515);
and U10682 (N_10682,N_9013,N_9052);
nand U10683 (N_10683,N_9741,N_9315);
nand U10684 (N_10684,N_9318,N_9089);
and U10685 (N_10685,N_9572,N_9777);
nor U10686 (N_10686,N_9429,N_9783);
nor U10687 (N_10687,N_9727,N_9235);
nand U10688 (N_10688,N_9921,N_9501);
nor U10689 (N_10689,N_9058,N_9510);
or U10690 (N_10690,N_9047,N_9553);
nor U10691 (N_10691,N_9496,N_9552);
and U10692 (N_10692,N_9519,N_9880);
nor U10693 (N_10693,N_9852,N_9680);
nor U10694 (N_10694,N_9063,N_9892);
and U10695 (N_10695,N_9787,N_9680);
nand U10696 (N_10696,N_9383,N_9187);
nor U10697 (N_10697,N_9861,N_9302);
xnor U10698 (N_10698,N_9368,N_9641);
nand U10699 (N_10699,N_9943,N_9870);
and U10700 (N_10700,N_9103,N_9957);
and U10701 (N_10701,N_9795,N_9482);
or U10702 (N_10702,N_9577,N_9774);
and U10703 (N_10703,N_9615,N_9832);
nand U10704 (N_10704,N_9315,N_9421);
nor U10705 (N_10705,N_9454,N_9074);
xnor U10706 (N_10706,N_9130,N_9302);
nor U10707 (N_10707,N_9825,N_9402);
or U10708 (N_10708,N_9531,N_9086);
or U10709 (N_10709,N_9909,N_9132);
nor U10710 (N_10710,N_9299,N_9847);
nand U10711 (N_10711,N_9050,N_9273);
or U10712 (N_10712,N_9115,N_9653);
nand U10713 (N_10713,N_9919,N_9325);
or U10714 (N_10714,N_9758,N_9975);
or U10715 (N_10715,N_9591,N_9324);
or U10716 (N_10716,N_9378,N_9814);
xor U10717 (N_10717,N_9833,N_9807);
nand U10718 (N_10718,N_9351,N_9210);
nor U10719 (N_10719,N_9392,N_9224);
nor U10720 (N_10720,N_9180,N_9264);
xnor U10721 (N_10721,N_9813,N_9918);
or U10722 (N_10722,N_9701,N_9078);
xnor U10723 (N_10723,N_9337,N_9600);
nor U10724 (N_10724,N_9376,N_9397);
or U10725 (N_10725,N_9661,N_9759);
and U10726 (N_10726,N_9348,N_9531);
and U10727 (N_10727,N_9203,N_9602);
nor U10728 (N_10728,N_9828,N_9513);
or U10729 (N_10729,N_9697,N_9374);
or U10730 (N_10730,N_9195,N_9743);
and U10731 (N_10731,N_9820,N_9811);
nor U10732 (N_10732,N_9574,N_9373);
nand U10733 (N_10733,N_9119,N_9859);
nor U10734 (N_10734,N_9200,N_9176);
and U10735 (N_10735,N_9853,N_9210);
xnor U10736 (N_10736,N_9125,N_9620);
nor U10737 (N_10737,N_9100,N_9485);
and U10738 (N_10738,N_9584,N_9027);
or U10739 (N_10739,N_9877,N_9057);
nor U10740 (N_10740,N_9029,N_9099);
and U10741 (N_10741,N_9588,N_9739);
nor U10742 (N_10742,N_9335,N_9083);
xor U10743 (N_10743,N_9127,N_9288);
nand U10744 (N_10744,N_9785,N_9333);
or U10745 (N_10745,N_9973,N_9505);
and U10746 (N_10746,N_9248,N_9957);
and U10747 (N_10747,N_9141,N_9954);
nand U10748 (N_10748,N_9393,N_9637);
and U10749 (N_10749,N_9337,N_9014);
and U10750 (N_10750,N_9813,N_9064);
nor U10751 (N_10751,N_9249,N_9704);
xor U10752 (N_10752,N_9634,N_9827);
nand U10753 (N_10753,N_9525,N_9846);
nand U10754 (N_10754,N_9655,N_9426);
or U10755 (N_10755,N_9374,N_9855);
nor U10756 (N_10756,N_9411,N_9217);
or U10757 (N_10757,N_9917,N_9586);
nand U10758 (N_10758,N_9859,N_9772);
or U10759 (N_10759,N_9122,N_9082);
xnor U10760 (N_10760,N_9500,N_9545);
or U10761 (N_10761,N_9352,N_9384);
and U10762 (N_10762,N_9070,N_9710);
nor U10763 (N_10763,N_9766,N_9252);
nand U10764 (N_10764,N_9643,N_9724);
nor U10765 (N_10765,N_9815,N_9823);
and U10766 (N_10766,N_9221,N_9089);
nand U10767 (N_10767,N_9440,N_9195);
and U10768 (N_10768,N_9034,N_9240);
nand U10769 (N_10769,N_9723,N_9054);
and U10770 (N_10770,N_9559,N_9977);
and U10771 (N_10771,N_9529,N_9080);
nor U10772 (N_10772,N_9981,N_9781);
and U10773 (N_10773,N_9659,N_9076);
nor U10774 (N_10774,N_9874,N_9476);
and U10775 (N_10775,N_9769,N_9215);
xnor U10776 (N_10776,N_9171,N_9322);
nor U10777 (N_10777,N_9837,N_9063);
nor U10778 (N_10778,N_9239,N_9865);
and U10779 (N_10779,N_9187,N_9184);
xor U10780 (N_10780,N_9941,N_9025);
nand U10781 (N_10781,N_9990,N_9484);
nand U10782 (N_10782,N_9771,N_9596);
and U10783 (N_10783,N_9322,N_9983);
or U10784 (N_10784,N_9381,N_9275);
nand U10785 (N_10785,N_9859,N_9200);
xnor U10786 (N_10786,N_9036,N_9062);
nand U10787 (N_10787,N_9151,N_9938);
and U10788 (N_10788,N_9830,N_9826);
and U10789 (N_10789,N_9429,N_9513);
nor U10790 (N_10790,N_9548,N_9748);
xor U10791 (N_10791,N_9801,N_9359);
nand U10792 (N_10792,N_9586,N_9248);
nand U10793 (N_10793,N_9125,N_9406);
nor U10794 (N_10794,N_9590,N_9854);
xor U10795 (N_10795,N_9118,N_9426);
and U10796 (N_10796,N_9789,N_9837);
and U10797 (N_10797,N_9733,N_9784);
nor U10798 (N_10798,N_9820,N_9244);
and U10799 (N_10799,N_9059,N_9426);
or U10800 (N_10800,N_9215,N_9294);
or U10801 (N_10801,N_9769,N_9400);
or U10802 (N_10802,N_9092,N_9019);
nor U10803 (N_10803,N_9515,N_9614);
nor U10804 (N_10804,N_9378,N_9971);
nor U10805 (N_10805,N_9516,N_9969);
nor U10806 (N_10806,N_9879,N_9230);
and U10807 (N_10807,N_9362,N_9863);
nand U10808 (N_10808,N_9307,N_9722);
or U10809 (N_10809,N_9866,N_9062);
and U10810 (N_10810,N_9849,N_9188);
xor U10811 (N_10811,N_9337,N_9925);
or U10812 (N_10812,N_9561,N_9167);
nor U10813 (N_10813,N_9171,N_9503);
nand U10814 (N_10814,N_9274,N_9306);
nand U10815 (N_10815,N_9393,N_9512);
nor U10816 (N_10816,N_9623,N_9691);
nand U10817 (N_10817,N_9541,N_9299);
or U10818 (N_10818,N_9888,N_9072);
nor U10819 (N_10819,N_9377,N_9568);
or U10820 (N_10820,N_9784,N_9155);
nand U10821 (N_10821,N_9408,N_9283);
nor U10822 (N_10822,N_9830,N_9263);
nor U10823 (N_10823,N_9485,N_9566);
nor U10824 (N_10824,N_9482,N_9844);
and U10825 (N_10825,N_9240,N_9788);
nand U10826 (N_10826,N_9216,N_9124);
nor U10827 (N_10827,N_9286,N_9833);
and U10828 (N_10828,N_9464,N_9439);
or U10829 (N_10829,N_9857,N_9794);
or U10830 (N_10830,N_9573,N_9103);
and U10831 (N_10831,N_9347,N_9369);
or U10832 (N_10832,N_9195,N_9473);
nand U10833 (N_10833,N_9106,N_9554);
and U10834 (N_10834,N_9602,N_9519);
nor U10835 (N_10835,N_9065,N_9761);
or U10836 (N_10836,N_9836,N_9780);
nand U10837 (N_10837,N_9779,N_9431);
nand U10838 (N_10838,N_9813,N_9937);
or U10839 (N_10839,N_9380,N_9811);
nor U10840 (N_10840,N_9183,N_9372);
or U10841 (N_10841,N_9908,N_9219);
nor U10842 (N_10842,N_9732,N_9068);
and U10843 (N_10843,N_9583,N_9270);
nand U10844 (N_10844,N_9663,N_9767);
nand U10845 (N_10845,N_9437,N_9875);
nand U10846 (N_10846,N_9146,N_9359);
and U10847 (N_10847,N_9186,N_9940);
nand U10848 (N_10848,N_9184,N_9219);
and U10849 (N_10849,N_9297,N_9587);
nor U10850 (N_10850,N_9533,N_9794);
and U10851 (N_10851,N_9422,N_9347);
nand U10852 (N_10852,N_9485,N_9172);
and U10853 (N_10853,N_9772,N_9748);
nor U10854 (N_10854,N_9128,N_9210);
or U10855 (N_10855,N_9411,N_9070);
nand U10856 (N_10856,N_9290,N_9698);
xnor U10857 (N_10857,N_9196,N_9234);
xnor U10858 (N_10858,N_9154,N_9586);
nand U10859 (N_10859,N_9389,N_9139);
and U10860 (N_10860,N_9847,N_9147);
and U10861 (N_10861,N_9584,N_9718);
nor U10862 (N_10862,N_9922,N_9542);
or U10863 (N_10863,N_9574,N_9959);
nor U10864 (N_10864,N_9444,N_9145);
nand U10865 (N_10865,N_9716,N_9840);
nor U10866 (N_10866,N_9928,N_9698);
nor U10867 (N_10867,N_9349,N_9599);
nor U10868 (N_10868,N_9889,N_9959);
and U10869 (N_10869,N_9644,N_9744);
nor U10870 (N_10870,N_9622,N_9632);
nand U10871 (N_10871,N_9701,N_9262);
and U10872 (N_10872,N_9462,N_9723);
or U10873 (N_10873,N_9777,N_9066);
or U10874 (N_10874,N_9007,N_9428);
nand U10875 (N_10875,N_9072,N_9457);
and U10876 (N_10876,N_9639,N_9205);
or U10877 (N_10877,N_9222,N_9743);
nor U10878 (N_10878,N_9127,N_9836);
nor U10879 (N_10879,N_9997,N_9886);
xor U10880 (N_10880,N_9748,N_9304);
and U10881 (N_10881,N_9034,N_9227);
nand U10882 (N_10882,N_9651,N_9546);
or U10883 (N_10883,N_9622,N_9976);
or U10884 (N_10884,N_9355,N_9595);
nor U10885 (N_10885,N_9358,N_9531);
and U10886 (N_10886,N_9781,N_9656);
nand U10887 (N_10887,N_9721,N_9141);
nand U10888 (N_10888,N_9442,N_9291);
nand U10889 (N_10889,N_9207,N_9094);
and U10890 (N_10890,N_9540,N_9963);
or U10891 (N_10891,N_9044,N_9140);
nor U10892 (N_10892,N_9954,N_9079);
xnor U10893 (N_10893,N_9812,N_9913);
nor U10894 (N_10894,N_9251,N_9948);
nand U10895 (N_10895,N_9691,N_9275);
or U10896 (N_10896,N_9673,N_9232);
nor U10897 (N_10897,N_9187,N_9533);
nor U10898 (N_10898,N_9307,N_9801);
nand U10899 (N_10899,N_9575,N_9408);
or U10900 (N_10900,N_9348,N_9913);
nor U10901 (N_10901,N_9188,N_9580);
or U10902 (N_10902,N_9105,N_9108);
xnor U10903 (N_10903,N_9759,N_9977);
or U10904 (N_10904,N_9421,N_9672);
or U10905 (N_10905,N_9887,N_9546);
and U10906 (N_10906,N_9794,N_9727);
nand U10907 (N_10907,N_9930,N_9677);
nand U10908 (N_10908,N_9096,N_9401);
or U10909 (N_10909,N_9046,N_9245);
or U10910 (N_10910,N_9137,N_9757);
and U10911 (N_10911,N_9872,N_9314);
nand U10912 (N_10912,N_9837,N_9613);
nand U10913 (N_10913,N_9305,N_9190);
and U10914 (N_10914,N_9499,N_9947);
and U10915 (N_10915,N_9311,N_9355);
and U10916 (N_10916,N_9278,N_9132);
and U10917 (N_10917,N_9169,N_9031);
or U10918 (N_10918,N_9922,N_9439);
xnor U10919 (N_10919,N_9711,N_9199);
nor U10920 (N_10920,N_9013,N_9765);
nor U10921 (N_10921,N_9787,N_9002);
and U10922 (N_10922,N_9482,N_9144);
or U10923 (N_10923,N_9514,N_9204);
and U10924 (N_10924,N_9043,N_9653);
or U10925 (N_10925,N_9968,N_9156);
nor U10926 (N_10926,N_9830,N_9132);
nor U10927 (N_10927,N_9273,N_9686);
nand U10928 (N_10928,N_9308,N_9558);
xnor U10929 (N_10929,N_9698,N_9204);
nand U10930 (N_10930,N_9652,N_9208);
or U10931 (N_10931,N_9301,N_9241);
and U10932 (N_10932,N_9779,N_9100);
nand U10933 (N_10933,N_9111,N_9792);
nor U10934 (N_10934,N_9076,N_9552);
nand U10935 (N_10935,N_9876,N_9490);
and U10936 (N_10936,N_9016,N_9107);
and U10937 (N_10937,N_9011,N_9744);
nor U10938 (N_10938,N_9715,N_9969);
nand U10939 (N_10939,N_9658,N_9697);
nor U10940 (N_10940,N_9631,N_9945);
nand U10941 (N_10941,N_9247,N_9572);
nand U10942 (N_10942,N_9987,N_9255);
and U10943 (N_10943,N_9357,N_9408);
or U10944 (N_10944,N_9143,N_9941);
nand U10945 (N_10945,N_9869,N_9415);
nor U10946 (N_10946,N_9482,N_9832);
nand U10947 (N_10947,N_9304,N_9298);
xnor U10948 (N_10948,N_9825,N_9670);
nand U10949 (N_10949,N_9185,N_9821);
nand U10950 (N_10950,N_9848,N_9605);
nand U10951 (N_10951,N_9406,N_9643);
nand U10952 (N_10952,N_9612,N_9914);
nand U10953 (N_10953,N_9997,N_9027);
nand U10954 (N_10954,N_9131,N_9988);
nand U10955 (N_10955,N_9118,N_9029);
xnor U10956 (N_10956,N_9456,N_9681);
and U10957 (N_10957,N_9648,N_9871);
and U10958 (N_10958,N_9047,N_9606);
nor U10959 (N_10959,N_9072,N_9126);
nor U10960 (N_10960,N_9209,N_9345);
nor U10961 (N_10961,N_9908,N_9917);
or U10962 (N_10962,N_9705,N_9378);
nor U10963 (N_10963,N_9159,N_9491);
nor U10964 (N_10964,N_9910,N_9495);
xnor U10965 (N_10965,N_9370,N_9930);
or U10966 (N_10966,N_9379,N_9781);
or U10967 (N_10967,N_9245,N_9578);
or U10968 (N_10968,N_9323,N_9870);
or U10969 (N_10969,N_9115,N_9550);
nor U10970 (N_10970,N_9551,N_9521);
and U10971 (N_10971,N_9702,N_9112);
nor U10972 (N_10972,N_9776,N_9923);
or U10973 (N_10973,N_9103,N_9633);
xnor U10974 (N_10974,N_9314,N_9273);
or U10975 (N_10975,N_9923,N_9394);
and U10976 (N_10976,N_9298,N_9112);
nor U10977 (N_10977,N_9929,N_9037);
nor U10978 (N_10978,N_9588,N_9242);
and U10979 (N_10979,N_9453,N_9575);
nor U10980 (N_10980,N_9106,N_9561);
nor U10981 (N_10981,N_9486,N_9837);
or U10982 (N_10982,N_9691,N_9272);
nand U10983 (N_10983,N_9117,N_9799);
and U10984 (N_10984,N_9444,N_9178);
xnor U10985 (N_10985,N_9023,N_9049);
or U10986 (N_10986,N_9713,N_9234);
nor U10987 (N_10987,N_9449,N_9087);
xnor U10988 (N_10988,N_9494,N_9815);
and U10989 (N_10989,N_9044,N_9356);
and U10990 (N_10990,N_9583,N_9139);
or U10991 (N_10991,N_9559,N_9801);
nor U10992 (N_10992,N_9180,N_9398);
or U10993 (N_10993,N_9290,N_9243);
nor U10994 (N_10994,N_9879,N_9414);
nor U10995 (N_10995,N_9717,N_9494);
and U10996 (N_10996,N_9808,N_9529);
nor U10997 (N_10997,N_9146,N_9398);
nand U10998 (N_10998,N_9002,N_9859);
or U10999 (N_10999,N_9917,N_9308);
and U11000 (N_11000,N_10560,N_10120);
and U11001 (N_11001,N_10973,N_10235);
nor U11002 (N_11002,N_10159,N_10606);
nor U11003 (N_11003,N_10330,N_10852);
nor U11004 (N_11004,N_10699,N_10822);
nor U11005 (N_11005,N_10304,N_10201);
or U11006 (N_11006,N_10662,N_10217);
xnor U11007 (N_11007,N_10468,N_10811);
xor U11008 (N_11008,N_10173,N_10873);
xor U11009 (N_11009,N_10228,N_10910);
or U11010 (N_11010,N_10007,N_10947);
nand U11011 (N_11011,N_10067,N_10749);
nand U11012 (N_11012,N_10017,N_10506);
or U11013 (N_11013,N_10291,N_10970);
and U11014 (N_11014,N_10079,N_10729);
and U11015 (N_11015,N_10723,N_10820);
or U11016 (N_11016,N_10027,N_10510);
nand U11017 (N_11017,N_10272,N_10126);
or U11018 (N_11018,N_10100,N_10842);
or U11019 (N_11019,N_10562,N_10853);
or U11020 (N_11020,N_10222,N_10656);
and U11021 (N_11021,N_10630,N_10976);
nor U11022 (N_11022,N_10993,N_10406);
xor U11023 (N_11023,N_10798,N_10878);
nor U11024 (N_11024,N_10718,N_10472);
and U11025 (N_11025,N_10035,N_10755);
nor U11026 (N_11026,N_10646,N_10181);
and U11027 (N_11027,N_10554,N_10257);
and U11028 (N_11028,N_10380,N_10043);
or U11029 (N_11029,N_10887,N_10153);
or U11030 (N_11030,N_10770,N_10581);
nand U11031 (N_11031,N_10991,N_10174);
and U11032 (N_11032,N_10382,N_10183);
or U11033 (N_11033,N_10883,N_10907);
nand U11034 (N_11034,N_10195,N_10208);
or U11035 (N_11035,N_10081,N_10482);
and U11036 (N_11036,N_10545,N_10283);
nand U11037 (N_11037,N_10474,N_10941);
xnor U11038 (N_11038,N_10094,N_10564);
nor U11039 (N_11039,N_10525,N_10194);
nand U11040 (N_11040,N_10556,N_10899);
nand U11041 (N_11041,N_10660,N_10353);
nor U11042 (N_11042,N_10350,N_10744);
nand U11043 (N_11043,N_10867,N_10389);
nor U11044 (N_11044,N_10761,N_10651);
xor U11045 (N_11045,N_10552,N_10176);
nor U11046 (N_11046,N_10013,N_10689);
and U11047 (N_11047,N_10983,N_10050);
nor U11048 (N_11048,N_10819,N_10312);
nor U11049 (N_11049,N_10601,N_10693);
and U11050 (N_11050,N_10987,N_10597);
or U11051 (N_11051,N_10045,N_10727);
nand U11052 (N_11052,N_10609,N_10262);
or U11053 (N_11053,N_10835,N_10213);
nand U11054 (N_11054,N_10377,N_10197);
or U11055 (N_11055,N_10783,N_10487);
nand U11056 (N_11056,N_10064,N_10166);
nor U11057 (N_11057,N_10766,N_10704);
or U11058 (N_11058,N_10263,N_10860);
nand U11059 (N_11059,N_10369,N_10719);
or U11060 (N_11060,N_10955,N_10968);
xor U11061 (N_11061,N_10921,N_10354);
or U11062 (N_11062,N_10295,N_10300);
and U11063 (N_11063,N_10904,N_10908);
nand U11064 (N_11064,N_10703,N_10485);
or U11065 (N_11065,N_10521,N_10505);
nor U11066 (N_11066,N_10838,N_10072);
xnor U11067 (N_11067,N_10858,N_10490);
nor U11068 (N_11068,N_10573,N_10575);
nor U11069 (N_11069,N_10362,N_10401);
or U11070 (N_11070,N_10049,N_10368);
or U11071 (N_11071,N_10716,N_10998);
or U11072 (N_11072,N_10800,N_10239);
or U11073 (N_11073,N_10495,N_10163);
or U11074 (N_11074,N_10333,N_10306);
nor U11075 (N_11075,N_10781,N_10110);
nand U11076 (N_11076,N_10165,N_10958);
nor U11077 (N_11077,N_10203,N_10055);
and U11078 (N_11078,N_10636,N_10856);
and U11079 (N_11079,N_10548,N_10200);
or U11080 (N_11080,N_10150,N_10314);
and U11081 (N_11081,N_10956,N_10374);
or U11082 (N_11082,N_10850,N_10456);
nand U11083 (N_11083,N_10898,N_10501);
or U11084 (N_11084,N_10984,N_10315);
or U11085 (N_11085,N_10829,N_10011);
nand U11086 (N_11086,N_10642,N_10370);
nand U11087 (N_11087,N_10236,N_10441);
xnor U11088 (N_11088,N_10461,N_10765);
or U11089 (N_11089,N_10282,N_10204);
nand U11090 (N_11090,N_10386,N_10981);
nand U11091 (N_11091,N_10206,N_10894);
and U11092 (N_11092,N_10268,N_10182);
and U11093 (N_11093,N_10911,N_10445);
xor U11094 (N_11094,N_10667,N_10839);
and U11095 (N_11095,N_10298,N_10464);
xor U11096 (N_11096,N_10070,N_10435);
and U11097 (N_11097,N_10882,N_10058);
or U11098 (N_11098,N_10205,N_10982);
and U11099 (N_11099,N_10625,N_10613);
nor U11100 (N_11100,N_10476,N_10785);
xor U11101 (N_11101,N_10317,N_10791);
or U11102 (N_11102,N_10678,N_10149);
nor U11103 (N_11103,N_10226,N_10652);
xnor U11104 (N_11104,N_10683,N_10611);
xor U11105 (N_11105,N_10494,N_10713);
or U11106 (N_11106,N_10666,N_10457);
or U11107 (N_11107,N_10740,N_10881);
nand U11108 (N_11108,N_10837,N_10164);
or U11109 (N_11109,N_10021,N_10924);
and U11110 (N_11110,N_10534,N_10540);
and U11111 (N_11111,N_10864,N_10338);
and U11112 (N_11112,N_10014,N_10192);
nand U11113 (N_11113,N_10383,N_10877);
nor U11114 (N_11114,N_10057,N_10224);
nand U11115 (N_11115,N_10586,N_10722);
and U11116 (N_11116,N_10025,N_10539);
and U11117 (N_11117,N_10847,N_10780);
or U11118 (N_11118,N_10901,N_10020);
nor U11119 (N_11119,N_10367,N_10496);
or U11120 (N_11120,N_10786,N_10563);
nand U11121 (N_11121,N_10071,N_10391);
nand U11122 (N_11122,N_10725,N_10361);
or U11123 (N_11123,N_10331,N_10855);
nand U11124 (N_11124,N_10926,N_10509);
and U11125 (N_11125,N_10925,N_10458);
nor U11126 (N_11126,N_10797,N_10357);
nand U11127 (N_11127,N_10180,N_10107);
nand U11128 (N_11128,N_10433,N_10715);
or U11129 (N_11129,N_10516,N_10938);
and U11130 (N_11130,N_10591,N_10488);
nand U11131 (N_11131,N_10066,N_10913);
xnor U11132 (N_11132,N_10969,N_10570);
nor U11133 (N_11133,N_10615,N_10242);
or U11134 (N_11134,N_10631,N_10610);
xnor U11135 (N_11135,N_10426,N_10734);
nor U11136 (N_11136,N_10400,N_10264);
nor U11137 (N_11137,N_10408,N_10187);
nand U11138 (N_11138,N_10061,N_10019);
and U11139 (N_11139,N_10671,N_10604);
and U11140 (N_11140,N_10335,N_10274);
nand U11141 (N_11141,N_10479,N_10402);
xor U11142 (N_11142,N_10549,N_10674);
nand U11143 (N_11143,N_10161,N_10225);
or U11144 (N_11144,N_10238,N_10084);
nor U11145 (N_11145,N_10795,N_10395);
and U11146 (N_11146,N_10914,N_10717);
nand U11147 (N_11147,N_10568,N_10407);
or U11148 (N_11148,N_10919,N_10876);
nor U11149 (N_11149,N_10532,N_10831);
or U11150 (N_11150,N_10957,N_10828);
nor U11151 (N_11151,N_10483,N_10789);
and U11152 (N_11152,N_10909,N_10676);
nor U11153 (N_11153,N_10232,N_10720);
nor U11154 (N_11154,N_10305,N_10790);
or U11155 (N_11155,N_10207,N_10620);
or U11156 (N_11156,N_10841,N_10428);
and U11157 (N_11157,N_10307,N_10861);
xor U11158 (N_11158,N_10098,N_10945);
or U11159 (N_11159,N_10803,N_10088);
nor U11160 (N_11160,N_10612,N_10854);
or U11161 (N_11161,N_10296,N_10934);
and U11162 (N_11162,N_10470,N_10536);
nand U11163 (N_11163,N_10677,N_10246);
or U11164 (N_11164,N_10409,N_10808);
nor U11165 (N_11165,N_10352,N_10256);
nand U11166 (N_11166,N_10709,N_10275);
and U11167 (N_11167,N_10885,N_10292);
or U11168 (N_11168,N_10289,N_10348);
nand U11169 (N_11169,N_10942,N_10809);
nor U11170 (N_11170,N_10669,N_10608);
or U11171 (N_11171,N_10721,N_10139);
or U11172 (N_11172,N_10096,N_10845);
nor U11173 (N_11173,N_10451,N_10453);
nor U11174 (N_11174,N_10933,N_10245);
xor U11175 (N_11175,N_10134,N_10129);
and U11176 (N_11176,N_10221,N_10840);
or U11177 (N_11177,N_10237,N_10844);
or U11178 (N_11178,N_10138,N_10114);
and U11179 (N_11179,N_10497,N_10869);
or U11180 (N_11180,N_10290,N_10018);
nor U11181 (N_11181,N_10706,N_10574);
nand U11182 (N_11182,N_10069,N_10223);
and U11183 (N_11183,N_10321,N_10429);
and U11184 (N_11184,N_10042,N_10133);
xnor U11185 (N_11185,N_10392,N_10846);
or U11186 (N_11186,N_10452,N_10661);
and U11187 (N_11187,N_10424,N_10893);
or U11188 (N_11188,N_10123,N_10041);
and U11189 (N_11189,N_10896,N_10614);
or U11190 (N_11190,N_10737,N_10892);
nor U11191 (N_11191,N_10454,N_10710);
or U11192 (N_11192,N_10449,N_10818);
nor U11193 (N_11193,N_10147,N_10111);
or U11194 (N_11194,N_10437,N_10112);
nor U11195 (N_11195,N_10657,N_10022);
nor U11196 (N_11196,N_10310,N_10447);
and U11197 (N_11197,N_10641,N_10355);
or U11198 (N_11198,N_10588,N_10393);
and U11199 (N_11199,N_10448,N_10154);
or U11200 (N_11200,N_10169,N_10834);
nor U11201 (N_11201,N_10279,N_10028);
nor U11202 (N_11202,N_10439,N_10008);
and U11203 (N_11203,N_10253,N_10423);
nor U11204 (N_11204,N_10463,N_10210);
nand U11205 (N_11205,N_10682,N_10686);
and U11206 (N_11206,N_10879,N_10059);
xnor U11207 (N_11207,N_10137,N_10051);
or U11208 (N_11208,N_10503,N_10384);
nor U11209 (N_11209,N_10036,N_10168);
or U11210 (N_11210,N_10932,N_10280);
nor U11211 (N_11211,N_10813,N_10080);
and U11212 (N_11212,N_10623,N_10214);
nor U11213 (N_11213,N_10889,N_10326);
xnor U11214 (N_11214,N_10155,N_10076);
nor U11215 (N_11215,N_10171,N_10373);
nand U11216 (N_11216,N_10916,N_10178);
nor U11217 (N_11217,N_10594,N_10266);
and U11218 (N_11218,N_10915,N_10319);
nor U11219 (N_11219,N_10005,N_10190);
nor U11220 (N_11220,N_10775,N_10157);
nand U11221 (N_11221,N_10012,N_10985);
nor U11222 (N_11222,N_10696,N_10757);
nand U11223 (N_11223,N_10923,N_10986);
nor U11224 (N_11224,N_10052,N_10030);
and U11225 (N_11225,N_10273,N_10550);
xnor U11226 (N_11226,N_10705,N_10888);
and U11227 (N_11227,N_10640,N_10796);
nand U11228 (N_11228,N_10342,N_10471);
and U11229 (N_11229,N_10566,N_10989);
or U11230 (N_11230,N_10376,N_10927);
or U11231 (N_11231,N_10950,N_10607);
and U11232 (N_11232,N_10015,N_10799);
nor U11233 (N_11233,N_10432,N_10480);
or U11234 (N_11234,N_10996,N_10121);
or U11235 (N_11235,N_10438,N_10249);
and U11236 (N_11236,N_10443,N_10124);
and U11237 (N_11237,N_10978,N_10928);
and U11238 (N_11238,N_10177,N_10038);
nand U11239 (N_11239,N_10113,N_10430);
nor U11240 (N_11240,N_10587,N_10356);
and U11241 (N_11241,N_10068,N_10762);
or U11242 (N_11242,N_10959,N_10009);
and U11243 (N_11243,N_10427,N_10037);
and U11244 (N_11244,N_10465,N_10596);
nor U11245 (N_11245,N_10397,N_10824);
and U11246 (N_11246,N_10450,N_10106);
and U11247 (N_11247,N_10347,N_10087);
or U11248 (N_11248,N_10814,N_10833);
and U11249 (N_11249,N_10297,N_10742);
and U11250 (N_11250,N_10815,N_10507);
nor U11251 (N_11251,N_10118,N_10063);
and U11252 (N_11252,N_10329,N_10684);
nand U11253 (N_11253,N_10980,N_10672);
nand U11254 (N_11254,N_10000,N_10131);
nand U11255 (N_11255,N_10967,N_10621);
xor U11256 (N_11256,N_10936,N_10508);
nand U11257 (N_11257,N_10255,N_10364);
nand U11258 (N_11258,N_10579,N_10251);
or U11259 (N_11259,N_10880,N_10031);
xnor U11260 (N_11260,N_10387,N_10241);
nor U11261 (N_11261,N_10002,N_10416);
or U11262 (N_11262,N_10234,N_10431);
nor U11263 (N_11263,N_10125,N_10874);
or U11264 (N_11264,N_10240,N_10092);
and U11265 (N_11265,N_10086,N_10953);
or U11266 (N_11266,N_10460,N_10943);
or U11267 (N_11267,N_10977,N_10685);
nor U11268 (N_11268,N_10769,N_10590);
nand U11269 (N_11269,N_10931,N_10378);
and U11270 (N_11270,N_10743,N_10616);
nor U11271 (N_11271,N_10673,N_10363);
nand U11272 (N_11272,N_10692,N_10638);
nand U11273 (N_11273,N_10836,N_10862);
or U11274 (N_11274,N_10127,N_10412);
nor U11275 (N_11275,N_10645,N_10812);
nand U11276 (N_11276,N_10248,N_10475);
nor U11277 (N_11277,N_10848,N_10804);
or U11278 (N_11278,N_10542,N_10714);
nand U11279 (N_11279,N_10186,N_10884);
nor U11280 (N_11280,N_10261,N_10327);
or U11281 (N_11281,N_10140,N_10966);
xnor U11282 (N_11282,N_10425,N_10158);
and U11283 (N_11283,N_10083,N_10773);
or U11284 (N_11284,N_10229,N_10293);
nor U11285 (N_11285,N_10659,N_10128);
and U11286 (N_11286,N_10940,N_10039);
and U11287 (N_11287,N_10648,N_10738);
nor U11288 (N_11288,N_10951,N_10859);
and U11289 (N_11289,N_10593,N_10029);
or U11290 (N_11290,N_10336,N_10767);
or U11291 (N_11291,N_10250,N_10708);
or U11292 (N_11292,N_10422,N_10230);
and U11293 (N_11293,N_10857,N_10537);
nor U11294 (N_11294,N_10750,N_10351);
nor U11295 (N_11295,N_10371,N_10961);
nor U11296 (N_11296,N_10417,N_10477);
nand U11297 (N_11297,N_10849,N_10196);
and U11298 (N_11298,N_10414,N_10979);
or U11299 (N_11299,N_10481,N_10900);
or U11300 (N_11300,N_10584,N_10075);
nor U11301 (N_11301,N_10340,N_10366);
and U11302 (N_11302,N_10675,N_10325);
xnor U11303 (N_11303,N_10459,N_10466);
or U11304 (N_11304,N_10047,N_10776);
nor U11305 (N_11305,N_10269,N_10751);
or U11306 (N_11306,N_10191,N_10040);
nand U11307 (N_11307,N_10633,N_10258);
nor U11308 (N_11308,N_10992,N_10555);
or U11309 (N_11309,N_10130,N_10440);
nor U11310 (N_11310,N_10313,N_10152);
and U11311 (N_11311,N_10294,N_10572);
and U11312 (N_11312,N_10753,N_10632);
nand U11313 (N_11313,N_10654,N_10649);
and U11314 (N_11314,N_10394,N_10865);
xnor U11315 (N_11315,N_10247,N_10747);
xor U11316 (N_11316,N_10619,N_10054);
nand U11317 (N_11317,N_10895,N_10419);
xnor U11318 (N_11318,N_10082,N_10745);
xor U11319 (N_11319,N_10736,N_10023);
or U11320 (N_11320,N_10792,N_10135);
or U11321 (N_11321,N_10276,N_10694);
nand U11322 (N_11322,N_10920,N_10288);
nand U11323 (N_11323,N_10172,N_10341);
or U11324 (N_11324,N_10185,N_10965);
nand U11325 (N_11325,N_10949,N_10801);
and U11326 (N_11326,N_10974,N_10493);
nand U11327 (N_11327,N_10491,N_10418);
or U11328 (N_11328,N_10184,N_10870);
nor U11329 (N_11329,N_10639,N_10758);
xor U11330 (N_11330,N_10546,N_10323);
nor U11331 (N_11331,N_10498,N_10522);
nor U11332 (N_11332,N_10752,N_10148);
nand U11333 (N_11333,N_10700,N_10517);
nand U11334 (N_11334,N_10810,N_10379);
or U11335 (N_11335,N_10571,N_10193);
nand U11336 (N_11336,N_10115,N_10243);
nand U11337 (N_11337,N_10216,N_10089);
or U11338 (N_11338,N_10337,N_10284);
nor U11339 (N_11339,N_10697,N_10093);
nand U11340 (N_11340,N_10411,N_10658);
nand U11341 (N_11341,N_10772,N_10760);
and U11342 (N_11342,N_10175,N_10287);
nand U11343 (N_11343,N_10918,N_10444);
or U11344 (N_11344,N_10375,N_10102);
xor U11345 (N_11345,N_10360,N_10455);
nand U11346 (N_11346,N_10782,N_10599);
and U11347 (N_11347,N_10119,N_10167);
or U11348 (N_11348,N_10764,N_10954);
and U11349 (N_11349,N_10339,N_10467);
nand U11350 (N_11350,N_10567,N_10531);
xnor U11351 (N_11351,N_10866,N_10538);
nand U11352 (N_11352,N_10345,N_10144);
nand U11353 (N_11353,N_10917,N_10664);
xnor U11354 (N_11354,N_10141,N_10695);
or U11355 (N_11355,N_10891,N_10372);
or U11356 (N_11356,N_10502,N_10929);
nand U11357 (N_11357,N_10922,N_10711);
nor U11358 (N_11358,N_10712,N_10544);
nor U11359 (N_11359,N_10044,N_10099);
or U11360 (N_11360,N_10421,N_10944);
or U11361 (N_11361,N_10626,N_10589);
or U11362 (N_11362,N_10863,N_10504);
or U11363 (N_11363,N_10827,N_10142);
nor U11364 (N_11364,N_10647,N_10385);
or U11365 (N_11365,N_10033,N_10524);
and U11366 (N_11366,N_10930,N_10188);
and U11367 (N_11367,N_10543,N_10788);
nand U11368 (N_11368,N_10231,N_10787);
or U11369 (N_11369,N_10533,N_10730);
nor U11370 (N_11370,N_10309,N_10817);
nor U11371 (N_11371,N_10390,N_10077);
or U11372 (N_11372,N_10260,N_10964);
nand U11373 (N_11373,N_10301,N_10832);
and U11374 (N_11374,N_10644,N_10999);
nor U11375 (N_11375,N_10816,N_10806);
or U11376 (N_11376,N_10101,N_10592);
nand U11377 (N_11377,N_10060,N_10016);
and U11378 (N_11378,N_10048,N_10617);
nand U11379 (N_11379,N_10807,N_10062);
or U11380 (N_11380,N_10547,N_10605);
nor U11381 (N_11381,N_10344,N_10702);
nor U11382 (N_11382,N_10551,N_10117);
and U11383 (N_11383,N_10473,N_10523);
nand U11384 (N_11384,N_10558,N_10960);
nand U11385 (N_11385,N_10024,N_10270);
nor U11386 (N_11386,N_10988,N_10489);
or U11387 (N_11387,N_10436,N_10346);
or U11388 (N_11388,N_10332,N_10526);
xnor U11389 (N_11389,N_10687,N_10219);
nor U11390 (N_11390,N_10122,N_10939);
nor U11391 (N_11391,N_10872,N_10299);
nor U11392 (N_11392,N_10768,N_10146);
nand U11393 (N_11393,N_10034,N_10541);
nand U11394 (N_11394,N_10211,N_10320);
nor U11395 (N_11395,N_10726,N_10132);
or U11396 (N_11396,N_10629,N_10912);
and U11397 (N_11397,N_10267,N_10032);
nor U11398 (N_11398,N_10278,N_10316);
and U11399 (N_11399,N_10618,N_10583);
xor U11400 (N_11400,N_10212,N_10679);
nor U11401 (N_11401,N_10779,N_10784);
nor U11402 (N_11402,N_10759,N_10559);
nor U11403 (N_11403,N_10569,N_10830);
or U11404 (N_11404,N_10143,N_10162);
or U11405 (N_11405,N_10997,N_10868);
and U11406 (N_11406,N_10303,N_10793);
or U11407 (N_11407,N_10499,N_10655);
nand U11408 (N_11408,N_10359,N_10650);
and U11409 (N_11409,N_10680,N_10091);
nor U11410 (N_11410,N_10160,N_10688);
nand U11411 (N_11411,N_10511,N_10513);
or U11412 (N_11412,N_10553,N_10358);
nor U11413 (N_11413,N_10116,N_10199);
nor U11414 (N_11414,N_10001,N_10698);
nand U11415 (N_11415,N_10518,N_10681);
nand U11416 (N_11416,N_10906,N_10890);
nand U11417 (N_11417,N_10871,N_10886);
or U11418 (N_11418,N_10635,N_10156);
nor U11419 (N_11419,N_10622,N_10778);
or U11420 (N_11420,N_10771,N_10311);
and U11421 (N_11421,N_10582,N_10963);
nand U11422 (N_11422,N_10962,N_10410);
or U11423 (N_11423,N_10634,N_10946);
or U11424 (N_11424,N_10535,N_10090);
xnor U11425 (N_11425,N_10218,N_10794);
nand U11426 (N_11426,N_10302,N_10937);
and U11427 (N_11427,N_10690,N_10396);
nor U11428 (N_11428,N_10821,N_10281);
or U11429 (N_11429,N_10739,N_10561);
or U11430 (N_11430,N_10520,N_10971);
or U11431 (N_11431,N_10254,N_10073);
or U11432 (N_11432,N_10724,N_10046);
or U11433 (N_11433,N_10349,N_10732);
or U11434 (N_11434,N_10065,N_10434);
or U11435 (N_11435,N_10136,N_10565);
nand U11436 (N_11436,N_10628,N_10823);
nand U11437 (N_11437,N_10733,N_10670);
nor U11438 (N_11438,N_10209,N_10486);
nand U11439 (N_11439,N_10825,N_10994);
and U11440 (N_11440,N_10010,N_10668);
or U11441 (N_11441,N_10585,N_10665);
nand U11442 (N_11442,N_10515,N_10478);
or U11443 (N_11443,N_10624,N_10598);
or U11444 (N_11444,N_10442,N_10663);
and U11445 (N_11445,N_10577,N_10826);
nor U11446 (N_11446,N_10003,N_10578);
nand U11447 (N_11447,N_10420,N_10653);
nor U11448 (N_11448,N_10995,N_10843);
and U11449 (N_11449,N_10735,N_10691);
and U11450 (N_11450,N_10006,N_10602);
nor U11451 (N_11451,N_10948,N_10179);
nor U11452 (N_11452,N_10802,N_10603);
nor U11453 (N_11453,N_10286,N_10085);
nor U11454 (N_11454,N_10754,N_10056);
nor U11455 (N_11455,N_10170,N_10053);
and U11456 (N_11456,N_10756,N_10805);
nand U11457 (N_11457,N_10233,N_10381);
nand U11458 (N_11458,N_10728,N_10905);
and U11459 (N_11459,N_10469,N_10777);
nor U11460 (N_11460,N_10701,N_10519);
and U11461 (N_11461,N_10103,N_10271);
and U11462 (N_11462,N_10576,N_10202);
xnor U11463 (N_11463,N_10514,N_10935);
nor U11464 (N_11464,N_10500,N_10707);
nor U11465 (N_11465,N_10328,N_10198);
nor U11466 (N_11466,N_10600,N_10763);
and U11467 (N_11467,N_10415,N_10637);
xnor U11468 (N_11468,N_10902,N_10074);
and U11469 (N_11469,N_10026,N_10189);
nor U11470 (N_11470,N_10972,N_10643);
and U11471 (N_11471,N_10227,N_10215);
nor U11472 (N_11472,N_10952,N_10530);
nor U11473 (N_11473,N_10484,N_10151);
nor U11474 (N_11474,N_10557,N_10078);
nand U11475 (N_11475,N_10324,N_10975);
and U11476 (N_11476,N_10145,N_10108);
or U11477 (N_11477,N_10004,N_10741);
nand U11478 (N_11478,N_10109,N_10104);
nand U11479 (N_11479,N_10446,N_10595);
nor U11480 (N_11480,N_10244,N_10220);
nor U11481 (N_11481,N_10265,N_10095);
or U11482 (N_11482,N_10405,N_10851);
and U11483 (N_11483,N_10462,N_10399);
and U11484 (N_11484,N_10388,N_10748);
nand U11485 (N_11485,N_10990,N_10259);
nor U11486 (N_11486,N_10529,N_10403);
nor U11487 (N_11487,N_10334,N_10285);
nor U11488 (N_11488,N_10398,N_10252);
nor U11489 (N_11489,N_10413,N_10365);
nand U11490 (N_11490,N_10731,N_10322);
nand U11491 (N_11491,N_10746,N_10512);
nand U11492 (N_11492,N_10527,N_10404);
nand U11493 (N_11493,N_10580,N_10528);
nor U11494 (N_11494,N_10897,N_10492);
and U11495 (N_11495,N_10343,N_10774);
nand U11496 (N_11496,N_10308,N_10903);
and U11497 (N_11497,N_10627,N_10097);
nor U11498 (N_11498,N_10875,N_10105);
nand U11499 (N_11499,N_10318,N_10277);
and U11500 (N_11500,N_10879,N_10382);
xnor U11501 (N_11501,N_10374,N_10913);
or U11502 (N_11502,N_10863,N_10409);
or U11503 (N_11503,N_10572,N_10498);
nor U11504 (N_11504,N_10409,N_10032);
nor U11505 (N_11505,N_10065,N_10186);
and U11506 (N_11506,N_10552,N_10290);
and U11507 (N_11507,N_10044,N_10726);
xor U11508 (N_11508,N_10554,N_10627);
nand U11509 (N_11509,N_10228,N_10608);
xor U11510 (N_11510,N_10053,N_10321);
and U11511 (N_11511,N_10060,N_10017);
nor U11512 (N_11512,N_10909,N_10631);
nor U11513 (N_11513,N_10637,N_10189);
or U11514 (N_11514,N_10343,N_10589);
nor U11515 (N_11515,N_10294,N_10755);
and U11516 (N_11516,N_10373,N_10300);
and U11517 (N_11517,N_10932,N_10194);
and U11518 (N_11518,N_10439,N_10505);
nor U11519 (N_11519,N_10789,N_10383);
nor U11520 (N_11520,N_10738,N_10685);
xnor U11521 (N_11521,N_10023,N_10457);
xor U11522 (N_11522,N_10847,N_10974);
nor U11523 (N_11523,N_10748,N_10215);
nand U11524 (N_11524,N_10391,N_10270);
or U11525 (N_11525,N_10930,N_10091);
nand U11526 (N_11526,N_10604,N_10002);
or U11527 (N_11527,N_10836,N_10260);
and U11528 (N_11528,N_10555,N_10129);
and U11529 (N_11529,N_10643,N_10777);
nor U11530 (N_11530,N_10682,N_10377);
nand U11531 (N_11531,N_10111,N_10312);
nor U11532 (N_11532,N_10833,N_10777);
nand U11533 (N_11533,N_10080,N_10207);
or U11534 (N_11534,N_10655,N_10358);
and U11535 (N_11535,N_10160,N_10841);
and U11536 (N_11536,N_10787,N_10823);
and U11537 (N_11537,N_10462,N_10338);
nand U11538 (N_11538,N_10313,N_10052);
and U11539 (N_11539,N_10629,N_10816);
nand U11540 (N_11540,N_10292,N_10848);
nor U11541 (N_11541,N_10970,N_10487);
nand U11542 (N_11542,N_10335,N_10779);
nand U11543 (N_11543,N_10491,N_10902);
nor U11544 (N_11544,N_10550,N_10113);
nor U11545 (N_11545,N_10672,N_10143);
or U11546 (N_11546,N_10948,N_10574);
nor U11547 (N_11547,N_10950,N_10153);
or U11548 (N_11548,N_10968,N_10250);
or U11549 (N_11549,N_10692,N_10891);
and U11550 (N_11550,N_10404,N_10819);
or U11551 (N_11551,N_10102,N_10084);
nand U11552 (N_11552,N_10499,N_10736);
or U11553 (N_11553,N_10429,N_10008);
nor U11554 (N_11554,N_10760,N_10196);
and U11555 (N_11555,N_10688,N_10079);
nor U11556 (N_11556,N_10543,N_10578);
xor U11557 (N_11557,N_10983,N_10577);
nor U11558 (N_11558,N_10504,N_10198);
xnor U11559 (N_11559,N_10235,N_10334);
and U11560 (N_11560,N_10799,N_10105);
xor U11561 (N_11561,N_10443,N_10405);
and U11562 (N_11562,N_10709,N_10600);
and U11563 (N_11563,N_10463,N_10329);
or U11564 (N_11564,N_10934,N_10348);
nand U11565 (N_11565,N_10940,N_10481);
nor U11566 (N_11566,N_10442,N_10401);
xor U11567 (N_11567,N_10216,N_10236);
nand U11568 (N_11568,N_10195,N_10441);
or U11569 (N_11569,N_10767,N_10876);
and U11570 (N_11570,N_10597,N_10119);
and U11571 (N_11571,N_10289,N_10546);
nor U11572 (N_11572,N_10615,N_10937);
or U11573 (N_11573,N_10590,N_10322);
nand U11574 (N_11574,N_10394,N_10985);
nor U11575 (N_11575,N_10235,N_10372);
xor U11576 (N_11576,N_10092,N_10897);
and U11577 (N_11577,N_10447,N_10990);
or U11578 (N_11578,N_10879,N_10206);
nor U11579 (N_11579,N_10955,N_10127);
nand U11580 (N_11580,N_10824,N_10665);
or U11581 (N_11581,N_10463,N_10823);
nor U11582 (N_11582,N_10903,N_10331);
nand U11583 (N_11583,N_10866,N_10833);
nor U11584 (N_11584,N_10221,N_10342);
nand U11585 (N_11585,N_10719,N_10249);
and U11586 (N_11586,N_10469,N_10789);
nor U11587 (N_11587,N_10471,N_10001);
and U11588 (N_11588,N_10214,N_10567);
or U11589 (N_11589,N_10511,N_10115);
or U11590 (N_11590,N_10014,N_10601);
and U11591 (N_11591,N_10718,N_10541);
nor U11592 (N_11592,N_10858,N_10028);
or U11593 (N_11593,N_10589,N_10321);
nor U11594 (N_11594,N_10784,N_10253);
nor U11595 (N_11595,N_10077,N_10999);
or U11596 (N_11596,N_10053,N_10901);
nor U11597 (N_11597,N_10022,N_10689);
nand U11598 (N_11598,N_10414,N_10619);
nand U11599 (N_11599,N_10800,N_10618);
nor U11600 (N_11600,N_10185,N_10707);
or U11601 (N_11601,N_10459,N_10785);
and U11602 (N_11602,N_10187,N_10228);
nor U11603 (N_11603,N_10680,N_10116);
and U11604 (N_11604,N_10423,N_10908);
xnor U11605 (N_11605,N_10233,N_10296);
xor U11606 (N_11606,N_10876,N_10390);
xor U11607 (N_11607,N_10699,N_10278);
nand U11608 (N_11608,N_10045,N_10372);
and U11609 (N_11609,N_10701,N_10466);
or U11610 (N_11610,N_10016,N_10629);
nand U11611 (N_11611,N_10111,N_10744);
or U11612 (N_11612,N_10531,N_10700);
and U11613 (N_11613,N_10771,N_10770);
and U11614 (N_11614,N_10930,N_10947);
nand U11615 (N_11615,N_10444,N_10462);
or U11616 (N_11616,N_10569,N_10498);
nand U11617 (N_11617,N_10406,N_10568);
nor U11618 (N_11618,N_10941,N_10293);
and U11619 (N_11619,N_10967,N_10723);
nor U11620 (N_11620,N_10572,N_10325);
or U11621 (N_11621,N_10432,N_10813);
nand U11622 (N_11622,N_10468,N_10828);
or U11623 (N_11623,N_10280,N_10431);
nor U11624 (N_11624,N_10283,N_10185);
and U11625 (N_11625,N_10049,N_10486);
or U11626 (N_11626,N_10657,N_10061);
or U11627 (N_11627,N_10712,N_10723);
and U11628 (N_11628,N_10176,N_10954);
or U11629 (N_11629,N_10975,N_10699);
and U11630 (N_11630,N_10262,N_10384);
nand U11631 (N_11631,N_10679,N_10084);
or U11632 (N_11632,N_10275,N_10774);
or U11633 (N_11633,N_10365,N_10105);
nand U11634 (N_11634,N_10415,N_10913);
xnor U11635 (N_11635,N_10929,N_10967);
xor U11636 (N_11636,N_10954,N_10353);
nand U11637 (N_11637,N_10528,N_10932);
and U11638 (N_11638,N_10489,N_10687);
xnor U11639 (N_11639,N_10707,N_10611);
or U11640 (N_11640,N_10537,N_10791);
and U11641 (N_11641,N_10762,N_10674);
nor U11642 (N_11642,N_10656,N_10601);
nor U11643 (N_11643,N_10526,N_10046);
nand U11644 (N_11644,N_10569,N_10524);
nand U11645 (N_11645,N_10008,N_10241);
nand U11646 (N_11646,N_10821,N_10177);
and U11647 (N_11647,N_10163,N_10280);
nor U11648 (N_11648,N_10931,N_10884);
and U11649 (N_11649,N_10492,N_10394);
nand U11650 (N_11650,N_10556,N_10601);
or U11651 (N_11651,N_10027,N_10597);
and U11652 (N_11652,N_10710,N_10012);
nand U11653 (N_11653,N_10087,N_10120);
nand U11654 (N_11654,N_10184,N_10174);
and U11655 (N_11655,N_10400,N_10141);
and U11656 (N_11656,N_10070,N_10799);
and U11657 (N_11657,N_10243,N_10639);
nor U11658 (N_11658,N_10324,N_10587);
nor U11659 (N_11659,N_10876,N_10475);
and U11660 (N_11660,N_10243,N_10264);
or U11661 (N_11661,N_10943,N_10914);
or U11662 (N_11662,N_10569,N_10577);
nand U11663 (N_11663,N_10760,N_10164);
nand U11664 (N_11664,N_10943,N_10510);
xnor U11665 (N_11665,N_10130,N_10962);
nand U11666 (N_11666,N_10989,N_10794);
and U11667 (N_11667,N_10566,N_10332);
and U11668 (N_11668,N_10871,N_10890);
nand U11669 (N_11669,N_10628,N_10952);
or U11670 (N_11670,N_10344,N_10728);
and U11671 (N_11671,N_10263,N_10636);
nand U11672 (N_11672,N_10568,N_10878);
and U11673 (N_11673,N_10848,N_10673);
nor U11674 (N_11674,N_10906,N_10141);
and U11675 (N_11675,N_10878,N_10576);
nor U11676 (N_11676,N_10717,N_10807);
and U11677 (N_11677,N_10345,N_10436);
or U11678 (N_11678,N_10825,N_10446);
nor U11679 (N_11679,N_10588,N_10833);
nand U11680 (N_11680,N_10999,N_10187);
nor U11681 (N_11681,N_10254,N_10500);
nand U11682 (N_11682,N_10036,N_10914);
nand U11683 (N_11683,N_10892,N_10063);
xnor U11684 (N_11684,N_10041,N_10264);
and U11685 (N_11685,N_10467,N_10268);
and U11686 (N_11686,N_10203,N_10174);
xor U11687 (N_11687,N_10827,N_10120);
nand U11688 (N_11688,N_10005,N_10812);
nor U11689 (N_11689,N_10857,N_10507);
xor U11690 (N_11690,N_10158,N_10266);
nand U11691 (N_11691,N_10620,N_10938);
nand U11692 (N_11692,N_10855,N_10703);
xor U11693 (N_11693,N_10460,N_10107);
nand U11694 (N_11694,N_10426,N_10268);
and U11695 (N_11695,N_10550,N_10142);
nor U11696 (N_11696,N_10366,N_10711);
nor U11697 (N_11697,N_10845,N_10882);
or U11698 (N_11698,N_10004,N_10812);
or U11699 (N_11699,N_10265,N_10428);
nand U11700 (N_11700,N_10937,N_10437);
nand U11701 (N_11701,N_10360,N_10471);
and U11702 (N_11702,N_10998,N_10755);
xnor U11703 (N_11703,N_10048,N_10777);
or U11704 (N_11704,N_10884,N_10090);
and U11705 (N_11705,N_10330,N_10516);
or U11706 (N_11706,N_10446,N_10930);
nand U11707 (N_11707,N_10419,N_10421);
or U11708 (N_11708,N_10382,N_10960);
nor U11709 (N_11709,N_10990,N_10509);
or U11710 (N_11710,N_10872,N_10980);
or U11711 (N_11711,N_10820,N_10071);
nor U11712 (N_11712,N_10429,N_10739);
nor U11713 (N_11713,N_10469,N_10633);
or U11714 (N_11714,N_10619,N_10980);
nor U11715 (N_11715,N_10563,N_10395);
nand U11716 (N_11716,N_10570,N_10698);
xnor U11717 (N_11717,N_10899,N_10196);
or U11718 (N_11718,N_10938,N_10835);
and U11719 (N_11719,N_10085,N_10060);
nand U11720 (N_11720,N_10095,N_10524);
nand U11721 (N_11721,N_10480,N_10710);
nand U11722 (N_11722,N_10421,N_10863);
or U11723 (N_11723,N_10428,N_10719);
nand U11724 (N_11724,N_10813,N_10322);
nand U11725 (N_11725,N_10508,N_10340);
nand U11726 (N_11726,N_10079,N_10523);
or U11727 (N_11727,N_10252,N_10183);
xnor U11728 (N_11728,N_10454,N_10867);
or U11729 (N_11729,N_10736,N_10728);
and U11730 (N_11730,N_10910,N_10216);
nor U11731 (N_11731,N_10025,N_10151);
and U11732 (N_11732,N_10583,N_10953);
nor U11733 (N_11733,N_10951,N_10382);
nor U11734 (N_11734,N_10061,N_10892);
nand U11735 (N_11735,N_10330,N_10522);
nand U11736 (N_11736,N_10531,N_10893);
xor U11737 (N_11737,N_10906,N_10763);
and U11738 (N_11738,N_10655,N_10066);
or U11739 (N_11739,N_10284,N_10589);
and U11740 (N_11740,N_10895,N_10558);
and U11741 (N_11741,N_10179,N_10200);
nor U11742 (N_11742,N_10757,N_10893);
nor U11743 (N_11743,N_10492,N_10744);
nor U11744 (N_11744,N_10287,N_10758);
nand U11745 (N_11745,N_10799,N_10679);
or U11746 (N_11746,N_10174,N_10094);
or U11747 (N_11747,N_10263,N_10378);
and U11748 (N_11748,N_10351,N_10560);
or U11749 (N_11749,N_10726,N_10422);
and U11750 (N_11750,N_10157,N_10076);
nand U11751 (N_11751,N_10281,N_10324);
nand U11752 (N_11752,N_10442,N_10195);
and U11753 (N_11753,N_10457,N_10945);
nand U11754 (N_11754,N_10903,N_10645);
xor U11755 (N_11755,N_10847,N_10846);
nor U11756 (N_11756,N_10487,N_10404);
nor U11757 (N_11757,N_10223,N_10230);
nand U11758 (N_11758,N_10410,N_10340);
and U11759 (N_11759,N_10817,N_10580);
and U11760 (N_11760,N_10466,N_10714);
and U11761 (N_11761,N_10118,N_10572);
and U11762 (N_11762,N_10606,N_10594);
or U11763 (N_11763,N_10429,N_10559);
xor U11764 (N_11764,N_10169,N_10163);
or U11765 (N_11765,N_10736,N_10539);
and U11766 (N_11766,N_10891,N_10224);
and U11767 (N_11767,N_10763,N_10968);
or U11768 (N_11768,N_10580,N_10999);
or U11769 (N_11769,N_10803,N_10881);
nor U11770 (N_11770,N_10805,N_10564);
nor U11771 (N_11771,N_10718,N_10416);
and U11772 (N_11772,N_10400,N_10448);
and U11773 (N_11773,N_10295,N_10944);
nor U11774 (N_11774,N_10373,N_10614);
or U11775 (N_11775,N_10300,N_10002);
nor U11776 (N_11776,N_10484,N_10853);
or U11777 (N_11777,N_10816,N_10194);
nand U11778 (N_11778,N_10877,N_10257);
nand U11779 (N_11779,N_10817,N_10365);
and U11780 (N_11780,N_10420,N_10241);
or U11781 (N_11781,N_10344,N_10868);
nand U11782 (N_11782,N_10164,N_10447);
and U11783 (N_11783,N_10415,N_10720);
and U11784 (N_11784,N_10925,N_10402);
or U11785 (N_11785,N_10642,N_10589);
nor U11786 (N_11786,N_10525,N_10783);
nand U11787 (N_11787,N_10815,N_10804);
and U11788 (N_11788,N_10800,N_10830);
nand U11789 (N_11789,N_10589,N_10550);
nand U11790 (N_11790,N_10050,N_10410);
nor U11791 (N_11791,N_10624,N_10810);
and U11792 (N_11792,N_10732,N_10042);
or U11793 (N_11793,N_10131,N_10725);
or U11794 (N_11794,N_10109,N_10296);
nand U11795 (N_11795,N_10175,N_10230);
or U11796 (N_11796,N_10474,N_10436);
nor U11797 (N_11797,N_10227,N_10199);
nand U11798 (N_11798,N_10312,N_10636);
xor U11799 (N_11799,N_10490,N_10110);
and U11800 (N_11800,N_10166,N_10481);
and U11801 (N_11801,N_10904,N_10705);
nor U11802 (N_11802,N_10720,N_10493);
nor U11803 (N_11803,N_10544,N_10328);
nor U11804 (N_11804,N_10825,N_10657);
and U11805 (N_11805,N_10695,N_10162);
nor U11806 (N_11806,N_10736,N_10993);
or U11807 (N_11807,N_10438,N_10555);
nor U11808 (N_11808,N_10006,N_10335);
nor U11809 (N_11809,N_10755,N_10646);
xor U11810 (N_11810,N_10342,N_10491);
and U11811 (N_11811,N_10511,N_10048);
nand U11812 (N_11812,N_10196,N_10996);
xor U11813 (N_11813,N_10298,N_10985);
nor U11814 (N_11814,N_10161,N_10306);
and U11815 (N_11815,N_10303,N_10458);
nand U11816 (N_11816,N_10362,N_10300);
nand U11817 (N_11817,N_10431,N_10370);
nand U11818 (N_11818,N_10089,N_10367);
and U11819 (N_11819,N_10595,N_10895);
and U11820 (N_11820,N_10446,N_10689);
or U11821 (N_11821,N_10250,N_10526);
nand U11822 (N_11822,N_10015,N_10082);
or U11823 (N_11823,N_10077,N_10940);
or U11824 (N_11824,N_10490,N_10347);
or U11825 (N_11825,N_10629,N_10845);
and U11826 (N_11826,N_10237,N_10525);
xor U11827 (N_11827,N_10076,N_10605);
nor U11828 (N_11828,N_10896,N_10637);
nand U11829 (N_11829,N_10877,N_10991);
or U11830 (N_11830,N_10872,N_10199);
nand U11831 (N_11831,N_10024,N_10428);
nor U11832 (N_11832,N_10914,N_10565);
and U11833 (N_11833,N_10318,N_10915);
nor U11834 (N_11834,N_10585,N_10555);
nor U11835 (N_11835,N_10961,N_10031);
or U11836 (N_11836,N_10428,N_10849);
xor U11837 (N_11837,N_10945,N_10545);
nand U11838 (N_11838,N_10259,N_10665);
nand U11839 (N_11839,N_10484,N_10075);
nor U11840 (N_11840,N_10230,N_10438);
xor U11841 (N_11841,N_10643,N_10385);
nand U11842 (N_11842,N_10779,N_10627);
or U11843 (N_11843,N_10836,N_10343);
or U11844 (N_11844,N_10433,N_10384);
nor U11845 (N_11845,N_10389,N_10957);
or U11846 (N_11846,N_10639,N_10880);
nand U11847 (N_11847,N_10506,N_10873);
nor U11848 (N_11848,N_10604,N_10896);
nand U11849 (N_11849,N_10156,N_10759);
nand U11850 (N_11850,N_10795,N_10108);
and U11851 (N_11851,N_10245,N_10637);
nor U11852 (N_11852,N_10921,N_10423);
nor U11853 (N_11853,N_10466,N_10487);
or U11854 (N_11854,N_10711,N_10496);
or U11855 (N_11855,N_10522,N_10863);
nor U11856 (N_11856,N_10497,N_10142);
and U11857 (N_11857,N_10544,N_10988);
nand U11858 (N_11858,N_10605,N_10670);
nand U11859 (N_11859,N_10666,N_10724);
or U11860 (N_11860,N_10984,N_10292);
or U11861 (N_11861,N_10025,N_10907);
nor U11862 (N_11862,N_10207,N_10068);
or U11863 (N_11863,N_10518,N_10870);
xor U11864 (N_11864,N_10045,N_10238);
and U11865 (N_11865,N_10523,N_10130);
xnor U11866 (N_11866,N_10638,N_10948);
and U11867 (N_11867,N_10742,N_10217);
nor U11868 (N_11868,N_10873,N_10667);
or U11869 (N_11869,N_10076,N_10192);
xnor U11870 (N_11870,N_10204,N_10427);
or U11871 (N_11871,N_10412,N_10691);
nor U11872 (N_11872,N_10430,N_10259);
and U11873 (N_11873,N_10156,N_10437);
or U11874 (N_11874,N_10790,N_10421);
or U11875 (N_11875,N_10316,N_10615);
or U11876 (N_11876,N_10522,N_10438);
nor U11877 (N_11877,N_10945,N_10560);
xor U11878 (N_11878,N_10552,N_10673);
and U11879 (N_11879,N_10664,N_10053);
and U11880 (N_11880,N_10654,N_10741);
or U11881 (N_11881,N_10087,N_10591);
nor U11882 (N_11882,N_10375,N_10303);
or U11883 (N_11883,N_10218,N_10081);
and U11884 (N_11884,N_10540,N_10271);
xnor U11885 (N_11885,N_10322,N_10879);
xor U11886 (N_11886,N_10896,N_10535);
or U11887 (N_11887,N_10260,N_10131);
nand U11888 (N_11888,N_10034,N_10878);
nand U11889 (N_11889,N_10091,N_10714);
nand U11890 (N_11890,N_10741,N_10573);
or U11891 (N_11891,N_10359,N_10162);
nand U11892 (N_11892,N_10459,N_10687);
or U11893 (N_11893,N_10888,N_10154);
nand U11894 (N_11894,N_10947,N_10904);
or U11895 (N_11895,N_10223,N_10112);
nand U11896 (N_11896,N_10278,N_10090);
or U11897 (N_11897,N_10356,N_10623);
or U11898 (N_11898,N_10584,N_10867);
and U11899 (N_11899,N_10008,N_10590);
and U11900 (N_11900,N_10203,N_10438);
nor U11901 (N_11901,N_10916,N_10498);
xor U11902 (N_11902,N_10026,N_10723);
nand U11903 (N_11903,N_10945,N_10715);
nor U11904 (N_11904,N_10553,N_10189);
and U11905 (N_11905,N_10704,N_10243);
and U11906 (N_11906,N_10137,N_10682);
nand U11907 (N_11907,N_10490,N_10515);
nor U11908 (N_11908,N_10366,N_10518);
and U11909 (N_11909,N_10585,N_10501);
nand U11910 (N_11910,N_10612,N_10793);
and U11911 (N_11911,N_10617,N_10858);
nor U11912 (N_11912,N_10786,N_10250);
nand U11913 (N_11913,N_10629,N_10233);
xor U11914 (N_11914,N_10263,N_10306);
nand U11915 (N_11915,N_10872,N_10538);
or U11916 (N_11916,N_10351,N_10925);
nor U11917 (N_11917,N_10845,N_10953);
and U11918 (N_11918,N_10759,N_10495);
or U11919 (N_11919,N_10617,N_10056);
nand U11920 (N_11920,N_10005,N_10502);
xnor U11921 (N_11921,N_10042,N_10312);
nand U11922 (N_11922,N_10011,N_10593);
and U11923 (N_11923,N_10992,N_10749);
or U11924 (N_11924,N_10180,N_10600);
or U11925 (N_11925,N_10713,N_10744);
or U11926 (N_11926,N_10174,N_10814);
and U11927 (N_11927,N_10852,N_10011);
and U11928 (N_11928,N_10445,N_10860);
or U11929 (N_11929,N_10137,N_10652);
nand U11930 (N_11930,N_10043,N_10375);
and U11931 (N_11931,N_10638,N_10325);
nor U11932 (N_11932,N_10754,N_10130);
or U11933 (N_11933,N_10589,N_10960);
xnor U11934 (N_11934,N_10483,N_10331);
and U11935 (N_11935,N_10247,N_10248);
and U11936 (N_11936,N_10610,N_10160);
and U11937 (N_11937,N_10564,N_10716);
or U11938 (N_11938,N_10205,N_10701);
nor U11939 (N_11939,N_10552,N_10114);
and U11940 (N_11940,N_10424,N_10555);
nand U11941 (N_11941,N_10071,N_10801);
and U11942 (N_11942,N_10299,N_10245);
or U11943 (N_11943,N_10718,N_10088);
and U11944 (N_11944,N_10259,N_10352);
nand U11945 (N_11945,N_10796,N_10811);
nand U11946 (N_11946,N_10402,N_10997);
nor U11947 (N_11947,N_10174,N_10759);
nor U11948 (N_11948,N_10838,N_10498);
or U11949 (N_11949,N_10617,N_10340);
nor U11950 (N_11950,N_10710,N_10295);
nand U11951 (N_11951,N_10490,N_10087);
nand U11952 (N_11952,N_10932,N_10372);
nand U11953 (N_11953,N_10130,N_10239);
and U11954 (N_11954,N_10344,N_10110);
nand U11955 (N_11955,N_10072,N_10388);
nand U11956 (N_11956,N_10501,N_10586);
nand U11957 (N_11957,N_10005,N_10151);
or U11958 (N_11958,N_10754,N_10935);
or U11959 (N_11959,N_10367,N_10792);
nand U11960 (N_11960,N_10185,N_10553);
or U11961 (N_11961,N_10112,N_10405);
and U11962 (N_11962,N_10347,N_10789);
nor U11963 (N_11963,N_10694,N_10251);
or U11964 (N_11964,N_10385,N_10257);
or U11965 (N_11965,N_10755,N_10404);
nor U11966 (N_11966,N_10639,N_10993);
nor U11967 (N_11967,N_10992,N_10580);
and U11968 (N_11968,N_10222,N_10437);
xnor U11969 (N_11969,N_10862,N_10728);
nor U11970 (N_11970,N_10584,N_10720);
xor U11971 (N_11971,N_10609,N_10630);
or U11972 (N_11972,N_10418,N_10325);
nand U11973 (N_11973,N_10631,N_10806);
and U11974 (N_11974,N_10536,N_10330);
or U11975 (N_11975,N_10236,N_10649);
nor U11976 (N_11976,N_10291,N_10406);
xor U11977 (N_11977,N_10899,N_10475);
or U11978 (N_11978,N_10960,N_10625);
nor U11979 (N_11979,N_10180,N_10641);
or U11980 (N_11980,N_10311,N_10834);
and U11981 (N_11981,N_10025,N_10430);
nand U11982 (N_11982,N_10074,N_10080);
nor U11983 (N_11983,N_10284,N_10437);
nand U11984 (N_11984,N_10725,N_10067);
nor U11985 (N_11985,N_10637,N_10640);
or U11986 (N_11986,N_10864,N_10659);
or U11987 (N_11987,N_10983,N_10293);
nand U11988 (N_11988,N_10598,N_10728);
nor U11989 (N_11989,N_10863,N_10843);
and U11990 (N_11990,N_10737,N_10815);
nor U11991 (N_11991,N_10805,N_10418);
or U11992 (N_11992,N_10016,N_10400);
nand U11993 (N_11993,N_10980,N_10518);
or U11994 (N_11994,N_10862,N_10708);
and U11995 (N_11995,N_10860,N_10414);
nor U11996 (N_11996,N_10636,N_10409);
nand U11997 (N_11997,N_10228,N_10578);
nor U11998 (N_11998,N_10141,N_10083);
nand U11999 (N_11999,N_10011,N_10687);
nand U12000 (N_12000,N_11328,N_11780);
or U12001 (N_12001,N_11673,N_11297);
and U12002 (N_12002,N_11921,N_11934);
nor U12003 (N_12003,N_11338,N_11126);
nor U12004 (N_12004,N_11665,N_11103);
or U12005 (N_12005,N_11269,N_11987);
or U12006 (N_12006,N_11979,N_11664);
or U12007 (N_12007,N_11282,N_11090);
nand U12008 (N_12008,N_11005,N_11607);
or U12009 (N_12009,N_11738,N_11332);
nand U12010 (N_12010,N_11339,N_11751);
and U12011 (N_12011,N_11764,N_11550);
and U12012 (N_12012,N_11777,N_11937);
or U12013 (N_12013,N_11346,N_11027);
nor U12014 (N_12014,N_11374,N_11417);
xnor U12015 (N_12015,N_11713,N_11152);
nand U12016 (N_12016,N_11265,N_11067);
nand U12017 (N_12017,N_11766,N_11678);
nand U12018 (N_12018,N_11836,N_11118);
xor U12019 (N_12019,N_11365,N_11641);
nand U12020 (N_12020,N_11014,N_11349);
nand U12021 (N_12021,N_11096,N_11649);
and U12022 (N_12022,N_11476,N_11320);
and U12023 (N_12023,N_11444,N_11393);
xnor U12024 (N_12024,N_11864,N_11489);
nor U12025 (N_12025,N_11988,N_11160);
nor U12026 (N_12026,N_11286,N_11547);
nand U12027 (N_12027,N_11405,N_11782);
nor U12028 (N_12028,N_11735,N_11565);
nand U12029 (N_12029,N_11443,N_11380);
nand U12030 (N_12030,N_11151,N_11206);
or U12031 (N_12031,N_11769,N_11926);
and U12032 (N_12032,N_11885,N_11425);
nor U12033 (N_12033,N_11671,N_11133);
nand U12034 (N_12034,N_11331,N_11079);
xor U12035 (N_12035,N_11931,N_11849);
or U12036 (N_12036,N_11288,N_11431);
xnor U12037 (N_12037,N_11589,N_11889);
and U12038 (N_12038,N_11150,N_11855);
nand U12039 (N_12039,N_11870,N_11852);
nor U12040 (N_12040,N_11064,N_11483);
nand U12041 (N_12041,N_11705,N_11469);
or U12042 (N_12042,N_11826,N_11451);
nor U12043 (N_12043,N_11539,N_11490);
nor U12044 (N_12044,N_11504,N_11778);
or U12045 (N_12045,N_11413,N_11841);
or U12046 (N_12046,N_11553,N_11364);
and U12047 (N_12047,N_11527,N_11801);
and U12048 (N_12048,N_11971,N_11440);
nand U12049 (N_12049,N_11403,N_11189);
or U12050 (N_12050,N_11045,N_11868);
xor U12051 (N_12051,N_11268,N_11129);
and U12052 (N_12052,N_11397,N_11519);
nand U12053 (N_12053,N_11991,N_11740);
xor U12054 (N_12054,N_11244,N_11406);
and U12055 (N_12055,N_11140,N_11367);
or U12056 (N_12056,N_11372,N_11568);
or U12057 (N_12057,N_11668,N_11585);
and U12058 (N_12058,N_11570,N_11640);
nor U12059 (N_12059,N_11691,N_11376);
nand U12060 (N_12060,N_11977,N_11128);
or U12061 (N_12061,N_11960,N_11871);
nand U12062 (N_12062,N_11312,N_11694);
nand U12063 (N_12063,N_11322,N_11314);
nand U12064 (N_12064,N_11121,N_11615);
nor U12065 (N_12065,N_11588,N_11993);
nand U12066 (N_12066,N_11882,N_11813);
or U12067 (N_12067,N_11806,N_11952);
and U12068 (N_12068,N_11420,N_11051);
xnor U12069 (N_12069,N_11373,N_11355);
and U12070 (N_12070,N_11422,N_11911);
nor U12071 (N_12071,N_11449,N_11283);
nor U12072 (N_12072,N_11060,N_11513);
xnor U12073 (N_12073,N_11935,N_11226);
and U12074 (N_12074,N_11657,N_11784);
nor U12075 (N_12075,N_11234,N_11028);
and U12076 (N_12076,N_11454,N_11273);
and U12077 (N_12077,N_11672,N_11566);
or U12078 (N_12078,N_11591,N_11158);
nand U12079 (N_12079,N_11390,N_11618);
or U12080 (N_12080,N_11517,N_11626);
or U12081 (N_12081,N_11492,N_11468);
and U12082 (N_12082,N_11084,N_11962);
nand U12083 (N_12083,N_11613,N_11630);
and U12084 (N_12084,N_11295,N_11036);
or U12085 (N_12085,N_11486,N_11088);
and U12086 (N_12086,N_11395,N_11202);
nor U12087 (N_12087,N_11131,N_11767);
or U12088 (N_12088,N_11956,N_11359);
nand U12089 (N_12089,N_11856,N_11388);
nand U12090 (N_12090,N_11939,N_11839);
nor U12091 (N_12091,N_11765,N_11307);
and U12092 (N_12092,N_11019,N_11007);
nor U12093 (N_12093,N_11501,N_11333);
xor U12094 (N_12094,N_11964,N_11974);
and U12095 (N_12095,N_11018,N_11185);
xor U12096 (N_12096,N_11894,N_11632);
and U12097 (N_12097,N_11854,N_11434);
nor U12098 (N_12098,N_11238,N_11032);
or U12099 (N_12099,N_11267,N_11512);
nand U12100 (N_12100,N_11879,N_11230);
or U12101 (N_12101,N_11368,N_11264);
and U12102 (N_12102,N_11802,N_11191);
and U12103 (N_12103,N_11003,N_11736);
and U12104 (N_12104,N_11195,N_11592);
nand U12105 (N_12105,N_11464,N_11946);
nor U12106 (N_12106,N_11670,N_11199);
nor U12107 (N_12107,N_11627,N_11085);
and U12108 (N_12108,N_11033,N_11201);
xnor U12109 (N_12109,N_11594,N_11772);
or U12110 (N_12110,N_11680,N_11139);
and U12111 (N_12111,N_11272,N_11159);
or U12112 (N_12112,N_11633,N_11990);
and U12113 (N_12113,N_11052,N_11537);
nor U12114 (N_12114,N_11162,N_11276);
xor U12115 (N_12115,N_11254,N_11345);
and U12116 (N_12116,N_11203,N_11301);
and U12117 (N_12117,N_11429,N_11781);
nand U12118 (N_12118,N_11721,N_11351);
nor U12119 (N_12119,N_11916,N_11034);
nand U12120 (N_12120,N_11194,N_11240);
and U12121 (N_12121,N_11072,N_11334);
and U12122 (N_12122,N_11091,N_11969);
and U12123 (N_12123,N_11893,N_11498);
and U12124 (N_12124,N_11681,N_11843);
nor U12125 (N_12125,N_11912,N_11795);
and U12126 (N_12126,N_11810,N_11366);
nand U12127 (N_12127,N_11614,N_11847);
and U12128 (N_12128,N_11989,N_11107);
and U12129 (N_12129,N_11686,N_11207);
nand U12130 (N_12130,N_11722,N_11447);
xor U12131 (N_12131,N_11883,N_11002);
xor U12132 (N_12132,N_11808,N_11508);
xnor U12133 (N_12133,N_11462,N_11621);
and U12134 (N_12134,N_11009,N_11563);
nand U12135 (N_12135,N_11510,N_11947);
or U12136 (N_12136,N_11506,N_11166);
and U12137 (N_12137,N_11940,N_11190);
nor U12138 (N_12138,N_11699,N_11726);
and U12139 (N_12139,N_11433,N_11361);
nand U12140 (N_12140,N_11915,N_11284);
or U12141 (N_12141,N_11082,N_11574);
xor U12142 (N_12142,N_11904,N_11482);
nor U12143 (N_12143,N_11992,N_11610);
nand U12144 (N_12144,N_11905,N_11292);
nand U12145 (N_12145,N_11712,N_11541);
and U12146 (N_12146,N_11768,N_11436);
and U12147 (N_12147,N_11493,N_11456);
or U12148 (N_12148,N_11676,N_11573);
and U12149 (N_12149,N_11168,N_11996);
nor U12150 (N_12150,N_11500,N_11628);
xnor U12151 (N_12151,N_11774,N_11289);
and U12152 (N_12152,N_11783,N_11310);
nor U12153 (N_12153,N_11677,N_11816);
xnor U12154 (N_12154,N_11844,N_11799);
nand U12155 (N_12155,N_11529,N_11938);
nor U12156 (N_12156,N_11688,N_11685);
and U12157 (N_12157,N_11706,N_11170);
nor U12158 (N_12158,N_11695,N_11171);
xnor U12159 (N_12159,N_11581,N_11119);
nand U12160 (N_12160,N_11344,N_11907);
nor U12161 (N_12161,N_11210,N_11898);
nand U12162 (N_12162,N_11277,N_11930);
nand U12163 (N_12163,N_11176,N_11184);
and U12164 (N_12164,N_11270,N_11467);
xnor U12165 (N_12165,N_11579,N_11619);
nand U12166 (N_12166,N_11378,N_11950);
or U12167 (N_12167,N_11427,N_11475);
or U12168 (N_12168,N_11723,N_11817);
nor U12169 (N_12169,N_11488,N_11616);
or U12170 (N_12170,N_11995,N_11976);
nand U12171 (N_12171,N_11561,N_11667);
and U12172 (N_12172,N_11154,N_11653);
nor U12173 (N_12173,N_11421,N_11652);
nand U12174 (N_12174,N_11714,N_11731);
nand U12175 (N_12175,N_11143,N_11701);
nand U12176 (N_12176,N_11304,N_11635);
xor U12177 (N_12177,N_11900,N_11381);
nor U12178 (N_12178,N_11326,N_11290);
and U12179 (N_12179,N_11875,N_11941);
or U12180 (N_12180,N_11316,N_11329);
nand U12181 (N_12181,N_11880,N_11183);
nand U12182 (N_12182,N_11258,N_11169);
and U12183 (N_12183,N_11865,N_11318);
nor U12184 (N_12184,N_11822,N_11148);
and U12185 (N_12185,N_11384,N_11697);
and U12186 (N_12186,N_11982,N_11303);
or U12187 (N_12187,N_11038,N_11655);
and U12188 (N_12188,N_11061,N_11845);
and U12189 (N_12189,N_11944,N_11984);
nand U12190 (N_12190,N_11216,N_11580);
xor U12191 (N_12191,N_11549,N_11457);
or U12192 (N_12192,N_11967,N_11229);
or U12193 (N_12193,N_11347,N_11021);
nor U12194 (N_12194,N_11639,N_11544);
and U12195 (N_12195,N_11603,N_11902);
xor U12196 (N_12196,N_11400,N_11980);
and U12197 (N_12197,N_11656,N_11629);
and U12198 (N_12198,N_11037,N_11704);
and U12199 (N_12199,N_11016,N_11411);
and U12200 (N_12200,N_11961,N_11948);
nand U12201 (N_12201,N_11227,N_11505);
or U12202 (N_12202,N_11149,N_11077);
nand U12203 (N_12203,N_11105,N_11584);
or U12204 (N_12204,N_11602,N_11070);
and U12205 (N_12205,N_11918,N_11192);
nor U12206 (N_12206,N_11785,N_11658);
and U12207 (N_12207,N_11514,N_11287);
or U12208 (N_12208,N_11903,N_11834);
and U12209 (N_12209,N_11050,N_11000);
and U12210 (N_12210,N_11908,N_11398);
nand U12211 (N_12211,N_11410,N_11873);
nand U12212 (N_12212,N_11246,N_11773);
and U12213 (N_12213,N_11545,N_11293);
and U12214 (N_12214,N_11430,N_11642);
nor U12215 (N_12215,N_11354,N_11963);
nand U12216 (N_12216,N_11362,N_11625);
or U12217 (N_12217,N_11259,N_11385);
or U12218 (N_12218,N_11336,N_11881);
nor U12219 (N_12219,N_11858,N_11127);
nor U12220 (N_12220,N_11474,N_11074);
nor U12221 (N_12221,N_11920,N_11583);
nand U12222 (N_12222,N_11942,N_11555);
nor U12223 (N_12223,N_11306,N_11375);
nor U12224 (N_12224,N_11919,N_11484);
or U12225 (N_12225,N_11308,N_11526);
and U12226 (N_12226,N_11675,N_11648);
xnor U12227 (N_12227,N_11460,N_11222);
nor U12228 (N_12228,N_11524,N_11231);
nor U12229 (N_12229,N_11205,N_11132);
nand U12230 (N_12230,N_11554,N_11687);
or U12231 (N_12231,N_11728,N_11142);
xor U12232 (N_12232,N_11453,N_11771);
nand U12233 (N_12233,N_11209,N_11204);
nor U12234 (N_12234,N_11059,N_11624);
nand U12235 (N_12235,N_11383,N_11369);
and U12236 (N_12236,N_11445,N_11901);
nand U12237 (N_12237,N_11487,N_11634);
or U12238 (N_12238,N_11812,N_11465);
nand U12239 (N_12239,N_11718,N_11927);
xnor U12240 (N_12240,N_11178,N_11754);
xnor U12241 (N_12241,N_11761,N_11008);
nor U12242 (N_12242,N_11913,N_11720);
nor U12243 (N_12243,N_11636,N_11896);
nand U12244 (N_12244,N_11011,N_11805);
nand U12245 (N_12245,N_11266,N_11788);
and U12246 (N_12246,N_11075,N_11387);
and U12247 (N_12247,N_11887,N_11606);
and U12248 (N_12248,N_11787,N_11975);
and U12249 (N_12249,N_11859,N_11605);
nor U12250 (N_12250,N_11237,N_11224);
nand U12251 (N_12251,N_11315,N_11569);
and U12252 (N_12252,N_11054,N_11832);
nor U12253 (N_12253,N_11041,N_11057);
nand U12254 (N_12254,N_11571,N_11679);
nand U12255 (N_12255,N_11559,N_11323);
nor U12256 (N_12256,N_11186,N_11876);
and U12257 (N_12257,N_11660,N_11543);
nor U12258 (N_12258,N_11596,N_11144);
and U12259 (N_12259,N_11730,N_11407);
or U12260 (N_12260,N_11120,N_11593);
or U12261 (N_12261,N_11340,N_11111);
nand U12262 (N_12262,N_11049,N_11156);
nor U12263 (N_12263,N_11485,N_11756);
or U12264 (N_12264,N_11208,N_11622);
nor U12265 (N_12265,N_11114,N_11495);
and U12266 (N_12266,N_11071,N_11848);
nand U12267 (N_12267,N_11755,N_11217);
xor U12268 (N_12268,N_11760,N_11092);
xnor U12269 (N_12269,N_11179,N_11983);
nor U12270 (N_12270,N_11062,N_11827);
or U12271 (N_12271,N_11707,N_11327);
or U12272 (N_12272,N_11775,N_11167);
nand U12273 (N_12273,N_11572,N_11542);
nand U12274 (N_12274,N_11753,N_11352);
and U12275 (N_12275,N_11499,N_11392);
and U12276 (N_12276,N_11609,N_11026);
nand U12277 (N_12277,N_11598,N_11225);
or U12278 (N_12278,N_11762,N_11862);
and U12279 (N_12279,N_11533,N_11748);
and U12280 (N_12280,N_11099,N_11214);
nand U12281 (N_12281,N_11412,N_11708);
nand U12282 (N_12282,N_11389,N_11432);
nand U12283 (N_12283,N_11115,N_11164);
nor U12284 (N_12284,N_11325,N_11530);
or U12285 (N_12285,N_11558,N_11418);
and U12286 (N_12286,N_11155,N_11604);
or U12287 (N_12287,N_11525,N_11069);
nand U12288 (N_12288,N_11219,N_11145);
and U12289 (N_12289,N_11239,N_11507);
or U12290 (N_12290,N_11047,N_11313);
or U12291 (N_12291,N_11892,N_11577);
nand U12292 (N_12292,N_11698,N_11663);
or U12293 (N_12293,N_11895,N_11260);
and U12294 (N_12294,N_11452,N_11044);
or U12295 (N_12295,N_11319,N_11350);
nand U12296 (N_12296,N_11953,N_11025);
xnor U12297 (N_12297,N_11818,N_11102);
and U12298 (N_12298,N_11046,N_11824);
and U12299 (N_12299,N_11248,N_11015);
nor U12300 (N_12300,N_11497,N_11343);
and U12301 (N_12301,N_11776,N_11874);
or U12302 (N_12302,N_11846,N_11620);
and U12303 (N_12303,N_11104,N_11357);
nor U12304 (N_12304,N_11794,N_11035);
nor U12305 (N_12305,N_11548,N_11100);
and U12306 (N_12306,N_11157,N_11857);
and U12307 (N_12307,N_11448,N_11779);
or U12308 (N_12308,N_11884,N_11494);
and U12309 (N_12309,N_11094,N_11236);
and U12310 (N_12310,N_11043,N_11068);
nand U12311 (N_12311,N_11564,N_11757);
or U12312 (N_12312,N_11985,N_11394);
or U12313 (N_12313,N_11480,N_11745);
nor U12314 (N_12314,N_11263,N_11710);
and U12315 (N_12315,N_11851,N_11823);
nor U12316 (N_12316,N_11978,N_11409);
and U12317 (N_12317,N_11644,N_11481);
xor U12318 (N_12318,N_11163,N_11321);
and U12319 (N_12319,N_11382,N_11053);
and U12320 (N_12320,N_11479,N_11280);
or U12321 (N_12321,N_11838,N_11386);
or U12322 (N_12322,N_11377,N_11623);
and U12323 (N_12323,N_11285,N_11943);
nor U12324 (N_12324,N_11994,N_11211);
xor U12325 (N_12325,N_11973,N_11419);
nand U12326 (N_12326,N_11279,N_11257);
xor U12327 (N_12327,N_11599,N_11968);
nor U12328 (N_12328,N_11408,N_11428);
and U12329 (N_12329,N_11337,N_11123);
nor U12330 (N_12330,N_11249,N_11029);
and U12331 (N_12331,N_11715,N_11175);
nand U12332 (N_12332,N_11693,N_11466);
nor U12333 (N_12333,N_11305,N_11717);
nor U12334 (N_12334,N_11039,N_11897);
or U12335 (N_12335,N_11017,N_11470);
and U12336 (N_12336,N_11954,N_11491);
nor U12337 (N_12337,N_11786,N_11198);
or U12338 (N_12338,N_11423,N_11330);
nand U12339 (N_12339,N_11098,N_11741);
nand U12340 (N_12340,N_11750,N_11117);
or U12341 (N_12341,N_11030,N_11278);
nor U12342 (N_12342,N_11651,N_11650);
or U12343 (N_12343,N_11890,N_11733);
nand U12344 (N_12344,N_11010,N_11252);
nand U12345 (N_12345,N_11137,N_11924);
nor U12346 (N_12346,N_11110,N_11752);
nor U12347 (N_12347,N_11909,N_11055);
and U12348 (N_12348,N_11804,N_11957);
and U12349 (N_12349,N_11809,N_11116);
and U12350 (N_12350,N_11821,N_11274);
nor U12351 (N_12351,N_11877,N_11637);
or U12352 (N_12352,N_11560,N_11540);
nor U12353 (N_12353,N_11177,N_11684);
and U12354 (N_12354,N_11065,N_11661);
nor U12355 (N_12355,N_11473,N_11441);
or U12356 (N_12356,N_11811,N_11477);
and U12357 (N_12357,N_11013,N_11595);
xor U12358 (N_12358,N_11134,N_11125);
xor U12359 (N_12359,N_11578,N_11188);
nand U12360 (N_12360,N_11792,N_11562);
nand U12361 (N_12361,N_11122,N_11551);
and U12362 (N_12362,N_11820,N_11643);
and U12363 (N_12363,N_11414,N_11590);
nor U12364 (N_12364,N_11081,N_11582);
nand U12365 (N_12365,N_11600,N_11972);
or U12366 (N_12366,N_11702,N_11024);
xnor U12367 (N_12367,N_11829,N_11317);
nand U12368 (N_12368,N_11022,N_11997);
nor U12369 (N_12369,N_11749,N_11727);
nor U12370 (N_12370,N_11415,N_11136);
nor U12371 (N_12371,N_11097,N_11796);
or U12372 (N_12372,N_11797,N_11180);
and U12373 (N_12373,N_11575,N_11763);
and U12374 (N_12374,N_11471,N_11342);
and U12375 (N_12375,N_11669,N_11732);
nor U12376 (N_12376,N_11725,N_11531);
nand U12377 (N_12377,N_11233,N_11215);
or U12378 (N_12378,N_11523,N_11970);
and U12379 (N_12379,N_11770,N_11638);
or U12380 (N_12380,N_11302,N_11012);
nor U12381 (N_12381,N_11245,N_11791);
nand U12382 (N_12382,N_11965,N_11608);
xnor U12383 (N_12383,N_11212,N_11866);
or U12384 (N_12384,N_11746,N_11353);
and U12385 (N_12385,N_11251,N_11793);
nand U12386 (N_12386,N_11161,N_11682);
nand U12387 (N_12387,N_11891,N_11446);
and U12388 (N_12388,N_11951,N_11299);
or U12389 (N_12389,N_11986,N_11744);
and U12390 (N_12390,N_11173,N_11703);
or U12391 (N_12391,N_11556,N_11348);
xnor U12392 (N_12392,N_11089,N_11709);
and U12393 (N_12393,N_11869,N_11020);
nor U12394 (N_12394,N_11528,N_11416);
xnor U12395 (N_12395,N_11910,N_11509);
xor U12396 (N_12396,N_11261,N_11929);
nand U12397 (N_12397,N_11193,N_11576);
or U12398 (N_12398,N_11108,N_11478);
and U12399 (N_12399,N_11358,N_11631);
nand U12400 (N_12400,N_11789,N_11458);
xor U12401 (N_12401,N_11496,N_11196);
xor U12402 (N_12402,N_11141,N_11396);
xor U12403 (N_12403,N_11932,N_11101);
nor U12404 (N_12404,N_11700,N_11999);
and U12405 (N_12405,N_11031,N_11001);
or U12406 (N_12406,N_11850,N_11521);
nand U12407 (N_12407,N_11803,N_11516);
nand U12408 (N_12408,N_11724,N_11674);
xnor U12409 (N_12409,N_11587,N_11719);
and U12410 (N_12410,N_11404,N_11438);
nand U12411 (N_12411,N_11742,N_11109);
nand U12412 (N_12412,N_11511,N_11955);
nor U12413 (N_12413,N_11356,N_11959);
nor U12414 (N_12414,N_11842,N_11831);
nand U12415 (N_12415,N_11567,N_11853);
and U12416 (N_12416,N_11004,N_11172);
nand U12417 (N_12417,N_11689,N_11518);
nand U12418 (N_12418,N_11040,N_11335);
and U12419 (N_12419,N_11546,N_11439);
or U12420 (N_12420,N_11860,N_11341);
nand U12421 (N_12421,N_11253,N_11223);
xor U12422 (N_12422,N_11917,N_11213);
and U12423 (N_12423,N_11981,N_11886);
nand U12424 (N_12424,N_11232,N_11300);
and U12425 (N_12425,N_11086,N_11243);
or U12426 (N_12426,N_11683,N_11147);
or U12427 (N_12427,N_11645,N_11242);
and U12428 (N_12428,N_11165,N_11535);
xnor U12429 (N_12429,N_11463,N_11124);
nor U12430 (N_12430,N_11833,N_11363);
and U12431 (N_12431,N_11692,N_11455);
or U12432 (N_12432,N_11747,N_11058);
and U12433 (N_12433,N_11459,N_11153);
and U12434 (N_12434,N_11611,N_11424);
nand U12435 (N_12435,N_11042,N_11174);
or U12436 (N_12436,N_11729,N_11922);
nand U12437 (N_12437,N_11146,N_11534);
nand U12438 (N_12438,N_11662,N_11867);
or U12439 (N_12439,N_11023,N_11840);
or U12440 (N_12440,N_11371,N_11532);
nand U12441 (N_12441,N_11138,N_11666);
and U12442 (N_12442,N_11612,N_11503);
or U12443 (N_12443,N_11958,N_11250);
xnor U12444 (N_12444,N_11281,N_11262);
nor U12445 (N_12445,N_11743,N_11401);
and U12446 (N_12446,N_11048,N_11197);
xor U12447 (N_12447,N_11914,N_11221);
or U12448 (N_12448,N_11112,N_11899);
and U12449 (N_12449,N_11472,N_11402);
and U12450 (N_12450,N_11379,N_11716);
nor U12451 (N_12451,N_11814,N_11586);
xnor U12452 (N_12452,N_11056,N_11998);
or U12453 (N_12453,N_11063,N_11888);
and U12454 (N_12454,N_11399,N_11135);
and U12455 (N_12455,N_11828,N_11552);
xnor U12456 (N_12456,N_11837,N_11557);
or U12457 (N_12457,N_11181,N_11087);
or U12458 (N_12458,N_11872,N_11275);
and U12459 (N_12459,N_11095,N_11923);
nor U12460 (N_12460,N_11255,N_11437);
and U12461 (N_12461,N_11187,N_11966);
or U12462 (N_12462,N_11235,N_11835);
nand U12463 (N_12463,N_11928,N_11442);
and U12464 (N_12464,N_11739,N_11790);
or U12465 (N_12465,N_11861,N_11654);
and U12466 (N_12466,N_11228,N_11311);
nand U12467 (N_12467,N_11093,N_11291);
nor U12468 (N_12468,N_11646,N_11461);
nand U12469 (N_12469,N_11825,N_11130);
nand U12470 (N_12470,N_11106,N_11659);
nand U12471 (N_12471,N_11271,N_11690);
nor U12472 (N_12472,N_11597,N_11080);
nand U12473 (N_12473,N_11113,N_11758);
nand U12474 (N_12474,N_11878,N_11296);
nand U12475 (N_12475,N_11256,N_11536);
or U12476 (N_12476,N_11078,N_11734);
xor U12477 (N_12477,N_11538,N_11696);
nor U12478 (N_12478,N_11182,N_11073);
or U12479 (N_12479,N_11798,N_11435);
and U12480 (N_12480,N_11925,N_11391);
xor U12481 (N_12481,N_11647,N_11759);
or U12482 (N_12482,N_11220,N_11241);
and U12483 (N_12483,N_11815,N_11502);
or U12484 (N_12484,N_11936,N_11426);
or U12485 (N_12485,N_11298,N_11520);
nor U12486 (N_12486,N_11515,N_11006);
nor U12487 (N_12487,N_11370,N_11906);
xor U12488 (N_12488,N_11076,N_11450);
and U12489 (N_12489,N_11294,N_11949);
and U12490 (N_12490,N_11863,N_11360);
and U12491 (N_12491,N_11324,N_11830);
and U12492 (N_12492,N_11711,N_11247);
and U12493 (N_12493,N_11522,N_11737);
nand U12494 (N_12494,N_11066,N_11218);
or U12495 (N_12495,N_11601,N_11800);
nand U12496 (N_12496,N_11617,N_11083);
or U12497 (N_12497,N_11945,N_11819);
nand U12498 (N_12498,N_11200,N_11807);
nor U12499 (N_12499,N_11933,N_11309);
nor U12500 (N_12500,N_11673,N_11441);
nor U12501 (N_12501,N_11461,N_11208);
or U12502 (N_12502,N_11661,N_11759);
nand U12503 (N_12503,N_11524,N_11152);
nand U12504 (N_12504,N_11750,N_11100);
nor U12505 (N_12505,N_11127,N_11114);
nand U12506 (N_12506,N_11087,N_11512);
and U12507 (N_12507,N_11286,N_11128);
or U12508 (N_12508,N_11882,N_11578);
or U12509 (N_12509,N_11918,N_11797);
or U12510 (N_12510,N_11999,N_11085);
nor U12511 (N_12511,N_11790,N_11134);
or U12512 (N_12512,N_11528,N_11802);
nor U12513 (N_12513,N_11283,N_11509);
nor U12514 (N_12514,N_11460,N_11112);
nand U12515 (N_12515,N_11400,N_11753);
or U12516 (N_12516,N_11764,N_11236);
nand U12517 (N_12517,N_11097,N_11856);
and U12518 (N_12518,N_11123,N_11653);
nand U12519 (N_12519,N_11272,N_11930);
or U12520 (N_12520,N_11859,N_11234);
or U12521 (N_12521,N_11011,N_11660);
and U12522 (N_12522,N_11618,N_11831);
and U12523 (N_12523,N_11341,N_11229);
and U12524 (N_12524,N_11461,N_11123);
or U12525 (N_12525,N_11468,N_11821);
nor U12526 (N_12526,N_11093,N_11394);
nand U12527 (N_12527,N_11729,N_11391);
nor U12528 (N_12528,N_11917,N_11821);
nor U12529 (N_12529,N_11087,N_11049);
nor U12530 (N_12530,N_11800,N_11128);
nor U12531 (N_12531,N_11559,N_11051);
and U12532 (N_12532,N_11901,N_11208);
nor U12533 (N_12533,N_11850,N_11634);
or U12534 (N_12534,N_11973,N_11360);
or U12535 (N_12535,N_11017,N_11647);
nor U12536 (N_12536,N_11957,N_11215);
or U12537 (N_12537,N_11599,N_11531);
nor U12538 (N_12538,N_11710,N_11821);
nand U12539 (N_12539,N_11856,N_11281);
nor U12540 (N_12540,N_11542,N_11989);
nor U12541 (N_12541,N_11480,N_11768);
and U12542 (N_12542,N_11054,N_11621);
nand U12543 (N_12543,N_11208,N_11937);
nand U12544 (N_12544,N_11391,N_11762);
and U12545 (N_12545,N_11978,N_11227);
nor U12546 (N_12546,N_11102,N_11678);
and U12547 (N_12547,N_11042,N_11764);
or U12548 (N_12548,N_11303,N_11686);
nor U12549 (N_12549,N_11895,N_11729);
nor U12550 (N_12550,N_11987,N_11730);
xor U12551 (N_12551,N_11322,N_11599);
nand U12552 (N_12552,N_11104,N_11335);
nor U12553 (N_12553,N_11266,N_11322);
nand U12554 (N_12554,N_11319,N_11191);
and U12555 (N_12555,N_11843,N_11140);
nand U12556 (N_12556,N_11880,N_11585);
nor U12557 (N_12557,N_11437,N_11429);
and U12558 (N_12558,N_11927,N_11942);
nand U12559 (N_12559,N_11860,N_11026);
nand U12560 (N_12560,N_11924,N_11868);
nor U12561 (N_12561,N_11710,N_11542);
nor U12562 (N_12562,N_11167,N_11908);
nor U12563 (N_12563,N_11963,N_11546);
xnor U12564 (N_12564,N_11024,N_11880);
xor U12565 (N_12565,N_11556,N_11043);
nand U12566 (N_12566,N_11479,N_11715);
nand U12567 (N_12567,N_11472,N_11978);
nor U12568 (N_12568,N_11372,N_11270);
nand U12569 (N_12569,N_11731,N_11955);
nor U12570 (N_12570,N_11096,N_11456);
and U12571 (N_12571,N_11938,N_11759);
or U12572 (N_12572,N_11867,N_11887);
nand U12573 (N_12573,N_11177,N_11595);
nor U12574 (N_12574,N_11620,N_11136);
and U12575 (N_12575,N_11316,N_11153);
nor U12576 (N_12576,N_11475,N_11321);
and U12577 (N_12577,N_11840,N_11161);
and U12578 (N_12578,N_11338,N_11134);
or U12579 (N_12579,N_11564,N_11813);
or U12580 (N_12580,N_11364,N_11166);
nor U12581 (N_12581,N_11148,N_11673);
nand U12582 (N_12582,N_11314,N_11692);
nand U12583 (N_12583,N_11598,N_11975);
nand U12584 (N_12584,N_11179,N_11252);
nor U12585 (N_12585,N_11327,N_11572);
or U12586 (N_12586,N_11620,N_11842);
nor U12587 (N_12587,N_11413,N_11761);
or U12588 (N_12588,N_11089,N_11773);
and U12589 (N_12589,N_11819,N_11693);
nor U12590 (N_12590,N_11677,N_11122);
nand U12591 (N_12591,N_11569,N_11441);
or U12592 (N_12592,N_11875,N_11380);
and U12593 (N_12593,N_11410,N_11580);
or U12594 (N_12594,N_11931,N_11188);
or U12595 (N_12595,N_11196,N_11769);
nor U12596 (N_12596,N_11773,N_11459);
nand U12597 (N_12597,N_11065,N_11950);
and U12598 (N_12598,N_11472,N_11924);
xnor U12599 (N_12599,N_11388,N_11061);
and U12600 (N_12600,N_11142,N_11801);
or U12601 (N_12601,N_11126,N_11887);
and U12602 (N_12602,N_11584,N_11036);
or U12603 (N_12603,N_11373,N_11316);
and U12604 (N_12604,N_11653,N_11147);
nor U12605 (N_12605,N_11724,N_11895);
nor U12606 (N_12606,N_11277,N_11521);
nor U12607 (N_12607,N_11248,N_11308);
and U12608 (N_12608,N_11101,N_11483);
or U12609 (N_12609,N_11002,N_11574);
xnor U12610 (N_12610,N_11823,N_11229);
and U12611 (N_12611,N_11259,N_11632);
nand U12612 (N_12612,N_11339,N_11258);
nor U12613 (N_12613,N_11796,N_11061);
or U12614 (N_12614,N_11415,N_11587);
xor U12615 (N_12615,N_11594,N_11052);
nor U12616 (N_12616,N_11097,N_11539);
or U12617 (N_12617,N_11823,N_11160);
nand U12618 (N_12618,N_11999,N_11638);
nand U12619 (N_12619,N_11406,N_11885);
nand U12620 (N_12620,N_11250,N_11609);
nor U12621 (N_12621,N_11831,N_11615);
or U12622 (N_12622,N_11669,N_11439);
nand U12623 (N_12623,N_11922,N_11945);
or U12624 (N_12624,N_11279,N_11903);
nor U12625 (N_12625,N_11183,N_11258);
and U12626 (N_12626,N_11841,N_11808);
and U12627 (N_12627,N_11915,N_11098);
nand U12628 (N_12628,N_11195,N_11865);
or U12629 (N_12629,N_11912,N_11388);
or U12630 (N_12630,N_11441,N_11610);
xor U12631 (N_12631,N_11967,N_11533);
nor U12632 (N_12632,N_11614,N_11725);
nand U12633 (N_12633,N_11237,N_11077);
and U12634 (N_12634,N_11603,N_11613);
and U12635 (N_12635,N_11825,N_11637);
nor U12636 (N_12636,N_11624,N_11478);
or U12637 (N_12637,N_11925,N_11097);
and U12638 (N_12638,N_11359,N_11290);
nor U12639 (N_12639,N_11360,N_11375);
nor U12640 (N_12640,N_11564,N_11034);
or U12641 (N_12641,N_11216,N_11142);
or U12642 (N_12642,N_11267,N_11209);
xnor U12643 (N_12643,N_11058,N_11519);
nand U12644 (N_12644,N_11647,N_11959);
or U12645 (N_12645,N_11040,N_11772);
nand U12646 (N_12646,N_11222,N_11291);
and U12647 (N_12647,N_11830,N_11532);
and U12648 (N_12648,N_11467,N_11772);
nand U12649 (N_12649,N_11169,N_11965);
or U12650 (N_12650,N_11091,N_11909);
nand U12651 (N_12651,N_11811,N_11261);
nor U12652 (N_12652,N_11974,N_11311);
or U12653 (N_12653,N_11185,N_11657);
and U12654 (N_12654,N_11102,N_11920);
nor U12655 (N_12655,N_11814,N_11757);
nor U12656 (N_12656,N_11062,N_11088);
nand U12657 (N_12657,N_11922,N_11144);
and U12658 (N_12658,N_11784,N_11386);
nor U12659 (N_12659,N_11635,N_11792);
xor U12660 (N_12660,N_11448,N_11256);
nand U12661 (N_12661,N_11937,N_11288);
nor U12662 (N_12662,N_11803,N_11187);
nor U12663 (N_12663,N_11695,N_11833);
or U12664 (N_12664,N_11415,N_11073);
and U12665 (N_12665,N_11615,N_11067);
nor U12666 (N_12666,N_11108,N_11053);
xnor U12667 (N_12667,N_11794,N_11120);
nor U12668 (N_12668,N_11000,N_11615);
xor U12669 (N_12669,N_11008,N_11990);
nand U12670 (N_12670,N_11838,N_11856);
nand U12671 (N_12671,N_11644,N_11091);
xor U12672 (N_12672,N_11631,N_11952);
xnor U12673 (N_12673,N_11517,N_11442);
or U12674 (N_12674,N_11612,N_11791);
and U12675 (N_12675,N_11197,N_11848);
nor U12676 (N_12676,N_11630,N_11674);
and U12677 (N_12677,N_11431,N_11003);
and U12678 (N_12678,N_11560,N_11581);
nand U12679 (N_12679,N_11747,N_11793);
nor U12680 (N_12680,N_11797,N_11554);
nor U12681 (N_12681,N_11438,N_11684);
and U12682 (N_12682,N_11939,N_11595);
xor U12683 (N_12683,N_11448,N_11921);
or U12684 (N_12684,N_11607,N_11072);
and U12685 (N_12685,N_11881,N_11756);
nor U12686 (N_12686,N_11343,N_11389);
or U12687 (N_12687,N_11897,N_11198);
and U12688 (N_12688,N_11450,N_11587);
or U12689 (N_12689,N_11741,N_11284);
and U12690 (N_12690,N_11540,N_11128);
and U12691 (N_12691,N_11492,N_11316);
or U12692 (N_12692,N_11520,N_11620);
and U12693 (N_12693,N_11611,N_11725);
nand U12694 (N_12694,N_11240,N_11673);
nand U12695 (N_12695,N_11661,N_11923);
xnor U12696 (N_12696,N_11830,N_11331);
or U12697 (N_12697,N_11342,N_11049);
nor U12698 (N_12698,N_11929,N_11173);
and U12699 (N_12699,N_11959,N_11790);
nand U12700 (N_12700,N_11959,N_11685);
or U12701 (N_12701,N_11258,N_11689);
nand U12702 (N_12702,N_11420,N_11312);
or U12703 (N_12703,N_11482,N_11747);
nor U12704 (N_12704,N_11353,N_11218);
or U12705 (N_12705,N_11418,N_11697);
and U12706 (N_12706,N_11824,N_11407);
xor U12707 (N_12707,N_11974,N_11665);
and U12708 (N_12708,N_11921,N_11711);
or U12709 (N_12709,N_11940,N_11251);
nor U12710 (N_12710,N_11496,N_11434);
nand U12711 (N_12711,N_11408,N_11128);
nand U12712 (N_12712,N_11695,N_11792);
and U12713 (N_12713,N_11133,N_11147);
and U12714 (N_12714,N_11299,N_11831);
or U12715 (N_12715,N_11128,N_11892);
and U12716 (N_12716,N_11458,N_11589);
nor U12717 (N_12717,N_11510,N_11601);
nor U12718 (N_12718,N_11944,N_11102);
nor U12719 (N_12719,N_11102,N_11713);
nand U12720 (N_12720,N_11308,N_11548);
and U12721 (N_12721,N_11164,N_11624);
nand U12722 (N_12722,N_11964,N_11917);
nand U12723 (N_12723,N_11513,N_11924);
xnor U12724 (N_12724,N_11516,N_11505);
nand U12725 (N_12725,N_11085,N_11362);
or U12726 (N_12726,N_11540,N_11649);
or U12727 (N_12727,N_11555,N_11408);
nor U12728 (N_12728,N_11357,N_11679);
and U12729 (N_12729,N_11922,N_11283);
nand U12730 (N_12730,N_11685,N_11848);
nand U12731 (N_12731,N_11740,N_11704);
and U12732 (N_12732,N_11863,N_11588);
or U12733 (N_12733,N_11681,N_11087);
and U12734 (N_12734,N_11797,N_11304);
or U12735 (N_12735,N_11104,N_11454);
and U12736 (N_12736,N_11758,N_11827);
and U12737 (N_12737,N_11734,N_11804);
nand U12738 (N_12738,N_11615,N_11512);
nand U12739 (N_12739,N_11158,N_11007);
nand U12740 (N_12740,N_11699,N_11574);
or U12741 (N_12741,N_11966,N_11387);
or U12742 (N_12742,N_11056,N_11925);
and U12743 (N_12743,N_11391,N_11640);
and U12744 (N_12744,N_11589,N_11479);
xnor U12745 (N_12745,N_11537,N_11563);
or U12746 (N_12746,N_11268,N_11388);
or U12747 (N_12747,N_11040,N_11942);
or U12748 (N_12748,N_11216,N_11937);
nand U12749 (N_12749,N_11897,N_11025);
nand U12750 (N_12750,N_11334,N_11987);
nand U12751 (N_12751,N_11237,N_11158);
nand U12752 (N_12752,N_11221,N_11051);
or U12753 (N_12753,N_11135,N_11742);
xor U12754 (N_12754,N_11712,N_11349);
nand U12755 (N_12755,N_11534,N_11777);
or U12756 (N_12756,N_11646,N_11627);
nor U12757 (N_12757,N_11697,N_11395);
nand U12758 (N_12758,N_11616,N_11834);
nand U12759 (N_12759,N_11697,N_11609);
or U12760 (N_12760,N_11933,N_11287);
or U12761 (N_12761,N_11957,N_11002);
nor U12762 (N_12762,N_11930,N_11966);
nor U12763 (N_12763,N_11949,N_11493);
nand U12764 (N_12764,N_11767,N_11910);
nor U12765 (N_12765,N_11352,N_11765);
or U12766 (N_12766,N_11361,N_11075);
nand U12767 (N_12767,N_11394,N_11747);
nand U12768 (N_12768,N_11498,N_11701);
and U12769 (N_12769,N_11417,N_11406);
and U12770 (N_12770,N_11116,N_11570);
nand U12771 (N_12771,N_11898,N_11455);
and U12772 (N_12772,N_11591,N_11252);
or U12773 (N_12773,N_11896,N_11153);
nor U12774 (N_12774,N_11069,N_11383);
and U12775 (N_12775,N_11271,N_11125);
or U12776 (N_12776,N_11599,N_11339);
nor U12777 (N_12777,N_11767,N_11706);
nor U12778 (N_12778,N_11246,N_11974);
nor U12779 (N_12779,N_11874,N_11401);
nand U12780 (N_12780,N_11069,N_11611);
xor U12781 (N_12781,N_11554,N_11972);
and U12782 (N_12782,N_11838,N_11533);
nand U12783 (N_12783,N_11764,N_11281);
and U12784 (N_12784,N_11491,N_11650);
and U12785 (N_12785,N_11898,N_11954);
or U12786 (N_12786,N_11076,N_11233);
or U12787 (N_12787,N_11285,N_11398);
or U12788 (N_12788,N_11267,N_11741);
and U12789 (N_12789,N_11902,N_11265);
nor U12790 (N_12790,N_11326,N_11372);
nor U12791 (N_12791,N_11768,N_11569);
nor U12792 (N_12792,N_11442,N_11170);
and U12793 (N_12793,N_11864,N_11450);
xnor U12794 (N_12794,N_11697,N_11161);
or U12795 (N_12795,N_11456,N_11412);
nand U12796 (N_12796,N_11728,N_11001);
nand U12797 (N_12797,N_11420,N_11807);
nand U12798 (N_12798,N_11588,N_11439);
nand U12799 (N_12799,N_11495,N_11248);
and U12800 (N_12800,N_11833,N_11853);
xor U12801 (N_12801,N_11889,N_11377);
nand U12802 (N_12802,N_11527,N_11876);
nor U12803 (N_12803,N_11701,N_11658);
nor U12804 (N_12804,N_11695,N_11731);
nor U12805 (N_12805,N_11760,N_11026);
or U12806 (N_12806,N_11601,N_11771);
nor U12807 (N_12807,N_11874,N_11327);
nor U12808 (N_12808,N_11497,N_11896);
or U12809 (N_12809,N_11529,N_11665);
nand U12810 (N_12810,N_11444,N_11085);
and U12811 (N_12811,N_11525,N_11510);
xnor U12812 (N_12812,N_11175,N_11044);
nor U12813 (N_12813,N_11463,N_11042);
nor U12814 (N_12814,N_11186,N_11609);
or U12815 (N_12815,N_11287,N_11646);
xor U12816 (N_12816,N_11663,N_11566);
nand U12817 (N_12817,N_11313,N_11394);
nor U12818 (N_12818,N_11974,N_11591);
or U12819 (N_12819,N_11266,N_11992);
nand U12820 (N_12820,N_11795,N_11878);
nand U12821 (N_12821,N_11395,N_11720);
nor U12822 (N_12822,N_11167,N_11235);
or U12823 (N_12823,N_11001,N_11489);
and U12824 (N_12824,N_11288,N_11538);
or U12825 (N_12825,N_11236,N_11528);
nor U12826 (N_12826,N_11837,N_11061);
or U12827 (N_12827,N_11021,N_11609);
nor U12828 (N_12828,N_11838,N_11954);
xor U12829 (N_12829,N_11165,N_11308);
and U12830 (N_12830,N_11107,N_11221);
or U12831 (N_12831,N_11620,N_11784);
nor U12832 (N_12832,N_11650,N_11652);
and U12833 (N_12833,N_11788,N_11885);
nand U12834 (N_12834,N_11200,N_11256);
nor U12835 (N_12835,N_11802,N_11178);
nand U12836 (N_12836,N_11215,N_11669);
and U12837 (N_12837,N_11318,N_11249);
nand U12838 (N_12838,N_11293,N_11605);
and U12839 (N_12839,N_11575,N_11302);
and U12840 (N_12840,N_11772,N_11866);
nor U12841 (N_12841,N_11770,N_11412);
xor U12842 (N_12842,N_11498,N_11212);
nand U12843 (N_12843,N_11500,N_11639);
nor U12844 (N_12844,N_11385,N_11098);
or U12845 (N_12845,N_11956,N_11325);
or U12846 (N_12846,N_11772,N_11759);
nand U12847 (N_12847,N_11820,N_11346);
nand U12848 (N_12848,N_11815,N_11008);
nor U12849 (N_12849,N_11493,N_11314);
and U12850 (N_12850,N_11619,N_11107);
or U12851 (N_12851,N_11928,N_11862);
nand U12852 (N_12852,N_11690,N_11078);
nor U12853 (N_12853,N_11572,N_11222);
nor U12854 (N_12854,N_11249,N_11497);
nor U12855 (N_12855,N_11087,N_11576);
and U12856 (N_12856,N_11869,N_11108);
and U12857 (N_12857,N_11175,N_11398);
or U12858 (N_12858,N_11492,N_11909);
xnor U12859 (N_12859,N_11024,N_11350);
or U12860 (N_12860,N_11163,N_11146);
nand U12861 (N_12861,N_11940,N_11541);
nor U12862 (N_12862,N_11699,N_11673);
xor U12863 (N_12863,N_11516,N_11160);
nor U12864 (N_12864,N_11234,N_11172);
nor U12865 (N_12865,N_11481,N_11093);
and U12866 (N_12866,N_11767,N_11687);
nand U12867 (N_12867,N_11788,N_11273);
and U12868 (N_12868,N_11906,N_11098);
nor U12869 (N_12869,N_11450,N_11447);
and U12870 (N_12870,N_11448,N_11645);
or U12871 (N_12871,N_11494,N_11911);
nand U12872 (N_12872,N_11616,N_11004);
or U12873 (N_12873,N_11220,N_11753);
nor U12874 (N_12874,N_11894,N_11302);
or U12875 (N_12875,N_11045,N_11367);
and U12876 (N_12876,N_11017,N_11087);
nand U12877 (N_12877,N_11567,N_11101);
and U12878 (N_12878,N_11428,N_11535);
nand U12879 (N_12879,N_11323,N_11682);
nor U12880 (N_12880,N_11440,N_11990);
nand U12881 (N_12881,N_11251,N_11001);
and U12882 (N_12882,N_11357,N_11554);
nand U12883 (N_12883,N_11074,N_11656);
nor U12884 (N_12884,N_11754,N_11647);
nor U12885 (N_12885,N_11083,N_11445);
nand U12886 (N_12886,N_11152,N_11910);
or U12887 (N_12887,N_11905,N_11666);
and U12888 (N_12888,N_11164,N_11461);
or U12889 (N_12889,N_11725,N_11412);
nor U12890 (N_12890,N_11054,N_11175);
or U12891 (N_12891,N_11371,N_11189);
and U12892 (N_12892,N_11447,N_11095);
and U12893 (N_12893,N_11324,N_11944);
or U12894 (N_12894,N_11283,N_11437);
or U12895 (N_12895,N_11225,N_11934);
nand U12896 (N_12896,N_11364,N_11819);
and U12897 (N_12897,N_11419,N_11459);
or U12898 (N_12898,N_11443,N_11843);
nand U12899 (N_12899,N_11970,N_11503);
nand U12900 (N_12900,N_11401,N_11793);
nor U12901 (N_12901,N_11401,N_11268);
and U12902 (N_12902,N_11177,N_11954);
and U12903 (N_12903,N_11597,N_11439);
nand U12904 (N_12904,N_11155,N_11746);
or U12905 (N_12905,N_11082,N_11512);
or U12906 (N_12906,N_11689,N_11926);
and U12907 (N_12907,N_11820,N_11567);
and U12908 (N_12908,N_11009,N_11554);
nor U12909 (N_12909,N_11560,N_11946);
or U12910 (N_12910,N_11525,N_11924);
or U12911 (N_12911,N_11272,N_11475);
or U12912 (N_12912,N_11442,N_11788);
or U12913 (N_12913,N_11722,N_11376);
nor U12914 (N_12914,N_11983,N_11654);
nand U12915 (N_12915,N_11668,N_11641);
nand U12916 (N_12916,N_11276,N_11827);
nor U12917 (N_12917,N_11972,N_11127);
xor U12918 (N_12918,N_11568,N_11555);
and U12919 (N_12919,N_11636,N_11847);
or U12920 (N_12920,N_11841,N_11978);
nor U12921 (N_12921,N_11830,N_11779);
nor U12922 (N_12922,N_11342,N_11998);
nor U12923 (N_12923,N_11625,N_11893);
nor U12924 (N_12924,N_11664,N_11528);
nor U12925 (N_12925,N_11918,N_11039);
nor U12926 (N_12926,N_11975,N_11154);
and U12927 (N_12927,N_11642,N_11968);
and U12928 (N_12928,N_11564,N_11601);
and U12929 (N_12929,N_11392,N_11335);
nor U12930 (N_12930,N_11455,N_11533);
xnor U12931 (N_12931,N_11603,N_11412);
nand U12932 (N_12932,N_11163,N_11715);
xor U12933 (N_12933,N_11247,N_11328);
nand U12934 (N_12934,N_11573,N_11482);
xnor U12935 (N_12935,N_11213,N_11629);
nor U12936 (N_12936,N_11742,N_11329);
or U12937 (N_12937,N_11547,N_11204);
and U12938 (N_12938,N_11048,N_11240);
and U12939 (N_12939,N_11573,N_11771);
or U12940 (N_12940,N_11317,N_11179);
nand U12941 (N_12941,N_11725,N_11668);
nand U12942 (N_12942,N_11327,N_11233);
nand U12943 (N_12943,N_11343,N_11197);
xnor U12944 (N_12944,N_11869,N_11717);
or U12945 (N_12945,N_11519,N_11807);
and U12946 (N_12946,N_11732,N_11509);
or U12947 (N_12947,N_11367,N_11211);
nand U12948 (N_12948,N_11851,N_11853);
nand U12949 (N_12949,N_11829,N_11009);
xnor U12950 (N_12950,N_11438,N_11815);
and U12951 (N_12951,N_11677,N_11508);
nor U12952 (N_12952,N_11492,N_11049);
nor U12953 (N_12953,N_11630,N_11330);
and U12954 (N_12954,N_11362,N_11164);
xor U12955 (N_12955,N_11192,N_11785);
nand U12956 (N_12956,N_11128,N_11439);
xor U12957 (N_12957,N_11254,N_11285);
xor U12958 (N_12958,N_11464,N_11375);
nand U12959 (N_12959,N_11010,N_11439);
nor U12960 (N_12960,N_11387,N_11998);
nor U12961 (N_12961,N_11884,N_11341);
nand U12962 (N_12962,N_11457,N_11781);
and U12963 (N_12963,N_11601,N_11629);
nand U12964 (N_12964,N_11583,N_11569);
nand U12965 (N_12965,N_11399,N_11580);
nor U12966 (N_12966,N_11542,N_11183);
nand U12967 (N_12967,N_11055,N_11762);
or U12968 (N_12968,N_11710,N_11396);
or U12969 (N_12969,N_11809,N_11138);
or U12970 (N_12970,N_11507,N_11255);
and U12971 (N_12971,N_11783,N_11033);
or U12972 (N_12972,N_11109,N_11974);
nand U12973 (N_12973,N_11555,N_11980);
and U12974 (N_12974,N_11333,N_11196);
or U12975 (N_12975,N_11956,N_11091);
xnor U12976 (N_12976,N_11223,N_11689);
nor U12977 (N_12977,N_11831,N_11557);
and U12978 (N_12978,N_11638,N_11449);
nand U12979 (N_12979,N_11989,N_11866);
nor U12980 (N_12980,N_11994,N_11472);
or U12981 (N_12981,N_11686,N_11843);
xnor U12982 (N_12982,N_11615,N_11021);
nand U12983 (N_12983,N_11894,N_11099);
or U12984 (N_12984,N_11434,N_11362);
or U12985 (N_12985,N_11691,N_11710);
or U12986 (N_12986,N_11884,N_11654);
and U12987 (N_12987,N_11272,N_11633);
or U12988 (N_12988,N_11865,N_11067);
and U12989 (N_12989,N_11624,N_11554);
or U12990 (N_12990,N_11273,N_11975);
and U12991 (N_12991,N_11758,N_11442);
and U12992 (N_12992,N_11615,N_11889);
and U12993 (N_12993,N_11975,N_11582);
nor U12994 (N_12994,N_11066,N_11906);
nand U12995 (N_12995,N_11534,N_11189);
or U12996 (N_12996,N_11662,N_11301);
nor U12997 (N_12997,N_11066,N_11506);
or U12998 (N_12998,N_11886,N_11229);
nor U12999 (N_12999,N_11376,N_11188);
nand U13000 (N_13000,N_12979,N_12315);
nand U13001 (N_13001,N_12652,N_12058);
nand U13002 (N_13002,N_12413,N_12593);
nand U13003 (N_13003,N_12530,N_12487);
nor U13004 (N_13004,N_12578,N_12672);
or U13005 (N_13005,N_12909,N_12544);
or U13006 (N_13006,N_12818,N_12049);
and U13007 (N_13007,N_12395,N_12637);
nand U13008 (N_13008,N_12113,N_12545);
nand U13009 (N_13009,N_12639,N_12954);
or U13010 (N_13010,N_12101,N_12475);
and U13011 (N_13011,N_12032,N_12916);
nand U13012 (N_13012,N_12884,N_12951);
or U13013 (N_13013,N_12861,N_12329);
nand U13014 (N_13014,N_12536,N_12580);
and U13015 (N_13015,N_12133,N_12467);
nand U13016 (N_13016,N_12505,N_12619);
or U13017 (N_13017,N_12958,N_12276);
or U13018 (N_13018,N_12196,N_12826);
nor U13019 (N_13019,N_12649,N_12110);
nor U13020 (N_13020,N_12965,N_12633);
nor U13021 (N_13021,N_12848,N_12504);
nor U13022 (N_13022,N_12096,N_12805);
or U13023 (N_13023,N_12136,N_12941);
nor U13024 (N_13024,N_12959,N_12379);
nor U13025 (N_13025,N_12881,N_12699);
and U13026 (N_13026,N_12044,N_12134);
or U13027 (N_13027,N_12849,N_12460);
nand U13028 (N_13028,N_12953,N_12787);
and U13029 (N_13029,N_12500,N_12791);
nand U13030 (N_13030,N_12983,N_12710);
xor U13031 (N_13031,N_12236,N_12159);
nor U13032 (N_13032,N_12198,N_12254);
or U13033 (N_13033,N_12410,N_12636);
and U13034 (N_13034,N_12701,N_12081);
and U13035 (N_13035,N_12003,N_12083);
nor U13036 (N_13036,N_12822,N_12911);
xor U13037 (N_13037,N_12857,N_12321);
nand U13038 (N_13038,N_12675,N_12577);
or U13039 (N_13039,N_12510,N_12999);
nand U13040 (N_13040,N_12926,N_12713);
nor U13041 (N_13041,N_12042,N_12168);
nor U13042 (N_13042,N_12807,N_12751);
nor U13043 (N_13043,N_12529,N_12148);
nand U13044 (N_13044,N_12520,N_12219);
xnor U13045 (N_13045,N_12444,N_12497);
nand U13046 (N_13046,N_12535,N_12803);
xor U13047 (N_13047,N_12694,N_12476);
nand U13048 (N_13048,N_12714,N_12768);
and U13049 (N_13049,N_12839,N_12738);
nand U13050 (N_13050,N_12871,N_12456);
nor U13051 (N_13051,N_12440,N_12836);
xor U13052 (N_13052,N_12496,N_12925);
xnor U13053 (N_13053,N_12682,N_12345);
nand U13054 (N_13054,N_12245,N_12062);
nor U13055 (N_13055,N_12862,N_12235);
nand U13056 (N_13056,N_12721,N_12128);
nand U13057 (N_13057,N_12406,N_12119);
nand U13058 (N_13058,N_12455,N_12767);
xnor U13059 (N_13059,N_12877,N_12354);
or U13060 (N_13060,N_12673,N_12976);
nor U13061 (N_13061,N_12648,N_12463);
or U13062 (N_13062,N_12481,N_12437);
xor U13063 (N_13063,N_12609,N_12495);
xnor U13064 (N_13064,N_12452,N_12688);
or U13065 (N_13065,N_12163,N_12937);
or U13066 (N_13066,N_12603,N_12352);
nor U13067 (N_13067,N_12788,N_12125);
nand U13068 (N_13068,N_12108,N_12424);
nand U13069 (N_13069,N_12991,N_12224);
and U13070 (N_13070,N_12122,N_12080);
or U13071 (N_13071,N_12347,N_12392);
or U13072 (N_13072,N_12982,N_12160);
nor U13073 (N_13073,N_12888,N_12929);
nand U13074 (N_13074,N_12330,N_12383);
nand U13075 (N_13075,N_12170,N_12301);
nor U13076 (N_13076,N_12028,N_12720);
xnor U13077 (N_13077,N_12109,N_12284);
nor U13078 (N_13078,N_12450,N_12401);
and U13079 (N_13079,N_12311,N_12290);
xor U13080 (N_13080,N_12774,N_12970);
nand U13081 (N_13081,N_12506,N_12686);
nand U13082 (N_13082,N_12581,N_12928);
and U13083 (N_13083,N_12860,N_12555);
or U13084 (N_13084,N_12008,N_12033);
or U13085 (N_13085,N_12115,N_12375);
nor U13086 (N_13086,N_12422,N_12280);
and U13087 (N_13087,N_12069,N_12785);
or U13088 (N_13088,N_12945,N_12309);
or U13089 (N_13089,N_12575,N_12644);
and U13090 (N_13090,N_12182,N_12762);
xnor U13091 (N_13091,N_12854,N_12833);
nand U13092 (N_13092,N_12263,N_12146);
xor U13093 (N_13093,N_12723,N_12292);
and U13094 (N_13094,N_12709,N_12902);
nor U13095 (N_13095,N_12990,N_12297);
and U13096 (N_13096,N_12967,N_12327);
and U13097 (N_13097,N_12607,N_12835);
nand U13098 (N_13098,N_12149,N_12766);
or U13099 (N_13099,N_12055,N_12317);
and U13100 (N_13100,N_12678,N_12514);
or U13101 (N_13101,N_12606,N_12441);
nor U13102 (N_13102,N_12592,N_12576);
or U13103 (N_13103,N_12906,N_12409);
nor U13104 (N_13104,N_12795,N_12247);
or U13105 (N_13105,N_12433,N_12138);
and U13106 (N_13106,N_12800,N_12657);
nor U13107 (N_13107,N_12037,N_12980);
nor U13108 (N_13108,N_12621,N_12318);
or U13109 (N_13109,N_12391,N_12512);
and U13110 (N_13110,N_12377,N_12717);
xor U13111 (N_13111,N_12700,N_12869);
xnor U13112 (N_13112,N_12316,N_12057);
and U13113 (N_13113,N_12201,N_12761);
or U13114 (N_13114,N_12408,N_12564);
xnor U13115 (N_13115,N_12828,N_12977);
nand U13116 (N_13116,N_12640,N_12988);
or U13117 (N_13117,N_12732,N_12930);
nand U13118 (N_13118,N_12532,N_12322);
nand U13119 (N_13119,N_12540,N_12571);
nor U13120 (N_13120,N_12784,N_12842);
and U13121 (N_13121,N_12070,N_12104);
nor U13122 (N_13122,N_12656,N_12473);
nand U13123 (N_13123,N_12061,N_12563);
or U13124 (N_13124,N_12727,N_12708);
or U13125 (N_13125,N_12332,N_12974);
xnor U13126 (N_13126,N_12306,N_12390);
nand U13127 (N_13127,N_12211,N_12627);
or U13128 (N_13128,N_12030,N_12416);
nand U13129 (N_13129,N_12356,N_12915);
nand U13130 (N_13130,N_12060,N_12760);
or U13131 (N_13131,N_12089,N_12858);
xor U13132 (N_13132,N_12173,N_12283);
nor U13133 (N_13133,N_12430,N_12855);
nand U13134 (N_13134,N_12812,N_12882);
and U13135 (N_13135,N_12158,N_12259);
and U13136 (N_13136,N_12939,N_12502);
and U13137 (N_13137,N_12000,N_12396);
nand U13138 (N_13138,N_12194,N_12917);
or U13139 (N_13139,N_12400,N_12248);
nand U13140 (N_13140,N_12950,N_12852);
nor U13141 (N_13141,N_12658,N_12503);
nand U13142 (N_13142,N_12343,N_12013);
nand U13143 (N_13143,N_12667,N_12253);
nand U13144 (N_13144,N_12051,N_12489);
and U13145 (N_13145,N_12087,N_12695);
nor U13146 (N_13146,N_12479,N_12124);
or U13147 (N_13147,N_12689,N_12234);
xnor U13148 (N_13148,N_12781,N_12132);
or U13149 (N_13149,N_12419,N_12480);
or U13150 (N_13150,N_12217,N_12600);
nor U13151 (N_13151,N_12590,N_12517);
or U13152 (N_13152,N_12655,N_12866);
or U13153 (N_13153,N_12007,N_12046);
nand U13154 (N_13154,N_12940,N_12004);
and U13155 (N_13155,N_12078,N_12645);
or U13156 (N_13156,N_12300,N_12783);
nor U13157 (N_13157,N_12885,N_12670);
nand U13158 (N_13158,N_12048,N_12423);
nor U13159 (N_13159,N_12518,N_12207);
nand U13160 (N_13160,N_12523,N_12393);
nand U13161 (N_13161,N_12002,N_12741);
and U13162 (N_13162,N_12494,N_12439);
or U13163 (N_13163,N_12863,N_12955);
or U13164 (N_13164,N_12900,N_12746);
or U13165 (N_13165,N_12617,N_12735);
and U13166 (N_13166,N_12470,N_12522);
and U13167 (N_13167,N_12498,N_12039);
nor U13168 (N_13168,N_12326,N_12629);
nand U13169 (N_13169,N_12868,N_12432);
nor U13170 (N_13170,N_12985,N_12258);
and U13171 (N_13171,N_12829,N_12998);
nand U13172 (N_13172,N_12222,N_12521);
and U13173 (N_13173,N_12023,N_12230);
nor U13174 (N_13174,N_12483,N_12242);
and U13175 (N_13175,N_12105,N_12598);
nand U13176 (N_13176,N_12507,N_12696);
and U13177 (N_13177,N_12840,N_12759);
and U13178 (N_13178,N_12126,N_12485);
and U13179 (N_13179,N_12097,N_12385);
nor U13180 (N_13180,N_12140,N_12542);
and U13181 (N_13181,N_12750,N_12873);
or U13182 (N_13182,N_12334,N_12883);
or U13183 (N_13183,N_12978,N_12802);
nor U13184 (N_13184,N_12127,N_12511);
nand U13185 (N_13185,N_12891,N_12568);
or U13186 (N_13186,N_12734,N_12331);
or U13187 (N_13187,N_12045,N_12323);
nand U13188 (N_13188,N_12531,N_12528);
and U13189 (N_13189,N_12638,N_12583);
or U13190 (N_13190,N_12038,N_12887);
nor U13191 (N_13191,N_12265,N_12832);
and U13192 (N_13192,N_12449,N_12074);
nor U13193 (N_13193,N_12035,N_12252);
or U13194 (N_13194,N_12166,N_12348);
and U13195 (N_13195,N_12853,N_12993);
nand U13196 (N_13196,N_12626,N_12006);
or U13197 (N_13197,N_12421,N_12043);
nand U13198 (N_13198,N_12553,N_12556);
or U13199 (N_13199,N_12736,N_12777);
nor U13200 (N_13200,N_12691,N_12579);
or U13201 (N_13201,N_12756,N_12228);
and U13202 (N_13202,N_12956,N_12927);
and U13203 (N_13203,N_12962,N_12371);
nand U13204 (N_13204,N_12154,N_12015);
nand U13205 (N_13205,N_12091,N_12328);
xor U13206 (N_13206,N_12350,N_12693);
nor U13207 (N_13207,N_12223,N_12130);
nand U13208 (N_13208,N_12336,N_12183);
xnor U13209 (N_13209,N_12543,N_12561);
or U13210 (N_13210,N_12171,N_12031);
and U13211 (N_13211,N_12789,N_12403);
and U13212 (N_13212,N_12604,N_12139);
and U13213 (N_13213,N_12747,N_12373);
nand U13214 (N_13214,N_12359,N_12426);
and U13215 (N_13215,N_12973,N_12743);
or U13216 (N_13216,N_12968,N_12275);
and U13217 (N_13217,N_12680,N_12610);
nor U13218 (N_13218,N_12612,N_12066);
xnor U13219 (N_13219,N_12155,N_12303);
or U13220 (N_13220,N_12145,N_12548);
nand U13221 (N_13221,N_12492,N_12647);
nor U13222 (N_13222,N_12806,N_12402);
nor U13223 (N_13223,N_12079,N_12796);
and U13224 (N_13224,N_12907,N_12779);
and U13225 (N_13225,N_12067,N_12624);
nand U13226 (N_13226,N_12117,N_12608);
and U13227 (N_13227,N_12491,N_12856);
nand U13228 (N_13228,N_12341,N_12642);
and U13229 (N_13229,N_12794,N_12167);
nand U13230 (N_13230,N_12250,N_12466);
nand U13231 (N_13231,N_12308,N_12216);
nand U13232 (N_13232,N_12204,N_12454);
nand U13233 (N_13233,N_12244,N_12995);
nor U13234 (N_13234,N_12020,N_12804);
nor U13235 (N_13235,N_12305,N_12987);
or U13236 (N_13236,N_12464,N_12340);
nor U13237 (N_13237,N_12705,N_12560);
nand U13238 (N_13238,N_12256,N_12674);
nand U13239 (N_13239,N_12001,N_12525);
nand U13240 (N_13240,N_12009,N_12107);
xnor U13241 (N_13241,N_12394,N_12027);
nand U13242 (N_13242,N_12135,N_12143);
and U13243 (N_13243,N_12846,N_12792);
nor U13244 (N_13244,N_12809,N_12541);
nor U13245 (N_13245,N_12586,N_12770);
nand U13246 (N_13246,N_12274,N_12769);
xnor U13247 (N_13247,N_12195,N_12024);
nor U13248 (N_13248,N_12257,N_12239);
and U13249 (N_13249,N_12901,N_12462);
nor U13250 (N_13250,N_12844,N_12378);
xor U13251 (N_13251,N_12547,N_12029);
or U13252 (N_13252,N_12920,N_12093);
nor U13253 (N_13253,N_12989,N_12278);
nor U13254 (N_13254,N_12471,N_12838);
nor U13255 (N_13255,N_12914,N_12790);
nor U13256 (N_13256,N_12233,N_12716);
nand U13257 (N_13257,N_12073,N_12924);
nand U13258 (N_13258,N_12210,N_12212);
nand U13259 (N_13259,N_12427,N_12539);
or U13260 (N_13260,N_12273,N_12351);
or U13261 (N_13261,N_12650,N_12519);
nand U13262 (N_13262,N_12552,N_12773);
and U13263 (N_13263,N_12499,N_12251);
nor U13264 (N_13264,N_12227,N_12921);
or U13265 (N_13265,N_12095,N_12823);
nand U13266 (N_13266,N_12279,N_12342);
or U13267 (N_13267,N_12615,N_12411);
and U13268 (N_13268,N_12942,N_12076);
and U13269 (N_13269,N_12588,N_12116);
and U13270 (N_13270,N_12690,N_12960);
nand U13271 (N_13271,N_12684,N_12515);
and U13272 (N_13272,N_12362,N_12156);
nor U13273 (N_13273,N_12185,N_12438);
or U13274 (N_13274,N_12753,N_12214);
nand U13275 (N_13275,N_12249,N_12918);
nand U13276 (N_13276,N_12509,N_12706);
nor U13277 (N_13277,N_12053,N_12824);
nor U13278 (N_13278,N_12874,N_12090);
nor U13279 (N_13279,N_12022,N_12152);
xor U13280 (N_13280,N_12289,N_12559);
nor U13281 (N_13281,N_12034,N_12875);
or U13282 (N_13282,N_12641,N_12669);
xnor U13283 (N_13283,N_12014,N_12103);
or U13284 (N_13284,N_12739,N_12616);
or U13285 (N_13285,N_12890,N_12905);
nor U13286 (N_13286,N_12819,N_12246);
nor U13287 (N_13287,N_12360,N_12952);
or U13288 (N_13288,N_12845,N_12215);
and U13289 (N_13289,N_12338,N_12623);
or U13290 (N_13290,N_12546,N_12851);
nor U13291 (N_13291,N_12646,N_12268);
and U13292 (N_13292,N_12948,N_12238);
and U13293 (N_13293,N_12801,N_12932);
nor U13294 (N_13294,N_12816,N_12724);
and U13295 (N_13295,N_12389,N_12635);
nor U13296 (N_13296,N_12896,N_12237);
nand U13297 (N_13297,N_12831,N_12431);
and U13298 (N_13298,N_12188,N_12808);
xnor U13299 (N_13299,N_12262,N_12963);
nand U13300 (N_13300,N_12772,N_12165);
nand U13301 (N_13301,N_12704,N_12526);
or U13302 (N_13302,N_12661,N_12241);
nand U13303 (N_13303,N_12404,N_12825);
or U13304 (N_13304,N_12744,N_12021);
or U13305 (N_13305,N_12469,N_12298);
and U13306 (N_13306,N_12975,N_12407);
and U13307 (N_13307,N_12562,N_12969);
xnor U13308 (N_13308,N_12277,N_12361);
nand U13309 (N_13309,N_12077,N_12382);
xor U13310 (N_13310,N_12010,N_12782);
nand U13311 (N_13311,N_12663,N_12333);
or U13312 (N_13312,N_12012,N_12933);
nand U13313 (N_13313,N_12793,N_12313);
nor U13314 (N_13314,N_12414,N_12374);
and U13315 (N_13315,N_12162,N_12075);
xnor U13316 (N_13316,N_12558,N_12372);
or U13317 (N_13317,N_12111,N_12320);
and U13318 (N_13318,N_12981,N_12474);
nor U13319 (N_13319,N_12458,N_12453);
nor U13320 (N_13320,N_12179,N_12036);
nand U13321 (N_13321,N_12944,N_12550);
and U13322 (N_13322,N_12086,N_12209);
nor U13323 (N_13323,N_12484,N_12923);
nand U13324 (N_13324,N_12886,N_12820);
xnor U13325 (N_13325,N_12364,N_12304);
nand U13326 (N_13326,N_12018,N_12567);
xnor U13327 (N_13327,N_12731,N_12757);
and U13328 (N_13328,N_12765,N_12418);
nor U13329 (N_13329,N_12059,N_12112);
and U13330 (N_13330,N_12200,N_12026);
and U13331 (N_13331,N_12630,N_12936);
nor U13332 (N_13332,N_12711,N_12436);
xor U13333 (N_13333,N_12596,N_12570);
xor U13334 (N_13334,N_12798,N_12443);
and U13335 (N_13335,N_12837,N_12810);
nand U13336 (N_13336,N_12733,N_12821);
nand U13337 (N_13337,N_12919,N_12225);
or U13338 (N_13338,N_12533,N_12434);
xor U13339 (N_13339,N_12019,N_12368);
or U13340 (N_13340,N_12141,N_12270);
nor U13341 (N_13341,N_12972,N_12722);
nor U13342 (N_13342,N_12964,N_12755);
nand U13343 (N_13343,N_12282,N_12310);
nor U13344 (N_13344,N_12551,N_12063);
and U13345 (N_13345,N_12387,N_12879);
and U13346 (N_13346,N_12415,N_12557);
xor U13347 (N_13347,N_12703,N_12712);
xnor U13348 (N_13348,N_12082,N_12231);
nand U13349 (N_13349,N_12175,N_12817);
nand U13350 (N_13350,N_12870,N_12574);
or U13351 (N_13351,N_12643,N_12363);
nand U13352 (N_13352,N_12666,N_12177);
nand U13353 (N_13353,N_12589,N_12565);
nor U13354 (N_13354,N_12748,N_12346);
and U13355 (N_13355,N_12946,N_12388);
and U13356 (N_13356,N_12516,N_12584);
nor U13357 (N_13357,N_12813,N_12157);
and U13358 (N_13358,N_12786,N_12631);
and U13359 (N_13359,N_12448,N_12676);
or U13360 (N_13360,N_12996,N_12005);
xnor U13361 (N_13361,N_12100,N_12490);
and U13362 (N_13362,N_12611,N_12572);
xnor U13363 (N_13363,N_12120,N_12662);
xnor U13364 (N_13364,N_12653,N_12827);
or U13365 (N_13365,N_12065,N_12957);
nand U13366 (N_13366,N_12595,N_12737);
or U13367 (N_13367,N_12291,N_12938);
nor U13368 (N_13368,N_12478,N_12834);
or U13369 (N_13369,N_12671,N_12961);
nand U13370 (N_13370,N_12587,N_12754);
nor U13371 (N_13371,N_12594,N_12685);
nor U13372 (N_13372,N_12660,N_12084);
nand U13373 (N_13373,N_12072,N_12651);
nand U13374 (N_13374,N_12205,N_12319);
nand U13375 (N_13375,N_12047,N_12707);
and U13376 (N_13376,N_12880,N_12186);
xor U13377 (N_13377,N_12174,N_12266);
nor U13378 (N_13378,N_12295,N_12614);
nor U13379 (N_13379,N_12098,N_12420);
nor U13380 (N_13380,N_12730,N_12847);
and U13381 (N_13381,N_12445,N_12294);
or U13382 (N_13382,N_12221,N_12632);
nor U13383 (N_13383,N_12085,N_12935);
nand U13384 (N_13384,N_12203,N_12366);
nor U13385 (N_13385,N_12137,N_12399);
or U13386 (N_13386,N_12613,N_12698);
xnor U13387 (N_13387,N_12740,N_12355);
nand U13388 (N_13388,N_12878,N_12269);
xor U13389 (N_13389,N_12229,N_12011);
xnor U13390 (N_13390,N_12573,N_12524);
xnor U13391 (N_13391,N_12240,N_12050);
xnor U13392 (N_13392,N_12697,N_12190);
nand U13393 (N_13393,N_12293,N_12056);
nand U13394 (N_13394,N_12797,N_12850);
and U13395 (N_13395,N_12199,N_12908);
and U13396 (N_13396,N_12147,N_12226);
or U13397 (N_13397,N_12380,N_12771);
or U13398 (N_13398,N_12349,N_12859);
nand U13399 (N_13399,N_12465,N_12264);
nor U13400 (N_13400,N_12193,N_12742);
nor U13401 (N_13401,N_12202,N_12068);
or U13402 (N_13402,N_12634,N_12129);
and U13403 (N_13403,N_12367,N_12106);
nor U13404 (N_13404,N_12830,N_12071);
nor U13405 (N_13405,N_12429,N_12114);
or U13406 (N_13406,N_12865,N_12272);
nand U13407 (N_13407,N_12243,N_12161);
xor U13408 (N_13408,N_12312,N_12417);
nand U13409 (N_13409,N_12934,N_12679);
nor U13410 (N_13410,N_12017,N_12131);
nor U13411 (N_13411,N_12527,N_12447);
or U13412 (N_13412,N_12446,N_12435);
nand U13413 (N_13413,N_12534,N_12867);
and U13414 (N_13414,N_12370,N_12041);
or U13415 (N_13415,N_12687,N_12997);
or U13416 (N_13416,N_12016,N_12442);
xnor U13417 (N_13417,N_12745,N_12189);
nor U13418 (N_13418,N_12913,N_12181);
or U13419 (N_13419,N_12299,N_12943);
nand U13420 (N_13420,N_12052,N_12457);
and U13421 (N_13421,N_12752,N_12776);
nor U13422 (N_13422,N_12549,N_12285);
or U13423 (N_13423,N_12296,N_12513);
nor U13424 (N_13424,N_12984,N_12889);
nand U13425 (N_13425,N_12728,N_12267);
and U13426 (N_13426,N_12151,N_12715);
and U13427 (N_13427,N_12625,N_12287);
or U13428 (N_13428,N_12054,N_12729);
and U13429 (N_13429,N_12893,N_12582);
nor U13430 (N_13430,N_12213,N_12898);
xnor U13431 (N_13431,N_12337,N_12585);
nand U13432 (N_13432,N_12628,N_12099);
nor U13433 (N_13433,N_12904,N_12654);
nand U13434 (N_13434,N_12261,N_12064);
or U13435 (N_13435,N_12620,N_12398);
nor U13436 (N_13436,N_12597,N_12659);
and U13437 (N_13437,N_12899,N_12092);
and U13438 (N_13438,N_12922,N_12903);
or U13439 (N_13439,N_12702,N_12187);
and U13440 (N_13440,N_12947,N_12508);
nor U13441 (N_13441,N_12425,N_12488);
or U13442 (N_13442,N_12569,N_12949);
or U13443 (N_13443,N_12232,N_12286);
nand U13444 (N_13444,N_12208,N_12986);
or U13445 (N_13445,N_12314,N_12353);
or U13446 (N_13446,N_12386,N_12472);
nand U13447 (N_13447,N_12566,N_12271);
nand U13448 (N_13448,N_12864,N_12895);
nor U13449 (N_13449,N_12144,N_12780);
or U13450 (N_13450,N_12405,N_12477);
or U13451 (N_13451,N_12601,N_12622);
xnor U13452 (N_13452,N_12538,N_12335);
nor U13453 (N_13453,N_12554,N_12912);
nor U13454 (N_13454,N_12381,N_12220);
nor U13455 (N_13455,N_12384,N_12180);
and U13456 (N_13456,N_12118,N_12164);
nor U13457 (N_13457,N_12365,N_12339);
nand U13458 (N_13458,N_12843,N_12142);
or U13459 (N_13459,N_12094,N_12197);
or U13460 (N_13460,N_12599,N_12811);
nor U13461 (N_13461,N_12677,N_12357);
nand U13462 (N_13462,N_12176,N_12537);
and U13463 (N_13463,N_12994,N_12665);
nand U13464 (N_13464,N_12681,N_12764);
or U13465 (N_13465,N_12664,N_12025);
or U13466 (N_13466,N_12178,N_12501);
and U13467 (N_13467,N_12897,N_12692);
or U13468 (N_13468,N_12778,N_12892);
or U13469 (N_13469,N_12260,N_12992);
and U13470 (N_13470,N_12894,N_12121);
nand U13471 (N_13471,N_12758,N_12325);
or U13472 (N_13472,N_12344,N_12281);
or U13473 (N_13473,N_12971,N_12482);
nor U13474 (N_13474,N_12369,N_12169);
or U13475 (N_13475,N_12966,N_12428);
nor U13476 (N_13476,N_12397,N_12876);
xor U13477 (N_13477,N_12088,N_12872);
or U13478 (N_13478,N_12123,N_12451);
nor U13479 (N_13479,N_12493,N_12461);
nand U13480 (N_13480,N_12206,N_12931);
nor U13481 (N_13481,N_12725,N_12668);
and U13482 (N_13482,N_12719,N_12815);
or U13483 (N_13483,N_12172,N_12288);
nor U13484 (N_13484,N_12605,N_12153);
nor U13485 (N_13485,N_12102,N_12763);
and U13486 (N_13486,N_12184,N_12618);
and U13487 (N_13487,N_12718,N_12468);
nand U13488 (N_13488,N_12683,N_12799);
xor U13489 (N_13489,N_12412,N_12602);
nor U13490 (N_13490,N_12192,N_12255);
and U13491 (N_13491,N_12040,N_12302);
or U13492 (N_13492,N_12910,N_12307);
and U13493 (N_13493,N_12459,N_12150);
and U13494 (N_13494,N_12814,N_12324);
nand U13495 (N_13495,N_12191,N_12841);
nand U13496 (N_13496,N_12749,N_12726);
nor U13497 (N_13497,N_12486,N_12591);
or U13498 (N_13498,N_12358,N_12775);
and U13499 (N_13499,N_12376,N_12218);
and U13500 (N_13500,N_12232,N_12148);
or U13501 (N_13501,N_12531,N_12285);
or U13502 (N_13502,N_12093,N_12991);
nor U13503 (N_13503,N_12637,N_12002);
and U13504 (N_13504,N_12906,N_12049);
or U13505 (N_13505,N_12653,N_12924);
nand U13506 (N_13506,N_12045,N_12011);
nand U13507 (N_13507,N_12752,N_12722);
nand U13508 (N_13508,N_12903,N_12646);
nor U13509 (N_13509,N_12146,N_12973);
or U13510 (N_13510,N_12125,N_12731);
nor U13511 (N_13511,N_12381,N_12143);
or U13512 (N_13512,N_12616,N_12180);
nand U13513 (N_13513,N_12530,N_12439);
nor U13514 (N_13514,N_12635,N_12344);
nor U13515 (N_13515,N_12238,N_12532);
nand U13516 (N_13516,N_12323,N_12974);
nor U13517 (N_13517,N_12723,N_12284);
and U13518 (N_13518,N_12950,N_12245);
or U13519 (N_13519,N_12676,N_12992);
xnor U13520 (N_13520,N_12296,N_12430);
nor U13521 (N_13521,N_12314,N_12460);
and U13522 (N_13522,N_12437,N_12736);
and U13523 (N_13523,N_12361,N_12620);
xnor U13524 (N_13524,N_12829,N_12254);
and U13525 (N_13525,N_12573,N_12346);
or U13526 (N_13526,N_12800,N_12530);
and U13527 (N_13527,N_12533,N_12098);
nor U13528 (N_13528,N_12143,N_12028);
nand U13529 (N_13529,N_12929,N_12714);
nand U13530 (N_13530,N_12729,N_12366);
nor U13531 (N_13531,N_12583,N_12688);
and U13532 (N_13532,N_12771,N_12268);
nor U13533 (N_13533,N_12757,N_12491);
and U13534 (N_13534,N_12764,N_12931);
nand U13535 (N_13535,N_12715,N_12824);
or U13536 (N_13536,N_12674,N_12657);
and U13537 (N_13537,N_12225,N_12437);
xnor U13538 (N_13538,N_12022,N_12885);
and U13539 (N_13539,N_12821,N_12370);
nor U13540 (N_13540,N_12235,N_12185);
or U13541 (N_13541,N_12662,N_12779);
nand U13542 (N_13542,N_12132,N_12919);
or U13543 (N_13543,N_12213,N_12035);
nand U13544 (N_13544,N_12538,N_12971);
nor U13545 (N_13545,N_12508,N_12929);
nand U13546 (N_13546,N_12441,N_12573);
nor U13547 (N_13547,N_12889,N_12708);
nor U13548 (N_13548,N_12362,N_12126);
or U13549 (N_13549,N_12090,N_12015);
nand U13550 (N_13550,N_12297,N_12868);
or U13551 (N_13551,N_12620,N_12856);
nor U13552 (N_13552,N_12710,N_12570);
xor U13553 (N_13553,N_12456,N_12676);
nor U13554 (N_13554,N_12774,N_12050);
and U13555 (N_13555,N_12425,N_12137);
nand U13556 (N_13556,N_12302,N_12309);
nor U13557 (N_13557,N_12184,N_12463);
nand U13558 (N_13558,N_12641,N_12566);
nor U13559 (N_13559,N_12487,N_12650);
and U13560 (N_13560,N_12469,N_12906);
nand U13561 (N_13561,N_12485,N_12678);
nor U13562 (N_13562,N_12867,N_12187);
and U13563 (N_13563,N_12555,N_12688);
or U13564 (N_13564,N_12415,N_12205);
nor U13565 (N_13565,N_12660,N_12439);
nor U13566 (N_13566,N_12399,N_12798);
nand U13567 (N_13567,N_12082,N_12854);
or U13568 (N_13568,N_12447,N_12055);
nand U13569 (N_13569,N_12793,N_12608);
xor U13570 (N_13570,N_12454,N_12302);
nor U13571 (N_13571,N_12808,N_12267);
or U13572 (N_13572,N_12765,N_12614);
nand U13573 (N_13573,N_12723,N_12136);
and U13574 (N_13574,N_12624,N_12192);
or U13575 (N_13575,N_12726,N_12351);
and U13576 (N_13576,N_12447,N_12362);
nand U13577 (N_13577,N_12288,N_12383);
nand U13578 (N_13578,N_12306,N_12728);
and U13579 (N_13579,N_12891,N_12682);
or U13580 (N_13580,N_12250,N_12541);
nand U13581 (N_13581,N_12938,N_12129);
xnor U13582 (N_13582,N_12469,N_12387);
or U13583 (N_13583,N_12542,N_12751);
nand U13584 (N_13584,N_12741,N_12305);
or U13585 (N_13585,N_12048,N_12998);
and U13586 (N_13586,N_12173,N_12818);
and U13587 (N_13587,N_12224,N_12302);
nand U13588 (N_13588,N_12100,N_12528);
or U13589 (N_13589,N_12963,N_12118);
and U13590 (N_13590,N_12473,N_12900);
or U13591 (N_13591,N_12908,N_12527);
nor U13592 (N_13592,N_12901,N_12204);
nand U13593 (N_13593,N_12216,N_12200);
nor U13594 (N_13594,N_12151,N_12771);
nand U13595 (N_13595,N_12989,N_12956);
and U13596 (N_13596,N_12880,N_12287);
nor U13597 (N_13597,N_12098,N_12531);
or U13598 (N_13598,N_12574,N_12382);
and U13599 (N_13599,N_12469,N_12639);
nor U13600 (N_13600,N_12438,N_12017);
or U13601 (N_13601,N_12566,N_12153);
and U13602 (N_13602,N_12192,N_12318);
and U13603 (N_13603,N_12476,N_12769);
xor U13604 (N_13604,N_12724,N_12274);
or U13605 (N_13605,N_12889,N_12652);
xnor U13606 (N_13606,N_12675,N_12779);
or U13607 (N_13607,N_12694,N_12010);
nor U13608 (N_13608,N_12825,N_12858);
or U13609 (N_13609,N_12065,N_12487);
and U13610 (N_13610,N_12057,N_12265);
xor U13611 (N_13611,N_12863,N_12978);
and U13612 (N_13612,N_12540,N_12328);
or U13613 (N_13613,N_12052,N_12557);
xor U13614 (N_13614,N_12425,N_12643);
nor U13615 (N_13615,N_12515,N_12397);
and U13616 (N_13616,N_12228,N_12443);
nor U13617 (N_13617,N_12463,N_12436);
or U13618 (N_13618,N_12342,N_12590);
and U13619 (N_13619,N_12015,N_12832);
or U13620 (N_13620,N_12345,N_12559);
xor U13621 (N_13621,N_12426,N_12738);
xnor U13622 (N_13622,N_12042,N_12758);
or U13623 (N_13623,N_12904,N_12636);
or U13624 (N_13624,N_12679,N_12541);
nand U13625 (N_13625,N_12557,N_12791);
nor U13626 (N_13626,N_12481,N_12365);
nor U13627 (N_13627,N_12229,N_12012);
and U13628 (N_13628,N_12358,N_12790);
or U13629 (N_13629,N_12352,N_12110);
nor U13630 (N_13630,N_12688,N_12093);
nand U13631 (N_13631,N_12025,N_12655);
or U13632 (N_13632,N_12982,N_12800);
or U13633 (N_13633,N_12178,N_12619);
and U13634 (N_13634,N_12542,N_12106);
nor U13635 (N_13635,N_12916,N_12570);
and U13636 (N_13636,N_12959,N_12935);
nor U13637 (N_13637,N_12467,N_12090);
and U13638 (N_13638,N_12246,N_12304);
nor U13639 (N_13639,N_12345,N_12783);
nor U13640 (N_13640,N_12375,N_12018);
and U13641 (N_13641,N_12777,N_12007);
and U13642 (N_13642,N_12397,N_12201);
nor U13643 (N_13643,N_12220,N_12841);
nor U13644 (N_13644,N_12629,N_12702);
and U13645 (N_13645,N_12478,N_12611);
and U13646 (N_13646,N_12971,N_12041);
or U13647 (N_13647,N_12337,N_12750);
nand U13648 (N_13648,N_12010,N_12044);
nand U13649 (N_13649,N_12267,N_12806);
or U13650 (N_13650,N_12732,N_12767);
nand U13651 (N_13651,N_12831,N_12621);
nor U13652 (N_13652,N_12582,N_12305);
nor U13653 (N_13653,N_12706,N_12791);
nand U13654 (N_13654,N_12427,N_12489);
nand U13655 (N_13655,N_12263,N_12682);
and U13656 (N_13656,N_12749,N_12826);
or U13657 (N_13657,N_12461,N_12152);
nand U13658 (N_13658,N_12181,N_12614);
xor U13659 (N_13659,N_12152,N_12653);
nor U13660 (N_13660,N_12495,N_12298);
and U13661 (N_13661,N_12723,N_12862);
or U13662 (N_13662,N_12658,N_12706);
nor U13663 (N_13663,N_12348,N_12129);
and U13664 (N_13664,N_12359,N_12165);
nor U13665 (N_13665,N_12572,N_12390);
and U13666 (N_13666,N_12005,N_12155);
or U13667 (N_13667,N_12972,N_12789);
or U13668 (N_13668,N_12684,N_12888);
nor U13669 (N_13669,N_12123,N_12950);
or U13670 (N_13670,N_12212,N_12929);
or U13671 (N_13671,N_12413,N_12276);
and U13672 (N_13672,N_12584,N_12007);
nor U13673 (N_13673,N_12677,N_12781);
or U13674 (N_13674,N_12257,N_12411);
or U13675 (N_13675,N_12072,N_12591);
xnor U13676 (N_13676,N_12808,N_12631);
or U13677 (N_13677,N_12646,N_12377);
or U13678 (N_13678,N_12089,N_12588);
or U13679 (N_13679,N_12592,N_12449);
nand U13680 (N_13680,N_12940,N_12554);
and U13681 (N_13681,N_12965,N_12973);
xnor U13682 (N_13682,N_12257,N_12753);
nor U13683 (N_13683,N_12512,N_12438);
and U13684 (N_13684,N_12011,N_12175);
nor U13685 (N_13685,N_12767,N_12200);
nor U13686 (N_13686,N_12362,N_12745);
nor U13687 (N_13687,N_12364,N_12046);
xnor U13688 (N_13688,N_12972,N_12595);
or U13689 (N_13689,N_12610,N_12336);
or U13690 (N_13690,N_12482,N_12355);
nor U13691 (N_13691,N_12913,N_12815);
xnor U13692 (N_13692,N_12743,N_12107);
nand U13693 (N_13693,N_12906,N_12691);
or U13694 (N_13694,N_12990,N_12565);
nand U13695 (N_13695,N_12491,N_12685);
xnor U13696 (N_13696,N_12456,N_12575);
nand U13697 (N_13697,N_12835,N_12740);
and U13698 (N_13698,N_12995,N_12439);
and U13699 (N_13699,N_12449,N_12636);
xor U13700 (N_13700,N_12848,N_12520);
and U13701 (N_13701,N_12287,N_12227);
and U13702 (N_13702,N_12424,N_12846);
nor U13703 (N_13703,N_12761,N_12821);
nor U13704 (N_13704,N_12407,N_12682);
or U13705 (N_13705,N_12978,N_12098);
or U13706 (N_13706,N_12291,N_12548);
xnor U13707 (N_13707,N_12221,N_12394);
xnor U13708 (N_13708,N_12731,N_12832);
and U13709 (N_13709,N_12686,N_12181);
nand U13710 (N_13710,N_12347,N_12224);
or U13711 (N_13711,N_12656,N_12815);
xor U13712 (N_13712,N_12558,N_12592);
and U13713 (N_13713,N_12161,N_12056);
and U13714 (N_13714,N_12139,N_12581);
nor U13715 (N_13715,N_12514,N_12220);
and U13716 (N_13716,N_12534,N_12947);
nor U13717 (N_13717,N_12325,N_12799);
nand U13718 (N_13718,N_12857,N_12511);
nand U13719 (N_13719,N_12379,N_12250);
nor U13720 (N_13720,N_12897,N_12057);
or U13721 (N_13721,N_12079,N_12194);
or U13722 (N_13722,N_12860,N_12658);
or U13723 (N_13723,N_12199,N_12860);
xor U13724 (N_13724,N_12492,N_12450);
nand U13725 (N_13725,N_12244,N_12318);
nand U13726 (N_13726,N_12526,N_12377);
and U13727 (N_13727,N_12369,N_12198);
xnor U13728 (N_13728,N_12433,N_12720);
nand U13729 (N_13729,N_12664,N_12640);
xnor U13730 (N_13730,N_12946,N_12094);
xnor U13731 (N_13731,N_12179,N_12646);
and U13732 (N_13732,N_12340,N_12193);
nand U13733 (N_13733,N_12941,N_12792);
xor U13734 (N_13734,N_12213,N_12922);
nor U13735 (N_13735,N_12349,N_12591);
or U13736 (N_13736,N_12731,N_12628);
nand U13737 (N_13737,N_12198,N_12498);
xor U13738 (N_13738,N_12304,N_12722);
and U13739 (N_13739,N_12752,N_12536);
or U13740 (N_13740,N_12385,N_12444);
nor U13741 (N_13741,N_12068,N_12394);
nand U13742 (N_13742,N_12533,N_12805);
nor U13743 (N_13743,N_12403,N_12148);
nor U13744 (N_13744,N_12927,N_12528);
nand U13745 (N_13745,N_12727,N_12679);
nor U13746 (N_13746,N_12436,N_12743);
xnor U13747 (N_13747,N_12729,N_12580);
nor U13748 (N_13748,N_12708,N_12089);
nand U13749 (N_13749,N_12204,N_12660);
or U13750 (N_13750,N_12173,N_12264);
or U13751 (N_13751,N_12369,N_12196);
and U13752 (N_13752,N_12563,N_12107);
nor U13753 (N_13753,N_12259,N_12624);
nor U13754 (N_13754,N_12079,N_12774);
or U13755 (N_13755,N_12831,N_12987);
nand U13756 (N_13756,N_12872,N_12370);
and U13757 (N_13757,N_12839,N_12648);
nor U13758 (N_13758,N_12219,N_12187);
and U13759 (N_13759,N_12499,N_12517);
or U13760 (N_13760,N_12896,N_12444);
and U13761 (N_13761,N_12717,N_12389);
nor U13762 (N_13762,N_12820,N_12503);
nand U13763 (N_13763,N_12627,N_12761);
xnor U13764 (N_13764,N_12975,N_12451);
nand U13765 (N_13765,N_12007,N_12971);
nor U13766 (N_13766,N_12347,N_12854);
nor U13767 (N_13767,N_12223,N_12400);
and U13768 (N_13768,N_12133,N_12143);
and U13769 (N_13769,N_12705,N_12631);
and U13770 (N_13770,N_12926,N_12541);
nand U13771 (N_13771,N_12173,N_12306);
nand U13772 (N_13772,N_12116,N_12072);
nor U13773 (N_13773,N_12670,N_12990);
nand U13774 (N_13774,N_12059,N_12122);
nor U13775 (N_13775,N_12164,N_12485);
and U13776 (N_13776,N_12496,N_12320);
xnor U13777 (N_13777,N_12874,N_12970);
nand U13778 (N_13778,N_12465,N_12044);
nand U13779 (N_13779,N_12962,N_12743);
and U13780 (N_13780,N_12882,N_12901);
or U13781 (N_13781,N_12008,N_12577);
or U13782 (N_13782,N_12101,N_12374);
or U13783 (N_13783,N_12484,N_12892);
nor U13784 (N_13784,N_12540,N_12588);
nand U13785 (N_13785,N_12173,N_12595);
or U13786 (N_13786,N_12062,N_12418);
and U13787 (N_13787,N_12654,N_12236);
or U13788 (N_13788,N_12981,N_12990);
and U13789 (N_13789,N_12054,N_12819);
or U13790 (N_13790,N_12592,N_12184);
nand U13791 (N_13791,N_12138,N_12271);
and U13792 (N_13792,N_12850,N_12727);
or U13793 (N_13793,N_12711,N_12693);
and U13794 (N_13794,N_12600,N_12614);
and U13795 (N_13795,N_12871,N_12673);
or U13796 (N_13796,N_12912,N_12402);
nand U13797 (N_13797,N_12696,N_12025);
xnor U13798 (N_13798,N_12387,N_12358);
and U13799 (N_13799,N_12861,N_12150);
or U13800 (N_13800,N_12511,N_12501);
nand U13801 (N_13801,N_12623,N_12287);
xnor U13802 (N_13802,N_12349,N_12006);
nor U13803 (N_13803,N_12492,N_12506);
or U13804 (N_13804,N_12197,N_12561);
and U13805 (N_13805,N_12148,N_12313);
nor U13806 (N_13806,N_12792,N_12956);
nor U13807 (N_13807,N_12473,N_12722);
and U13808 (N_13808,N_12614,N_12206);
nand U13809 (N_13809,N_12222,N_12378);
nand U13810 (N_13810,N_12277,N_12898);
nand U13811 (N_13811,N_12929,N_12222);
nand U13812 (N_13812,N_12804,N_12928);
nor U13813 (N_13813,N_12986,N_12694);
and U13814 (N_13814,N_12694,N_12597);
nor U13815 (N_13815,N_12592,N_12112);
and U13816 (N_13816,N_12044,N_12114);
or U13817 (N_13817,N_12479,N_12946);
nor U13818 (N_13818,N_12395,N_12064);
or U13819 (N_13819,N_12391,N_12212);
and U13820 (N_13820,N_12516,N_12079);
or U13821 (N_13821,N_12106,N_12083);
nand U13822 (N_13822,N_12747,N_12662);
and U13823 (N_13823,N_12507,N_12603);
xnor U13824 (N_13824,N_12394,N_12643);
nor U13825 (N_13825,N_12601,N_12504);
or U13826 (N_13826,N_12337,N_12145);
nand U13827 (N_13827,N_12571,N_12341);
nor U13828 (N_13828,N_12445,N_12616);
and U13829 (N_13829,N_12569,N_12436);
nand U13830 (N_13830,N_12901,N_12233);
nand U13831 (N_13831,N_12851,N_12163);
and U13832 (N_13832,N_12985,N_12881);
nand U13833 (N_13833,N_12803,N_12954);
nor U13834 (N_13834,N_12725,N_12431);
xor U13835 (N_13835,N_12505,N_12303);
nand U13836 (N_13836,N_12171,N_12776);
and U13837 (N_13837,N_12919,N_12009);
nor U13838 (N_13838,N_12291,N_12524);
nor U13839 (N_13839,N_12355,N_12211);
nand U13840 (N_13840,N_12509,N_12521);
nor U13841 (N_13841,N_12787,N_12062);
xor U13842 (N_13842,N_12985,N_12024);
nand U13843 (N_13843,N_12491,N_12741);
or U13844 (N_13844,N_12513,N_12057);
nand U13845 (N_13845,N_12782,N_12912);
and U13846 (N_13846,N_12472,N_12785);
or U13847 (N_13847,N_12690,N_12182);
xnor U13848 (N_13848,N_12871,N_12607);
nor U13849 (N_13849,N_12552,N_12544);
and U13850 (N_13850,N_12802,N_12606);
or U13851 (N_13851,N_12572,N_12477);
and U13852 (N_13852,N_12900,N_12856);
or U13853 (N_13853,N_12257,N_12166);
nor U13854 (N_13854,N_12219,N_12487);
or U13855 (N_13855,N_12429,N_12523);
nor U13856 (N_13856,N_12397,N_12786);
or U13857 (N_13857,N_12572,N_12874);
and U13858 (N_13858,N_12909,N_12434);
nor U13859 (N_13859,N_12743,N_12375);
nor U13860 (N_13860,N_12927,N_12386);
nand U13861 (N_13861,N_12233,N_12411);
nand U13862 (N_13862,N_12330,N_12531);
or U13863 (N_13863,N_12786,N_12117);
nor U13864 (N_13864,N_12944,N_12104);
nor U13865 (N_13865,N_12858,N_12640);
nand U13866 (N_13866,N_12820,N_12967);
nor U13867 (N_13867,N_12509,N_12091);
nor U13868 (N_13868,N_12928,N_12767);
nand U13869 (N_13869,N_12390,N_12448);
or U13870 (N_13870,N_12509,N_12000);
nand U13871 (N_13871,N_12311,N_12647);
or U13872 (N_13872,N_12929,N_12780);
and U13873 (N_13873,N_12686,N_12826);
xor U13874 (N_13874,N_12220,N_12716);
nor U13875 (N_13875,N_12986,N_12087);
nor U13876 (N_13876,N_12801,N_12460);
nand U13877 (N_13877,N_12233,N_12906);
nand U13878 (N_13878,N_12844,N_12673);
and U13879 (N_13879,N_12019,N_12862);
and U13880 (N_13880,N_12574,N_12752);
nand U13881 (N_13881,N_12744,N_12909);
nor U13882 (N_13882,N_12647,N_12733);
or U13883 (N_13883,N_12486,N_12519);
and U13884 (N_13884,N_12409,N_12047);
nand U13885 (N_13885,N_12595,N_12535);
nor U13886 (N_13886,N_12554,N_12018);
nor U13887 (N_13887,N_12488,N_12805);
nand U13888 (N_13888,N_12401,N_12875);
and U13889 (N_13889,N_12885,N_12272);
nor U13890 (N_13890,N_12815,N_12967);
nor U13891 (N_13891,N_12803,N_12610);
or U13892 (N_13892,N_12271,N_12864);
or U13893 (N_13893,N_12890,N_12564);
and U13894 (N_13894,N_12867,N_12676);
nor U13895 (N_13895,N_12076,N_12656);
xor U13896 (N_13896,N_12241,N_12398);
and U13897 (N_13897,N_12897,N_12736);
or U13898 (N_13898,N_12375,N_12241);
and U13899 (N_13899,N_12126,N_12607);
nor U13900 (N_13900,N_12452,N_12984);
and U13901 (N_13901,N_12509,N_12819);
nand U13902 (N_13902,N_12986,N_12478);
or U13903 (N_13903,N_12881,N_12465);
xnor U13904 (N_13904,N_12122,N_12789);
nor U13905 (N_13905,N_12680,N_12050);
or U13906 (N_13906,N_12489,N_12275);
or U13907 (N_13907,N_12583,N_12858);
and U13908 (N_13908,N_12464,N_12747);
nand U13909 (N_13909,N_12413,N_12368);
or U13910 (N_13910,N_12046,N_12331);
nor U13911 (N_13911,N_12230,N_12700);
xnor U13912 (N_13912,N_12879,N_12933);
nor U13913 (N_13913,N_12079,N_12524);
or U13914 (N_13914,N_12821,N_12669);
nand U13915 (N_13915,N_12885,N_12665);
and U13916 (N_13916,N_12433,N_12526);
nand U13917 (N_13917,N_12989,N_12362);
nor U13918 (N_13918,N_12799,N_12939);
nor U13919 (N_13919,N_12641,N_12560);
xor U13920 (N_13920,N_12780,N_12548);
or U13921 (N_13921,N_12053,N_12286);
nor U13922 (N_13922,N_12426,N_12443);
nor U13923 (N_13923,N_12134,N_12642);
nand U13924 (N_13924,N_12948,N_12356);
xor U13925 (N_13925,N_12173,N_12776);
and U13926 (N_13926,N_12589,N_12007);
xor U13927 (N_13927,N_12262,N_12276);
or U13928 (N_13928,N_12223,N_12148);
xor U13929 (N_13929,N_12812,N_12045);
xnor U13930 (N_13930,N_12174,N_12582);
xor U13931 (N_13931,N_12456,N_12595);
or U13932 (N_13932,N_12064,N_12610);
nand U13933 (N_13933,N_12306,N_12908);
nand U13934 (N_13934,N_12949,N_12883);
nor U13935 (N_13935,N_12961,N_12000);
or U13936 (N_13936,N_12459,N_12590);
or U13937 (N_13937,N_12308,N_12821);
and U13938 (N_13938,N_12367,N_12978);
and U13939 (N_13939,N_12881,N_12361);
nand U13940 (N_13940,N_12627,N_12531);
and U13941 (N_13941,N_12717,N_12683);
nand U13942 (N_13942,N_12881,N_12857);
or U13943 (N_13943,N_12918,N_12324);
and U13944 (N_13944,N_12763,N_12163);
or U13945 (N_13945,N_12642,N_12762);
and U13946 (N_13946,N_12729,N_12744);
nor U13947 (N_13947,N_12899,N_12413);
or U13948 (N_13948,N_12421,N_12584);
nor U13949 (N_13949,N_12080,N_12745);
nand U13950 (N_13950,N_12664,N_12083);
or U13951 (N_13951,N_12462,N_12209);
and U13952 (N_13952,N_12978,N_12487);
nor U13953 (N_13953,N_12238,N_12676);
or U13954 (N_13954,N_12521,N_12928);
nor U13955 (N_13955,N_12940,N_12570);
and U13956 (N_13956,N_12362,N_12879);
or U13957 (N_13957,N_12910,N_12630);
nor U13958 (N_13958,N_12160,N_12060);
or U13959 (N_13959,N_12875,N_12595);
or U13960 (N_13960,N_12045,N_12610);
or U13961 (N_13961,N_12736,N_12028);
xnor U13962 (N_13962,N_12376,N_12962);
nor U13963 (N_13963,N_12072,N_12381);
nand U13964 (N_13964,N_12420,N_12000);
and U13965 (N_13965,N_12681,N_12721);
xor U13966 (N_13966,N_12674,N_12066);
nand U13967 (N_13967,N_12027,N_12660);
nand U13968 (N_13968,N_12867,N_12705);
or U13969 (N_13969,N_12348,N_12624);
nor U13970 (N_13970,N_12173,N_12236);
nand U13971 (N_13971,N_12090,N_12173);
or U13972 (N_13972,N_12365,N_12374);
nor U13973 (N_13973,N_12187,N_12179);
and U13974 (N_13974,N_12438,N_12912);
or U13975 (N_13975,N_12970,N_12867);
nand U13976 (N_13976,N_12932,N_12039);
and U13977 (N_13977,N_12423,N_12620);
and U13978 (N_13978,N_12508,N_12998);
and U13979 (N_13979,N_12880,N_12283);
and U13980 (N_13980,N_12167,N_12124);
or U13981 (N_13981,N_12296,N_12391);
nor U13982 (N_13982,N_12033,N_12342);
nand U13983 (N_13983,N_12778,N_12369);
nor U13984 (N_13984,N_12362,N_12336);
and U13985 (N_13985,N_12861,N_12814);
nand U13986 (N_13986,N_12351,N_12783);
xnor U13987 (N_13987,N_12249,N_12925);
nor U13988 (N_13988,N_12010,N_12432);
and U13989 (N_13989,N_12534,N_12884);
nor U13990 (N_13990,N_12850,N_12593);
nor U13991 (N_13991,N_12711,N_12969);
xnor U13992 (N_13992,N_12804,N_12500);
nor U13993 (N_13993,N_12767,N_12207);
and U13994 (N_13994,N_12637,N_12834);
and U13995 (N_13995,N_12431,N_12281);
and U13996 (N_13996,N_12343,N_12374);
nand U13997 (N_13997,N_12649,N_12225);
and U13998 (N_13998,N_12926,N_12884);
xnor U13999 (N_13999,N_12988,N_12289);
nor U14000 (N_14000,N_13072,N_13176);
or U14001 (N_14001,N_13167,N_13573);
nand U14002 (N_14002,N_13878,N_13467);
nor U14003 (N_14003,N_13985,N_13171);
and U14004 (N_14004,N_13928,N_13858);
nand U14005 (N_14005,N_13016,N_13104);
and U14006 (N_14006,N_13914,N_13463);
and U14007 (N_14007,N_13099,N_13163);
nand U14008 (N_14008,N_13220,N_13863);
nor U14009 (N_14009,N_13867,N_13379);
nand U14010 (N_14010,N_13081,N_13014);
nand U14011 (N_14011,N_13726,N_13101);
nor U14012 (N_14012,N_13635,N_13653);
or U14013 (N_14013,N_13775,N_13260);
nor U14014 (N_14014,N_13699,N_13695);
xnor U14015 (N_14015,N_13901,N_13701);
xnor U14016 (N_14016,N_13918,N_13788);
nor U14017 (N_14017,N_13694,N_13668);
nand U14018 (N_14018,N_13426,N_13462);
nor U14019 (N_14019,N_13307,N_13091);
and U14020 (N_14020,N_13690,N_13142);
nor U14021 (N_14021,N_13786,N_13905);
nand U14022 (N_14022,N_13980,N_13283);
and U14023 (N_14023,N_13444,N_13195);
nand U14024 (N_14024,N_13006,N_13616);
nand U14025 (N_14025,N_13951,N_13380);
and U14026 (N_14026,N_13738,N_13080);
or U14027 (N_14027,N_13231,N_13923);
or U14028 (N_14028,N_13249,N_13355);
and U14029 (N_14029,N_13100,N_13465);
nor U14030 (N_14030,N_13737,N_13636);
nor U14031 (N_14031,N_13791,N_13102);
nor U14032 (N_14032,N_13145,N_13671);
nand U14033 (N_14033,N_13257,N_13489);
and U14034 (N_14034,N_13531,N_13178);
and U14035 (N_14035,N_13766,N_13261);
and U14036 (N_14036,N_13621,N_13057);
nand U14037 (N_14037,N_13446,N_13326);
nor U14038 (N_14038,N_13772,N_13764);
or U14039 (N_14039,N_13824,N_13857);
and U14040 (N_14040,N_13188,N_13069);
nor U14041 (N_14041,N_13957,N_13480);
nor U14042 (N_14042,N_13950,N_13181);
nand U14043 (N_14043,N_13973,N_13684);
and U14044 (N_14044,N_13812,N_13902);
nor U14045 (N_14045,N_13472,N_13817);
and U14046 (N_14046,N_13855,N_13981);
and U14047 (N_14047,N_13744,N_13784);
xnor U14048 (N_14048,N_13953,N_13998);
xnor U14049 (N_14049,N_13316,N_13344);
and U14050 (N_14050,N_13753,N_13849);
nor U14051 (N_14051,N_13656,N_13606);
xnor U14052 (N_14052,N_13043,N_13797);
or U14053 (N_14053,N_13956,N_13023);
and U14054 (N_14054,N_13537,N_13510);
or U14055 (N_14055,N_13652,N_13230);
nor U14056 (N_14056,N_13036,N_13556);
nand U14057 (N_14057,N_13443,N_13946);
and U14058 (N_14058,N_13093,N_13209);
nand U14059 (N_14059,N_13810,N_13869);
nand U14060 (N_14060,N_13938,N_13617);
nor U14061 (N_14061,N_13292,N_13280);
and U14062 (N_14062,N_13777,N_13172);
nand U14063 (N_14063,N_13708,N_13148);
nand U14064 (N_14064,N_13174,N_13053);
or U14065 (N_14065,N_13854,N_13034);
or U14066 (N_14066,N_13245,N_13755);
nand U14067 (N_14067,N_13440,N_13015);
nor U14068 (N_14068,N_13763,N_13890);
xor U14069 (N_14069,N_13376,N_13156);
or U14070 (N_14070,N_13021,N_13412);
and U14071 (N_14071,N_13113,N_13235);
or U14072 (N_14072,N_13612,N_13525);
nand U14073 (N_14073,N_13203,N_13648);
and U14074 (N_14074,N_13494,N_13182);
nor U14075 (N_14075,N_13927,N_13720);
or U14076 (N_14076,N_13602,N_13765);
nand U14077 (N_14077,N_13128,N_13536);
and U14078 (N_14078,N_13618,N_13975);
and U14079 (N_14079,N_13555,N_13448);
or U14080 (N_14080,N_13518,N_13868);
and U14081 (N_14081,N_13255,N_13248);
nand U14082 (N_14082,N_13563,N_13048);
nor U14083 (N_14083,N_13627,N_13825);
nor U14084 (N_14084,N_13971,N_13592);
and U14085 (N_14085,N_13962,N_13466);
nand U14086 (N_14086,N_13075,N_13453);
nand U14087 (N_14087,N_13157,N_13488);
xnor U14088 (N_14088,N_13153,N_13709);
nor U14089 (N_14089,N_13512,N_13007);
nor U14090 (N_14090,N_13915,N_13207);
nand U14091 (N_14091,N_13013,N_13793);
or U14092 (N_14092,N_13364,N_13175);
and U14093 (N_14093,N_13374,N_13277);
xor U14094 (N_14094,N_13809,N_13143);
nand U14095 (N_14095,N_13588,N_13638);
and U14096 (N_14096,N_13524,N_13187);
and U14097 (N_14097,N_13967,N_13136);
nand U14098 (N_14098,N_13345,N_13286);
or U14099 (N_14099,N_13437,N_13039);
or U14100 (N_14100,N_13986,N_13820);
xor U14101 (N_14101,N_13404,N_13441);
nand U14102 (N_14102,N_13900,N_13632);
nor U14103 (N_14103,N_13599,N_13945);
and U14104 (N_14104,N_13415,N_13598);
or U14105 (N_14105,N_13949,N_13146);
or U14106 (N_14106,N_13659,N_13089);
or U14107 (N_14107,N_13138,N_13680);
nand U14108 (N_14108,N_13503,N_13672);
and U14109 (N_14109,N_13217,N_13803);
and U14110 (N_14110,N_13582,N_13645);
and U14111 (N_14111,N_13562,N_13071);
or U14112 (N_14112,N_13881,N_13430);
nand U14113 (N_14113,N_13508,N_13743);
and U14114 (N_14114,N_13455,N_13523);
nor U14115 (N_14115,N_13271,N_13700);
xor U14116 (N_14116,N_13999,N_13916);
nand U14117 (N_14117,N_13169,N_13578);
or U14118 (N_14118,N_13078,N_13432);
nand U14119 (N_14119,N_13600,N_13974);
nand U14120 (N_14120,N_13517,N_13377);
nand U14121 (N_14121,N_13527,N_13968);
nor U14122 (N_14122,N_13657,N_13875);
nor U14123 (N_14123,N_13164,N_13162);
and U14124 (N_14124,N_13533,N_13068);
xor U14125 (N_14125,N_13678,N_13689);
nand U14126 (N_14126,N_13633,N_13514);
nor U14127 (N_14127,N_13540,N_13077);
xnor U14128 (N_14128,N_13276,N_13674);
nand U14129 (N_14129,N_13628,N_13387);
nor U14130 (N_14130,N_13827,N_13543);
nand U14131 (N_14131,N_13464,N_13239);
and U14132 (N_14132,N_13196,N_13692);
nor U14133 (N_14133,N_13392,N_13356);
and U14134 (N_14134,N_13870,N_13570);
nor U14135 (N_14135,N_13714,N_13227);
xor U14136 (N_14136,N_13879,N_13587);
and U14137 (N_14137,N_13400,N_13368);
nand U14138 (N_14138,N_13579,N_13816);
or U14139 (N_14139,N_13988,N_13213);
xor U14140 (N_14140,N_13724,N_13727);
or U14141 (N_14141,N_13076,N_13808);
or U14142 (N_14142,N_13389,N_13688);
and U14143 (N_14143,N_13240,N_13061);
nand U14144 (N_14144,N_13740,N_13650);
nor U14145 (N_14145,N_13995,N_13409);
nor U14146 (N_14146,N_13212,N_13427);
nor U14147 (N_14147,N_13484,N_13353);
or U14148 (N_14148,N_13572,N_13060);
nand U14149 (N_14149,N_13112,N_13906);
nand U14150 (N_14150,N_13780,N_13848);
or U14151 (N_14151,N_13940,N_13521);
or U14152 (N_14152,N_13746,N_13917);
nand U14153 (N_14153,N_13574,N_13776);
and U14154 (N_14154,N_13913,N_13712);
nor U14155 (N_14155,N_13044,N_13370);
and U14156 (N_14156,N_13706,N_13086);
xnor U14157 (N_14157,N_13530,N_13329);
and U14158 (N_14158,N_13752,N_13711);
nor U14159 (N_14159,N_13228,N_13046);
nand U14160 (N_14160,N_13384,N_13482);
xnor U14161 (N_14161,N_13281,N_13982);
nor U14162 (N_14162,N_13256,N_13681);
and U14163 (N_14163,N_13095,N_13305);
or U14164 (N_14164,N_13876,N_13019);
nor U14165 (N_14165,N_13954,N_13382);
and U14166 (N_14166,N_13568,N_13017);
and U14167 (N_14167,N_13054,N_13223);
or U14168 (N_14168,N_13383,N_13126);
nor U14169 (N_14169,N_13114,N_13047);
xnor U14170 (N_14170,N_13334,N_13130);
and U14171 (N_14171,N_13972,N_13544);
xnor U14172 (N_14172,N_13522,N_13559);
nand U14173 (N_14173,N_13297,N_13904);
nand U14174 (N_14174,N_13566,N_13070);
nand U14175 (N_14175,N_13815,N_13147);
and U14176 (N_14176,N_13894,N_13924);
and U14177 (N_14177,N_13087,N_13272);
nor U14178 (N_14178,N_13651,N_13375);
xnor U14179 (N_14179,N_13042,N_13670);
nand U14180 (N_14180,N_13590,N_13832);
nor U14181 (N_14181,N_13614,N_13330);
and U14182 (N_14182,N_13964,N_13736);
xnor U14183 (N_14183,N_13603,N_13251);
nand U14184 (N_14184,N_13634,N_13677);
nand U14185 (N_14185,N_13492,N_13381);
and U14186 (N_14186,N_13713,N_13702);
nor U14187 (N_14187,N_13921,N_13298);
and U14188 (N_14188,N_13507,N_13885);
and U14189 (N_14189,N_13862,N_13996);
nor U14190 (N_14190,N_13760,N_13253);
and U14191 (N_14191,N_13269,N_13168);
or U14192 (N_14192,N_13367,N_13605);
nand U14193 (N_14193,N_13360,N_13408);
xor U14194 (N_14194,N_13205,N_13004);
nor U14195 (N_14195,N_13654,N_13853);
nand U14196 (N_14196,N_13515,N_13177);
nor U14197 (N_14197,N_13796,N_13058);
nand U14198 (N_14198,N_13062,N_13667);
nor U14199 (N_14199,N_13293,N_13122);
or U14200 (N_14200,N_13378,N_13411);
or U14201 (N_14201,N_13748,N_13696);
and U14202 (N_14202,N_13675,N_13139);
xor U14203 (N_14203,N_13703,N_13872);
nor U14204 (N_14204,N_13770,N_13655);
and U14205 (N_14205,N_13350,N_13557);
and U14206 (N_14206,N_13939,N_13871);
nor U14207 (N_14207,N_13814,N_13313);
or U14208 (N_14208,N_13718,N_13561);
and U14209 (N_14209,N_13020,N_13351);
nor U14210 (N_14210,N_13247,N_13424);
nor U14211 (N_14211,N_13179,N_13641);
nand U14212 (N_14212,N_13640,N_13476);
and U14213 (N_14213,N_13050,N_13545);
nor U14214 (N_14214,N_13516,N_13813);
and U14215 (N_14215,N_13026,N_13798);
and U14216 (N_14216,N_13952,N_13073);
xnor U14217 (N_14217,N_13622,N_13742);
nand U14218 (N_14218,N_13850,N_13541);
and U14219 (N_14219,N_13989,N_13390);
nor U14220 (N_14220,N_13098,N_13421);
xor U14221 (N_14221,N_13500,N_13719);
nand U14222 (N_14222,N_13338,N_13941);
and U14223 (N_14223,N_13843,N_13229);
and U14224 (N_14224,N_13059,N_13647);
and U14225 (N_14225,N_13417,N_13201);
nor U14226 (N_14226,N_13761,N_13586);
nor U14227 (N_14227,N_13236,N_13639);
or U14228 (N_14228,N_13083,N_13001);
or U14229 (N_14229,N_13925,N_13420);
or U14230 (N_14230,N_13238,N_13274);
nor U14231 (N_14231,N_13210,N_13082);
nand U14232 (N_14232,N_13133,N_13535);
nor U14233 (N_14233,N_13216,N_13513);
nor U14234 (N_14234,N_13342,N_13221);
or U14235 (N_14235,N_13486,N_13722);
nor U14236 (N_14236,N_13037,N_13581);
or U14237 (N_14237,N_13747,N_13434);
or U14238 (N_14238,N_13856,N_13629);
nor U14239 (N_14239,N_13285,N_13698);
nand U14240 (N_14240,N_13140,N_13830);
nor U14241 (N_14241,N_13222,N_13977);
nor U14242 (N_14242,N_13357,N_13937);
or U14243 (N_14243,N_13154,N_13790);
xor U14244 (N_14244,N_13644,N_13040);
or U14245 (N_14245,N_13505,N_13189);
xnor U14246 (N_14246,N_13385,N_13859);
and U14247 (N_14247,N_13926,N_13135);
xor U14248 (N_14248,N_13301,N_13252);
or U14249 (N_14249,N_13929,N_13309);
nor U14250 (N_14250,N_13308,N_13822);
or U14251 (N_14251,N_13818,N_13837);
nand U14252 (N_14252,N_13451,N_13150);
nor U14253 (N_14253,N_13284,N_13243);
or U14254 (N_14254,N_13619,N_13932);
nor U14255 (N_14255,N_13388,N_13435);
nand U14256 (N_14256,N_13294,N_13686);
nand U14257 (N_14257,N_13456,N_13646);
xor U14258 (N_14258,N_13774,N_13922);
nand U14259 (N_14259,N_13406,N_13413);
xor U14260 (N_14260,N_13802,N_13733);
nor U14261 (N_14261,N_13085,N_13771);
xnor U14262 (N_14262,N_13845,N_13767);
or U14263 (N_14263,N_13232,N_13613);
nand U14264 (N_14264,N_13109,N_13643);
nor U14265 (N_14265,N_13852,N_13275);
nor U14266 (N_14266,N_13960,N_13707);
xor U14267 (N_14267,N_13299,N_13200);
or U14268 (N_14268,N_13961,N_13027);
nand U14269 (N_14269,N_13219,N_13834);
or U14270 (N_14270,N_13642,N_13314);
or U14271 (N_14271,N_13165,N_13237);
and U14272 (N_14272,N_13436,N_13593);
and U14273 (N_14273,N_13679,N_13637);
or U14274 (N_14274,N_13288,N_13410);
nor U14275 (N_14275,N_13211,N_13778);
or U14276 (N_14276,N_13501,N_13754);
nand U14277 (N_14277,N_13829,N_13161);
nor U14278 (N_14278,N_13403,N_13963);
and U14279 (N_14279,N_13729,N_13429);
xor U14280 (N_14280,N_13012,N_13206);
and U14281 (N_14281,N_13511,N_13401);
or U14282 (N_14282,N_13439,N_13886);
xnor U14283 (N_14283,N_13250,N_13458);
xnor U14284 (N_14284,N_13107,N_13584);
or U14285 (N_14285,N_13880,N_13475);
or U14286 (N_14286,N_13631,N_13947);
xnor U14287 (N_14287,N_13395,N_13123);
or U14288 (N_14288,N_13282,N_13558);
xnor U14289 (N_14289,N_13805,N_13315);
and U14290 (N_14290,N_13844,N_13959);
nor U14291 (N_14291,N_13811,N_13676);
nand U14292 (N_14292,N_13225,N_13341);
and U14293 (N_14293,N_13477,N_13660);
xnor U14294 (N_14294,N_13839,N_13550);
nand U14295 (N_14295,N_13129,N_13366);
and U14296 (N_14296,N_13337,N_13860);
nor U14297 (N_14297,N_13673,N_13149);
xnor U14298 (N_14298,N_13666,N_13504);
and U14299 (N_14299,N_13576,N_13152);
or U14300 (N_14300,N_13866,N_13358);
and U14301 (N_14301,N_13608,N_13897);
and U14302 (N_14302,N_13625,N_13317);
nand U14303 (N_14303,N_13710,N_13549);
nor U14304 (N_14304,N_13892,N_13166);
nand U14305 (N_14305,N_13359,N_13262);
nand U14306 (N_14306,N_13910,N_13116);
nand U14307 (N_14307,N_13496,N_13433);
nor U14308 (N_14308,N_13214,N_13571);
xor U14309 (N_14309,N_13009,N_13131);
nor U14310 (N_14310,N_13396,N_13090);
nand U14311 (N_14311,N_13662,N_13155);
nor U14312 (N_14312,N_13615,N_13033);
or U14313 (N_14313,N_13903,N_13197);
or U14314 (N_14314,N_13597,N_13851);
xor U14315 (N_14315,N_13198,N_13296);
xnor U14316 (N_14316,N_13762,N_13891);
nand U14317 (N_14317,N_13984,N_13721);
xnor U14318 (N_14318,N_13041,N_13028);
nor U14319 (N_14319,N_13741,N_13226);
nor U14320 (N_14320,N_13942,N_13993);
nor U14321 (N_14321,N_13399,N_13056);
nor U14322 (N_14322,N_13506,N_13369);
and U14323 (N_14323,N_13119,N_13490);
nor U14324 (N_14324,N_13626,N_13750);
and U14325 (N_14325,N_13691,N_13785);
nor U14326 (N_14326,N_13978,N_13474);
nand U14327 (N_14327,N_13425,N_13199);
or U14328 (N_14328,N_13819,N_13528);
nor U14329 (N_14329,N_13783,N_13723);
xor U14330 (N_14330,N_13567,N_13121);
nor U14331 (N_14331,N_13287,N_13279);
nand U14332 (N_14332,N_13454,N_13705);
or U14333 (N_14333,N_13547,N_13186);
nor U14334 (N_14334,N_13336,N_13717);
and U14335 (N_14335,N_13170,N_13664);
or U14336 (N_14336,N_13318,N_13920);
and U14337 (N_14337,N_13273,N_13526);
and U14338 (N_14338,N_13029,N_13704);
or U14339 (N_14339,N_13888,N_13609);
and U14340 (N_14340,N_13185,N_13883);
and U14341 (N_14341,N_13930,N_13063);
nand U14342 (N_14342,N_13304,N_13473);
or U14343 (N_14343,N_13779,N_13184);
and U14344 (N_14344,N_13983,N_13665);
and U14345 (N_14345,N_13335,N_13663);
or U14346 (N_14346,N_13332,N_13265);
nand U14347 (N_14347,N_13934,N_13111);
and U14348 (N_14348,N_13303,N_13716);
nor U14349 (N_14349,N_13291,N_13327);
nand U14350 (N_14350,N_13661,N_13328);
nand U14351 (N_14351,N_13339,N_13757);
and U14352 (N_14352,N_13539,N_13936);
nor U14353 (N_14353,N_13290,N_13173);
xnor U14354 (N_14354,N_13751,N_13127);
or U14355 (N_14355,N_13005,N_13944);
or U14356 (N_14356,N_13577,N_13895);
and U14357 (N_14357,N_13589,N_13349);
xnor U14358 (N_14358,N_13320,N_13120);
nand U14359 (N_14359,N_13117,N_13519);
and U14360 (N_14360,N_13487,N_13909);
nor U14361 (N_14361,N_13066,N_13097);
nand U14362 (N_14362,N_13180,N_13846);
or U14363 (N_14363,N_13781,N_13452);
xnor U14364 (N_14364,N_13580,N_13397);
nand U14365 (N_14365,N_13244,N_13354);
or U14366 (N_14366,N_13835,N_13493);
nand U14367 (N_14367,N_13792,N_13838);
or U14368 (N_14368,N_13191,N_13624);
xor U14369 (N_14369,N_13534,N_13365);
nor U14370 (N_14370,N_13758,N_13125);
and U14371 (N_14371,N_13051,N_13302);
nor U14372 (N_14372,N_13300,N_13734);
and U14373 (N_14373,N_13943,N_13363);
nand U14374 (N_14374,N_13595,N_13144);
nor U14375 (N_14375,N_13479,N_13782);
or U14376 (N_14376,N_13030,N_13509);
nand U14377 (N_14377,N_13575,N_13884);
nor U14378 (N_14378,N_13485,N_13735);
and U14379 (N_14379,N_13976,N_13134);
nand U14380 (N_14380,N_13491,N_13874);
nor U14381 (N_14381,N_13789,N_13343);
and U14382 (N_14382,N_13052,N_13324);
and U14383 (N_14383,N_13459,N_13987);
or U14384 (N_14384,N_13495,N_13604);
xnor U14385 (N_14385,N_13032,N_13630);
nand U14386 (N_14386,N_13442,N_13003);
and U14387 (N_14387,N_13732,N_13074);
and U14388 (N_14388,N_13428,N_13794);
nand U14389 (N_14389,N_13997,N_13124);
and U14390 (N_14390,N_13478,N_13769);
or U14391 (N_14391,N_13450,N_13067);
and U14392 (N_14392,N_13800,N_13088);
nand U14393 (N_14393,N_13192,N_13554);
and U14394 (N_14394,N_13414,N_13548);
nand U14395 (N_14395,N_13045,N_13552);
nand U14396 (N_14396,N_13969,N_13160);
and U14397 (N_14397,N_13683,N_13725);
and U14398 (N_14398,N_13049,N_13911);
or U14399 (N_14399,N_13105,N_13931);
nor U14400 (N_14400,N_13799,N_13730);
and U14401 (N_14401,N_13669,N_13224);
nand U14402 (N_14402,N_13268,N_13873);
or U14403 (N_14403,N_13898,N_13907);
nand U14404 (N_14404,N_13979,N_13094);
xnor U14405 (N_14405,N_13546,N_13000);
xnor U14406 (N_14406,N_13394,N_13241);
nor U14407 (N_14407,N_13687,N_13319);
nor U14408 (N_14408,N_13110,N_13011);
or U14409 (N_14409,N_13591,N_13965);
nand U14410 (N_14410,N_13266,N_13826);
or U14411 (N_14411,N_13398,N_13118);
or U14412 (N_14412,N_13865,N_13115);
nor U14413 (N_14413,N_13682,N_13233);
or U14414 (N_14414,N_13759,N_13151);
nand U14415 (N_14415,N_13215,N_13407);
nand U14416 (N_14416,N_13352,N_13594);
xor U14417 (N_14417,N_13502,N_13306);
nor U14418 (N_14418,N_13468,N_13106);
nor U14419 (N_14419,N_13333,N_13312);
and U14420 (N_14420,N_13481,N_13560);
nor U14421 (N_14421,N_13348,N_13419);
and U14422 (N_14422,N_13623,N_13542);
nor U14423 (N_14423,N_13731,N_13806);
nor U14424 (N_14424,N_13994,N_13393);
or U14425 (N_14425,N_13532,N_13295);
and U14426 (N_14426,N_13569,N_13096);
nor U14427 (N_14427,N_13749,N_13877);
and U14428 (N_14428,N_13137,N_13035);
nor U14429 (N_14429,N_13190,N_13202);
nor U14430 (N_14430,N_13831,N_13899);
xor U14431 (N_14431,N_13372,N_13064);
and U14432 (N_14432,N_13431,N_13254);
or U14433 (N_14433,N_13234,N_13310);
or U14434 (N_14434,N_13861,N_13084);
nand U14435 (N_14435,N_13193,N_13361);
nor U14436 (N_14436,N_13025,N_13847);
nand U14437 (N_14437,N_13728,N_13919);
or U14438 (N_14438,N_13801,N_13218);
nand U14439 (N_14439,N_13499,N_13990);
xor U14440 (N_14440,N_13325,N_13323);
and U14441 (N_14441,N_13912,N_13159);
nor U14442 (N_14442,N_13773,N_13264);
nor U14443 (N_14443,N_13620,N_13322);
and U14444 (N_14444,N_13079,N_13371);
and U14445 (N_14445,N_13896,N_13821);
and U14446 (N_14446,N_13787,N_13024);
xnor U14447 (N_14447,N_13208,N_13108);
nand U14448 (N_14448,N_13311,N_13373);
xnor U14449 (N_14449,N_13887,N_13055);
nand U14450 (N_14450,N_13565,N_13457);
nand U14451 (N_14451,N_13242,N_13804);
xnor U14452 (N_14452,N_13611,N_13183);
and U14453 (N_14453,N_13970,N_13795);
nor U14454 (N_14454,N_13889,N_13422);
nand U14455 (N_14455,N_13649,N_13610);
or U14456 (N_14456,N_13948,N_13445);
nor U14457 (N_14457,N_13693,N_13418);
and U14458 (N_14458,N_13447,N_13391);
nor U14459 (N_14459,N_13278,N_13258);
nor U14460 (N_14460,N_13461,N_13022);
and U14461 (N_14461,N_13460,N_13132);
nand U14462 (N_14462,N_13893,N_13347);
and U14463 (N_14463,N_13259,N_13715);
or U14464 (N_14464,N_13520,N_13828);
nand U14465 (N_14465,N_13038,N_13010);
nand U14466 (N_14466,N_13103,N_13346);
or U14467 (N_14467,N_13194,N_13841);
or U14468 (N_14468,N_13002,N_13992);
or U14469 (N_14469,N_13263,N_13018);
nand U14470 (N_14470,N_13497,N_13483);
and U14471 (N_14471,N_13416,N_13933);
and U14472 (N_14472,N_13966,N_13538);
or U14473 (N_14473,N_13955,N_13842);
nand U14474 (N_14474,N_13469,N_13362);
nand U14475 (N_14475,N_13658,N_13423);
and U14476 (N_14476,N_13158,N_13470);
or U14477 (N_14477,N_13340,N_13596);
or U14478 (N_14478,N_13289,N_13270);
nor U14479 (N_14479,N_13141,N_13697);
or U14480 (N_14480,N_13498,N_13756);
nand U14481 (N_14481,N_13551,N_13768);
nor U14482 (N_14482,N_13601,N_13438);
and U14483 (N_14483,N_13065,N_13991);
or U14484 (N_14484,N_13267,N_13331);
nand U14485 (N_14485,N_13405,N_13739);
and U14486 (N_14486,N_13607,N_13833);
or U14487 (N_14487,N_13092,N_13321);
nand U14488 (N_14488,N_13908,N_13204);
xor U14489 (N_14489,N_13958,N_13745);
or U14490 (N_14490,N_13008,N_13882);
nand U14491 (N_14491,N_13553,N_13583);
or U14492 (N_14492,N_13685,N_13807);
and U14493 (N_14493,N_13935,N_13585);
and U14494 (N_14494,N_13246,N_13402);
xor U14495 (N_14495,N_13823,N_13471);
nand U14496 (N_14496,N_13864,N_13840);
nand U14497 (N_14497,N_13836,N_13449);
and U14498 (N_14498,N_13031,N_13386);
nor U14499 (N_14499,N_13564,N_13529);
nand U14500 (N_14500,N_13860,N_13750);
nand U14501 (N_14501,N_13406,N_13128);
nor U14502 (N_14502,N_13176,N_13016);
or U14503 (N_14503,N_13614,N_13048);
xnor U14504 (N_14504,N_13395,N_13142);
or U14505 (N_14505,N_13045,N_13589);
xor U14506 (N_14506,N_13449,N_13074);
and U14507 (N_14507,N_13252,N_13247);
or U14508 (N_14508,N_13064,N_13084);
or U14509 (N_14509,N_13423,N_13446);
nand U14510 (N_14510,N_13016,N_13981);
nand U14511 (N_14511,N_13514,N_13753);
xnor U14512 (N_14512,N_13520,N_13370);
xor U14513 (N_14513,N_13791,N_13017);
nor U14514 (N_14514,N_13546,N_13360);
nand U14515 (N_14515,N_13593,N_13456);
and U14516 (N_14516,N_13695,N_13200);
nor U14517 (N_14517,N_13896,N_13904);
or U14518 (N_14518,N_13042,N_13703);
or U14519 (N_14519,N_13876,N_13995);
nor U14520 (N_14520,N_13952,N_13541);
or U14521 (N_14521,N_13340,N_13909);
nor U14522 (N_14522,N_13699,N_13245);
or U14523 (N_14523,N_13772,N_13680);
nor U14524 (N_14524,N_13865,N_13511);
nand U14525 (N_14525,N_13528,N_13628);
nor U14526 (N_14526,N_13095,N_13195);
nand U14527 (N_14527,N_13327,N_13487);
nand U14528 (N_14528,N_13809,N_13368);
or U14529 (N_14529,N_13970,N_13725);
nand U14530 (N_14530,N_13809,N_13444);
nor U14531 (N_14531,N_13994,N_13202);
and U14532 (N_14532,N_13555,N_13841);
nor U14533 (N_14533,N_13291,N_13735);
or U14534 (N_14534,N_13773,N_13858);
and U14535 (N_14535,N_13307,N_13309);
nand U14536 (N_14536,N_13275,N_13382);
and U14537 (N_14537,N_13615,N_13747);
and U14538 (N_14538,N_13226,N_13724);
or U14539 (N_14539,N_13748,N_13263);
xnor U14540 (N_14540,N_13532,N_13315);
or U14541 (N_14541,N_13999,N_13295);
nor U14542 (N_14542,N_13558,N_13670);
nand U14543 (N_14543,N_13190,N_13395);
nand U14544 (N_14544,N_13710,N_13900);
nand U14545 (N_14545,N_13808,N_13251);
and U14546 (N_14546,N_13416,N_13547);
xnor U14547 (N_14547,N_13772,N_13969);
nor U14548 (N_14548,N_13372,N_13435);
and U14549 (N_14549,N_13993,N_13342);
or U14550 (N_14550,N_13267,N_13125);
or U14551 (N_14551,N_13494,N_13469);
and U14552 (N_14552,N_13852,N_13513);
or U14553 (N_14553,N_13719,N_13993);
xnor U14554 (N_14554,N_13119,N_13235);
nor U14555 (N_14555,N_13513,N_13034);
and U14556 (N_14556,N_13077,N_13054);
or U14557 (N_14557,N_13253,N_13716);
or U14558 (N_14558,N_13068,N_13227);
and U14559 (N_14559,N_13582,N_13410);
nand U14560 (N_14560,N_13647,N_13167);
nor U14561 (N_14561,N_13946,N_13907);
nor U14562 (N_14562,N_13134,N_13652);
nand U14563 (N_14563,N_13228,N_13118);
nand U14564 (N_14564,N_13642,N_13679);
nor U14565 (N_14565,N_13775,N_13091);
nor U14566 (N_14566,N_13290,N_13157);
and U14567 (N_14567,N_13420,N_13028);
or U14568 (N_14568,N_13833,N_13261);
nor U14569 (N_14569,N_13475,N_13294);
nor U14570 (N_14570,N_13803,N_13778);
xnor U14571 (N_14571,N_13947,N_13165);
nor U14572 (N_14572,N_13756,N_13893);
nand U14573 (N_14573,N_13776,N_13414);
nand U14574 (N_14574,N_13902,N_13302);
nor U14575 (N_14575,N_13349,N_13508);
xor U14576 (N_14576,N_13642,N_13304);
nand U14577 (N_14577,N_13814,N_13485);
nor U14578 (N_14578,N_13183,N_13403);
nor U14579 (N_14579,N_13885,N_13666);
or U14580 (N_14580,N_13171,N_13314);
nand U14581 (N_14581,N_13914,N_13551);
or U14582 (N_14582,N_13523,N_13469);
or U14583 (N_14583,N_13684,N_13865);
nor U14584 (N_14584,N_13412,N_13782);
nand U14585 (N_14585,N_13013,N_13877);
nand U14586 (N_14586,N_13581,N_13819);
and U14587 (N_14587,N_13305,N_13225);
nand U14588 (N_14588,N_13184,N_13774);
or U14589 (N_14589,N_13040,N_13014);
or U14590 (N_14590,N_13293,N_13715);
or U14591 (N_14591,N_13274,N_13747);
nor U14592 (N_14592,N_13637,N_13502);
nand U14593 (N_14593,N_13099,N_13800);
or U14594 (N_14594,N_13758,N_13676);
nand U14595 (N_14595,N_13077,N_13082);
nand U14596 (N_14596,N_13685,N_13703);
or U14597 (N_14597,N_13827,N_13667);
and U14598 (N_14598,N_13215,N_13042);
nor U14599 (N_14599,N_13403,N_13247);
nand U14600 (N_14600,N_13948,N_13341);
or U14601 (N_14601,N_13615,N_13107);
nand U14602 (N_14602,N_13084,N_13629);
xor U14603 (N_14603,N_13141,N_13260);
or U14604 (N_14604,N_13075,N_13877);
or U14605 (N_14605,N_13777,N_13539);
and U14606 (N_14606,N_13404,N_13594);
and U14607 (N_14607,N_13733,N_13940);
xnor U14608 (N_14608,N_13235,N_13613);
and U14609 (N_14609,N_13471,N_13292);
nand U14610 (N_14610,N_13514,N_13923);
nor U14611 (N_14611,N_13987,N_13521);
or U14612 (N_14612,N_13132,N_13908);
and U14613 (N_14613,N_13929,N_13856);
xnor U14614 (N_14614,N_13891,N_13038);
nand U14615 (N_14615,N_13419,N_13605);
nand U14616 (N_14616,N_13618,N_13444);
nor U14617 (N_14617,N_13919,N_13661);
or U14618 (N_14618,N_13677,N_13669);
and U14619 (N_14619,N_13815,N_13659);
nor U14620 (N_14620,N_13443,N_13359);
or U14621 (N_14621,N_13056,N_13665);
and U14622 (N_14622,N_13508,N_13716);
or U14623 (N_14623,N_13425,N_13224);
nor U14624 (N_14624,N_13869,N_13607);
nand U14625 (N_14625,N_13744,N_13656);
and U14626 (N_14626,N_13238,N_13110);
nand U14627 (N_14627,N_13078,N_13210);
or U14628 (N_14628,N_13963,N_13388);
nor U14629 (N_14629,N_13741,N_13828);
xor U14630 (N_14630,N_13783,N_13005);
nand U14631 (N_14631,N_13092,N_13101);
and U14632 (N_14632,N_13503,N_13377);
and U14633 (N_14633,N_13907,N_13090);
nand U14634 (N_14634,N_13903,N_13566);
or U14635 (N_14635,N_13327,N_13514);
nand U14636 (N_14636,N_13269,N_13871);
nand U14637 (N_14637,N_13574,N_13940);
nand U14638 (N_14638,N_13722,N_13648);
nand U14639 (N_14639,N_13851,N_13805);
and U14640 (N_14640,N_13750,N_13343);
nor U14641 (N_14641,N_13204,N_13260);
and U14642 (N_14642,N_13702,N_13622);
nand U14643 (N_14643,N_13034,N_13013);
and U14644 (N_14644,N_13028,N_13251);
and U14645 (N_14645,N_13900,N_13085);
nor U14646 (N_14646,N_13100,N_13445);
xnor U14647 (N_14647,N_13013,N_13264);
xor U14648 (N_14648,N_13301,N_13010);
and U14649 (N_14649,N_13951,N_13931);
or U14650 (N_14650,N_13465,N_13085);
and U14651 (N_14651,N_13616,N_13636);
or U14652 (N_14652,N_13466,N_13638);
xnor U14653 (N_14653,N_13787,N_13998);
or U14654 (N_14654,N_13495,N_13520);
and U14655 (N_14655,N_13283,N_13822);
xor U14656 (N_14656,N_13953,N_13977);
nor U14657 (N_14657,N_13531,N_13244);
nand U14658 (N_14658,N_13687,N_13593);
xor U14659 (N_14659,N_13123,N_13492);
and U14660 (N_14660,N_13065,N_13649);
and U14661 (N_14661,N_13244,N_13056);
nor U14662 (N_14662,N_13127,N_13204);
xnor U14663 (N_14663,N_13163,N_13046);
or U14664 (N_14664,N_13628,N_13142);
nor U14665 (N_14665,N_13818,N_13732);
xnor U14666 (N_14666,N_13276,N_13453);
nand U14667 (N_14667,N_13653,N_13921);
nand U14668 (N_14668,N_13761,N_13135);
and U14669 (N_14669,N_13160,N_13787);
nor U14670 (N_14670,N_13305,N_13853);
or U14671 (N_14671,N_13081,N_13782);
nor U14672 (N_14672,N_13910,N_13820);
xor U14673 (N_14673,N_13479,N_13361);
and U14674 (N_14674,N_13778,N_13758);
nand U14675 (N_14675,N_13843,N_13823);
nand U14676 (N_14676,N_13005,N_13950);
and U14677 (N_14677,N_13437,N_13297);
or U14678 (N_14678,N_13744,N_13183);
or U14679 (N_14679,N_13190,N_13813);
and U14680 (N_14680,N_13038,N_13964);
and U14681 (N_14681,N_13019,N_13522);
xor U14682 (N_14682,N_13118,N_13975);
nand U14683 (N_14683,N_13874,N_13045);
nand U14684 (N_14684,N_13149,N_13508);
or U14685 (N_14685,N_13578,N_13463);
nand U14686 (N_14686,N_13791,N_13772);
or U14687 (N_14687,N_13151,N_13987);
and U14688 (N_14688,N_13477,N_13445);
nor U14689 (N_14689,N_13593,N_13890);
or U14690 (N_14690,N_13495,N_13419);
nor U14691 (N_14691,N_13393,N_13788);
and U14692 (N_14692,N_13688,N_13921);
and U14693 (N_14693,N_13862,N_13899);
nand U14694 (N_14694,N_13157,N_13091);
xnor U14695 (N_14695,N_13984,N_13433);
nor U14696 (N_14696,N_13012,N_13751);
nand U14697 (N_14697,N_13471,N_13667);
and U14698 (N_14698,N_13015,N_13675);
nor U14699 (N_14699,N_13561,N_13555);
and U14700 (N_14700,N_13500,N_13370);
nor U14701 (N_14701,N_13469,N_13414);
nand U14702 (N_14702,N_13991,N_13362);
nor U14703 (N_14703,N_13309,N_13667);
or U14704 (N_14704,N_13499,N_13914);
xor U14705 (N_14705,N_13496,N_13934);
nor U14706 (N_14706,N_13125,N_13403);
and U14707 (N_14707,N_13647,N_13304);
nor U14708 (N_14708,N_13681,N_13734);
nand U14709 (N_14709,N_13121,N_13199);
or U14710 (N_14710,N_13701,N_13870);
nand U14711 (N_14711,N_13428,N_13382);
xnor U14712 (N_14712,N_13882,N_13941);
and U14713 (N_14713,N_13594,N_13975);
or U14714 (N_14714,N_13827,N_13059);
and U14715 (N_14715,N_13760,N_13941);
nor U14716 (N_14716,N_13360,N_13821);
nor U14717 (N_14717,N_13487,N_13381);
nor U14718 (N_14718,N_13198,N_13348);
nand U14719 (N_14719,N_13114,N_13936);
and U14720 (N_14720,N_13301,N_13952);
and U14721 (N_14721,N_13346,N_13020);
nand U14722 (N_14722,N_13290,N_13881);
nand U14723 (N_14723,N_13582,N_13043);
nand U14724 (N_14724,N_13712,N_13093);
nand U14725 (N_14725,N_13382,N_13595);
nand U14726 (N_14726,N_13118,N_13461);
and U14727 (N_14727,N_13232,N_13739);
nand U14728 (N_14728,N_13624,N_13087);
nand U14729 (N_14729,N_13511,N_13045);
or U14730 (N_14730,N_13395,N_13387);
nand U14731 (N_14731,N_13707,N_13467);
nor U14732 (N_14732,N_13666,N_13843);
and U14733 (N_14733,N_13988,N_13001);
nand U14734 (N_14734,N_13605,N_13543);
nand U14735 (N_14735,N_13831,N_13093);
and U14736 (N_14736,N_13215,N_13242);
nor U14737 (N_14737,N_13477,N_13456);
or U14738 (N_14738,N_13413,N_13521);
or U14739 (N_14739,N_13261,N_13792);
nand U14740 (N_14740,N_13832,N_13574);
nand U14741 (N_14741,N_13162,N_13377);
or U14742 (N_14742,N_13209,N_13592);
nand U14743 (N_14743,N_13000,N_13572);
nor U14744 (N_14744,N_13548,N_13618);
xnor U14745 (N_14745,N_13531,N_13648);
nand U14746 (N_14746,N_13593,N_13447);
nand U14747 (N_14747,N_13337,N_13930);
nor U14748 (N_14748,N_13076,N_13102);
nand U14749 (N_14749,N_13880,N_13167);
or U14750 (N_14750,N_13567,N_13325);
nor U14751 (N_14751,N_13067,N_13373);
or U14752 (N_14752,N_13467,N_13475);
nor U14753 (N_14753,N_13726,N_13949);
nor U14754 (N_14754,N_13974,N_13328);
nand U14755 (N_14755,N_13432,N_13611);
nor U14756 (N_14756,N_13623,N_13226);
and U14757 (N_14757,N_13419,N_13395);
nor U14758 (N_14758,N_13237,N_13460);
or U14759 (N_14759,N_13798,N_13919);
and U14760 (N_14760,N_13752,N_13723);
and U14761 (N_14761,N_13398,N_13170);
nor U14762 (N_14762,N_13559,N_13967);
nor U14763 (N_14763,N_13454,N_13472);
xnor U14764 (N_14764,N_13819,N_13272);
nor U14765 (N_14765,N_13280,N_13897);
nor U14766 (N_14766,N_13963,N_13156);
xnor U14767 (N_14767,N_13087,N_13179);
nor U14768 (N_14768,N_13924,N_13686);
nand U14769 (N_14769,N_13293,N_13393);
nand U14770 (N_14770,N_13468,N_13154);
and U14771 (N_14771,N_13994,N_13183);
nor U14772 (N_14772,N_13422,N_13166);
nand U14773 (N_14773,N_13433,N_13247);
or U14774 (N_14774,N_13771,N_13379);
nor U14775 (N_14775,N_13161,N_13002);
nor U14776 (N_14776,N_13189,N_13932);
xnor U14777 (N_14777,N_13316,N_13260);
nor U14778 (N_14778,N_13050,N_13202);
xnor U14779 (N_14779,N_13367,N_13797);
nand U14780 (N_14780,N_13543,N_13271);
and U14781 (N_14781,N_13476,N_13836);
nand U14782 (N_14782,N_13497,N_13840);
nor U14783 (N_14783,N_13127,N_13598);
or U14784 (N_14784,N_13149,N_13588);
and U14785 (N_14785,N_13005,N_13323);
and U14786 (N_14786,N_13240,N_13045);
nor U14787 (N_14787,N_13964,N_13450);
and U14788 (N_14788,N_13850,N_13625);
and U14789 (N_14789,N_13354,N_13427);
and U14790 (N_14790,N_13024,N_13813);
or U14791 (N_14791,N_13834,N_13318);
and U14792 (N_14792,N_13771,N_13604);
xnor U14793 (N_14793,N_13386,N_13313);
xor U14794 (N_14794,N_13296,N_13148);
and U14795 (N_14795,N_13652,N_13602);
nor U14796 (N_14796,N_13439,N_13212);
nand U14797 (N_14797,N_13686,N_13895);
or U14798 (N_14798,N_13941,N_13200);
nor U14799 (N_14799,N_13398,N_13531);
and U14800 (N_14800,N_13408,N_13596);
and U14801 (N_14801,N_13622,N_13046);
or U14802 (N_14802,N_13347,N_13870);
xnor U14803 (N_14803,N_13472,N_13697);
xnor U14804 (N_14804,N_13292,N_13631);
or U14805 (N_14805,N_13575,N_13188);
or U14806 (N_14806,N_13786,N_13244);
xnor U14807 (N_14807,N_13782,N_13681);
and U14808 (N_14808,N_13588,N_13924);
nor U14809 (N_14809,N_13308,N_13165);
xnor U14810 (N_14810,N_13639,N_13734);
or U14811 (N_14811,N_13941,N_13152);
and U14812 (N_14812,N_13305,N_13633);
nand U14813 (N_14813,N_13768,N_13209);
nand U14814 (N_14814,N_13387,N_13847);
xnor U14815 (N_14815,N_13777,N_13280);
and U14816 (N_14816,N_13545,N_13717);
xnor U14817 (N_14817,N_13962,N_13351);
nor U14818 (N_14818,N_13470,N_13016);
xnor U14819 (N_14819,N_13101,N_13831);
nand U14820 (N_14820,N_13583,N_13926);
nor U14821 (N_14821,N_13359,N_13468);
and U14822 (N_14822,N_13309,N_13576);
nand U14823 (N_14823,N_13244,N_13303);
or U14824 (N_14824,N_13215,N_13217);
xnor U14825 (N_14825,N_13705,N_13945);
nor U14826 (N_14826,N_13003,N_13110);
nand U14827 (N_14827,N_13804,N_13887);
xor U14828 (N_14828,N_13217,N_13600);
nor U14829 (N_14829,N_13974,N_13041);
nand U14830 (N_14830,N_13847,N_13704);
nand U14831 (N_14831,N_13071,N_13594);
nand U14832 (N_14832,N_13934,N_13663);
nand U14833 (N_14833,N_13522,N_13284);
and U14834 (N_14834,N_13781,N_13608);
nand U14835 (N_14835,N_13402,N_13805);
and U14836 (N_14836,N_13944,N_13549);
and U14837 (N_14837,N_13426,N_13312);
nand U14838 (N_14838,N_13955,N_13983);
and U14839 (N_14839,N_13162,N_13813);
or U14840 (N_14840,N_13540,N_13264);
nand U14841 (N_14841,N_13810,N_13546);
or U14842 (N_14842,N_13437,N_13354);
and U14843 (N_14843,N_13026,N_13645);
and U14844 (N_14844,N_13730,N_13484);
or U14845 (N_14845,N_13202,N_13004);
and U14846 (N_14846,N_13406,N_13356);
and U14847 (N_14847,N_13533,N_13134);
or U14848 (N_14848,N_13909,N_13331);
and U14849 (N_14849,N_13280,N_13827);
nor U14850 (N_14850,N_13013,N_13684);
or U14851 (N_14851,N_13639,N_13778);
or U14852 (N_14852,N_13219,N_13938);
or U14853 (N_14853,N_13572,N_13787);
nand U14854 (N_14854,N_13724,N_13037);
or U14855 (N_14855,N_13337,N_13233);
nand U14856 (N_14856,N_13119,N_13584);
xor U14857 (N_14857,N_13997,N_13767);
nor U14858 (N_14858,N_13012,N_13514);
or U14859 (N_14859,N_13972,N_13889);
or U14860 (N_14860,N_13256,N_13793);
and U14861 (N_14861,N_13121,N_13057);
nor U14862 (N_14862,N_13424,N_13951);
or U14863 (N_14863,N_13301,N_13334);
or U14864 (N_14864,N_13878,N_13541);
nand U14865 (N_14865,N_13169,N_13937);
and U14866 (N_14866,N_13572,N_13991);
nor U14867 (N_14867,N_13923,N_13484);
nor U14868 (N_14868,N_13077,N_13295);
and U14869 (N_14869,N_13264,N_13796);
nand U14870 (N_14870,N_13943,N_13463);
nor U14871 (N_14871,N_13360,N_13893);
nor U14872 (N_14872,N_13467,N_13543);
or U14873 (N_14873,N_13384,N_13194);
and U14874 (N_14874,N_13299,N_13402);
nand U14875 (N_14875,N_13350,N_13669);
and U14876 (N_14876,N_13189,N_13993);
xnor U14877 (N_14877,N_13276,N_13747);
and U14878 (N_14878,N_13298,N_13074);
and U14879 (N_14879,N_13867,N_13741);
nor U14880 (N_14880,N_13531,N_13280);
nand U14881 (N_14881,N_13871,N_13539);
xor U14882 (N_14882,N_13532,N_13145);
and U14883 (N_14883,N_13175,N_13517);
and U14884 (N_14884,N_13809,N_13113);
or U14885 (N_14885,N_13858,N_13207);
or U14886 (N_14886,N_13872,N_13977);
or U14887 (N_14887,N_13493,N_13818);
nand U14888 (N_14888,N_13366,N_13919);
and U14889 (N_14889,N_13884,N_13496);
nand U14890 (N_14890,N_13879,N_13276);
and U14891 (N_14891,N_13904,N_13457);
and U14892 (N_14892,N_13873,N_13904);
nor U14893 (N_14893,N_13365,N_13332);
and U14894 (N_14894,N_13349,N_13989);
and U14895 (N_14895,N_13323,N_13622);
and U14896 (N_14896,N_13913,N_13953);
and U14897 (N_14897,N_13245,N_13435);
nor U14898 (N_14898,N_13956,N_13721);
or U14899 (N_14899,N_13229,N_13727);
nand U14900 (N_14900,N_13335,N_13652);
nor U14901 (N_14901,N_13305,N_13894);
or U14902 (N_14902,N_13957,N_13630);
nor U14903 (N_14903,N_13281,N_13087);
and U14904 (N_14904,N_13144,N_13934);
or U14905 (N_14905,N_13519,N_13748);
xnor U14906 (N_14906,N_13329,N_13963);
or U14907 (N_14907,N_13396,N_13415);
nor U14908 (N_14908,N_13854,N_13525);
or U14909 (N_14909,N_13028,N_13166);
nor U14910 (N_14910,N_13234,N_13995);
or U14911 (N_14911,N_13517,N_13991);
or U14912 (N_14912,N_13618,N_13149);
and U14913 (N_14913,N_13648,N_13428);
or U14914 (N_14914,N_13965,N_13539);
nor U14915 (N_14915,N_13855,N_13561);
and U14916 (N_14916,N_13733,N_13482);
nor U14917 (N_14917,N_13206,N_13340);
and U14918 (N_14918,N_13465,N_13062);
or U14919 (N_14919,N_13883,N_13461);
nand U14920 (N_14920,N_13236,N_13448);
or U14921 (N_14921,N_13911,N_13094);
nor U14922 (N_14922,N_13470,N_13198);
or U14923 (N_14923,N_13768,N_13745);
and U14924 (N_14924,N_13580,N_13062);
and U14925 (N_14925,N_13396,N_13528);
nand U14926 (N_14926,N_13831,N_13472);
nand U14927 (N_14927,N_13464,N_13387);
nor U14928 (N_14928,N_13579,N_13450);
and U14929 (N_14929,N_13715,N_13955);
nand U14930 (N_14930,N_13441,N_13850);
xor U14931 (N_14931,N_13925,N_13802);
xor U14932 (N_14932,N_13364,N_13707);
nand U14933 (N_14933,N_13050,N_13406);
or U14934 (N_14934,N_13576,N_13275);
or U14935 (N_14935,N_13232,N_13662);
nor U14936 (N_14936,N_13098,N_13286);
nand U14937 (N_14937,N_13197,N_13277);
and U14938 (N_14938,N_13178,N_13026);
nand U14939 (N_14939,N_13396,N_13591);
and U14940 (N_14940,N_13079,N_13240);
nand U14941 (N_14941,N_13416,N_13357);
nand U14942 (N_14942,N_13304,N_13650);
nand U14943 (N_14943,N_13553,N_13878);
or U14944 (N_14944,N_13325,N_13874);
nand U14945 (N_14945,N_13839,N_13151);
and U14946 (N_14946,N_13934,N_13775);
and U14947 (N_14947,N_13887,N_13642);
or U14948 (N_14948,N_13534,N_13991);
xor U14949 (N_14949,N_13083,N_13482);
or U14950 (N_14950,N_13676,N_13470);
nor U14951 (N_14951,N_13903,N_13861);
nor U14952 (N_14952,N_13351,N_13694);
nand U14953 (N_14953,N_13697,N_13103);
and U14954 (N_14954,N_13115,N_13214);
or U14955 (N_14955,N_13818,N_13371);
nand U14956 (N_14956,N_13091,N_13554);
and U14957 (N_14957,N_13632,N_13827);
nand U14958 (N_14958,N_13032,N_13232);
nor U14959 (N_14959,N_13663,N_13743);
nand U14960 (N_14960,N_13727,N_13364);
or U14961 (N_14961,N_13960,N_13501);
nor U14962 (N_14962,N_13633,N_13742);
nand U14963 (N_14963,N_13122,N_13133);
nor U14964 (N_14964,N_13894,N_13488);
and U14965 (N_14965,N_13051,N_13843);
nand U14966 (N_14966,N_13013,N_13582);
xnor U14967 (N_14967,N_13162,N_13144);
nand U14968 (N_14968,N_13615,N_13001);
nand U14969 (N_14969,N_13378,N_13512);
nand U14970 (N_14970,N_13848,N_13705);
or U14971 (N_14971,N_13483,N_13717);
and U14972 (N_14972,N_13552,N_13907);
xnor U14973 (N_14973,N_13202,N_13358);
nor U14974 (N_14974,N_13548,N_13241);
nor U14975 (N_14975,N_13166,N_13868);
nor U14976 (N_14976,N_13902,N_13854);
and U14977 (N_14977,N_13329,N_13724);
nand U14978 (N_14978,N_13485,N_13702);
nand U14979 (N_14979,N_13367,N_13139);
and U14980 (N_14980,N_13763,N_13754);
or U14981 (N_14981,N_13452,N_13680);
nor U14982 (N_14982,N_13515,N_13496);
nand U14983 (N_14983,N_13394,N_13940);
or U14984 (N_14984,N_13022,N_13567);
nand U14985 (N_14985,N_13004,N_13018);
or U14986 (N_14986,N_13306,N_13070);
and U14987 (N_14987,N_13171,N_13496);
nand U14988 (N_14988,N_13598,N_13029);
and U14989 (N_14989,N_13485,N_13155);
or U14990 (N_14990,N_13698,N_13721);
nor U14991 (N_14991,N_13522,N_13408);
or U14992 (N_14992,N_13571,N_13438);
or U14993 (N_14993,N_13055,N_13019);
nor U14994 (N_14994,N_13562,N_13130);
nor U14995 (N_14995,N_13020,N_13950);
and U14996 (N_14996,N_13096,N_13781);
nand U14997 (N_14997,N_13699,N_13329);
nor U14998 (N_14998,N_13596,N_13301);
nand U14999 (N_14999,N_13053,N_13890);
nor U15000 (N_15000,N_14360,N_14431);
xor U15001 (N_15001,N_14177,N_14068);
nor U15002 (N_15002,N_14058,N_14624);
nand U15003 (N_15003,N_14162,N_14894);
and U15004 (N_15004,N_14565,N_14548);
nor U15005 (N_15005,N_14997,N_14953);
xor U15006 (N_15006,N_14413,N_14229);
nor U15007 (N_15007,N_14044,N_14804);
or U15008 (N_15008,N_14402,N_14689);
or U15009 (N_15009,N_14064,N_14739);
or U15010 (N_15010,N_14764,N_14805);
nor U15011 (N_15011,N_14003,N_14424);
nor U15012 (N_15012,N_14555,N_14608);
or U15013 (N_15013,N_14279,N_14364);
nand U15014 (N_15014,N_14942,N_14949);
or U15015 (N_15015,N_14505,N_14966);
nor U15016 (N_15016,N_14420,N_14782);
nor U15017 (N_15017,N_14909,N_14952);
or U15018 (N_15018,N_14379,N_14538);
xor U15019 (N_15019,N_14595,N_14500);
nand U15020 (N_15020,N_14391,N_14770);
xor U15021 (N_15021,N_14336,N_14275);
nand U15022 (N_15022,N_14726,N_14877);
or U15023 (N_15023,N_14000,N_14258);
and U15024 (N_15024,N_14857,N_14117);
nor U15025 (N_15025,N_14491,N_14182);
or U15026 (N_15026,N_14612,N_14254);
and U15027 (N_15027,N_14015,N_14786);
nor U15028 (N_15028,N_14771,N_14376);
nor U15029 (N_15029,N_14511,N_14311);
xnor U15030 (N_15030,N_14674,N_14390);
or U15031 (N_15031,N_14193,N_14643);
or U15032 (N_15032,N_14762,N_14869);
or U15033 (N_15033,N_14546,N_14340);
and U15034 (N_15034,N_14658,N_14688);
nor U15035 (N_15035,N_14220,N_14242);
nand U15036 (N_15036,N_14063,N_14960);
or U15037 (N_15037,N_14825,N_14169);
and U15038 (N_15038,N_14774,N_14975);
and U15039 (N_15039,N_14002,N_14860);
xor U15040 (N_15040,N_14165,N_14647);
nand U15041 (N_15041,N_14350,N_14706);
xnor U15042 (N_15042,N_14089,N_14691);
or U15043 (N_15043,N_14284,N_14596);
and U15044 (N_15044,N_14702,N_14852);
xnor U15045 (N_15045,N_14125,N_14210);
and U15046 (N_15046,N_14400,N_14832);
and U15047 (N_15047,N_14056,N_14518);
nand U15048 (N_15048,N_14922,N_14432);
and U15049 (N_15049,N_14768,N_14365);
and U15050 (N_15050,N_14441,N_14497);
nor U15051 (N_15051,N_14031,N_14806);
or U15052 (N_15052,N_14423,N_14847);
nand U15053 (N_15053,N_14398,N_14455);
nand U15054 (N_15054,N_14013,N_14679);
and U15055 (N_15055,N_14054,N_14082);
and U15056 (N_15056,N_14260,N_14251);
and U15057 (N_15057,N_14584,N_14175);
nor U15058 (N_15058,N_14204,N_14628);
xnor U15059 (N_15059,N_14507,N_14591);
and U15060 (N_15060,N_14313,N_14623);
nand U15061 (N_15061,N_14813,N_14539);
nor U15062 (N_15062,N_14870,N_14905);
nand U15063 (N_15063,N_14032,N_14247);
nand U15064 (N_15064,N_14589,N_14038);
nand U15065 (N_15065,N_14467,N_14659);
nand U15066 (N_15066,N_14844,N_14701);
and U15067 (N_15067,N_14327,N_14456);
or U15068 (N_15068,N_14334,N_14202);
nor U15069 (N_15069,N_14508,N_14041);
xor U15070 (N_15070,N_14373,N_14824);
xor U15071 (N_15071,N_14920,N_14235);
and U15072 (N_15072,N_14208,N_14673);
or U15073 (N_15073,N_14009,N_14959);
xor U15074 (N_15074,N_14304,N_14040);
nand U15075 (N_15075,N_14447,N_14100);
or U15076 (N_15076,N_14337,N_14822);
nand U15077 (N_15077,N_14719,N_14819);
xor U15078 (N_15078,N_14614,N_14338);
or U15079 (N_15079,N_14914,N_14910);
nand U15080 (N_15080,N_14600,N_14599);
xor U15081 (N_15081,N_14622,N_14401);
nor U15082 (N_15082,N_14918,N_14085);
nand U15083 (N_15083,N_14541,N_14722);
or U15084 (N_15084,N_14296,N_14199);
or U15085 (N_15085,N_14881,N_14629);
nand U15086 (N_15086,N_14371,N_14069);
and U15087 (N_15087,N_14273,N_14903);
xnor U15088 (N_15088,N_14106,N_14223);
xor U15089 (N_15089,N_14131,N_14936);
and U15090 (N_15090,N_14707,N_14862);
nand U15091 (N_15091,N_14471,N_14249);
or U15092 (N_15092,N_14154,N_14195);
xnor U15093 (N_15093,N_14527,N_14409);
and U15094 (N_15094,N_14494,N_14542);
nand U15095 (N_15095,N_14639,N_14670);
and U15096 (N_15096,N_14246,N_14683);
or U15097 (N_15097,N_14482,N_14529);
or U15098 (N_15098,N_14377,N_14236);
nand U15099 (N_15099,N_14607,N_14644);
nand U15100 (N_15100,N_14641,N_14983);
or U15101 (N_15101,N_14461,N_14797);
or U15102 (N_15102,N_14167,N_14119);
and U15103 (N_15103,N_14536,N_14462);
xnor U15104 (N_15104,N_14744,N_14159);
nand U15105 (N_15105,N_14325,N_14287);
xnor U15106 (N_15106,N_14958,N_14451);
or U15107 (N_15107,N_14776,N_14004);
xnor U15108 (N_15108,N_14562,N_14685);
nand U15109 (N_15109,N_14501,N_14924);
or U15110 (N_15110,N_14238,N_14171);
nand U15111 (N_15111,N_14986,N_14289);
nor U15112 (N_15112,N_14713,N_14662);
or U15113 (N_15113,N_14577,N_14381);
xor U15114 (N_15114,N_14605,N_14809);
nand U15115 (N_15115,N_14502,N_14829);
nand U15116 (N_15116,N_14459,N_14152);
nor U15117 (N_15117,N_14704,N_14256);
nand U15118 (N_15118,N_14074,N_14642);
and U15119 (N_15119,N_14603,N_14457);
and U15120 (N_15120,N_14653,N_14439);
nor U15121 (N_15121,N_14687,N_14887);
nor U15122 (N_15122,N_14493,N_14964);
xnor U15123 (N_15123,N_14445,N_14084);
nand U15124 (N_15124,N_14102,N_14933);
nor U15125 (N_15125,N_14522,N_14323);
nand U15126 (N_15126,N_14593,N_14873);
nor U15127 (N_15127,N_14686,N_14876);
nand U15128 (N_15128,N_14524,N_14579);
or U15129 (N_15129,N_14427,N_14521);
and U15130 (N_15130,N_14245,N_14648);
and U15131 (N_15131,N_14792,N_14477);
xnor U15132 (N_15132,N_14791,N_14950);
nor U15133 (N_15133,N_14135,N_14341);
nand U15134 (N_15134,N_14884,N_14594);
nand U15135 (N_15135,N_14332,N_14855);
and U15136 (N_15136,N_14333,N_14987);
nor U15137 (N_15137,N_14517,N_14556);
nor U15138 (N_15138,N_14422,N_14863);
nor U15139 (N_15139,N_14026,N_14788);
and U15140 (N_15140,N_14209,N_14071);
and U15141 (N_15141,N_14228,N_14990);
and U15142 (N_15142,N_14039,N_14488);
and U15143 (N_15143,N_14853,N_14740);
nor U15144 (N_15144,N_14028,N_14898);
nand U15145 (N_15145,N_14928,N_14230);
or U15146 (N_15146,N_14720,N_14277);
and U15147 (N_15147,N_14576,N_14976);
and U15148 (N_15148,N_14144,N_14292);
and U15149 (N_15149,N_14328,N_14440);
xnor U15150 (N_15150,N_14170,N_14370);
nor U15151 (N_15151,N_14879,N_14295);
xor U15152 (N_15152,N_14145,N_14940);
nor U15153 (N_15153,N_14549,N_14231);
nor U15154 (N_15154,N_14259,N_14951);
nand U15155 (N_15155,N_14601,N_14742);
nand U15156 (N_15156,N_14318,N_14753);
and U15157 (N_15157,N_14465,N_14087);
and U15158 (N_15158,N_14808,N_14161);
nor U15159 (N_15159,N_14225,N_14317);
nor U15160 (N_15160,N_14344,N_14394);
nand U15161 (N_15161,N_14970,N_14160);
or U15162 (N_15162,N_14078,N_14885);
nor U15163 (N_15163,N_14414,N_14769);
nand U15164 (N_15164,N_14925,N_14967);
and U15165 (N_15165,N_14257,N_14785);
or U15166 (N_15166,N_14417,N_14005);
and U15167 (N_15167,N_14592,N_14757);
and U15168 (N_15168,N_14570,N_14790);
or U15169 (N_15169,N_14961,N_14977);
or U15170 (N_15170,N_14814,N_14906);
and U15171 (N_15171,N_14046,N_14429);
or U15172 (N_15172,N_14018,N_14416);
nor U15173 (N_15173,N_14891,N_14203);
and U15174 (N_15174,N_14682,N_14811);
nand U15175 (N_15175,N_14834,N_14554);
and U15176 (N_15176,N_14897,N_14916);
nand U15177 (N_15177,N_14267,N_14405);
or U15178 (N_15178,N_14120,N_14619);
nand U15179 (N_15179,N_14319,N_14205);
and U15180 (N_15180,N_14871,N_14481);
and U15181 (N_15181,N_14047,N_14567);
nand U15182 (N_15182,N_14676,N_14315);
or U15183 (N_15183,N_14303,N_14866);
and U15184 (N_15184,N_14915,N_14627);
or U15185 (N_15185,N_14290,N_14184);
xor U15186 (N_15186,N_14557,N_14362);
nand U15187 (N_15187,N_14859,N_14331);
nand U15188 (N_15188,N_14540,N_14351);
nor U15189 (N_15189,N_14842,N_14307);
or U15190 (N_15190,N_14930,N_14008);
or U15191 (N_15191,N_14566,N_14727);
xor U15192 (N_15192,N_14052,N_14750);
nand U15193 (N_15193,N_14248,N_14343);
xnor U15194 (N_15194,N_14001,N_14393);
nor U15195 (N_15195,N_14291,N_14618);
nand U15196 (N_15196,N_14140,N_14412);
and U15197 (N_15197,N_14178,N_14868);
and U15198 (N_15198,N_14191,N_14712);
nor U15199 (N_15199,N_14219,N_14094);
xor U15200 (N_15200,N_14747,N_14474);
and U15201 (N_15201,N_14748,N_14559);
nor U15202 (N_15202,N_14124,N_14478);
nand U15203 (N_15203,N_14156,N_14901);
nand U15204 (N_15204,N_14252,N_14407);
nand U15205 (N_15205,N_14514,N_14569);
nor U15206 (N_15206,N_14316,N_14011);
or U15207 (N_15207,N_14543,N_14227);
or U15208 (N_15208,N_14921,N_14148);
nand U15209 (N_15209,N_14388,N_14992);
nor U15210 (N_15210,N_14288,N_14198);
nand U15211 (N_15211,N_14941,N_14312);
xnor U15212 (N_15212,N_14787,N_14649);
nand U15213 (N_15213,N_14993,N_14587);
nor U15214 (N_15214,N_14616,N_14356);
nand U15215 (N_15215,N_14820,N_14646);
xnor U15216 (N_15216,N_14262,N_14929);
nor U15217 (N_15217,N_14021,N_14982);
nor U15218 (N_15218,N_14446,N_14515);
nor U15219 (N_15219,N_14904,N_14525);
or U15220 (N_15220,N_14127,N_14783);
and U15221 (N_15221,N_14080,N_14263);
or U15222 (N_15222,N_14359,N_14917);
nand U15223 (N_15223,N_14489,N_14985);
or U15224 (N_15224,N_14544,N_14705);
and U15225 (N_15225,N_14573,N_14907);
nor U15226 (N_15226,N_14947,N_14664);
and U15227 (N_15227,N_14865,N_14133);
or U15228 (N_15228,N_14828,N_14221);
and U15229 (N_15229,N_14116,N_14610);
nor U15230 (N_15230,N_14025,N_14217);
nor U15231 (N_15231,N_14716,N_14758);
or U15232 (N_15232,N_14314,N_14483);
xnor U15233 (N_15233,N_14807,N_14794);
and U15234 (N_15234,N_14123,N_14927);
and U15235 (N_15235,N_14437,N_14850);
xnor U15236 (N_15236,N_14112,N_14751);
and U15237 (N_15237,N_14433,N_14572);
xor U15238 (N_15238,N_14968,N_14956);
nor U15239 (N_15239,N_14625,N_14972);
or U15240 (N_15240,N_14157,N_14717);
and U15241 (N_15241,N_14974,N_14900);
and U15242 (N_15242,N_14597,N_14732);
nor U15243 (N_15243,N_14721,N_14265);
or U15244 (N_15244,N_14841,N_14272);
xor U15245 (N_15245,N_14070,N_14837);
nand U15246 (N_15246,N_14931,N_14519);
nand U15247 (N_15247,N_14324,N_14406);
and U15248 (N_15248,N_14139,N_14954);
nor U15249 (N_15249,N_14656,N_14419);
or U15250 (N_15250,N_14428,N_14241);
nor U15251 (N_15251,N_14746,N_14874);
and U15252 (N_15252,N_14669,N_14697);
nor U15253 (N_15253,N_14151,N_14410);
or U15254 (N_15254,N_14113,N_14654);
nand U15255 (N_15255,N_14613,N_14269);
or U15256 (N_15256,N_14476,N_14346);
nor U15257 (N_15257,N_14633,N_14189);
or U15258 (N_15258,N_14700,N_14609);
nand U15259 (N_15259,N_14763,N_14411);
and U15260 (N_15260,N_14963,N_14239);
or U15261 (N_15261,N_14066,N_14839);
and U15262 (N_15262,N_14743,N_14073);
nor U15263 (N_15263,N_14014,N_14196);
nand U15264 (N_15264,N_14023,N_14183);
or U15265 (N_15265,N_14201,N_14128);
nand U15266 (N_15266,N_14109,N_14270);
and U15267 (N_15267,N_14766,N_14564);
nand U15268 (N_15268,N_14108,N_14784);
nand U15269 (N_15269,N_14382,N_14163);
nor U15270 (N_15270,N_14075,N_14092);
nand U15271 (N_15271,N_14838,N_14551);
nor U15272 (N_15272,N_14492,N_14077);
or U15273 (N_15273,N_14661,N_14297);
and U15274 (N_15274,N_14999,N_14043);
nand U15275 (N_15275,N_14093,N_14735);
or U15276 (N_15276,N_14458,N_14244);
and U15277 (N_15277,N_14660,N_14798);
and U15278 (N_15278,N_14114,N_14053);
nor U15279 (N_15279,N_14442,N_14450);
nor U15280 (N_15280,N_14728,N_14192);
nand U15281 (N_15281,N_14215,N_14520);
and U15282 (N_15282,N_14197,N_14979);
xor U15283 (N_15283,N_14283,N_14761);
or U15284 (N_15284,N_14655,N_14115);
and U15285 (N_15285,N_14060,N_14715);
xnor U15286 (N_15286,N_14583,N_14438);
xor U15287 (N_15287,N_14725,N_14155);
nand U15288 (N_15288,N_14981,N_14752);
nand U15289 (N_15289,N_14734,N_14578);
or U15290 (N_15290,N_14965,N_14306);
nor U15291 (N_15291,N_14590,N_14361);
nor U15292 (N_15292,N_14472,N_14878);
and U15293 (N_15293,N_14250,N_14435);
or U15294 (N_15294,N_14090,N_14872);
nand U15295 (N_15295,N_14888,N_14765);
nand U15296 (N_15296,N_14848,N_14464);
nand U15297 (N_15297,N_14380,N_14321);
nor U15298 (N_15298,N_14368,N_14532);
and U15299 (N_15299,N_14640,N_14358);
nor U15300 (N_15300,N_14062,N_14935);
or U15301 (N_15301,N_14759,N_14799);
nor U15302 (N_15302,N_14158,N_14330);
and U15303 (N_15303,N_14946,N_14449);
or U15304 (N_15304,N_14430,N_14998);
xnor U15305 (N_15305,N_14523,N_14657);
nor U15306 (N_15306,N_14582,N_14234);
nand U15307 (N_15307,N_14988,N_14767);
or U15308 (N_15308,N_14126,N_14281);
nor U15309 (N_15309,N_14187,N_14487);
nor U15310 (N_15310,N_14190,N_14937);
and U15311 (N_15311,N_14086,N_14301);
and U15312 (N_15312,N_14280,N_14996);
xor U15313 (N_15313,N_14867,N_14448);
nand U15314 (N_15314,N_14232,N_14694);
nor U15315 (N_15315,N_14233,N_14035);
nor U15316 (N_15316,N_14835,N_14995);
or U15317 (N_15317,N_14347,N_14237);
and U15318 (N_15318,N_14718,N_14635);
nor U15319 (N_15319,N_14348,N_14059);
and U15320 (N_15320,N_14699,N_14800);
and U15321 (N_15321,N_14504,N_14938);
nand U15322 (N_15322,N_14285,N_14030);
or U15323 (N_15323,N_14650,N_14096);
and U15324 (N_15324,N_14027,N_14989);
nand U15325 (N_15325,N_14072,N_14469);
or U15326 (N_15326,N_14695,N_14580);
or U15327 (N_15327,N_14206,N_14810);
and U15328 (N_15328,N_14268,N_14733);
nand U15329 (N_15329,N_14374,N_14530);
xnor U15330 (N_15330,N_14948,N_14710);
or U15331 (N_15331,N_14385,N_14255);
nor U15332 (N_15332,N_14286,N_14369);
xnor U15333 (N_15333,N_14463,N_14741);
nor U15334 (N_15334,N_14378,N_14499);
nor U15335 (N_15335,N_14355,N_14353);
nand U15336 (N_15336,N_14994,N_14802);
nand U15337 (N_15337,N_14711,N_14496);
or U15338 (N_15338,N_14668,N_14226);
xor U15339 (N_15339,N_14083,N_14545);
nor U15340 (N_15340,N_14147,N_14984);
and U15341 (N_15341,N_14651,N_14991);
nor U15342 (N_15342,N_14218,N_14065);
nor U15343 (N_15343,N_14632,N_14150);
nor U15344 (N_15344,N_14383,N_14864);
nor U15345 (N_15345,N_14444,N_14480);
and U15346 (N_15346,N_14626,N_14007);
and U15347 (N_15347,N_14773,N_14425);
nor U15348 (N_15348,N_14051,N_14121);
nand U15349 (N_15349,N_14076,N_14194);
nor U15350 (N_15350,N_14923,N_14172);
nand U15351 (N_15351,N_14851,N_14266);
or U15352 (N_15352,N_14558,N_14146);
and U15353 (N_15353,N_14561,N_14781);
xnor U15354 (N_15354,N_14261,N_14278);
and U15355 (N_15355,N_14528,N_14585);
and U15356 (N_15356,N_14602,N_14470);
or U15357 (N_15357,N_14436,N_14403);
nand U15358 (N_15358,N_14029,N_14200);
nor U15359 (N_15359,N_14854,N_14510);
nand U15360 (N_15360,N_14034,N_14738);
and U15361 (N_15361,N_14902,N_14132);
and U15362 (N_15362,N_14858,N_14138);
and U15363 (N_15363,N_14253,N_14443);
nor U15364 (N_15364,N_14421,N_14957);
and U15365 (N_15365,N_14775,N_14375);
xor U15366 (N_15366,N_14693,N_14274);
or U15367 (N_15367,N_14534,N_14944);
nand U15368 (N_15368,N_14088,N_14971);
and U15369 (N_15369,N_14479,N_14067);
nand U15370 (N_15370,N_14908,N_14620);
nor U15371 (N_15371,N_14690,N_14598);
nand U15372 (N_15372,N_14216,N_14310);
nand U15373 (N_15373,N_14883,N_14207);
xor U15374 (N_15374,N_14962,N_14755);
and U15375 (N_15375,N_14550,N_14498);
or U15376 (N_15376,N_14892,N_14271);
or U15377 (N_15377,N_14815,N_14042);
nand U15378 (N_15378,N_14434,N_14387);
nor U15379 (N_15379,N_14495,N_14553);
nand U15380 (N_15380,N_14037,N_14389);
and U15381 (N_15381,N_14017,N_14777);
nand U15382 (N_15382,N_14033,N_14836);
or U15383 (N_15383,N_14454,N_14631);
and U15384 (N_15384,N_14022,N_14484);
or U15385 (N_15385,N_14045,N_14506);
xor U15386 (N_15386,N_14696,N_14778);
nand U15387 (N_15387,N_14714,N_14095);
nor U15388 (N_15388,N_14490,N_14919);
nor U15389 (N_15389,N_14104,N_14130);
xor U15390 (N_15390,N_14723,N_14934);
nand U15391 (N_15391,N_14049,N_14667);
nor U15392 (N_15392,N_14845,N_14675);
and U15393 (N_15393,N_14560,N_14932);
nand U15394 (N_15394,N_14335,N_14418);
xor U15395 (N_15395,N_14955,N_14637);
and U15396 (N_15396,N_14212,N_14166);
and U15397 (N_15397,N_14342,N_14680);
nor U15398 (N_15398,N_14760,N_14415);
and U15399 (N_15399,N_14136,N_14081);
and U15400 (N_15400,N_14293,N_14574);
nand U15401 (N_15401,N_14575,N_14945);
nand U15402 (N_15402,N_14475,N_14912);
nand U15403 (N_15403,N_14509,N_14621);
and U15404 (N_15404,N_14731,N_14173);
or U15405 (N_15405,N_14737,N_14552);
nand U15406 (N_15406,N_14322,N_14816);
or U15407 (N_15407,N_14010,N_14392);
nor U15408 (N_15408,N_14408,N_14535);
and U15409 (N_15409,N_14630,N_14396);
or U15410 (N_15410,N_14168,N_14666);
or U15411 (N_15411,N_14973,N_14186);
nor U15412 (N_15412,N_14404,N_14181);
and U15413 (N_15413,N_14856,N_14386);
xnor U15414 (N_15414,N_14357,N_14305);
nor U15415 (N_15415,N_14754,N_14188);
nor U15416 (N_15416,N_14512,N_14213);
xnor U15417 (N_15417,N_14048,N_14818);
nor U15418 (N_15418,N_14745,N_14730);
nor U15419 (N_15419,N_14243,N_14533);
xnor U15420 (N_15420,N_14830,N_14547);
nand U15421 (N_15421,N_14638,N_14012);
nor U15422 (N_15422,N_14309,N_14671);
nand U15423 (N_15423,N_14122,N_14796);
nand U15424 (N_15424,N_14672,N_14354);
or U15425 (N_15425,N_14320,N_14882);
nor U15426 (N_15426,N_14397,N_14276);
and U15427 (N_15427,N_14895,N_14185);
or U15428 (N_15428,N_14061,N_14019);
and U15429 (N_15429,N_14645,N_14568);
and U15430 (N_15430,N_14843,N_14665);
or U15431 (N_15431,N_14789,N_14692);
and U15432 (N_15432,N_14604,N_14681);
nand U15433 (N_15433,N_14345,N_14055);
or U15434 (N_15434,N_14893,N_14849);
or U15435 (N_15435,N_14174,N_14801);
nor U15436 (N_15436,N_14142,N_14372);
xor U15437 (N_15437,N_14890,N_14298);
xnor U15438 (N_15438,N_14329,N_14101);
or U15439 (N_15439,N_14780,N_14817);
xnor U15440 (N_15440,N_14240,N_14282);
or U15441 (N_15441,N_14363,N_14833);
or U15442 (N_15442,N_14006,N_14164);
or U15443 (N_15443,N_14098,N_14978);
nor U15444 (N_15444,N_14826,N_14980);
and U15445 (N_15445,N_14485,N_14803);
nand U15446 (N_15446,N_14516,N_14581);
nor U15447 (N_15447,N_14107,N_14308);
or U15448 (N_15448,N_14452,N_14137);
or U15449 (N_15449,N_14020,N_14339);
xnor U15450 (N_15450,N_14468,N_14176);
and U15451 (N_15451,N_14831,N_14846);
nor U15452 (N_15452,N_14036,N_14326);
nand U15453 (N_15453,N_14821,N_14677);
or U15454 (N_15454,N_14460,N_14143);
xnor U15455 (N_15455,N_14611,N_14103);
nor U15456 (N_15456,N_14615,N_14703);
and U15457 (N_15457,N_14636,N_14503);
and U15458 (N_15458,N_14724,N_14652);
and U15459 (N_15459,N_14264,N_14097);
nor U15460 (N_15460,N_14708,N_14110);
and U15461 (N_15461,N_14526,N_14889);
nor U15462 (N_15462,N_14211,N_14663);
nor U15463 (N_15463,N_14861,N_14367);
or U15464 (N_15464,N_14793,N_14466);
nor U15465 (N_15465,N_14840,N_14453);
or U15466 (N_15466,N_14099,N_14299);
and U15467 (N_15467,N_14823,N_14016);
and U15468 (N_15468,N_14426,N_14756);
or U15469 (N_15469,N_14926,N_14024);
nor U15470 (N_15470,N_14827,N_14729);
or U15471 (N_15471,N_14079,N_14179);
or U15472 (N_15472,N_14886,N_14709);
nand U15473 (N_15473,N_14913,N_14606);
xnor U15474 (N_15474,N_14779,N_14294);
or U15475 (N_15475,N_14875,N_14105);
and U15476 (N_15476,N_14588,N_14634);
and U15477 (N_15477,N_14129,N_14224);
nor U15478 (N_15478,N_14513,N_14911);
nand U15479 (N_15479,N_14772,N_14698);
nand U15480 (N_15480,N_14486,N_14684);
xnor U15481 (N_15481,N_14091,N_14352);
nor U15482 (N_15482,N_14395,N_14749);
nand U15483 (N_15483,N_14399,N_14563);
nor U15484 (N_15484,N_14222,N_14214);
nand U15485 (N_15485,N_14943,N_14180);
and U15486 (N_15486,N_14678,N_14969);
nand U15487 (N_15487,N_14111,N_14473);
or U15488 (N_15488,N_14302,N_14349);
nor U15489 (N_15489,N_14896,N_14300);
or U15490 (N_15490,N_14057,N_14617);
nand U15491 (N_15491,N_14899,N_14134);
or U15492 (N_15492,N_14050,N_14118);
or U15493 (N_15493,N_14795,N_14366);
nor U15494 (N_15494,N_14537,N_14149);
or U15495 (N_15495,N_14586,N_14736);
and U15496 (N_15496,N_14880,N_14571);
or U15497 (N_15497,N_14939,N_14153);
nor U15498 (N_15498,N_14141,N_14531);
or U15499 (N_15499,N_14812,N_14384);
xnor U15500 (N_15500,N_14723,N_14136);
nand U15501 (N_15501,N_14705,N_14158);
or U15502 (N_15502,N_14641,N_14120);
or U15503 (N_15503,N_14397,N_14789);
and U15504 (N_15504,N_14837,N_14169);
and U15505 (N_15505,N_14425,N_14358);
or U15506 (N_15506,N_14842,N_14577);
xnor U15507 (N_15507,N_14949,N_14088);
nand U15508 (N_15508,N_14345,N_14551);
or U15509 (N_15509,N_14243,N_14364);
nor U15510 (N_15510,N_14002,N_14438);
nand U15511 (N_15511,N_14253,N_14577);
nor U15512 (N_15512,N_14333,N_14168);
nor U15513 (N_15513,N_14893,N_14892);
nand U15514 (N_15514,N_14978,N_14162);
nand U15515 (N_15515,N_14943,N_14840);
nand U15516 (N_15516,N_14767,N_14713);
or U15517 (N_15517,N_14183,N_14464);
nor U15518 (N_15518,N_14807,N_14932);
or U15519 (N_15519,N_14031,N_14346);
or U15520 (N_15520,N_14020,N_14296);
nand U15521 (N_15521,N_14273,N_14742);
or U15522 (N_15522,N_14969,N_14282);
or U15523 (N_15523,N_14311,N_14961);
nand U15524 (N_15524,N_14411,N_14111);
nand U15525 (N_15525,N_14088,N_14460);
or U15526 (N_15526,N_14876,N_14027);
and U15527 (N_15527,N_14960,N_14784);
nor U15528 (N_15528,N_14537,N_14994);
and U15529 (N_15529,N_14859,N_14588);
or U15530 (N_15530,N_14316,N_14504);
or U15531 (N_15531,N_14786,N_14100);
nand U15532 (N_15532,N_14261,N_14156);
nand U15533 (N_15533,N_14336,N_14092);
or U15534 (N_15534,N_14185,N_14923);
xnor U15535 (N_15535,N_14553,N_14231);
and U15536 (N_15536,N_14638,N_14090);
or U15537 (N_15537,N_14891,N_14283);
nor U15538 (N_15538,N_14147,N_14909);
nand U15539 (N_15539,N_14130,N_14353);
or U15540 (N_15540,N_14782,N_14802);
or U15541 (N_15541,N_14910,N_14662);
xnor U15542 (N_15542,N_14098,N_14950);
or U15543 (N_15543,N_14917,N_14532);
xnor U15544 (N_15544,N_14727,N_14678);
nand U15545 (N_15545,N_14627,N_14894);
nor U15546 (N_15546,N_14391,N_14997);
and U15547 (N_15547,N_14383,N_14741);
nand U15548 (N_15548,N_14046,N_14819);
or U15549 (N_15549,N_14498,N_14353);
nand U15550 (N_15550,N_14386,N_14288);
or U15551 (N_15551,N_14682,N_14869);
nor U15552 (N_15552,N_14173,N_14945);
nand U15553 (N_15553,N_14910,N_14343);
or U15554 (N_15554,N_14368,N_14462);
nand U15555 (N_15555,N_14039,N_14254);
xnor U15556 (N_15556,N_14155,N_14800);
nor U15557 (N_15557,N_14475,N_14579);
or U15558 (N_15558,N_14234,N_14777);
nand U15559 (N_15559,N_14122,N_14988);
or U15560 (N_15560,N_14715,N_14730);
and U15561 (N_15561,N_14051,N_14604);
nor U15562 (N_15562,N_14132,N_14107);
and U15563 (N_15563,N_14348,N_14990);
or U15564 (N_15564,N_14145,N_14921);
or U15565 (N_15565,N_14239,N_14679);
nor U15566 (N_15566,N_14949,N_14516);
nand U15567 (N_15567,N_14116,N_14424);
nand U15568 (N_15568,N_14320,N_14590);
and U15569 (N_15569,N_14223,N_14924);
or U15570 (N_15570,N_14030,N_14953);
or U15571 (N_15571,N_14444,N_14528);
and U15572 (N_15572,N_14264,N_14208);
and U15573 (N_15573,N_14669,N_14059);
or U15574 (N_15574,N_14640,N_14905);
and U15575 (N_15575,N_14248,N_14296);
xnor U15576 (N_15576,N_14091,N_14143);
nor U15577 (N_15577,N_14722,N_14922);
nand U15578 (N_15578,N_14968,N_14484);
nor U15579 (N_15579,N_14567,N_14421);
nor U15580 (N_15580,N_14003,N_14774);
or U15581 (N_15581,N_14183,N_14393);
nor U15582 (N_15582,N_14363,N_14463);
nor U15583 (N_15583,N_14549,N_14425);
and U15584 (N_15584,N_14277,N_14066);
and U15585 (N_15585,N_14944,N_14974);
or U15586 (N_15586,N_14552,N_14042);
nor U15587 (N_15587,N_14576,N_14375);
nand U15588 (N_15588,N_14853,N_14348);
nor U15589 (N_15589,N_14262,N_14324);
or U15590 (N_15590,N_14766,N_14568);
nand U15591 (N_15591,N_14518,N_14849);
or U15592 (N_15592,N_14584,N_14088);
and U15593 (N_15593,N_14286,N_14005);
nor U15594 (N_15594,N_14436,N_14311);
xnor U15595 (N_15595,N_14496,N_14105);
or U15596 (N_15596,N_14083,N_14770);
or U15597 (N_15597,N_14327,N_14013);
and U15598 (N_15598,N_14514,N_14978);
and U15599 (N_15599,N_14535,N_14933);
or U15600 (N_15600,N_14698,N_14911);
and U15601 (N_15601,N_14233,N_14200);
nand U15602 (N_15602,N_14872,N_14340);
nand U15603 (N_15603,N_14600,N_14763);
or U15604 (N_15604,N_14153,N_14735);
nand U15605 (N_15605,N_14919,N_14757);
xor U15606 (N_15606,N_14788,N_14525);
or U15607 (N_15607,N_14869,N_14142);
nand U15608 (N_15608,N_14439,N_14445);
or U15609 (N_15609,N_14634,N_14815);
and U15610 (N_15610,N_14799,N_14974);
nor U15611 (N_15611,N_14050,N_14892);
nor U15612 (N_15612,N_14785,N_14673);
nand U15613 (N_15613,N_14498,N_14715);
or U15614 (N_15614,N_14155,N_14440);
and U15615 (N_15615,N_14658,N_14220);
or U15616 (N_15616,N_14213,N_14393);
and U15617 (N_15617,N_14625,N_14927);
or U15618 (N_15618,N_14717,N_14804);
nor U15619 (N_15619,N_14870,N_14927);
or U15620 (N_15620,N_14628,N_14920);
and U15621 (N_15621,N_14206,N_14883);
xnor U15622 (N_15622,N_14127,N_14545);
or U15623 (N_15623,N_14355,N_14104);
or U15624 (N_15624,N_14751,N_14035);
nor U15625 (N_15625,N_14246,N_14476);
nand U15626 (N_15626,N_14947,N_14358);
or U15627 (N_15627,N_14692,N_14660);
nor U15628 (N_15628,N_14958,N_14788);
and U15629 (N_15629,N_14373,N_14104);
or U15630 (N_15630,N_14869,N_14848);
nand U15631 (N_15631,N_14988,N_14873);
and U15632 (N_15632,N_14247,N_14895);
and U15633 (N_15633,N_14187,N_14091);
or U15634 (N_15634,N_14856,N_14770);
xor U15635 (N_15635,N_14230,N_14057);
or U15636 (N_15636,N_14539,N_14802);
or U15637 (N_15637,N_14290,N_14051);
or U15638 (N_15638,N_14327,N_14299);
or U15639 (N_15639,N_14931,N_14452);
nand U15640 (N_15640,N_14210,N_14769);
xnor U15641 (N_15641,N_14148,N_14541);
nand U15642 (N_15642,N_14082,N_14621);
or U15643 (N_15643,N_14599,N_14239);
and U15644 (N_15644,N_14366,N_14840);
or U15645 (N_15645,N_14279,N_14935);
xnor U15646 (N_15646,N_14508,N_14339);
nor U15647 (N_15647,N_14178,N_14273);
or U15648 (N_15648,N_14523,N_14194);
or U15649 (N_15649,N_14950,N_14803);
and U15650 (N_15650,N_14059,N_14407);
and U15651 (N_15651,N_14514,N_14428);
xnor U15652 (N_15652,N_14969,N_14816);
nand U15653 (N_15653,N_14973,N_14615);
nor U15654 (N_15654,N_14021,N_14427);
nor U15655 (N_15655,N_14090,N_14216);
nor U15656 (N_15656,N_14428,N_14711);
or U15657 (N_15657,N_14622,N_14020);
and U15658 (N_15658,N_14729,N_14942);
and U15659 (N_15659,N_14098,N_14130);
xnor U15660 (N_15660,N_14716,N_14929);
and U15661 (N_15661,N_14224,N_14849);
nor U15662 (N_15662,N_14992,N_14782);
nand U15663 (N_15663,N_14524,N_14775);
and U15664 (N_15664,N_14939,N_14820);
nand U15665 (N_15665,N_14888,N_14462);
or U15666 (N_15666,N_14402,N_14460);
nand U15667 (N_15667,N_14559,N_14442);
and U15668 (N_15668,N_14092,N_14870);
xor U15669 (N_15669,N_14619,N_14528);
xnor U15670 (N_15670,N_14073,N_14146);
nor U15671 (N_15671,N_14259,N_14343);
nand U15672 (N_15672,N_14984,N_14530);
nand U15673 (N_15673,N_14951,N_14772);
xnor U15674 (N_15674,N_14667,N_14887);
nor U15675 (N_15675,N_14715,N_14913);
and U15676 (N_15676,N_14930,N_14655);
or U15677 (N_15677,N_14893,N_14261);
or U15678 (N_15678,N_14041,N_14415);
or U15679 (N_15679,N_14590,N_14083);
and U15680 (N_15680,N_14205,N_14076);
nand U15681 (N_15681,N_14488,N_14600);
and U15682 (N_15682,N_14536,N_14157);
or U15683 (N_15683,N_14829,N_14247);
or U15684 (N_15684,N_14486,N_14265);
and U15685 (N_15685,N_14307,N_14974);
nand U15686 (N_15686,N_14152,N_14402);
nor U15687 (N_15687,N_14373,N_14712);
xnor U15688 (N_15688,N_14704,N_14828);
or U15689 (N_15689,N_14492,N_14004);
nor U15690 (N_15690,N_14477,N_14239);
nand U15691 (N_15691,N_14443,N_14467);
nor U15692 (N_15692,N_14355,N_14370);
or U15693 (N_15693,N_14165,N_14814);
and U15694 (N_15694,N_14623,N_14962);
nor U15695 (N_15695,N_14973,N_14422);
xnor U15696 (N_15696,N_14915,N_14474);
xor U15697 (N_15697,N_14611,N_14567);
nand U15698 (N_15698,N_14965,N_14270);
nand U15699 (N_15699,N_14996,N_14639);
and U15700 (N_15700,N_14656,N_14585);
or U15701 (N_15701,N_14243,N_14749);
and U15702 (N_15702,N_14440,N_14579);
nand U15703 (N_15703,N_14107,N_14936);
or U15704 (N_15704,N_14842,N_14385);
or U15705 (N_15705,N_14025,N_14775);
or U15706 (N_15706,N_14263,N_14230);
and U15707 (N_15707,N_14672,N_14407);
or U15708 (N_15708,N_14146,N_14851);
nand U15709 (N_15709,N_14274,N_14154);
or U15710 (N_15710,N_14099,N_14418);
nor U15711 (N_15711,N_14688,N_14470);
or U15712 (N_15712,N_14783,N_14576);
nand U15713 (N_15713,N_14822,N_14364);
and U15714 (N_15714,N_14877,N_14984);
and U15715 (N_15715,N_14713,N_14240);
and U15716 (N_15716,N_14658,N_14093);
and U15717 (N_15717,N_14806,N_14477);
or U15718 (N_15718,N_14771,N_14845);
and U15719 (N_15719,N_14688,N_14281);
or U15720 (N_15720,N_14131,N_14817);
or U15721 (N_15721,N_14814,N_14690);
nand U15722 (N_15722,N_14883,N_14062);
nand U15723 (N_15723,N_14422,N_14833);
and U15724 (N_15724,N_14596,N_14784);
nor U15725 (N_15725,N_14505,N_14140);
nor U15726 (N_15726,N_14291,N_14995);
and U15727 (N_15727,N_14894,N_14595);
xnor U15728 (N_15728,N_14562,N_14438);
nand U15729 (N_15729,N_14214,N_14838);
nand U15730 (N_15730,N_14422,N_14403);
nand U15731 (N_15731,N_14422,N_14955);
nand U15732 (N_15732,N_14568,N_14849);
nand U15733 (N_15733,N_14185,N_14943);
nand U15734 (N_15734,N_14086,N_14106);
xor U15735 (N_15735,N_14543,N_14980);
nor U15736 (N_15736,N_14778,N_14577);
nor U15737 (N_15737,N_14961,N_14330);
nand U15738 (N_15738,N_14434,N_14749);
nor U15739 (N_15739,N_14667,N_14061);
nand U15740 (N_15740,N_14932,N_14586);
or U15741 (N_15741,N_14842,N_14250);
and U15742 (N_15742,N_14791,N_14273);
and U15743 (N_15743,N_14343,N_14449);
nand U15744 (N_15744,N_14812,N_14605);
nand U15745 (N_15745,N_14592,N_14734);
and U15746 (N_15746,N_14464,N_14945);
and U15747 (N_15747,N_14420,N_14914);
and U15748 (N_15748,N_14770,N_14218);
nor U15749 (N_15749,N_14414,N_14346);
nand U15750 (N_15750,N_14924,N_14960);
and U15751 (N_15751,N_14227,N_14681);
nand U15752 (N_15752,N_14828,N_14244);
nor U15753 (N_15753,N_14861,N_14947);
and U15754 (N_15754,N_14593,N_14506);
nor U15755 (N_15755,N_14312,N_14153);
and U15756 (N_15756,N_14308,N_14813);
nor U15757 (N_15757,N_14178,N_14478);
and U15758 (N_15758,N_14522,N_14217);
nand U15759 (N_15759,N_14624,N_14449);
and U15760 (N_15760,N_14957,N_14920);
nor U15761 (N_15761,N_14671,N_14396);
nand U15762 (N_15762,N_14811,N_14403);
nor U15763 (N_15763,N_14321,N_14991);
nand U15764 (N_15764,N_14825,N_14164);
nor U15765 (N_15765,N_14963,N_14123);
nor U15766 (N_15766,N_14366,N_14550);
nand U15767 (N_15767,N_14376,N_14272);
nor U15768 (N_15768,N_14532,N_14690);
nand U15769 (N_15769,N_14783,N_14978);
nor U15770 (N_15770,N_14559,N_14736);
nor U15771 (N_15771,N_14424,N_14914);
nor U15772 (N_15772,N_14133,N_14351);
and U15773 (N_15773,N_14347,N_14387);
and U15774 (N_15774,N_14248,N_14466);
nand U15775 (N_15775,N_14785,N_14316);
or U15776 (N_15776,N_14353,N_14945);
nor U15777 (N_15777,N_14105,N_14797);
and U15778 (N_15778,N_14463,N_14444);
or U15779 (N_15779,N_14277,N_14663);
xor U15780 (N_15780,N_14074,N_14944);
nand U15781 (N_15781,N_14548,N_14036);
nor U15782 (N_15782,N_14194,N_14487);
xnor U15783 (N_15783,N_14940,N_14262);
nor U15784 (N_15784,N_14433,N_14689);
xnor U15785 (N_15785,N_14544,N_14832);
and U15786 (N_15786,N_14889,N_14736);
or U15787 (N_15787,N_14846,N_14532);
or U15788 (N_15788,N_14895,N_14658);
nor U15789 (N_15789,N_14323,N_14788);
and U15790 (N_15790,N_14691,N_14416);
or U15791 (N_15791,N_14010,N_14623);
and U15792 (N_15792,N_14264,N_14592);
xnor U15793 (N_15793,N_14724,N_14655);
nor U15794 (N_15794,N_14349,N_14672);
nor U15795 (N_15795,N_14472,N_14350);
nand U15796 (N_15796,N_14187,N_14929);
nor U15797 (N_15797,N_14241,N_14989);
xnor U15798 (N_15798,N_14116,N_14089);
or U15799 (N_15799,N_14546,N_14552);
or U15800 (N_15800,N_14439,N_14981);
nor U15801 (N_15801,N_14301,N_14839);
or U15802 (N_15802,N_14465,N_14622);
or U15803 (N_15803,N_14730,N_14993);
xor U15804 (N_15804,N_14810,N_14084);
or U15805 (N_15805,N_14775,N_14099);
and U15806 (N_15806,N_14703,N_14810);
or U15807 (N_15807,N_14641,N_14606);
and U15808 (N_15808,N_14172,N_14594);
and U15809 (N_15809,N_14281,N_14080);
xor U15810 (N_15810,N_14741,N_14700);
nor U15811 (N_15811,N_14765,N_14017);
and U15812 (N_15812,N_14045,N_14232);
or U15813 (N_15813,N_14659,N_14979);
xor U15814 (N_15814,N_14884,N_14438);
and U15815 (N_15815,N_14493,N_14615);
or U15816 (N_15816,N_14990,N_14820);
nor U15817 (N_15817,N_14207,N_14390);
nor U15818 (N_15818,N_14933,N_14001);
nor U15819 (N_15819,N_14600,N_14151);
nand U15820 (N_15820,N_14150,N_14619);
or U15821 (N_15821,N_14882,N_14819);
nor U15822 (N_15822,N_14090,N_14882);
or U15823 (N_15823,N_14569,N_14715);
or U15824 (N_15824,N_14960,N_14524);
nor U15825 (N_15825,N_14865,N_14010);
or U15826 (N_15826,N_14189,N_14617);
nor U15827 (N_15827,N_14821,N_14313);
and U15828 (N_15828,N_14215,N_14906);
nor U15829 (N_15829,N_14046,N_14085);
nand U15830 (N_15830,N_14469,N_14549);
and U15831 (N_15831,N_14813,N_14270);
and U15832 (N_15832,N_14352,N_14514);
or U15833 (N_15833,N_14290,N_14816);
xnor U15834 (N_15834,N_14807,N_14194);
and U15835 (N_15835,N_14343,N_14086);
or U15836 (N_15836,N_14211,N_14589);
and U15837 (N_15837,N_14406,N_14967);
nor U15838 (N_15838,N_14333,N_14732);
nor U15839 (N_15839,N_14492,N_14421);
xor U15840 (N_15840,N_14875,N_14814);
and U15841 (N_15841,N_14876,N_14503);
nand U15842 (N_15842,N_14463,N_14181);
nor U15843 (N_15843,N_14911,N_14259);
nand U15844 (N_15844,N_14872,N_14104);
nor U15845 (N_15845,N_14694,N_14644);
nand U15846 (N_15846,N_14126,N_14571);
and U15847 (N_15847,N_14172,N_14340);
nand U15848 (N_15848,N_14327,N_14497);
and U15849 (N_15849,N_14570,N_14093);
nand U15850 (N_15850,N_14621,N_14083);
nand U15851 (N_15851,N_14381,N_14288);
nand U15852 (N_15852,N_14810,N_14316);
and U15853 (N_15853,N_14896,N_14867);
nand U15854 (N_15854,N_14397,N_14889);
nand U15855 (N_15855,N_14021,N_14985);
nand U15856 (N_15856,N_14811,N_14417);
and U15857 (N_15857,N_14612,N_14537);
nand U15858 (N_15858,N_14796,N_14741);
or U15859 (N_15859,N_14432,N_14056);
and U15860 (N_15860,N_14025,N_14893);
or U15861 (N_15861,N_14128,N_14066);
nand U15862 (N_15862,N_14427,N_14456);
or U15863 (N_15863,N_14476,N_14073);
or U15864 (N_15864,N_14556,N_14932);
and U15865 (N_15865,N_14557,N_14180);
or U15866 (N_15866,N_14483,N_14219);
nand U15867 (N_15867,N_14140,N_14036);
nor U15868 (N_15868,N_14537,N_14695);
nand U15869 (N_15869,N_14830,N_14738);
nor U15870 (N_15870,N_14436,N_14884);
nand U15871 (N_15871,N_14731,N_14863);
nor U15872 (N_15872,N_14891,N_14197);
nand U15873 (N_15873,N_14909,N_14936);
nand U15874 (N_15874,N_14024,N_14662);
and U15875 (N_15875,N_14648,N_14246);
and U15876 (N_15876,N_14841,N_14160);
and U15877 (N_15877,N_14364,N_14278);
or U15878 (N_15878,N_14954,N_14687);
nor U15879 (N_15879,N_14440,N_14006);
and U15880 (N_15880,N_14987,N_14162);
or U15881 (N_15881,N_14576,N_14463);
and U15882 (N_15882,N_14709,N_14050);
and U15883 (N_15883,N_14041,N_14279);
and U15884 (N_15884,N_14353,N_14653);
nand U15885 (N_15885,N_14468,N_14593);
or U15886 (N_15886,N_14158,N_14570);
or U15887 (N_15887,N_14130,N_14122);
and U15888 (N_15888,N_14554,N_14885);
and U15889 (N_15889,N_14320,N_14504);
nor U15890 (N_15890,N_14226,N_14403);
nand U15891 (N_15891,N_14480,N_14384);
nand U15892 (N_15892,N_14021,N_14069);
and U15893 (N_15893,N_14125,N_14934);
xnor U15894 (N_15894,N_14846,N_14379);
xor U15895 (N_15895,N_14026,N_14475);
nor U15896 (N_15896,N_14554,N_14254);
and U15897 (N_15897,N_14248,N_14968);
and U15898 (N_15898,N_14114,N_14560);
or U15899 (N_15899,N_14034,N_14953);
or U15900 (N_15900,N_14469,N_14597);
or U15901 (N_15901,N_14832,N_14316);
nand U15902 (N_15902,N_14857,N_14758);
and U15903 (N_15903,N_14202,N_14922);
and U15904 (N_15904,N_14577,N_14746);
xor U15905 (N_15905,N_14816,N_14017);
and U15906 (N_15906,N_14977,N_14027);
nor U15907 (N_15907,N_14009,N_14136);
nor U15908 (N_15908,N_14191,N_14467);
nor U15909 (N_15909,N_14706,N_14800);
nor U15910 (N_15910,N_14838,N_14076);
and U15911 (N_15911,N_14431,N_14302);
and U15912 (N_15912,N_14308,N_14069);
or U15913 (N_15913,N_14725,N_14732);
or U15914 (N_15914,N_14791,N_14010);
or U15915 (N_15915,N_14920,N_14052);
and U15916 (N_15916,N_14494,N_14989);
nor U15917 (N_15917,N_14138,N_14332);
nand U15918 (N_15918,N_14200,N_14306);
nor U15919 (N_15919,N_14063,N_14805);
nand U15920 (N_15920,N_14982,N_14520);
and U15921 (N_15921,N_14925,N_14143);
nor U15922 (N_15922,N_14860,N_14334);
or U15923 (N_15923,N_14691,N_14321);
or U15924 (N_15924,N_14506,N_14794);
or U15925 (N_15925,N_14590,N_14867);
nor U15926 (N_15926,N_14132,N_14457);
xnor U15927 (N_15927,N_14555,N_14167);
nand U15928 (N_15928,N_14969,N_14973);
or U15929 (N_15929,N_14722,N_14887);
nor U15930 (N_15930,N_14270,N_14804);
xor U15931 (N_15931,N_14795,N_14458);
and U15932 (N_15932,N_14000,N_14599);
nor U15933 (N_15933,N_14401,N_14086);
nand U15934 (N_15934,N_14177,N_14030);
and U15935 (N_15935,N_14078,N_14261);
or U15936 (N_15936,N_14512,N_14850);
nor U15937 (N_15937,N_14074,N_14605);
or U15938 (N_15938,N_14181,N_14396);
nor U15939 (N_15939,N_14969,N_14032);
and U15940 (N_15940,N_14705,N_14578);
xnor U15941 (N_15941,N_14392,N_14023);
xnor U15942 (N_15942,N_14721,N_14506);
nor U15943 (N_15943,N_14202,N_14574);
nand U15944 (N_15944,N_14563,N_14660);
nand U15945 (N_15945,N_14445,N_14092);
or U15946 (N_15946,N_14556,N_14842);
nor U15947 (N_15947,N_14176,N_14373);
or U15948 (N_15948,N_14717,N_14407);
or U15949 (N_15949,N_14494,N_14232);
or U15950 (N_15950,N_14986,N_14211);
and U15951 (N_15951,N_14579,N_14138);
or U15952 (N_15952,N_14146,N_14820);
nor U15953 (N_15953,N_14021,N_14922);
or U15954 (N_15954,N_14457,N_14109);
or U15955 (N_15955,N_14409,N_14044);
xnor U15956 (N_15956,N_14320,N_14066);
nor U15957 (N_15957,N_14289,N_14506);
and U15958 (N_15958,N_14866,N_14847);
or U15959 (N_15959,N_14721,N_14697);
or U15960 (N_15960,N_14238,N_14307);
or U15961 (N_15961,N_14883,N_14402);
or U15962 (N_15962,N_14882,N_14642);
nand U15963 (N_15963,N_14153,N_14038);
nor U15964 (N_15964,N_14326,N_14870);
and U15965 (N_15965,N_14755,N_14432);
and U15966 (N_15966,N_14274,N_14356);
nand U15967 (N_15967,N_14456,N_14338);
nand U15968 (N_15968,N_14043,N_14445);
and U15969 (N_15969,N_14715,N_14081);
and U15970 (N_15970,N_14590,N_14594);
or U15971 (N_15971,N_14069,N_14489);
or U15972 (N_15972,N_14120,N_14151);
nand U15973 (N_15973,N_14415,N_14237);
nand U15974 (N_15974,N_14495,N_14949);
xnor U15975 (N_15975,N_14695,N_14010);
and U15976 (N_15976,N_14749,N_14644);
nand U15977 (N_15977,N_14878,N_14710);
or U15978 (N_15978,N_14246,N_14638);
or U15979 (N_15979,N_14876,N_14956);
nor U15980 (N_15980,N_14657,N_14973);
and U15981 (N_15981,N_14720,N_14861);
and U15982 (N_15982,N_14514,N_14284);
nor U15983 (N_15983,N_14762,N_14425);
nor U15984 (N_15984,N_14897,N_14333);
nor U15985 (N_15985,N_14765,N_14035);
and U15986 (N_15986,N_14706,N_14587);
and U15987 (N_15987,N_14611,N_14921);
nand U15988 (N_15988,N_14564,N_14891);
nand U15989 (N_15989,N_14565,N_14244);
xor U15990 (N_15990,N_14592,N_14761);
and U15991 (N_15991,N_14092,N_14685);
nor U15992 (N_15992,N_14161,N_14719);
or U15993 (N_15993,N_14496,N_14244);
or U15994 (N_15994,N_14636,N_14575);
nor U15995 (N_15995,N_14537,N_14565);
nand U15996 (N_15996,N_14173,N_14751);
and U15997 (N_15997,N_14594,N_14462);
and U15998 (N_15998,N_14806,N_14127);
or U15999 (N_15999,N_14196,N_14726);
and U16000 (N_16000,N_15032,N_15282);
nand U16001 (N_16001,N_15676,N_15996);
and U16002 (N_16002,N_15432,N_15056);
nand U16003 (N_16003,N_15465,N_15208);
or U16004 (N_16004,N_15808,N_15659);
xor U16005 (N_16005,N_15956,N_15289);
or U16006 (N_16006,N_15527,N_15174);
nand U16007 (N_16007,N_15256,N_15895);
nand U16008 (N_16008,N_15684,N_15169);
nand U16009 (N_16009,N_15078,N_15991);
or U16010 (N_16010,N_15495,N_15955);
or U16011 (N_16011,N_15624,N_15625);
nand U16012 (N_16012,N_15013,N_15711);
xnor U16013 (N_16013,N_15091,N_15209);
nor U16014 (N_16014,N_15845,N_15016);
and U16015 (N_16015,N_15844,N_15574);
or U16016 (N_16016,N_15482,N_15747);
nand U16017 (N_16017,N_15558,N_15001);
or U16018 (N_16018,N_15542,N_15366);
or U16019 (N_16019,N_15930,N_15245);
and U16020 (N_16020,N_15925,N_15132);
and U16021 (N_16021,N_15769,N_15846);
nand U16022 (N_16022,N_15860,N_15553);
nor U16023 (N_16023,N_15573,N_15251);
nor U16024 (N_16024,N_15834,N_15405);
nand U16025 (N_16025,N_15678,N_15960);
and U16026 (N_16026,N_15487,N_15488);
nor U16027 (N_16027,N_15997,N_15265);
and U16028 (N_16028,N_15296,N_15621);
and U16029 (N_16029,N_15902,N_15555);
nor U16030 (N_16030,N_15236,N_15445);
nand U16031 (N_16031,N_15517,N_15328);
nand U16032 (N_16032,N_15157,N_15373);
nor U16033 (N_16033,N_15514,N_15655);
nor U16034 (N_16034,N_15752,N_15191);
nand U16035 (N_16035,N_15535,N_15428);
xor U16036 (N_16036,N_15400,N_15258);
nor U16037 (N_16037,N_15184,N_15021);
nand U16038 (N_16038,N_15719,N_15429);
nand U16039 (N_16039,N_15628,N_15789);
nor U16040 (N_16040,N_15604,N_15903);
nand U16041 (N_16041,N_15733,N_15434);
nand U16042 (N_16042,N_15513,N_15440);
and U16043 (N_16043,N_15564,N_15937);
or U16044 (N_16044,N_15461,N_15855);
or U16045 (N_16045,N_15199,N_15315);
or U16046 (N_16046,N_15213,N_15504);
nand U16047 (N_16047,N_15494,N_15350);
nand U16048 (N_16048,N_15252,N_15335);
and U16049 (N_16049,N_15088,N_15283);
or U16050 (N_16050,N_15363,N_15891);
and U16051 (N_16051,N_15919,N_15581);
nand U16052 (N_16052,N_15675,N_15337);
or U16053 (N_16053,N_15850,N_15076);
and U16054 (N_16054,N_15133,N_15051);
xor U16055 (N_16055,N_15302,N_15090);
or U16056 (N_16056,N_15112,N_15129);
nor U16057 (N_16057,N_15582,N_15713);
nand U16058 (N_16058,N_15660,N_15990);
nor U16059 (N_16059,N_15836,N_15444);
nand U16060 (N_16060,N_15475,N_15641);
or U16061 (N_16061,N_15153,N_15830);
or U16062 (N_16062,N_15921,N_15623);
and U16063 (N_16063,N_15222,N_15831);
nand U16064 (N_16064,N_15848,N_15668);
xnor U16065 (N_16065,N_15785,N_15520);
nor U16066 (N_16066,N_15234,N_15339);
nor U16067 (N_16067,N_15230,N_15111);
or U16068 (N_16068,N_15726,N_15094);
nor U16069 (N_16069,N_15261,N_15462);
nor U16070 (N_16070,N_15031,N_15588);
xnor U16071 (N_16071,N_15196,N_15124);
and U16072 (N_16072,N_15687,N_15704);
nor U16073 (N_16073,N_15398,N_15364);
nand U16074 (N_16074,N_15944,N_15647);
nand U16075 (N_16075,N_15097,N_15086);
and U16076 (N_16076,N_15409,N_15198);
and U16077 (N_16077,N_15320,N_15454);
nand U16078 (N_16078,N_15083,N_15767);
xor U16079 (N_16079,N_15970,N_15994);
nor U16080 (N_16080,N_15092,N_15468);
or U16081 (N_16081,N_15110,N_15404);
nand U16082 (N_16082,N_15765,N_15382);
nor U16083 (N_16083,N_15596,N_15880);
and U16084 (N_16084,N_15269,N_15499);
nor U16085 (N_16085,N_15701,N_15244);
and U16086 (N_16086,N_15760,N_15182);
and U16087 (N_16087,N_15414,N_15722);
or U16088 (N_16088,N_15065,N_15672);
nand U16089 (N_16089,N_15390,N_15699);
or U16090 (N_16090,N_15598,N_15763);
nand U16091 (N_16091,N_15489,N_15976);
nor U16092 (N_16092,N_15346,N_15501);
nor U16093 (N_16093,N_15000,N_15703);
and U16094 (N_16094,N_15332,N_15591);
nand U16095 (N_16095,N_15290,N_15833);
or U16096 (N_16096,N_15962,N_15368);
xor U16097 (N_16097,N_15317,N_15464);
xnor U16098 (N_16098,N_15419,N_15240);
nor U16099 (N_16099,N_15353,N_15562);
nor U16100 (N_16100,N_15478,N_15927);
and U16101 (N_16101,N_15255,N_15399);
and U16102 (N_16102,N_15149,N_15139);
or U16103 (N_16103,N_15497,N_15805);
nor U16104 (N_16104,N_15786,N_15305);
nand U16105 (N_16105,N_15045,N_15951);
nand U16106 (N_16106,N_15904,N_15796);
or U16107 (N_16107,N_15941,N_15273);
and U16108 (N_16108,N_15274,N_15742);
xnor U16109 (N_16109,N_15971,N_15714);
nor U16110 (N_16110,N_15246,N_15579);
or U16111 (N_16111,N_15532,N_15540);
or U16112 (N_16112,N_15757,N_15349);
nand U16113 (N_16113,N_15220,N_15635);
or U16114 (N_16114,N_15841,N_15663);
and U16115 (N_16115,N_15677,N_15972);
and U16116 (N_16116,N_15068,N_15797);
nand U16117 (N_16117,N_15717,N_15916);
or U16118 (N_16118,N_15686,N_15616);
nand U16119 (N_16119,N_15826,N_15248);
and U16120 (N_16120,N_15818,N_15882);
nor U16121 (N_16121,N_15073,N_15259);
and U16122 (N_16122,N_15508,N_15799);
and U16123 (N_16123,N_15963,N_15197);
nor U16124 (N_16124,N_15662,N_15568);
xnor U16125 (N_16125,N_15226,N_15351);
xor U16126 (N_16126,N_15721,N_15879);
or U16127 (N_16127,N_15044,N_15416);
or U16128 (N_16128,N_15551,N_15069);
nor U16129 (N_16129,N_15740,N_15896);
nand U16130 (N_16130,N_15384,N_15819);
nand U16131 (N_16131,N_15036,N_15585);
nand U16132 (N_16132,N_15840,N_15657);
or U16133 (N_16133,N_15365,N_15378);
nor U16134 (N_16134,N_15141,N_15566);
nand U16135 (N_16135,N_15062,N_15122);
and U16136 (N_16136,N_15974,N_15518);
nand U16137 (N_16137,N_15874,N_15753);
or U16138 (N_16138,N_15887,N_15295);
and U16139 (N_16139,N_15696,N_15225);
nor U16140 (N_16140,N_15838,N_15093);
nand U16141 (N_16141,N_15357,N_15966);
and U16142 (N_16142,N_15355,N_15533);
xor U16143 (N_16143,N_15820,N_15734);
nor U16144 (N_16144,N_15233,N_15803);
nand U16145 (N_16145,N_15374,N_15807);
nor U16146 (N_16146,N_15082,N_15651);
and U16147 (N_16147,N_15402,N_15691);
and U16148 (N_16148,N_15643,N_15053);
xnor U16149 (N_16149,N_15529,N_15777);
and U16150 (N_16150,N_15816,N_15938);
nor U16151 (N_16151,N_15606,N_15783);
xor U16152 (N_16152,N_15388,N_15219);
and U16153 (N_16153,N_15430,N_15125);
and U16154 (N_16154,N_15254,N_15424);
nor U16155 (N_16155,N_15814,N_15089);
and U16156 (N_16156,N_15872,N_15716);
and U16157 (N_16157,N_15652,N_15449);
or U16158 (N_16158,N_15864,N_15381);
and U16159 (N_16159,N_15999,N_15135);
or U16160 (N_16160,N_15193,N_15017);
nor U16161 (N_16161,N_15544,N_15324);
nand U16162 (N_16162,N_15806,N_15291);
nand U16163 (N_16163,N_15035,N_15521);
nand U16164 (N_16164,N_15018,N_15952);
and U16165 (N_16165,N_15341,N_15866);
nor U16166 (N_16166,N_15165,N_15791);
and U16167 (N_16167,N_15048,N_15561);
nand U16168 (N_16168,N_15050,N_15969);
nand U16169 (N_16169,N_15476,N_15026);
nand U16170 (N_16170,N_15171,N_15206);
and U16171 (N_16171,N_15654,N_15644);
and U16172 (N_16172,N_15988,N_15859);
or U16173 (N_16173,N_15762,N_15695);
or U16174 (N_16174,N_15656,N_15801);
and U16175 (N_16175,N_15728,N_15965);
or U16176 (N_16176,N_15812,N_15474);
nand U16177 (N_16177,N_15204,N_15731);
and U16178 (N_16178,N_15195,N_15912);
xor U16179 (N_16179,N_15002,N_15602);
nor U16180 (N_16180,N_15718,N_15372);
and U16181 (N_16181,N_15415,N_15732);
and U16182 (N_16182,N_15739,N_15237);
nand U16183 (N_16183,N_15027,N_15639);
and U16184 (N_16184,N_15493,N_15995);
and U16185 (N_16185,N_15485,N_15940);
nand U16186 (N_16186,N_15189,N_15427);
and U16187 (N_16187,N_15298,N_15804);
or U16188 (N_16188,N_15809,N_15072);
nor U16189 (N_16189,N_15375,N_15817);
xor U16190 (N_16190,N_15933,N_15539);
xnor U16191 (N_16191,N_15205,N_15853);
or U16192 (N_16192,N_15126,N_15435);
nand U16193 (N_16193,N_15115,N_15705);
or U16194 (N_16194,N_15342,N_15674);
nand U16195 (N_16195,N_15395,N_15594);
and U16196 (N_16196,N_15438,N_15232);
nand U16197 (N_16197,N_15473,N_15109);
nor U16198 (N_16198,N_15263,N_15217);
nand U16199 (N_16199,N_15058,N_15852);
and U16200 (N_16200,N_15610,N_15778);
or U16201 (N_16201,N_15839,N_15934);
nand U16202 (N_16202,N_15707,N_15064);
or U16203 (N_16203,N_15978,N_15500);
and U16204 (N_16204,N_15280,N_15330);
nand U16205 (N_16205,N_15505,N_15619);
nand U16206 (N_16206,N_15312,N_15385);
or U16207 (N_16207,N_15067,N_15446);
xor U16208 (N_16208,N_15229,N_15710);
and U16209 (N_16209,N_15890,N_15557);
or U16210 (N_16210,N_15570,N_15509);
nor U16211 (N_16211,N_15571,N_15775);
nand U16212 (N_16212,N_15671,N_15774);
and U16213 (N_16213,N_15877,N_15743);
nor U16214 (N_16214,N_15615,N_15892);
nand U16215 (N_16215,N_15851,N_15242);
and U16216 (N_16216,N_15583,N_15525);
and U16217 (N_16217,N_15422,N_15979);
or U16218 (N_16218,N_15413,N_15608);
and U16219 (N_16219,N_15463,N_15913);
or U16220 (N_16220,N_15356,N_15792);
or U16221 (N_16221,N_15071,N_15723);
and U16222 (N_16222,N_15689,N_15100);
and U16223 (N_16223,N_15159,N_15523);
nand U16224 (N_16224,N_15648,N_15709);
nand U16225 (N_16225,N_15943,N_15620);
nand U16226 (N_16226,N_15469,N_15957);
xor U16227 (N_16227,N_15528,N_15288);
xnor U16228 (N_16228,N_15099,N_15649);
nor U16229 (N_16229,N_15175,N_15712);
nor U16230 (N_16230,N_15776,N_15854);
or U16231 (N_16231,N_15004,N_15824);
nor U16232 (N_16232,N_15745,N_15055);
and U16233 (N_16233,N_15294,N_15140);
or U16234 (N_16234,N_15790,N_15168);
nor U16235 (N_16235,N_15599,N_15322);
and U16236 (N_16236,N_15340,N_15549);
nand U16237 (N_16237,N_15006,N_15188);
and U16238 (N_16238,N_15210,N_15172);
nand U16239 (N_16239,N_15681,N_15759);
or U16240 (N_16240,N_15466,N_15052);
and U16241 (N_16241,N_15862,N_15151);
nand U16242 (N_16242,N_15005,N_15572);
nor U16243 (N_16243,N_15143,N_15560);
xnor U16244 (N_16244,N_15456,N_15683);
nand U16245 (N_16245,N_15034,N_15452);
or U16246 (N_16246,N_15128,N_15267);
or U16247 (N_16247,N_15074,N_15603);
and U16248 (N_16248,N_15391,N_15313);
nand U16249 (N_16249,N_15441,N_15386);
and U16250 (N_16250,N_15595,N_15418);
nand U16251 (N_16251,N_15486,N_15519);
nor U16252 (N_16252,N_15737,N_15827);
nand U16253 (N_16253,N_15609,N_15334);
xnor U16254 (N_16254,N_15632,N_15347);
or U16255 (N_16255,N_15284,N_15578);
or U16256 (N_16256,N_15228,N_15116);
and U16257 (N_16257,N_15865,N_15344);
and U16258 (N_16258,N_15479,N_15144);
and U16259 (N_16259,N_15694,N_15439);
xor U16260 (N_16260,N_15319,N_15764);
nand U16261 (N_16261,N_15811,N_15915);
xor U16262 (N_16262,N_15370,N_15531);
and U16263 (N_16263,N_15047,N_15876);
and U16264 (N_16264,N_15243,N_15155);
nand U16265 (N_16265,N_15936,N_15019);
nor U16266 (N_16266,N_15888,N_15973);
nor U16267 (N_16267,N_15271,N_15190);
nor U16268 (N_16268,N_15396,N_15868);
and U16269 (N_16269,N_15627,N_15387);
and U16270 (N_16270,N_15918,N_15307);
nand U16271 (N_16271,N_15618,N_15024);
and U16272 (N_16272,N_15455,N_15642);
nor U16273 (N_16273,N_15362,N_15114);
and U16274 (N_16274,N_15448,N_15148);
and U16275 (N_16275,N_15761,N_15343);
nand U16276 (N_16276,N_15407,N_15967);
nand U16277 (N_16277,N_15645,N_15498);
and U16278 (N_16278,N_15301,N_15040);
nor U16279 (N_16279,N_15985,N_15325);
and U16280 (N_16280,N_15526,N_15569);
nand U16281 (N_16281,N_15946,N_15054);
or U16282 (N_16282,N_15276,N_15829);
nor U16283 (N_16283,N_15688,N_15867);
and U16284 (N_16284,N_15984,N_15942);
and U16285 (N_16285,N_15898,N_15300);
or U16286 (N_16286,N_15425,N_15730);
nand U16287 (N_16287,N_15308,N_15950);
or U16288 (N_16288,N_15137,N_15336);
or U16289 (N_16289,N_15238,N_15629);
nand U16290 (N_16290,N_15700,N_15393);
or U16291 (N_16291,N_15630,N_15795);
and U16292 (N_16292,N_15008,N_15828);
xor U16293 (N_16293,N_15412,N_15345);
nor U16294 (N_16294,N_15939,N_15534);
and U16295 (N_16295,N_15889,N_15870);
and U16296 (N_16296,N_15861,N_15613);
and U16297 (N_16297,N_15057,N_15751);
and U16298 (N_16298,N_15247,N_15239);
nor U16299 (N_16299,N_15593,N_15450);
or U16300 (N_16300,N_15471,N_15536);
nand U16301 (N_16301,N_15297,N_15857);
and U16302 (N_16302,N_15741,N_15164);
and U16303 (N_16303,N_15426,N_15309);
and U16304 (N_16304,N_15161,N_15772);
and U16305 (N_16305,N_15843,N_15788);
and U16306 (N_16306,N_15748,N_15964);
nor U16307 (N_16307,N_15029,N_15279);
xor U16308 (N_16308,N_15359,N_15025);
or U16309 (N_16309,N_15924,N_15156);
and U16310 (N_16310,N_15945,N_15634);
nor U16311 (N_16311,N_15079,N_15264);
or U16312 (N_16312,N_15975,N_15186);
and U16313 (N_16313,N_15825,N_15947);
nor U16314 (N_16314,N_15215,N_15200);
nand U16315 (N_16315,N_15154,N_15235);
nand U16316 (N_16316,N_15117,N_15060);
and U16317 (N_16317,N_15886,N_15147);
and U16318 (N_16318,N_15081,N_15881);
nand U16319 (N_16319,N_15272,N_15163);
or U16320 (N_16320,N_15545,N_15884);
nand U16321 (N_16321,N_15266,N_15477);
nand U16322 (N_16322,N_15420,N_15007);
or U16323 (N_16323,N_15022,N_15626);
and U16324 (N_16324,N_15953,N_15037);
nand U16325 (N_16325,N_15589,N_15858);
and U16326 (N_16326,N_15253,N_15401);
and U16327 (N_16327,N_15736,N_15311);
nand U16328 (N_16328,N_15869,N_15262);
or U16329 (N_16329,N_15910,N_15192);
nand U16330 (N_16330,N_15697,N_15453);
xnor U16331 (N_16331,N_15331,N_15959);
xor U16332 (N_16332,N_15813,N_15798);
nor U16333 (N_16333,N_15397,N_15637);
or U16334 (N_16334,N_15510,N_15842);
nor U16335 (N_16335,N_15436,N_15431);
nor U16336 (N_16336,N_15152,N_15685);
xnor U16337 (N_16337,N_15323,N_15906);
nand U16338 (N_16338,N_15287,N_15231);
or U16339 (N_16339,N_15693,N_15666);
nor U16340 (N_16340,N_15667,N_15077);
or U16341 (N_16341,N_15640,N_15856);
nand U16342 (N_16342,N_15015,N_15490);
nor U16343 (N_16343,N_15556,N_15358);
or U16344 (N_16344,N_15746,N_15905);
and U16345 (N_16345,N_15878,N_15389);
and U16346 (N_16346,N_15920,N_15014);
nor U16347 (N_16347,N_15756,N_15376);
xor U16348 (N_16348,N_15166,N_15720);
or U16349 (N_16349,N_15038,N_15367);
nor U16350 (N_16350,N_15622,N_15281);
nor U16351 (N_16351,N_15983,N_15847);
nor U16352 (N_16352,N_15075,N_15692);
nand U16353 (N_16353,N_15729,N_15780);
xor U16354 (N_16354,N_15607,N_15121);
and U16355 (N_16355,N_15958,N_15770);
nor U16356 (N_16356,N_15961,N_15894);
nor U16357 (N_16357,N_15897,N_15749);
and U16358 (N_16358,N_15216,N_15929);
and U16359 (N_16359,N_15802,N_15650);
nand U16360 (N_16360,N_15664,N_15554);
nand U16361 (N_16361,N_15102,N_15515);
or U16362 (N_16362,N_15145,N_15981);
nand U16363 (N_16363,N_15547,N_15725);
or U16364 (N_16364,N_15020,N_15059);
or U16365 (N_16365,N_15914,N_15530);
and U16366 (N_16366,N_15443,N_15104);
nor U16367 (N_16367,N_15278,N_15113);
and U16368 (N_16368,N_15863,N_15522);
nor U16369 (N_16369,N_15754,N_15948);
nor U16370 (N_16370,N_15212,N_15931);
or U16371 (N_16371,N_15541,N_15011);
nor U16372 (N_16372,N_15457,N_15750);
nand U16373 (N_16373,N_15636,N_15046);
xor U16374 (N_16374,N_15241,N_15010);
nor U16375 (N_16375,N_15543,N_15131);
and U16376 (N_16376,N_15275,N_15218);
nor U16377 (N_16377,N_15548,N_15755);
nor U16378 (N_16378,N_15080,N_15782);
or U16379 (N_16379,N_15333,N_15875);
and U16380 (N_16380,N_15160,N_15326);
or U16381 (N_16381,N_15360,N_15986);
or U16382 (N_16382,N_15822,N_15907);
nor U16383 (N_16383,N_15576,N_15923);
or U16384 (N_16384,N_15631,N_15917);
and U16385 (N_16385,N_15392,N_15181);
xnor U16386 (N_16386,N_15658,N_15039);
or U16387 (N_16387,N_15134,N_15665);
and U16388 (N_16388,N_15552,N_15614);
nor U16389 (N_16389,N_15977,N_15257);
or U16390 (N_16390,N_15095,N_15771);
nand U16391 (N_16391,N_15185,N_15661);
or U16392 (N_16392,N_15584,N_15577);
or U16393 (N_16393,N_15524,N_15823);
nand U16394 (N_16394,N_15177,N_15442);
nand U16395 (N_16395,N_15041,N_15118);
nor U16396 (N_16396,N_15794,N_15009);
or U16397 (N_16397,N_15893,N_15277);
and U16398 (N_16398,N_15546,N_15070);
nor U16399 (N_16399,N_15849,N_15180);
and U16400 (N_16400,N_15162,N_15690);
nand U16401 (N_16401,N_15706,N_15087);
and U16402 (N_16402,N_15480,N_15030);
or U16403 (N_16403,N_15327,N_15063);
or U16404 (N_16404,N_15421,N_15835);
xnor U16405 (N_16405,N_15638,N_15909);
nand U16406 (N_16406,N_15911,N_15987);
or U16407 (N_16407,N_15680,N_15481);
and U16408 (N_16408,N_15187,N_15098);
nor U16409 (N_16409,N_15871,N_15066);
nand U16410 (N_16410,N_15176,N_15601);
and U16411 (N_16411,N_15033,N_15669);
and U16412 (N_16412,N_15227,N_15735);
nand U16413 (N_16413,N_15101,N_15394);
nand U16414 (N_16414,N_15928,N_15178);
xnor U16415 (N_16415,N_15460,N_15538);
or U16416 (N_16416,N_15968,N_15354);
nor U16417 (N_16417,N_15106,N_15800);
and U16418 (N_16418,N_15484,N_15214);
or U16419 (N_16419,N_15611,N_15361);
xnor U16420 (N_16420,N_15511,N_15567);
or U16421 (N_16421,N_15433,N_15592);
xor U16422 (N_16422,N_15586,N_15314);
nor U16423 (N_16423,N_15837,N_15491);
nor U16424 (N_16424,N_15003,N_15982);
nor U16425 (N_16425,N_15096,N_15023);
and U16426 (N_16426,N_15459,N_15908);
nand U16427 (N_16427,N_15467,N_15646);
nand U16428 (N_16428,N_15673,N_15377);
nand U16429 (N_16429,N_15268,N_15506);
and U16430 (N_16430,N_15173,N_15992);
and U16431 (N_16431,N_15348,N_15369);
nand U16432 (N_16432,N_15224,N_15084);
xor U16433 (N_16433,N_15167,N_15316);
or U16434 (N_16434,N_15612,N_15049);
and U16435 (N_16435,N_15221,N_15458);
or U16436 (N_16436,N_15105,N_15285);
nand U16437 (N_16437,N_15380,N_15885);
and U16438 (N_16438,N_15781,N_15158);
nor U16439 (N_16439,N_15423,N_15451);
or U16440 (N_16440,N_15411,N_15304);
xor U16441 (N_16441,N_15123,N_15119);
nor U16442 (N_16442,N_15136,N_15873);
nor U16443 (N_16443,N_15203,N_15043);
nand U16444 (N_16444,N_15447,N_15142);
nor U16445 (N_16445,N_15922,N_15507);
or U16446 (N_16446,N_15403,N_15286);
xnor U16447 (N_16447,N_15042,N_15698);
or U16448 (N_16448,N_15926,N_15103);
and U16449 (N_16449,N_15299,N_15954);
nand U16450 (N_16450,N_15516,N_15223);
nor U16451 (N_16451,N_15787,N_15012);
nor U16452 (N_16452,N_15550,N_15492);
nor U16453 (N_16453,N_15900,N_15779);
nand U16454 (N_16454,N_15194,N_15605);
xnor U16455 (N_16455,N_15653,N_15179);
nand U16456 (N_16456,N_15496,N_15587);
and U16457 (N_16457,N_15183,N_15310);
nand U16458 (N_16458,N_15437,N_15883);
nand U16459 (N_16459,N_15170,N_15633);
nor U16460 (N_16460,N_15130,N_15702);
nor U16461 (N_16461,N_15207,N_15682);
xor U16462 (N_16462,N_15408,N_15138);
nor U16463 (N_16463,N_15832,N_15590);
or U16464 (N_16464,N_15670,N_15768);
nand U16465 (N_16465,N_15949,N_15303);
and U16466 (N_16466,N_15901,N_15993);
and U16467 (N_16467,N_15406,N_15932);
nand U16468 (N_16468,N_15371,N_15108);
and U16469 (N_16469,N_15410,N_15318);
nand U16470 (N_16470,N_15338,N_15085);
nand U16471 (N_16471,N_15899,N_15028);
nor U16472 (N_16472,N_15483,N_15744);
xor U16473 (N_16473,N_15150,N_15211);
or U16474 (N_16474,N_15470,N_15306);
and U16475 (N_16475,N_15250,N_15503);
and U16476 (N_16476,N_15810,N_15270);
or U16477 (N_16477,N_15249,N_15472);
or U16478 (N_16478,N_15352,N_15715);
and U16479 (N_16479,N_15260,N_15815);
nor U16480 (N_16480,N_15597,N_15575);
and U16481 (N_16481,N_15998,N_15793);
and U16482 (N_16482,N_15559,N_15758);
or U16483 (N_16483,N_15512,N_15821);
nor U16484 (N_16484,N_15679,N_15935);
nor U16485 (N_16485,N_15727,N_15766);
xnor U16486 (N_16486,N_15292,N_15563);
nor U16487 (N_16487,N_15120,N_15329);
and U16488 (N_16488,N_15537,N_15724);
nor U16489 (N_16489,N_15600,N_15417);
nor U16490 (N_16490,N_15293,N_15321);
and U16491 (N_16491,N_15565,N_15502);
or U16492 (N_16492,N_15784,N_15383);
nor U16493 (N_16493,N_15201,N_15773);
and U16494 (N_16494,N_15127,N_15202);
nand U16495 (N_16495,N_15061,N_15738);
nand U16496 (N_16496,N_15989,N_15379);
nand U16497 (N_16497,N_15107,N_15580);
and U16498 (N_16498,N_15708,N_15617);
nand U16499 (N_16499,N_15146,N_15980);
or U16500 (N_16500,N_15102,N_15555);
or U16501 (N_16501,N_15507,N_15878);
nor U16502 (N_16502,N_15382,N_15984);
nand U16503 (N_16503,N_15991,N_15150);
nor U16504 (N_16504,N_15198,N_15927);
nor U16505 (N_16505,N_15609,N_15089);
and U16506 (N_16506,N_15078,N_15772);
nand U16507 (N_16507,N_15850,N_15509);
nand U16508 (N_16508,N_15462,N_15202);
and U16509 (N_16509,N_15668,N_15089);
and U16510 (N_16510,N_15548,N_15855);
or U16511 (N_16511,N_15506,N_15483);
or U16512 (N_16512,N_15884,N_15029);
nand U16513 (N_16513,N_15638,N_15035);
nor U16514 (N_16514,N_15160,N_15705);
xor U16515 (N_16515,N_15840,N_15855);
nand U16516 (N_16516,N_15464,N_15182);
and U16517 (N_16517,N_15137,N_15520);
nand U16518 (N_16518,N_15842,N_15626);
nand U16519 (N_16519,N_15763,N_15804);
and U16520 (N_16520,N_15469,N_15690);
or U16521 (N_16521,N_15717,N_15344);
nand U16522 (N_16522,N_15338,N_15380);
or U16523 (N_16523,N_15834,N_15631);
xor U16524 (N_16524,N_15014,N_15770);
and U16525 (N_16525,N_15787,N_15926);
nor U16526 (N_16526,N_15968,N_15952);
nand U16527 (N_16527,N_15539,N_15186);
or U16528 (N_16528,N_15996,N_15633);
nand U16529 (N_16529,N_15664,N_15283);
nor U16530 (N_16530,N_15466,N_15293);
nor U16531 (N_16531,N_15095,N_15602);
nand U16532 (N_16532,N_15569,N_15337);
nand U16533 (N_16533,N_15081,N_15730);
and U16534 (N_16534,N_15967,N_15483);
or U16535 (N_16535,N_15581,N_15394);
nor U16536 (N_16536,N_15025,N_15026);
and U16537 (N_16537,N_15474,N_15939);
and U16538 (N_16538,N_15247,N_15853);
nand U16539 (N_16539,N_15303,N_15215);
xor U16540 (N_16540,N_15404,N_15458);
nand U16541 (N_16541,N_15766,N_15547);
nor U16542 (N_16542,N_15533,N_15149);
and U16543 (N_16543,N_15970,N_15368);
nor U16544 (N_16544,N_15648,N_15272);
and U16545 (N_16545,N_15007,N_15035);
nor U16546 (N_16546,N_15462,N_15842);
and U16547 (N_16547,N_15951,N_15233);
nor U16548 (N_16548,N_15947,N_15648);
nand U16549 (N_16549,N_15411,N_15813);
xnor U16550 (N_16550,N_15530,N_15160);
or U16551 (N_16551,N_15848,N_15659);
or U16552 (N_16552,N_15751,N_15314);
and U16553 (N_16553,N_15047,N_15557);
nor U16554 (N_16554,N_15814,N_15147);
nand U16555 (N_16555,N_15508,N_15630);
nand U16556 (N_16556,N_15115,N_15539);
and U16557 (N_16557,N_15681,N_15064);
nor U16558 (N_16558,N_15376,N_15829);
and U16559 (N_16559,N_15060,N_15842);
nor U16560 (N_16560,N_15794,N_15582);
xnor U16561 (N_16561,N_15024,N_15881);
nor U16562 (N_16562,N_15588,N_15520);
nor U16563 (N_16563,N_15717,N_15141);
nor U16564 (N_16564,N_15094,N_15651);
nor U16565 (N_16565,N_15973,N_15861);
nand U16566 (N_16566,N_15088,N_15153);
nand U16567 (N_16567,N_15372,N_15185);
and U16568 (N_16568,N_15732,N_15024);
or U16569 (N_16569,N_15963,N_15496);
nor U16570 (N_16570,N_15557,N_15957);
nor U16571 (N_16571,N_15549,N_15811);
and U16572 (N_16572,N_15058,N_15874);
and U16573 (N_16573,N_15414,N_15726);
nand U16574 (N_16574,N_15906,N_15057);
xnor U16575 (N_16575,N_15571,N_15074);
or U16576 (N_16576,N_15652,N_15638);
and U16577 (N_16577,N_15963,N_15428);
nor U16578 (N_16578,N_15706,N_15035);
or U16579 (N_16579,N_15049,N_15654);
nand U16580 (N_16580,N_15012,N_15297);
nand U16581 (N_16581,N_15972,N_15271);
nor U16582 (N_16582,N_15045,N_15263);
or U16583 (N_16583,N_15199,N_15831);
and U16584 (N_16584,N_15724,N_15474);
nor U16585 (N_16585,N_15276,N_15775);
nand U16586 (N_16586,N_15885,N_15733);
or U16587 (N_16587,N_15397,N_15710);
nand U16588 (N_16588,N_15641,N_15854);
nor U16589 (N_16589,N_15762,N_15619);
or U16590 (N_16590,N_15804,N_15451);
and U16591 (N_16591,N_15841,N_15915);
nor U16592 (N_16592,N_15071,N_15701);
or U16593 (N_16593,N_15027,N_15686);
nor U16594 (N_16594,N_15875,N_15749);
and U16595 (N_16595,N_15378,N_15914);
nor U16596 (N_16596,N_15820,N_15596);
or U16597 (N_16597,N_15265,N_15730);
and U16598 (N_16598,N_15947,N_15137);
xor U16599 (N_16599,N_15129,N_15983);
nand U16600 (N_16600,N_15994,N_15120);
xnor U16601 (N_16601,N_15941,N_15331);
nor U16602 (N_16602,N_15015,N_15632);
and U16603 (N_16603,N_15657,N_15022);
nor U16604 (N_16604,N_15243,N_15528);
xnor U16605 (N_16605,N_15160,N_15247);
xor U16606 (N_16606,N_15757,N_15857);
nor U16607 (N_16607,N_15777,N_15950);
and U16608 (N_16608,N_15534,N_15332);
and U16609 (N_16609,N_15438,N_15508);
and U16610 (N_16610,N_15055,N_15814);
nand U16611 (N_16611,N_15721,N_15286);
xor U16612 (N_16612,N_15816,N_15040);
or U16613 (N_16613,N_15160,N_15687);
xor U16614 (N_16614,N_15688,N_15319);
nor U16615 (N_16615,N_15616,N_15510);
or U16616 (N_16616,N_15992,N_15473);
nor U16617 (N_16617,N_15607,N_15554);
nor U16618 (N_16618,N_15161,N_15751);
and U16619 (N_16619,N_15266,N_15112);
and U16620 (N_16620,N_15195,N_15708);
nor U16621 (N_16621,N_15313,N_15518);
nor U16622 (N_16622,N_15987,N_15826);
xor U16623 (N_16623,N_15755,N_15323);
nor U16624 (N_16624,N_15545,N_15067);
xnor U16625 (N_16625,N_15010,N_15376);
nor U16626 (N_16626,N_15788,N_15366);
or U16627 (N_16627,N_15098,N_15452);
xnor U16628 (N_16628,N_15711,N_15004);
or U16629 (N_16629,N_15722,N_15327);
and U16630 (N_16630,N_15734,N_15547);
or U16631 (N_16631,N_15941,N_15740);
and U16632 (N_16632,N_15459,N_15519);
or U16633 (N_16633,N_15925,N_15897);
xor U16634 (N_16634,N_15336,N_15475);
xor U16635 (N_16635,N_15768,N_15910);
nor U16636 (N_16636,N_15702,N_15717);
nand U16637 (N_16637,N_15900,N_15234);
xnor U16638 (N_16638,N_15967,N_15947);
nor U16639 (N_16639,N_15856,N_15144);
or U16640 (N_16640,N_15310,N_15341);
nor U16641 (N_16641,N_15052,N_15479);
or U16642 (N_16642,N_15282,N_15856);
nand U16643 (N_16643,N_15093,N_15754);
xnor U16644 (N_16644,N_15251,N_15030);
or U16645 (N_16645,N_15405,N_15111);
nand U16646 (N_16646,N_15181,N_15567);
and U16647 (N_16647,N_15412,N_15133);
xnor U16648 (N_16648,N_15819,N_15111);
or U16649 (N_16649,N_15886,N_15553);
nand U16650 (N_16650,N_15196,N_15664);
xnor U16651 (N_16651,N_15695,N_15838);
and U16652 (N_16652,N_15066,N_15440);
and U16653 (N_16653,N_15539,N_15795);
or U16654 (N_16654,N_15198,N_15314);
nand U16655 (N_16655,N_15294,N_15307);
nor U16656 (N_16656,N_15680,N_15280);
or U16657 (N_16657,N_15419,N_15202);
xor U16658 (N_16658,N_15930,N_15180);
xnor U16659 (N_16659,N_15465,N_15988);
nor U16660 (N_16660,N_15095,N_15066);
or U16661 (N_16661,N_15161,N_15336);
xnor U16662 (N_16662,N_15811,N_15443);
nor U16663 (N_16663,N_15271,N_15246);
and U16664 (N_16664,N_15482,N_15966);
nand U16665 (N_16665,N_15519,N_15336);
nand U16666 (N_16666,N_15104,N_15159);
and U16667 (N_16667,N_15481,N_15033);
and U16668 (N_16668,N_15204,N_15007);
xor U16669 (N_16669,N_15292,N_15052);
nand U16670 (N_16670,N_15633,N_15332);
or U16671 (N_16671,N_15224,N_15128);
or U16672 (N_16672,N_15113,N_15421);
and U16673 (N_16673,N_15232,N_15453);
nor U16674 (N_16674,N_15153,N_15523);
nand U16675 (N_16675,N_15213,N_15310);
nor U16676 (N_16676,N_15631,N_15170);
nor U16677 (N_16677,N_15196,N_15448);
nand U16678 (N_16678,N_15947,N_15112);
nand U16679 (N_16679,N_15647,N_15997);
nor U16680 (N_16680,N_15734,N_15246);
nor U16681 (N_16681,N_15109,N_15645);
or U16682 (N_16682,N_15228,N_15413);
and U16683 (N_16683,N_15833,N_15149);
nand U16684 (N_16684,N_15262,N_15889);
or U16685 (N_16685,N_15234,N_15079);
nor U16686 (N_16686,N_15792,N_15287);
nand U16687 (N_16687,N_15482,N_15768);
and U16688 (N_16688,N_15479,N_15266);
xnor U16689 (N_16689,N_15627,N_15083);
xor U16690 (N_16690,N_15503,N_15251);
xor U16691 (N_16691,N_15377,N_15620);
nand U16692 (N_16692,N_15269,N_15558);
xnor U16693 (N_16693,N_15820,N_15424);
or U16694 (N_16694,N_15334,N_15624);
or U16695 (N_16695,N_15914,N_15675);
nor U16696 (N_16696,N_15856,N_15989);
nand U16697 (N_16697,N_15919,N_15930);
nand U16698 (N_16698,N_15262,N_15489);
and U16699 (N_16699,N_15252,N_15205);
nor U16700 (N_16700,N_15065,N_15181);
nor U16701 (N_16701,N_15099,N_15525);
nand U16702 (N_16702,N_15610,N_15023);
nor U16703 (N_16703,N_15061,N_15202);
and U16704 (N_16704,N_15460,N_15879);
or U16705 (N_16705,N_15439,N_15196);
nor U16706 (N_16706,N_15505,N_15850);
or U16707 (N_16707,N_15054,N_15144);
nand U16708 (N_16708,N_15128,N_15618);
nand U16709 (N_16709,N_15255,N_15402);
or U16710 (N_16710,N_15241,N_15337);
or U16711 (N_16711,N_15669,N_15779);
nor U16712 (N_16712,N_15571,N_15163);
or U16713 (N_16713,N_15737,N_15217);
xor U16714 (N_16714,N_15418,N_15120);
or U16715 (N_16715,N_15575,N_15285);
or U16716 (N_16716,N_15823,N_15129);
xnor U16717 (N_16717,N_15489,N_15193);
or U16718 (N_16718,N_15955,N_15973);
nand U16719 (N_16719,N_15543,N_15450);
nand U16720 (N_16720,N_15365,N_15034);
and U16721 (N_16721,N_15965,N_15689);
xnor U16722 (N_16722,N_15585,N_15239);
nor U16723 (N_16723,N_15752,N_15382);
nand U16724 (N_16724,N_15398,N_15566);
nand U16725 (N_16725,N_15165,N_15414);
nand U16726 (N_16726,N_15916,N_15086);
nor U16727 (N_16727,N_15858,N_15146);
nand U16728 (N_16728,N_15238,N_15979);
nand U16729 (N_16729,N_15517,N_15645);
or U16730 (N_16730,N_15353,N_15865);
and U16731 (N_16731,N_15771,N_15109);
nor U16732 (N_16732,N_15315,N_15290);
nor U16733 (N_16733,N_15329,N_15238);
nand U16734 (N_16734,N_15866,N_15813);
nand U16735 (N_16735,N_15139,N_15803);
and U16736 (N_16736,N_15377,N_15601);
nor U16737 (N_16737,N_15038,N_15478);
xor U16738 (N_16738,N_15570,N_15564);
and U16739 (N_16739,N_15151,N_15765);
nor U16740 (N_16740,N_15778,N_15478);
xor U16741 (N_16741,N_15061,N_15032);
or U16742 (N_16742,N_15694,N_15244);
nand U16743 (N_16743,N_15696,N_15061);
or U16744 (N_16744,N_15766,N_15913);
nand U16745 (N_16745,N_15833,N_15673);
nor U16746 (N_16746,N_15756,N_15575);
and U16747 (N_16747,N_15520,N_15540);
nor U16748 (N_16748,N_15427,N_15083);
and U16749 (N_16749,N_15860,N_15600);
nor U16750 (N_16750,N_15196,N_15208);
xnor U16751 (N_16751,N_15221,N_15204);
and U16752 (N_16752,N_15815,N_15629);
nand U16753 (N_16753,N_15345,N_15406);
and U16754 (N_16754,N_15110,N_15309);
and U16755 (N_16755,N_15169,N_15367);
xor U16756 (N_16756,N_15116,N_15005);
nand U16757 (N_16757,N_15980,N_15347);
nand U16758 (N_16758,N_15177,N_15211);
and U16759 (N_16759,N_15155,N_15348);
nand U16760 (N_16760,N_15951,N_15339);
and U16761 (N_16761,N_15330,N_15784);
nand U16762 (N_16762,N_15749,N_15407);
nor U16763 (N_16763,N_15864,N_15140);
xor U16764 (N_16764,N_15965,N_15000);
and U16765 (N_16765,N_15034,N_15127);
nor U16766 (N_16766,N_15464,N_15706);
nor U16767 (N_16767,N_15408,N_15737);
nand U16768 (N_16768,N_15794,N_15220);
or U16769 (N_16769,N_15532,N_15192);
xor U16770 (N_16770,N_15373,N_15312);
nor U16771 (N_16771,N_15845,N_15863);
nand U16772 (N_16772,N_15759,N_15818);
and U16773 (N_16773,N_15055,N_15592);
nand U16774 (N_16774,N_15312,N_15070);
xnor U16775 (N_16775,N_15475,N_15517);
nand U16776 (N_16776,N_15427,N_15038);
or U16777 (N_16777,N_15861,N_15331);
nand U16778 (N_16778,N_15964,N_15777);
and U16779 (N_16779,N_15583,N_15204);
or U16780 (N_16780,N_15920,N_15335);
and U16781 (N_16781,N_15970,N_15738);
or U16782 (N_16782,N_15597,N_15201);
or U16783 (N_16783,N_15295,N_15348);
nor U16784 (N_16784,N_15387,N_15117);
nand U16785 (N_16785,N_15319,N_15680);
or U16786 (N_16786,N_15121,N_15977);
nor U16787 (N_16787,N_15381,N_15528);
nand U16788 (N_16788,N_15444,N_15300);
and U16789 (N_16789,N_15596,N_15415);
and U16790 (N_16790,N_15645,N_15736);
nor U16791 (N_16791,N_15948,N_15929);
and U16792 (N_16792,N_15274,N_15283);
or U16793 (N_16793,N_15516,N_15606);
nor U16794 (N_16794,N_15680,N_15335);
and U16795 (N_16795,N_15720,N_15119);
nor U16796 (N_16796,N_15524,N_15716);
nor U16797 (N_16797,N_15850,N_15804);
and U16798 (N_16798,N_15128,N_15717);
and U16799 (N_16799,N_15649,N_15498);
xnor U16800 (N_16800,N_15701,N_15813);
nor U16801 (N_16801,N_15750,N_15939);
or U16802 (N_16802,N_15490,N_15064);
nor U16803 (N_16803,N_15472,N_15845);
or U16804 (N_16804,N_15656,N_15969);
and U16805 (N_16805,N_15183,N_15710);
nor U16806 (N_16806,N_15148,N_15689);
or U16807 (N_16807,N_15742,N_15159);
or U16808 (N_16808,N_15136,N_15848);
and U16809 (N_16809,N_15552,N_15474);
nor U16810 (N_16810,N_15371,N_15154);
nand U16811 (N_16811,N_15977,N_15489);
and U16812 (N_16812,N_15472,N_15407);
or U16813 (N_16813,N_15006,N_15349);
nor U16814 (N_16814,N_15771,N_15969);
nor U16815 (N_16815,N_15091,N_15504);
nor U16816 (N_16816,N_15159,N_15110);
or U16817 (N_16817,N_15336,N_15497);
or U16818 (N_16818,N_15412,N_15997);
nor U16819 (N_16819,N_15615,N_15195);
and U16820 (N_16820,N_15210,N_15003);
and U16821 (N_16821,N_15339,N_15676);
nand U16822 (N_16822,N_15721,N_15428);
nand U16823 (N_16823,N_15682,N_15811);
xor U16824 (N_16824,N_15768,N_15038);
nor U16825 (N_16825,N_15135,N_15465);
xor U16826 (N_16826,N_15708,N_15183);
nand U16827 (N_16827,N_15681,N_15029);
or U16828 (N_16828,N_15403,N_15889);
and U16829 (N_16829,N_15100,N_15753);
or U16830 (N_16830,N_15282,N_15340);
nor U16831 (N_16831,N_15204,N_15316);
and U16832 (N_16832,N_15124,N_15634);
and U16833 (N_16833,N_15273,N_15935);
nor U16834 (N_16834,N_15212,N_15354);
and U16835 (N_16835,N_15554,N_15978);
nand U16836 (N_16836,N_15410,N_15122);
xnor U16837 (N_16837,N_15380,N_15495);
and U16838 (N_16838,N_15001,N_15946);
nor U16839 (N_16839,N_15013,N_15973);
nor U16840 (N_16840,N_15511,N_15524);
or U16841 (N_16841,N_15740,N_15885);
and U16842 (N_16842,N_15535,N_15548);
or U16843 (N_16843,N_15577,N_15830);
and U16844 (N_16844,N_15934,N_15678);
and U16845 (N_16845,N_15170,N_15253);
or U16846 (N_16846,N_15621,N_15948);
xnor U16847 (N_16847,N_15012,N_15409);
nor U16848 (N_16848,N_15711,N_15901);
nand U16849 (N_16849,N_15767,N_15486);
xnor U16850 (N_16850,N_15987,N_15155);
nor U16851 (N_16851,N_15578,N_15795);
nand U16852 (N_16852,N_15745,N_15465);
and U16853 (N_16853,N_15671,N_15443);
nor U16854 (N_16854,N_15458,N_15951);
and U16855 (N_16855,N_15656,N_15213);
nor U16856 (N_16856,N_15333,N_15393);
or U16857 (N_16857,N_15135,N_15317);
and U16858 (N_16858,N_15026,N_15563);
xor U16859 (N_16859,N_15927,N_15790);
or U16860 (N_16860,N_15321,N_15730);
nor U16861 (N_16861,N_15807,N_15222);
or U16862 (N_16862,N_15392,N_15600);
xor U16863 (N_16863,N_15220,N_15171);
and U16864 (N_16864,N_15376,N_15075);
and U16865 (N_16865,N_15070,N_15355);
and U16866 (N_16866,N_15770,N_15337);
and U16867 (N_16867,N_15398,N_15702);
or U16868 (N_16868,N_15099,N_15329);
and U16869 (N_16869,N_15104,N_15309);
nor U16870 (N_16870,N_15737,N_15071);
and U16871 (N_16871,N_15236,N_15320);
or U16872 (N_16872,N_15722,N_15027);
nor U16873 (N_16873,N_15563,N_15296);
nor U16874 (N_16874,N_15232,N_15185);
nor U16875 (N_16875,N_15775,N_15102);
xor U16876 (N_16876,N_15180,N_15952);
xor U16877 (N_16877,N_15443,N_15004);
nand U16878 (N_16878,N_15287,N_15900);
or U16879 (N_16879,N_15974,N_15005);
nor U16880 (N_16880,N_15933,N_15982);
and U16881 (N_16881,N_15037,N_15801);
and U16882 (N_16882,N_15672,N_15325);
and U16883 (N_16883,N_15352,N_15532);
xnor U16884 (N_16884,N_15996,N_15794);
and U16885 (N_16885,N_15708,N_15833);
nand U16886 (N_16886,N_15614,N_15118);
nor U16887 (N_16887,N_15021,N_15502);
nand U16888 (N_16888,N_15123,N_15772);
nor U16889 (N_16889,N_15003,N_15731);
and U16890 (N_16890,N_15476,N_15025);
nor U16891 (N_16891,N_15000,N_15722);
or U16892 (N_16892,N_15489,N_15966);
nand U16893 (N_16893,N_15522,N_15254);
nor U16894 (N_16894,N_15075,N_15742);
and U16895 (N_16895,N_15334,N_15921);
or U16896 (N_16896,N_15161,N_15342);
nor U16897 (N_16897,N_15023,N_15576);
and U16898 (N_16898,N_15033,N_15443);
or U16899 (N_16899,N_15040,N_15999);
nor U16900 (N_16900,N_15834,N_15433);
nand U16901 (N_16901,N_15692,N_15061);
xnor U16902 (N_16902,N_15302,N_15446);
nand U16903 (N_16903,N_15859,N_15172);
or U16904 (N_16904,N_15060,N_15836);
nor U16905 (N_16905,N_15425,N_15141);
or U16906 (N_16906,N_15826,N_15694);
or U16907 (N_16907,N_15126,N_15892);
nor U16908 (N_16908,N_15344,N_15724);
xnor U16909 (N_16909,N_15285,N_15599);
or U16910 (N_16910,N_15105,N_15595);
or U16911 (N_16911,N_15223,N_15145);
and U16912 (N_16912,N_15345,N_15668);
and U16913 (N_16913,N_15264,N_15498);
nand U16914 (N_16914,N_15170,N_15610);
and U16915 (N_16915,N_15768,N_15928);
nand U16916 (N_16916,N_15048,N_15070);
nand U16917 (N_16917,N_15017,N_15281);
or U16918 (N_16918,N_15515,N_15791);
xnor U16919 (N_16919,N_15007,N_15015);
and U16920 (N_16920,N_15116,N_15584);
nor U16921 (N_16921,N_15657,N_15030);
nor U16922 (N_16922,N_15678,N_15004);
and U16923 (N_16923,N_15984,N_15070);
xor U16924 (N_16924,N_15470,N_15571);
and U16925 (N_16925,N_15780,N_15737);
nor U16926 (N_16926,N_15217,N_15749);
nand U16927 (N_16927,N_15685,N_15941);
and U16928 (N_16928,N_15966,N_15583);
nor U16929 (N_16929,N_15083,N_15649);
nor U16930 (N_16930,N_15410,N_15963);
or U16931 (N_16931,N_15176,N_15201);
or U16932 (N_16932,N_15967,N_15291);
or U16933 (N_16933,N_15365,N_15086);
or U16934 (N_16934,N_15384,N_15498);
nand U16935 (N_16935,N_15936,N_15634);
and U16936 (N_16936,N_15726,N_15531);
or U16937 (N_16937,N_15802,N_15092);
and U16938 (N_16938,N_15941,N_15349);
nor U16939 (N_16939,N_15763,N_15080);
nor U16940 (N_16940,N_15800,N_15203);
nand U16941 (N_16941,N_15215,N_15642);
or U16942 (N_16942,N_15589,N_15780);
or U16943 (N_16943,N_15766,N_15319);
nor U16944 (N_16944,N_15738,N_15370);
xor U16945 (N_16945,N_15454,N_15725);
nand U16946 (N_16946,N_15595,N_15905);
nor U16947 (N_16947,N_15749,N_15405);
or U16948 (N_16948,N_15538,N_15924);
or U16949 (N_16949,N_15032,N_15955);
nand U16950 (N_16950,N_15425,N_15924);
nor U16951 (N_16951,N_15841,N_15724);
or U16952 (N_16952,N_15921,N_15411);
and U16953 (N_16953,N_15472,N_15495);
nor U16954 (N_16954,N_15521,N_15834);
and U16955 (N_16955,N_15710,N_15561);
or U16956 (N_16956,N_15929,N_15204);
nand U16957 (N_16957,N_15425,N_15998);
and U16958 (N_16958,N_15953,N_15271);
or U16959 (N_16959,N_15321,N_15771);
nand U16960 (N_16960,N_15579,N_15619);
nand U16961 (N_16961,N_15145,N_15176);
or U16962 (N_16962,N_15893,N_15412);
nand U16963 (N_16963,N_15948,N_15291);
and U16964 (N_16964,N_15230,N_15213);
and U16965 (N_16965,N_15617,N_15582);
nand U16966 (N_16966,N_15859,N_15276);
or U16967 (N_16967,N_15942,N_15269);
nor U16968 (N_16968,N_15695,N_15194);
or U16969 (N_16969,N_15926,N_15394);
or U16970 (N_16970,N_15786,N_15788);
and U16971 (N_16971,N_15167,N_15105);
xnor U16972 (N_16972,N_15432,N_15804);
and U16973 (N_16973,N_15136,N_15440);
or U16974 (N_16974,N_15748,N_15746);
nand U16975 (N_16975,N_15339,N_15650);
and U16976 (N_16976,N_15202,N_15363);
xnor U16977 (N_16977,N_15557,N_15671);
and U16978 (N_16978,N_15160,N_15555);
and U16979 (N_16979,N_15308,N_15971);
nand U16980 (N_16980,N_15262,N_15263);
and U16981 (N_16981,N_15570,N_15845);
nor U16982 (N_16982,N_15107,N_15505);
nand U16983 (N_16983,N_15052,N_15665);
nand U16984 (N_16984,N_15402,N_15182);
or U16985 (N_16985,N_15616,N_15359);
xor U16986 (N_16986,N_15571,N_15500);
and U16987 (N_16987,N_15337,N_15004);
nor U16988 (N_16988,N_15524,N_15502);
nand U16989 (N_16989,N_15772,N_15636);
or U16990 (N_16990,N_15669,N_15565);
nor U16991 (N_16991,N_15339,N_15965);
or U16992 (N_16992,N_15477,N_15245);
and U16993 (N_16993,N_15426,N_15832);
nand U16994 (N_16994,N_15531,N_15052);
nor U16995 (N_16995,N_15439,N_15927);
nand U16996 (N_16996,N_15752,N_15400);
xor U16997 (N_16997,N_15297,N_15534);
xor U16998 (N_16998,N_15866,N_15507);
or U16999 (N_16999,N_15306,N_15880);
nand U17000 (N_17000,N_16906,N_16045);
xor U17001 (N_17001,N_16099,N_16357);
or U17002 (N_17002,N_16120,N_16915);
and U17003 (N_17003,N_16017,N_16929);
and U17004 (N_17004,N_16966,N_16565);
xor U17005 (N_17005,N_16257,N_16475);
or U17006 (N_17006,N_16215,N_16234);
nand U17007 (N_17007,N_16289,N_16247);
or U17008 (N_17008,N_16599,N_16607);
nand U17009 (N_17009,N_16146,N_16067);
nand U17010 (N_17010,N_16582,N_16135);
nand U17011 (N_17011,N_16974,N_16577);
and U17012 (N_17012,N_16155,N_16388);
or U17013 (N_17013,N_16941,N_16277);
or U17014 (N_17014,N_16191,N_16773);
xnor U17015 (N_17015,N_16212,N_16389);
nor U17016 (N_17016,N_16794,N_16148);
nor U17017 (N_17017,N_16575,N_16503);
and U17018 (N_17018,N_16226,N_16953);
xnor U17019 (N_17019,N_16428,N_16029);
nor U17020 (N_17020,N_16973,N_16827);
nor U17021 (N_17021,N_16819,N_16840);
or U17022 (N_17022,N_16544,N_16442);
nand U17023 (N_17023,N_16649,N_16805);
xnor U17024 (N_17024,N_16139,N_16309);
nand U17025 (N_17025,N_16820,N_16816);
nor U17026 (N_17026,N_16824,N_16458);
and U17027 (N_17027,N_16437,N_16147);
nor U17028 (N_17028,N_16015,N_16101);
or U17029 (N_17029,N_16683,N_16720);
and U17030 (N_17030,N_16573,N_16164);
and U17031 (N_17031,N_16880,N_16087);
and U17032 (N_17032,N_16680,N_16774);
nor U17033 (N_17033,N_16498,N_16625);
or U17034 (N_17034,N_16732,N_16838);
or U17035 (N_17035,N_16763,N_16217);
nor U17036 (N_17036,N_16268,N_16627);
and U17037 (N_17037,N_16374,N_16399);
and U17038 (N_17038,N_16447,N_16008);
xor U17039 (N_17039,N_16831,N_16451);
and U17040 (N_17040,N_16515,N_16343);
and U17041 (N_17041,N_16991,N_16065);
or U17042 (N_17042,N_16651,N_16538);
or U17043 (N_17043,N_16292,N_16679);
and U17044 (N_17044,N_16492,N_16137);
nor U17045 (N_17045,N_16169,N_16982);
or U17046 (N_17046,N_16729,N_16128);
xnor U17047 (N_17047,N_16441,N_16747);
nand U17048 (N_17048,N_16452,N_16282);
or U17049 (N_17049,N_16299,N_16961);
and U17050 (N_17050,N_16020,N_16703);
and U17051 (N_17051,N_16914,N_16295);
nor U17052 (N_17052,N_16330,N_16984);
or U17053 (N_17053,N_16699,N_16211);
or U17054 (N_17054,N_16052,N_16832);
and U17055 (N_17055,N_16843,N_16671);
nand U17056 (N_17056,N_16993,N_16286);
or U17057 (N_17057,N_16193,N_16287);
and U17058 (N_17058,N_16377,N_16409);
or U17059 (N_17059,N_16587,N_16788);
nor U17060 (N_17060,N_16779,N_16957);
and U17061 (N_17061,N_16686,N_16829);
nor U17062 (N_17062,N_16116,N_16163);
and U17063 (N_17063,N_16221,N_16172);
nand U17064 (N_17064,N_16753,N_16631);
or U17065 (N_17065,N_16823,N_16668);
xor U17066 (N_17066,N_16770,N_16010);
and U17067 (N_17067,N_16913,N_16907);
nand U17068 (N_17068,N_16333,N_16460);
and U17069 (N_17069,N_16356,N_16596);
xnor U17070 (N_17070,N_16310,N_16855);
nor U17071 (N_17071,N_16078,N_16902);
nand U17072 (N_17072,N_16734,N_16465);
nor U17073 (N_17073,N_16934,N_16612);
and U17074 (N_17074,N_16250,N_16351);
and U17075 (N_17075,N_16134,N_16537);
nor U17076 (N_17076,N_16195,N_16050);
nor U17077 (N_17077,N_16887,N_16814);
nor U17078 (N_17078,N_16580,N_16383);
xnor U17079 (N_17079,N_16862,N_16856);
or U17080 (N_17080,N_16711,N_16943);
nor U17081 (N_17081,N_16700,N_16690);
or U17082 (N_17082,N_16534,N_16345);
or U17083 (N_17083,N_16509,N_16822);
or U17084 (N_17084,N_16233,N_16329);
and U17085 (N_17085,N_16270,N_16477);
and U17086 (N_17086,N_16549,N_16617);
or U17087 (N_17087,N_16808,N_16661);
xor U17088 (N_17088,N_16893,N_16244);
nand U17089 (N_17089,N_16996,N_16904);
and U17090 (N_17090,N_16117,N_16076);
nor U17091 (N_17091,N_16639,N_16618);
or U17092 (N_17092,N_16103,N_16558);
nor U17093 (N_17093,N_16007,N_16712);
or U17094 (N_17094,N_16884,N_16523);
or U17095 (N_17095,N_16200,N_16157);
or U17096 (N_17096,N_16610,N_16896);
or U17097 (N_17097,N_16983,N_16531);
or U17098 (N_17098,N_16804,N_16886);
and U17099 (N_17099,N_16249,N_16371);
nand U17100 (N_17100,N_16694,N_16153);
and U17101 (N_17101,N_16294,N_16380);
or U17102 (N_17102,N_16293,N_16888);
or U17103 (N_17103,N_16815,N_16072);
or U17104 (N_17104,N_16317,N_16311);
nand U17105 (N_17105,N_16179,N_16279);
nor U17106 (N_17106,N_16208,N_16240);
xor U17107 (N_17107,N_16325,N_16791);
nand U17108 (N_17108,N_16159,N_16266);
xor U17109 (N_17109,N_16574,N_16536);
and U17110 (N_17110,N_16825,N_16021);
xnor U17111 (N_17111,N_16336,N_16263);
nand U17112 (N_17112,N_16992,N_16496);
and U17113 (N_17113,N_16848,N_16821);
nand U17114 (N_17114,N_16059,N_16413);
or U17115 (N_17115,N_16083,N_16977);
or U17116 (N_17116,N_16787,N_16043);
or U17117 (N_17117,N_16946,N_16568);
or U17118 (N_17118,N_16801,N_16528);
xor U17119 (N_17119,N_16497,N_16433);
xnor U17120 (N_17120,N_16173,N_16865);
or U17121 (N_17121,N_16207,N_16707);
and U17122 (N_17122,N_16921,N_16667);
nand U17123 (N_17123,N_16382,N_16901);
or U17124 (N_17124,N_16811,N_16968);
or U17125 (N_17125,N_16201,N_16005);
nand U17126 (N_17126,N_16346,N_16341);
or U17127 (N_17127,N_16404,N_16192);
or U17128 (N_17128,N_16620,N_16889);
or U17129 (N_17129,N_16635,N_16272);
xor U17130 (N_17130,N_16402,N_16571);
nor U17131 (N_17131,N_16924,N_16954);
nand U17132 (N_17132,N_16416,N_16485);
nand U17133 (N_17133,N_16047,N_16459);
nand U17134 (N_17134,N_16364,N_16557);
or U17135 (N_17135,N_16533,N_16362);
and U17136 (N_17136,N_16105,N_16669);
and U17137 (N_17137,N_16323,N_16235);
or U17138 (N_17138,N_16259,N_16487);
nand U17139 (N_17139,N_16367,N_16919);
nand U17140 (N_17140,N_16198,N_16600);
or U17141 (N_17141,N_16554,N_16253);
and U17142 (N_17142,N_16303,N_16036);
nand U17143 (N_17143,N_16740,N_16301);
and U17144 (N_17144,N_16425,N_16097);
and U17145 (N_17145,N_16952,N_16644);
and U17146 (N_17146,N_16520,N_16202);
xor U17147 (N_17147,N_16419,N_16813);
nor U17148 (N_17148,N_16062,N_16188);
or U17149 (N_17149,N_16909,N_16931);
and U17150 (N_17150,N_16641,N_16755);
or U17151 (N_17151,N_16353,N_16390);
xor U17152 (N_17152,N_16717,N_16204);
nor U17153 (N_17153,N_16781,N_16181);
and U17154 (N_17154,N_16741,N_16265);
nor U17155 (N_17155,N_16916,N_16115);
and U17156 (N_17156,N_16938,N_16456);
nand U17157 (N_17157,N_16104,N_16632);
or U17158 (N_17158,N_16776,N_16553);
and U17159 (N_17159,N_16489,N_16305);
nand U17160 (N_17160,N_16742,N_16347);
nand U17161 (N_17161,N_16970,N_16567);
nor U17162 (N_17162,N_16276,N_16559);
nand U17163 (N_17163,N_16547,N_16678);
nand U17164 (N_17164,N_16611,N_16189);
and U17165 (N_17165,N_16145,N_16354);
and U17166 (N_17166,N_16307,N_16463);
xor U17167 (N_17167,N_16502,N_16344);
nand U17168 (N_17168,N_16057,N_16950);
nand U17169 (N_17169,N_16339,N_16844);
nor U17170 (N_17170,N_16878,N_16715);
and U17171 (N_17171,N_16972,N_16025);
xnor U17172 (N_17172,N_16006,N_16415);
nor U17173 (N_17173,N_16752,N_16594);
xor U17174 (N_17174,N_16216,N_16900);
nand U17175 (N_17175,N_16174,N_16028);
and U17176 (N_17176,N_16702,N_16312);
xor U17177 (N_17177,N_16422,N_16521);
nand U17178 (N_17178,N_16114,N_16677);
or U17179 (N_17179,N_16803,N_16593);
and U17180 (N_17180,N_16784,N_16236);
nor U17181 (N_17181,N_16942,N_16569);
nand U17182 (N_17182,N_16109,N_16190);
nand U17183 (N_17183,N_16466,N_16255);
nand U17184 (N_17184,N_16876,N_16629);
xnor U17185 (N_17185,N_16060,N_16443);
and U17186 (N_17186,N_16423,N_16508);
nand U17187 (N_17187,N_16845,N_16278);
nand U17188 (N_17188,N_16836,N_16892);
xor U17189 (N_17189,N_16242,N_16472);
nor U17190 (N_17190,N_16424,N_16733);
and U17191 (N_17191,N_16161,N_16370);
and U17192 (N_17192,N_16239,N_16030);
or U17193 (N_17193,N_16910,N_16939);
or U17194 (N_17194,N_16727,N_16857);
xnor U17195 (N_17195,N_16802,N_16512);
or U17196 (N_17196,N_16655,N_16144);
nor U17197 (N_17197,N_16863,N_16918);
or U17198 (N_17198,N_16228,N_16049);
or U17199 (N_17199,N_16879,N_16518);
or U17200 (N_17200,N_16142,N_16895);
or U17201 (N_17201,N_16556,N_16633);
nor U17202 (N_17202,N_16427,N_16967);
nor U17203 (N_17203,N_16187,N_16316);
and U17204 (N_17204,N_16870,N_16360);
or U17205 (N_17205,N_16933,N_16387);
or U17206 (N_17206,N_16483,N_16074);
and U17207 (N_17207,N_16385,N_16348);
nand U17208 (N_17208,N_16578,N_16721);
or U17209 (N_17209,N_16897,N_16042);
and U17210 (N_17210,N_16948,N_16846);
nor U17211 (N_17211,N_16800,N_16051);
or U17212 (N_17212,N_16839,N_16636);
nand U17213 (N_17213,N_16165,N_16665);
or U17214 (N_17214,N_16541,N_16698);
or U17215 (N_17215,N_16602,N_16874);
or U17216 (N_17216,N_16183,N_16697);
xnor U17217 (N_17217,N_16684,N_16724);
nor U17218 (N_17218,N_16118,N_16994);
and U17219 (N_17219,N_16230,N_16737);
nor U17220 (N_17220,N_16156,N_16969);
nand U17221 (N_17221,N_16545,N_16149);
xor U17222 (N_17222,N_16396,N_16407);
and U17223 (N_17223,N_16999,N_16761);
or U17224 (N_17224,N_16053,N_16642);
nor U17225 (N_17225,N_16435,N_16513);
nor U17226 (N_17226,N_16658,N_16936);
or U17227 (N_17227,N_16468,N_16368);
or U17228 (N_17228,N_16524,N_16335);
and U17229 (N_17229,N_16764,N_16622);
nand U17230 (N_17230,N_16760,N_16511);
and U17231 (N_17231,N_16772,N_16754);
nor U17232 (N_17232,N_16517,N_16171);
nor U17233 (N_17233,N_16361,N_16795);
nand U17234 (N_17234,N_16659,N_16003);
nor U17235 (N_17235,N_16797,N_16177);
xnor U17236 (N_17236,N_16759,N_16530);
nand U17237 (N_17237,N_16245,N_16673);
nand U17238 (N_17238,N_16218,N_16762);
and U17239 (N_17239,N_16643,N_16064);
and U17240 (N_17240,N_16735,N_16089);
xnor U17241 (N_17241,N_16670,N_16132);
xnor U17242 (N_17242,N_16350,N_16514);
nand U17243 (N_17243,N_16657,N_16626);
xnor U17244 (N_17244,N_16454,N_16038);
and U17245 (N_17245,N_16340,N_16981);
or U17246 (N_17246,N_16113,N_16584);
and U17247 (N_17247,N_16790,N_16229);
nor U17248 (N_17248,N_16562,N_16860);
and U17249 (N_17249,N_16692,N_16237);
or U17250 (N_17250,N_16778,N_16883);
and U17251 (N_17251,N_16873,N_16432);
nand U17252 (N_17252,N_16854,N_16662);
nor U17253 (N_17253,N_16522,N_16925);
and U17254 (N_17254,N_16012,N_16719);
nand U17255 (N_17255,N_16792,N_16248);
nor U17256 (N_17256,N_16318,N_16081);
xor U17257 (N_17257,N_16372,N_16903);
or U17258 (N_17258,N_16841,N_16809);
or U17259 (N_17259,N_16619,N_16068);
xnor U17260 (N_17260,N_16393,N_16001);
nand U17261 (N_17261,N_16040,N_16152);
nor U17262 (N_17262,N_16725,N_16400);
nand U17263 (N_17263,N_16535,N_16041);
and U17264 (N_17264,N_16696,N_16640);
and U17265 (N_17265,N_16647,N_16638);
and U17266 (N_17266,N_16092,N_16098);
nand U17267 (N_17267,N_16780,N_16449);
nor U17268 (N_17268,N_16789,N_16826);
or U17269 (N_17269,N_16525,N_16231);
nand U17270 (N_17270,N_16453,N_16833);
and U17271 (N_17271,N_16995,N_16765);
or U17272 (N_17272,N_16960,N_16405);
nor U17273 (N_17273,N_16736,N_16935);
nand U17274 (N_17274,N_16975,N_16793);
nand U17275 (N_17275,N_16663,N_16920);
or U17276 (N_17276,N_16395,N_16392);
nand U17277 (N_17277,N_16757,N_16094);
nor U17278 (N_17278,N_16751,N_16429);
xnor U17279 (N_17279,N_16979,N_16771);
nand U17280 (N_17280,N_16927,N_16024);
nand U17281 (N_17281,N_16408,N_16455);
or U17282 (N_17282,N_16471,N_16180);
and U17283 (N_17283,N_16546,N_16328);
nand U17284 (N_17284,N_16125,N_16685);
nor U17285 (N_17285,N_16154,N_16223);
nor U17286 (N_17286,N_16258,N_16718);
or U17287 (N_17287,N_16591,N_16519);
nor U17288 (N_17288,N_16532,N_16606);
or U17289 (N_17289,N_16168,N_16529);
nor U17290 (N_17290,N_16123,N_16100);
xnor U17291 (N_17291,N_16426,N_16786);
nand U17292 (N_17292,N_16675,N_16758);
or U17293 (N_17293,N_16714,N_16366);
nand U17294 (N_17294,N_16828,N_16767);
nor U17295 (N_17295,N_16476,N_16071);
nor U17296 (N_17296,N_16646,N_16281);
xnor U17297 (N_17297,N_16959,N_16652);
and U17298 (N_17298,N_16796,N_16023);
or U17299 (N_17299,N_16160,N_16444);
nand U17300 (N_17300,N_16777,N_16989);
nor U17301 (N_17301,N_16491,N_16296);
and U17302 (N_17302,N_16019,N_16084);
or U17303 (N_17303,N_16194,N_16990);
or U17304 (N_17304,N_16327,N_16872);
and U17305 (N_17305,N_16085,N_16911);
nand U17306 (N_17306,N_16614,N_16550);
or U17307 (N_17307,N_16457,N_16016);
nor U17308 (N_17308,N_16868,N_16598);
nor U17309 (N_17309,N_16997,N_16197);
and U17310 (N_17310,N_16785,N_16381);
nand U17311 (N_17311,N_16298,N_16342);
and U17312 (N_17312,N_16958,N_16107);
nor U17313 (N_17313,N_16313,N_16131);
xor U17314 (N_17314,N_16031,N_16806);
xor U17315 (N_17315,N_16176,N_16436);
and U17316 (N_17316,N_16923,N_16881);
nor U17317 (N_17317,N_16273,N_16501);
nor U17318 (N_17318,N_16420,N_16486);
or U17319 (N_17319,N_16570,N_16945);
nand U17320 (N_17320,N_16069,N_16937);
nor U17321 (N_17321,N_16812,N_16716);
xnor U17322 (N_17322,N_16608,N_16170);
or U17323 (N_17323,N_16130,N_16319);
and U17324 (N_17324,N_16564,N_16133);
nor U17325 (N_17325,N_16013,N_16728);
and U17326 (N_17326,N_16412,N_16138);
nor U17327 (N_17327,N_16613,N_16241);
or U17328 (N_17328,N_16267,N_16418);
xor U17329 (N_17329,N_16908,N_16058);
or U17330 (N_17330,N_16363,N_16681);
nand U17331 (N_17331,N_16499,N_16032);
nand U17332 (N_17332,N_16127,N_16110);
and U17333 (N_17333,N_16666,N_16688);
or U17334 (N_17334,N_16516,N_16810);
xor U17335 (N_17335,N_16158,N_16222);
nor U17336 (N_17336,N_16912,N_16280);
nor U17337 (N_17337,N_16738,N_16075);
nand U17338 (N_17338,N_16750,N_16440);
or U17339 (N_17339,N_16136,N_16850);
or U17340 (N_17340,N_16858,N_16175);
xor U17341 (N_17341,N_16332,N_16205);
nor U17342 (N_17342,N_16232,N_16080);
xnor U17343 (N_17343,N_16243,N_16705);
and U17344 (N_17344,N_16956,N_16359);
nand U17345 (N_17345,N_16349,N_16506);
or U17346 (N_17346,N_16830,N_16885);
and U17347 (N_17347,N_16551,N_16184);
xnor U17348 (N_17348,N_16386,N_16121);
nand U17349 (N_17349,N_16585,N_16849);
or U17350 (N_17350,N_16434,N_16082);
or U17351 (N_17351,N_16141,N_16710);
nor U17352 (N_17352,N_16143,N_16300);
xnor U17353 (N_17353,N_16899,N_16527);
and U17354 (N_17354,N_16645,N_16039);
or U17355 (N_17355,N_16086,N_16473);
nor U17356 (N_17356,N_16691,N_16213);
or U17357 (N_17357,N_16398,N_16930);
nor U17358 (N_17358,N_16150,N_16224);
and U17359 (N_17359,N_16034,N_16766);
xnor U17360 (N_17360,N_16616,N_16004);
or U17361 (N_17361,N_16726,N_16648);
and U17362 (N_17362,N_16871,N_16621);
nor U17363 (N_17363,N_16256,N_16009);
nor U17364 (N_17364,N_16706,N_16140);
or U17365 (N_17365,N_16479,N_16552);
and U17366 (N_17366,N_16769,N_16572);
and U17367 (N_17367,N_16448,N_16352);
or U17368 (N_17368,N_16891,N_16601);
nor U17369 (N_17369,N_16401,N_16589);
xnor U17370 (N_17370,N_16209,N_16238);
or U17371 (N_17371,N_16615,N_16106);
and U17372 (N_17372,N_16731,N_16604);
and U17373 (N_17373,N_16482,N_16922);
nand U17374 (N_17374,N_16251,N_16947);
or U17375 (N_17375,N_16384,N_16940);
and U17376 (N_17376,N_16539,N_16971);
nor U17377 (N_17377,N_16056,N_16196);
nand U17378 (N_17378,N_16932,N_16421);
xor U17379 (N_17379,N_16102,N_16331);
and U17380 (N_17380,N_16011,N_16583);
and U17381 (N_17381,N_16976,N_16851);
nor U17382 (N_17382,N_16186,N_16151);
nand U17383 (N_17383,N_16847,N_16166);
nand U17384 (N_17384,N_16355,N_16837);
nand U17385 (N_17385,N_16748,N_16949);
nand U17386 (N_17386,N_16875,N_16022);
nand U17387 (N_17387,N_16093,N_16561);
or U17388 (N_17388,N_16484,N_16708);
and U17389 (N_17389,N_16542,N_16262);
nor U17390 (N_17390,N_16315,N_16091);
or U17391 (N_17391,N_16035,N_16687);
or U17392 (N_17392,N_16246,N_16410);
and U17393 (N_17393,N_16112,N_16185);
nand U17394 (N_17394,N_16061,N_16713);
nand U17395 (N_17395,N_16817,N_16905);
xor U17396 (N_17396,N_16676,N_16581);
or U17397 (N_17397,N_16403,N_16650);
nor U17398 (N_17398,N_16337,N_16220);
and U17399 (N_17399,N_16859,N_16861);
nand U17400 (N_17400,N_16037,N_16882);
nor U17401 (N_17401,N_16199,N_16695);
or U17402 (N_17402,N_16304,N_16126);
nand U17403 (N_17403,N_16749,N_16744);
nor U17404 (N_17404,N_16369,N_16963);
or U17405 (N_17405,N_16033,N_16579);
and U17406 (N_17406,N_16709,N_16704);
nor U17407 (N_17407,N_16500,N_16926);
nor U17408 (N_17408,N_16798,N_16674);
and U17409 (N_17409,N_16807,N_16073);
nand U17410 (N_17410,N_16182,N_16890);
and U17411 (N_17411,N_16210,N_16637);
nor U17412 (N_17412,N_16672,N_16693);
or U17413 (N_17413,N_16417,N_16739);
xor U17414 (N_17414,N_16469,N_16206);
xnor U17415 (N_17415,N_16129,N_16162);
or U17416 (N_17416,N_16634,N_16054);
nand U17417 (N_17417,N_16624,N_16654);
nand U17418 (N_17418,N_16988,N_16254);
nor U17419 (N_17419,N_16438,N_16306);
or U17420 (N_17420,N_16066,N_16998);
or U17421 (N_17421,N_16623,N_16227);
or U17422 (N_17422,N_16743,N_16450);
nor U17423 (N_17423,N_16510,N_16964);
nand U17424 (N_17424,N_16505,N_16334);
and U17425 (N_17425,N_16495,N_16756);
nor U17426 (N_17426,N_16504,N_16096);
nor U17427 (N_17427,N_16063,N_16470);
xnor U17428 (N_17428,N_16978,N_16324);
and U17429 (N_17429,N_16782,N_16320);
nor U17430 (N_17430,N_16167,N_16783);
nand U17431 (N_17431,N_16842,N_16302);
nand U17432 (N_17432,N_16026,N_16252);
or U17433 (N_17433,N_16944,N_16664);
and U17434 (N_17434,N_16818,N_16775);
and U17435 (N_17435,N_16326,N_16480);
or U17436 (N_17436,N_16481,N_16869);
and U17437 (N_17437,N_16628,N_16070);
or U17438 (N_17438,N_16595,N_16297);
and U17439 (N_17439,N_16338,N_16046);
and U17440 (N_17440,N_16214,N_16048);
nand U17441 (N_17441,N_16285,N_16260);
nand U17442 (N_17442,N_16493,N_16365);
or U17443 (N_17443,N_16768,N_16321);
or U17444 (N_17444,N_16866,N_16745);
nor U17445 (N_17445,N_16079,N_16376);
nor U17446 (N_17446,N_16464,N_16284);
or U17447 (N_17447,N_16490,N_16002);
or U17448 (N_17448,N_16264,N_16379);
nand U17449 (N_17449,N_16088,N_16090);
nor U17450 (N_17450,N_16000,N_16955);
and U17451 (N_17451,N_16555,N_16586);
xor U17452 (N_17452,N_16462,N_16275);
xor U17453 (N_17453,N_16111,N_16507);
or U17454 (N_17454,N_16119,N_16576);
nor U17455 (N_17455,N_16799,N_16917);
nand U17456 (N_17456,N_16397,N_16391);
nor U17457 (N_17457,N_16867,N_16291);
and U17458 (N_17458,N_16986,N_16322);
or U17459 (N_17459,N_16965,N_16894);
nand U17460 (N_17460,N_16378,N_16701);
and U17461 (N_17461,N_16414,N_16055);
or U17462 (N_17462,N_16445,N_16430);
nor U17463 (N_17463,N_16590,N_16225);
nand U17464 (N_17464,N_16864,N_16375);
nor U17465 (N_17465,N_16609,N_16203);
and U17466 (N_17466,N_16898,N_16461);
or U17467 (N_17467,N_16018,N_16014);
and U17468 (N_17468,N_16219,N_16108);
and U17469 (N_17469,N_16077,N_16411);
nand U17470 (N_17470,N_16723,N_16951);
xor U17471 (N_17471,N_16124,N_16271);
xnor U17472 (N_17472,N_16730,N_16603);
or U17473 (N_17473,N_16439,N_16928);
xnor U17474 (N_17474,N_16834,N_16835);
nor U17475 (N_17475,N_16985,N_16431);
or U17476 (N_17476,N_16274,N_16566);
or U17477 (N_17477,N_16494,N_16373);
or U17478 (N_17478,N_16560,N_16980);
nor U17479 (N_17479,N_16563,N_16588);
nand U17480 (N_17480,N_16358,N_16592);
nor U17481 (N_17481,N_16853,N_16178);
nor U17482 (N_17482,N_16852,N_16656);
xor U17483 (N_17483,N_16722,N_16987);
or U17484 (N_17484,N_16308,N_16467);
nor U17485 (N_17485,N_16548,N_16526);
nand U17486 (N_17486,N_16877,N_16290);
xor U17487 (N_17487,N_16283,N_16394);
or U17488 (N_17488,N_16478,N_16653);
or U17489 (N_17489,N_16446,N_16962);
nand U17490 (N_17490,N_16543,N_16689);
nor U17491 (N_17491,N_16597,N_16746);
and U17492 (N_17492,N_16406,N_16682);
nor U17493 (N_17493,N_16474,N_16269);
and U17494 (N_17494,N_16488,N_16540);
or U17495 (N_17495,N_16660,N_16630);
and U17496 (N_17496,N_16122,N_16095);
and U17497 (N_17497,N_16288,N_16027);
nand U17498 (N_17498,N_16605,N_16314);
and U17499 (N_17499,N_16261,N_16044);
or U17500 (N_17500,N_16884,N_16095);
nor U17501 (N_17501,N_16274,N_16547);
or U17502 (N_17502,N_16861,N_16076);
xnor U17503 (N_17503,N_16180,N_16702);
xor U17504 (N_17504,N_16849,N_16099);
nand U17505 (N_17505,N_16220,N_16463);
nor U17506 (N_17506,N_16437,N_16501);
nand U17507 (N_17507,N_16828,N_16444);
xnor U17508 (N_17508,N_16932,N_16663);
nand U17509 (N_17509,N_16360,N_16571);
and U17510 (N_17510,N_16453,N_16591);
nor U17511 (N_17511,N_16616,N_16332);
and U17512 (N_17512,N_16527,N_16673);
or U17513 (N_17513,N_16585,N_16506);
and U17514 (N_17514,N_16709,N_16163);
or U17515 (N_17515,N_16288,N_16539);
or U17516 (N_17516,N_16063,N_16223);
and U17517 (N_17517,N_16860,N_16621);
and U17518 (N_17518,N_16010,N_16151);
nor U17519 (N_17519,N_16771,N_16046);
xor U17520 (N_17520,N_16459,N_16077);
and U17521 (N_17521,N_16700,N_16984);
xor U17522 (N_17522,N_16567,N_16245);
and U17523 (N_17523,N_16956,N_16589);
nand U17524 (N_17524,N_16155,N_16182);
nor U17525 (N_17525,N_16732,N_16974);
nor U17526 (N_17526,N_16781,N_16630);
nor U17527 (N_17527,N_16598,N_16439);
nor U17528 (N_17528,N_16268,N_16391);
nor U17529 (N_17529,N_16245,N_16628);
nor U17530 (N_17530,N_16213,N_16684);
xor U17531 (N_17531,N_16413,N_16410);
and U17532 (N_17532,N_16976,N_16609);
and U17533 (N_17533,N_16572,N_16526);
and U17534 (N_17534,N_16514,N_16529);
or U17535 (N_17535,N_16346,N_16876);
nand U17536 (N_17536,N_16778,N_16211);
nand U17537 (N_17537,N_16816,N_16148);
nor U17538 (N_17538,N_16956,N_16662);
xor U17539 (N_17539,N_16352,N_16888);
xor U17540 (N_17540,N_16524,N_16937);
or U17541 (N_17541,N_16146,N_16367);
nor U17542 (N_17542,N_16486,N_16246);
and U17543 (N_17543,N_16726,N_16192);
nor U17544 (N_17544,N_16613,N_16412);
xor U17545 (N_17545,N_16033,N_16211);
or U17546 (N_17546,N_16383,N_16767);
xor U17547 (N_17547,N_16905,N_16532);
nand U17548 (N_17548,N_16210,N_16276);
and U17549 (N_17549,N_16046,N_16375);
nor U17550 (N_17550,N_16559,N_16973);
xor U17551 (N_17551,N_16232,N_16683);
nor U17552 (N_17552,N_16748,N_16532);
xor U17553 (N_17553,N_16257,N_16234);
nand U17554 (N_17554,N_16701,N_16636);
or U17555 (N_17555,N_16473,N_16116);
nand U17556 (N_17556,N_16410,N_16788);
nor U17557 (N_17557,N_16300,N_16169);
nor U17558 (N_17558,N_16802,N_16379);
or U17559 (N_17559,N_16893,N_16599);
and U17560 (N_17560,N_16855,N_16909);
or U17561 (N_17561,N_16437,N_16993);
nor U17562 (N_17562,N_16048,N_16805);
nand U17563 (N_17563,N_16573,N_16574);
and U17564 (N_17564,N_16434,N_16022);
and U17565 (N_17565,N_16543,N_16382);
nor U17566 (N_17566,N_16916,N_16179);
nand U17567 (N_17567,N_16695,N_16739);
or U17568 (N_17568,N_16807,N_16293);
or U17569 (N_17569,N_16723,N_16813);
nand U17570 (N_17570,N_16621,N_16603);
nand U17571 (N_17571,N_16280,N_16772);
and U17572 (N_17572,N_16387,N_16187);
xor U17573 (N_17573,N_16415,N_16734);
and U17574 (N_17574,N_16162,N_16614);
or U17575 (N_17575,N_16357,N_16613);
nand U17576 (N_17576,N_16427,N_16823);
xnor U17577 (N_17577,N_16898,N_16025);
and U17578 (N_17578,N_16874,N_16846);
nor U17579 (N_17579,N_16611,N_16714);
or U17580 (N_17580,N_16010,N_16978);
nand U17581 (N_17581,N_16269,N_16060);
nor U17582 (N_17582,N_16147,N_16335);
nand U17583 (N_17583,N_16959,N_16510);
nor U17584 (N_17584,N_16782,N_16406);
and U17585 (N_17585,N_16670,N_16265);
nor U17586 (N_17586,N_16191,N_16347);
or U17587 (N_17587,N_16968,N_16128);
nand U17588 (N_17588,N_16123,N_16994);
xor U17589 (N_17589,N_16091,N_16070);
nor U17590 (N_17590,N_16675,N_16973);
nor U17591 (N_17591,N_16807,N_16770);
nand U17592 (N_17592,N_16184,N_16236);
nor U17593 (N_17593,N_16963,N_16667);
and U17594 (N_17594,N_16482,N_16999);
nor U17595 (N_17595,N_16183,N_16350);
or U17596 (N_17596,N_16977,N_16119);
nand U17597 (N_17597,N_16816,N_16259);
nor U17598 (N_17598,N_16201,N_16391);
or U17599 (N_17599,N_16515,N_16044);
and U17600 (N_17600,N_16114,N_16017);
or U17601 (N_17601,N_16982,N_16901);
nor U17602 (N_17602,N_16040,N_16544);
nor U17603 (N_17603,N_16335,N_16378);
nand U17604 (N_17604,N_16513,N_16877);
or U17605 (N_17605,N_16943,N_16421);
nor U17606 (N_17606,N_16317,N_16041);
and U17607 (N_17607,N_16452,N_16003);
and U17608 (N_17608,N_16688,N_16238);
nor U17609 (N_17609,N_16491,N_16036);
nand U17610 (N_17610,N_16417,N_16661);
nor U17611 (N_17611,N_16228,N_16260);
nor U17612 (N_17612,N_16756,N_16046);
nor U17613 (N_17613,N_16005,N_16561);
and U17614 (N_17614,N_16397,N_16675);
or U17615 (N_17615,N_16645,N_16547);
xor U17616 (N_17616,N_16665,N_16701);
and U17617 (N_17617,N_16883,N_16613);
nand U17618 (N_17618,N_16264,N_16679);
and U17619 (N_17619,N_16556,N_16694);
or U17620 (N_17620,N_16168,N_16078);
nor U17621 (N_17621,N_16635,N_16672);
nor U17622 (N_17622,N_16450,N_16003);
nand U17623 (N_17623,N_16675,N_16866);
and U17624 (N_17624,N_16846,N_16351);
and U17625 (N_17625,N_16844,N_16044);
xnor U17626 (N_17626,N_16953,N_16429);
nor U17627 (N_17627,N_16182,N_16165);
xnor U17628 (N_17628,N_16076,N_16993);
or U17629 (N_17629,N_16846,N_16957);
xnor U17630 (N_17630,N_16869,N_16478);
nor U17631 (N_17631,N_16237,N_16655);
xor U17632 (N_17632,N_16871,N_16136);
nor U17633 (N_17633,N_16428,N_16630);
nand U17634 (N_17634,N_16528,N_16775);
nand U17635 (N_17635,N_16411,N_16003);
and U17636 (N_17636,N_16584,N_16429);
and U17637 (N_17637,N_16915,N_16723);
and U17638 (N_17638,N_16664,N_16238);
nor U17639 (N_17639,N_16334,N_16294);
nand U17640 (N_17640,N_16759,N_16420);
and U17641 (N_17641,N_16286,N_16848);
or U17642 (N_17642,N_16607,N_16964);
nand U17643 (N_17643,N_16313,N_16251);
nand U17644 (N_17644,N_16138,N_16661);
or U17645 (N_17645,N_16841,N_16911);
and U17646 (N_17646,N_16892,N_16377);
and U17647 (N_17647,N_16267,N_16695);
or U17648 (N_17648,N_16297,N_16278);
xor U17649 (N_17649,N_16437,N_16933);
nand U17650 (N_17650,N_16101,N_16104);
and U17651 (N_17651,N_16043,N_16245);
xnor U17652 (N_17652,N_16201,N_16470);
and U17653 (N_17653,N_16244,N_16009);
or U17654 (N_17654,N_16213,N_16173);
nand U17655 (N_17655,N_16671,N_16886);
and U17656 (N_17656,N_16579,N_16752);
or U17657 (N_17657,N_16360,N_16892);
and U17658 (N_17658,N_16556,N_16872);
or U17659 (N_17659,N_16513,N_16440);
xor U17660 (N_17660,N_16747,N_16153);
or U17661 (N_17661,N_16736,N_16247);
and U17662 (N_17662,N_16183,N_16514);
nor U17663 (N_17663,N_16541,N_16652);
nor U17664 (N_17664,N_16093,N_16148);
nor U17665 (N_17665,N_16259,N_16511);
and U17666 (N_17666,N_16222,N_16905);
and U17667 (N_17667,N_16366,N_16676);
nor U17668 (N_17668,N_16718,N_16465);
and U17669 (N_17669,N_16730,N_16306);
nand U17670 (N_17670,N_16746,N_16067);
and U17671 (N_17671,N_16873,N_16583);
nand U17672 (N_17672,N_16248,N_16791);
and U17673 (N_17673,N_16150,N_16826);
or U17674 (N_17674,N_16430,N_16043);
and U17675 (N_17675,N_16130,N_16799);
nand U17676 (N_17676,N_16480,N_16969);
nor U17677 (N_17677,N_16669,N_16573);
and U17678 (N_17678,N_16266,N_16890);
or U17679 (N_17679,N_16417,N_16790);
and U17680 (N_17680,N_16455,N_16010);
nand U17681 (N_17681,N_16965,N_16378);
nor U17682 (N_17682,N_16000,N_16550);
or U17683 (N_17683,N_16327,N_16325);
nand U17684 (N_17684,N_16067,N_16456);
xor U17685 (N_17685,N_16807,N_16402);
or U17686 (N_17686,N_16731,N_16318);
or U17687 (N_17687,N_16496,N_16588);
nor U17688 (N_17688,N_16900,N_16316);
nor U17689 (N_17689,N_16127,N_16915);
or U17690 (N_17690,N_16201,N_16393);
nand U17691 (N_17691,N_16105,N_16946);
and U17692 (N_17692,N_16795,N_16976);
or U17693 (N_17693,N_16962,N_16626);
and U17694 (N_17694,N_16796,N_16083);
nor U17695 (N_17695,N_16373,N_16071);
xnor U17696 (N_17696,N_16024,N_16986);
xor U17697 (N_17697,N_16126,N_16547);
or U17698 (N_17698,N_16829,N_16811);
or U17699 (N_17699,N_16953,N_16472);
nand U17700 (N_17700,N_16302,N_16162);
nor U17701 (N_17701,N_16507,N_16993);
and U17702 (N_17702,N_16755,N_16943);
nand U17703 (N_17703,N_16764,N_16308);
xnor U17704 (N_17704,N_16652,N_16290);
nand U17705 (N_17705,N_16731,N_16704);
xnor U17706 (N_17706,N_16036,N_16562);
and U17707 (N_17707,N_16230,N_16746);
nor U17708 (N_17708,N_16978,N_16187);
or U17709 (N_17709,N_16133,N_16385);
or U17710 (N_17710,N_16624,N_16569);
or U17711 (N_17711,N_16531,N_16576);
nand U17712 (N_17712,N_16089,N_16043);
nor U17713 (N_17713,N_16851,N_16416);
and U17714 (N_17714,N_16031,N_16640);
xnor U17715 (N_17715,N_16362,N_16867);
xor U17716 (N_17716,N_16324,N_16972);
or U17717 (N_17717,N_16519,N_16257);
or U17718 (N_17718,N_16069,N_16931);
nand U17719 (N_17719,N_16437,N_16256);
xnor U17720 (N_17720,N_16032,N_16570);
nor U17721 (N_17721,N_16320,N_16917);
and U17722 (N_17722,N_16118,N_16561);
nand U17723 (N_17723,N_16584,N_16032);
or U17724 (N_17724,N_16143,N_16142);
nor U17725 (N_17725,N_16348,N_16480);
nand U17726 (N_17726,N_16723,N_16029);
nor U17727 (N_17727,N_16679,N_16266);
nand U17728 (N_17728,N_16644,N_16600);
or U17729 (N_17729,N_16812,N_16535);
and U17730 (N_17730,N_16711,N_16286);
or U17731 (N_17731,N_16136,N_16602);
nor U17732 (N_17732,N_16256,N_16616);
or U17733 (N_17733,N_16662,N_16201);
nor U17734 (N_17734,N_16042,N_16864);
and U17735 (N_17735,N_16955,N_16938);
nand U17736 (N_17736,N_16674,N_16877);
nor U17737 (N_17737,N_16299,N_16037);
nand U17738 (N_17738,N_16908,N_16059);
nor U17739 (N_17739,N_16301,N_16747);
xnor U17740 (N_17740,N_16732,N_16513);
or U17741 (N_17741,N_16014,N_16720);
and U17742 (N_17742,N_16233,N_16451);
nor U17743 (N_17743,N_16524,N_16200);
nand U17744 (N_17744,N_16262,N_16779);
and U17745 (N_17745,N_16842,N_16743);
nand U17746 (N_17746,N_16443,N_16021);
nand U17747 (N_17747,N_16226,N_16112);
nand U17748 (N_17748,N_16583,N_16892);
or U17749 (N_17749,N_16630,N_16585);
xor U17750 (N_17750,N_16284,N_16828);
and U17751 (N_17751,N_16421,N_16065);
and U17752 (N_17752,N_16639,N_16630);
or U17753 (N_17753,N_16499,N_16022);
or U17754 (N_17754,N_16516,N_16914);
nor U17755 (N_17755,N_16822,N_16479);
and U17756 (N_17756,N_16194,N_16602);
and U17757 (N_17757,N_16838,N_16538);
nor U17758 (N_17758,N_16992,N_16386);
and U17759 (N_17759,N_16187,N_16382);
nand U17760 (N_17760,N_16078,N_16852);
xor U17761 (N_17761,N_16563,N_16672);
xor U17762 (N_17762,N_16651,N_16203);
or U17763 (N_17763,N_16742,N_16335);
xor U17764 (N_17764,N_16634,N_16891);
nand U17765 (N_17765,N_16973,N_16552);
nor U17766 (N_17766,N_16985,N_16835);
nor U17767 (N_17767,N_16515,N_16274);
and U17768 (N_17768,N_16152,N_16710);
nand U17769 (N_17769,N_16621,N_16458);
or U17770 (N_17770,N_16369,N_16198);
xnor U17771 (N_17771,N_16711,N_16833);
or U17772 (N_17772,N_16507,N_16694);
nand U17773 (N_17773,N_16387,N_16808);
nand U17774 (N_17774,N_16648,N_16090);
xnor U17775 (N_17775,N_16022,N_16435);
and U17776 (N_17776,N_16911,N_16149);
or U17777 (N_17777,N_16002,N_16771);
nor U17778 (N_17778,N_16317,N_16642);
or U17779 (N_17779,N_16631,N_16380);
and U17780 (N_17780,N_16786,N_16571);
nor U17781 (N_17781,N_16281,N_16198);
xnor U17782 (N_17782,N_16757,N_16557);
or U17783 (N_17783,N_16450,N_16052);
and U17784 (N_17784,N_16083,N_16999);
and U17785 (N_17785,N_16073,N_16591);
nand U17786 (N_17786,N_16982,N_16400);
and U17787 (N_17787,N_16222,N_16575);
xnor U17788 (N_17788,N_16219,N_16198);
nor U17789 (N_17789,N_16421,N_16860);
and U17790 (N_17790,N_16083,N_16577);
and U17791 (N_17791,N_16627,N_16803);
nor U17792 (N_17792,N_16951,N_16806);
or U17793 (N_17793,N_16090,N_16688);
nand U17794 (N_17794,N_16131,N_16737);
nand U17795 (N_17795,N_16459,N_16505);
nor U17796 (N_17796,N_16562,N_16460);
and U17797 (N_17797,N_16564,N_16208);
xnor U17798 (N_17798,N_16300,N_16218);
and U17799 (N_17799,N_16325,N_16289);
nor U17800 (N_17800,N_16123,N_16727);
xor U17801 (N_17801,N_16015,N_16167);
nand U17802 (N_17802,N_16002,N_16215);
and U17803 (N_17803,N_16579,N_16206);
and U17804 (N_17804,N_16505,N_16913);
and U17805 (N_17805,N_16997,N_16064);
and U17806 (N_17806,N_16835,N_16384);
nand U17807 (N_17807,N_16881,N_16942);
and U17808 (N_17808,N_16338,N_16418);
nor U17809 (N_17809,N_16193,N_16662);
nand U17810 (N_17810,N_16818,N_16127);
nor U17811 (N_17811,N_16723,N_16080);
nor U17812 (N_17812,N_16426,N_16750);
xor U17813 (N_17813,N_16609,N_16168);
and U17814 (N_17814,N_16235,N_16225);
xnor U17815 (N_17815,N_16916,N_16324);
or U17816 (N_17816,N_16263,N_16914);
nor U17817 (N_17817,N_16434,N_16604);
nand U17818 (N_17818,N_16115,N_16464);
xor U17819 (N_17819,N_16198,N_16971);
xor U17820 (N_17820,N_16718,N_16515);
nor U17821 (N_17821,N_16295,N_16094);
or U17822 (N_17822,N_16327,N_16304);
nor U17823 (N_17823,N_16669,N_16465);
or U17824 (N_17824,N_16514,N_16485);
and U17825 (N_17825,N_16714,N_16042);
and U17826 (N_17826,N_16693,N_16626);
or U17827 (N_17827,N_16954,N_16318);
and U17828 (N_17828,N_16906,N_16477);
xnor U17829 (N_17829,N_16170,N_16642);
nor U17830 (N_17830,N_16778,N_16344);
and U17831 (N_17831,N_16436,N_16149);
or U17832 (N_17832,N_16410,N_16635);
or U17833 (N_17833,N_16291,N_16056);
nor U17834 (N_17834,N_16991,N_16609);
or U17835 (N_17835,N_16065,N_16353);
and U17836 (N_17836,N_16333,N_16080);
and U17837 (N_17837,N_16280,N_16703);
or U17838 (N_17838,N_16409,N_16586);
nand U17839 (N_17839,N_16633,N_16227);
and U17840 (N_17840,N_16777,N_16818);
and U17841 (N_17841,N_16518,N_16188);
nand U17842 (N_17842,N_16529,N_16437);
nand U17843 (N_17843,N_16655,N_16130);
xor U17844 (N_17844,N_16813,N_16383);
nand U17845 (N_17845,N_16295,N_16027);
and U17846 (N_17846,N_16090,N_16493);
and U17847 (N_17847,N_16797,N_16951);
nand U17848 (N_17848,N_16973,N_16173);
or U17849 (N_17849,N_16516,N_16983);
and U17850 (N_17850,N_16374,N_16571);
nor U17851 (N_17851,N_16074,N_16887);
xnor U17852 (N_17852,N_16381,N_16742);
nor U17853 (N_17853,N_16460,N_16656);
nand U17854 (N_17854,N_16317,N_16313);
and U17855 (N_17855,N_16563,N_16726);
or U17856 (N_17856,N_16255,N_16526);
xnor U17857 (N_17857,N_16346,N_16423);
and U17858 (N_17858,N_16184,N_16180);
and U17859 (N_17859,N_16299,N_16920);
and U17860 (N_17860,N_16510,N_16659);
or U17861 (N_17861,N_16912,N_16861);
or U17862 (N_17862,N_16343,N_16072);
nor U17863 (N_17863,N_16782,N_16823);
nor U17864 (N_17864,N_16300,N_16639);
and U17865 (N_17865,N_16154,N_16855);
or U17866 (N_17866,N_16483,N_16361);
and U17867 (N_17867,N_16496,N_16927);
nor U17868 (N_17868,N_16038,N_16285);
nor U17869 (N_17869,N_16420,N_16343);
or U17870 (N_17870,N_16867,N_16315);
and U17871 (N_17871,N_16027,N_16325);
and U17872 (N_17872,N_16489,N_16727);
and U17873 (N_17873,N_16503,N_16256);
or U17874 (N_17874,N_16335,N_16240);
or U17875 (N_17875,N_16350,N_16357);
nor U17876 (N_17876,N_16744,N_16216);
nor U17877 (N_17877,N_16684,N_16191);
and U17878 (N_17878,N_16702,N_16125);
or U17879 (N_17879,N_16703,N_16015);
nand U17880 (N_17880,N_16102,N_16242);
and U17881 (N_17881,N_16096,N_16090);
nand U17882 (N_17882,N_16224,N_16222);
nor U17883 (N_17883,N_16350,N_16017);
nor U17884 (N_17884,N_16093,N_16625);
nor U17885 (N_17885,N_16884,N_16073);
or U17886 (N_17886,N_16231,N_16815);
and U17887 (N_17887,N_16261,N_16837);
nand U17888 (N_17888,N_16759,N_16044);
or U17889 (N_17889,N_16493,N_16228);
nor U17890 (N_17890,N_16375,N_16031);
nor U17891 (N_17891,N_16306,N_16701);
xnor U17892 (N_17892,N_16710,N_16712);
nand U17893 (N_17893,N_16696,N_16320);
and U17894 (N_17894,N_16813,N_16412);
nand U17895 (N_17895,N_16699,N_16447);
nor U17896 (N_17896,N_16603,N_16298);
and U17897 (N_17897,N_16894,N_16754);
or U17898 (N_17898,N_16542,N_16284);
and U17899 (N_17899,N_16736,N_16111);
nor U17900 (N_17900,N_16174,N_16935);
nand U17901 (N_17901,N_16995,N_16383);
nand U17902 (N_17902,N_16934,N_16145);
and U17903 (N_17903,N_16729,N_16751);
nand U17904 (N_17904,N_16586,N_16696);
xnor U17905 (N_17905,N_16954,N_16987);
nor U17906 (N_17906,N_16252,N_16597);
nor U17907 (N_17907,N_16106,N_16950);
nand U17908 (N_17908,N_16735,N_16822);
or U17909 (N_17909,N_16673,N_16660);
nor U17910 (N_17910,N_16587,N_16943);
xnor U17911 (N_17911,N_16413,N_16487);
and U17912 (N_17912,N_16495,N_16421);
or U17913 (N_17913,N_16588,N_16192);
nand U17914 (N_17914,N_16033,N_16397);
nor U17915 (N_17915,N_16193,N_16488);
and U17916 (N_17916,N_16144,N_16025);
nor U17917 (N_17917,N_16922,N_16874);
and U17918 (N_17918,N_16772,N_16433);
nand U17919 (N_17919,N_16440,N_16448);
or U17920 (N_17920,N_16975,N_16476);
nor U17921 (N_17921,N_16720,N_16136);
nor U17922 (N_17922,N_16166,N_16092);
nand U17923 (N_17923,N_16876,N_16734);
nor U17924 (N_17924,N_16561,N_16994);
nand U17925 (N_17925,N_16343,N_16898);
and U17926 (N_17926,N_16780,N_16671);
xor U17927 (N_17927,N_16495,N_16341);
nand U17928 (N_17928,N_16175,N_16890);
nor U17929 (N_17929,N_16656,N_16812);
and U17930 (N_17930,N_16041,N_16801);
nor U17931 (N_17931,N_16723,N_16933);
nand U17932 (N_17932,N_16126,N_16708);
nand U17933 (N_17933,N_16673,N_16147);
nand U17934 (N_17934,N_16207,N_16526);
xor U17935 (N_17935,N_16634,N_16429);
or U17936 (N_17936,N_16490,N_16537);
xor U17937 (N_17937,N_16419,N_16685);
and U17938 (N_17938,N_16343,N_16230);
nand U17939 (N_17939,N_16117,N_16812);
nand U17940 (N_17940,N_16320,N_16527);
or U17941 (N_17941,N_16521,N_16442);
and U17942 (N_17942,N_16636,N_16397);
nor U17943 (N_17943,N_16582,N_16842);
and U17944 (N_17944,N_16139,N_16979);
nor U17945 (N_17945,N_16738,N_16367);
nand U17946 (N_17946,N_16498,N_16448);
or U17947 (N_17947,N_16714,N_16098);
and U17948 (N_17948,N_16827,N_16021);
and U17949 (N_17949,N_16871,N_16276);
and U17950 (N_17950,N_16720,N_16866);
or U17951 (N_17951,N_16842,N_16696);
or U17952 (N_17952,N_16648,N_16276);
xor U17953 (N_17953,N_16000,N_16264);
and U17954 (N_17954,N_16790,N_16354);
nor U17955 (N_17955,N_16828,N_16432);
and U17956 (N_17956,N_16324,N_16425);
and U17957 (N_17957,N_16398,N_16140);
nand U17958 (N_17958,N_16164,N_16406);
and U17959 (N_17959,N_16895,N_16292);
or U17960 (N_17960,N_16348,N_16070);
nand U17961 (N_17961,N_16851,N_16799);
or U17962 (N_17962,N_16219,N_16805);
nor U17963 (N_17963,N_16891,N_16440);
xnor U17964 (N_17964,N_16236,N_16090);
or U17965 (N_17965,N_16400,N_16256);
nand U17966 (N_17966,N_16518,N_16077);
nand U17967 (N_17967,N_16071,N_16287);
or U17968 (N_17968,N_16924,N_16205);
and U17969 (N_17969,N_16594,N_16558);
and U17970 (N_17970,N_16576,N_16729);
and U17971 (N_17971,N_16034,N_16504);
nand U17972 (N_17972,N_16761,N_16017);
or U17973 (N_17973,N_16247,N_16123);
and U17974 (N_17974,N_16519,N_16338);
or U17975 (N_17975,N_16384,N_16444);
and U17976 (N_17976,N_16823,N_16737);
nand U17977 (N_17977,N_16487,N_16889);
nand U17978 (N_17978,N_16860,N_16643);
nand U17979 (N_17979,N_16562,N_16136);
nor U17980 (N_17980,N_16363,N_16365);
nor U17981 (N_17981,N_16315,N_16378);
nor U17982 (N_17982,N_16141,N_16441);
and U17983 (N_17983,N_16889,N_16642);
nand U17984 (N_17984,N_16387,N_16248);
or U17985 (N_17985,N_16716,N_16706);
and U17986 (N_17986,N_16902,N_16074);
and U17987 (N_17987,N_16119,N_16327);
nor U17988 (N_17988,N_16341,N_16193);
nor U17989 (N_17989,N_16583,N_16752);
or U17990 (N_17990,N_16581,N_16633);
nor U17991 (N_17991,N_16930,N_16595);
nor U17992 (N_17992,N_16253,N_16403);
xor U17993 (N_17993,N_16036,N_16938);
nand U17994 (N_17994,N_16809,N_16465);
and U17995 (N_17995,N_16265,N_16983);
xor U17996 (N_17996,N_16170,N_16965);
nor U17997 (N_17997,N_16926,N_16397);
nand U17998 (N_17998,N_16857,N_16272);
xor U17999 (N_17999,N_16911,N_16517);
nand U18000 (N_18000,N_17451,N_17139);
nor U18001 (N_18001,N_17741,N_17997);
and U18002 (N_18002,N_17745,N_17879);
and U18003 (N_18003,N_17898,N_17551);
xor U18004 (N_18004,N_17172,N_17821);
nor U18005 (N_18005,N_17310,N_17459);
nor U18006 (N_18006,N_17543,N_17570);
and U18007 (N_18007,N_17647,N_17592);
nor U18008 (N_18008,N_17642,N_17807);
nor U18009 (N_18009,N_17627,N_17864);
nor U18010 (N_18010,N_17010,N_17129);
xnor U18011 (N_18011,N_17230,N_17372);
nor U18012 (N_18012,N_17845,N_17078);
and U18013 (N_18013,N_17262,N_17524);
and U18014 (N_18014,N_17107,N_17303);
or U18015 (N_18015,N_17430,N_17605);
nand U18016 (N_18016,N_17818,N_17380);
nand U18017 (N_18017,N_17410,N_17335);
nand U18018 (N_18018,N_17921,N_17813);
nor U18019 (N_18019,N_17527,N_17508);
nand U18020 (N_18020,N_17757,N_17203);
nor U18021 (N_18021,N_17977,N_17175);
and U18022 (N_18022,N_17098,N_17406);
nor U18023 (N_18023,N_17790,N_17987);
nand U18024 (N_18024,N_17924,N_17952);
nand U18025 (N_18025,N_17258,N_17479);
or U18026 (N_18026,N_17374,N_17734);
and U18027 (N_18027,N_17160,N_17170);
and U18028 (N_18028,N_17296,N_17948);
nand U18029 (N_18029,N_17168,N_17827);
nand U18030 (N_18030,N_17616,N_17249);
nor U18031 (N_18031,N_17135,N_17243);
and U18032 (N_18032,N_17962,N_17283);
and U18033 (N_18033,N_17097,N_17018);
nand U18034 (N_18034,N_17448,N_17193);
or U18035 (N_18035,N_17884,N_17210);
xnor U18036 (N_18036,N_17201,N_17587);
and U18037 (N_18037,N_17783,N_17279);
or U18038 (N_18038,N_17370,N_17221);
xor U18039 (N_18039,N_17971,N_17390);
and U18040 (N_18040,N_17694,N_17309);
nand U18041 (N_18041,N_17225,N_17589);
nor U18042 (N_18042,N_17081,N_17763);
nand U18043 (N_18043,N_17331,N_17738);
and U18044 (N_18044,N_17939,N_17941);
nand U18045 (N_18045,N_17811,N_17732);
nand U18046 (N_18046,N_17231,N_17393);
and U18047 (N_18047,N_17874,N_17689);
nor U18048 (N_18048,N_17151,N_17253);
nand U18049 (N_18049,N_17252,N_17747);
xor U18050 (N_18050,N_17405,N_17163);
nand U18051 (N_18051,N_17892,N_17979);
nand U18052 (N_18052,N_17715,N_17241);
nand U18053 (N_18053,N_17314,N_17391);
nor U18054 (N_18054,N_17313,N_17700);
nand U18055 (N_18055,N_17463,N_17164);
nor U18056 (N_18056,N_17623,N_17523);
and U18057 (N_18057,N_17974,N_17565);
and U18058 (N_18058,N_17782,N_17349);
and U18059 (N_18059,N_17156,N_17533);
nand U18060 (N_18060,N_17057,N_17737);
or U18061 (N_18061,N_17348,N_17597);
and U18062 (N_18062,N_17909,N_17115);
and U18063 (N_18063,N_17556,N_17434);
nand U18064 (N_18064,N_17121,N_17145);
nand U18065 (N_18065,N_17658,N_17644);
xor U18066 (N_18066,N_17481,N_17529);
or U18067 (N_18067,N_17820,N_17970);
nand U18068 (N_18068,N_17166,N_17504);
nor U18069 (N_18069,N_17588,N_17542);
nand U18070 (N_18070,N_17000,N_17350);
and U18071 (N_18071,N_17831,N_17574);
xor U18072 (N_18072,N_17944,N_17246);
xor U18073 (N_18073,N_17891,N_17340);
or U18074 (N_18074,N_17361,N_17438);
or U18075 (N_18075,N_17618,N_17158);
and U18076 (N_18076,N_17263,N_17698);
and U18077 (N_18077,N_17213,N_17223);
nor U18078 (N_18078,N_17080,N_17612);
nor U18079 (N_18079,N_17104,N_17701);
or U18080 (N_18080,N_17334,N_17999);
or U18081 (N_18081,N_17815,N_17969);
or U18082 (N_18082,N_17007,N_17048);
and U18083 (N_18083,N_17111,N_17034);
or U18084 (N_18084,N_17282,N_17596);
or U18085 (N_18085,N_17559,N_17880);
or U18086 (N_18086,N_17105,N_17912);
or U18087 (N_18087,N_17431,N_17887);
nor U18088 (N_18088,N_17278,N_17413);
or U18089 (N_18089,N_17134,N_17379);
nor U18090 (N_18090,N_17452,N_17710);
nand U18091 (N_18091,N_17803,N_17106);
xnor U18092 (N_18092,N_17245,N_17595);
and U18093 (N_18093,N_17507,N_17005);
nor U18094 (N_18094,N_17625,N_17454);
nor U18095 (N_18095,N_17639,N_17049);
and U18096 (N_18096,N_17847,N_17522);
or U18097 (N_18097,N_17840,N_17960);
nand U18098 (N_18098,N_17159,N_17495);
nand U18099 (N_18099,N_17538,N_17001);
nand U18100 (N_18100,N_17916,N_17301);
nor U18101 (N_18101,N_17731,N_17345);
xor U18102 (N_18102,N_17101,N_17086);
or U18103 (N_18103,N_17179,N_17656);
nand U18104 (N_18104,N_17752,N_17494);
and U18105 (N_18105,N_17687,N_17852);
nor U18106 (N_18106,N_17011,N_17472);
and U18107 (N_18107,N_17548,N_17118);
nand U18108 (N_18108,N_17009,N_17268);
or U18109 (N_18109,N_17267,N_17855);
and U18110 (N_18110,N_17674,N_17445);
nand U18111 (N_18111,N_17711,N_17006);
nand U18112 (N_18112,N_17265,N_17103);
nand U18113 (N_18113,N_17401,N_17186);
nor U18114 (N_18114,N_17753,N_17774);
or U18115 (N_18115,N_17281,N_17904);
and U18116 (N_18116,N_17358,N_17581);
or U18117 (N_18117,N_17931,N_17383);
and U18118 (N_18118,N_17728,N_17469);
nand U18119 (N_18119,N_17675,N_17893);
and U18120 (N_18120,N_17403,N_17560);
or U18121 (N_18121,N_17141,N_17387);
or U18122 (N_18122,N_17718,N_17980);
nand U18123 (N_18123,N_17399,N_17363);
and U18124 (N_18124,N_17446,N_17464);
or U18125 (N_18125,N_17211,N_17462);
nand U18126 (N_18126,N_17315,N_17482);
nor U18127 (N_18127,N_17515,N_17549);
and U18128 (N_18128,N_17228,N_17222);
or U18129 (N_18129,N_17032,N_17835);
nor U18130 (N_18130,N_17247,N_17502);
nand U18131 (N_18131,N_17044,N_17470);
and U18132 (N_18132,N_17720,N_17829);
or U18133 (N_18133,N_17302,N_17087);
xor U18134 (N_18134,N_17802,N_17951);
nor U18135 (N_18135,N_17306,N_17501);
xor U18136 (N_18136,N_17863,N_17419);
nor U18137 (N_18137,N_17217,N_17337);
nor U18138 (N_18138,N_17229,N_17045);
and U18139 (N_18139,N_17365,N_17503);
nor U18140 (N_18140,N_17376,N_17695);
nor U18141 (N_18141,N_17795,N_17090);
nor U18142 (N_18142,N_17037,N_17900);
nand U18143 (N_18143,N_17284,N_17322);
and U18144 (N_18144,N_17113,N_17534);
and U18145 (N_18145,N_17610,N_17359);
xor U18146 (N_18146,N_17773,N_17713);
or U18147 (N_18147,N_17063,N_17418);
nand U18148 (N_18148,N_17318,N_17295);
or U18149 (N_18149,N_17841,N_17513);
or U18150 (N_18150,N_17577,N_17993);
nand U18151 (N_18151,N_17860,N_17338);
or U18152 (N_18152,N_17137,N_17120);
or U18153 (N_18153,N_17266,N_17788);
nor U18154 (N_18154,N_17708,N_17071);
nand U18155 (N_18155,N_17759,N_17865);
nor U18156 (N_18156,N_17292,N_17084);
nand U18157 (N_18157,N_17456,N_17927);
or U18158 (N_18158,N_17466,N_17958);
and U18159 (N_18159,N_17339,N_17509);
nand U18160 (N_18160,N_17846,N_17122);
and U18161 (N_18161,N_17308,N_17885);
and U18162 (N_18162,N_17575,N_17794);
nor U18163 (N_18163,N_17594,N_17636);
nor U18164 (N_18164,N_17780,N_17729);
and U18165 (N_18165,N_17136,N_17461);
or U18166 (N_18166,N_17959,N_17259);
and U18167 (N_18167,N_17169,N_17116);
nor U18168 (N_18168,N_17050,N_17521);
nor U18169 (N_18169,N_17812,N_17260);
xnor U18170 (N_18170,N_17490,N_17157);
nand U18171 (N_18171,N_17027,N_17740);
or U18172 (N_18172,N_17785,N_17473);
nand U18173 (N_18173,N_17460,N_17917);
and U18174 (N_18174,N_17199,N_17765);
and U18175 (N_18175,N_17366,N_17545);
xnor U18176 (N_18176,N_17664,N_17070);
nand U18177 (N_18177,N_17415,N_17660);
or U18178 (N_18178,N_17060,N_17746);
or U18179 (N_18179,N_17065,N_17777);
or U18180 (N_18180,N_17304,N_17019);
nand U18181 (N_18181,N_17953,N_17657);
nand U18182 (N_18182,N_17510,N_17843);
or U18183 (N_18183,N_17930,N_17998);
and U18184 (N_18184,N_17603,N_17882);
and U18185 (N_18185,N_17442,N_17068);
nor U18186 (N_18186,N_17233,N_17447);
nand U18187 (N_18187,N_17127,N_17877);
or U18188 (N_18188,N_17300,N_17085);
nand U18189 (N_18189,N_17663,N_17385);
nand U18190 (N_18190,N_17427,N_17102);
and U18191 (N_18191,N_17723,N_17305);
nand U18192 (N_18192,N_17554,N_17218);
or U18193 (N_18193,N_17798,N_17076);
and U18194 (N_18194,N_17580,N_17978);
nand U18195 (N_18195,N_17149,N_17192);
and U18196 (N_18196,N_17784,N_17176);
and U18197 (N_18197,N_17051,N_17069);
and U18198 (N_18198,N_17957,N_17561);
or U18199 (N_18199,N_17458,N_17789);
xnor U18200 (N_18200,N_17576,N_17681);
or U18201 (N_18201,N_17117,N_17205);
nor U18202 (N_18202,N_17095,N_17319);
nor U18203 (N_18203,N_17209,N_17404);
or U18204 (N_18204,N_17735,N_17058);
and U18205 (N_18205,N_17493,N_17398);
or U18206 (N_18206,N_17352,N_17329);
and U18207 (N_18207,N_17333,N_17547);
nand U18208 (N_18208,N_17356,N_17035);
or U18209 (N_18209,N_17641,N_17760);
nand U18210 (N_18210,N_17025,N_17796);
and U18211 (N_18211,N_17683,N_17629);
or U18212 (N_18212,N_17566,N_17407);
or U18213 (N_18213,N_17686,N_17029);
and U18214 (N_18214,N_17806,N_17722);
and U18215 (N_18215,N_17726,N_17367);
or U18216 (N_18216,N_17219,N_17600);
or U18217 (N_18217,N_17272,N_17441);
and U18218 (N_18218,N_17299,N_17234);
xor U18219 (N_18219,N_17326,N_17584);
nand U18220 (N_18220,N_17804,N_17008);
and U18221 (N_18221,N_17054,N_17637);
xor U18222 (N_18222,N_17981,N_17130);
nand U18223 (N_18223,N_17119,N_17950);
or U18224 (N_18224,N_17604,N_17653);
xor U18225 (N_18225,N_17922,N_17808);
nand U18226 (N_18226,N_17291,N_17388);
and U18227 (N_18227,N_17633,N_17215);
nand U18228 (N_18228,N_17643,N_17270);
and U18229 (N_18229,N_17832,N_17138);
nand U18230 (N_18230,N_17975,N_17615);
or U18231 (N_18231,N_17769,N_17934);
xor U18232 (N_18232,N_17856,N_17435);
or U18233 (N_18233,N_17862,N_17440);
and U18234 (N_18234,N_17347,N_17679);
and U18235 (N_18235,N_17341,N_17437);
nor U18236 (N_18236,N_17992,N_17132);
and U18237 (N_18237,N_17449,N_17346);
and U18238 (N_18238,N_17355,N_17188);
nand U18239 (N_18239,N_17850,N_17572);
nor U18240 (N_18240,N_17825,N_17411);
nor U18241 (N_18241,N_17506,N_17582);
or U18242 (N_18242,N_17499,N_17800);
xnor U18243 (N_18243,N_17598,N_17894);
xnor U18244 (N_18244,N_17108,N_17364);
nand U18245 (N_18245,N_17162,N_17667);
and U18246 (N_18246,N_17770,N_17420);
nand U18247 (N_18247,N_17013,N_17567);
and U18248 (N_18248,N_17244,N_17640);
nor U18249 (N_18249,N_17954,N_17724);
nor U18250 (N_18250,N_17421,N_17038);
and U18251 (N_18251,N_17609,N_17943);
and U18252 (N_18252,N_17532,N_17896);
nor U18253 (N_18253,N_17526,N_17467);
or U18254 (N_18254,N_17328,N_17429);
xor U18255 (N_18255,N_17226,N_17949);
xnor U18256 (N_18256,N_17191,N_17381);
or U18257 (N_18257,N_17492,N_17607);
nand U18258 (N_18258,N_17457,N_17235);
or U18259 (N_18259,N_17839,N_17167);
or U18260 (N_18260,N_17918,N_17854);
nand U18261 (N_18261,N_17714,N_17743);
nand U18262 (N_18262,N_17028,N_17327);
or U18263 (N_18263,N_17195,N_17408);
nand U18264 (N_18264,N_17455,N_17703);
nand U18265 (N_18265,N_17725,N_17692);
or U18266 (N_18266,N_17336,N_17497);
or U18267 (N_18267,N_17059,N_17342);
xor U18268 (N_18268,N_17064,N_17183);
nand U18269 (N_18269,N_17212,N_17312);
nand U18270 (N_18270,N_17220,N_17091);
and U18271 (N_18271,N_17238,N_17094);
nor U18272 (N_18272,N_17500,N_17654);
or U18273 (N_18273,N_17083,N_17956);
nand U18274 (N_18274,N_17991,N_17748);
or U18275 (N_18275,N_17061,N_17465);
nand U18276 (N_18276,N_17040,N_17125);
xor U18277 (N_18277,N_17989,N_17739);
nand U18278 (N_18278,N_17932,N_17423);
nand U18279 (N_18279,N_17126,N_17810);
nor U18280 (N_18280,N_17453,N_17919);
and U18281 (N_18281,N_17669,N_17635);
or U18282 (N_18282,N_17144,N_17535);
or U18283 (N_18283,N_17432,N_17276);
or U18284 (N_18284,N_17148,N_17004);
and U18285 (N_18285,N_17907,N_17870);
and U18286 (N_18286,N_17428,N_17444);
nand U18287 (N_18287,N_17859,N_17571);
and U18288 (N_18288,N_17965,N_17539);
or U18289 (N_18289,N_17828,N_17389);
xor U18290 (N_18290,N_17072,N_17416);
nor U18291 (N_18291,N_17867,N_17801);
nand U18292 (N_18292,N_17142,N_17471);
and U18293 (N_18293,N_17673,N_17661);
and U18294 (N_18294,N_17593,N_17198);
nand U18295 (N_18295,N_17776,N_17848);
nor U18296 (N_18296,N_17995,N_17255);
nor U18297 (N_18297,N_17002,N_17324);
nor U18298 (N_18298,N_17540,N_17206);
xor U18299 (N_18299,N_17286,N_17298);
nor U18300 (N_18300,N_17964,N_17377);
nand U18301 (N_18301,N_17632,N_17585);
or U18302 (N_18302,N_17146,N_17173);
and U18303 (N_18303,N_17178,N_17323);
or U18304 (N_18304,N_17869,N_17171);
or U18305 (N_18305,N_17133,N_17696);
or U18306 (N_18306,N_17074,N_17277);
xnor U18307 (N_18307,N_17751,N_17307);
nand U18308 (N_18308,N_17152,N_17766);
nand U18309 (N_18309,N_17189,N_17638);
and U18310 (N_18310,N_17516,N_17395);
and U18311 (N_18311,N_17237,N_17412);
or U18312 (N_18312,N_17311,N_17787);
and U18313 (N_18313,N_17242,N_17705);
nor U18314 (N_18314,N_17131,N_17878);
xnor U18315 (N_18315,N_17020,N_17631);
nand U18316 (N_18316,N_17645,N_17207);
nor U18317 (N_18317,N_17239,N_17622);
nand U18318 (N_18318,N_17288,N_17426);
or U18319 (N_18319,N_17897,N_17023);
nor U18320 (N_18320,N_17414,N_17704);
nor U18321 (N_18321,N_17053,N_17823);
or U18322 (N_18322,N_17041,N_17396);
nor U18323 (N_18323,N_17180,N_17986);
and U18324 (N_18324,N_17177,N_17293);
xnor U18325 (N_18325,N_17520,N_17486);
nand U18326 (N_18326,N_17611,N_17990);
and U18327 (N_18327,N_17824,N_17409);
nor U18328 (N_18328,N_17519,N_17089);
nand U18329 (N_18329,N_17474,N_17662);
and U18330 (N_18330,N_17947,N_17764);
xor U18331 (N_18331,N_17982,N_17161);
nand U18332 (N_18332,N_17264,N_17208);
nand U18333 (N_18333,N_17214,N_17275);
or U18334 (N_18334,N_17988,N_17563);
or U18335 (N_18335,N_17143,N_17805);
and U18336 (N_18336,N_17826,N_17942);
nor U18337 (N_18337,N_17400,N_17558);
nor U18338 (N_18338,N_17923,N_17197);
nor U18339 (N_18339,N_17778,N_17256);
and U18340 (N_18340,N_17727,N_17392);
or U18341 (N_18341,N_17320,N_17749);
and U18342 (N_18342,N_17903,N_17280);
and U18343 (N_18343,N_17905,N_17926);
or U18344 (N_18344,N_17294,N_17354);
nand U18345 (N_18345,N_17634,N_17961);
xor U18346 (N_18346,N_17668,N_17216);
nor U18347 (N_18347,N_17996,N_17402);
or U18348 (N_18348,N_17343,N_17833);
nand U18349 (N_18349,N_17709,N_17837);
and U18350 (N_18350,N_17369,N_17688);
or U18351 (N_18351,N_17021,N_17140);
and U18352 (N_18352,N_17886,N_17517);
nand U18353 (N_18353,N_17099,N_17066);
nand U18354 (N_18354,N_17697,N_17344);
xnor U18355 (N_18355,N_17672,N_17531);
nor U18356 (N_18356,N_17250,N_17541);
nor U18357 (N_18357,N_17477,N_17047);
or U18358 (N_18358,N_17088,N_17489);
and U18359 (N_18359,N_17933,N_17883);
or U18360 (N_18360,N_17614,N_17583);
nor U18361 (N_18361,N_17913,N_17792);
or U18362 (N_18362,N_17822,N_17190);
nand U18363 (N_18363,N_17676,N_17297);
or U18364 (N_18364,N_17578,N_17666);
and U18365 (N_18365,N_17251,N_17911);
and U18366 (N_18366,N_17797,N_17012);
nand U18367 (N_18367,N_17791,N_17976);
and U18368 (N_18368,N_17450,N_17851);
and U18369 (N_18369,N_17124,N_17966);
or U18370 (N_18370,N_17649,N_17373);
or U18371 (N_18371,N_17677,N_17648);
and U18372 (N_18372,N_17849,N_17736);
xor U18373 (N_18373,N_17039,N_17202);
nand U18374 (N_18374,N_17601,N_17325);
or U18375 (N_18375,N_17733,N_17382);
nor U18376 (N_18376,N_17973,N_17204);
xor U18377 (N_18377,N_17651,N_17353);
and U18378 (N_18378,N_17036,N_17834);
nor U18379 (N_18379,N_17368,N_17552);
or U18380 (N_18380,N_17371,N_17684);
or U18381 (N_18381,N_17174,N_17602);
nor U18382 (N_18382,N_17685,N_17553);
xnor U18383 (N_18383,N_17015,N_17853);
or U18384 (N_18384,N_17109,N_17397);
xor U18385 (N_18385,N_17809,N_17599);
nand U18386 (N_18386,N_17817,N_17755);
or U18387 (N_18387,N_17902,N_17985);
or U18388 (N_18388,N_17123,N_17055);
or U18389 (N_18389,N_17868,N_17562);
nor U18390 (N_18390,N_17691,N_17196);
or U18391 (N_18391,N_17768,N_17569);
nor U18392 (N_18392,N_17154,N_17274);
nor U18393 (N_18393,N_17092,N_17200);
and U18394 (N_18394,N_17875,N_17935);
and U18395 (N_18395,N_17014,N_17240);
and U18396 (N_18396,N_17257,N_17536);
xor U18397 (N_18397,N_17968,N_17033);
nand U18398 (N_18398,N_17754,N_17920);
or U18399 (N_18399,N_17290,N_17484);
nand U18400 (N_18400,N_17659,N_17937);
nand U18401 (N_18401,N_17756,N_17042);
and U18402 (N_18402,N_17617,N_17518);
and U18403 (N_18403,N_17699,N_17384);
nand U18404 (N_18404,N_17682,N_17591);
nand U18405 (N_18405,N_17967,N_17557);
nor U18406 (N_18406,N_17248,N_17719);
nor U18407 (N_18407,N_17670,N_17287);
and U18408 (N_18408,N_17606,N_17628);
nor U18409 (N_18409,N_17706,N_17873);
xnor U18410 (N_18410,N_17814,N_17436);
or U18411 (N_18411,N_17910,N_17003);
nand U18412 (N_18412,N_17185,N_17889);
nor U18413 (N_18413,N_17761,N_17112);
or U18414 (N_18414,N_17514,N_17906);
nand U18415 (N_18415,N_17512,N_17908);
and U18416 (N_18416,N_17716,N_17052);
nand U18417 (N_18417,N_17678,N_17945);
nor U18418 (N_18418,N_17983,N_17480);
nor U18419 (N_18419,N_17836,N_17351);
and U18420 (N_18420,N_17488,N_17062);
and U18421 (N_18421,N_17082,N_17586);
xnor U18422 (N_18422,N_17762,N_17316);
or U18423 (N_18423,N_17895,N_17043);
nand U18424 (N_18424,N_17443,N_17608);
nor U18425 (N_18425,N_17680,N_17114);
and U18426 (N_18426,N_17194,N_17955);
xnor U18427 (N_18427,N_17530,N_17771);
and U18428 (N_18428,N_17525,N_17232);
xor U18429 (N_18429,N_17332,N_17779);
and U18430 (N_18430,N_17498,N_17793);
nand U18431 (N_18431,N_17439,N_17394);
nor U18432 (N_18432,N_17022,N_17671);
nor U18433 (N_18433,N_17857,N_17758);
and U18434 (N_18434,N_17046,N_17100);
or U18435 (N_18435,N_17079,N_17620);
nand U18436 (N_18436,N_17750,N_17528);
nand U18437 (N_18437,N_17424,N_17925);
and U18438 (N_18438,N_17433,N_17227);
or U18439 (N_18439,N_17707,N_17946);
and U18440 (N_18440,N_17690,N_17254);
or U18441 (N_18441,N_17816,N_17321);
or U18442 (N_18442,N_17485,N_17187);
xnor U18443 (N_18443,N_17269,N_17786);
and U18444 (N_18444,N_17096,N_17936);
xor U18445 (N_18445,N_17702,N_17972);
nand U18446 (N_18446,N_17505,N_17858);
or U18447 (N_18447,N_17273,N_17546);
xor U18448 (N_18448,N_17646,N_17422);
nor U18449 (N_18449,N_17555,N_17590);
xor U18450 (N_18450,N_17914,N_17184);
or U18451 (N_18451,N_17357,N_17153);
nand U18452 (N_18452,N_17417,N_17624);
and U18453 (N_18453,N_17650,N_17181);
nand U18454 (N_18454,N_17742,N_17077);
nand U18455 (N_18455,N_17155,N_17017);
and U18456 (N_18456,N_17693,N_17929);
nand U18457 (N_18457,N_17799,N_17375);
xnor U18458 (N_18458,N_17075,N_17819);
nand U18459 (N_18459,N_17861,N_17838);
nor U18460 (N_18460,N_17881,N_17468);
nand U18461 (N_18461,N_17067,N_17621);
or U18462 (N_18462,N_17665,N_17940);
nor U18463 (N_18463,N_17031,N_17537);
or U18464 (N_18464,N_17317,N_17491);
nor U18465 (N_18465,N_17721,N_17717);
xnor U18466 (N_18466,N_17165,N_17844);
xnor U18467 (N_18467,N_17478,N_17425);
and U18468 (N_18468,N_17994,N_17872);
xnor U18469 (N_18469,N_17362,N_17767);
nor U18470 (N_18470,N_17261,N_17026);
nand U18471 (N_18471,N_17568,N_17866);
and U18472 (N_18472,N_17772,N_17928);
nand U18473 (N_18473,N_17888,N_17652);
nand U18474 (N_18474,N_17871,N_17579);
nand U18475 (N_18475,N_17496,N_17744);
or U18476 (N_18476,N_17781,N_17730);
or U18477 (N_18477,N_17511,N_17842);
nor U18478 (N_18478,N_17285,N_17150);
nor U18479 (N_18479,N_17110,N_17626);
nand U18480 (N_18480,N_17550,N_17487);
or U18481 (N_18481,N_17712,N_17630);
xnor U18482 (N_18482,N_17271,N_17386);
and U18483 (N_18483,N_17901,N_17573);
nand U18484 (N_18484,N_17963,N_17016);
nor U18485 (N_18485,N_17378,N_17476);
nor U18486 (N_18486,N_17147,N_17236);
nand U18487 (N_18487,N_17984,N_17544);
nor U18488 (N_18488,N_17564,N_17899);
nand U18489 (N_18489,N_17483,N_17475);
or U18490 (N_18490,N_17330,N_17938);
xor U18491 (N_18491,N_17830,N_17093);
nor U18492 (N_18492,N_17915,N_17289);
nor U18493 (N_18493,N_17655,N_17619);
nor U18494 (N_18494,N_17056,N_17876);
nor U18495 (N_18495,N_17182,N_17073);
or U18496 (N_18496,N_17224,N_17890);
and U18497 (N_18497,N_17128,N_17030);
nand U18498 (N_18498,N_17775,N_17360);
nand U18499 (N_18499,N_17024,N_17613);
and U18500 (N_18500,N_17688,N_17515);
and U18501 (N_18501,N_17608,N_17378);
nand U18502 (N_18502,N_17782,N_17854);
xor U18503 (N_18503,N_17693,N_17350);
xor U18504 (N_18504,N_17606,N_17521);
and U18505 (N_18505,N_17271,N_17278);
nor U18506 (N_18506,N_17423,N_17657);
nand U18507 (N_18507,N_17285,N_17740);
and U18508 (N_18508,N_17879,N_17657);
xor U18509 (N_18509,N_17774,N_17845);
nor U18510 (N_18510,N_17325,N_17324);
nand U18511 (N_18511,N_17407,N_17642);
and U18512 (N_18512,N_17013,N_17183);
or U18513 (N_18513,N_17468,N_17363);
and U18514 (N_18514,N_17775,N_17664);
or U18515 (N_18515,N_17333,N_17550);
nor U18516 (N_18516,N_17765,N_17178);
xor U18517 (N_18517,N_17509,N_17342);
nand U18518 (N_18518,N_17954,N_17030);
nor U18519 (N_18519,N_17600,N_17619);
nand U18520 (N_18520,N_17907,N_17155);
nand U18521 (N_18521,N_17115,N_17114);
or U18522 (N_18522,N_17148,N_17953);
or U18523 (N_18523,N_17306,N_17132);
or U18524 (N_18524,N_17262,N_17694);
and U18525 (N_18525,N_17511,N_17556);
or U18526 (N_18526,N_17441,N_17936);
or U18527 (N_18527,N_17490,N_17125);
and U18528 (N_18528,N_17136,N_17216);
nor U18529 (N_18529,N_17874,N_17181);
or U18530 (N_18530,N_17226,N_17889);
or U18531 (N_18531,N_17044,N_17610);
and U18532 (N_18532,N_17250,N_17103);
nand U18533 (N_18533,N_17137,N_17715);
nand U18534 (N_18534,N_17039,N_17683);
and U18535 (N_18535,N_17671,N_17388);
nand U18536 (N_18536,N_17597,N_17058);
or U18537 (N_18537,N_17161,N_17391);
or U18538 (N_18538,N_17571,N_17534);
or U18539 (N_18539,N_17809,N_17961);
and U18540 (N_18540,N_17449,N_17737);
or U18541 (N_18541,N_17110,N_17322);
and U18542 (N_18542,N_17427,N_17515);
nand U18543 (N_18543,N_17176,N_17585);
nor U18544 (N_18544,N_17936,N_17829);
or U18545 (N_18545,N_17700,N_17061);
nor U18546 (N_18546,N_17867,N_17531);
and U18547 (N_18547,N_17141,N_17272);
and U18548 (N_18548,N_17608,N_17611);
and U18549 (N_18549,N_17372,N_17636);
xor U18550 (N_18550,N_17845,N_17812);
and U18551 (N_18551,N_17549,N_17294);
or U18552 (N_18552,N_17147,N_17115);
or U18553 (N_18553,N_17888,N_17040);
or U18554 (N_18554,N_17317,N_17111);
and U18555 (N_18555,N_17117,N_17970);
nor U18556 (N_18556,N_17182,N_17710);
nor U18557 (N_18557,N_17982,N_17994);
nor U18558 (N_18558,N_17381,N_17900);
xor U18559 (N_18559,N_17652,N_17614);
or U18560 (N_18560,N_17200,N_17678);
nor U18561 (N_18561,N_17475,N_17675);
xor U18562 (N_18562,N_17912,N_17272);
or U18563 (N_18563,N_17829,N_17856);
or U18564 (N_18564,N_17175,N_17643);
nand U18565 (N_18565,N_17835,N_17862);
xnor U18566 (N_18566,N_17136,N_17668);
nor U18567 (N_18567,N_17690,N_17553);
xor U18568 (N_18568,N_17871,N_17893);
nand U18569 (N_18569,N_17822,N_17724);
nor U18570 (N_18570,N_17217,N_17716);
nor U18571 (N_18571,N_17620,N_17881);
or U18572 (N_18572,N_17561,N_17752);
nor U18573 (N_18573,N_17492,N_17335);
nor U18574 (N_18574,N_17067,N_17822);
nand U18575 (N_18575,N_17181,N_17446);
or U18576 (N_18576,N_17688,N_17589);
or U18577 (N_18577,N_17032,N_17058);
nand U18578 (N_18578,N_17064,N_17806);
and U18579 (N_18579,N_17013,N_17912);
nor U18580 (N_18580,N_17265,N_17075);
nor U18581 (N_18581,N_17357,N_17775);
or U18582 (N_18582,N_17346,N_17266);
nor U18583 (N_18583,N_17027,N_17136);
nor U18584 (N_18584,N_17163,N_17034);
nor U18585 (N_18585,N_17558,N_17883);
nand U18586 (N_18586,N_17583,N_17680);
nor U18587 (N_18587,N_17419,N_17732);
or U18588 (N_18588,N_17801,N_17414);
nor U18589 (N_18589,N_17393,N_17512);
nor U18590 (N_18590,N_17364,N_17535);
and U18591 (N_18591,N_17509,N_17744);
or U18592 (N_18592,N_17314,N_17247);
and U18593 (N_18593,N_17611,N_17452);
or U18594 (N_18594,N_17950,N_17230);
xor U18595 (N_18595,N_17341,N_17580);
and U18596 (N_18596,N_17680,N_17881);
nand U18597 (N_18597,N_17626,N_17386);
nand U18598 (N_18598,N_17460,N_17177);
and U18599 (N_18599,N_17061,N_17659);
xnor U18600 (N_18600,N_17719,N_17876);
nor U18601 (N_18601,N_17483,N_17264);
nand U18602 (N_18602,N_17650,N_17955);
nor U18603 (N_18603,N_17529,N_17243);
or U18604 (N_18604,N_17948,N_17347);
nand U18605 (N_18605,N_17334,N_17888);
nor U18606 (N_18606,N_17479,N_17310);
nor U18607 (N_18607,N_17758,N_17141);
or U18608 (N_18608,N_17266,N_17572);
nor U18609 (N_18609,N_17410,N_17666);
xor U18610 (N_18610,N_17603,N_17482);
or U18611 (N_18611,N_17862,N_17576);
nor U18612 (N_18612,N_17384,N_17458);
and U18613 (N_18613,N_17243,N_17921);
nor U18614 (N_18614,N_17367,N_17157);
or U18615 (N_18615,N_17057,N_17799);
nand U18616 (N_18616,N_17680,N_17637);
and U18617 (N_18617,N_17769,N_17290);
nor U18618 (N_18618,N_17921,N_17478);
or U18619 (N_18619,N_17562,N_17656);
or U18620 (N_18620,N_17507,N_17602);
and U18621 (N_18621,N_17214,N_17008);
nand U18622 (N_18622,N_17901,N_17560);
nand U18623 (N_18623,N_17496,N_17995);
and U18624 (N_18624,N_17605,N_17167);
or U18625 (N_18625,N_17048,N_17732);
or U18626 (N_18626,N_17713,N_17200);
and U18627 (N_18627,N_17190,N_17175);
or U18628 (N_18628,N_17563,N_17070);
nand U18629 (N_18629,N_17535,N_17076);
or U18630 (N_18630,N_17549,N_17869);
xor U18631 (N_18631,N_17402,N_17367);
nand U18632 (N_18632,N_17813,N_17072);
nor U18633 (N_18633,N_17186,N_17931);
nor U18634 (N_18634,N_17313,N_17040);
nor U18635 (N_18635,N_17856,N_17413);
or U18636 (N_18636,N_17224,N_17824);
and U18637 (N_18637,N_17220,N_17055);
nor U18638 (N_18638,N_17486,N_17587);
xor U18639 (N_18639,N_17733,N_17402);
or U18640 (N_18640,N_17263,N_17227);
nand U18641 (N_18641,N_17061,N_17142);
nand U18642 (N_18642,N_17491,N_17706);
or U18643 (N_18643,N_17176,N_17788);
nor U18644 (N_18644,N_17460,N_17559);
or U18645 (N_18645,N_17476,N_17035);
or U18646 (N_18646,N_17415,N_17724);
or U18647 (N_18647,N_17160,N_17988);
xor U18648 (N_18648,N_17039,N_17778);
and U18649 (N_18649,N_17282,N_17946);
nand U18650 (N_18650,N_17173,N_17744);
nor U18651 (N_18651,N_17676,N_17237);
nor U18652 (N_18652,N_17460,N_17601);
nor U18653 (N_18653,N_17130,N_17110);
and U18654 (N_18654,N_17760,N_17471);
nand U18655 (N_18655,N_17898,N_17764);
nand U18656 (N_18656,N_17143,N_17549);
nand U18657 (N_18657,N_17496,N_17913);
nand U18658 (N_18658,N_17885,N_17905);
nor U18659 (N_18659,N_17581,N_17128);
nand U18660 (N_18660,N_17047,N_17713);
nand U18661 (N_18661,N_17045,N_17703);
or U18662 (N_18662,N_17876,N_17470);
and U18663 (N_18663,N_17776,N_17056);
nand U18664 (N_18664,N_17448,N_17462);
or U18665 (N_18665,N_17012,N_17135);
and U18666 (N_18666,N_17806,N_17945);
nor U18667 (N_18667,N_17894,N_17773);
xnor U18668 (N_18668,N_17719,N_17685);
nor U18669 (N_18669,N_17920,N_17513);
or U18670 (N_18670,N_17519,N_17785);
or U18671 (N_18671,N_17238,N_17720);
and U18672 (N_18672,N_17164,N_17611);
and U18673 (N_18673,N_17918,N_17584);
xnor U18674 (N_18674,N_17325,N_17639);
nand U18675 (N_18675,N_17627,N_17131);
nor U18676 (N_18676,N_17005,N_17682);
nand U18677 (N_18677,N_17988,N_17197);
or U18678 (N_18678,N_17696,N_17374);
and U18679 (N_18679,N_17894,N_17642);
or U18680 (N_18680,N_17184,N_17904);
nor U18681 (N_18681,N_17385,N_17305);
nor U18682 (N_18682,N_17723,N_17766);
nand U18683 (N_18683,N_17313,N_17769);
nand U18684 (N_18684,N_17030,N_17649);
nor U18685 (N_18685,N_17851,N_17418);
nor U18686 (N_18686,N_17305,N_17234);
and U18687 (N_18687,N_17411,N_17637);
and U18688 (N_18688,N_17867,N_17313);
or U18689 (N_18689,N_17966,N_17349);
xor U18690 (N_18690,N_17670,N_17473);
nand U18691 (N_18691,N_17655,N_17486);
nand U18692 (N_18692,N_17935,N_17679);
and U18693 (N_18693,N_17248,N_17029);
or U18694 (N_18694,N_17780,N_17598);
and U18695 (N_18695,N_17017,N_17543);
or U18696 (N_18696,N_17846,N_17596);
and U18697 (N_18697,N_17366,N_17850);
and U18698 (N_18698,N_17213,N_17593);
nand U18699 (N_18699,N_17111,N_17389);
nand U18700 (N_18700,N_17966,N_17116);
and U18701 (N_18701,N_17162,N_17556);
nand U18702 (N_18702,N_17922,N_17389);
or U18703 (N_18703,N_17223,N_17912);
or U18704 (N_18704,N_17947,N_17402);
and U18705 (N_18705,N_17094,N_17112);
nand U18706 (N_18706,N_17277,N_17015);
nor U18707 (N_18707,N_17499,N_17796);
nand U18708 (N_18708,N_17213,N_17641);
nand U18709 (N_18709,N_17032,N_17026);
and U18710 (N_18710,N_17329,N_17971);
or U18711 (N_18711,N_17625,N_17114);
xnor U18712 (N_18712,N_17922,N_17964);
and U18713 (N_18713,N_17084,N_17816);
nor U18714 (N_18714,N_17401,N_17578);
or U18715 (N_18715,N_17001,N_17217);
and U18716 (N_18716,N_17047,N_17053);
or U18717 (N_18717,N_17263,N_17709);
or U18718 (N_18718,N_17854,N_17168);
or U18719 (N_18719,N_17678,N_17428);
xor U18720 (N_18720,N_17822,N_17735);
nand U18721 (N_18721,N_17094,N_17236);
xnor U18722 (N_18722,N_17655,N_17733);
or U18723 (N_18723,N_17663,N_17745);
and U18724 (N_18724,N_17166,N_17631);
or U18725 (N_18725,N_17573,N_17226);
nand U18726 (N_18726,N_17125,N_17174);
or U18727 (N_18727,N_17245,N_17628);
and U18728 (N_18728,N_17131,N_17454);
nand U18729 (N_18729,N_17491,N_17606);
nor U18730 (N_18730,N_17245,N_17330);
nand U18731 (N_18731,N_17961,N_17040);
nor U18732 (N_18732,N_17588,N_17418);
xor U18733 (N_18733,N_17233,N_17706);
nand U18734 (N_18734,N_17495,N_17179);
and U18735 (N_18735,N_17263,N_17348);
nor U18736 (N_18736,N_17546,N_17262);
or U18737 (N_18737,N_17668,N_17769);
nor U18738 (N_18738,N_17527,N_17798);
or U18739 (N_18739,N_17561,N_17037);
nor U18740 (N_18740,N_17505,N_17313);
nand U18741 (N_18741,N_17731,N_17074);
or U18742 (N_18742,N_17029,N_17779);
nand U18743 (N_18743,N_17477,N_17679);
and U18744 (N_18744,N_17341,N_17837);
or U18745 (N_18745,N_17774,N_17417);
nor U18746 (N_18746,N_17852,N_17866);
nand U18747 (N_18747,N_17877,N_17707);
nor U18748 (N_18748,N_17243,N_17975);
nor U18749 (N_18749,N_17177,N_17715);
nor U18750 (N_18750,N_17341,N_17897);
or U18751 (N_18751,N_17243,N_17354);
or U18752 (N_18752,N_17602,N_17249);
or U18753 (N_18753,N_17588,N_17831);
or U18754 (N_18754,N_17549,N_17968);
and U18755 (N_18755,N_17900,N_17157);
nor U18756 (N_18756,N_17137,N_17834);
nor U18757 (N_18757,N_17046,N_17712);
nand U18758 (N_18758,N_17123,N_17547);
or U18759 (N_18759,N_17786,N_17979);
nor U18760 (N_18760,N_17843,N_17087);
or U18761 (N_18761,N_17291,N_17347);
and U18762 (N_18762,N_17681,N_17647);
nor U18763 (N_18763,N_17099,N_17130);
nor U18764 (N_18764,N_17782,N_17915);
or U18765 (N_18765,N_17815,N_17638);
nand U18766 (N_18766,N_17143,N_17423);
and U18767 (N_18767,N_17973,N_17615);
nand U18768 (N_18768,N_17715,N_17101);
and U18769 (N_18769,N_17409,N_17701);
nand U18770 (N_18770,N_17971,N_17910);
nor U18771 (N_18771,N_17342,N_17722);
and U18772 (N_18772,N_17417,N_17749);
nand U18773 (N_18773,N_17144,N_17092);
xor U18774 (N_18774,N_17369,N_17496);
and U18775 (N_18775,N_17785,N_17964);
xnor U18776 (N_18776,N_17782,N_17507);
and U18777 (N_18777,N_17296,N_17519);
nor U18778 (N_18778,N_17069,N_17127);
and U18779 (N_18779,N_17836,N_17702);
or U18780 (N_18780,N_17379,N_17800);
and U18781 (N_18781,N_17974,N_17951);
or U18782 (N_18782,N_17738,N_17335);
nand U18783 (N_18783,N_17353,N_17149);
and U18784 (N_18784,N_17583,N_17134);
nand U18785 (N_18785,N_17497,N_17075);
nand U18786 (N_18786,N_17055,N_17311);
nor U18787 (N_18787,N_17476,N_17111);
xor U18788 (N_18788,N_17442,N_17328);
and U18789 (N_18789,N_17295,N_17473);
or U18790 (N_18790,N_17502,N_17204);
nand U18791 (N_18791,N_17807,N_17434);
nor U18792 (N_18792,N_17960,N_17273);
or U18793 (N_18793,N_17203,N_17382);
nor U18794 (N_18794,N_17035,N_17674);
nor U18795 (N_18795,N_17507,N_17260);
nor U18796 (N_18796,N_17958,N_17190);
nor U18797 (N_18797,N_17313,N_17755);
nor U18798 (N_18798,N_17929,N_17205);
or U18799 (N_18799,N_17517,N_17259);
or U18800 (N_18800,N_17911,N_17923);
nor U18801 (N_18801,N_17111,N_17933);
nor U18802 (N_18802,N_17116,N_17984);
or U18803 (N_18803,N_17461,N_17114);
or U18804 (N_18804,N_17804,N_17812);
nor U18805 (N_18805,N_17984,N_17783);
and U18806 (N_18806,N_17706,N_17705);
and U18807 (N_18807,N_17512,N_17025);
nor U18808 (N_18808,N_17029,N_17873);
or U18809 (N_18809,N_17477,N_17855);
nor U18810 (N_18810,N_17983,N_17197);
nand U18811 (N_18811,N_17219,N_17154);
and U18812 (N_18812,N_17324,N_17241);
nor U18813 (N_18813,N_17633,N_17826);
or U18814 (N_18814,N_17290,N_17130);
nand U18815 (N_18815,N_17415,N_17983);
xor U18816 (N_18816,N_17507,N_17826);
nor U18817 (N_18817,N_17374,N_17457);
nand U18818 (N_18818,N_17958,N_17706);
or U18819 (N_18819,N_17108,N_17492);
or U18820 (N_18820,N_17030,N_17274);
and U18821 (N_18821,N_17420,N_17812);
and U18822 (N_18822,N_17564,N_17113);
and U18823 (N_18823,N_17003,N_17955);
nand U18824 (N_18824,N_17628,N_17921);
xor U18825 (N_18825,N_17577,N_17733);
xnor U18826 (N_18826,N_17544,N_17668);
xor U18827 (N_18827,N_17398,N_17856);
nand U18828 (N_18828,N_17611,N_17526);
or U18829 (N_18829,N_17957,N_17970);
nand U18830 (N_18830,N_17648,N_17540);
nor U18831 (N_18831,N_17168,N_17660);
xor U18832 (N_18832,N_17923,N_17990);
or U18833 (N_18833,N_17293,N_17684);
nor U18834 (N_18834,N_17428,N_17172);
and U18835 (N_18835,N_17240,N_17222);
nor U18836 (N_18836,N_17226,N_17892);
or U18837 (N_18837,N_17034,N_17317);
and U18838 (N_18838,N_17835,N_17044);
and U18839 (N_18839,N_17367,N_17177);
nor U18840 (N_18840,N_17909,N_17700);
nand U18841 (N_18841,N_17894,N_17029);
and U18842 (N_18842,N_17692,N_17661);
or U18843 (N_18843,N_17867,N_17983);
nor U18844 (N_18844,N_17690,N_17772);
nor U18845 (N_18845,N_17252,N_17803);
and U18846 (N_18846,N_17937,N_17397);
nor U18847 (N_18847,N_17049,N_17364);
nand U18848 (N_18848,N_17892,N_17666);
and U18849 (N_18849,N_17578,N_17594);
and U18850 (N_18850,N_17215,N_17016);
xnor U18851 (N_18851,N_17391,N_17025);
and U18852 (N_18852,N_17787,N_17519);
and U18853 (N_18853,N_17372,N_17832);
and U18854 (N_18854,N_17419,N_17299);
or U18855 (N_18855,N_17153,N_17659);
and U18856 (N_18856,N_17068,N_17665);
and U18857 (N_18857,N_17186,N_17975);
and U18858 (N_18858,N_17025,N_17794);
and U18859 (N_18859,N_17625,N_17265);
nand U18860 (N_18860,N_17783,N_17293);
or U18861 (N_18861,N_17851,N_17293);
and U18862 (N_18862,N_17782,N_17461);
and U18863 (N_18863,N_17653,N_17708);
nand U18864 (N_18864,N_17346,N_17106);
nor U18865 (N_18865,N_17807,N_17368);
and U18866 (N_18866,N_17668,N_17104);
and U18867 (N_18867,N_17538,N_17520);
nand U18868 (N_18868,N_17952,N_17353);
and U18869 (N_18869,N_17649,N_17658);
or U18870 (N_18870,N_17626,N_17248);
nand U18871 (N_18871,N_17764,N_17002);
and U18872 (N_18872,N_17318,N_17027);
and U18873 (N_18873,N_17438,N_17793);
nor U18874 (N_18874,N_17115,N_17383);
nand U18875 (N_18875,N_17595,N_17115);
or U18876 (N_18876,N_17504,N_17984);
nand U18877 (N_18877,N_17744,N_17718);
and U18878 (N_18878,N_17223,N_17986);
nand U18879 (N_18879,N_17866,N_17065);
and U18880 (N_18880,N_17184,N_17836);
or U18881 (N_18881,N_17818,N_17848);
and U18882 (N_18882,N_17894,N_17229);
xnor U18883 (N_18883,N_17997,N_17632);
and U18884 (N_18884,N_17204,N_17719);
and U18885 (N_18885,N_17249,N_17982);
and U18886 (N_18886,N_17154,N_17020);
or U18887 (N_18887,N_17403,N_17358);
or U18888 (N_18888,N_17233,N_17777);
and U18889 (N_18889,N_17516,N_17155);
xor U18890 (N_18890,N_17692,N_17357);
or U18891 (N_18891,N_17461,N_17196);
nand U18892 (N_18892,N_17570,N_17211);
nand U18893 (N_18893,N_17316,N_17019);
nor U18894 (N_18894,N_17253,N_17405);
nor U18895 (N_18895,N_17333,N_17472);
and U18896 (N_18896,N_17930,N_17418);
nand U18897 (N_18897,N_17651,N_17308);
nor U18898 (N_18898,N_17566,N_17079);
or U18899 (N_18899,N_17883,N_17763);
nor U18900 (N_18900,N_17600,N_17339);
nor U18901 (N_18901,N_17120,N_17197);
nand U18902 (N_18902,N_17214,N_17928);
and U18903 (N_18903,N_17064,N_17237);
or U18904 (N_18904,N_17541,N_17781);
xor U18905 (N_18905,N_17842,N_17135);
nor U18906 (N_18906,N_17429,N_17049);
nand U18907 (N_18907,N_17088,N_17552);
and U18908 (N_18908,N_17231,N_17281);
nand U18909 (N_18909,N_17346,N_17080);
and U18910 (N_18910,N_17300,N_17210);
xnor U18911 (N_18911,N_17635,N_17001);
and U18912 (N_18912,N_17209,N_17750);
nand U18913 (N_18913,N_17996,N_17604);
and U18914 (N_18914,N_17476,N_17102);
or U18915 (N_18915,N_17015,N_17278);
and U18916 (N_18916,N_17458,N_17502);
nand U18917 (N_18917,N_17330,N_17170);
nor U18918 (N_18918,N_17340,N_17401);
and U18919 (N_18919,N_17559,N_17736);
or U18920 (N_18920,N_17905,N_17874);
nand U18921 (N_18921,N_17170,N_17306);
nor U18922 (N_18922,N_17928,N_17219);
nand U18923 (N_18923,N_17186,N_17275);
or U18924 (N_18924,N_17912,N_17806);
nand U18925 (N_18925,N_17515,N_17074);
nand U18926 (N_18926,N_17267,N_17289);
nand U18927 (N_18927,N_17497,N_17795);
nor U18928 (N_18928,N_17583,N_17032);
nand U18929 (N_18929,N_17529,N_17196);
nand U18930 (N_18930,N_17926,N_17400);
nor U18931 (N_18931,N_17629,N_17500);
and U18932 (N_18932,N_17643,N_17185);
nand U18933 (N_18933,N_17460,N_17369);
and U18934 (N_18934,N_17770,N_17169);
or U18935 (N_18935,N_17451,N_17564);
and U18936 (N_18936,N_17415,N_17496);
nor U18937 (N_18937,N_17777,N_17704);
and U18938 (N_18938,N_17853,N_17568);
nand U18939 (N_18939,N_17524,N_17601);
nor U18940 (N_18940,N_17492,N_17254);
nand U18941 (N_18941,N_17975,N_17690);
or U18942 (N_18942,N_17659,N_17243);
nor U18943 (N_18943,N_17556,N_17488);
or U18944 (N_18944,N_17543,N_17762);
nor U18945 (N_18945,N_17904,N_17418);
nor U18946 (N_18946,N_17351,N_17357);
and U18947 (N_18947,N_17625,N_17093);
nand U18948 (N_18948,N_17642,N_17050);
and U18949 (N_18949,N_17466,N_17618);
nor U18950 (N_18950,N_17659,N_17033);
xor U18951 (N_18951,N_17768,N_17601);
nor U18952 (N_18952,N_17920,N_17093);
xor U18953 (N_18953,N_17702,N_17299);
and U18954 (N_18954,N_17820,N_17572);
nand U18955 (N_18955,N_17065,N_17654);
nor U18956 (N_18956,N_17374,N_17612);
and U18957 (N_18957,N_17526,N_17146);
or U18958 (N_18958,N_17472,N_17561);
and U18959 (N_18959,N_17425,N_17299);
or U18960 (N_18960,N_17701,N_17950);
nand U18961 (N_18961,N_17974,N_17837);
nand U18962 (N_18962,N_17381,N_17278);
or U18963 (N_18963,N_17224,N_17367);
or U18964 (N_18964,N_17970,N_17424);
or U18965 (N_18965,N_17741,N_17936);
nand U18966 (N_18966,N_17300,N_17279);
nand U18967 (N_18967,N_17424,N_17703);
or U18968 (N_18968,N_17736,N_17516);
and U18969 (N_18969,N_17124,N_17700);
nand U18970 (N_18970,N_17112,N_17480);
or U18971 (N_18971,N_17902,N_17264);
nand U18972 (N_18972,N_17994,N_17643);
xor U18973 (N_18973,N_17421,N_17957);
and U18974 (N_18974,N_17516,N_17554);
xor U18975 (N_18975,N_17807,N_17280);
nor U18976 (N_18976,N_17647,N_17311);
and U18977 (N_18977,N_17176,N_17073);
nand U18978 (N_18978,N_17085,N_17993);
or U18979 (N_18979,N_17540,N_17451);
and U18980 (N_18980,N_17489,N_17662);
nor U18981 (N_18981,N_17201,N_17040);
xor U18982 (N_18982,N_17016,N_17104);
nor U18983 (N_18983,N_17746,N_17687);
nor U18984 (N_18984,N_17443,N_17166);
and U18985 (N_18985,N_17609,N_17373);
nand U18986 (N_18986,N_17746,N_17217);
and U18987 (N_18987,N_17994,N_17259);
nand U18988 (N_18988,N_17576,N_17267);
nand U18989 (N_18989,N_17839,N_17127);
nor U18990 (N_18990,N_17551,N_17230);
nor U18991 (N_18991,N_17135,N_17070);
or U18992 (N_18992,N_17342,N_17638);
nand U18993 (N_18993,N_17322,N_17872);
nand U18994 (N_18994,N_17807,N_17518);
or U18995 (N_18995,N_17410,N_17362);
and U18996 (N_18996,N_17300,N_17644);
xor U18997 (N_18997,N_17161,N_17691);
nor U18998 (N_18998,N_17983,N_17424);
nand U18999 (N_18999,N_17957,N_17842);
or U19000 (N_19000,N_18215,N_18315);
nor U19001 (N_19001,N_18988,N_18271);
or U19002 (N_19002,N_18930,N_18054);
or U19003 (N_19003,N_18593,N_18322);
nor U19004 (N_19004,N_18479,N_18784);
xnor U19005 (N_19005,N_18824,N_18006);
nand U19006 (N_19006,N_18401,N_18073);
and U19007 (N_19007,N_18901,N_18502);
nand U19008 (N_19008,N_18413,N_18772);
xnor U19009 (N_19009,N_18122,N_18009);
nor U19010 (N_19010,N_18704,N_18022);
or U19011 (N_19011,N_18735,N_18426);
or U19012 (N_19012,N_18695,N_18480);
and U19013 (N_19013,N_18746,N_18703);
or U19014 (N_19014,N_18339,N_18814);
nand U19015 (N_19015,N_18437,N_18892);
nor U19016 (N_19016,N_18218,N_18420);
and U19017 (N_19017,N_18485,N_18312);
nand U19018 (N_19018,N_18700,N_18782);
or U19019 (N_19019,N_18893,N_18591);
nor U19020 (N_19020,N_18273,N_18499);
or U19021 (N_19021,N_18369,N_18962);
and U19022 (N_19022,N_18622,N_18920);
or U19023 (N_19023,N_18257,N_18002);
nor U19024 (N_19024,N_18136,N_18840);
nor U19025 (N_19025,N_18759,N_18974);
nor U19026 (N_19026,N_18605,N_18826);
and U19027 (N_19027,N_18590,N_18142);
nor U19028 (N_19028,N_18262,N_18167);
nor U19029 (N_19029,N_18965,N_18344);
and U19030 (N_19030,N_18579,N_18847);
or U19031 (N_19031,N_18155,N_18790);
nand U19032 (N_19032,N_18395,N_18302);
nand U19033 (N_19033,N_18056,N_18690);
or U19034 (N_19034,N_18752,N_18186);
or U19035 (N_19035,N_18099,N_18564);
nor U19036 (N_19036,N_18329,N_18554);
nor U19037 (N_19037,N_18280,N_18341);
nor U19038 (N_19038,N_18209,N_18323);
nor U19039 (N_19039,N_18392,N_18786);
and U19040 (N_19040,N_18873,N_18774);
xnor U19041 (N_19041,N_18190,N_18545);
or U19042 (N_19042,N_18130,N_18069);
or U19043 (N_19043,N_18906,N_18515);
or U19044 (N_19044,N_18574,N_18614);
nor U19045 (N_19045,N_18512,N_18184);
or U19046 (N_19046,N_18823,N_18958);
or U19047 (N_19047,N_18491,N_18366);
and U19048 (N_19048,N_18345,N_18368);
and U19049 (N_19049,N_18381,N_18351);
nor U19050 (N_19050,N_18060,N_18405);
nand U19051 (N_19051,N_18693,N_18361);
and U19052 (N_19052,N_18792,N_18469);
or U19053 (N_19053,N_18033,N_18898);
nand U19054 (N_19054,N_18818,N_18318);
or U19055 (N_19055,N_18720,N_18173);
nor U19056 (N_19056,N_18441,N_18769);
nor U19057 (N_19057,N_18585,N_18394);
nand U19058 (N_19058,N_18278,N_18996);
or U19059 (N_19059,N_18596,N_18043);
xor U19060 (N_19060,N_18749,N_18047);
or U19061 (N_19061,N_18178,N_18011);
or U19062 (N_19062,N_18269,N_18014);
and U19063 (N_19063,N_18087,N_18194);
nor U19064 (N_19064,N_18643,N_18866);
nand U19065 (N_19065,N_18737,N_18507);
or U19066 (N_19066,N_18994,N_18125);
nor U19067 (N_19067,N_18148,N_18003);
or U19068 (N_19068,N_18683,N_18147);
nor U19069 (N_19069,N_18295,N_18227);
xnor U19070 (N_19070,N_18281,N_18832);
xnor U19071 (N_19071,N_18694,N_18844);
xnor U19072 (N_19072,N_18985,N_18386);
nand U19073 (N_19073,N_18428,N_18000);
nand U19074 (N_19074,N_18553,N_18598);
and U19075 (N_19075,N_18955,N_18275);
and U19076 (N_19076,N_18251,N_18114);
or U19077 (N_19077,N_18421,N_18384);
or U19078 (N_19078,N_18740,N_18686);
nor U19079 (N_19079,N_18036,N_18570);
and U19080 (N_19080,N_18243,N_18012);
nor U19081 (N_19081,N_18868,N_18748);
nor U19082 (N_19082,N_18317,N_18933);
nor U19083 (N_19083,N_18645,N_18017);
nand U19084 (N_19084,N_18666,N_18102);
nand U19085 (N_19085,N_18264,N_18037);
nor U19086 (N_19086,N_18468,N_18617);
nor U19087 (N_19087,N_18313,N_18723);
nand U19088 (N_19088,N_18482,N_18050);
and U19089 (N_19089,N_18846,N_18358);
or U19090 (N_19090,N_18821,N_18621);
and U19091 (N_19091,N_18766,N_18217);
nor U19092 (N_19092,N_18374,N_18795);
and U19093 (N_19093,N_18532,N_18279);
nor U19094 (N_19094,N_18623,N_18228);
nor U19095 (N_19095,N_18088,N_18884);
or U19096 (N_19096,N_18870,N_18926);
and U19097 (N_19097,N_18602,N_18747);
and U19098 (N_19098,N_18980,N_18013);
and U19099 (N_19099,N_18350,N_18265);
nor U19100 (N_19100,N_18454,N_18536);
and U19101 (N_19101,N_18908,N_18914);
nand U19102 (N_19102,N_18696,N_18547);
nand U19103 (N_19103,N_18411,N_18078);
nand U19104 (N_19104,N_18116,N_18449);
and U19105 (N_19105,N_18293,N_18803);
nor U19106 (N_19106,N_18673,N_18081);
and U19107 (N_19107,N_18342,N_18314);
and U19108 (N_19108,N_18305,N_18815);
nand U19109 (N_19109,N_18038,N_18352);
nor U19110 (N_19110,N_18164,N_18612);
or U19111 (N_19111,N_18885,N_18245);
nand U19112 (N_19112,N_18944,N_18326);
or U19113 (N_19113,N_18524,N_18562);
nor U19114 (N_19114,N_18438,N_18462);
or U19115 (N_19115,N_18927,N_18195);
nor U19116 (N_19116,N_18877,N_18229);
nor U19117 (N_19117,N_18058,N_18647);
nand U19118 (N_19118,N_18918,N_18519);
nor U19119 (N_19119,N_18239,N_18788);
or U19120 (N_19120,N_18583,N_18200);
xnor U19121 (N_19121,N_18939,N_18586);
or U19122 (N_19122,N_18198,N_18144);
nand U19123 (N_19123,N_18961,N_18811);
and U19124 (N_19124,N_18231,N_18722);
or U19125 (N_19125,N_18377,N_18283);
or U19126 (N_19126,N_18500,N_18387);
and U19127 (N_19127,N_18382,N_18808);
xor U19128 (N_19128,N_18890,N_18991);
nor U19129 (N_19129,N_18838,N_18005);
or U19130 (N_19130,N_18303,N_18616);
xor U19131 (N_19131,N_18842,N_18543);
and U19132 (N_19132,N_18340,N_18135);
or U19133 (N_19133,N_18767,N_18850);
and U19134 (N_19134,N_18389,N_18355);
nand U19135 (N_19135,N_18573,N_18796);
nand U19136 (N_19136,N_18169,N_18233);
nor U19137 (N_19137,N_18530,N_18242);
or U19138 (N_19138,N_18565,N_18743);
nor U19139 (N_19139,N_18813,N_18670);
xnor U19140 (N_19140,N_18127,N_18652);
and U19141 (N_19141,N_18529,N_18765);
xnor U19142 (N_19142,N_18959,N_18097);
nand U19143 (N_19143,N_18165,N_18268);
and U19144 (N_19144,N_18453,N_18249);
or U19145 (N_19145,N_18697,N_18456);
nor U19146 (N_19146,N_18076,N_18895);
nand U19147 (N_19147,N_18336,N_18535);
or U19148 (N_19148,N_18285,N_18220);
and U19149 (N_19149,N_18497,N_18781);
and U19150 (N_19150,N_18839,N_18856);
nand U19151 (N_19151,N_18396,N_18806);
or U19152 (N_19152,N_18379,N_18131);
xnor U19153 (N_19153,N_18637,N_18109);
or U19154 (N_19154,N_18849,N_18091);
or U19155 (N_19155,N_18051,N_18348);
nor U19156 (N_19156,N_18522,N_18121);
or U19157 (N_19157,N_18800,N_18124);
nor U19158 (N_19158,N_18653,N_18603);
xor U19159 (N_19159,N_18705,N_18223);
xnor U19160 (N_19160,N_18915,N_18455);
nand U19161 (N_19161,N_18618,N_18990);
nor U19162 (N_19162,N_18309,N_18301);
or U19163 (N_19163,N_18858,N_18646);
nor U19164 (N_19164,N_18947,N_18662);
and U19165 (N_19165,N_18129,N_18082);
or U19166 (N_19166,N_18756,N_18658);
and U19167 (N_19167,N_18070,N_18161);
nand U19168 (N_19168,N_18297,N_18528);
or U19169 (N_19169,N_18668,N_18357);
nand U19170 (N_19170,N_18913,N_18816);
nand U19171 (N_19171,N_18909,N_18044);
nor U19172 (N_19172,N_18648,N_18578);
nor U19173 (N_19173,N_18791,N_18773);
or U19174 (N_19174,N_18595,N_18065);
nor U19175 (N_19175,N_18584,N_18882);
and U19176 (N_19176,N_18942,N_18261);
and U19177 (N_19177,N_18968,N_18607);
nand U19178 (N_19178,N_18175,N_18707);
nand U19179 (N_19179,N_18534,N_18624);
nor U19180 (N_19180,N_18708,N_18887);
nand U19181 (N_19181,N_18140,N_18197);
and U19182 (N_19182,N_18644,N_18817);
or U19183 (N_19183,N_18483,N_18189);
nand U19184 (N_19184,N_18434,N_18032);
xnor U19185 (N_19185,N_18429,N_18030);
or U19186 (N_19186,N_18172,N_18879);
or U19187 (N_19187,N_18599,N_18236);
and U19188 (N_19188,N_18308,N_18291);
xnor U19189 (N_19189,N_18953,N_18508);
and U19190 (N_19190,N_18146,N_18202);
nand U19191 (N_19191,N_18829,N_18298);
nor U19192 (N_19192,N_18225,N_18853);
xor U19193 (N_19193,N_18831,N_18857);
nor U19194 (N_19194,N_18970,N_18098);
and U19195 (N_19195,N_18635,N_18779);
or U19196 (N_19196,N_18798,N_18698);
and U19197 (N_19197,N_18582,N_18263);
and U19198 (N_19198,N_18244,N_18042);
xor U19199 (N_19199,N_18610,N_18092);
or U19200 (N_19200,N_18477,N_18007);
nand U19201 (N_19201,N_18592,N_18992);
or U19202 (N_19202,N_18435,N_18799);
nand U19203 (N_19203,N_18110,N_18237);
and U19204 (N_19204,N_18094,N_18090);
nand U19205 (N_19205,N_18544,N_18728);
and U19206 (N_19206,N_18465,N_18692);
nand U19207 (N_19207,N_18932,N_18450);
xor U19208 (N_19208,N_18559,N_18423);
nor U19209 (N_19209,N_18075,N_18260);
nand U19210 (N_19210,N_18360,N_18810);
xnor U19211 (N_19211,N_18656,N_18675);
nor U19212 (N_19212,N_18928,N_18577);
nor U19213 (N_19213,N_18212,N_18805);
nand U19214 (N_19214,N_18201,N_18677);
and U19215 (N_19215,N_18757,N_18581);
nand U19216 (N_19216,N_18706,N_18134);
nor U19217 (N_19217,N_18923,N_18487);
nand U19218 (N_19218,N_18048,N_18936);
or U19219 (N_19219,N_18993,N_18967);
nor U19220 (N_19220,N_18112,N_18886);
xor U19221 (N_19221,N_18952,N_18398);
and U19222 (N_19222,N_18138,N_18203);
and U19223 (N_19223,N_18780,N_18270);
or U19224 (N_19224,N_18505,N_18854);
and U19225 (N_19225,N_18213,N_18654);
and U19226 (N_19226,N_18983,N_18383);
and U19227 (N_19227,N_18071,N_18179);
nand U19228 (N_19228,N_18035,N_18332);
nand U19229 (N_19229,N_18687,N_18630);
nor U19230 (N_19230,N_18207,N_18444);
and U19231 (N_19231,N_18163,N_18029);
or U19232 (N_19232,N_18316,N_18661);
nor U19233 (N_19233,N_18409,N_18682);
nor U19234 (N_19234,N_18074,N_18680);
nor U19235 (N_19235,N_18966,N_18981);
and U19236 (N_19236,N_18797,N_18860);
nand U19237 (N_19237,N_18376,N_18170);
and U19238 (N_19238,N_18555,N_18230);
and U19239 (N_19239,N_18615,N_18372);
nand U19240 (N_19240,N_18896,N_18594);
or U19241 (N_19241,N_18843,N_18496);
or U19242 (N_19242,N_18362,N_18427);
nor U19243 (N_19243,N_18182,N_18294);
nor U19244 (N_19244,N_18390,N_18328);
nand U19245 (N_19245,N_18253,N_18568);
and U19246 (N_19246,N_18222,N_18393);
nor U19247 (N_19247,N_18095,N_18904);
xor U19248 (N_19248,N_18715,N_18370);
or U19249 (N_19249,N_18168,N_18546);
nor U19250 (N_19250,N_18971,N_18324);
nor U19251 (N_19251,N_18567,N_18556);
and U19252 (N_19252,N_18008,N_18679);
nand U19253 (N_19253,N_18067,N_18123);
nor U19254 (N_19254,N_18558,N_18495);
nor U19255 (N_19255,N_18474,N_18712);
nor U19256 (N_19256,N_18059,N_18511);
and U19257 (N_19257,N_18457,N_18820);
and U19258 (N_19258,N_18149,N_18733);
xor U19259 (N_19259,N_18561,N_18141);
nand U19260 (N_19260,N_18721,N_18331);
nor U19261 (N_19261,N_18830,N_18763);
nor U19262 (N_19262,N_18311,N_18028);
and U19263 (N_19263,N_18986,N_18925);
and U19264 (N_19264,N_18284,N_18064);
nor U19265 (N_19265,N_18246,N_18948);
or U19266 (N_19266,N_18776,N_18041);
and U19267 (N_19267,N_18589,N_18957);
or U19268 (N_19268,N_18062,N_18256);
and U19269 (N_19269,N_18804,N_18717);
or U19270 (N_19270,N_18649,N_18196);
nand U19271 (N_19271,N_18629,N_18750);
or U19272 (N_19272,N_18288,N_18964);
and U19273 (N_19273,N_18335,N_18902);
nand U19274 (N_19274,N_18490,N_18922);
nor U19275 (N_19275,N_18688,N_18461);
and U19276 (N_19276,N_18601,N_18631);
or U19277 (N_19277,N_18825,N_18158);
or U19278 (N_19278,N_18040,N_18852);
or U19279 (N_19279,N_18373,N_18880);
xor U19280 (N_19280,N_18299,N_18151);
or U19281 (N_19281,N_18604,N_18995);
nor U19282 (N_19282,N_18481,N_18210);
nand U19283 (N_19283,N_18464,N_18118);
nor U19284 (N_19284,N_18533,N_18492);
nand U19285 (N_19285,N_18354,N_18083);
nor U19286 (N_19286,N_18793,N_18600);
or U19287 (N_19287,N_18470,N_18636);
and U19288 (N_19288,N_18476,N_18691);
xnor U19289 (N_19289,N_18641,N_18219);
xor U19290 (N_19290,N_18319,N_18527);
nor U19291 (N_19291,N_18126,N_18552);
or U19292 (N_19292,N_18451,N_18024);
nor U19293 (N_19293,N_18171,N_18238);
nand U19294 (N_19294,N_18224,N_18452);
and U19295 (N_19295,N_18199,N_18878);
nor U19296 (N_19296,N_18910,N_18183);
nand U19297 (N_19297,N_18388,N_18760);
xor U19298 (N_19298,N_18247,N_18180);
or U19299 (N_19299,N_18115,N_18204);
nand U19300 (N_19300,N_18979,N_18775);
and U19301 (N_19301,N_18053,N_18611);
or U19302 (N_19302,N_18874,N_18267);
nor U19303 (N_19303,N_18638,N_18105);
or U19304 (N_19304,N_18976,N_18912);
and U19305 (N_19305,N_18517,N_18848);
nor U19306 (N_19306,N_18214,N_18550);
nand U19307 (N_19307,N_18232,N_18977);
xor U19308 (N_19308,N_18055,N_18120);
nand U19309 (N_19309,N_18785,N_18447);
nor U19310 (N_19310,N_18021,N_18835);
and U19311 (N_19311,N_18248,N_18259);
nor U19312 (N_19312,N_18137,N_18888);
or U19313 (N_19313,N_18881,N_18191);
xnor U19314 (N_19314,N_18606,N_18272);
nor U19315 (N_19315,N_18745,N_18108);
or U19316 (N_19316,N_18557,N_18819);
or U19317 (N_19317,N_18783,N_18068);
nor U19318 (N_19318,N_18551,N_18221);
and U19319 (N_19319,N_18537,N_18520);
nor U19320 (N_19320,N_18758,N_18891);
nand U19321 (N_19321,N_18439,N_18346);
and U19322 (N_19322,N_18506,N_18563);
or U19323 (N_19323,N_18514,N_18949);
or U19324 (N_19324,N_18077,N_18406);
nand U19325 (N_19325,N_18531,N_18699);
nor U19326 (N_19326,N_18963,N_18713);
nand U19327 (N_19327,N_18106,N_18987);
or U19328 (N_19328,N_18425,N_18408);
nor U19329 (N_19329,N_18103,N_18730);
nand U19330 (N_19330,N_18572,N_18755);
nand U19331 (N_19331,N_18632,N_18150);
or U19332 (N_19332,N_18883,N_18681);
and U19333 (N_19333,N_18588,N_18861);
nor U19334 (N_19334,N_18625,N_18241);
nor U19335 (N_19335,N_18768,N_18789);
or U19336 (N_19336,N_18252,N_18837);
and U19337 (N_19337,N_18801,N_18430);
nand U19338 (N_19338,N_18938,N_18973);
nor U19339 (N_19339,N_18422,N_18982);
or U19340 (N_19340,N_18741,N_18419);
nor U19341 (N_19341,N_18145,N_18046);
or U19342 (N_19342,N_18538,N_18841);
and U19343 (N_19343,N_18080,N_18061);
nand U19344 (N_19344,N_18863,N_18872);
and U19345 (N_19345,N_18010,N_18894);
nand U19346 (N_19346,N_18509,N_18113);
xor U19347 (N_19347,N_18119,N_18665);
and U19348 (N_19348,N_18296,N_18347);
and U19349 (N_19349,N_18542,N_18240);
or U19350 (N_19350,N_18655,N_18978);
nand U19351 (N_19351,N_18946,N_18467);
and U19352 (N_19352,N_18802,N_18540);
xnor U19353 (N_19353,N_18049,N_18541);
nand U19354 (N_19354,N_18385,N_18188);
nand U19355 (N_19355,N_18525,N_18905);
or U19356 (N_19356,N_18597,N_18031);
nand U19357 (N_19357,N_18415,N_18628);
xnor U19358 (N_19358,N_18436,N_18463);
or U19359 (N_19359,N_18166,N_18117);
and U19360 (N_19360,N_18206,N_18101);
nor U19361 (N_19361,N_18751,N_18216);
or U19362 (N_19362,N_18651,N_18187);
nand U19363 (N_19363,N_18096,N_18139);
or U19364 (N_19364,N_18159,N_18777);
nand U19365 (N_19365,N_18489,N_18828);
nand U19366 (N_19366,N_18917,N_18417);
and U19367 (N_19367,N_18445,N_18865);
nor U19368 (N_19368,N_18156,N_18689);
nand U19369 (N_19369,N_18764,N_18701);
nand U19370 (N_19370,N_18086,N_18724);
nor U19371 (N_19371,N_18128,N_18292);
nor U19372 (N_19372,N_18057,N_18205);
nand U19373 (N_19373,N_18711,N_18807);
or U19374 (N_19374,N_18432,N_18663);
nor U19375 (N_19375,N_18851,N_18433);
nand U19376 (N_19376,N_18334,N_18440);
or U19377 (N_19377,N_18587,N_18424);
nand U19378 (N_19378,N_18753,N_18363);
or U19379 (N_19379,N_18153,N_18400);
or U19380 (N_19380,N_18619,N_18989);
and U19381 (N_19381,N_18999,N_18513);
and U19382 (N_19382,N_18954,N_18626);
and U19383 (N_19383,N_18181,N_18685);
or U19384 (N_19384,N_18320,N_18907);
nand U19385 (N_19385,N_18903,N_18504);
or U19386 (N_19386,N_18063,N_18093);
nand U19387 (N_19387,N_18325,N_18466);
nor U19388 (N_19388,N_18732,N_18869);
or U19389 (N_19389,N_18833,N_18018);
xnor U19390 (N_19390,N_18950,N_18472);
or U19391 (N_19391,N_18193,N_18020);
and U19392 (N_19392,N_18684,N_18157);
nor U19393 (N_19393,N_18162,N_18575);
and U19394 (N_19394,N_18338,N_18079);
or U19395 (N_19395,N_18871,N_18459);
or U19396 (N_19396,N_18997,N_18015);
nor U19397 (N_19397,N_18276,N_18034);
nand U19398 (N_19398,N_18660,N_18493);
or U19399 (N_19399,N_18761,N_18378);
nand U19400 (N_19400,N_18475,N_18669);
nor U19401 (N_19401,N_18027,N_18089);
and U19402 (N_19402,N_18107,N_18343);
xor U19403 (N_19403,N_18460,N_18211);
and U19404 (N_19404,N_18403,N_18359);
nand U19405 (N_19405,N_18277,N_18608);
and U19406 (N_19406,N_18640,N_18412);
or U19407 (N_19407,N_18812,N_18956);
or U19408 (N_19408,N_18580,N_18185);
nor U19409 (N_19409,N_18609,N_18274);
or U19410 (N_19410,N_18998,N_18407);
and U19411 (N_19411,N_18613,N_18867);
or U19412 (N_19412,N_18356,N_18945);
nand U19413 (N_19413,N_18576,N_18431);
nand U19414 (N_19414,N_18521,N_18951);
or U19415 (N_19415,N_18719,N_18864);
or U19416 (N_19416,N_18143,N_18714);
nor U19417 (N_19417,N_18498,N_18458);
or U19418 (N_19418,N_18667,N_18494);
and U19419 (N_19419,N_18726,N_18085);
nor U19420 (N_19420,N_18488,N_18754);
and U19421 (N_19421,N_18286,N_18718);
nor U19422 (N_19422,N_18716,N_18725);
or U19423 (N_19423,N_18672,N_18526);
nor U19424 (N_19424,N_18152,N_18943);
or U19425 (N_19425,N_18001,N_18486);
or U19426 (N_19426,N_18709,N_18052);
and U19427 (N_19427,N_18380,N_18025);
nand U19428 (N_19428,N_18855,N_18226);
or U19429 (N_19429,N_18282,N_18935);
nor U19430 (N_19430,N_18787,N_18333);
xor U19431 (N_19431,N_18627,N_18862);
nor U19432 (N_19432,N_18307,N_18330);
nor U19433 (N_19433,N_18924,N_18235);
or U19434 (N_19434,N_18921,N_18367);
and U19435 (N_19435,N_18365,N_18739);
nand U19436 (N_19436,N_18836,N_18710);
nor U19437 (N_19437,N_18975,N_18448);
xnor U19438 (N_19438,N_18016,N_18039);
and U19439 (N_19439,N_18084,N_18727);
nor U19440 (N_19440,N_18327,N_18742);
and U19441 (N_19441,N_18931,N_18897);
and U19442 (N_19442,N_18289,N_18650);
nor U19443 (N_19443,N_18664,N_18484);
or U19444 (N_19444,N_18778,N_18300);
nand U19445 (N_19445,N_18501,N_18304);
or U19446 (N_19446,N_18414,N_18734);
nor U19447 (N_19447,N_18177,N_18876);
nand U19448 (N_19448,N_18416,N_18176);
nor U19449 (N_19449,N_18702,N_18916);
and U19450 (N_19450,N_18510,N_18941);
and U19451 (N_19451,N_18523,N_18321);
nor U19452 (N_19452,N_18004,N_18875);
or U19453 (N_19453,N_18889,N_18642);
nand U19454 (N_19454,N_18960,N_18566);
nand U19455 (N_19455,N_18402,N_18337);
and U19456 (N_19456,N_18738,N_18478);
nor U19457 (N_19457,N_18633,N_18349);
nor U19458 (N_19458,N_18258,N_18744);
or U19459 (N_19459,N_18306,N_18762);
or U19460 (N_19460,N_18548,N_18934);
nor U19461 (N_19461,N_18919,N_18154);
nor U19462 (N_19462,N_18571,N_18900);
or U19463 (N_19463,N_18290,N_18671);
nor U19464 (N_19464,N_18104,N_18827);
xor U19465 (N_19465,N_18972,N_18729);
or U19466 (N_19466,N_18657,N_18473);
nor U19467 (N_19467,N_18287,N_18026);
or U19468 (N_19468,N_18731,N_18560);
and U19469 (N_19469,N_18418,N_18192);
nand U19470 (N_19470,N_18549,N_18659);
or U19471 (N_19471,N_18397,N_18899);
nor U19472 (N_19472,N_18404,N_18174);
nand U19473 (N_19473,N_18111,N_18516);
nor U19474 (N_19474,N_18160,N_18503);
and U19475 (N_19475,N_18266,N_18937);
xnor U19476 (N_19476,N_18208,N_18539);
and U19477 (N_19477,N_18375,N_18471);
or U19478 (N_19478,N_18674,N_18771);
or U19479 (N_19479,N_18391,N_18234);
xnor U19480 (N_19480,N_18620,N_18446);
or U19481 (N_19481,N_18794,N_18371);
and U19482 (N_19482,N_18353,N_18634);
or U19483 (N_19483,N_18364,N_18133);
nand U19484 (N_19484,N_18678,N_18443);
nor U19485 (N_19485,N_18639,N_18399);
nand U19486 (N_19486,N_18770,N_18736);
or U19487 (N_19487,N_18969,N_18929);
or U19488 (N_19488,N_18250,N_18442);
nand U19489 (N_19489,N_18822,N_18410);
nor U19490 (N_19490,N_18569,N_18859);
nand U19491 (N_19491,N_18072,N_18100);
nor U19492 (N_19492,N_18254,N_18255);
nor U19493 (N_19493,N_18834,N_18045);
nor U19494 (N_19494,N_18809,N_18518);
and U19495 (N_19495,N_18310,N_18940);
nand U19496 (N_19496,N_18132,N_18676);
nand U19497 (N_19497,N_18911,N_18023);
and U19498 (N_19498,N_18845,N_18019);
nand U19499 (N_19499,N_18066,N_18984);
or U19500 (N_19500,N_18931,N_18368);
nor U19501 (N_19501,N_18947,N_18647);
nor U19502 (N_19502,N_18928,N_18718);
or U19503 (N_19503,N_18675,N_18691);
and U19504 (N_19504,N_18643,N_18871);
nand U19505 (N_19505,N_18992,N_18092);
nand U19506 (N_19506,N_18472,N_18616);
nor U19507 (N_19507,N_18981,N_18965);
xnor U19508 (N_19508,N_18790,N_18157);
or U19509 (N_19509,N_18175,N_18533);
nor U19510 (N_19510,N_18082,N_18498);
and U19511 (N_19511,N_18887,N_18800);
nor U19512 (N_19512,N_18133,N_18979);
nor U19513 (N_19513,N_18386,N_18182);
xnor U19514 (N_19514,N_18511,N_18137);
and U19515 (N_19515,N_18587,N_18175);
and U19516 (N_19516,N_18218,N_18260);
or U19517 (N_19517,N_18590,N_18402);
nor U19518 (N_19518,N_18989,N_18002);
nor U19519 (N_19519,N_18056,N_18283);
xor U19520 (N_19520,N_18382,N_18610);
or U19521 (N_19521,N_18796,N_18975);
nand U19522 (N_19522,N_18964,N_18322);
nand U19523 (N_19523,N_18422,N_18417);
nand U19524 (N_19524,N_18479,N_18322);
or U19525 (N_19525,N_18524,N_18833);
nand U19526 (N_19526,N_18413,N_18151);
and U19527 (N_19527,N_18136,N_18825);
nor U19528 (N_19528,N_18668,N_18610);
nand U19529 (N_19529,N_18133,N_18811);
or U19530 (N_19530,N_18715,N_18056);
nor U19531 (N_19531,N_18423,N_18756);
and U19532 (N_19532,N_18606,N_18520);
and U19533 (N_19533,N_18592,N_18295);
nor U19534 (N_19534,N_18260,N_18597);
nor U19535 (N_19535,N_18510,N_18361);
xor U19536 (N_19536,N_18355,N_18123);
nand U19537 (N_19537,N_18861,N_18198);
nand U19538 (N_19538,N_18420,N_18826);
nor U19539 (N_19539,N_18261,N_18112);
or U19540 (N_19540,N_18164,N_18243);
nand U19541 (N_19541,N_18262,N_18085);
or U19542 (N_19542,N_18472,N_18203);
xnor U19543 (N_19543,N_18748,N_18690);
and U19544 (N_19544,N_18759,N_18373);
xor U19545 (N_19545,N_18807,N_18873);
and U19546 (N_19546,N_18571,N_18657);
or U19547 (N_19547,N_18597,N_18396);
or U19548 (N_19548,N_18721,N_18844);
nand U19549 (N_19549,N_18620,N_18754);
xor U19550 (N_19550,N_18138,N_18927);
nand U19551 (N_19551,N_18048,N_18746);
and U19552 (N_19552,N_18235,N_18555);
nand U19553 (N_19553,N_18764,N_18920);
nor U19554 (N_19554,N_18953,N_18325);
nor U19555 (N_19555,N_18374,N_18669);
nand U19556 (N_19556,N_18027,N_18951);
nand U19557 (N_19557,N_18447,N_18000);
nor U19558 (N_19558,N_18755,N_18167);
and U19559 (N_19559,N_18051,N_18993);
nor U19560 (N_19560,N_18312,N_18790);
xor U19561 (N_19561,N_18568,N_18975);
or U19562 (N_19562,N_18208,N_18832);
and U19563 (N_19563,N_18370,N_18917);
and U19564 (N_19564,N_18131,N_18016);
nor U19565 (N_19565,N_18628,N_18181);
or U19566 (N_19566,N_18236,N_18608);
xor U19567 (N_19567,N_18415,N_18730);
and U19568 (N_19568,N_18722,N_18909);
nand U19569 (N_19569,N_18623,N_18653);
nand U19570 (N_19570,N_18107,N_18788);
nor U19571 (N_19571,N_18091,N_18913);
and U19572 (N_19572,N_18452,N_18900);
nand U19573 (N_19573,N_18358,N_18441);
nor U19574 (N_19574,N_18034,N_18535);
nand U19575 (N_19575,N_18796,N_18977);
or U19576 (N_19576,N_18116,N_18600);
or U19577 (N_19577,N_18494,N_18174);
and U19578 (N_19578,N_18941,N_18036);
nand U19579 (N_19579,N_18892,N_18721);
or U19580 (N_19580,N_18702,N_18402);
nand U19581 (N_19581,N_18517,N_18042);
nand U19582 (N_19582,N_18840,N_18362);
xor U19583 (N_19583,N_18295,N_18586);
xor U19584 (N_19584,N_18367,N_18914);
xor U19585 (N_19585,N_18036,N_18836);
and U19586 (N_19586,N_18346,N_18373);
and U19587 (N_19587,N_18010,N_18582);
and U19588 (N_19588,N_18658,N_18096);
and U19589 (N_19589,N_18587,N_18295);
nand U19590 (N_19590,N_18978,N_18016);
nand U19591 (N_19591,N_18602,N_18768);
and U19592 (N_19592,N_18851,N_18316);
or U19593 (N_19593,N_18023,N_18216);
nand U19594 (N_19594,N_18108,N_18648);
nand U19595 (N_19595,N_18558,N_18770);
nor U19596 (N_19596,N_18854,N_18109);
and U19597 (N_19597,N_18186,N_18003);
and U19598 (N_19598,N_18344,N_18155);
nand U19599 (N_19599,N_18622,N_18944);
or U19600 (N_19600,N_18804,N_18842);
and U19601 (N_19601,N_18544,N_18939);
or U19602 (N_19602,N_18908,N_18975);
or U19603 (N_19603,N_18049,N_18477);
nor U19604 (N_19604,N_18247,N_18146);
or U19605 (N_19605,N_18385,N_18659);
or U19606 (N_19606,N_18267,N_18987);
xnor U19607 (N_19607,N_18705,N_18775);
nor U19608 (N_19608,N_18448,N_18810);
or U19609 (N_19609,N_18048,N_18321);
or U19610 (N_19610,N_18730,N_18298);
and U19611 (N_19611,N_18890,N_18387);
or U19612 (N_19612,N_18968,N_18565);
or U19613 (N_19613,N_18671,N_18362);
and U19614 (N_19614,N_18216,N_18729);
and U19615 (N_19615,N_18890,N_18778);
nor U19616 (N_19616,N_18377,N_18295);
and U19617 (N_19617,N_18976,N_18460);
nand U19618 (N_19618,N_18608,N_18359);
or U19619 (N_19619,N_18528,N_18481);
or U19620 (N_19620,N_18087,N_18046);
and U19621 (N_19621,N_18034,N_18043);
and U19622 (N_19622,N_18018,N_18982);
and U19623 (N_19623,N_18895,N_18990);
and U19624 (N_19624,N_18369,N_18979);
and U19625 (N_19625,N_18128,N_18322);
and U19626 (N_19626,N_18292,N_18131);
nand U19627 (N_19627,N_18311,N_18648);
nand U19628 (N_19628,N_18425,N_18068);
nand U19629 (N_19629,N_18105,N_18906);
and U19630 (N_19630,N_18891,N_18166);
nor U19631 (N_19631,N_18837,N_18278);
nand U19632 (N_19632,N_18456,N_18810);
nand U19633 (N_19633,N_18432,N_18856);
or U19634 (N_19634,N_18219,N_18786);
nor U19635 (N_19635,N_18081,N_18192);
or U19636 (N_19636,N_18593,N_18326);
nand U19637 (N_19637,N_18765,N_18152);
xor U19638 (N_19638,N_18668,N_18966);
and U19639 (N_19639,N_18742,N_18534);
nand U19640 (N_19640,N_18271,N_18495);
nor U19641 (N_19641,N_18466,N_18411);
nor U19642 (N_19642,N_18926,N_18929);
nor U19643 (N_19643,N_18897,N_18899);
and U19644 (N_19644,N_18913,N_18598);
nand U19645 (N_19645,N_18209,N_18003);
nand U19646 (N_19646,N_18832,N_18260);
and U19647 (N_19647,N_18622,N_18008);
xnor U19648 (N_19648,N_18890,N_18040);
and U19649 (N_19649,N_18104,N_18149);
nand U19650 (N_19650,N_18903,N_18585);
nand U19651 (N_19651,N_18637,N_18873);
nand U19652 (N_19652,N_18743,N_18471);
or U19653 (N_19653,N_18593,N_18889);
xor U19654 (N_19654,N_18347,N_18571);
nor U19655 (N_19655,N_18459,N_18682);
nand U19656 (N_19656,N_18463,N_18053);
nand U19657 (N_19657,N_18034,N_18200);
or U19658 (N_19658,N_18673,N_18168);
nor U19659 (N_19659,N_18050,N_18245);
and U19660 (N_19660,N_18049,N_18660);
and U19661 (N_19661,N_18588,N_18862);
or U19662 (N_19662,N_18771,N_18490);
or U19663 (N_19663,N_18369,N_18388);
xor U19664 (N_19664,N_18419,N_18416);
nand U19665 (N_19665,N_18319,N_18524);
nand U19666 (N_19666,N_18767,N_18649);
or U19667 (N_19667,N_18277,N_18476);
xnor U19668 (N_19668,N_18492,N_18923);
xnor U19669 (N_19669,N_18955,N_18963);
nand U19670 (N_19670,N_18473,N_18502);
nand U19671 (N_19671,N_18530,N_18570);
nor U19672 (N_19672,N_18997,N_18360);
nand U19673 (N_19673,N_18111,N_18250);
xnor U19674 (N_19674,N_18811,N_18962);
or U19675 (N_19675,N_18085,N_18235);
or U19676 (N_19676,N_18407,N_18262);
or U19677 (N_19677,N_18354,N_18897);
xor U19678 (N_19678,N_18224,N_18790);
or U19679 (N_19679,N_18432,N_18387);
nor U19680 (N_19680,N_18507,N_18750);
and U19681 (N_19681,N_18784,N_18913);
or U19682 (N_19682,N_18003,N_18318);
or U19683 (N_19683,N_18741,N_18912);
nor U19684 (N_19684,N_18084,N_18287);
nand U19685 (N_19685,N_18225,N_18426);
nand U19686 (N_19686,N_18324,N_18829);
or U19687 (N_19687,N_18220,N_18893);
xnor U19688 (N_19688,N_18006,N_18924);
nor U19689 (N_19689,N_18950,N_18353);
nor U19690 (N_19690,N_18663,N_18067);
nand U19691 (N_19691,N_18368,N_18828);
xnor U19692 (N_19692,N_18701,N_18952);
and U19693 (N_19693,N_18665,N_18002);
nand U19694 (N_19694,N_18122,N_18293);
nand U19695 (N_19695,N_18323,N_18735);
and U19696 (N_19696,N_18747,N_18877);
nand U19697 (N_19697,N_18722,N_18604);
or U19698 (N_19698,N_18185,N_18547);
and U19699 (N_19699,N_18161,N_18246);
nor U19700 (N_19700,N_18352,N_18091);
or U19701 (N_19701,N_18725,N_18387);
or U19702 (N_19702,N_18885,N_18067);
nor U19703 (N_19703,N_18101,N_18172);
or U19704 (N_19704,N_18941,N_18411);
nand U19705 (N_19705,N_18023,N_18942);
nand U19706 (N_19706,N_18314,N_18157);
and U19707 (N_19707,N_18348,N_18726);
nor U19708 (N_19708,N_18636,N_18390);
or U19709 (N_19709,N_18760,N_18356);
and U19710 (N_19710,N_18507,N_18939);
nand U19711 (N_19711,N_18899,N_18339);
or U19712 (N_19712,N_18328,N_18794);
nand U19713 (N_19713,N_18403,N_18829);
and U19714 (N_19714,N_18924,N_18539);
nand U19715 (N_19715,N_18050,N_18530);
and U19716 (N_19716,N_18759,N_18935);
nand U19717 (N_19717,N_18371,N_18144);
or U19718 (N_19718,N_18317,N_18083);
and U19719 (N_19719,N_18000,N_18830);
xor U19720 (N_19720,N_18147,N_18756);
nor U19721 (N_19721,N_18817,N_18407);
or U19722 (N_19722,N_18105,N_18085);
xor U19723 (N_19723,N_18887,N_18828);
nor U19724 (N_19724,N_18518,N_18301);
nand U19725 (N_19725,N_18666,N_18271);
or U19726 (N_19726,N_18298,N_18683);
nor U19727 (N_19727,N_18784,N_18127);
nand U19728 (N_19728,N_18114,N_18426);
xnor U19729 (N_19729,N_18362,N_18031);
nand U19730 (N_19730,N_18767,N_18523);
or U19731 (N_19731,N_18202,N_18965);
nor U19732 (N_19732,N_18843,N_18972);
or U19733 (N_19733,N_18281,N_18663);
or U19734 (N_19734,N_18171,N_18380);
and U19735 (N_19735,N_18782,N_18206);
or U19736 (N_19736,N_18518,N_18899);
or U19737 (N_19737,N_18418,N_18638);
nand U19738 (N_19738,N_18604,N_18451);
nor U19739 (N_19739,N_18549,N_18115);
nand U19740 (N_19740,N_18979,N_18859);
nand U19741 (N_19741,N_18209,N_18064);
nand U19742 (N_19742,N_18586,N_18929);
nor U19743 (N_19743,N_18995,N_18085);
nand U19744 (N_19744,N_18668,N_18848);
and U19745 (N_19745,N_18288,N_18162);
or U19746 (N_19746,N_18017,N_18482);
and U19747 (N_19747,N_18205,N_18214);
nor U19748 (N_19748,N_18723,N_18514);
and U19749 (N_19749,N_18944,N_18015);
nand U19750 (N_19750,N_18901,N_18431);
nand U19751 (N_19751,N_18937,N_18949);
xnor U19752 (N_19752,N_18697,N_18588);
and U19753 (N_19753,N_18826,N_18567);
nor U19754 (N_19754,N_18019,N_18302);
nand U19755 (N_19755,N_18720,N_18804);
nand U19756 (N_19756,N_18504,N_18737);
nand U19757 (N_19757,N_18985,N_18664);
xor U19758 (N_19758,N_18567,N_18787);
and U19759 (N_19759,N_18313,N_18673);
nor U19760 (N_19760,N_18683,N_18387);
nor U19761 (N_19761,N_18845,N_18330);
and U19762 (N_19762,N_18131,N_18938);
nor U19763 (N_19763,N_18728,N_18548);
or U19764 (N_19764,N_18520,N_18848);
and U19765 (N_19765,N_18020,N_18699);
nand U19766 (N_19766,N_18894,N_18130);
and U19767 (N_19767,N_18717,N_18150);
or U19768 (N_19768,N_18828,N_18824);
nand U19769 (N_19769,N_18472,N_18627);
nand U19770 (N_19770,N_18321,N_18543);
nor U19771 (N_19771,N_18433,N_18421);
xor U19772 (N_19772,N_18310,N_18390);
or U19773 (N_19773,N_18608,N_18561);
or U19774 (N_19774,N_18650,N_18772);
or U19775 (N_19775,N_18813,N_18867);
nor U19776 (N_19776,N_18560,N_18540);
nand U19777 (N_19777,N_18280,N_18435);
and U19778 (N_19778,N_18938,N_18805);
nor U19779 (N_19779,N_18922,N_18681);
nand U19780 (N_19780,N_18449,N_18982);
nor U19781 (N_19781,N_18939,N_18128);
or U19782 (N_19782,N_18612,N_18873);
or U19783 (N_19783,N_18912,N_18339);
and U19784 (N_19784,N_18888,N_18770);
nand U19785 (N_19785,N_18374,N_18476);
or U19786 (N_19786,N_18540,N_18857);
or U19787 (N_19787,N_18914,N_18570);
and U19788 (N_19788,N_18675,N_18410);
nand U19789 (N_19789,N_18560,N_18401);
xor U19790 (N_19790,N_18342,N_18437);
or U19791 (N_19791,N_18423,N_18654);
and U19792 (N_19792,N_18806,N_18731);
and U19793 (N_19793,N_18666,N_18019);
nand U19794 (N_19794,N_18178,N_18707);
and U19795 (N_19795,N_18133,N_18895);
or U19796 (N_19796,N_18655,N_18053);
and U19797 (N_19797,N_18976,N_18969);
nor U19798 (N_19798,N_18493,N_18212);
or U19799 (N_19799,N_18862,N_18060);
nand U19800 (N_19800,N_18802,N_18590);
nor U19801 (N_19801,N_18129,N_18261);
nand U19802 (N_19802,N_18806,N_18242);
or U19803 (N_19803,N_18339,N_18123);
nand U19804 (N_19804,N_18425,N_18718);
nand U19805 (N_19805,N_18677,N_18713);
and U19806 (N_19806,N_18351,N_18449);
and U19807 (N_19807,N_18929,N_18542);
or U19808 (N_19808,N_18255,N_18297);
and U19809 (N_19809,N_18982,N_18170);
and U19810 (N_19810,N_18164,N_18839);
or U19811 (N_19811,N_18701,N_18101);
and U19812 (N_19812,N_18041,N_18974);
nor U19813 (N_19813,N_18845,N_18593);
nor U19814 (N_19814,N_18321,N_18732);
and U19815 (N_19815,N_18214,N_18841);
or U19816 (N_19816,N_18016,N_18748);
nor U19817 (N_19817,N_18226,N_18206);
or U19818 (N_19818,N_18213,N_18544);
or U19819 (N_19819,N_18802,N_18297);
or U19820 (N_19820,N_18699,N_18755);
nand U19821 (N_19821,N_18914,N_18927);
nand U19822 (N_19822,N_18827,N_18999);
and U19823 (N_19823,N_18247,N_18267);
or U19824 (N_19824,N_18488,N_18923);
nand U19825 (N_19825,N_18299,N_18884);
xor U19826 (N_19826,N_18162,N_18336);
nand U19827 (N_19827,N_18371,N_18159);
and U19828 (N_19828,N_18237,N_18018);
xor U19829 (N_19829,N_18965,N_18030);
xnor U19830 (N_19830,N_18699,N_18156);
nor U19831 (N_19831,N_18269,N_18869);
nand U19832 (N_19832,N_18332,N_18961);
and U19833 (N_19833,N_18751,N_18383);
or U19834 (N_19834,N_18218,N_18180);
and U19835 (N_19835,N_18143,N_18996);
or U19836 (N_19836,N_18630,N_18600);
nand U19837 (N_19837,N_18911,N_18575);
and U19838 (N_19838,N_18170,N_18929);
and U19839 (N_19839,N_18228,N_18257);
nor U19840 (N_19840,N_18793,N_18339);
nor U19841 (N_19841,N_18005,N_18897);
nand U19842 (N_19842,N_18745,N_18934);
and U19843 (N_19843,N_18377,N_18288);
nor U19844 (N_19844,N_18145,N_18835);
and U19845 (N_19845,N_18286,N_18823);
and U19846 (N_19846,N_18092,N_18650);
or U19847 (N_19847,N_18163,N_18912);
and U19848 (N_19848,N_18134,N_18551);
nor U19849 (N_19849,N_18051,N_18828);
or U19850 (N_19850,N_18062,N_18637);
nor U19851 (N_19851,N_18144,N_18158);
nand U19852 (N_19852,N_18786,N_18762);
nand U19853 (N_19853,N_18576,N_18699);
xnor U19854 (N_19854,N_18814,N_18884);
or U19855 (N_19855,N_18424,N_18900);
and U19856 (N_19856,N_18791,N_18310);
and U19857 (N_19857,N_18674,N_18853);
or U19858 (N_19858,N_18128,N_18194);
nand U19859 (N_19859,N_18372,N_18517);
nand U19860 (N_19860,N_18221,N_18696);
nor U19861 (N_19861,N_18119,N_18635);
or U19862 (N_19862,N_18653,N_18768);
nor U19863 (N_19863,N_18173,N_18462);
or U19864 (N_19864,N_18677,N_18037);
xnor U19865 (N_19865,N_18146,N_18765);
and U19866 (N_19866,N_18589,N_18918);
and U19867 (N_19867,N_18094,N_18777);
nor U19868 (N_19868,N_18346,N_18248);
and U19869 (N_19869,N_18716,N_18630);
nand U19870 (N_19870,N_18991,N_18198);
or U19871 (N_19871,N_18687,N_18826);
nand U19872 (N_19872,N_18176,N_18060);
nand U19873 (N_19873,N_18851,N_18551);
nand U19874 (N_19874,N_18264,N_18620);
nand U19875 (N_19875,N_18373,N_18476);
or U19876 (N_19876,N_18786,N_18883);
and U19877 (N_19877,N_18068,N_18177);
or U19878 (N_19878,N_18240,N_18865);
or U19879 (N_19879,N_18104,N_18728);
nor U19880 (N_19880,N_18825,N_18562);
nand U19881 (N_19881,N_18272,N_18548);
and U19882 (N_19882,N_18367,N_18916);
or U19883 (N_19883,N_18227,N_18885);
and U19884 (N_19884,N_18653,N_18617);
nor U19885 (N_19885,N_18245,N_18274);
nand U19886 (N_19886,N_18350,N_18672);
nand U19887 (N_19887,N_18762,N_18337);
nand U19888 (N_19888,N_18285,N_18106);
nor U19889 (N_19889,N_18990,N_18025);
nand U19890 (N_19890,N_18612,N_18215);
nor U19891 (N_19891,N_18105,N_18587);
nor U19892 (N_19892,N_18748,N_18977);
and U19893 (N_19893,N_18374,N_18229);
nand U19894 (N_19894,N_18125,N_18615);
or U19895 (N_19895,N_18968,N_18661);
nand U19896 (N_19896,N_18522,N_18009);
and U19897 (N_19897,N_18731,N_18516);
nor U19898 (N_19898,N_18967,N_18391);
and U19899 (N_19899,N_18493,N_18983);
and U19900 (N_19900,N_18218,N_18757);
nand U19901 (N_19901,N_18850,N_18708);
or U19902 (N_19902,N_18078,N_18726);
and U19903 (N_19903,N_18999,N_18437);
nand U19904 (N_19904,N_18779,N_18409);
or U19905 (N_19905,N_18340,N_18787);
nor U19906 (N_19906,N_18293,N_18377);
nand U19907 (N_19907,N_18129,N_18920);
nand U19908 (N_19908,N_18443,N_18882);
nor U19909 (N_19909,N_18285,N_18714);
nand U19910 (N_19910,N_18412,N_18924);
nand U19911 (N_19911,N_18870,N_18490);
and U19912 (N_19912,N_18207,N_18536);
and U19913 (N_19913,N_18286,N_18292);
nand U19914 (N_19914,N_18154,N_18242);
or U19915 (N_19915,N_18687,N_18914);
and U19916 (N_19916,N_18486,N_18085);
or U19917 (N_19917,N_18620,N_18330);
nor U19918 (N_19918,N_18001,N_18757);
or U19919 (N_19919,N_18994,N_18319);
xor U19920 (N_19920,N_18924,N_18219);
xor U19921 (N_19921,N_18331,N_18944);
and U19922 (N_19922,N_18760,N_18189);
or U19923 (N_19923,N_18964,N_18464);
or U19924 (N_19924,N_18612,N_18022);
or U19925 (N_19925,N_18063,N_18982);
or U19926 (N_19926,N_18414,N_18425);
and U19927 (N_19927,N_18108,N_18567);
nor U19928 (N_19928,N_18550,N_18543);
xor U19929 (N_19929,N_18152,N_18738);
nor U19930 (N_19930,N_18668,N_18662);
nand U19931 (N_19931,N_18311,N_18907);
xor U19932 (N_19932,N_18871,N_18439);
and U19933 (N_19933,N_18013,N_18631);
and U19934 (N_19934,N_18149,N_18337);
and U19935 (N_19935,N_18797,N_18310);
and U19936 (N_19936,N_18422,N_18078);
xnor U19937 (N_19937,N_18956,N_18198);
xnor U19938 (N_19938,N_18657,N_18849);
or U19939 (N_19939,N_18427,N_18181);
or U19940 (N_19940,N_18208,N_18859);
and U19941 (N_19941,N_18934,N_18434);
xnor U19942 (N_19942,N_18505,N_18887);
or U19943 (N_19943,N_18816,N_18714);
nor U19944 (N_19944,N_18103,N_18450);
or U19945 (N_19945,N_18777,N_18125);
nor U19946 (N_19946,N_18853,N_18378);
and U19947 (N_19947,N_18073,N_18215);
and U19948 (N_19948,N_18139,N_18289);
xnor U19949 (N_19949,N_18078,N_18121);
or U19950 (N_19950,N_18340,N_18440);
nand U19951 (N_19951,N_18818,N_18689);
nand U19952 (N_19952,N_18696,N_18916);
nand U19953 (N_19953,N_18627,N_18201);
nor U19954 (N_19954,N_18406,N_18391);
nor U19955 (N_19955,N_18813,N_18192);
nor U19956 (N_19956,N_18284,N_18001);
nand U19957 (N_19957,N_18861,N_18731);
or U19958 (N_19958,N_18152,N_18365);
nor U19959 (N_19959,N_18750,N_18528);
or U19960 (N_19960,N_18201,N_18939);
nand U19961 (N_19961,N_18876,N_18207);
nor U19962 (N_19962,N_18632,N_18688);
nand U19963 (N_19963,N_18921,N_18790);
or U19964 (N_19964,N_18654,N_18114);
or U19965 (N_19965,N_18103,N_18868);
nor U19966 (N_19966,N_18705,N_18211);
nand U19967 (N_19967,N_18313,N_18687);
nor U19968 (N_19968,N_18797,N_18500);
nand U19969 (N_19969,N_18708,N_18011);
and U19970 (N_19970,N_18515,N_18165);
nor U19971 (N_19971,N_18069,N_18736);
or U19972 (N_19972,N_18220,N_18109);
xor U19973 (N_19973,N_18720,N_18457);
nand U19974 (N_19974,N_18571,N_18659);
and U19975 (N_19975,N_18533,N_18508);
nand U19976 (N_19976,N_18699,N_18509);
nor U19977 (N_19977,N_18435,N_18124);
nor U19978 (N_19978,N_18879,N_18878);
nand U19979 (N_19979,N_18758,N_18353);
or U19980 (N_19980,N_18042,N_18282);
or U19981 (N_19981,N_18655,N_18767);
or U19982 (N_19982,N_18900,N_18559);
and U19983 (N_19983,N_18643,N_18037);
and U19984 (N_19984,N_18481,N_18304);
nand U19985 (N_19985,N_18579,N_18710);
or U19986 (N_19986,N_18646,N_18715);
xor U19987 (N_19987,N_18796,N_18844);
nor U19988 (N_19988,N_18842,N_18682);
nor U19989 (N_19989,N_18666,N_18989);
nand U19990 (N_19990,N_18522,N_18841);
or U19991 (N_19991,N_18549,N_18401);
nand U19992 (N_19992,N_18769,N_18433);
xnor U19993 (N_19993,N_18703,N_18196);
and U19994 (N_19994,N_18830,N_18930);
and U19995 (N_19995,N_18372,N_18089);
and U19996 (N_19996,N_18561,N_18751);
nor U19997 (N_19997,N_18413,N_18522);
nand U19998 (N_19998,N_18548,N_18652);
and U19999 (N_19999,N_18533,N_18380);
or UO_0 (O_0,N_19978,N_19621);
or UO_1 (O_1,N_19710,N_19331);
and UO_2 (O_2,N_19376,N_19823);
or UO_3 (O_3,N_19240,N_19944);
xor UO_4 (O_4,N_19193,N_19887);
nor UO_5 (O_5,N_19706,N_19549);
nand UO_6 (O_6,N_19624,N_19210);
xnor UO_7 (O_7,N_19440,N_19363);
nor UO_8 (O_8,N_19943,N_19081);
nor UO_9 (O_9,N_19687,N_19370);
xor UO_10 (O_10,N_19326,N_19134);
nand UO_11 (O_11,N_19428,N_19760);
nand UO_12 (O_12,N_19358,N_19026);
nand UO_13 (O_13,N_19521,N_19028);
xnor UO_14 (O_14,N_19939,N_19762);
and UO_15 (O_15,N_19531,N_19498);
and UO_16 (O_16,N_19647,N_19133);
or UO_17 (O_17,N_19861,N_19115);
or UO_18 (O_18,N_19786,N_19323);
nand UO_19 (O_19,N_19812,N_19962);
or UO_20 (O_20,N_19073,N_19538);
nor UO_21 (O_21,N_19524,N_19041);
nand UO_22 (O_22,N_19622,N_19456);
xnor UO_23 (O_23,N_19930,N_19686);
nor UO_24 (O_24,N_19131,N_19122);
or UO_25 (O_25,N_19731,N_19774);
nor UO_26 (O_26,N_19699,N_19576);
nand UO_27 (O_27,N_19889,N_19352);
and UO_28 (O_28,N_19671,N_19529);
nor UO_29 (O_29,N_19664,N_19043);
or UO_30 (O_30,N_19533,N_19246);
and UO_31 (O_31,N_19644,N_19534);
or UO_32 (O_32,N_19905,N_19274);
and UO_33 (O_33,N_19884,N_19171);
nand UO_34 (O_34,N_19215,N_19221);
nor UO_35 (O_35,N_19393,N_19799);
nand UO_36 (O_36,N_19196,N_19142);
or UO_37 (O_37,N_19255,N_19491);
or UO_38 (O_38,N_19360,N_19670);
nor UO_39 (O_39,N_19234,N_19497);
or UO_40 (O_40,N_19660,N_19727);
and UO_41 (O_41,N_19803,N_19174);
xor UO_42 (O_42,N_19044,N_19135);
xnor UO_43 (O_43,N_19751,N_19233);
nand UO_44 (O_44,N_19249,N_19024);
nand UO_45 (O_45,N_19633,N_19172);
xor UO_46 (O_46,N_19828,N_19779);
and UO_47 (O_47,N_19749,N_19941);
or UO_48 (O_48,N_19409,N_19958);
xnor UO_49 (O_49,N_19318,N_19975);
and UO_50 (O_50,N_19207,N_19981);
or UO_51 (O_51,N_19665,N_19213);
nand UO_52 (O_52,N_19150,N_19219);
nand UO_53 (O_53,N_19679,N_19175);
or UO_54 (O_54,N_19220,N_19801);
or UO_55 (O_55,N_19047,N_19381);
nor UO_56 (O_56,N_19940,N_19334);
and UO_57 (O_57,N_19238,N_19503);
nor UO_58 (O_58,N_19663,N_19987);
nand UO_59 (O_59,N_19296,N_19407);
nand UO_60 (O_60,N_19276,N_19645);
nand UO_61 (O_61,N_19906,N_19227);
and UO_62 (O_62,N_19566,N_19232);
nor UO_63 (O_63,N_19514,N_19139);
or UO_64 (O_64,N_19528,N_19190);
nor UO_65 (O_65,N_19230,N_19925);
xor UO_66 (O_66,N_19748,N_19372);
and UO_67 (O_67,N_19753,N_19103);
nand UO_68 (O_68,N_19369,N_19490);
nor UO_69 (O_69,N_19895,N_19713);
or UO_70 (O_70,N_19181,N_19502);
nor UO_71 (O_71,N_19855,N_19085);
nand UO_72 (O_72,N_19452,N_19886);
nor UO_73 (O_73,N_19766,N_19253);
nor UO_74 (O_74,N_19705,N_19904);
and UO_75 (O_75,N_19020,N_19265);
nand UO_76 (O_76,N_19197,N_19011);
nor UO_77 (O_77,N_19775,N_19515);
nor UO_78 (O_78,N_19821,N_19894);
and UO_79 (O_79,N_19165,N_19319);
nor UO_80 (O_80,N_19587,N_19031);
and UO_81 (O_81,N_19540,N_19720);
or UO_82 (O_82,N_19877,N_19025);
nor UO_83 (O_83,N_19991,N_19681);
and UO_84 (O_84,N_19864,N_19721);
nand UO_85 (O_85,N_19707,N_19982);
nor UO_86 (O_86,N_19101,N_19867);
or UO_87 (O_87,N_19283,N_19767);
and UO_88 (O_88,N_19120,N_19259);
xnor UO_89 (O_89,N_19160,N_19102);
and UO_90 (O_90,N_19859,N_19084);
nor UO_91 (O_91,N_19267,N_19494);
or UO_92 (O_92,N_19313,N_19386);
nor UO_93 (O_93,N_19863,N_19539);
or UO_94 (O_94,N_19790,N_19048);
and UO_95 (O_95,N_19537,N_19922);
and UO_96 (O_96,N_19194,N_19642);
nand UO_97 (O_97,N_19898,N_19076);
xor UO_98 (O_98,N_19034,N_19630);
nand UO_99 (O_99,N_19596,N_19408);
and UO_100 (O_100,N_19064,N_19050);
nand UO_101 (O_101,N_19287,N_19467);
xor UO_102 (O_102,N_19366,N_19817);
or UO_103 (O_103,N_19290,N_19154);
xnor UO_104 (O_104,N_19614,N_19564);
and UO_105 (O_105,N_19577,N_19619);
and UO_106 (O_106,N_19829,N_19075);
nor UO_107 (O_107,N_19784,N_19329);
nand UO_108 (O_108,N_19795,N_19033);
nand UO_109 (O_109,N_19873,N_19132);
and UO_110 (O_110,N_19737,N_19682);
or UO_111 (O_111,N_19109,N_19038);
nand UO_112 (O_112,N_19460,N_19239);
nor UO_113 (O_113,N_19170,N_19655);
nand UO_114 (O_114,N_19412,N_19099);
and UO_115 (O_115,N_19847,N_19377);
nand UO_116 (O_116,N_19743,N_19127);
or UO_117 (O_117,N_19579,N_19575);
xnor UO_118 (O_118,N_19559,N_19496);
and UO_119 (O_119,N_19717,N_19964);
nand UO_120 (O_120,N_19183,N_19422);
nand UO_121 (O_121,N_19554,N_19833);
or UO_122 (O_122,N_19164,N_19294);
nor UO_123 (O_123,N_19365,N_19486);
xnor UO_124 (O_124,N_19371,N_19696);
or UO_125 (O_125,N_19482,N_19923);
xnor UO_126 (O_126,N_19734,N_19545);
nor UO_127 (O_127,N_19914,N_19772);
or UO_128 (O_128,N_19505,N_19258);
and UO_129 (O_129,N_19680,N_19692);
nor UO_130 (O_130,N_19901,N_19136);
or UO_131 (O_131,N_19353,N_19493);
nor UO_132 (O_132,N_19688,N_19744);
xnor UO_133 (O_133,N_19001,N_19027);
nor UO_134 (O_134,N_19351,N_19045);
nor UO_135 (O_135,N_19634,N_19809);
and UO_136 (O_136,N_19454,N_19908);
nand UO_137 (O_137,N_19567,N_19338);
nand UO_138 (O_138,N_19957,N_19314);
nor UO_139 (O_139,N_19156,N_19588);
and UO_140 (O_140,N_19231,N_19333);
nand UO_141 (O_141,N_19956,N_19489);
nor UO_142 (O_142,N_19676,N_19969);
or UO_143 (O_143,N_19112,N_19455);
and UO_144 (O_144,N_19667,N_19184);
nor UO_145 (O_145,N_19427,N_19223);
nand UO_146 (O_146,N_19343,N_19677);
xor UO_147 (O_147,N_19469,N_19402);
and UO_148 (O_148,N_19017,N_19245);
nand UO_149 (O_149,N_19307,N_19752);
and UO_150 (O_150,N_19417,N_19060);
nand UO_151 (O_151,N_19029,N_19928);
or UO_152 (O_152,N_19461,N_19512);
nand UO_153 (O_153,N_19330,N_19780);
and UO_154 (O_154,N_19431,N_19598);
and UO_155 (O_155,N_19729,N_19548);
xnor UO_156 (O_156,N_19866,N_19899);
nand UO_157 (O_157,N_19989,N_19757);
or UO_158 (O_158,N_19865,N_19808);
xnor UO_159 (O_159,N_19040,N_19177);
xnor UO_160 (O_160,N_19854,N_19354);
or UO_161 (O_161,N_19214,N_19862);
nand UO_162 (O_162,N_19162,N_19993);
nor UO_163 (O_163,N_19931,N_19998);
and UO_164 (O_164,N_19104,N_19942);
nand UO_165 (O_165,N_19053,N_19921);
or UO_166 (O_166,N_19438,N_19617);
nor UO_167 (O_167,N_19690,N_19145);
or UO_168 (O_168,N_19945,N_19356);
nor UO_169 (O_169,N_19083,N_19740);
nor UO_170 (O_170,N_19643,N_19976);
and UO_171 (O_171,N_19845,N_19275);
nor UO_172 (O_172,N_19979,N_19247);
nand UO_173 (O_173,N_19244,N_19842);
nor UO_174 (O_174,N_19014,N_19445);
xor UO_175 (O_175,N_19069,N_19327);
nor UO_176 (O_176,N_19108,N_19892);
or UO_177 (O_177,N_19544,N_19810);
and UO_178 (O_178,N_19361,N_19201);
nor UO_179 (O_179,N_19202,N_19977);
or UO_180 (O_180,N_19096,N_19189);
nand UO_181 (O_181,N_19052,N_19320);
nand UO_182 (O_182,N_19712,N_19324);
nand UO_183 (O_183,N_19768,N_19441);
nand UO_184 (O_184,N_19144,N_19126);
or UO_185 (O_185,N_19387,N_19794);
or UO_186 (O_186,N_19209,N_19763);
xor UO_187 (O_187,N_19789,N_19517);
or UO_188 (O_188,N_19718,N_19432);
nor UO_189 (O_189,N_19565,N_19668);
nor UO_190 (O_190,N_19986,N_19303);
or UO_191 (O_191,N_19610,N_19997);
or UO_192 (O_192,N_19450,N_19019);
nor UO_193 (O_193,N_19543,N_19755);
nand UO_194 (O_194,N_19278,N_19462);
nor UO_195 (O_195,N_19777,N_19403);
or UO_196 (O_196,N_19423,N_19967);
or UO_197 (O_197,N_19728,N_19272);
xor UO_198 (O_198,N_19693,N_19530);
nand UO_199 (O_199,N_19604,N_19382);
and UO_200 (O_200,N_19268,N_19394);
xnor UO_201 (O_201,N_19954,N_19155);
or UO_202 (O_202,N_19913,N_19058);
nand UO_203 (O_203,N_19100,N_19030);
or UO_204 (O_204,N_19242,N_19008);
or UO_205 (O_205,N_19225,N_19953);
nor UO_206 (O_206,N_19556,N_19002);
nand UO_207 (O_207,N_19439,N_19088);
xnor UO_208 (O_208,N_19947,N_19250);
nand UO_209 (O_209,N_19012,N_19813);
and UO_210 (O_210,N_19414,N_19869);
and UO_211 (O_211,N_19148,N_19446);
and UO_212 (O_212,N_19536,N_19846);
nor UO_213 (O_213,N_19678,N_19153);
nor UO_214 (O_214,N_19988,N_19616);
nand UO_215 (O_215,N_19094,N_19091);
nor UO_216 (O_216,N_19827,N_19335);
nor UO_217 (O_217,N_19235,N_19128);
or UO_218 (O_218,N_19893,N_19036);
nand UO_219 (O_219,N_19107,N_19241);
and UO_220 (O_220,N_19658,N_19373);
nor UO_221 (O_221,N_19054,N_19649);
xnor UO_222 (O_222,N_19695,N_19342);
or UO_223 (O_223,N_19117,N_19581);
and UO_224 (O_224,N_19016,N_19437);
nor UO_225 (O_225,N_19228,N_19385);
and UO_226 (O_226,N_19723,N_19746);
nor UO_227 (O_227,N_19625,N_19613);
xor UO_228 (O_228,N_19355,N_19442);
nand UO_229 (O_229,N_19822,N_19811);
and UO_230 (O_230,N_19764,N_19015);
and UO_231 (O_231,N_19023,N_19130);
xnor UO_232 (O_232,N_19648,N_19295);
nand UO_233 (O_233,N_19800,N_19281);
and UO_234 (O_234,N_19972,N_19310);
nand UO_235 (O_235,N_19282,N_19032);
xnor UO_236 (O_236,N_19602,N_19123);
nand UO_237 (O_237,N_19637,N_19451);
or UO_238 (O_238,N_19555,N_19546);
and UO_239 (O_239,N_19237,N_19594);
or UO_240 (O_240,N_19137,N_19035);
xnor UO_241 (O_241,N_19878,N_19158);
and UO_242 (O_242,N_19735,N_19492);
and UO_243 (O_243,N_19896,N_19420);
nor UO_244 (O_244,N_19345,N_19909);
and UO_245 (O_245,N_19968,N_19708);
nand UO_246 (O_246,N_19405,N_19631);
and UO_247 (O_247,N_19284,N_19971);
nor UO_248 (O_248,N_19669,N_19114);
xor UO_249 (O_249,N_19316,N_19443);
nor UO_250 (O_250,N_19071,N_19483);
and UO_251 (O_251,N_19413,N_19191);
nor UO_252 (O_252,N_19018,N_19252);
and UO_253 (O_253,N_19638,N_19879);
nand UO_254 (O_254,N_19912,N_19951);
xnor UO_255 (O_255,N_19325,N_19583);
and UO_256 (O_256,N_19698,N_19349);
nor UO_257 (O_257,N_19985,N_19357);
or UO_258 (O_258,N_19806,N_19666);
and UO_259 (O_259,N_19599,N_19725);
nand UO_260 (O_260,N_19541,N_19858);
or UO_261 (O_261,N_19632,N_19820);
and UO_262 (O_262,N_19124,N_19066);
nor UO_263 (O_263,N_19419,N_19902);
and UO_264 (O_264,N_19433,N_19261);
and UO_265 (O_265,N_19778,N_19297);
and UO_266 (O_266,N_19856,N_19042);
or UO_267 (O_267,N_19662,N_19063);
nand UO_268 (O_268,N_19340,N_19870);
nand UO_269 (O_269,N_19691,N_19410);
nand UO_270 (O_270,N_19121,N_19169);
and UO_271 (O_271,N_19871,N_19759);
and UO_272 (O_272,N_19163,N_19785);
and UO_273 (O_273,N_19618,N_19472);
or UO_274 (O_274,N_19157,N_19138);
and UO_275 (O_275,N_19525,N_19920);
and UO_276 (O_276,N_19756,N_19974);
nor UO_277 (O_277,N_19570,N_19176);
and UO_278 (O_278,N_19983,N_19933);
and UO_279 (O_279,N_19211,N_19262);
nand UO_280 (O_280,N_19118,N_19558);
and UO_281 (O_281,N_19346,N_19584);
and UO_282 (O_282,N_19640,N_19733);
nor UO_283 (O_283,N_19955,N_19673);
or UO_284 (O_284,N_19994,N_19203);
nand UO_285 (O_285,N_19390,N_19398);
xnor UO_286 (O_286,N_19504,N_19519);
and UO_287 (O_287,N_19585,N_19092);
or UO_288 (O_288,N_19661,N_19830);
and UO_289 (O_289,N_19990,N_19222);
and UO_290 (O_290,N_19021,N_19654);
nor UO_291 (O_291,N_19783,N_19814);
nand UO_292 (O_292,N_19111,N_19070);
xor UO_293 (O_293,N_19747,N_19341);
and UO_294 (O_294,N_19623,N_19694);
nand UO_295 (O_295,N_19459,N_19271);
and UO_296 (O_296,N_19273,N_19046);
nor UO_297 (O_297,N_19093,N_19919);
nor UO_298 (O_298,N_19257,N_19890);
and UO_299 (O_299,N_19980,N_19831);
nand UO_300 (O_300,N_19119,N_19569);
or UO_301 (O_301,N_19832,N_19416);
nand UO_302 (O_302,N_19105,N_19178);
and UO_303 (O_303,N_19507,N_19736);
nand UO_304 (O_304,N_19949,N_19580);
or UO_305 (O_305,N_19309,N_19348);
or UO_306 (O_306,N_19900,N_19885);
nor UO_307 (O_307,N_19315,N_19636);
nand UO_308 (O_308,N_19097,N_19264);
or UO_309 (O_309,N_19824,N_19500);
xnor UO_310 (O_310,N_19430,N_19627);
or UO_311 (O_311,N_19473,N_19010);
or UO_312 (O_312,N_19595,N_19819);
nand UO_313 (O_313,N_19875,N_19639);
or UO_314 (O_314,N_19788,N_19470);
xor UO_315 (O_315,N_19269,N_19391);
and UO_316 (O_316,N_19797,N_19406);
and UO_317 (O_317,N_19802,N_19719);
and UO_318 (O_318,N_19600,N_19605);
nor UO_319 (O_319,N_19350,N_19798);
xor UO_320 (O_320,N_19383,N_19840);
nor UO_321 (O_321,N_19098,N_19301);
nand UO_322 (O_322,N_19347,N_19805);
nand UO_323 (O_323,N_19306,N_19204);
or UO_324 (O_324,N_19090,N_19603);
xnor UO_325 (O_325,N_19876,N_19198);
nand UO_326 (O_326,N_19161,N_19151);
and UO_327 (O_327,N_19911,N_19488);
or UO_328 (O_328,N_19750,N_19844);
nor UO_329 (O_329,N_19321,N_19304);
or UO_330 (O_330,N_19336,N_19765);
nor UO_331 (O_331,N_19952,N_19995);
nand UO_332 (O_332,N_19984,N_19841);
and UO_333 (O_333,N_19730,N_19463);
and UO_334 (O_334,N_19224,N_19464);
nor UO_335 (O_335,N_19037,N_19448);
nor UO_336 (O_336,N_19078,N_19966);
and UO_337 (O_337,N_19129,N_19738);
or UO_338 (O_338,N_19551,N_19970);
nand UO_339 (O_339,N_19560,N_19641);
nor UO_340 (O_340,N_19305,N_19068);
or UO_341 (O_341,N_19080,N_19963);
or UO_342 (O_342,N_19792,N_19557);
nand UO_343 (O_343,N_19839,N_19055);
nor UO_344 (O_344,N_19293,N_19888);
nand UO_345 (O_345,N_19770,N_19049);
or UO_346 (O_346,N_19339,N_19149);
xnor UO_347 (O_347,N_19650,N_19476);
nand UO_348 (O_348,N_19948,N_19518);
and UO_349 (O_349,N_19552,N_19843);
nand UO_350 (O_350,N_19095,N_19251);
or UO_351 (O_351,N_19714,N_19005);
nor UO_352 (O_352,N_19368,N_19672);
xnor UO_353 (O_353,N_19513,N_19961);
nand UO_354 (O_354,N_19742,N_19447);
xor UO_355 (O_355,N_19004,N_19179);
and UO_356 (O_356,N_19615,N_19086);
nor UO_357 (O_357,N_19110,N_19838);
or UO_358 (O_358,N_19180,N_19480);
nor UO_359 (O_359,N_19266,N_19837);
or UO_360 (O_360,N_19199,N_19999);
or UO_361 (O_361,N_19166,N_19192);
nor UO_362 (O_362,N_19429,N_19563);
nor UO_363 (O_363,N_19415,N_19256);
or UO_364 (O_364,N_19485,N_19374);
and UO_365 (O_365,N_19411,N_19769);
nor UO_366 (O_366,N_19270,N_19860);
and UO_367 (O_367,N_19499,N_19444);
and UO_368 (O_368,N_19188,N_19773);
nand UO_369 (O_369,N_19629,N_19849);
nand UO_370 (O_370,N_19061,N_19726);
and UO_371 (O_371,N_19932,N_19289);
nand UO_372 (O_372,N_19152,N_19960);
or UO_373 (O_373,N_19125,N_19881);
nand UO_374 (O_374,N_19397,N_19973);
or UO_375 (O_375,N_19816,N_19950);
nor UO_376 (O_376,N_19479,N_19187);
and UO_377 (O_377,N_19051,N_19704);
nor UO_378 (O_378,N_19520,N_19572);
or UO_379 (O_379,N_19299,N_19147);
or UO_380 (O_380,N_19703,N_19378);
and UO_381 (O_381,N_19701,N_19685);
and UO_382 (O_382,N_19300,N_19079);
nor UO_383 (O_383,N_19635,N_19597);
or UO_384 (O_384,N_19426,N_19791);
or UO_385 (O_385,N_19140,N_19586);
nor UO_386 (O_386,N_19173,N_19850);
nor UO_387 (O_387,N_19526,N_19481);
nor UO_388 (O_388,N_19826,N_19651);
or UO_389 (O_389,N_19487,N_19946);
nand UO_390 (O_390,N_19523,N_19868);
and UO_391 (O_391,N_19522,N_19907);
and UO_392 (O_392,N_19167,N_19065);
nor UO_393 (O_393,N_19607,N_19206);
and UO_394 (O_394,N_19146,N_19626);
nand UO_395 (O_395,N_19421,N_19280);
and UO_396 (O_396,N_19916,N_19609);
xor UO_397 (O_397,N_19396,N_19815);
or UO_398 (O_398,N_19186,N_19317);
or UO_399 (O_399,N_19601,N_19308);
and UO_400 (O_400,N_19684,N_19359);
or UO_401 (O_401,N_19722,N_19217);
and UO_402 (O_402,N_19996,N_19754);
xnor UO_403 (O_403,N_19836,N_19535);
or UO_404 (O_404,N_19574,N_19506);
and UO_405 (O_405,N_19475,N_19776);
or UO_406 (O_406,N_19796,N_19057);
nor UO_407 (O_407,N_19659,N_19547);
nor UO_408 (O_408,N_19400,N_19236);
and UO_409 (O_409,N_19388,N_19562);
nor UO_410 (O_410,N_19200,N_19077);
and UO_411 (O_411,N_19573,N_19457);
and UO_412 (O_412,N_19364,N_19477);
nand UO_413 (O_413,N_19938,N_19715);
xor UO_414 (O_414,N_19022,N_19700);
and UO_415 (O_415,N_19185,N_19612);
nor UO_416 (O_416,N_19761,N_19807);
or UO_417 (O_417,N_19380,N_19062);
and UO_418 (O_418,N_19910,N_19656);
and UO_419 (O_419,N_19782,N_19006);
xor UO_420 (O_420,N_19007,N_19424);
or UO_421 (O_421,N_19883,N_19322);
nor UO_422 (O_422,N_19834,N_19711);
nor UO_423 (O_423,N_19279,N_19652);
nor UO_424 (O_424,N_19067,N_19298);
nand UO_425 (O_425,N_19697,N_19468);
nand UO_426 (O_426,N_19592,N_19362);
and UO_427 (O_427,N_19229,N_19291);
or UO_428 (O_428,N_19288,N_19702);
and UO_429 (O_429,N_19510,N_19745);
xnor UO_430 (O_430,N_19495,N_19474);
or UO_431 (O_431,N_19392,N_19003);
and UO_432 (O_432,N_19216,N_19218);
nor UO_433 (O_433,N_19818,N_19992);
nor UO_434 (O_434,N_19182,N_19263);
or UO_435 (O_435,N_19484,N_19732);
or UO_436 (O_436,N_19606,N_19466);
nor UO_437 (O_437,N_19787,N_19226);
nand UO_438 (O_438,N_19918,N_19337);
xor UO_439 (O_439,N_19113,N_19965);
and UO_440 (O_440,N_19260,N_19399);
xor UO_441 (O_441,N_19248,N_19561);
nor UO_442 (O_442,N_19212,N_19926);
xor UO_443 (O_443,N_19292,N_19059);
xor UO_444 (O_444,N_19542,N_19509);
and UO_445 (O_445,N_19825,N_19929);
or UO_446 (O_446,N_19143,N_19401);
and UO_447 (O_447,N_19683,N_19891);
or UO_448 (O_448,N_19243,N_19312);
nor UO_449 (O_449,N_19302,N_19013);
or UO_450 (O_450,N_19646,N_19771);
nor UO_451 (O_451,N_19880,N_19449);
and UO_452 (O_452,N_19082,N_19591);
or UO_453 (O_453,N_19195,N_19072);
and UO_454 (O_454,N_19674,N_19168);
nand UO_455 (O_455,N_19959,N_19897);
and UO_456 (O_456,N_19628,N_19328);
and UO_457 (O_457,N_19872,N_19675);
nand UO_458 (O_458,N_19501,N_19578);
nor UO_459 (O_459,N_19436,N_19924);
xor UO_460 (O_460,N_19367,N_19254);
nor UO_461 (O_461,N_19159,N_19435);
and UO_462 (O_462,N_19590,N_19571);
and UO_463 (O_463,N_19286,N_19532);
and UO_464 (O_464,N_19508,N_19009);
and UO_465 (O_465,N_19384,N_19936);
and UO_466 (O_466,N_19106,N_19848);
xor UO_467 (O_467,N_19582,N_19471);
or UO_468 (O_468,N_19395,N_19709);
and UO_469 (O_469,N_19285,N_19934);
or UO_470 (O_470,N_19593,N_19375);
nor UO_471 (O_471,N_19089,N_19379);
and UO_472 (O_472,N_19389,N_19653);
xnor UO_473 (O_473,N_19344,N_19857);
or UO_474 (O_474,N_19453,N_19418);
and UO_475 (O_475,N_19332,N_19425);
nor UO_476 (O_476,N_19087,N_19937);
or UO_477 (O_477,N_19458,N_19516);
or UO_478 (O_478,N_19874,N_19716);
nor UO_479 (O_479,N_19000,N_19758);
and UO_480 (O_480,N_19404,N_19852);
and UO_481 (O_481,N_19589,N_19739);
or UO_482 (O_482,N_19657,N_19208);
and UO_483 (O_483,N_19478,N_19205);
or UO_484 (O_484,N_19903,N_19568);
nor UO_485 (O_485,N_19039,N_19935);
and UO_486 (O_486,N_19141,N_19511);
or UO_487 (O_487,N_19311,N_19527);
xor UO_488 (O_488,N_19277,N_19434);
nand UO_489 (O_489,N_19882,N_19465);
and UO_490 (O_490,N_19074,N_19793);
or UO_491 (O_491,N_19724,N_19853);
nor UO_492 (O_492,N_19620,N_19917);
and UO_493 (O_493,N_19550,N_19056);
nor UO_494 (O_494,N_19608,N_19927);
and UO_495 (O_495,N_19611,N_19915);
nor UO_496 (O_496,N_19553,N_19835);
nand UO_497 (O_497,N_19781,N_19689);
nand UO_498 (O_498,N_19851,N_19116);
or UO_499 (O_499,N_19804,N_19741);
xor UO_500 (O_500,N_19143,N_19156);
xor UO_501 (O_501,N_19149,N_19440);
nor UO_502 (O_502,N_19117,N_19768);
or UO_503 (O_503,N_19293,N_19546);
and UO_504 (O_504,N_19859,N_19026);
nor UO_505 (O_505,N_19811,N_19761);
and UO_506 (O_506,N_19074,N_19443);
or UO_507 (O_507,N_19093,N_19670);
xor UO_508 (O_508,N_19055,N_19728);
or UO_509 (O_509,N_19180,N_19935);
and UO_510 (O_510,N_19322,N_19950);
nor UO_511 (O_511,N_19553,N_19296);
and UO_512 (O_512,N_19679,N_19887);
nand UO_513 (O_513,N_19287,N_19583);
and UO_514 (O_514,N_19458,N_19002);
nand UO_515 (O_515,N_19411,N_19825);
xnor UO_516 (O_516,N_19109,N_19450);
and UO_517 (O_517,N_19740,N_19957);
or UO_518 (O_518,N_19336,N_19029);
nor UO_519 (O_519,N_19525,N_19200);
nor UO_520 (O_520,N_19543,N_19227);
nand UO_521 (O_521,N_19723,N_19507);
or UO_522 (O_522,N_19031,N_19230);
and UO_523 (O_523,N_19753,N_19892);
nor UO_524 (O_524,N_19467,N_19126);
and UO_525 (O_525,N_19824,N_19873);
nor UO_526 (O_526,N_19417,N_19347);
or UO_527 (O_527,N_19373,N_19069);
or UO_528 (O_528,N_19553,N_19188);
and UO_529 (O_529,N_19024,N_19463);
nand UO_530 (O_530,N_19058,N_19794);
xor UO_531 (O_531,N_19023,N_19891);
or UO_532 (O_532,N_19209,N_19478);
nor UO_533 (O_533,N_19140,N_19602);
nor UO_534 (O_534,N_19656,N_19348);
or UO_535 (O_535,N_19952,N_19156);
nor UO_536 (O_536,N_19816,N_19896);
nand UO_537 (O_537,N_19904,N_19816);
or UO_538 (O_538,N_19787,N_19598);
nor UO_539 (O_539,N_19108,N_19379);
and UO_540 (O_540,N_19945,N_19197);
or UO_541 (O_541,N_19071,N_19014);
or UO_542 (O_542,N_19796,N_19635);
nor UO_543 (O_543,N_19386,N_19920);
or UO_544 (O_544,N_19171,N_19453);
nor UO_545 (O_545,N_19037,N_19713);
nand UO_546 (O_546,N_19550,N_19856);
or UO_547 (O_547,N_19243,N_19764);
nor UO_548 (O_548,N_19149,N_19627);
or UO_549 (O_549,N_19882,N_19021);
and UO_550 (O_550,N_19706,N_19247);
and UO_551 (O_551,N_19431,N_19591);
xor UO_552 (O_552,N_19333,N_19147);
nor UO_553 (O_553,N_19245,N_19529);
and UO_554 (O_554,N_19735,N_19630);
nor UO_555 (O_555,N_19626,N_19765);
nor UO_556 (O_556,N_19696,N_19309);
and UO_557 (O_557,N_19845,N_19724);
nand UO_558 (O_558,N_19808,N_19404);
and UO_559 (O_559,N_19057,N_19107);
and UO_560 (O_560,N_19286,N_19118);
nand UO_561 (O_561,N_19527,N_19095);
nor UO_562 (O_562,N_19762,N_19842);
nor UO_563 (O_563,N_19644,N_19634);
nor UO_564 (O_564,N_19878,N_19940);
nor UO_565 (O_565,N_19667,N_19041);
xor UO_566 (O_566,N_19266,N_19224);
xnor UO_567 (O_567,N_19125,N_19468);
and UO_568 (O_568,N_19014,N_19243);
nand UO_569 (O_569,N_19144,N_19167);
nor UO_570 (O_570,N_19346,N_19287);
and UO_571 (O_571,N_19344,N_19199);
and UO_572 (O_572,N_19833,N_19520);
and UO_573 (O_573,N_19539,N_19445);
nor UO_574 (O_574,N_19211,N_19203);
and UO_575 (O_575,N_19226,N_19441);
or UO_576 (O_576,N_19457,N_19423);
nand UO_577 (O_577,N_19100,N_19934);
and UO_578 (O_578,N_19700,N_19944);
nor UO_579 (O_579,N_19313,N_19762);
nor UO_580 (O_580,N_19619,N_19680);
nor UO_581 (O_581,N_19837,N_19533);
and UO_582 (O_582,N_19267,N_19949);
nand UO_583 (O_583,N_19879,N_19693);
or UO_584 (O_584,N_19323,N_19032);
or UO_585 (O_585,N_19165,N_19884);
xnor UO_586 (O_586,N_19444,N_19455);
or UO_587 (O_587,N_19453,N_19760);
nand UO_588 (O_588,N_19222,N_19401);
nor UO_589 (O_589,N_19037,N_19231);
and UO_590 (O_590,N_19378,N_19824);
nand UO_591 (O_591,N_19944,N_19346);
or UO_592 (O_592,N_19449,N_19491);
or UO_593 (O_593,N_19036,N_19497);
and UO_594 (O_594,N_19483,N_19033);
and UO_595 (O_595,N_19500,N_19532);
nand UO_596 (O_596,N_19284,N_19556);
and UO_597 (O_597,N_19427,N_19112);
nor UO_598 (O_598,N_19788,N_19119);
and UO_599 (O_599,N_19877,N_19787);
or UO_600 (O_600,N_19039,N_19561);
or UO_601 (O_601,N_19799,N_19440);
xnor UO_602 (O_602,N_19470,N_19904);
or UO_603 (O_603,N_19519,N_19399);
xor UO_604 (O_604,N_19308,N_19920);
nor UO_605 (O_605,N_19604,N_19611);
or UO_606 (O_606,N_19883,N_19308);
nor UO_607 (O_607,N_19837,N_19534);
or UO_608 (O_608,N_19929,N_19746);
or UO_609 (O_609,N_19388,N_19638);
xor UO_610 (O_610,N_19645,N_19562);
nor UO_611 (O_611,N_19711,N_19376);
nand UO_612 (O_612,N_19910,N_19759);
or UO_613 (O_613,N_19863,N_19636);
or UO_614 (O_614,N_19524,N_19717);
nor UO_615 (O_615,N_19925,N_19218);
xnor UO_616 (O_616,N_19195,N_19864);
nor UO_617 (O_617,N_19827,N_19324);
nand UO_618 (O_618,N_19649,N_19606);
nor UO_619 (O_619,N_19460,N_19620);
or UO_620 (O_620,N_19619,N_19763);
nand UO_621 (O_621,N_19165,N_19215);
nand UO_622 (O_622,N_19722,N_19347);
xnor UO_623 (O_623,N_19750,N_19846);
nand UO_624 (O_624,N_19478,N_19043);
nand UO_625 (O_625,N_19675,N_19660);
or UO_626 (O_626,N_19313,N_19614);
and UO_627 (O_627,N_19474,N_19135);
or UO_628 (O_628,N_19255,N_19137);
xnor UO_629 (O_629,N_19995,N_19950);
nor UO_630 (O_630,N_19423,N_19589);
nor UO_631 (O_631,N_19397,N_19870);
or UO_632 (O_632,N_19021,N_19854);
nor UO_633 (O_633,N_19420,N_19659);
nor UO_634 (O_634,N_19958,N_19550);
nand UO_635 (O_635,N_19700,N_19063);
nor UO_636 (O_636,N_19408,N_19227);
nor UO_637 (O_637,N_19099,N_19669);
nand UO_638 (O_638,N_19128,N_19865);
nor UO_639 (O_639,N_19314,N_19615);
or UO_640 (O_640,N_19075,N_19583);
nor UO_641 (O_641,N_19866,N_19064);
and UO_642 (O_642,N_19625,N_19433);
and UO_643 (O_643,N_19904,N_19932);
or UO_644 (O_644,N_19433,N_19246);
nor UO_645 (O_645,N_19185,N_19459);
and UO_646 (O_646,N_19817,N_19043);
nor UO_647 (O_647,N_19521,N_19774);
and UO_648 (O_648,N_19763,N_19434);
nor UO_649 (O_649,N_19243,N_19273);
or UO_650 (O_650,N_19436,N_19789);
xnor UO_651 (O_651,N_19496,N_19927);
nor UO_652 (O_652,N_19427,N_19739);
nor UO_653 (O_653,N_19003,N_19515);
or UO_654 (O_654,N_19485,N_19661);
nand UO_655 (O_655,N_19153,N_19796);
nor UO_656 (O_656,N_19494,N_19034);
nand UO_657 (O_657,N_19421,N_19603);
nand UO_658 (O_658,N_19855,N_19073);
xor UO_659 (O_659,N_19456,N_19457);
or UO_660 (O_660,N_19498,N_19270);
nand UO_661 (O_661,N_19722,N_19750);
and UO_662 (O_662,N_19148,N_19841);
nand UO_663 (O_663,N_19171,N_19696);
and UO_664 (O_664,N_19935,N_19315);
nor UO_665 (O_665,N_19767,N_19198);
or UO_666 (O_666,N_19003,N_19696);
or UO_667 (O_667,N_19521,N_19169);
nand UO_668 (O_668,N_19870,N_19117);
or UO_669 (O_669,N_19197,N_19784);
xor UO_670 (O_670,N_19008,N_19001);
xnor UO_671 (O_671,N_19669,N_19782);
or UO_672 (O_672,N_19637,N_19674);
or UO_673 (O_673,N_19099,N_19303);
nand UO_674 (O_674,N_19168,N_19596);
and UO_675 (O_675,N_19481,N_19329);
nand UO_676 (O_676,N_19434,N_19513);
nor UO_677 (O_677,N_19352,N_19623);
xnor UO_678 (O_678,N_19273,N_19486);
nor UO_679 (O_679,N_19205,N_19835);
or UO_680 (O_680,N_19042,N_19011);
xnor UO_681 (O_681,N_19104,N_19686);
xnor UO_682 (O_682,N_19362,N_19699);
and UO_683 (O_683,N_19462,N_19029);
nand UO_684 (O_684,N_19908,N_19924);
nand UO_685 (O_685,N_19928,N_19660);
and UO_686 (O_686,N_19148,N_19557);
or UO_687 (O_687,N_19168,N_19784);
and UO_688 (O_688,N_19008,N_19231);
nor UO_689 (O_689,N_19458,N_19913);
and UO_690 (O_690,N_19448,N_19027);
and UO_691 (O_691,N_19730,N_19852);
nand UO_692 (O_692,N_19317,N_19401);
nand UO_693 (O_693,N_19261,N_19309);
or UO_694 (O_694,N_19493,N_19375);
nand UO_695 (O_695,N_19049,N_19438);
or UO_696 (O_696,N_19583,N_19013);
nand UO_697 (O_697,N_19321,N_19179);
and UO_698 (O_698,N_19078,N_19095);
or UO_699 (O_699,N_19151,N_19261);
xor UO_700 (O_700,N_19789,N_19932);
or UO_701 (O_701,N_19276,N_19374);
nand UO_702 (O_702,N_19004,N_19725);
and UO_703 (O_703,N_19097,N_19709);
nand UO_704 (O_704,N_19218,N_19451);
nand UO_705 (O_705,N_19950,N_19903);
nand UO_706 (O_706,N_19246,N_19635);
or UO_707 (O_707,N_19578,N_19776);
nor UO_708 (O_708,N_19028,N_19984);
nor UO_709 (O_709,N_19214,N_19320);
nor UO_710 (O_710,N_19079,N_19834);
nand UO_711 (O_711,N_19232,N_19376);
and UO_712 (O_712,N_19366,N_19671);
and UO_713 (O_713,N_19149,N_19873);
nor UO_714 (O_714,N_19898,N_19929);
and UO_715 (O_715,N_19015,N_19100);
nor UO_716 (O_716,N_19191,N_19653);
and UO_717 (O_717,N_19397,N_19232);
or UO_718 (O_718,N_19859,N_19704);
or UO_719 (O_719,N_19992,N_19018);
nor UO_720 (O_720,N_19486,N_19604);
nand UO_721 (O_721,N_19329,N_19155);
and UO_722 (O_722,N_19750,N_19455);
or UO_723 (O_723,N_19233,N_19473);
or UO_724 (O_724,N_19307,N_19774);
nand UO_725 (O_725,N_19412,N_19709);
nand UO_726 (O_726,N_19564,N_19899);
and UO_727 (O_727,N_19664,N_19268);
nand UO_728 (O_728,N_19572,N_19914);
nand UO_729 (O_729,N_19588,N_19978);
or UO_730 (O_730,N_19772,N_19706);
and UO_731 (O_731,N_19429,N_19059);
nand UO_732 (O_732,N_19717,N_19447);
nand UO_733 (O_733,N_19181,N_19323);
and UO_734 (O_734,N_19902,N_19953);
nor UO_735 (O_735,N_19172,N_19335);
or UO_736 (O_736,N_19989,N_19685);
or UO_737 (O_737,N_19719,N_19616);
nor UO_738 (O_738,N_19102,N_19973);
nor UO_739 (O_739,N_19831,N_19620);
or UO_740 (O_740,N_19054,N_19714);
or UO_741 (O_741,N_19229,N_19701);
or UO_742 (O_742,N_19825,N_19161);
nand UO_743 (O_743,N_19950,N_19344);
or UO_744 (O_744,N_19617,N_19687);
or UO_745 (O_745,N_19937,N_19212);
or UO_746 (O_746,N_19677,N_19153);
and UO_747 (O_747,N_19954,N_19817);
and UO_748 (O_748,N_19924,N_19882);
nand UO_749 (O_749,N_19038,N_19724);
or UO_750 (O_750,N_19042,N_19137);
nor UO_751 (O_751,N_19731,N_19017);
xnor UO_752 (O_752,N_19170,N_19989);
nand UO_753 (O_753,N_19067,N_19043);
and UO_754 (O_754,N_19067,N_19303);
and UO_755 (O_755,N_19402,N_19392);
nor UO_756 (O_756,N_19671,N_19242);
nand UO_757 (O_757,N_19918,N_19506);
or UO_758 (O_758,N_19263,N_19608);
xor UO_759 (O_759,N_19392,N_19005);
and UO_760 (O_760,N_19965,N_19430);
nand UO_761 (O_761,N_19322,N_19175);
nor UO_762 (O_762,N_19951,N_19271);
nor UO_763 (O_763,N_19136,N_19721);
nand UO_764 (O_764,N_19146,N_19650);
and UO_765 (O_765,N_19376,N_19732);
nor UO_766 (O_766,N_19313,N_19435);
nor UO_767 (O_767,N_19865,N_19211);
or UO_768 (O_768,N_19446,N_19930);
nor UO_769 (O_769,N_19819,N_19000);
nand UO_770 (O_770,N_19604,N_19983);
nor UO_771 (O_771,N_19315,N_19724);
and UO_772 (O_772,N_19972,N_19738);
nor UO_773 (O_773,N_19890,N_19438);
nand UO_774 (O_774,N_19246,N_19477);
or UO_775 (O_775,N_19064,N_19288);
or UO_776 (O_776,N_19412,N_19175);
and UO_777 (O_777,N_19379,N_19994);
xor UO_778 (O_778,N_19267,N_19376);
nand UO_779 (O_779,N_19111,N_19329);
xor UO_780 (O_780,N_19620,N_19149);
nand UO_781 (O_781,N_19077,N_19933);
and UO_782 (O_782,N_19974,N_19405);
and UO_783 (O_783,N_19817,N_19468);
nor UO_784 (O_784,N_19233,N_19014);
and UO_785 (O_785,N_19497,N_19737);
or UO_786 (O_786,N_19455,N_19240);
or UO_787 (O_787,N_19287,N_19305);
or UO_788 (O_788,N_19877,N_19655);
nor UO_789 (O_789,N_19934,N_19858);
and UO_790 (O_790,N_19092,N_19261);
nand UO_791 (O_791,N_19797,N_19565);
nand UO_792 (O_792,N_19466,N_19402);
nand UO_793 (O_793,N_19879,N_19715);
nand UO_794 (O_794,N_19695,N_19040);
xor UO_795 (O_795,N_19984,N_19766);
nor UO_796 (O_796,N_19215,N_19320);
and UO_797 (O_797,N_19463,N_19894);
nand UO_798 (O_798,N_19325,N_19699);
or UO_799 (O_799,N_19900,N_19570);
and UO_800 (O_800,N_19301,N_19499);
nand UO_801 (O_801,N_19495,N_19613);
nand UO_802 (O_802,N_19438,N_19032);
and UO_803 (O_803,N_19098,N_19278);
and UO_804 (O_804,N_19591,N_19411);
and UO_805 (O_805,N_19020,N_19854);
or UO_806 (O_806,N_19897,N_19751);
nor UO_807 (O_807,N_19248,N_19752);
nor UO_808 (O_808,N_19631,N_19504);
nor UO_809 (O_809,N_19280,N_19255);
xor UO_810 (O_810,N_19427,N_19083);
nor UO_811 (O_811,N_19503,N_19909);
nor UO_812 (O_812,N_19218,N_19144);
nand UO_813 (O_813,N_19789,N_19678);
and UO_814 (O_814,N_19631,N_19626);
nor UO_815 (O_815,N_19746,N_19013);
or UO_816 (O_816,N_19625,N_19392);
or UO_817 (O_817,N_19257,N_19658);
nand UO_818 (O_818,N_19099,N_19165);
and UO_819 (O_819,N_19431,N_19144);
nand UO_820 (O_820,N_19656,N_19454);
or UO_821 (O_821,N_19260,N_19569);
nor UO_822 (O_822,N_19689,N_19904);
xnor UO_823 (O_823,N_19889,N_19494);
nor UO_824 (O_824,N_19137,N_19706);
nand UO_825 (O_825,N_19803,N_19410);
or UO_826 (O_826,N_19020,N_19621);
xnor UO_827 (O_827,N_19623,N_19072);
nor UO_828 (O_828,N_19228,N_19812);
nor UO_829 (O_829,N_19007,N_19809);
nor UO_830 (O_830,N_19992,N_19569);
nor UO_831 (O_831,N_19158,N_19025);
nand UO_832 (O_832,N_19508,N_19450);
or UO_833 (O_833,N_19123,N_19076);
nand UO_834 (O_834,N_19390,N_19616);
nand UO_835 (O_835,N_19716,N_19049);
or UO_836 (O_836,N_19965,N_19389);
nand UO_837 (O_837,N_19441,N_19663);
or UO_838 (O_838,N_19949,N_19321);
nand UO_839 (O_839,N_19451,N_19759);
or UO_840 (O_840,N_19740,N_19905);
or UO_841 (O_841,N_19856,N_19084);
and UO_842 (O_842,N_19582,N_19392);
xnor UO_843 (O_843,N_19492,N_19843);
nor UO_844 (O_844,N_19931,N_19860);
or UO_845 (O_845,N_19320,N_19250);
nor UO_846 (O_846,N_19471,N_19860);
nand UO_847 (O_847,N_19069,N_19838);
or UO_848 (O_848,N_19621,N_19405);
nand UO_849 (O_849,N_19255,N_19251);
or UO_850 (O_850,N_19426,N_19568);
xnor UO_851 (O_851,N_19422,N_19061);
xnor UO_852 (O_852,N_19268,N_19902);
or UO_853 (O_853,N_19872,N_19768);
and UO_854 (O_854,N_19443,N_19486);
or UO_855 (O_855,N_19375,N_19923);
nor UO_856 (O_856,N_19885,N_19296);
xor UO_857 (O_857,N_19429,N_19466);
or UO_858 (O_858,N_19302,N_19512);
nand UO_859 (O_859,N_19232,N_19525);
nor UO_860 (O_860,N_19825,N_19326);
or UO_861 (O_861,N_19738,N_19003);
or UO_862 (O_862,N_19381,N_19914);
nor UO_863 (O_863,N_19600,N_19925);
or UO_864 (O_864,N_19265,N_19763);
nand UO_865 (O_865,N_19681,N_19419);
nor UO_866 (O_866,N_19033,N_19354);
and UO_867 (O_867,N_19273,N_19400);
nor UO_868 (O_868,N_19767,N_19844);
or UO_869 (O_869,N_19636,N_19793);
and UO_870 (O_870,N_19226,N_19217);
nor UO_871 (O_871,N_19093,N_19885);
xor UO_872 (O_872,N_19390,N_19297);
nand UO_873 (O_873,N_19130,N_19120);
nor UO_874 (O_874,N_19088,N_19404);
nor UO_875 (O_875,N_19037,N_19716);
xnor UO_876 (O_876,N_19322,N_19434);
or UO_877 (O_877,N_19831,N_19556);
and UO_878 (O_878,N_19023,N_19121);
nor UO_879 (O_879,N_19732,N_19238);
nand UO_880 (O_880,N_19739,N_19569);
and UO_881 (O_881,N_19452,N_19014);
or UO_882 (O_882,N_19756,N_19000);
and UO_883 (O_883,N_19957,N_19321);
xnor UO_884 (O_884,N_19774,N_19368);
xor UO_885 (O_885,N_19207,N_19841);
nor UO_886 (O_886,N_19424,N_19242);
or UO_887 (O_887,N_19486,N_19332);
and UO_888 (O_888,N_19410,N_19051);
nor UO_889 (O_889,N_19104,N_19936);
and UO_890 (O_890,N_19580,N_19355);
nand UO_891 (O_891,N_19800,N_19075);
xnor UO_892 (O_892,N_19705,N_19651);
and UO_893 (O_893,N_19331,N_19681);
nand UO_894 (O_894,N_19475,N_19900);
and UO_895 (O_895,N_19103,N_19839);
nand UO_896 (O_896,N_19862,N_19699);
or UO_897 (O_897,N_19957,N_19766);
nand UO_898 (O_898,N_19828,N_19745);
and UO_899 (O_899,N_19901,N_19232);
or UO_900 (O_900,N_19695,N_19348);
xor UO_901 (O_901,N_19127,N_19480);
and UO_902 (O_902,N_19760,N_19899);
nand UO_903 (O_903,N_19723,N_19334);
nor UO_904 (O_904,N_19278,N_19421);
nand UO_905 (O_905,N_19118,N_19571);
nand UO_906 (O_906,N_19151,N_19729);
nand UO_907 (O_907,N_19515,N_19739);
nor UO_908 (O_908,N_19073,N_19632);
and UO_909 (O_909,N_19093,N_19023);
nand UO_910 (O_910,N_19104,N_19325);
or UO_911 (O_911,N_19838,N_19642);
nor UO_912 (O_912,N_19696,N_19008);
and UO_913 (O_913,N_19903,N_19314);
nand UO_914 (O_914,N_19517,N_19023);
nor UO_915 (O_915,N_19460,N_19838);
nor UO_916 (O_916,N_19841,N_19652);
or UO_917 (O_917,N_19161,N_19455);
nand UO_918 (O_918,N_19574,N_19413);
nand UO_919 (O_919,N_19871,N_19791);
or UO_920 (O_920,N_19148,N_19759);
or UO_921 (O_921,N_19213,N_19045);
nand UO_922 (O_922,N_19431,N_19867);
nor UO_923 (O_923,N_19596,N_19823);
or UO_924 (O_924,N_19672,N_19528);
or UO_925 (O_925,N_19268,N_19783);
nor UO_926 (O_926,N_19013,N_19826);
or UO_927 (O_927,N_19311,N_19869);
nor UO_928 (O_928,N_19258,N_19477);
or UO_929 (O_929,N_19286,N_19551);
and UO_930 (O_930,N_19005,N_19218);
nor UO_931 (O_931,N_19841,N_19222);
nor UO_932 (O_932,N_19068,N_19198);
or UO_933 (O_933,N_19019,N_19890);
xnor UO_934 (O_934,N_19014,N_19500);
and UO_935 (O_935,N_19466,N_19018);
nand UO_936 (O_936,N_19529,N_19024);
and UO_937 (O_937,N_19842,N_19779);
or UO_938 (O_938,N_19702,N_19052);
nand UO_939 (O_939,N_19612,N_19999);
nand UO_940 (O_940,N_19608,N_19820);
and UO_941 (O_941,N_19800,N_19141);
nor UO_942 (O_942,N_19105,N_19477);
nand UO_943 (O_943,N_19785,N_19770);
or UO_944 (O_944,N_19272,N_19074);
nand UO_945 (O_945,N_19355,N_19161);
and UO_946 (O_946,N_19513,N_19466);
xnor UO_947 (O_947,N_19079,N_19715);
nor UO_948 (O_948,N_19716,N_19833);
nor UO_949 (O_949,N_19639,N_19706);
or UO_950 (O_950,N_19515,N_19445);
xnor UO_951 (O_951,N_19477,N_19233);
and UO_952 (O_952,N_19475,N_19694);
or UO_953 (O_953,N_19232,N_19995);
nand UO_954 (O_954,N_19585,N_19719);
nor UO_955 (O_955,N_19946,N_19235);
nand UO_956 (O_956,N_19590,N_19454);
or UO_957 (O_957,N_19573,N_19143);
nor UO_958 (O_958,N_19890,N_19970);
nand UO_959 (O_959,N_19856,N_19092);
nand UO_960 (O_960,N_19603,N_19305);
and UO_961 (O_961,N_19336,N_19664);
or UO_962 (O_962,N_19785,N_19956);
nor UO_963 (O_963,N_19258,N_19019);
xor UO_964 (O_964,N_19058,N_19300);
and UO_965 (O_965,N_19041,N_19597);
nor UO_966 (O_966,N_19457,N_19300);
and UO_967 (O_967,N_19045,N_19324);
or UO_968 (O_968,N_19379,N_19768);
or UO_969 (O_969,N_19388,N_19845);
or UO_970 (O_970,N_19211,N_19398);
and UO_971 (O_971,N_19697,N_19945);
nand UO_972 (O_972,N_19703,N_19558);
xnor UO_973 (O_973,N_19213,N_19229);
xnor UO_974 (O_974,N_19772,N_19139);
and UO_975 (O_975,N_19007,N_19241);
nand UO_976 (O_976,N_19511,N_19978);
xnor UO_977 (O_977,N_19339,N_19096);
nand UO_978 (O_978,N_19177,N_19516);
xnor UO_979 (O_979,N_19054,N_19961);
nand UO_980 (O_980,N_19532,N_19080);
and UO_981 (O_981,N_19178,N_19555);
or UO_982 (O_982,N_19886,N_19375);
nor UO_983 (O_983,N_19005,N_19119);
nor UO_984 (O_984,N_19897,N_19930);
and UO_985 (O_985,N_19956,N_19646);
xnor UO_986 (O_986,N_19028,N_19505);
and UO_987 (O_987,N_19327,N_19934);
and UO_988 (O_988,N_19044,N_19140);
nor UO_989 (O_989,N_19066,N_19807);
and UO_990 (O_990,N_19020,N_19454);
or UO_991 (O_991,N_19385,N_19506);
nand UO_992 (O_992,N_19163,N_19530);
nor UO_993 (O_993,N_19081,N_19632);
nand UO_994 (O_994,N_19653,N_19694);
and UO_995 (O_995,N_19393,N_19777);
xnor UO_996 (O_996,N_19682,N_19931);
nand UO_997 (O_997,N_19072,N_19553);
nand UO_998 (O_998,N_19643,N_19264);
and UO_999 (O_999,N_19319,N_19254);
nor UO_1000 (O_1000,N_19823,N_19632);
nor UO_1001 (O_1001,N_19957,N_19985);
xor UO_1002 (O_1002,N_19822,N_19634);
or UO_1003 (O_1003,N_19057,N_19791);
and UO_1004 (O_1004,N_19031,N_19835);
nand UO_1005 (O_1005,N_19094,N_19175);
and UO_1006 (O_1006,N_19899,N_19844);
or UO_1007 (O_1007,N_19598,N_19008);
xnor UO_1008 (O_1008,N_19144,N_19822);
nand UO_1009 (O_1009,N_19908,N_19244);
and UO_1010 (O_1010,N_19823,N_19344);
nor UO_1011 (O_1011,N_19913,N_19071);
or UO_1012 (O_1012,N_19363,N_19085);
nor UO_1013 (O_1013,N_19329,N_19453);
and UO_1014 (O_1014,N_19260,N_19778);
nor UO_1015 (O_1015,N_19991,N_19745);
and UO_1016 (O_1016,N_19011,N_19525);
and UO_1017 (O_1017,N_19367,N_19101);
or UO_1018 (O_1018,N_19364,N_19358);
and UO_1019 (O_1019,N_19557,N_19295);
or UO_1020 (O_1020,N_19055,N_19100);
nand UO_1021 (O_1021,N_19779,N_19535);
or UO_1022 (O_1022,N_19149,N_19408);
nor UO_1023 (O_1023,N_19478,N_19581);
nor UO_1024 (O_1024,N_19743,N_19593);
nor UO_1025 (O_1025,N_19317,N_19236);
nand UO_1026 (O_1026,N_19116,N_19175);
and UO_1027 (O_1027,N_19510,N_19578);
xnor UO_1028 (O_1028,N_19270,N_19728);
nand UO_1029 (O_1029,N_19000,N_19530);
and UO_1030 (O_1030,N_19498,N_19122);
xor UO_1031 (O_1031,N_19910,N_19473);
nor UO_1032 (O_1032,N_19513,N_19328);
and UO_1033 (O_1033,N_19641,N_19660);
xnor UO_1034 (O_1034,N_19888,N_19189);
or UO_1035 (O_1035,N_19915,N_19525);
or UO_1036 (O_1036,N_19112,N_19222);
or UO_1037 (O_1037,N_19868,N_19571);
xnor UO_1038 (O_1038,N_19522,N_19046);
nor UO_1039 (O_1039,N_19708,N_19186);
nand UO_1040 (O_1040,N_19048,N_19017);
nor UO_1041 (O_1041,N_19623,N_19496);
or UO_1042 (O_1042,N_19698,N_19699);
or UO_1043 (O_1043,N_19453,N_19553);
or UO_1044 (O_1044,N_19033,N_19458);
xnor UO_1045 (O_1045,N_19976,N_19561);
nand UO_1046 (O_1046,N_19030,N_19448);
nand UO_1047 (O_1047,N_19963,N_19677);
nor UO_1048 (O_1048,N_19873,N_19991);
and UO_1049 (O_1049,N_19494,N_19726);
nor UO_1050 (O_1050,N_19801,N_19442);
nor UO_1051 (O_1051,N_19259,N_19610);
or UO_1052 (O_1052,N_19042,N_19723);
nand UO_1053 (O_1053,N_19086,N_19563);
xnor UO_1054 (O_1054,N_19142,N_19660);
nand UO_1055 (O_1055,N_19912,N_19639);
or UO_1056 (O_1056,N_19678,N_19890);
nand UO_1057 (O_1057,N_19058,N_19676);
and UO_1058 (O_1058,N_19338,N_19509);
and UO_1059 (O_1059,N_19010,N_19196);
nor UO_1060 (O_1060,N_19382,N_19465);
nand UO_1061 (O_1061,N_19686,N_19369);
and UO_1062 (O_1062,N_19403,N_19079);
nand UO_1063 (O_1063,N_19412,N_19361);
nand UO_1064 (O_1064,N_19419,N_19190);
or UO_1065 (O_1065,N_19070,N_19113);
nand UO_1066 (O_1066,N_19928,N_19897);
xnor UO_1067 (O_1067,N_19517,N_19573);
xnor UO_1068 (O_1068,N_19000,N_19213);
or UO_1069 (O_1069,N_19119,N_19553);
nor UO_1070 (O_1070,N_19977,N_19680);
nor UO_1071 (O_1071,N_19897,N_19206);
or UO_1072 (O_1072,N_19712,N_19751);
and UO_1073 (O_1073,N_19154,N_19840);
and UO_1074 (O_1074,N_19773,N_19626);
nor UO_1075 (O_1075,N_19075,N_19469);
and UO_1076 (O_1076,N_19899,N_19138);
nand UO_1077 (O_1077,N_19081,N_19090);
nor UO_1078 (O_1078,N_19295,N_19160);
nand UO_1079 (O_1079,N_19656,N_19539);
nor UO_1080 (O_1080,N_19552,N_19265);
xor UO_1081 (O_1081,N_19584,N_19900);
or UO_1082 (O_1082,N_19711,N_19946);
or UO_1083 (O_1083,N_19910,N_19226);
nand UO_1084 (O_1084,N_19014,N_19522);
xnor UO_1085 (O_1085,N_19820,N_19338);
xor UO_1086 (O_1086,N_19451,N_19920);
and UO_1087 (O_1087,N_19160,N_19742);
and UO_1088 (O_1088,N_19671,N_19900);
or UO_1089 (O_1089,N_19983,N_19469);
and UO_1090 (O_1090,N_19303,N_19543);
and UO_1091 (O_1091,N_19944,N_19256);
nor UO_1092 (O_1092,N_19364,N_19354);
xnor UO_1093 (O_1093,N_19954,N_19423);
xor UO_1094 (O_1094,N_19476,N_19028);
and UO_1095 (O_1095,N_19811,N_19023);
nand UO_1096 (O_1096,N_19698,N_19959);
and UO_1097 (O_1097,N_19561,N_19526);
nand UO_1098 (O_1098,N_19319,N_19171);
nor UO_1099 (O_1099,N_19023,N_19383);
nor UO_1100 (O_1100,N_19929,N_19419);
and UO_1101 (O_1101,N_19806,N_19992);
xnor UO_1102 (O_1102,N_19042,N_19443);
xor UO_1103 (O_1103,N_19889,N_19661);
nand UO_1104 (O_1104,N_19190,N_19216);
and UO_1105 (O_1105,N_19360,N_19361);
nand UO_1106 (O_1106,N_19747,N_19551);
and UO_1107 (O_1107,N_19038,N_19074);
and UO_1108 (O_1108,N_19167,N_19114);
nor UO_1109 (O_1109,N_19440,N_19805);
and UO_1110 (O_1110,N_19603,N_19910);
or UO_1111 (O_1111,N_19537,N_19985);
nand UO_1112 (O_1112,N_19205,N_19841);
nor UO_1113 (O_1113,N_19051,N_19828);
nand UO_1114 (O_1114,N_19493,N_19325);
and UO_1115 (O_1115,N_19340,N_19587);
nand UO_1116 (O_1116,N_19353,N_19231);
xnor UO_1117 (O_1117,N_19170,N_19940);
nor UO_1118 (O_1118,N_19629,N_19903);
and UO_1119 (O_1119,N_19438,N_19247);
and UO_1120 (O_1120,N_19449,N_19558);
nor UO_1121 (O_1121,N_19622,N_19940);
nand UO_1122 (O_1122,N_19360,N_19364);
and UO_1123 (O_1123,N_19722,N_19324);
and UO_1124 (O_1124,N_19791,N_19776);
and UO_1125 (O_1125,N_19905,N_19966);
nor UO_1126 (O_1126,N_19328,N_19878);
nor UO_1127 (O_1127,N_19897,N_19329);
nor UO_1128 (O_1128,N_19603,N_19819);
xor UO_1129 (O_1129,N_19000,N_19144);
nor UO_1130 (O_1130,N_19714,N_19053);
nor UO_1131 (O_1131,N_19034,N_19429);
or UO_1132 (O_1132,N_19508,N_19007);
xor UO_1133 (O_1133,N_19821,N_19114);
nand UO_1134 (O_1134,N_19372,N_19149);
nor UO_1135 (O_1135,N_19004,N_19133);
nor UO_1136 (O_1136,N_19147,N_19443);
or UO_1137 (O_1137,N_19858,N_19760);
or UO_1138 (O_1138,N_19832,N_19713);
nor UO_1139 (O_1139,N_19398,N_19444);
nor UO_1140 (O_1140,N_19798,N_19632);
or UO_1141 (O_1141,N_19447,N_19882);
nor UO_1142 (O_1142,N_19332,N_19349);
nand UO_1143 (O_1143,N_19622,N_19954);
nor UO_1144 (O_1144,N_19505,N_19922);
and UO_1145 (O_1145,N_19162,N_19863);
nor UO_1146 (O_1146,N_19560,N_19308);
and UO_1147 (O_1147,N_19878,N_19247);
or UO_1148 (O_1148,N_19885,N_19776);
or UO_1149 (O_1149,N_19342,N_19443);
xor UO_1150 (O_1150,N_19422,N_19737);
or UO_1151 (O_1151,N_19923,N_19169);
nand UO_1152 (O_1152,N_19908,N_19751);
nand UO_1153 (O_1153,N_19292,N_19750);
nor UO_1154 (O_1154,N_19819,N_19720);
nand UO_1155 (O_1155,N_19070,N_19200);
and UO_1156 (O_1156,N_19707,N_19566);
nor UO_1157 (O_1157,N_19038,N_19652);
or UO_1158 (O_1158,N_19602,N_19724);
nand UO_1159 (O_1159,N_19596,N_19231);
and UO_1160 (O_1160,N_19175,N_19574);
nor UO_1161 (O_1161,N_19184,N_19950);
nor UO_1162 (O_1162,N_19604,N_19680);
or UO_1163 (O_1163,N_19545,N_19025);
nor UO_1164 (O_1164,N_19294,N_19688);
or UO_1165 (O_1165,N_19585,N_19504);
nand UO_1166 (O_1166,N_19865,N_19518);
or UO_1167 (O_1167,N_19044,N_19051);
nand UO_1168 (O_1168,N_19368,N_19054);
nor UO_1169 (O_1169,N_19614,N_19243);
xor UO_1170 (O_1170,N_19267,N_19036);
xnor UO_1171 (O_1171,N_19374,N_19574);
nand UO_1172 (O_1172,N_19796,N_19637);
nand UO_1173 (O_1173,N_19028,N_19229);
xor UO_1174 (O_1174,N_19433,N_19519);
nand UO_1175 (O_1175,N_19193,N_19943);
and UO_1176 (O_1176,N_19096,N_19687);
nand UO_1177 (O_1177,N_19341,N_19777);
and UO_1178 (O_1178,N_19974,N_19503);
and UO_1179 (O_1179,N_19796,N_19961);
nor UO_1180 (O_1180,N_19010,N_19388);
or UO_1181 (O_1181,N_19955,N_19349);
and UO_1182 (O_1182,N_19752,N_19351);
xnor UO_1183 (O_1183,N_19664,N_19368);
nand UO_1184 (O_1184,N_19524,N_19423);
nand UO_1185 (O_1185,N_19330,N_19640);
xnor UO_1186 (O_1186,N_19279,N_19427);
and UO_1187 (O_1187,N_19601,N_19594);
and UO_1188 (O_1188,N_19000,N_19268);
and UO_1189 (O_1189,N_19546,N_19405);
and UO_1190 (O_1190,N_19762,N_19722);
nand UO_1191 (O_1191,N_19887,N_19429);
nand UO_1192 (O_1192,N_19855,N_19650);
or UO_1193 (O_1193,N_19040,N_19337);
nand UO_1194 (O_1194,N_19589,N_19061);
nor UO_1195 (O_1195,N_19919,N_19448);
or UO_1196 (O_1196,N_19769,N_19814);
and UO_1197 (O_1197,N_19584,N_19807);
xnor UO_1198 (O_1198,N_19840,N_19357);
and UO_1199 (O_1199,N_19476,N_19645);
nor UO_1200 (O_1200,N_19071,N_19581);
or UO_1201 (O_1201,N_19869,N_19239);
nor UO_1202 (O_1202,N_19511,N_19818);
and UO_1203 (O_1203,N_19266,N_19618);
or UO_1204 (O_1204,N_19815,N_19184);
nand UO_1205 (O_1205,N_19885,N_19549);
and UO_1206 (O_1206,N_19411,N_19600);
nand UO_1207 (O_1207,N_19938,N_19493);
and UO_1208 (O_1208,N_19802,N_19436);
xnor UO_1209 (O_1209,N_19980,N_19178);
and UO_1210 (O_1210,N_19257,N_19552);
nand UO_1211 (O_1211,N_19643,N_19513);
nor UO_1212 (O_1212,N_19196,N_19153);
xor UO_1213 (O_1213,N_19442,N_19972);
or UO_1214 (O_1214,N_19678,N_19804);
nor UO_1215 (O_1215,N_19921,N_19016);
nor UO_1216 (O_1216,N_19811,N_19478);
nand UO_1217 (O_1217,N_19090,N_19466);
nor UO_1218 (O_1218,N_19641,N_19906);
nand UO_1219 (O_1219,N_19249,N_19295);
and UO_1220 (O_1220,N_19714,N_19943);
and UO_1221 (O_1221,N_19326,N_19477);
nand UO_1222 (O_1222,N_19505,N_19784);
nand UO_1223 (O_1223,N_19462,N_19800);
or UO_1224 (O_1224,N_19827,N_19690);
and UO_1225 (O_1225,N_19897,N_19344);
and UO_1226 (O_1226,N_19673,N_19337);
nand UO_1227 (O_1227,N_19001,N_19071);
or UO_1228 (O_1228,N_19941,N_19246);
nand UO_1229 (O_1229,N_19627,N_19897);
nand UO_1230 (O_1230,N_19735,N_19274);
and UO_1231 (O_1231,N_19621,N_19319);
and UO_1232 (O_1232,N_19823,N_19040);
nor UO_1233 (O_1233,N_19865,N_19061);
nor UO_1234 (O_1234,N_19877,N_19724);
nand UO_1235 (O_1235,N_19281,N_19380);
or UO_1236 (O_1236,N_19763,N_19472);
nand UO_1237 (O_1237,N_19187,N_19986);
or UO_1238 (O_1238,N_19763,N_19150);
or UO_1239 (O_1239,N_19435,N_19949);
nand UO_1240 (O_1240,N_19809,N_19050);
nor UO_1241 (O_1241,N_19607,N_19639);
nor UO_1242 (O_1242,N_19641,N_19152);
or UO_1243 (O_1243,N_19184,N_19888);
nor UO_1244 (O_1244,N_19580,N_19411);
and UO_1245 (O_1245,N_19743,N_19375);
and UO_1246 (O_1246,N_19931,N_19395);
nor UO_1247 (O_1247,N_19551,N_19542);
xor UO_1248 (O_1248,N_19241,N_19352);
and UO_1249 (O_1249,N_19898,N_19008);
or UO_1250 (O_1250,N_19421,N_19384);
or UO_1251 (O_1251,N_19431,N_19401);
or UO_1252 (O_1252,N_19710,N_19829);
nor UO_1253 (O_1253,N_19761,N_19515);
xnor UO_1254 (O_1254,N_19339,N_19850);
and UO_1255 (O_1255,N_19930,N_19739);
or UO_1256 (O_1256,N_19615,N_19573);
nor UO_1257 (O_1257,N_19019,N_19884);
nand UO_1258 (O_1258,N_19315,N_19664);
and UO_1259 (O_1259,N_19195,N_19934);
xnor UO_1260 (O_1260,N_19433,N_19059);
and UO_1261 (O_1261,N_19297,N_19950);
and UO_1262 (O_1262,N_19155,N_19656);
or UO_1263 (O_1263,N_19895,N_19176);
nand UO_1264 (O_1264,N_19495,N_19997);
nand UO_1265 (O_1265,N_19970,N_19988);
or UO_1266 (O_1266,N_19295,N_19264);
xor UO_1267 (O_1267,N_19559,N_19823);
and UO_1268 (O_1268,N_19844,N_19629);
or UO_1269 (O_1269,N_19395,N_19057);
or UO_1270 (O_1270,N_19674,N_19777);
or UO_1271 (O_1271,N_19840,N_19444);
nand UO_1272 (O_1272,N_19096,N_19114);
nor UO_1273 (O_1273,N_19826,N_19312);
and UO_1274 (O_1274,N_19299,N_19616);
and UO_1275 (O_1275,N_19607,N_19299);
nand UO_1276 (O_1276,N_19518,N_19093);
or UO_1277 (O_1277,N_19572,N_19266);
and UO_1278 (O_1278,N_19936,N_19692);
or UO_1279 (O_1279,N_19088,N_19347);
and UO_1280 (O_1280,N_19565,N_19452);
nand UO_1281 (O_1281,N_19800,N_19054);
nand UO_1282 (O_1282,N_19211,N_19365);
nand UO_1283 (O_1283,N_19827,N_19615);
or UO_1284 (O_1284,N_19109,N_19842);
nor UO_1285 (O_1285,N_19547,N_19056);
and UO_1286 (O_1286,N_19654,N_19300);
xnor UO_1287 (O_1287,N_19969,N_19447);
or UO_1288 (O_1288,N_19981,N_19074);
nand UO_1289 (O_1289,N_19080,N_19917);
nor UO_1290 (O_1290,N_19912,N_19122);
nor UO_1291 (O_1291,N_19722,N_19915);
xor UO_1292 (O_1292,N_19574,N_19163);
and UO_1293 (O_1293,N_19207,N_19457);
nand UO_1294 (O_1294,N_19000,N_19880);
nand UO_1295 (O_1295,N_19927,N_19402);
xnor UO_1296 (O_1296,N_19525,N_19823);
nand UO_1297 (O_1297,N_19091,N_19236);
nor UO_1298 (O_1298,N_19697,N_19771);
or UO_1299 (O_1299,N_19243,N_19181);
and UO_1300 (O_1300,N_19364,N_19117);
and UO_1301 (O_1301,N_19945,N_19227);
and UO_1302 (O_1302,N_19961,N_19481);
nand UO_1303 (O_1303,N_19886,N_19583);
xor UO_1304 (O_1304,N_19645,N_19731);
or UO_1305 (O_1305,N_19073,N_19146);
nand UO_1306 (O_1306,N_19119,N_19261);
and UO_1307 (O_1307,N_19985,N_19113);
nor UO_1308 (O_1308,N_19290,N_19162);
and UO_1309 (O_1309,N_19840,N_19842);
xnor UO_1310 (O_1310,N_19665,N_19503);
and UO_1311 (O_1311,N_19493,N_19268);
or UO_1312 (O_1312,N_19638,N_19755);
nand UO_1313 (O_1313,N_19976,N_19716);
and UO_1314 (O_1314,N_19584,N_19358);
or UO_1315 (O_1315,N_19806,N_19687);
xnor UO_1316 (O_1316,N_19764,N_19668);
and UO_1317 (O_1317,N_19009,N_19490);
nor UO_1318 (O_1318,N_19310,N_19304);
or UO_1319 (O_1319,N_19883,N_19455);
or UO_1320 (O_1320,N_19983,N_19443);
and UO_1321 (O_1321,N_19595,N_19091);
or UO_1322 (O_1322,N_19972,N_19489);
nor UO_1323 (O_1323,N_19515,N_19325);
xor UO_1324 (O_1324,N_19638,N_19507);
and UO_1325 (O_1325,N_19119,N_19297);
nand UO_1326 (O_1326,N_19089,N_19536);
and UO_1327 (O_1327,N_19613,N_19338);
nor UO_1328 (O_1328,N_19197,N_19262);
and UO_1329 (O_1329,N_19958,N_19967);
nand UO_1330 (O_1330,N_19345,N_19157);
nand UO_1331 (O_1331,N_19343,N_19364);
or UO_1332 (O_1332,N_19128,N_19336);
nand UO_1333 (O_1333,N_19634,N_19913);
xor UO_1334 (O_1334,N_19412,N_19422);
and UO_1335 (O_1335,N_19056,N_19257);
or UO_1336 (O_1336,N_19496,N_19719);
nor UO_1337 (O_1337,N_19930,N_19711);
xnor UO_1338 (O_1338,N_19766,N_19353);
or UO_1339 (O_1339,N_19944,N_19752);
nor UO_1340 (O_1340,N_19826,N_19261);
nor UO_1341 (O_1341,N_19062,N_19882);
or UO_1342 (O_1342,N_19295,N_19758);
and UO_1343 (O_1343,N_19772,N_19638);
nor UO_1344 (O_1344,N_19585,N_19161);
nor UO_1345 (O_1345,N_19307,N_19784);
xnor UO_1346 (O_1346,N_19601,N_19926);
nand UO_1347 (O_1347,N_19686,N_19417);
or UO_1348 (O_1348,N_19437,N_19178);
xor UO_1349 (O_1349,N_19823,N_19972);
and UO_1350 (O_1350,N_19127,N_19021);
nor UO_1351 (O_1351,N_19577,N_19682);
or UO_1352 (O_1352,N_19479,N_19480);
nand UO_1353 (O_1353,N_19285,N_19157);
xor UO_1354 (O_1354,N_19371,N_19100);
or UO_1355 (O_1355,N_19084,N_19065);
nor UO_1356 (O_1356,N_19027,N_19843);
nand UO_1357 (O_1357,N_19347,N_19586);
xnor UO_1358 (O_1358,N_19224,N_19123);
nand UO_1359 (O_1359,N_19742,N_19200);
and UO_1360 (O_1360,N_19126,N_19112);
nor UO_1361 (O_1361,N_19904,N_19483);
or UO_1362 (O_1362,N_19089,N_19485);
and UO_1363 (O_1363,N_19145,N_19781);
nand UO_1364 (O_1364,N_19868,N_19718);
nor UO_1365 (O_1365,N_19359,N_19414);
or UO_1366 (O_1366,N_19241,N_19568);
nand UO_1367 (O_1367,N_19284,N_19280);
and UO_1368 (O_1368,N_19886,N_19820);
or UO_1369 (O_1369,N_19601,N_19785);
and UO_1370 (O_1370,N_19036,N_19095);
or UO_1371 (O_1371,N_19668,N_19747);
xor UO_1372 (O_1372,N_19769,N_19555);
and UO_1373 (O_1373,N_19632,N_19360);
and UO_1374 (O_1374,N_19556,N_19584);
xnor UO_1375 (O_1375,N_19466,N_19251);
or UO_1376 (O_1376,N_19406,N_19960);
and UO_1377 (O_1377,N_19964,N_19124);
or UO_1378 (O_1378,N_19003,N_19478);
nor UO_1379 (O_1379,N_19724,N_19551);
nor UO_1380 (O_1380,N_19783,N_19135);
nand UO_1381 (O_1381,N_19722,N_19299);
nand UO_1382 (O_1382,N_19977,N_19898);
or UO_1383 (O_1383,N_19007,N_19586);
and UO_1384 (O_1384,N_19852,N_19847);
and UO_1385 (O_1385,N_19759,N_19773);
nand UO_1386 (O_1386,N_19525,N_19831);
and UO_1387 (O_1387,N_19532,N_19827);
and UO_1388 (O_1388,N_19424,N_19815);
xor UO_1389 (O_1389,N_19691,N_19705);
nand UO_1390 (O_1390,N_19527,N_19501);
or UO_1391 (O_1391,N_19031,N_19482);
and UO_1392 (O_1392,N_19379,N_19362);
or UO_1393 (O_1393,N_19897,N_19233);
nand UO_1394 (O_1394,N_19967,N_19419);
nor UO_1395 (O_1395,N_19038,N_19202);
nand UO_1396 (O_1396,N_19331,N_19414);
and UO_1397 (O_1397,N_19626,N_19599);
nor UO_1398 (O_1398,N_19516,N_19253);
nor UO_1399 (O_1399,N_19640,N_19065);
xor UO_1400 (O_1400,N_19421,N_19291);
nand UO_1401 (O_1401,N_19008,N_19939);
nand UO_1402 (O_1402,N_19068,N_19278);
nand UO_1403 (O_1403,N_19339,N_19914);
or UO_1404 (O_1404,N_19517,N_19250);
and UO_1405 (O_1405,N_19097,N_19631);
nand UO_1406 (O_1406,N_19463,N_19782);
and UO_1407 (O_1407,N_19171,N_19118);
xor UO_1408 (O_1408,N_19059,N_19789);
xnor UO_1409 (O_1409,N_19256,N_19582);
and UO_1410 (O_1410,N_19586,N_19403);
nor UO_1411 (O_1411,N_19320,N_19363);
xnor UO_1412 (O_1412,N_19159,N_19083);
nand UO_1413 (O_1413,N_19191,N_19458);
nand UO_1414 (O_1414,N_19617,N_19499);
nand UO_1415 (O_1415,N_19776,N_19554);
and UO_1416 (O_1416,N_19669,N_19445);
xnor UO_1417 (O_1417,N_19082,N_19404);
and UO_1418 (O_1418,N_19205,N_19559);
nand UO_1419 (O_1419,N_19316,N_19367);
xnor UO_1420 (O_1420,N_19998,N_19878);
nand UO_1421 (O_1421,N_19444,N_19772);
and UO_1422 (O_1422,N_19471,N_19322);
or UO_1423 (O_1423,N_19842,N_19326);
xor UO_1424 (O_1424,N_19821,N_19745);
nand UO_1425 (O_1425,N_19948,N_19240);
or UO_1426 (O_1426,N_19477,N_19979);
nor UO_1427 (O_1427,N_19399,N_19527);
or UO_1428 (O_1428,N_19230,N_19282);
and UO_1429 (O_1429,N_19593,N_19885);
nand UO_1430 (O_1430,N_19025,N_19492);
or UO_1431 (O_1431,N_19922,N_19507);
nand UO_1432 (O_1432,N_19342,N_19180);
nor UO_1433 (O_1433,N_19332,N_19459);
and UO_1434 (O_1434,N_19411,N_19694);
and UO_1435 (O_1435,N_19453,N_19332);
nand UO_1436 (O_1436,N_19555,N_19041);
nand UO_1437 (O_1437,N_19163,N_19970);
nand UO_1438 (O_1438,N_19047,N_19037);
and UO_1439 (O_1439,N_19896,N_19492);
nand UO_1440 (O_1440,N_19822,N_19969);
nand UO_1441 (O_1441,N_19737,N_19493);
nor UO_1442 (O_1442,N_19460,N_19650);
and UO_1443 (O_1443,N_19652,N_19192);
or UO_1444 (O_1444,N_19011,N_19735);
nor UO_1445 (O_1445,N_19856,N_19015);
nor UO_1446 (O_1446,N_19631,N_19493);
or UO_1447 (O_1447,N_19963,N_19902);
and UO_1448 (O_1448,N_19264,N_19730);
and UO_1449 (O_1449,N_19939,N_19116);
nand UO_1450 (O_1450,N_19265,N_19912);
nor UO_1451 (O_1451,N_19150,N_19910);
nand UO_1452 (O_1452,N_19487,N_19812);
nand UO_1453 (O_1453,N_19693,N_19463);
or UO_1454 (O_1454,N_19506,N_19943);
or UO_1455 (O_1455,N_19993,N_19943);
or UO_1456 (O_1456,N_19792,N_19338);
nor UO_1457 (O_1457,N_19011,N_19333);
xnor UO_1458 (O_1458,N_19023,N_19349);
nor UO_1459 (O_1459,N_19993,N_19574);
nand UO_1460 (O_1460,N_19654,N_19204);
xor UO_1461 (O_1461,N_19838,N_19371);
and UO_1462 (O_1462,N_19481,N_19498);
nand UO_1463 (O_1463,N_19994,N_19892);
nand UO_1464 (O_1464,N_19162,N_19195);
or UO_1465 (O_1465,N_19081,N_19146);
nand UO_1466 (O_1466,N_19789,N_19572);
nor UO_1467 (O_1467,N_19321,N_19410);
or UO_1468 (O_1468,N_19072,N_19703);
nand UO_1469 (O_1469,N_19474,N_19928);
or UO_1470 (O_1470,N_19872,N_19394);
nor UO_1471 (O_1471,N_19310,N_19676);
and UO_1472 (O_1472,N_19467,N_19870);
nor UO_1473 (O_1473,N_19771,N_19854);
xnor UO_1474 (O_1474,N_19305,N_19596);
nor UO_1475 (O_1475,N_19645,N_19121);
nor UO_1476 (O_1476,N_19591,N_19748);
xnor UO_1477 (O_1477,N_19744,N_19827);
nand UO_1478 (O_1478,N_19472,N_19929);
or UO_1479 (O_1479,N_19366,N_19561);
nor UO_1480 (O_1480,N_19222,N_19776);
xor UO_1481 (O_1481,N_19189,N_19405);
nor UO_1482 (O_1482,N_19844,N_19082);
and UO_1483 (O_1483,N_19257,N_19838);
and UO_1484 (O_1484,N_19346,N_19372);
xor UO_1485 (O_1485,N_19195,N_19006);
or UO_1486 (O_1486,N_19018,N_19095);
nand UO_1487 (O_1487,N_19205,N_19489);
nand UO_1488 (O_1488,N_19638,N_19079);
nand UO_1489 (O_1489,N_19169,N_19036);
nor UO_1490 (O_1490,N_19364,N_19757);
or UO_1491 (O_1491,N_19346,N_19255);
xor UO_1492 (O_1492,N_19980,N_19868);
nor UO_1493 (O_1493,N_19962,N_19448);
nand UO_1494 (O_1494,N_19264,N_19900);
and UO_1495 (O_1495,N_19706,N_19954);
nor UO_1496 (O_1496,N_19536,N_19036);
or UO_1497 (O_1497,N_19524,N_19358);
xnor UO_1498 (O_1498,N_19824,N_19272);
nor UO_1499 (O_1499,N_19385,N_19029);
and UO_1500 (O_1500,N_19011,N_19052);
and UO_1501 (O_1501,N_19340,N_19172);
and UO_1502 (O_1502,N_19013,N_19681);
and UO_1503 (O_1503,N_19859,N_19749);
nor UO_1504 (O_1504,N_19643,N_19763);
nand UO_1505 (O_1505,N_19079,N_19095);
and UO_1506 (O_1506,N_19888,N_19264);
and UO_1507 (O_1507,N_19540,N_19172);
nor UO_1508 (O_1508,N_19136,N_19992);
xnor UO_1509 (O_1509,N_19665,N_19825);
nor UO_1510 (O_1510,N_19586,N_19886);
nor UO_1511 (O_1511,N_19509,N_19388);
or UO_1512 (O_1512,N_19382,N_19896);
or UO_1513 (O_1513,N_19647,N_19069);
or UO_1514 (O_1514,N_19413,N_19389);
nand UO_1515 (O_1515,N_19277,N_19218);
nor UO_1516 (O_1516,N_19766,N_19826);
xor UO_1517 (O_1517,N_19484,N_19966);
or UO_1518 (O_1518,N_19356,N_19283);
xor UO_1519 (O_1519,N_19621,N_19454);
nor UO_1520 (O_1520,N_19127,N_19110);
xor UO_1521 (O_1521,N_19912,N_19002);
and UO_1522 (O_1522,N_19250,N_19681);
xor UO_1523 (O_1523,N_19416,N_19830);
and UO_1524 (O_1524,N_19913,N_19077);
nand UO_1525 (O_1525,N_19182,N_19769);
nor UO_1526 (O_1526,N_19600,N_19151);
nor UO_1527 (O_1527,N_19364,N_19671);
nand UO_1528 (O_1528,N_19567,N_19648);
nor UO_1529 (O_1529,N_19312,N_19774);
nor UO_1530 (O_1530,N_19093,N_19135);
nor UO_1531 (O_1531,N_19231,N_19093);
nor UO_1532 (O_1532,N_19447,N_19783);
xnor UO_1533 (O_1533,N_19366,N_19712);
nand UO_1534 (O_1534,N_19367,N_19872);
nand UO_1535 (O_1535,N_19345,N_19223);
nor UO_1536 (O_1536,N_19817,N_19938);
and UO_1537 (O_1537,N_19350,N_19670);
and UO_1538 (O_1538,N_19544,N_19537);
nand UO_1539 (O_1539,N_19689,N_19220);
or UO_1540 (O_1540,N_19396,N_19977);
and UO_1541 (O_1541,N_19170,N_19112);
nor UO_1542 (O_1542,N_19450,N_19855);
xor UO_1543 (O_1543,N_19946,N_19928);
and UO_1544 (O_1544,N_19749,N_19102);
nand UO_1545 (O_1545,N_19217,N_19358);
or UO_1546 (O_1546,N_19122,N_19808);
or UO_1547 (O_1547,N_19920,N_19422);
or UO_1548 (O_1548,N_19645,N_19989);
and UO_1549 (O_1549,N_19196,N_19729);
xnor UO_1550 (O_1550,N_19321,N_19567);
nand UO_1551 (O_1551,N_19248,N_19567);
nor UO_1552 (O_1552,N_19136,N_19200);
nor UO_1553 (O_1553,N_19103,N_19895);
and UO_1554 (O_1554,N_19365,N_19371);
and UO_1555 (O_1555,N_19578,N_19970);
nand UO_1556 (O_1556,N_19267,N_19937);
nor UO_1557 (O_1557,N_19878,N_19807);
and UO_1558 (O_1558,N_19501,N_19854);
nor UO_1559 (O_1559,N_19698,N_19374);
or UO_1560 (O_1560,N_19502,N_19550);
nor UO_1561 (O_1561,N_19417,N_19540);
or UO_1562 (O_1562,N_19082,N_19740);
nand UO_1563 (O_1563,N_19189,N_19320);
nor UO_1564 (O_1564,N_19296,N_19515);
nand UO_1565 (O_1565,N_19693,N_19464);
and UO_1566 (O_1566,N_19184,N_19036);
and UO_1567 (O_1567,N_19525,N_19853);
or UO_1568 (O_1568,N_19488,N_19382);
xor UO_1569 (O_1569,N_19026,N_19197);
nand UO_1570 (O_1570,N_19729,N_19365);
xnor UO_1571 (O_1571,N_19251,N_19543);
and UO_1572 (O_1572,N_19948,N_19277);
or UO_1573 (O_1573,N_19143,N_19154);
nand UO_1574 (O_1574,N_19171,N_19678);
nor UO_1575 (O_1575,N_19737,N_19351);
or UO_1576 (O_1576,N_19940,N_19571);
xor UO_1577 (O_1577,N_19291,N_19863);
xnor UO_1578 (O_1578,N_19761,N_19224);
or UO_1579 (O_1579,N_19486,N_19962);
or UO_1580 (O_1580,N_19265,N_19463);
and UO_1581 (O_1581,N_19297,N_19932);
nand UO_1582 (O_1582,N_19077,N_19821);
xnor UO_1583 (O_1583,N_19310,N_19632);
and UO_1584 (O_1584,N_19961,N_19362);
or UO_1585 (O_1585,N_19469,N_19224);
nor UO_1586 (O_1586,N_19389,N_19167);
or UO_1587 (O_1587,N_19112,N_19492);
nor UO_1588 (O_1588,N_19111,N_19877);
and UO_1589 (O_1589,N_19072,N_19067);
and UO_1590 (O_1590,N_19320,N_19049);
and UO_1591 (O_1591,N_19183,N_19784);
or UO_1592 (O_1592,N_19123,N_19584);
nand UO_1593 (O_1593,N_19427,N_19484);
and UO_1594 (O_1594,N_19565,N_19250);
xnor UO_1595 (O_1595,N_19985,N_19398);
and UO_1596 (O_1596,N_19655,N_19196);
nor UO_1597 (O_1597,N_19469,N_19130);
nand UO_1598 (O_1598,N_19494,N_19785);
nand UO_1599 (O_1599,N_19310,N_19769);
and UO_1600 (O_1600,N_19468,N_19255);
nand UO_1601 (O_1601,N_19415,N_19435);
and UO_1602 (O_1602,N_19315,N_19702);
nor UO_1603 (O_1603,N_19475,N_19338);
and UO_1604 (O_1604,N_19676,N_19508);
and UO_1605 (O_1605,N_19354,N_19602);
nand UO_1606 (O_1606,N_19037,N_19458);
or UO_1607 (O_1607,N_19124,N_19010);
and UO_1608 (O_1608,N_19192,N_19332);
nand UO_1609 (O_1609,N_19972,N_19524);
nor UO_1610 (O_1610,N_19070,N_19151);
and UO_1611 (O_1611,N_19401,N_19849);
or UO_1612 (O_1612,N_19132,N_19242);
nor UO_1613 (O_1613,N_19201,N_19567);
nand UO_1614 (O_1614,N_19211,N_19282);
or UO_1615 (O_1615,N_19265,N_19432);
xor UO_1616 (O_1616,N_19489,N_19696);
and UO_1617 (O_1617,N_19155,N_19396);
nor UO_1618 (O_1618,N_19322,N_19432);
nor UO_1619 (O_1619,N_19944,N_19986);
nand UO_1620 (O_1620,N_19245,N_19722);
and UO_1621 (O_1621,N_19057,N_19204);
and UO_1622 (O_1622,N_19951,N_19981);
and UO_1623 (O_1623,N_19883,N_19631);
xor UO_1624 (O_1624,N_19013,N_19571);
and UO_1625 (O_1625,N_19743,N_19436);
nor UO_1626 (O_1626,N_19213,N_19823);
or UO_1627 (O_1627,N_19352,N_19655);
xnor UO_1628 (O_1628,N_19621,N_19667);
or UO_1629 (O_1629,N_19929,N_19263);
nand UO_1630 (O_1630,N_19243,N_19298);
or UO_1631 (O_1631,N_19981,N_19167);
nor UO_1632 (O_1632,N_19988,N_19879);
and UO_1633 (O_1633,N_19842,N_19179);
or UO_1634 (O_1634,N_19831,N_19522);
nor UO_1635 (O_1635,N_19590,N_19852);
nand UO_1636 (O_1636,N_19510,N_19659);
nand UO_1637 (O_1637,N_19925,N_19532);
and UO_1638 (O_1638,N_19819,N_19063);
nor UO_1639 (O_1639,N_19127,N_19510);
and UO_1640 (O_1640,N_19743,N_19028);
xnor UO_1641 (O_1641,N_19759,N_19801);
and UO_1642 (O_1642,N_19178,N_19765);
or UO_1643 (O_1643,N_19937,N_19402);
xnor UO_1644 (O_1644,N_19122,N_19774);
or UO_1645 (O_1645,N_19888,N_19997);
and UO_1646 (O_1646,N_19748,N_19637);
nand UO_1647 (O_1647,N_19751,N_19998);
nand UO_1648 (O_1648,N_19454,N_19031);
nor UO_1649 (O_1649,N_19135,N_19600);
nand UO_1650 (O_1650,N_19624,N_19879);
or UO_1651 (O_1651,N_19307,N_19532);
nor UO_1652 (O_1652,N_19244,N_19949);
nor UO_1653 (O_1653,N_19126,N_19994);
and UO_1654 (O_1654,N_19086,N_19538);
nand UO_1655 (O_1655,N_19041,N_19574);
nand UO_1656 (O_1656,N_19161,N_19885);
nor UO_1657 (O_1657,N_19122,N_19214);
nor UO_1658 (O_1658,N_19283,N_19058);
nand UO_1659 (O_1659,N_19814,N_19072);
nand UO_1660 (O_1660,N_19881,N_19368);
nand UO_1661 (O_1661,N_19285,N_19992);
nand UO_1662 (O_1662,N_19733,N_19890);
and UO_1663 (O_1663,N_19589,N_19060);
nand UO_1664 (O_1664,N_19301,N_19644);
and UO_1665 (O_1665,N_19327,N_19594);
and UO_1666 (O_1666,N_19285,N_19373);
nor UO_1667 (O_1667,N_19697,N_19658);
nor UO_1668 (O_1668,N_19182,N_19860);
nand UO_1669 (O_1669,N_19749,N_19848);
nand UO_1670 (O_1670,N_19434,N_19968);
or UO_1671 (O_1671,N_19531,N_19637);
nor UO_1672 (O_1672,N_19220,N_19345);
and UO_1673 (O_1673,N_19618,N_19614);
nand UO_1674 (O_1674,N_19695,N_19140);
nand UO_1675 (O_1675,N_19598,N_19390);
or UO_1676 (O_1676,N_19859,N_19908);
nand UO_1677 (O_1677,N_19008,N_19714);
nand UO_1678 (O_1678,N_19704,N_19108);
or UO_1679 (O_1679,N_19288,N_19895);
or UO_1680 (O_1680,N_19277,N_19762);
or UO_1681 (O_1681,N_19907,N_19161);
and UO_1682 (O_1682,N_19066,N_19736);
and UO_1683 (O_1683,N_19543,N_19142);
and UO_1684 (O_1684,N_19915,N_19644);
nand UO_1685 (O_1685,N_19975,N_19252);
nand UO_1686 (O_1686,N_19412,N_19384);
and UO_1687 (O_1687,N_19424,N_19856);
nand UO_1688 (O_1688,N_19049,N_19090);
and UO_1689 (O_1689,N_19745,N_19725);
or UO_1690 (O_1690,N_19414,N_19639);
xor UO_1691 (O_1691,N_19528,N_19403);
or UO_1692 (O_1692,N_19884,N_19870);
or UO_1693 (O_1693,N_19881,N_19461);
and UO_1694 (O_1694,N_19305,N_19114);
or UO_1695 (O_1695,N_19745,N_19244);
nand UO_1696 (O_1696,N_19073,N_19691);
nor UO_1697 (O_1697,N_19453,N_19327);
nor UO_1698 (O_1698,N_19511,N_19215);
nand UO_1699 (O_1699,N_19368,N_19990);
nand UO_1700 (O_1700,N_19828,N_19996);
or UO_1701 (O_1701,N_19562,N_19686);
or UO_1702 (O_1702,N_19814,N_19686);
or UO_1703 (O_1703,N_19187,N_19713);
nand UO_1704 (O_1704,N_19887,N_19623);
or UO_1705 (O_1705,N_19107,N_19380);
nand UO_1706 (O_1706,N_19238,N_19400);
and UO_1707 (O_1707,N_19769,N_19492);
nand UO_1708 (O_1708,N_19063,N_19457);
nand UO_1709 (O_1709,N_19618,N_19236);
xor UO_1710 (O_1710,N_19906,N_19505);
and UO_1711 (O_1711,N_19889,N_19432);
nor UO_1712 (O_1712,N_19087,N_19295);
or UO_1713 (O_1713,N_19045,N_19021);
xnor UO_1714 (O_1714,N_19508,N_19478);
nand UO_1715 (O_1715,N_19937,N_19183);
and UO_1716 (O_1716,N_19227,N_19649);
and UO_1717 (O_1717,N_19161,N_19813);
xnor UO_1718 (O_1718,N_19266,N_19280);
xor UO_1719 (O_1719,N_19966,N_19911);
nand UO_1720 (O_1720,N_19859,N_19465);
or UO_1721 (O_1721,N_19505,N_19676);
nand UO_1722 (O_1722,N_19730,N_19217);
nand UO_1723 (O_1723,N_19662,N_19976);
nor UO_1724 (O_1724,N_19812,N_19659);
or UO_1725 (O_1725,N_19613,N_19585);
nor UO_1726 (O_1726,N_19826,N_19160);
or UO_1727 (O_1727,N_19490,N_19715);
nor UO_1728 (O_1728,N_19078,N_19330);
nand UO_1729 (O_1729,N_19302,N_19853);
or UO_1730 (O_1730,N_19917,N_19054);
or UO_1731 (O_1731,N_19887,N_19901);
or UO_1732 (O_1732,N_19260,N_19002);
nand UO_1733 (O_1733,N_19439,N_19052);
nor UO_1734 (O_1734,N_19521,N_19928);
and UO_1735 (O_1735,N_19040,N_19474);
xor UO_1736 (O_1736,N_19575,N_19898);
nand UO_1737 (O_1737,N_19417,N_19823);
nor UO_1738 (O_1738,N_19872,N_19028);
or UO_1739 (O_1739,N_19522,N_19025);
and UO_1740 (O_1740,N_19713,N_19072);
nor UO_1741 (O_1741,N_19479,N_19968);
or UO_1742 (O_1742,N_19976,N_19081);
xnor UO_1743 (O_1743,N_19261,N_19767);
nand UO_1744 (O_1744,N_19470,N_19944);
or UO_1745 (O_1745,N_19083,N_19874);
nand UO_1746 (O_1746,N_19029,N_19439);
nand UO_1747 (O_1747,N_19266,N_19708);
nand UO_1748 (O_1748,N_19339,N_19265);
nand UO_1749 (O_1749,N_19966,N_19374);
nand UO_1750 (O_1750,N_19194,N_19755);
xor UO_1751 (O_1751,N_19753,N_19547);
nor UO_1752 (O_1752,N_19050,N_19046);
and UO_1753 (O_1753,N_19939,N_19076);
and UO_1754 (O_1754,N_19225,N_19481);
and UO_1755 (O_1755,N_19982,N_19867);
or UO_1756 (O_1756,N_19164,N_19114);
nor UO_1757 (O_1757,N_19439,N_19950);
nor UO_1758 (O_1758,N_19500,N_19488);
nor UO_1759 (O_1759,N_19800,N_19916);
or UO_1760 (O_1760,N_19884,N_19951);
and UO_1761 (O_1761,N_19853,N_19118);
and UO_1762 (O_1762,N_19571,N_19552);
and UO_1763 (O_1763,N_19284,N_19918);
or UO_1764 (O_1764,N_19678,N_19222);
nand UO_1765 (O_1765,N_19737,N_19903);
or UO_1766 (O_1766,N_19545,N_19066);
nor UO_1767 (O_1767,N_19210,N_19880);
nor UO_1768 (O_1768,N_19185,N_19274);
nand UO_1769 (O_1769,N_19040,N_19168);
nand UO_1770 (O_1770,N_19960,N_19254);
or UO_1771 (O_1771,N_19097,N_19745);
or UO_1772 (O_1772,N_19844,N_19951);
nand UO_1773 (O_1773,N_19080,N_19299);
or UO_1774 (O_1774,N_19876,N_19887);
nand UO_1775 (O_1775,N_19268,N_19639);
or UO_1776 (O_1776,N_19773,N_19100);
xor UO_1777 (O_1777,N_19950,N_19088);
nor UO_1778 (O_1778,N_19091,N_19825);
nand UO_1779 (O_1779,N_19902,N_19420);
nor UO_1780 (O_1780,N_19588,N_19812);
or UO_1781 (O_1781,N_19790,N_19329);
or UO_1782 (O_1782,N_19994,N_19350);
and UO_1783 (O_1783,N_19095,N_19659);
nor UO_1784 (O_1784,N_19426,N_19808);
nor UO_1785 (O_1785,N_19734,N_19430);
xor UO_1786 (O_1786,N_19034,N_19283);
or UO_1787 (O_1787,N_19790,N_19639);
nor UO_1788 (O_1788,N_19814,N_19209);
nor UO_1789 (O_1789,N_19934,N_19342);
and UO_1790 (O_1790,N_19010,N_19465);
or UO_1791 (O_1791,N_19858,N_19875);
and UO_1792 (O_1792,N_19397,N_19529);
nor UO_1793 (O_1793,N_19839,N_19538);
nand UO_1794 (O_1794,N_19914,N_19031);
and UO_1795 (O_1795,N_19316,N_19491);
nor UO_1796 (O_1796,N_19518,N_19530);
nand UO_1797 (O_1797,N_19103,N_19298);
and UO_1798 (O_1798,N_19716,N_19766);
nand UO_1799 (O_1799,N_19955,N_19562);
xnor UO_1800 (O_1800,N_19119,N_19821);
xnor UO_1801 (O_1801,N_19803,N_19122);
nand UO_1802 (O_1802,N_19564,N_19291);
nor UO_1803 (O_1803,N_19313,N_19674);
and UO_1804 (O_1804,N_19344,N_19926);
or UO_1805 (O_1805,N_19831,N_19858);
nand UO_1806 (O_1806,N_19211,N_19478);
nand UO_1807 (O_1807,N_19049,N_19333);
or UO_1808 (O_1808,N_19074,N_19747);
xnor UO_1809 (O_1809,N_19858,N_19043);
or UO_1810 (O_1810,N_19382,N_19874);
or UO_1811 (O_1811,N_19901,N_19024);
or UO_1812 (O_1812,N_19301,N_19473);
and UO_1813 (O_1813,N_19378,N_19868);
nor UO_1814 (O_1814,N_19640,N_19676);
nor UO_1815 (O_1815,N_19764,N_19138);
or UO_1816 (O_1816,N_19375,N_19986);
or UO_1817 (O_1817,N_19682,N_19157);
and UO_1818 (O_1818,N_19272,N_19342);
nand UO_1819 (O_1819,N_19040,N_19531);
and UO_1820 (O_1820,N_19389,N_19949);
nand UO_1821 (O_1821,N_19044,N_19830);
xor UO_1822 (O_1822,N_19225,N_19664);
or UO_1823 (O_1823,N_19894,N_19633);
nand UO_1824 (O_1824,N_19863,N_19436);
nand UO_1825 (O_1825,N_19226,N_19343);
nand UO_1826 (O_1826,N_19631,N_19869);
nand UO_1827 (O_1827,N_19997,N_19498);
nand UO_1828 (O_1828,N_19876,N_19744);
nor UO_1829 (O_1829,N_19623,N_19258);
nand UO_1830 (O_1830,N_19651,N_19294);
and UO_1831 (O_1831,N_19168,N_19148);
nand UO_1832 (O_1832,N_19443,N_19848);
xnor UO_1833 (O_1833,N_19544,N_19026);
xor UO_1834 (O_1834,N_19576,N_19656);
nor UO_1835 (O_1835,N_19162,N_19452);
and UO_1836 (O_1836,N_19551,N_19838);
and UO_1837 (O_1837,N_19968,N_19212);
or UO_1838 (O_1838,N_19377,N_19497);
nor UO_1839 (O_1839,N_19592,N_19405);
nand UO_1840 (O_1840,N_19312,N_19599);
or UO_1841 (O_1841,N_19742,N_19900);
or UO_1842 (O_1842,N_19150,N_19560);
xor UO_1843 (O_1843,N_19608,N_19656);
and UO_1844 (O_1844,N_19604,N_19192);
nand UO_1845 (O_1845,N_19852,N_19139);
xor UO_1846 (O_1846,N_19977,N_19710);
nand UO_1847 (O_1847,N_19889,N_19031);
nand UO_1848 (O_1848,N_19190,N_19533);
nor UO_1849 (O_1849,N_19235,N_19182);
nor UO_1850 (O_1850,N_19100,N_19917);
nand UO_1851 (O_1851,N_19491,N_19371);
and UO_1852 (O_1852,N_19677,N_19967);
nand UO_1853 (O_1853,N_19284,N_19447);
nor UO_1854 (O_1854,N_19219,N_19531);
and UO_1855 (O_1855,N_19290,N_19600);
nor UO_1856 (O_1856,N_19471,N_19110);
or UO_1857 (O_1857,N_19782,N_19075);
nor UO_1858 (O_1858,N_19559,N_19682);
or UO_1859 (O_1859,N_19957,N_19959);
nand UO_1860 (O_1860,N_19964,N_19414);
nand UO_1861 (O_1861,N_19378,N_19202);
or UO_1862 (O_1862,N_19043,N_19966);
nor UO_1863 (O_1863,N_19864,N_19825);
and UO_1864 (O_1864,N_19916,N_19943);
xnor UO_1865 (O_1865,N_19045,N_19272);
or UO_1866 (O_1866,N_19106,N_19516);
nand UO_1867 (O_1867,N_19514,N_19523);
nand UO_1868 (O_1868,N_19469,N_19348);
xor UO_1869 (O_1869,N_19573,N_19886);
or UO_1870 (O_1870,N_19590,N_19755);
nor UO_1871 (O_1871,N_19858,N_19665);
nor UO_1872 (O_1872,N_19553,N_19077);
xor UO_1873 (O_1873,N_19946,N_19603);
or UO_1874 (O_1874,N_19892,N_19822);
xnor UO_1875 (O_1875,N_19498,N_19986);
or UO_1876 (O_1876,N_19747,N_19774);
and UO_1877 (O_1877,N_19848,N_19065);
nand UO_1878 (O_1878,N_19141,N_19312);
or UO_1879 (O_1879,N_19428,N_19696);
and UO_1880 (O_1880,N_19105,N_19084);
and UO_1881 (O_1881,N_19099,N_19688);
nor UO_1882 (O_1882,N_19734,N_19163);
nand UO_1883 (O_1883,N_19547,N_19310);
xor UO_1884 (O_1884,N_19911,N_19865);
nor UO_1885 (O_1885,N_19374,N_19845);
nor UO_1886 (O_1886,N_19369,N_19749);
and UO_1887 (O_1887,N_19397,N_19913);
and UO_1888 (O_1888,N_19666,N_19665);
nand UO_1889 (O_1889,N_19447,N_19232);
nand UO_1890 (O_1890,N_19963,N_19262);
nand UO_1891 (O_1891,N_19748,N_19093);
nand UO_1892 (O_1892,N_19684,N_19743);
nor UO_1893 (O_1893,N_19460,N_19779);
or UO_1894 (O_1894,N_19833,N_19862);
nor UO_1895 (O_1895,N_19634,N_19786);
nand UO_1896 (O_1896,N_19134,N_19570);
nand UO_1897 (O_1897,N_19481,N_19916);
nand UO_1898 (O_1898,N_19681,N_19867);
and UO_1899 (O_1899,N_19813,N_19015);
or UO_1900 (O_1900,N_19011,N_19683);
nor UO_1901 (O_1901,N_19661,N_19688);
nand UO_1902 (O_1902,N_19018,N_19376);
nand UO_1903 (O_1903,N_19347,N_19141);
xor UO_1904 (O_1904,N_19588,N_19303);
and UO_1905 (O_1905,N_19935,N_19791);
or UO_1906 (O_1906,N_19671,N_19028);
nor UO_1907 (O_1907,N_19356,N_19105);
or UO_1908 (O_1908,N_19146,N_19682);
nor UO_1909 (O_1909,N_19267,N_19979);
nand UO_1910 (O_1910,N_19060,N_19179);
or UO_1911 (O_1911,N_19086,N_19513);
nor UO_1912 (O_1912,N_19638,N_19373);
nand UO_1913 (O_1913,N_19525,N_19053);
and UO_1914 (O_1914,N_19733,N_19738);
nand UO_1915 (O_1915,N_19219,N_19611);
or UO_1916 (O_1916,N_19904,N_19913);
and UO_1917 (O_1917,N_19711,N_19416);
nor UO_1918 (O_1918,N_19922,N_19039);
nand UO_1919 (O_1919,N_19891,N_19980);
nand UO_1920 (O_1920,N_19209,N_19085);
xor UO_1921 (O_1921,N_19160,N_19967);
or UO_1922 (O_1922,N_19303,N_19032);
and UO_1923 (O_1923,N_19774,N_19627);
nand UO_1924 (O_1924,N_19950,N_19003);
xor UO_1925 (O_1925,N_19610,N_19155);
or UO_1926 (O_1926,N_19328,N_19777);
and UO_1927 (O_1927,N_19260,N_19540);
xnor UO_1928 (O_1928,N_19692,N_19431);
xor UO_1929 (O_1929,N_19752,N_19797);
and UO_1930 (O_1930,N_19854,N_19452);
nor UO_1931 (O_1931,N_19160,N_19692);
nor UO_1932 (O_1932,N_19694,N_19754);
and UO_1933 (O_1933,N_19083,N_19854);
or UO_1934 (O_1934,N_19849,N_19538);
or UO_1935 (O_1935,N_19961,N_19223);
nand UO_1936 (O_1936,N_19171,N_19747);
nor UO_1937 (O_1937,N_19821,N_19791);
or UO_1938 (O_1938,N_19720,N_19886);
xnor UO_1939 (O_1939,N_19907,N_19244);
nand UO_1940 (O_1940,N_19858,N_19654);
nor UO_1941 (O_1941,N_19126,N_19695);
nand UO_1942 (O_1942,N_19760,N_19761);
and UO_1943 (O_1943,N_19855,N_19145);
nor UO_1944 (O_1944,N_19608,N_19645);
and UO_1945 (O_1945,N_19391,N_19078);
xnor UO_1946 (O_1946,N_19936,N_19376);
nand UO_1947 (O_1947,N_19851,N_19163);
or UO_1948 (O_1948,N_19875,N_19924);
or UO_1949 (O_1949,N_19431,N_19332);
and UO_1950 (O_1950,N_19455,N_19695);
nand UO_1951 (O_1951,N_19111,N_19666);
and UO_1952 (O_1952,N_19289,N_19924);
or UO_1953 (O_1953,N_19908,N_19258);
and UO_1954 (O_1954,N_19909,N_19355);
nand UO_1955 (O_1955,N_19810,N_19199);
or UO_1956 (O_1956,N_19296,N_19934);
nand UO_1957 (O_1957,N_19203,N_19416);
nand UO_1958 (O_1958,N_19695,N_19453);
and UO_1959 (O_1959,N_19299,N_19656);
or UO_1960 (O_1960,N_19143,N_19941);
or UO_1961 (O_1961,N_19104,N_19869);
and UO_1962 (O_1962,N_19248,N_19207);
nor UO_1963 (O_1963,N_19130,N_19194);
nor UO_1964 (O_1964,N_19724,N_19467);
and UO_1965 (O_1965,N_19438,N_19678);
and UO_1966 (O_1966,N_19047,N_19915);
and UO_1967 (O_1967,N_19162,N_19928);
and UO_1968 (O_1968,N_19634,N_19194);
nor UO_1969 (O_1969,N_19629,N_19701);
and UO_1970 (O_1970,N_19969,N_19905);
and UO_1971 (O_1971,N_19012,N_19985);
xnor UO_1972 (O_1972,N_19212,N_19638);
xor UO_1973 (O_1973,N_19441,N_19180);
and UO_1974 (O_1974,N_19709,N_19833);
and UO_1975 (O_1975,N_19049,N_19958);
nor UO_1976 (O_1976,N_19280,N_19667);
and UO_1977 (O_1977,N_19966,N_19530);
nand UO_1978 (O_1978,N_19307,N_19498);
xor UO_1979 (O_1979,N_19516,N_19128);
and UO_1980 (O_1980,N_19417,N_19362);
xor UO_1981 (O_1981,N_19651,N_19971);
xnor UO_1982 (O_1982,N_19080,N_19513);
or UO_1983 (O_1983,N_19236,N_19786);
and UO_1984 (O_1984,N_19564,N_19190);
nand UO_1985 (O_1985,N_19558,N_19968);
nand UO_1986 (O_1986,N_19112,N_19801);
xor UO_1987 (O_1987,N_19990,N_19214);
xnor UO_1988 (O_1988,N_19793,N_19908);
and UO_1989 (O_1989,N_19266,N_19957);
nor UO_1990 (O_1990,N_19632,N_19760);
or UO_1991 (O_1991,N_19943,N_19615);
nor UO_1992 (O_1992,N_19673,N_19045);
nor UO_1993 (O_1993,N_19831,N_19050);
and UO_1994 (O_1994,N_19291,N_19636);
and UO_1995 (O_1995,N_19146,N_19493);
nand UO_1996 (O_1996,N_19762,N_19030);
xor UO_1997 (O_1997,N_19123,N_19333);
xor UO_1998 (O_1998,N_19499,N_19968);
or UO_1999 (O_1999,N_19750,N_19441);
and UO_2000 (O_2000,N_19058,N_19697);
and UO_2001 (O_2001,N_19794,N_19941);
and UO_2002 (O_2002,N_19143,N_19207);
or UO_2003 (O_2003,N_19560,N_19857);
or UO_2004 (O_2004,N_19416,N_19231);
xor UO_2005 (O_2005,N_19717,N_19792);
or UO_2006 (O_2006,N_19228,N_19331);
or UO_2007 (O_2007,N_19192,N_19915);
or UO_2008 (O_2008,N_19832,N_19068);
and UO_2009 (O_2009,N_19928,N_19160);
and UO_2010 (O_2010,N_19232,N_19390);
nor UO_2011 (O_2011,N_19071,N_19249);
and UO_2012 (O_2012,N_19063,N_19195);
nor UO_2013 (O_2013,N_19996,N_19843);
or UO_2014 (O_2014,N_19634,N_19187);
nand UO_2015 (O_2015,N_19253,N_19043);
nor UO_2016 (O_2016,N_19483,N_19262);
and UO_2017 (O_2017,N_19775,N_19756);
nand UO_2018 (O_2018,N_19236,N_19277);
nand UO_2019 (O_2019,N_19748,N_19082);
xnor UO_2020 (O_2020,N_19330,N_19311);
or UO_2021 (O_2021,N_19804,N_19009);
and UO_2022 (O_2022,N_19448,N_19032);
xnor UO_2023 (O_2023,N_19354,N_19010);
nand UO_2024 (O_2024,N_19584,N_19919);
nand UO_2025 (O_2025,N_19590,N_19875);
or UO_2026 (O_2026,N_19294,N_19275);
nor UO_2027 (O_2027,N_19773,N_19383);
xnor UO_2028 (O_2028,N_19850,N_19649);
nand UO_2029 (O_2029,N_19487,N_19676);
or UO_2030 (O_2030,N_19432,N_19379);
and UO_2031 (O_2031,N_19258,N_19099);
xor UO_2032 (O_2032,N_19032,N_19710);
or UO_2033 (O_2033,N_19851,N_19720);
nand UO_2034 (O_2034,N_19815,N_19112);
nand UO_2035 (O_2035,N_19874,N_19726);
xor UO_2036 (O_2036,N_19321,N_19793);
xnor UO_2037 (O_2037,N_19240,N_19995);
nand UO_2038 (O_2038,N_19448,N_19708);
nand UO_2039 (O_2039,N_19279,N_19448);
and UO_2040 (O_2040,N_19173,N_19461);
nor UO_2041 (O_2041,N_19709,N_19923);
nand UO_2042 (O_2042,N_19524,N_19518);
and UO_2043 (O_2043,N_19165,N_19635);
nand UO_2044 (O_2044,N_19479,N_19990);
nor UO_2045 (O_2045,N_19263,N_19442);
nor UO_2046 (O_2046,N_19112,N_19330);
xor UO_2047 (O_2047,N_19880,N_19466);
nand UO_2048 (O_2048,N_19241,N_19213);
xnor UO_2049 (O_2049,N_19313,N_19652);
nor UO_2050 (O_2050,N_19885,N_19529);
xnor UO_2051 (O_2051,N_19789,N_19680);
and UO_2052 (O_2052,N_19429,N_19739);
or UO_2053 (O_2053,N_19516,N_19167);
nor UO_2054 (O_2054,N_19105,N_19836);
and UO_2055 (O_2055,N_19808,N_19367);
or UO_2056 (O_2056,N_19682,N_19105);
nand UO_2057 (O_2057,N_19093,N_19583);
and UO_2058 (O_2058,N_19555,N_19930);
or UO_2059 (O_2059,N_19589,N_19028);
and UO_2060 (O_2060,N_19719,N_19768);
or UO_2061 (O_2061,N_19250,N_19729);
and UO_2062 (O_2062,N_19556,N_19615);
or UO_2063 (O_2063,N_19245,N_19310);
or UO_2064 (O_2064,N_19169,N_19297);
nor UO_2065 (O_2065,N_19067,N_19224);
or UO_2066 (O_2066,N_19717,N_19621);
nor UO_2067 (O_2067,N_19098,N_19102);
xnor UO_2068 (O_2068,N_19860,N_19016);
nor UO_2069 (O_2069,N_19317,N_19898);
nor UO_2070 (O_2070,N_19984,N_19879);
or UO_2071 (O_2071,N_19985,N_19519);
xnor UO_2072 (O_2072,N_19532,N_19738);
nor UO_2073 (O_2073,N_19636,N_19630);
or UO_2074 (O_2074,N_19284,N_19019);
and UO_2075 (O_2075,N_19388,N_19438);
nor UO_2076 (O_2076,N_19304,N_19525);
xnor UO_2077 (O_2077,N_19440,N_19909);
xnor UO_2078 (O_2078,N_19501,N_19662);
nand UO_2079 (O_2079,N_19159,N_19840);
or UO_2080 (O_2080,N_19668,N_19657);
and UO_2081 (O_2081,N_19847,N_19199);
nor UO_2082 (O_2082,N_19914,N_19367);
or UO_2083 (O_2083,N_19343,N_19455);
and UO_2084 (O_2084,N_19470,N_19818);
nor UO_2085 (O_2085,N_19815,N_19256);
or UO_2086 (O_2086,N_19737,N_19999);
nor UO_2087 (O_2087,N_19315,N_19353);
xnor UO_2088 (O_2088,N_19315,N_19492);
and UO_2089 (O_2089,N_19016,N_19442);
nand UO_2090 (O_2090,N_19488,N_19813);
nor UO_2091 (O_2091,N_19057,N_19139);
nand UO_2092 (O_2092,N_19217,N_19232);
or UO_2093 (O_2093,N_19379,N_19436);
xor UO_2094 (O_2094,N_19172,N_19738);
or UO_2095 (O_2095,N_19349,N_19203);
nor UO_2096 (O_2096,N_19073,N_19493);
nor UO_2097 (O_2097,N_19215,N_19724);
nor UO_2098 (O_2098,N_19513,N_19209);
or UO_2099 (O_2099,N_19448,N_19300);
nand UO_2100 (O_2100,N_19089,N_19383);
or UO_2101 (O_2101,N_19762,N_19468);
nor UO_2102 (O_2102,N_19171,N_19776);
nor UO_2103 (O_2103,N_19459,N_19961);
nand UO_2104 (O_2104,N_19694,N_19039);
or UO_2105 (O_2105,N_19922,N_19275);
nand UO_2106 (O_2106,N_19088,N_19219);
nor UO_2107 (O_2107,N_19284,N_19147);
nor UO_2108 (O_2108,N_19716,N_19747);
and UO_2109 (O_2109,N_19327,N_19787);
and UO_2110 (O_2110,N_19394,N_19530);
or UO_2111 (O_2111,N_19308,N_19417);
nand UO_2112 (O_2112,N_19900,N_19145);
and UO_2113 (O_2113,N_19344,N_19000);
and UO_2114 (O_2114,N_19470,N_19984);
or UO_2115 (O_2115,N_19881,N_19084);
or UO_2116 (O_2116,N_19951,N_19865);
or UO_2117 (O_2117,N_19404,N_19365);
and UO_2118 (O_2118,N_19846,N_19679);
or UO_2119 (O_2119,N_19910,N_19364);
and UO_2120 (O_2120,N_19814,N_19702);
and UO_2121 (O_2121,N_19918,N_19293);
or UO_2122 (O_2122,N_19612,N_19851);
nor UO_2123 (O_2123,N_19897,N_19508);
and UO_2124 (O_2124,N_19382,N_19437);
or UO_2125 (O_2125,N_19013,N_19574);
nor UO_2126 (O_2126,N_19871,N_19500);
nor UO_2127 (O_2127,N_19031,N_19281);
nand UO_2128 (O_2128,N_19273,N_19502);
or UO_2129 (O_2129,N_19943,N_19829);
or UO_2130 (O_2130,N_19578,N_19178);
nor UO_2131 (O_2131,N_19981,N_19533);
and UO_2132 (O_2132,N_19257,N_19667);
and UO_2133 (O_2133,N_19302,N_19392);
nand UO_2134 (O_2134,N_19922,N_19897);
and UO_2135 (O_2135,N_19718,N_19984);
nand UO_2136 (O_2136,N_19789,N_19569);
or UO_2137 (O_2137,N_19017,N_19898);
and UO_2138 (O_2138,N_19786,N_19154);
xor UO_2139 (O_2139,N_19005,N_19600);
nand UO_2140 (O_2140,N_19389,N_19269);
and UO_2141 (O_2141,N_19501,N_19563);
or UO_2142 (O_2142,N_19057,N_19346);
and UO_2143 (O_2143,N_19599,N_19341);
nor UO_2144 (O_2144,N_19462,N_19197);
and UO_2145 (O_2145,N_19695,N_19614);
and UO_2146 (O_2146,N_19332,N_19917);
nand UO_2147 (O_2147,N_19608,N_19416);
nand UO_2148 (O_2148,N_19099,N_19213);
or UO_2149 (O_2149,N_19006,N_19223);
nor UO_2150 (O_2150,N_19679,N_19395);
and UO_2151 (O_2151,N_19854,N_19446);
or UO_2152 (O_2152,N_19131,N_19050);
nor UO_2153 (O_2153,N_19026,N_19317);
nor UO_2154 (O_2154,N_19297,N_19981);
or UO_2155 (O_2155,N_19234,N_19129);
nor UO_2156 (O_2156,N_19063,N_19112);
and UO_2157 (O_2157,N_19831,N_19312);
nand UO_2158 (O_2158,N_19882,N_19695);
nor UO_2159 (O_2159,N_19617,N_19231);
and UO_2160 (O_2160,N_19307,N_19270);
xor UO_2161 (O_2161,N_19744,N_19973);
nor UO_2162 (O_2162,N_19057,N_19593);
and UO_2163 (O_2163,N_19235,N_19785);
and UO_2164 (O_2164,N_19453,N_19260);
nand UO_2165 (O_2165,N_19489,N_19114);
or UO_2166 (O_2166,N_19776,N_19060);
or UO_2167 (O_2167,N_19295,N_19541);
nor UO_2168 (O_2168,N_19737,N_19374);
nor UO_2169 (O_2169,N_19235,N_19096);
nor UO_2170 (O_2170,N_19930,N_19276);
nand UO_2171 (O_2171,N_19721,N_19121);
nor UO_2172 (O_2172,N_19907,N_19338);
xnor UO_2173 (O_2173,N_19212,N_19276);
nand UO_2174 (O_2174,N_19090,N_19924);
and UO_2175 (O_2175,N_19587,N_19885);
xor UO_2176 (O_2176,N_19601,N_19560);
nor UO_2177 (O_2177,N_19786,N_19848);
nand UO_2178 (O_2178,N_19629,N_19673);
or UO_2179 (O_2179,N_19611,N_19999);
or UO_2180 (O_2180,N_19370,N_19184);
and UO_2181 (O_2181,N_19180,N_19348);
or UO_2182 (O_2182,N_19671,N_19227);
nor UO_2183 (O_2183,N_19862,N_19515);
nand UO_2184 (O_2184,N_19851,N_19697);
nand UO_2185 (O_2185,N_19430,N_19071);
nand UO_2186 (O_2186,N_19309,N_19484);
nor UO_2187 (O_2187,N_19396,N_19622);
and UO_2188 (O_2188,N_19945,N_19066);
or UO_2189 (O_2189,N_19137,N_19800);
and UO_2190 (O_2190,N_19530,N_19531);
nand UO_2191 (O_2191,N_19329,N_19301);
and UO_2192 (O_2192,N_19140,N_19272);
or UO_2193 (O_2193,N_19545,N_19574);
or UO_2194 (O_2194,N_19719,N_19518);
or UO_2195 (O_2195,N_19733,N_19988);
and UO_2196 (O_2196,N_19204,N_19880);
nand UO_2197 (O_2197,N_19420,N_19864);
or UO_2198 (O_2198,N_19456,N_19016);
and UO_2199 (O_2199,N_19320,N_19644);
nor UO_2200 (O_2200,N_19565,N_19577);
or UO_2201 (O_2201,N_19613,N_19788);
xnor UO_2202 (O_2202,N_19986,N_19010);
xor UO_2203 (O_2203,N_19603,N_19730);
nor UO_2204 (O_2204,N_19785,N_19013);
and UO_2205 (O_2205,N_19527,N_19384);
nor UO_2206 (O_2206,N_19954,N_19503);
nor UO_2207 (O_2207,N_19084,N_19614);
and UO_2208 (O_2208,N_19353,N_19424);
or UO_2209 (O_2209,N_19095,N_19843);
nand UO_2210 (O_2210,N_19748,N_19946);
or UO_2211 (O_2211,N_19797,N_19266);
nor UO_2212 (O_2212,N_19279,N_19335);
and UO_2213 (O_2213,N_19242,N_19944);
and UO_2214 (O_2214,N_19355,N_19633);
and UO_2215 (O_2215,N_19910,N_19527);
xnor UO_2216 (O_2216,N_19310,N_19102);
and UO_2217 (O_2217,N_19292,N_19489);
nand UO_2218 (O_2218,N_19711,N_19027);
nand UO_2219 (O_2219,N_19910,N_19352);
nor UO_2220 (O_2220,N_19523,N_19037);
or UO_2221 (O_2221,N_19726,N_19054);
nor UO_2222 (O_2222,N_19341,N_19942);
nor UO_2223 (O_2223,N_19890,N_19441);
or UO_2224 (O_2224,N_19979,N_19592);
and UO_2225 (O_2225,N_19186,N_19798);
nand UO_2226 (O_2226,N_19329,N_19183);
nor UO_2227 (O_2227,N_19479,N_19535);
or UO_2228 (O_2228,N_19687,N_19090);
nand UO_2229 (O_2229,N_19048,N_19557);
nor UO_2230 (O_2230,N_19085,N_19036);
or UO_2231 (O_2231,N_19599,N_19168);
nand UO_2232 (O_2232,N_19600,N_19559);
or UO_2233 (O_2233,N_19988,N_19207);
nor UO_2234 (O_2234,N_19746,N_19520);
nand UO_2235 (O_2235,N_19803,N_19038);
or UO_2236 (O_2236,N_19140,N_19493);
nand UO_2237 (O_2237,N_19934,N_19031);
or UO_2238 (O_2238,N_19111,N_19054);
and UO_2239 (O_2239,N_19868,N_19001);
nand UO_2240 (O_2240,N_19692,N_19596);
or UO_2241 (O_2241,N_19689,N_19081);
nor UO_2242 (O_2242,N_19088,N_19959);
nor UO_2243 (O_2243,N_19654,N_19458);
or UO_2244 (O_2244,N_19769,N_19802);
and UO_2245 (O_2245,N_19594,N_19778);
and UO_2246 (O_2246,N_19334,N_19043);
nand UO_2247 (O_2247,N_19588,N_19010);
nor UO_2248 (O_2248,N_19975,N_19759);
xnor UO_2249 (O_2249,N_19581,N_19045);
and UO_2250 (O_2250,N_19893,N_19283);
nor UO_2251 (O_2251,N_19977,N_19653);
or UO_2252 (O_2252,N_19337,N_19085);
nor UO_2253 (O_2253,N_19372,N_19133);
or UO_2254 (O_2254,N_19722,N_19032);
nor UO_2255 (O_2255,N_19742,N_19158);
nand UO_2256 (O_2256,N_19125,N_19573);
and UO_2257 (O_2257,N_19092,N_19531);
or UO_2258 (O_2258,N_19864,N_19223);
nand UO_2259 (O_2259,N_19124,N_19521);
nor UO_2260 (O_2260,N_19533,N_19032);
and UO_2261 (O_2261,N_19753,N_19876);
nor UO_2262 (O_2262,N_19821,N_19544);
nand UO_2263 (O_2263,N_19057,N_19012);
nand UO_2264 (O_2264,N_19270,N_19695);
and UO_2265 (O_2265,N_19836,N_19967);
nand UO_2266 (O_2266,N_19290,N_19816);
and UO_2267 (O_2267,N_19894,N_19595);
nor UO_2268 (O_2268,N_19417,N_19410);
xnor UO_2269 (O_2269,N_19474,N_19706);
or UO_2270 (O_2270,N_19209,N_19033);
and UO_2271 (O_2271,N_19259,N_19106);
nor UO_2272 (O_2272,N_19437,N_19397);
nor UO_2273 (O_2273,N_19111,N_19951);
nand UO_2274 (O_2274,N_19216,N_19151);
xnor UO_2275 (O_2275,N_19292,N_19231);
nor UO_2276 (O_2276,N_19242,N_19037);
or UO_2277 (O_2277,N_19980,N_19304);
nand UO_2278 (O_2278,N_19408,N_19661);
nor UO_2279 (O_2279,N_19609,N_19992);
or UO_2280 (O_2280,N_19102,N_19038);
and UO_2281 (O_2281,N_19933,N_19047);
and UO_2282 (O_2282,N_19504,N_19559);
xnor UO_2283 (O_2283,N_19296,N_19369);
or UO_2284 (O_2284,N_19024,N_19649);
or UO_2285 (O_2285,N_19531,N_19323);
nand UO_2286 (O_2286,N_19074,N_19839);
nand UO_2287 (O_2287,N_19597,N_19096);
and UO_2288 (O_2288,N_19766,N_19819);
nand UO_2289 (O_2289,N_19169,N_19029);
or UO_2290 (O_2290,N_19131,N_19522);
and UO_2291 (O_2291,N_19602,N_19598);
xor UO_2292 (O_2292,N_19097,N_19523);
and UO_2293 (O_2293,N_19720,N_19408);
or UO_2294 (O_2294,N_19951,N_19964);
xnor UO_2295 (O_2295,N_19213,N_19183);
nand UO_2296 (O_2296,N_19609,N_19855);
or UO_2297 (O_2297,N_19600,N_19312);
nor UO_2298 (O_2298,N_19944,N_19738);
or UO_2299 (O_2299,N_19666,N_19388);
nand UO_2300 (O_2300,N_19074,N_19399);
and UO_2301 (O_2301,N_19440,N_19519);
nor UO_2302 (O_2302,N_19936,N_19612);
or UO_2303 (O_2303,N_19089,N_19769);
xnor UO_2304 (O_2304,N_19601,N_19205);
xnor UO_2305 (O_2305,N_19002,N_19859);
nand UO_2306 (O_2306,N_19315,N_19735);
xor UO_2307 (O_2307,N_19729,N_19591);
nor UO_2308 (O_2308,N_19295,N_19353);
and UO_2309 (O_2309,N_19989,N_19593);
and UO_2310 (O_2310,N_19932,N_19795);
nor UO_2311 (O_2311,N_19503,N_19034);
nor UO_2312 (O_2312,N_19876,N_19465);
or UO_2313 (O_2313,N_19175,N_19805);
nor UO_2314 (O_2314,N_19838,N_19700);
or UO_2315 (O_2315,N_19477,N_19667);
or UO_2316 (O_2316,N_19324,N_19235);
nor UO_2317 (O_2317,N_19882,N_19162);
nor UO_2318 (O_2318,N_19411,N_19465);
nand UO_2319 (O_2319,N_19852,N_19344);
xor UO_2320 (O_2320,N_19029,N_19445);
nor UO_2321 (O_2321,N_19349,N_19700);
or UO_2322 (O_2322,N_19543,N_19093);
and UO_2323 (O_2323,N_19205,N_19966);
and UO_2324 (O_2324,N_19117,N_19182);
nand UO_2325 (O_2325,N_19734,N_19827);
or UO_2326 (O_2326,N_19127,N_19145);
nor UO_2327 (O_2327,N_19029,N_19330);
xor UO_2328 (O_2328,N_19725,N_19034);
nand UO_2329 (O_2329,N_19033,N_19699);
nor UO_2330 (O_2330,N_19868,N_19916);
and UO_2331 (O_2331,N_19052,N_19458);
and UO_2332 (O_2332,N_19101,N_19725);
nand UO_2333 (O_2333,N_19126,N_19743);
nand UO_2334 (O_2334,N_19338,N_19558);
or UO_2335 (O_2335,N_19840,N_19459);
nand UO_2336 (O_2336,N_19151,N_19673);
nand UO_2337 (O_2337,N_19728,N_19492);
or UO_2338 (O_2338,N_19314,N_19202);
or UO_2339 (O_2339,N_19268,N_19085);
nor UO_2340 (O_2340,N_19378,N_19107);
nand UO_2341 (O_2341,N_19845,N_19292);
nand UO_2342 (O_2342,N_19837,N_19891);
and UO_2343 (O_2343,N_19449,N_19300);
or UO_2344 (O_2344,N_19136,N_19931);
nand UO_2345 (O_2345,N_19529,N_19379);
and UO_2346 (O_2346,N_19122,N_19177);
nor UO_2347 (O_2347,N_19439,N_19467);
or UO_2348 (O_2348,N_19591,N_19745);
nor UO_2349 (O_2349,N_19699,N_19382);
nor UO_2350 (O_2350,N_19933,N_19848);
nor UO_2351 (O_2351,N_19794,N_19524);
nor UO_2352 (O_2352,N_19109,N_19958);
xnor UO_2353 (O_2353,N_19214,N_19086);
or UO_2354 (O_2354,N_19970,N_19941);
nor UO_2355 (O_2355,N_19652,N_19085);
nor UO_2356 (O_2356,N_19107,N_19326);
or UO_2357 (O_2357,N_19856,N_19060);
nand UO_2358 (O_2358,N_19578,N_19196);
and UO_2359 (O_2359,N_19295,N_19236);
or UO_2360 (O_2360,N_19114,N_19380);
nand UO_2361 (O_2361,N_19257,N_19500);
and UO_2362 (O_2362,N_19815,N_19458);
and UO_2363 (O_2363,N_19621,N_19105);
nand UO_2364 (O_2364,N_19533,N_19663);
nand UO_2365 (O_2365,N_19928,N_19274);
or UO_2366 (O_2366,N_19241,N_19075);
nand UO_2367 (O_2367,N_19218,N_19672);
xor UO_2368 (O_2368,N_19214,N_19874);
and UO_2369 (O_2369,N_19759,N_19701);
nand UO_2370 (O_2370,N_19378,N_19898);
or UO_2371 (O_2371,N_19404,N_19925);
or UO_2372 (O_2372,N_19343,N_19818);
nand UO_2373 (O_2373,N_19743,N_19320);
nor UO_2374 (O_2374,N_19854,N_19500);
nand UO_2375 (O_2375,N_19467,N_19497);
or UO_2376 (O_2376,N_19345,N_19122);
nand UO_2377 (O_2377,N_19810,N_19682);
xnor UO_2378 (O_2378,N_19071,N_19327);
nand UO_2379 (O_2379,N_19184,N_19418);
and UO_2380 (O_2380,N_19133,N_19458);
xnor UO_2381 (O_2381,N_19137,N_19208);
xor UO_2382 (O_2382,N_19584,N_19789);
nand UO_2383 (O_2383,N_19276,N_19489);
or UO_2384 (O_2384,N_19321,N_19208);
nand UO_2385 (O_2385,N_19753,N_19336);
nand UO_2386 (O_2386,N_19878,N_19075);
nor UO_2387 (O_2387,N_19297,N_19593);
nor UO_2388 (O_2388,N_19840,N_19765);
nand UO_2389 (O_2389,N_19004,N_19003);
nor UO_2390 (O_2390,N_19556,N_19222);
and UO_2391 (O_2391,N_19637,N_19085);
nor UO_2392 (O_2392,N_19003,N_19263);
xor UO_2393 (O_2393,N_19353,N_19785);
nand UO_2394 (O_2394,N_19761,N_19986);
nor UO_2395 (O_2395,N_19013,N_19227);
nor UO_2396 (O_2396,N_19841,N_19908);
and UO_2397 (O_2397,N_19325,N_19562);
and UO_2398 (O_2398,N_19490,N_19635);
nand UO_2399 (O_2399,N_19680,N_19482);
nand UO_2400 (O_2400,N_19724,N_19106);
and UO_2401 (O_2401,N_19185,N_19552);
nand UO_2402 (O_2402,N_19383,N_19298);
nor UO_2403 (O_2403,N_19355,N_19667);
nand UO_2404 (O_2404,N_19803,N_19613);
nand UO_2405 (O_2405,N_19652,N_19324);
and UO_2406 (O_2406,N_19346,N_19572);
and UO_2407 (O_2407,N_19271,N_19047);
and UO_2408 (O_2408,N_19126,N_19074);
or UO_2409 (O_2409,N_19968,N_19534);
nand UO_2410 (O_2410,N_19403,N_19411);
nor UO_2411 (O_2411,N_19047,N_19941);
nor UO_2412 (O_2412,N_19484,N_19391);
or UO_2413 (O_2413,N_19751,N_19495);
and UO_2414 (O_2414,N_19969,N_19383);
nand UO_2415 (O_2415,N_19132,N_19771);
nor UO_2416 (O_2416,N_19567,N_19708);
nor UO_2417 (O_2417,N_19800,N_19286);
and UO_2418 (O_2418,N_19187,N_19180);
and UO_2419 (O_2419,N_19255,N_19872);
or UO_2420 (O_2420,N_19436,N_19169);
xor UO_2421 (O_2421,N_19411,N_19452);
or UO_2422 (O_2422,N_19275,N_19732);
or UO_2423 (O_2423,N_19559,N_19783);
nor UO_2424 (O_2424,N_19746,N_19970);
or UO_2425 (O_2425,N_19053,N_19746);
or UO_2426 (O_2426,N_19601,N_19537);
or UO_2427 (O_2427,N_19689,N_19193);
nor UO_2428 (O_2428,N_19704,N_19133);
and UO_2429 (O_2429,N_19628,N_19595);
xnor UO_2430 (O_2430,N_19113,N_19068);
and UO_2431 (O_2431,N_19374,N_19628);
and UO_2432 (O_2432,N_19290,N_19423);
or UO_2433 (O_2433,N_19562,N_19403);
xor UO_2434 (O_2434,N_19228,N_19726);
or UO_2435 (O_2435,N_19666,N_19746);
or UO_2436 (O_2436,N_19076,N_19345);
nand UO_2437 (O_2437,N_19046,N_19617);
nand UO_2438 (O_2438,N_19899,N_19615);
nor UO_2439 (O_2439,N_19279,N_19207);
nor UO_2440 (O_2440,N_19324,N_19374);
nor UO_2441 (O_2441,N_19383,N_19068);
nand UO_2442 (O_2442,N_19947,N_19430);
nand UO_2443 (O_2443,N_19103,N_19011);
nand UO_2444 (O_2444,N_19594,N_19206);
nand UO_2445 (O_2445,N_19395,N_19701);
and UO_2446 (O_2446,N_19521,N_19419);
nand UO_2447 (O_2447,N_19213,N_19643);
and UO_2448 (O_2448,N_19527,N_19236);
or UO_2449 (O_2449,N_19159,N_19576);
or UO_2450 (O_2450,N_19186,N_19807);
nand UO_2451 (O_2451,N_19324,N_19087);
and UO_2452 (O_2452,N_19099,N_19807);
and UO_2453 (O_2453,N_19484,N_19070);
or UO_2454 (O_2454,N_19181,N_19725);
nor UO_2455 (O_2455,N_19764,N_19020);
and UO_2456 (O_2456,N_19587,N_19525);
or UO_2457 (O_2457,N_19467,N_19683);
and UO_2458 (O_2458,N_19928,N_19356);
and UO_2459 (O_2459,N_19235,N_19461);
and UO_2460 (O_2460,N_19543,N_19903);
nand UO_2461 (O_2461,N_19392,N_19011);
or UO_2462 (O_2462,N_19902,N_19075);
nor UO_2463 (O_2463,N_19197,N_19036);
nor UO_2464 (O_2464,N_19622,N_19807);
nor UO_2465 (O_2465,N_19012,N_19397);
and UO_2466 (O_2466,N_19611,N_19546);
or UO_2467 (O_2467,N_19633,N_19245);
and UO_2468 (O_2468,N_19835,N_19675);
or UO_2469 (O_2469,N_19784,N_19786);
or UO_2470 (O_2470,N_19108,N_19885);
or UO_2471 (O_2471,N_19303,N_19888);
nand UO_2472 (O_2472,N_19191,N_19536);
nor UO_2473 (O_2473,N_19587,N_19518);
or UO_2474 (O_2474,N_19325,N_19388);
nand UO_2475 (O_2475,N_19349,N_19377);
and UO_2476 (O_2476,N_19511,N_19735);
and UO_2477 (O_2477,N_19329,N_19741);
or UO_2478 (O_2478,N_19643,N_19367);
xor UO_2479 (O_2479,N_19802,N_19207);
or UO_2480 (O_2480,N_19367,N_19990);
and UO_2481 (O_2481,N_19680,N_19266);
and UO_2482 (O_2482,N_19558,N_19967);
nor UO_2483 (O_2483,N_19308,N_19963);
xor UO_2484 (O_2484,N_19974,N_19395);
or UO_2485 (O_2485,N_19286,N_19300);
or UO_2486 (O_2486,N_19991,N_19836);
or UO_2487 (O_2487,N_19530,N_19220);
nor UO_2488 (O_2488,N_19647,N_19752);
and UO_2489 (O_2489,N_19955,N_19438);
nor UO_2490 (O_2490,N_19253,N_19250);
or UO_2491 (O_2491,N_19503,N_19105);
nor UO_2492 (O_2492,N_19484,N_19211);
or UO_2493 (O_2493,N_19430,N_19817);
and UO_2494 (O_2494,N_19215,N_19986);
and UO_2495 (O_2495,N_19550,N_19254);
or UO_2496 (O_2496,N_19192,N_19634);
nor UO_2497 (O_2497,N_19200,N_19629);
or UO_2498 (O_2498,N_19476,N_19850);
or UO_2499 (O_2499,N_19037,N_19749);
endmodule