module basic_3000_30000_3500_50_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
and U0 (N_0,In_2891,In_1987);
nand U1 (N_1,In_650,In_198);
or U2 (N_2,In_760,In_1335);
nand U3 (N_3,In_291,In_739);
nand U4 (N_4,In_507,In_848);
xor U5 (N_5,In_1149,In_1884);
xnor U6 (N_6,In_831,In_280);
or U7 (N_7,In_384,In_2397);
or U8 (N_8,In_56,In_2443);
or U9 (N_9,In_75,In_2263);
and U10 (N_10,In_1808,In_1915);
nor U11 (N_11,In_196,In_1762);
nand U12 (N_12,In_2220,In_844);
nor U13 (N_13,In_2919,In_407);
and U14 (N_14,In_1395,In_1879);
nand U15 (N_15,In_2608,In_2520);
nand U16 (N_16,In_2474,In_1301);
or U17 (N_17,In_2649,In_780);
or U18 (N_18,In_2136,In_1455);
or U19 (N_19,In_2002,In_911);
nor U20 (N_20,In_2395,In_921);
and U21 (N_21,In_1948,In_2344);
nand U22 (N_22,In_1347,In_1264);
nor U23 (N_23,In_2752,In_2498);
nand U24 (N_24,In_1393,In_615);
nor U25 (N_25,In_2989,In_2431);
or U26 (N_26,In_2529,In_2749);
xnor U27 (N_27,In_1878,In_1910);
xnor U28 (N_28,In_467,In_2177);
nor U29 (N_29,In_2051,In_1868);
xnor U30 (N_30,In_1578,In_1599);
nor U31 (N_31,In_547,In_1867);
or U32 (N_32,In_2437,In_2483);
nor U33 (N_33,In_40,In_614);
nand U34 (N_34,In_445,In_2281);
and U35 (N_35,In_2698,In_1709);
nand U36 (N_36,In_689,In_1000);
or U37 (N_37,In_1161,In_1354);
xnor U38 (N_38,In_1257,In_853);
nand U39 (N_39,In_569,In_664);
xor U40 (N_40,In_769,In_428);
xnor U41 (N_41,In_1827,In_954);
or U42 (N_42,In_2473,In_907);
nand U43 (N_43,In_157,In_341);
and U44 (N_44,In_1453,In_394);
or U45 (N_45,In_1986,In_457);
nand U46 (N_46,In_1289,In_2554);
and U47 (N_47,In_1816,In_2037);
and U48 (N_48,In_22,In_2417);
nand U49 (N_49,In_1267,In_1861);
nand U50 (N_50,In_402,In_826);
or U51 (N_51,In_2134,In_78);
and U52 (N_52,In_540,In_1359);
xnor U53 (N_53,In_1083,In_2075);
xor U54 (N_54,In_275,In_434);
and U55 (N_55,In_2700,In_1026);
xnor U56 (N_56,In_2476,In_1725);
and U57 (N_57,In_2238,In_2560);
xnor U58 (N_58,In_1413,In_1869);
or U59 (N_59,In_2696,In_1263);
nand U60 (N_60,In_2944,In_970);
nand U61 (N_61,In_711,In_2192);
nor U62 (N_62,In_1760,In_509);
or U63 (N_63,In_890,In_1014);
nor U64 (N_64,In_82,In_2772);
xor U65 (N_65,In_2092,In_68);
xnor U66 (N_66,In_1520,In_997);
nand U67 (N_67,In_251,In_2224);
and U68 (N_68,In_1602,In_1936);
and U69 (N_69,In_1387,In_583);
or U70 (N_70,In_2769,In_2506);
and U71 (N_71,In_2874,In_2949);
or U72 (N_72,In_1082,In_316);
and U73 (N_73,In_1767,In_795);
or U74 (N_74,In_1744,In_2633);
nor U75 (N_75,In_2499,In_260);
nor U76 (N_76,In_107,In_436);
or U77 (N_77,In_2124,In_70);
nand U78 (N_78,In_1484,In_2314);
xor U79 (N_79,In_192,In_2083);
nor U80 (N_80,In_1142,In_723);
nand U81 (N_81,In_2973,In_2068);
and U82 (N_82,In_466,In_863);
and U83 (N_83,In_370,In_726);
nor U84 (N_84,In_50,In_2343);
xor U85 (N_85,In_1045,In_1848);
nor U86 (N_86,In_2105,In_2807);
and U87 (N_87,In_1600,In_1670);
or U88 (N_88,In_1231,In_2577);
xnor U89 (N_89,In_1636,In_142);
and U90 (N_90,In_1841,In_2928);
nand U91 (N_91,In_2298,In_354);
xnor U92 (N_92,In_2315,In_824);
nand U93 (N_93,In_2370,In_715);
nand U94 (N_94,In_918,In_2492);
nand U95 (N_95,In_496,In_1889);
nor U96 (N_96,In_745,In_506);
xor U97 (N_97,In_2864,In_1182);
or U98 (N_98,In_1888,In_1729);
or U99 (N_99,In_1732,In_1351);
nor U100 (N_100,In_2182,In_1047);
and U101 (N_101,In_654,In_2272);
nor U102 (N_102,In_986,In_1819);
nand U103 (N_103,In_1156,In_95);
nand U104 (N_104,In_2023,In_1079);
nand U105 (N_105,In_253,In_2440);
nand U106 (N_106,In_1394,In_2328);
xor U107 (N_107,In_2941,In_1807);
nor U108 (N_108,In_1803,In_1653);
nand U109 (N_109,In_164,In_2494);
nand U110 (N_110,In_2674,In_1200);
nor U111 (N_111,In_543,In_1739);
and U112 (N_112,In_2463,In_173);
or U113 (N_113,In_9,In_1718);
and U114 (N_114,In_38,In_893);
xor U115 (N_115,In_1569,In_1356);
or U116 (N_116,In_1136,In_1642);
nand U117 (N_117,In_630,In_1877);
xor U118 (N_118,In_1315,In_2384);
xor U119 (N_119,In_2525,In_221);
xor U120 (N_120,In_1728,In_313);
nand U121 (N_121,In_1557,In_659);
nand U122 (N_122,In_1857,In_597);
nand U123 (N_123,In_1780,In_2717);
or U124 (N_124,In_1781,In_936);
nor U125 (N_125,In_2726,In_1518);
xor U126 (N_126,In_2273,In_1839);
and U127 (N_127,In_1917,In_1032);
nand U128 (N_128,In_287,In_2042);
and U129 (N_129,In_2122,In_2974);
and U130 (N_130,In_380,In_2838);
nor U131 (N_131,In_2318,In_2833);
nor U132 (N_132,In_411,In_812);
and U133 (N_133,In_660,In_2945);
and U134 (N_134,In_1421,In_2996);
xnor U135 (N_135,In_1914,In_111);
nor U136 (N_136,In_976,In_1285);
nand U137 (N_137,In_2363,In_533);
xor U138 (N_138,In_2196,In_2537);
xor U139 (N_139,In_1514,In_1988);
or U140 (N_140,In_2713,In_299);
nand U141 (N_141,In_560,In_1522);
and U142 (N_142,In_2208,In_1939);
nor U143 (N_143,In_63,In_74);
xor U144 (N_144,In_1517,In_1903);
xor U145 (N_145,In_869,In_1958);
and U146 (N_146,In_1445,In_2541);
nor U147 (N_147,In_2994,In_351);
xor U148 (N_148,In_1234,In_2894);
xnor U149 (N_149,In_2046,In_237);
and U150 (N_150,In_1570,In_2360);
and U151 (N_151,In_105,In_1225);
or U152 (N_152,In_1253,In_602);
xor U153 (N_153,In_2236,In_1761);
xor U154 (N_154,In_2140,In_2151);
nand U155 (N_155,In_1168,In_1710);
or U156 (N_156,In_725,In_2362);
and U157 (N_157,In_2732,In_2968);
nor U158 (N_158,In_1496,In_594);
xor U159 (N_159,In_216,In_2148);
and U160 (N_160,In_2561,In_1194);
xnor U161 (N_161,In_1740,In_2670);
or U162 (N_162,In_1478,In_931);
and U163 (N_163,In_1148,In_1959);
or U164 (N_164,In_668,In_2606);
and U165 (N_165,In_989,In_152);
nand U166 (N_166,In_185,In_1124);
nand U167 (N_167,In_2706,In_2993);
nor U168 (N_168,In_2867,In_666);
nor U169 (N_169,In_2321,In_209);
nor U170 (N_170,In_2286,In_749);
nand U171 (N_171,In_2767,In_1992);
and U172 (N_172,In_2840,In_218);
or U173 (N_173,In_952,In_545);
or U174 (N_174,In_1108,In_2985);
nor U175 (N_175,In_1126,In_383);
or U176 (N_176,In_2578,In_1458);
nor U177 (N_177,In_1985,In_203);
nand U178 (N_178,In_461,In_1070);
xor U179 (N_179,In_1392,In_2672);
nor U180 (N_180,In_127,In_317);
nor U181 (N_181,In_2695,In_1817);
nor U182 (N_182,In_1037,In_2789);
xnor U183 (N_183,In_1115,In_1409);
or U184 (N_184,In_2609,In_1286);
nor U185 (N_185,In_870,In_493);
and U186 (N_186,In_1707,In_2442);
nand U187 (N_187,In_2623,In_2511);
nand U188 (N_188,In_2091,In_2123);
or U189 (N_189,In_1691,In_1436);
and U190 (N_190,In_2802,In_1620);
or U191 (N_191,In_1287,In_2354);
xor U192 (N_192,In_191,In_2803);
or U193 (N_193,In_153,In_514);
nor U194 (N_194,In_2116,In_1947);
nand U195 (N_195,In_2175,In_2256);
or U196 (N_196,In_2358,In_2830);
and U197 (N_197,In_1030,In_2636);
nor U198 (N_198,In_1088,In_311);
nor U199 (N_199,In_2518,In_499);
and U200 (N_200,In_994,In_42);
nor U201 (N_201,In_1127,In_1308);
nor U202 (N_202,In_410,In_1317);
xnor U203 (N_203,In_2795,In_1934);
and U204 (N_204,In_2898,In_2304);
and U205 (N_205,In_12,In_1318);
or U206 (N_206,In_43,In_71);
and U207 (N_207,In_2504,In_1971);
nor U208 (N_208,In_451,In_2992);
nor U209 (N_209,In_1454,In_632);
nand U210 (N_210,In_913,In_2762);
nand U211 (N_211,In_558,In_1306);
xnor U212 (N_212,In_1275,In_991);
xor U213 (N_213,In_643,In_2013);
and U214 (N_214,In_678,In_2591);
and U215 (N_215,In_995,In_638);
xor U216 (N_216,In_2248,In_2163);
nand U217 (N_217,In_2459,In_2820);
xor U218 (N_218,In_1577,In_782);
xor U219 (N_219,In_2173,In_1391);
xor U220 (N_220,In_945,In_549);
xnor U221 (N_221,In_1104,In_141);
and U222 (N_222,In_2188,In_690);
and U223 (N_223,In_2157,In_752);
nand U224 (N_224,In_2438,In_1622);
and U225 (N_225,In_683,In_2559);
and U226 (N_226,In_1506,In_160);
nand U227 (N_227,In_2382,In_339);
nor U228 (N_228,In_1831,In_2794);
nor U229 (N_229,In_2491,In_1349);
nand U230 (N_230,In_940,In_372);
and U231 (N_231,In_1751,In_1292);
or U232 (N_232,In_548,In_2667);
nand U233 (N_233,In_817,In_733);
nor U234 (N_234,In_695,In_1820);
and U235 (N_235,In_1724,In_629);
xnor U236 (N_236,In_842,In_1470);
or U237 (N_237,In_401,In_770);
nor U238 (N_238,In_2813,In_1446);
or U239 (N_239,In_2966,In_2290);
nor U240 (N_240,In_2793,In_590);
xnor U241 (N_241,In_2643,In_1702);
nand U242 (N_242,In_892,In_2509);
xnor U243 (N_243,In_2065,In_2688);
nand U244 (N_244,In_1012,In_1175);
xnor U245 (N_245,In_1615,In_1103);
and U246 (N_246,In_1313,In_967);
xor U247 (N_247,In_2579,In_132);
xnor U248 (N_248,In_101,In_778);
and U249 (N_249,In_1573,In_1399);
nor U250 (N_250,In_292,In_811);
and U251 (N_251,In_958,In_2255);
nand U252 (N_252,In_279,In_2927);
and U253 (N_253,In_2675,In_1850);
nand U254 (N_254,In_1278,In_2661);
nand U255 (N_255,In_357,In_308);
and U256 (N_256,In_1303,In_1906);
xor U257 (N_257,In_462,In_577);
nor U258 (N_258,In_1009,In_2405);
nand U259 (N_259,In_828,In_2741);
and U260 (N_260,In_1525,In_228);
and U261 (N_261,In_1945,In_150);
and U262 (N_262,In_2436,In_1558);
nand U263 (N_263,In_2102,In_163);
nand U264 (N_264,In_1534,In_2333);
and U265 (N_265,In_347,In_2621);
nand U266 (N_266,In_2630,In_1466);
and U267 (N_267,In_737,In_2656);
nand U268 (N_268,In_667,In_2378);
or U269 (N_269,In_2441,In_2233);
nor U270 (N_270,In_523,In_821);
and U271 (N_271,In_102,In_786);
nand U272 (N_272,In_2082,In_1552);
xor U273 (N_273,In_2217,In_1430);
or U274 (N_274,In_2510,In_1960);
xnor U275 (N_275,In_2508,In_246);
xnor U276 (N_276,In_2612,In_1941);
or U277 (N_277,In_367,In_2266);
xnor U278 (N_278,In_2486,In_1684);
xnor U279 (N_279,In_2189,In_2409);
nor U280 (N_280,In_2193,In_1655);
xnor U281 (N_281,In_147,In_2393);
xor U282 (N_282,In_1633,In_727);
and U283 (N_283,In_2635,In_2740);
xor U284 (N_284,In_2539,In_2770);
or U285 (N_285,In_1475,In_106);
or U286 (N_286,In_485,In_2357);
or U287 (N_287,In_1482,In_2756);
nand U288 (N_288,In_882,In_2368);
nor U289 (N_289,In_1976,In_1288);
nor U290 (N_290,In_1645,In_1626);
and U291 (N_291,In_712,In_2070);
nor U292 (N_292,In_2212,In_60);
or U293 (N_293,In_2811,In_2753);
xnor U294 (N_294,In_1016,In_646);
nor U295 (N_295,In_1251,In_1450);
nand U296 (N_296,In_242,In_883);
xor U297 (N_297,In_1711,In_1488);
nor U298 (N_298,In_2061,In_529);
or U299 (N_299,In_333,In_110);
and U300 (N_300,In_1297,In_1134);
xor U301 (N_301,In_1102,In_943);
or U302 (N_302,In_2089,In_1172);
nor U303 (N_303,In_2191,In_765);
nand U304 (N_304,In_1069,In_2285);
nor U305 (N_305,In_399,In_5);
or U306 (N_306,In_2638,In_2462);
nand U307 (N_307,In_1266,In_1374);
or U308 (N_308,In_2352,In_28);
or U309 (N_309,In_1597,In_187);
nor U310 (N_310,In_184,In_2844);
nor U311 (N_311,In_2214,In_1058);
or U312 (N_312,In_416,In_2341);
nand U313 (N_313,In_2758,In_2129);
or U314 (N_314,In_413,In_645);
xor U315 (N_315,In_1311,In_793);
nand U316 (N_316,In_2654,In_1050);
nor U317 (N_317,In_2781,In_2015);
nand U318 (N_318,In_1205,In_2871);
and U319 (N_319,In_1222,In_790);
or U320 (N_320,In_1511,In_1426);
xnor U321 (N_321,In_2748,In_677);
nand U322 (N_322,In_956,In_2745);
nand U323 (N_323,In_2077,In_2955);
nor U324 (N_324,In_1899,In_79);
nand U325 (N_325,In_31,In_2587);
xnor U326 (N_326,In_2154,In_584);
xnor U327 (N_327,In_2307,In_125);
nand U328 (N_328,In_942,In_2109);
and U329 (N_329,In_1706,In_2785);
nor U330 (N_330,In_591,In_1801);
xnor U331 (N_331,In_1591,In_2495);
and U332 (N_332,In_709,In_2020);
nand U333 (N_333,In_1556,In_1893);
or U334 (N_334,In_2467,In_2144);
nor U335 (N_335,In_2975,In_2637);
nor U336 (N_336,In_2917,In_2104);
and U337 (N_337,In_1408,In_1838);
or U338 (N_338,In_774,In_2359);
nand U339 (N_339,In_1386,In_1494);
xnor U340 (N_340,In_1840,In_131);
xor U341 (N_341,In_1646,In_1679);
or U342 (N_342,In_2006,In_290);
and U343 (N_343,In_532,In_2569);
xor U344 (N_344,In_2062,In_1871);
nand U345 (N_345,In_2736,In_2260);
and U346 (N_346,In_338,In_877);
and U347 (N_347,In_2800,In_24);
xnor U348 (N_348,In_2774,In_2283);
nor U349 (N_349,In_644,In_2589);
xor U350 (N_350,In_2567,In_2270);
nor U351 (N_351,In_949,In_694);
nand U352 (N_352,In_801,In_1923);
or U353 (N_353,In_2149,In_620);
or U354 (N_354,In_562,In_2950);
nand U355 (N_355,In_1117,In_2646);
and U356 (N_356,In_2161,In_1330);
nand U357 (N_357,In_2117,In_1063);
nand U358 (N_358,In_623,In_1953);
or U359 (N_359,In_775,In_621);
nand U360 (N_360,In_2399,In_957);
or U361 (N_361,In_1262,In_2484);
nand U362 (N_362,In_1485,In_1084);
or U363 (N_363,In_2538,In_139);
nor U364 (N_364,In_2288,In_1737);
and U365 (N_365,In_318,In_2414);
nand U366 (N_366,In_2863,In_1324);
nand U367 (N_367,In_252,In_787);
and U368 (N_368,In_208,In_463);
or U369 (N_369,In_1252,In_1398);
nor U370 (N_370,In_2592,In_406);
xnor U371 (N_371,In_2766,In_996);
nor U372 (N_372,In_705,In_2961);
nor U373 (N_373,In_753,In_1554);
nor U374 (N_374,In_839,In_1087);
nand U375 (N_375,In_47,In_1510);
nand U376 (N_376,In_2948,In_2045);
xor U377 (N_377,In_61,In_2296);
or U378 (N_378,In_1241,In_1774);
or U379 (N_379,In_1362,In_1943);
xnor U380 (N_380,In_323,In_433);
nor U381 (N_381,In_1894,In_206);
nand U382 (N_382,In_1814,In_1442);
and U383 (N_383,In_360,In_2223);
xnor U384 (N_384,In_567,In_264);
nor U385 (N_385,In_2058,In_914);
and U386 (N_386,In_137,In_2433);
and U387 (N_387,In_1457,In_2870);
and U388 (N_388,In_980,In_321);
and U389 (N_389,In_2522,In_2166);
xnor U390 (N_390,In_2365,In_1590);
xor U391 (N_391,In_1340,In_2531);
nor U392 (N_392,In_220,In_2097);
or U393 (N_393,In_1926,In_2044);
and U394 (N_394,In_1750,In_2216);
and U395 (N_395,In_1049,In_767);
and U396 (N_396,In_2682,In_306);
nor U397 (N_397,In_2297,In_2241);
xnor U398 (N_398,In_2012,In_1130);
nor U399 (N_399,In_2095,In_55);
nor U400 (N_400,In_1388,In_754);
nand U401 (N_401,In_1833,In_2711);
nand U402 (N_402,In_2849,In_856);
xor U403 (N_403,In_2703,In_186);
and U404 (N_404,In_438,In_2856);
nand U405 (N_405,In_570,In_2435);
and U406 (N_406,In_1428,In_1298);
nand U407 (N_407,In_1585,In_2502);
or U408 (N_408,In_2905,In_478);
nand U409 (N_409,In_1563,In_86);
or U410 (N_410,In_2664,In_2827);
nor U411 (N_411,In_1162,In_2596);
nor U412 (N_412,In_2648,In_1304);
and U413 (N_413,In_681,In_1190);
xor U414 (N_414,In_2930,In_2824);
nand U415 (N_415,In_315,In_2316);
nand U416 (N_416,In_682,In_2049);
xor U417 (N_417,In_2516,In_494);
xor U418 (N_418,In_2171,In_80);
nand U419 (N_419,In_271,In_1497);
nand U420 (N_420,In_447,In_2330);
nor U421 (N_421,In_30,In_335);
nand U422 (N_422,In_1197,In_1280);
or U423 (N_423,In_1619,In_1248);
xor U424 (N_424,In_2876,In_302);
or U425 (N_425,In_205,In_508);
or U426 (N_426,In_922,In_2660);
and U427 (N_427,In_219,In_2055);
nand U428 (N_428,In_1876,In_103);
xnor U429 (N_429,In_707,In_2331);
or U430 (N_430,In_1477,In_2059);
nor U431 (N_431,In_674,In_272);
nor U432 (N_432,In_895,In_2852);
or U433 (N_433,In_2195,In_1361);
nand U434 (N_434,In_87,In_1595);
nand U435 (N_435,In_2025,In_751);
xor U436 (N_436,In_649,In_2555);
or U437 (N_437,In_2977,In_2501);
nor U438 (N_438,In_1238,In_959);
and U439 (N_439,In_868,In_199);
xnor U440 (N_440,In_21,In_1532);
xnor U441 (N_441,In_1765,In_2323);
and U442 (N_442,In_1696,In_1309);
xnor U443 (N_443,In_982,In_721);
nand U444 (N_444,In_200,In_1464);
or U445 (N_445,In_1571,In_1424);
nand U446 (N_446,In_2746,In_2910);
or U447 (N_447,In_1255,In_766);
nand U448 (N_448,In_917,In_1748);
or U449 (N_449,In_229,In_444);
nand U450 (N_450,In_983,In_885);
nor U451 (N_451,In_901,In_1203);
or U452 (N_452,In_2477,In_2470);
nand U453 (N_453,In_1813,In_1325);
or U454 (N_454,In_2312,In_1284);
and U455 (N_455,In_2086,In_2207);
and U456 (N_456,In_100,In_2375);
xor U457 (N_457,In_1053,In_953);
nand U458 (N_458,In_303,In_2201);
nand U459 (N_459,In_1766,In_2907);
xor U460 (N_460,In_2835,In_288);
nor U461 (N_461,In_2653,In_939);
nand U462 (N_462,In_1783,In_1400);
nor U463 (N_463,In_2535,In_1671);
and U464 (N_464,In_500,In_1528);
xor U465 (N_465,In_553,In_1666);
or U466 (N_466,In_2797,In_802);
nor U467 (N_467,In_1358,In_119);
nor U468 (N_468,In_617,In_641);
or U469 (N_469,In_1931,In_1060);
nor U470 (N_470,In_231,In_2112);
or U471 (N_471,In_85,In_679);
and U472 (N_472,In_431,In_1860);
nor U473 (N_473,In_898,In_2167);
or U474 (N_474,In_430,In_1245);
xor U475 (N_475,In_1397,In_1193);
nand U476 (N_476,In_52,In_2458);
nor U477 (N_477,In_2530,In_194);
nand U478 (N_478,In_1199,In_1333);
xor U479 (N_479,In_656,In_2937);
xnor U480 (N_480,In_2760,In_2096);
nor U481 (N_481,In_415,In_1006);
xnor U482 (N_482,In_987,In_1777);
xor U483 (N_483,In_599,In_2213);
and U484 (N_484,In_1944,In_1900);
nor U485 (N_485,In_2553,In_806);
and U486 (N_486,In_2737,In_1523);
or U487 (N_487,In_2017,In_16);
xnor U488 (N_488,In_552,In_1021);
nor U489 (N_489,In_1085,In_435);
nor U490 (N_490,In_2187,In_1290);
and U491 (N_491,In_2651,In_2465);
nand U492 (N_492,In_2100,In_1961);
nand U493 (N_493,In_1598,In_376);
nand U494 (N_494,In_1742,In_2622);
xnor U495 (N_495,In_2957,In_2231);
and U496 (N_496,In_2366,In_1687);
nand U497 (N_497,In_1946,In_167);
and U498 (N_498,In_1295,In_2814);
xor U499 (N_499,In_175,In_2895);
and U500 (N_500,In_2963,In_93);
or U501 (N_501,In_489,In_2822);
xor U502 (N_502,In_2744,In_1091);
nor U503 (N_503,In_2593,In_155);
nand U504 (N_504,In_1970,In_366);
and U505 (N_505,In_2990,In_2731);
or U506 (N_506,In_248,In_1447);
nand U507 (N_507,In_2988,In_2407);
or U508 (N_508,In_2926,In_849);
and U509 (N_509,In_546,In_73);
nor U510 (N_510,In_1885,In_517);
or U511 (N_511,In_1845,In_2657);
nor U512 (N_512,In_25,In_193);
xor U513 (N_513,In_2598,In_796);
or U514 (N_514,In_1796,In_1089);
nor U515 (N_515,In_1828,In_2965);
nor U516 (N_516,In_2278,In_2727);
xnor U517 (N_517,In_2962,In_1073);
or U518 (N_518,In_14,In_2069);
and U519 (N_519,In_2970,In_2862);
or U520 (N_520,In_1972,In_420);
nor U521 (N_521,In_1112,In_2179);
xnor U522 (N_522,In_1339,In_2348);
nand U523 (N_523,In_244,In_2210);
and U524 (N_524,In_1076,In_2115);
xor U525 (N_525,In_2039,In_1180);
xor U526 (N_526,In_919,In_2480);
xor U527 (N_527,In_2707,In_655);
xor U528 (N_528,In_97,In_1133);
nand U529 (N_529,In_1404,In_822);
nor U530 (N_530,In_2558,In_2139);
and U531 (N_531,In_568,In_1240);
or U532 (N_532,In_1823,In_1165);
nor U533 (N_533,In_2235,In_932);
nand U534 (N_534,In_671,In_700);
nor U535 (N_535,In_1733,In_1071);
nand U536 (N_536,In_2935,In_1260);
nor U537 (N_537,In_563,In_2710);
xnor U538 (N_538,In_2137,In_2914);
nor U539 (N_539,In_1144,In_1995);
or U540 (N_540,In_44,In_1141);
or U541 (N_541,In_2739,In_2999);
or U542 (N_542,In_385,In_162);
or U543 (N_543,In_2971,In_2253);
xnor U544 (N_544,In_820,In_48);
or U545 (N_545,In_1650,In_1095);
or U546 (N_546,In_2728,In_1415);
or U547 (N_547,In_2088,In_72);
xor U548 (N_548,In_2572,In_295);
xnor U549 (N_549,In_2604,In_521);
xor U550 (N_550,In_736,In_1465);
xor U551 (N_551,In_1272,In_1815);
or U552 (N_552,In_665,In_1204);
or U553 (N_553,In_2426,In_748);
xnor U554 (N_554,In_889,In_1365);
xor U555 (N_555,In_1249,In_2056);
or U556 (N_556,In_146,In_116);
and U557 (N_557,In_1011,In_1625);
or U558 (N_558,In_2655,In_2460);
or U559 (N_559,In_2846,In_1100);
or U560 (N_560,In_884,In_1727);
nor U561 (N_561,In_1693,In_136);
nand U562 (N_562,In_2678,In_800);
or U563 (N_563,In_2447,In_1437);
xnor U564 (N_564,In_2563,In_1401);
and U565 (N_565,In_278,In_843);
and U566 (N_566,In_2311,In_326);
nor U567 (N_567,In_1772,In_993);
xor U568 (N_568,In_1639,In_329);
or U569 (N_569,In_2127,In_1773);
xor U570 (N_570,In_717,In_1847);
nand U571 (N_571,In_2743,In_1486);
nand U572 (N_572,In_2887,In_1492);
and U573 (N_573,In_2222,In_1033);
or U574 (N_574,In_2428,In_1039);
nor U575 (N_575,In_1348,In_2747);
nor U576 (N_576,In_1980,In_247);
and U577 (N_577,In_2582,In_1922);
and U578 (N_578,In_469,In_734);
xnor U579 (N_579,In_1508,In_1504);
nor U580 (N_580,In_1730,In_1575);
or U581 (N_581,In_2138,In_960);
and U582 (N_582,In_495,In_345);
or U583 (N_583,In_2503,In_2411);
nor U584 (N_584,In_1562,In_312);
xor U585 (N_585,In_2387,In_334);
or U586 (N_586,In_369,In_815);
or U587 (N_587,In_1364,In_239);
and U588 (N_588,In_910,In_352);
xor U589 (N_589,In_2228,In_1094);
and U590 (N_590,In_589,In_1024);
or U591 (N_591,In_809,In_2825);
and U592 (N_592,In_2854,In_2030);
nand U593 (N_593,In_1965,In_1254);
or U594 (N_594,In_1034,In_544);
xor U595 (N_595,In_1206,In_1270);
nor U596 (N_596,In_859,In_2274);
nor U597 (N_597,In_2584,In_2763);
xor U598 (N_598,In_2995,In_2714);
xnor U599 (N_599,In_2594,In_1256);
and U600 (N_600,In_2642,N_94);
and U601 (N_601,In_1319,In_2036);
or U602 (N_602,In_1700,In_1242);
and U603 (N_603,In_819,In_2346);
or U604 (N_604,In_1699,In_1469);
nor U605 (N_605,In_2615,N_234);
nand U606 (N_606,N_122,In_364);
nand U607 (N_607,N_335,In_2410);
xnor U608 (N_608,In_2374,In_1886);
or U609 (N_609,In_1822,In_1863);
and U610 (N_610,In_1681,In_933);
xnor U611 (N_611,N_434,N_106);
and U612 (N_612,In_524,N_119);
and U613 (N_613,In_1769,In_1676);
xnor U614 (N_614,N_392,In_2765);
xor U615 (N_615,In_580,N_99);
xnor U616 (N_616,In_2725,In_1129);
nor U617 (N_617,In_1826,N_214);
nor U618 (N_618,In_611,N_125);
or U619 (N_619,In_1326,In_1167);
and U620 (N_620,In_1657,N_213);
xnor U621 (N_621,In_2631,N_110);
nor U622 (N_622,In_2308,In_676);
nand U623 (N_623,N_535,In_551);
xnor U624 (N_624,N_302,In_1277);
nor U625 (N_625,In_2242,In_2673);
nor U626 (N_626,In_459,In_818);
and U627 (N_627,N_473,In_1367);
nand U628 (N_628,In_2881,In_286);
nor U629 (N_629,N_259,In_747);
nand U630 (N_630,In_1535,In_756);
or U631 (N_631,N_195,N_19);
and U632 (N_632,In_2901,In_1444);
xor U633 (N_633,In_1594,In_1935);
nand U634 (N_634,N_380,In_426);
xor U635 (N_635,In_988,N_478);
or U636 (N_636,In_1618,In_1081);
and U637 (N_637,N_591,In_832);
xor U638 (N_638,In_270,In_1451);
nor U639 (N_639,In_1539,N_536);
or U640 (N_640,In_525,In_3);
nor U641 (N_641,In_8,In_881);
and U642 (N_642,In_722,In_1540);
nor U643 (N_643,In_2276,In_1460);
nand U644 (N_644,In_1770,In_698);
nor U645 (N_645,In_2108,In_1064);
nand U646 (N_646,N_247,In_222);
xnor U647 (N_647,In_1758,In_935);
nor U648 (N_648,In_1332,N_484);
xor U649 (N_649,In_2369,In_2626);
xnor U650 (N_650,N_53,In_2540);
nor U651 (N_651,N_469,In_586);
or U652 (N_652,In_2932,N_486);
nand U653 (N_653,In_2066,In_1660);
nor U654 (N_654,In_2568,In_293);
nand U655 (N_655,In_2300,In_1481);
and U656 (N_656,In_1853,In_973);
nor U657 (N_657,In_2090,N_320);
or U658 (N_658,In_149,N_272);
nand U659 (N_659,In_210,In_2418);
nor U660 (N_660,In_224,In_808);
nand U661 (N_661,In_2427,In_1145);
nor U662 (N_662,In_1061,N_520);
nand U663 (N_663,N_246,In_2356);
or U664 (N_664,In_2913,In_177);
nor U665 (N_665,In_512,In_1726);
nand U666 (N_666,In_858,In_1370);
xnor U667 (N_667,N_578,In_300);
nand U668 (N_668,N_537,In_2512);
or U669 (N_669,N_428,In_1043);
and U670 (N_670,In_1782,In_374);
nor U671 (N_671,N_61,N_269);
or U672 (N_672,In_1157,In_1291);
or U673 (N_673,In_845,In_2237);
and U674 (N_674,N_14,In_2424);
xnor U675 (N_675,In_814,N_396);
and U676 (N_676,In_148,In_571);
xor U677 (N_677,In_2546,In_2419);
xnor U678 (N_678,N_514,In_1652);
xor U679 (N_679,In_2557,In_2034);
nor U680 (N_680,In_977,In_1759);
nand U681 (N_681,N_526,In_2351);
or U682 (N_682,In_2472,In_503);
nor U683 (N_683,In_699,In_750);
nor U684 (N_684,In_2038,N_471);
xor U685 (N_685,In_215,In_77);
nor U686 (N_686,N_80,N_204);
nand U687 (N_687,In_2203,N_144);
or U688 (N_688,N_345,In_2861);
nand U689 (N_689,N_185,In_365);
nor U690 (N_690,N_546,In_2218);
or U691 (N_691,In_607,In_1322);
and U692 (N_692,In_1346,In_841);
nand U693 (N_693,In_2668,N_583);
xnor U694 (N_694,In_2923,N_224);
nor U695 (N_695,In_759,N_340);
and U696 (N_696,In_691,In_1452);
or U697 (N_697,N_179,N_162);
xnor U698 (N_698,In_2094,In_2338);
xor U699 (N_699,In_233,In_1797);
xnor U700 (N_700,In_449,N_198);
and U701 (N_701,In_1989,In_2209);
xor U702 (N_702,In_1789,In_1459);
or U703 (N_703,In_207,In_2597);
and U704 (N_704,N_303,N_8);
xnor U705 (N_705,In_484,In_343);
or U706 (N_706,N_548,N_565);
and U707 (N_707,In_2939,In_2869);
nor U708 (N_708,In_2507,In_1090);
or U709 (N_709,In_1991,In_283);
nor U710 (N_710,In_2823,In_121);
nor U711 (N_711,In_1704,In_1183);
or U712 (N_712,In_62,In_658);
or U713 (N_713,In_2174,In_502);
nand U714 (N_714,N_132,In_1870);
nor U715 (N_715,In_2379,In_262);
nor U716 (N_716,In_835,In_2704);
nor U717 (N_717,In_1561,In_1235);
nor U718 (N_718,In_2946,In_140);
xor U719 (N_719,In_1153,In_1123);
or U720 (N_720,In_2377,In_1065);
or U721 (N_721,In_731,In_282);
xor U722 (N_722,N_333,N_491);
nor U723 (N_723,N_366,In_1835);
and U724 (N_724,In_2386,In_11);
xnor U725 (N_725,In_672,In_1406);
nor U726 (N_726,In_1927,In_6);
or U727 (N_727,In_720,In_2389);
and U728 (N_728,In_1631,In_1323);
xor U729 (N_729,In_1411,In_526);
or U730 (N_730,In_124,N_284);
xor U731 (N_731,In_1341,In_684);
and U732 (N_732,In_2843,N_124);
nor U733 (N_733,In_1334,In_1975);
nand U734 (N_734,In_1471,In_1668);
xor U735 (N_735,In_1589,In_473);
xor U736 (N_736,In_799,N_257);
nand U737 (N_737,In_1170,In_1320);
or U738 (N_738,In_1849,In_2074);
xnor U739 (N_739,In_762,N_190);
nand U740 (N_740,N_82,In_1821);
nand U741 (N_741,In_2873,In_1908);
xnor U742 (N_742,In_1842,In_109);
and U743 (N_743,N_300,N_101);
or U744 (N_744,In_2110,N_276);
or U745 (N_745,In_518,N_375);
xor U746 (N_746,In_862,In_2128);
nor U747 (N_747,In_636,N_193);
nor U748 (N_748,N_517,In_268);
xor U749 (N_749,N_560,N_38);
nor U750 (N_750,N_238,N_45);
nand U751 (N_751,N_358,In_1938);
nor U752 (N_752,N_438,In_1345);
nand U753 (N_753,In_1111,In_628);
and U754 (N_754,In_1271,N_441);
xnor U755 (N_755,In_2780,In_2326);
xnor U756 (N_756,In_1307,In_1013);
xnor U757 (N_757,N_160,In_66);
or U758 (N_758,In_2057,In_2644);
nand U759 (N_759,N_593,N_482);
and U760 (N_760,In_557,In_1434);
and U761 (N_761,In_2032,In_2875);
or U762 (N_762,N_63,In_114);
xor U763 (N_763,In_2866,In_1321);
and U764 (N_764,In_1512,In_1735);
and U765 (N_765,In_1360,In_15);
nor U766 (N_766,In_2295,N_381);
or U767 (N_767,In_609,In_961);
or U768 (N_768,N_25,In_2773);
or U769 (N_769,In_1865,In_742);
xor U770 (N_770,N_400,N_218);
nor U771 (N_771,In_2865,N_50);
xnor U772 (N_772,In_225,N_296);
and U773 (N_773,In_307,In_639);
nand U774 (N_774,N_468,In_2339);
nor U775 (N_775,In_1664,In_1213);
nand U776 (N_776,In_823,N_96);
nor U777 (N_777,In_2886,In_2860);
xnor U778 (N_778,In_1747,In_1674);
or U779 (N_779,In_771,N_498);
and U780 (N_780,In_1483,N_487);
and U781 (N_781,In_1612,In_400);
xnor U782 (N_782,In_2317,In_1553);
nor U783 (N_783,In_916,N_184);
nand U784 (N_784,In_601,N_343);
and U785 (N_785,In_608,N_362);
nand U786 (N_786,N_415,In_487);
nand U787 (N_787,In_1537,In_2444);
or U788 (N_788,In_2131,In_2831);
or U789 (N_789,N_389,In_274);
or U790 (N_790,In_470,In_1383);
or U791 (N_791,In_581,In_2259);
nor U792 (N_792,In_2391,In_158);
nor U793 (N_793,In_741,N_52);
or U794 (N_794,N_544,In_1719);
xnor U795 (N_795,N_57,In_2118);
and U796 (N_796,N_385,In_226);
and U797 (N_797,In_1810,In_1763);
xor U798 (N_798,N_505,In_1493);
nor U799 (N_799,In_2705,In_2685);
or U800 (N_800,In_2921,N_264);
and U801 (N_801,In_965,In_2219);
nand U802 (N_802,In_2603,In_2720);
xor U803 (N_803,In_133,In_183);
nand U804 (N_804,N_485,In_536);
nand U805 (N_805,In_1217,In_2422);
or U806 (N_806,In_772,In_2028);
nand U807 (N_807,N_146,In_2319);
nand U808 (N_808,In_1146,In_439);
nor U809 (N_809,In_2620,In_807);
nand U810 (N_810,In_1066,In_2420);
nor U811 (N_811,In_2851,In_240);
and U812 (N_812,In_1701,In_1858);
and U813 (N_813,In_2084,In_1312);
nor U814 (N_814,In_1930,In_2381);
nand U815 (N_815,N_558,In_2984);
or U816 (N_816,In_1196,In_135);
nor U817 (N_817,N_492,In_373);
xnor U818 (N_818,In_1046,N_566);
or U819 (N_819,In_2388,In_19);
or U820 (N_820,In_2570,In_250);
nor U821 (N_821,N_411,In_905);
nand U822 (N_822,In_1541,In_474);
or U823 (N_823,In_805,N_529);
or U824 (N_824,In_1501,In_685);
or U825 (N_825,N_550,In_83);
nor U826 (N_826,In_1029,In_2245);
nand U827 (N_827,In_925,In_1809);
and U828 (N_828,In_1439,In_1717);
xor U829 (N_829,In_2617,In_1649);
xnor U830 (N_830,In_1075,In_2790);
or U831 (N_831,In_1390,N_524);
or U832 (N_832,In_1169,N_3);
or U833 (N_833,In_1543,In_2521);
or U834 (N_834,In_2022,In_1405);
xnor U835 (N_835,N_113,In_1806);
xor U836 (N_836,In_115,In_482);
nand U837 (N_837,In_1448,In_2828);
nor U838 (N_838,In_837,In_1299);
and U839 (N_839,In_1191,In_296);
or U840 (N_840,N_332,In_1586);
nand U841 (N_841,N_424,N_105);
xnor U842 (N_842,In_2600,In_1099);
or U843 (N_843,In_1973,In_2933);
or U844 (N_844,N_115,In_1546);
nor U845 (N_845,In_574,N_406);
nand U846 (N_846,In_2956,In_1051);
nor U847 (N_847,In_472,N_453);
nand U848 (N_848,In_879,In_1881);
nor U849 (N_849,In_452,N_93);
or U850 (N_850,In_2334,In_2275);
or U851 (N_851,N_212,N_331);
nand U852 (N_852,In_1752,In_409);
and U853 (N_853,N_577,N_346);
nand U854 (N_854,In_564,In_2244);
xor U855 (N_855,In_1911,In_2980);
nor U856 (N_856,In_915,N_12);
and U857 (N_857,In_2010,In_2759);
nor U858 (N_858,N_467,N_265);
nor U859 (N_859,N_51,In_2987);
xnor U860 (N_860,N_48,N_326);
xor U861 (N_861,In_243,In_2225);
xnor U862 (N_862,N_433,In_2787);
nand U863 (N_863,In_937,In_861);
nor U864 (N_864,In_1982,N_425);
or U865 (N_865,In_1331,In_1638);
or U866 (N_866,In_405,In_2071);
nand U867 (N_867,In_2404,N_270);
and U868 (N_868,In_1778,In_477);
or U869 (N_869,In_188,In_1247);
xnor U870 (N_870,In_1220,In_145);
xor U871 (N_871,In_2526,In_1659);
xor U872 (N_872,In_2611,In_2859);
or U873 (N_873,In_1414,In_2452);
nor U874 (N_874,In_576,In_368);
or U875 (N_875,In_1138,In_2309);
nand U876 (N_876,In_169,In_337);
nand U877 (N_877,N_20,In_2960);
nor U878 (N_878,In_582,N_65);
xor U879 (N_879,In_2469,In_330);
nand U880 (N_880,N_598,In_2545);
nand U881 (N_881,In_539,In_661);
and U882 (N_882,In_1246,In_1596);
and U883 (N_883,In_2911,In_230);
nand U884 (N_884,N_169,N_445);
or U885 (N_885,N_180,N_245);
or U886 (N_886,In_2722,In_143);
nand U887 (N_887,N_252,N_472);
nand U888 (N_888,N_137,N_192);
nor U889 (N_889,In_1745,In_361);
nor U890 (N_890,In_854,In_2141);
and U891 (N_891,In_1978,In_276);
and U892 (N_892,In_1480,In_1966);
and U893 (N_893,In_1328,In_2406);
xnor U894 (N_894,N_495,In_968);
nand U895 (N_895,In_1579,In_1384);
nand U896 (N_896,In_362,In_2099);
nand U897 (N_897,In_381,In_2724);
nor U898 (N_898,N_545,In_696);
nor U899 (N_899,In_69,N_504);
and U900 (N_900,N_152,N_9);
xor U901 (N_901,In_2158,In_1300);
or U902 (N_902,In_2978,In_873);
nand U903 (N_903,In_1382,In_519);
xnor U904 (N_904,N_256,In_2479);
xor U905 (N_905,In_784,In_680);
nor U906 (N_906,N_31,N_443);
nor U907 (N_907,N_262,N_0);
nand U908 (N_908,N_280,In_2742);
nand U909 (N_909,N_89,N_477);
and U910 (N_910,In_2940,In_1529);
or U911 (N_911,N_350,In_1716);
nand U912 (N_912,N_412,N_288);
xor U913 (N_913,N_432,N_336);
nor U914 (N_914,In_2027,N_575);
or U915 (N_915,In_1651,In_1566);
or U916 (N_916,In_2380,N_496);
xnor U917 (N_917,N_390,In_353);
or U918 (N_918,N_103,In_2345);
and U919 (N_919,In_325,In_2402);
and U920 (N_920,In_2761,In_2053);
or U921 (N_921,In_1281,In_1227);
nand U922 (N_922,In_1097,In_2551);
or U923 (N_923,N_474,In_2337);
xnor U924 (N_924,In_2190,In_2536);
or U925 (N_925,N_464,N_519);
nor U926 (N_926,N_13,N_533);
nor U927 (N_927,In_2076,N_413);
and U928 (N_928,In_217,In_2114);
nand U929 (N_929,In_648,N_240);
and U930 (N_930,In_1463,In_2885);
or U931 (N_931,In_1377,In_460);
nor U932 (N_932,In_498,In_1219);
nand U933 (N_933,In_1342,In_156);
xor U934 (N_934,N_510,In_57);
nand U935 (N_935,In_2054,In_2544);
xnor U936 (N_936,In_2048,N_208);
nor U937 (N_937,In_600,N_305);
xnor U938 (N_938,In_2730,In_2816);
or U939 (N_939,In_972,N_236);
xor U940 (N_940,In_1440,In_1519);
nand U941 (N_941,In_950,N_493);
and U942 (N_942,N_68,In_26);
nand U943 (N_943,In_573,In_424);
xnor U944 (N_944,N_149,N_217);
nand U945 (N_945,In_610,In_2857);
or U946 (N_946,In_154,N_553);
and U947 (N_947,In_588,In_324);
nand U948 (N_948,In_2605,In_992);
nor U949 (N_949,N_248,In_834);
and U950 (N_950,N_293,In_2079);
nor U951 (N_951,N_261,In_2650);
or U952 (N_952,In_342,In_2680);
nor U953 (N_953,In_2712,In_126);
and U954 (N_954,In_2282,In_596);
nor U955 (N_955,N_186,In_2);
or U956 (N_956,In_1243,In_2976);
nor U957 (N_957,In_1140,In_29);
nand U958 (N_958,In_1174,N_509);
and U959 (N_959,In_2183,In_2000);
or U960 (N_960,In_2652,In_1962);
and U961 (N_961,In_1363,In_1181);
and U962 (N_962,N_237,In_2564);
xnor U963 (N_963,N_207,In_297);
nor U964 (N_964,In_2692,In_899);
or U965 (N_965,In_1036,N_356);
nor U966 (N_966,In_1896,In_2471);
nor U967 (N_967,In_2287,In_1467);
xor U968 (N_968,N_223,In_2299);
and U969 (N_969,N_243,In_585);
xnor U970 (N_970,N_573,In_423);
or U971 (N_971,N_90,N_489);
xor U972 (N_972,N_191,In_2602);
nand U973 (N_973,In_1265,N_225);
xnor U974 (N_974,In_1824,N_2);
nor U975 (N_975,In_1472,In_1276);
xor U976 (N_976,In_2616,N_244);
xnor U977 (N_977,N_232,N_312);
xnor U978 (N_978,In_2305,In_1186);
and U979 (N_979,In_598,In_327);
or U980 (N_980,N_290,N_449);
xnor U981 (N_981,In_640,In_516);
nor U982 (N_982,In_1924,In_1904);
nand U983 (N_983,In_168,In_1804);
nor U984 (N_984,In_2018,In_2967);
or U985 (N_985,In_2009,In_277);
and U986 (N_986,In_2750,In_1690);
or U987 (N_987,N_588,In_990);
nand U988 (N_988,N_286,In_2497);
or U989 (N_989,N_111,In_2896);
nor U990 (N_990,In_928,N_410);
xnor U991 (N_991,In_2697,N_58);
and U992 (N_992,In_1509,In_88);
nand U993 (N_993,N_462,In_1568);
nor U994 (N_994,N_273,In_2184);
nor U995 (N_995,In_719,In_975);
or U996 (N_996,In_2934,In_1592);
xor U997 (N_997,In_2280,In_1160);
nand U998 (N_998,In_2839,In_2841);
nand U999 (N_999,In_1379,In_2496);
xnor U1000 (N_1000,In_1555,In_604);
and U1001 (N_1001,In_1208,N_422);
nand U1002 (N_1002,N_576,In_816);
nand U1003 (N_1003,In_578,In_301);
xnor U1004 (N_1004,In_1994,In_2052);
nor U1005 (N_1005,In_1617,In_1329);
xnor U1006 (N_1006,N_398,N_481);
nor U1007 (N_1007,In_1274,In_1096);
xor U1008 (N_1008,N_499,In_1628);
or U1009 (N_1009,N_501,N_597);
xor U1010 (N_1010,In_1560,In_618);
and U1011 (N_1011,In_1956,In_1527);
and U1012 (N_1012,N_10,In_2211);
nand U1013 (N_1013,In_798,In_1654);
nor U1014 (N_1014,N_289,N_282);
and U1015 (N_1015,In_1113,N_33);
nand U1016 (N_1016,In_836,In_1802);
or U1017 (N_1017,N_11,In_1369);
nand U1018 (N_1018,In_1233,N_66);
xnor U1019 (N_1019,In_2997,In_1031);
or U1020 (N_1020,In_624,N_522);
and U1021 (N_1021,In_1125,In_998);
nand U1022 (N_1022,N_483,In_2837);
xnor U1023 (N_1023,In_537,In_593);
nand U1024 (N_1024,In_2699,In_930);
nand U1025 (N_1025,In_2466,N_364);
xnor U1026 (N_1026,In_1731,N_592);
and U1027 (N_1027,In_104,In_108);
and U1028 (N_1028,In_18,In_2639);
and U1029 (N_1029,In_1686,N_440);
xnor U1030 (N_1030,In_852,In_1507);
nor U1031 (N_1031,In_1672,In_2805);
xor U1032 (N_1032,In_542,In_1677);
or U1033 (N_1033,N_421,In_2169);
and U1034 (N_1034,In_730,In_2628);
nor U1035 (N_1035,In_2666,In_425);
nand U1036 (N_1036,N_490,N_292);
nand U1037 (N_1037,N_235,In_1192);
or U1038 (N_1038,N_221,N_161);
nand U1039 (N_1039,In_2478,In_1178);
nand U1040 (N_1040,In_1232,N_287);
nand U1041 (N_1041,In_2252,In_1705);
nand U1042 (N_1042,In_1608,In_1166);
or U1043 (N_1043,N_150,In_331);
nand U1044 (N_1044,In_2202,N_166);
and U1045 (N_1045,In_39,In_1407);
nand U1046 (N_1046,N_59,In_304);
and U1047 (N_1047,In_2979,In_1150);
nand U1048 (N_1048,N_182,In_718);
nor U1049 (N_1049,In_1244,N_507);
xor U1050 (N_1050,In_2416,In_1109);
nand U1051 (N_1051,In_2575,In_96);
nor U1052 (N_1052,In_1811,In_122);
nand U1053 (N_1053,In_371,In_1689);
and U1054 (N_1054,In_1818,In_1403);
nand U1055 (N_1055,N_176,In_979);
or U1056 (N_1056,In_634,N_134);
and U1057 (N_1057,In_1544,In_492);
and U1058 (N_1058,N_328,N_177);
or U1059 (N_1059,In_2249,N_126);
nand U1060 (N_1060,N_310,N_210);
nand U1061 (N_1061,In_633,N_98);
nor U1062 (N_1062,In_929,In_1042);
nor U1063 (N_1063,In_2063,In_54);
nor U1064 (N_1064,In_1714,N_116);
nand U1065 (N_1065,In_398,In_1372);
and U1066 (N_1066,In_2902,In_1226);
nor U1067 (N_1067,In_2170,In_2130);
xnor U1068 (N_1068,In_204,In_59);
nand U1069 (N_1069,In_2376,N_181);
nand U1070 (N_1070,In_2523,In_1606);
xnor U1071 (N_1071,In_1607,In_761);
nor U1072 (N_1072,In_1656,In_2777);
nor U1073 (N_1073,In_172,In_2532);
xnor U1074 (N_1074,In_864,In_2164);
xnor U1075 (N_1075,In_2576,In_2168);
nor U1076 (N_1076,In_2543,N_219);
xor U1077 (N_1077,N_35,In_418);
or U1078 (N_1078,In_2834,In_1137);
nand U1079 (N_1079,In_2258,N_266);
and U1080 (N_1080,In_1302,N_466);
nand U1081 (N_1081,In_1929,In_2085);
nand U1082 (N_1082,In_2007,In_2250);
and U1083 (N_1083,N_442,In_2172);
nand U1084 (N_1084,In_1549,In_1224);
or U1085 (N_1085,In_1468,In_421);
and U1086 (N_1086,N_164,In_554);
and U1087 (N_1087,In_2599,N_306);
nor U1088 (N_1088,N_171,N_112);
and U1089 (N_1089,In_1098,In_1999);
nor U1090 (N_1090,N_189,In_2832);
nor U1091 (N_1091,In_1536,N_15);
xnor U1092 (N_1092,In_1667,In_1023);
and U1093 (N_1093,In_1135,N_172);
and U1094 (N_1094,In_1353,In_2204);
nor U1095 (N_1095,N_402,N_158);
xor U1096 (N_1096,In_969,In_2791);
nand U1097 (N_1097,N_401,In_1059);
and U1098 (N_1098,N_383,In_2798);
xor U1099 (N_1099,In_2716,In_285);
nand U1100 (N_1100,In_1855,In_76);
xor U1101 (N_1101,In_827,N_317);
or U1102 (N_1102,In_1418,N_384);
nor U1103 (N_1103,N_596,In_2240);
and U1104 (N_1104,In_1420,In_92);
xnor U1105 (N_1105,In_1545,In_876);
nand U1106 (N_1106,In_227,In_403);
and U1107 (N_1107,In_1574,In_1337);
xor U1108 (N_1108,In_2904,In_1202);
nand U1109 (N_1109,N_579,In_1613);
nor U1110 (N_1110,N_321,In_2291);
nand U1111 (N_1111,In_2601,N_78);
xnor U1112 (N_1112,In_1283,N_405);
nor U1113 (N_1113,In_2900,In_2513);
nand U1114 (N_1114,In_1836,N_209);
or U1115 (N_1115,In_2581,In_1054);
nor U1116 (N_1116,In_1003,N_429);
or U1117 (N_1117,N_147,In_906);
and U1118 (N_1118,N_534,N_374);
and U1119 (N_1119,In_1741,In_1020);
nor U1120 (N_1120,In_1164,N_23);
and U1121 (N_1121,In_2342,In_89);
or U1122 (N_1122,N_382,In_1912);
and U1123 (N_1123,N_454,In_281);
or U1124 (N_1124,N_133,In_2490);
nand U1125 (N_1125,In_2145,In_1779);
nor U1126 (N_1126,In_627,In_1373);
xor U1127 (N_1127,N_74,In_941);
and U1128 (N_1128,In_1258,In_2423);
nand U1129 (N_1129,In_2181,In_2595);
xnor U1130 (N_1130,In_728,In_675);
nor U1131 (N_1131,N_203,In_651);
nor U1132 (N_1132,N_319,In_829);
xnor U1133 (N_1133,N_463,In_309);
xnor U1134 (N_1134,In_377,In_2033);
nor U1135 (N_1135,In_2810,In_259);
nand U1136 (N_1136,In_825,N_388);
xnor U1137 (N_1137,In_1830,In_2135);
or U1138 (N_1138,In_1019,In_2194);
or U1139 (N_1139,In_2829,N_100);
nand U1140 (N_1140,In_375,In_2585);
and U1141 (N_1141,In_2916,In_2373);
xor U1142 (N_1142,In_2884,N_64);
and U1143 (N_1143,N_580,N_136);
xor U1144 (N_1144,In_2771,In_803);
nor U1145 (N_1145,In_340,In_642);
or U1146 (N_1146,In_813,In_2445);
nor U1147 (N_1147,In_178,In_559);
or U1148 (N_1148,In_1981,In_794);
and U1149 (N_1149,N_196,In_2676);
or U1150 (N_1150,In_2848,In_1669);
nor U1151 (N_1151,In_10,In_2776);
and U1152 (N_1152,In_909,In_2858);
nand U1153 (N_1153,N_502,In_1461);
xor U1154 (N_1154,In_1158,In_1688);
xnor U1155 (N_1155,In_2721,In_2246);
xnor U1156 (N_1156,In_1792,In_468);
and U1157 (N_1157,In_2475,In_23);
nand U1158 (N_1158,In_64,In_963);
nand U1159 (N_1159,N_216,In_2796);
nor U1160 (N_1160,In_1580,In_1787);
nor U1161 (N_1161,In_1236,In_1310);
or U1162 (N_1162,N_22,In_2983);
xor U1163 (N_1163,In_33,N_518);
nor U1164 (N_1164,In_258,In_476);
xnor U1165 (N_1165,In_1587,N_556);
xor U1166 (N_1166,In_1022,N_316);
nor U1167 (N_1167,N_241,In_2826);
nor U1168 (N_1168,N_527,In_635);
xnor U1169 (N_1169,In_2931,N_92);
nand U1170 (N_1170,In_497,N_460);
nand U1171 (N_1171,In_2533,N_253);
nand U1172 (N_1172,In_788,In_1380);
and U1173 (N_1173,N_278,In_1775);
nor U1174 (N_1174,In_1925,In_2121);
xnor U1175 (N_1175,In_84,In_2398);
and U1176 (N_1176,In_764,N_5);
xor U1177 (N_1177,N_515,In_1572);
or U1178 (N_1178,In_704,In_2064);
nor U1179 (N_1179,N_377,In_1603);
and U1180 (N_1180,In_443,In_2681);
or U1181 (N_1181,In_2855,In_1355);
or U1182 (N_1182,In_1846,In_475);
xor U1183 (N_1183,In_396,In_404);
and U1184 (N_1184,In_1776,In_1005);
nor U1185 (N_1185,In_1490,In_1159);
nor U1186 (N_1186,In_2060,N_397);
and U1187 (N_1187,In_2590,In_702);
nor U1188 (N_1188,In_91,In_1344);
nand U1189 (N_1189,In_647,N_87);
and U1190 (N_1190,In_1212,In_530);
or U1191 (N_1191,In_1239,In_2001);
xor U1192 (N_1192,In_1584,In_1114);
and U1193 (N_1193,In_1502,N_450);
and U1194 (N_1194,In_2485,In_1952);
nand U1195 (N_1195,In_1887,In_211);
nor U1196 (N_1196,In_363,In_927);
nor U1197 (N_1197,N_408,In_2449);
or U1198 (N_1198,In_235,In_2645);
nand U1199 (N_1199,In_510,In_491);
nand U1200 (N_1200,In_1997,In_1025);
nor U1201 (N_1201,N_981,In_1957);
and U1202 (N_1202,In_2819,In_2815);
and U1203 (N_1203,In_2456,In_1834);
and U1204 (N_1204,N_1183,N_391);
nand U1205 (N_1205,In_151,In_273);
nand U1206 (N_1206,N_882,In_2782);
nor U1207 (N_1207,In_1749,In_2924);
and U1208 (N_1208,N_251,N_455);
and U1209 (N_1209,N_1043,In_1757);
nand U1210 (N_1210,N_367,In_432);
xnor U1211 (N_1211,In_897,In_1637);
nand U1212 (N_1212,N_379,In_2310);
nand U1213 (N_1213,In_2120,In_1698);
and U1214 (N_1214,N_145,N_826);
nand U1215 (N_1215,In_1343,N_129);
nor U1216 (N_1216,N_1128,In_1955);
nor U1217 (N_1217,N_996,In_2903);
or U1218 (N_1218,In_165,In_2350);
xnor U1219 (N_1219,N_788,N_655);
xnor U1220 (N_1220,In_1851,N_1074);
and U1221 (N_1221,In_515,In_830);
or U1222 (N_1222,N_1152,In_1476);
or U1223 (N_1223,In_779,In_900);
and U1224 (N_1224,N_600,In_2180);
nand U1225 (N_1225,In_117,In_2708);
nor U1226 (N_1226,N_718,In_2408);
xor U1227 (N_1227,N_776,N_848);
or U1228 (N_1228,In_1614,In_2783);
or U1229 (N_1229,N_1119,In_1423);
nor U1230 (N_1230,N_955,N_21);
and U1231 (N_1231,In_1143,In_538);
xor U1232 (N_1232,In_2390,N_142);
or U1233 (N_1233,N_295,In_804);
nor U1234 (N_1234,N_322,In_2920);
nor U1235 (N_1235,N_155,N_206);
and U1236 (N_1236,In_1950,In_1515);
nor U1237 (N_1237,In_1658,N_712);
and U1238 (N_1238,In_113,In_2488);
nor U1239 (N_1239,N_1137,N_971);
or U1240 (N_1240,In_1216,In_743);
or U1241 (N_1241,In_1967,N_807);
and U1242 (N_1242,N_844,N_891);
nand U1243 (N_1243,In_847,N_985);
nor U1244 (N_1244,In_1419,N_865);
and U1245 (N_1245,In_2632,N_615);
xor U1246 (N_1246,In_1793,N_915);
nor U1247 (N_1247,In_2268,In_2981);
and U1248 (N_1248,In_1798,In_850);
nand U1249 (N_1249,In_2723,N_920);
xnor U1250 (N_1250,N_1085,N_1009);
and U1251 (N_1251,N_202,N_298);
nand U1252 (N_1252,N_373,In_414);
xnor U1253 (N_1253,In_1984,N_81);
nand U1254 (N_1254,N_85,N_394);
and U1255 (N_1255,N_999,N_876);
xnor U1256 (N_1256,In_592,In_180);
xnor U1257 (N_1257,N_109,N_751);
nor U1258 (N_1258,In_2669,N_1091);
nor U1259 (N_1259,N_430,N_1070);
and U1260 (N_1260,N_353,N_717);
and U1261 (N_1261,In_161,N_966);
xor U1262 (N_1262,N_104,In_395);
nor U1263 (N_1263,N_564,N_685);
and U1264 (N_1264,In_2754,N_590);
nor U1265 (N_1265,In_781,In_1474);
nor U1266 (N_1266,In_2515,In_1605);
nor U1267 (N_1267,N_418,In_2176);
nor U1268 (N_1268,N_683,In_41);
nor U1269 (N_1269,N_780,In_2325);
and U1270 (N_1270,N_799,N_1122);
nor U1271 (N_1271,In_999,In_1431);
nor U1272 (N_1272,N_759,In_2279);
or U1273 (N_1273,In_129,In_878);
nor U1274 (N_1274,In_2412,N_461);
and U1275 (N_1275,In_2850,N_569);
or U1276 (N_1276,N_347,N_1156);
xor U1277 (N_1277,N_649,In_1722);
nor U1278 (N_1278,N_360,In_314);
and U1279 (N_1279,In_926,N_348);
nand U1280 (N_1280,In_2262,In_397);
xor U1281 (N_1281,In_1371,N_1109);
or U1282 (N_1282,In_1048,In_1983);
nand U1283 (N_1283,In_1784,N_902);
xor U1284 (N_1284,N_819,In_294);
or U1285 (N_1285,N_178,In_448);
nor U1286 (N_1286,N_1026,In_2313);
nor U1287 (N_1287,In_1576,In_2335);
and U1288 (N_1288,In_388,In_2454);
nand U1289 (N_1289,In_2527,In_1210);
nor U1290 (N_1290,In_1259,N_743);
xnor U1291 (N_1291,N_965,N_1101);
and U1292 (N_1292,N_810,N_386);
or U1293 (N_1293,N_95,N_523);
xor U1294 (N_1294,In_2019,In_2922);
and U1295 (N_1295,In_392,N_719);
xnor U1296 (N_1296,N_1098,In_170);
or U1297 (N_1297,N_1176,In_2016);
or U1298 (N_1298,N_633,N_291);
and U1299 (N_1299,N_986,In_1086);
xnor U1300 (N_1300,N_1158,In_1675);
nand U1301 (N_1301,In_1491,In_255);
and U1302 (N_1302,In_2450,N_541);
nand U1303 (N_1303,In_0,N_885);
nand U1304 (N_1304,N_121,N_1093);
xor U1305 (N_1305,N_830,N_71);
nand U1306 (N_1306,N_944,N_1067);
and U1307 (N_1307,In_214,N_341);
or U1308 (N_1308,In_1794,In_1314);
nor U1309 (N_1309,N_949,N_838);
xor U1310 (N_1310,In_886,In_755);
or U1311 (N_1311,In_2178,N_903);
nor U1312 (N_1312,N_1036,In_1875);
nor U1313 (N_1313,In_2093,In_1072);
xor U1314 (N_1314,N_907,In_2396);
or U1315 (N_1315,In_625,N_194);
or U1316 (N_1316,N_1102,N_849);
nand U1317 (N_1317,In_2684,N_959);
and U1318 (N_1318,In_1993,N_1112);
nor U1319 (N_1319,N_684,N_923);
or U1320 (N_1320,N_994,In_2430);
nor U1321 (N_1321,In_951,In_555);
nor U1322 (N_1322,N_1117,In_1524);
xor U1323 (N_1323,N_804,N_675);
and U1324 (N_1324,N_893,N_619);
nand U1325 (N_1325,N_653,N_957);
or U1326 (N_1326,N_120,In_1017);
xnor U1327 (N_1327,In_891,In_2041);
xor U1328 (N_1328,N_250,N_1058);
nand U1329 (N_1329,In_1110,In_350);
nor U1330 (N_1330,In_2757,In_1052);
nand U1331 (N_1331,N_139,N_945);
or U1332 (N_1332,N_79,N_1180);
xnor U1333 (N_1333,N_982,N_1167);
xor U1334 (N_1334,In_1008,N_439);
xnor U1335 (N_1335,N_839,In_1933);
xnor U1336 (N_1336,In_1825,In_1376);
nor U1337 (N_1337,In_1068,N_710);
xor U1338 (N_1338,In_1067,N_730);
and U1339 (N_1339,N_868,In_622);
xnor U1340 (N_1340,N_809,In_2734);
nor U1341 (N_1341,N_928,N_796);
nor U1342 (N_1342,In_595,In_955);
and U1343 (N_1343,N_637,N_837);
nand U1344 (N_1344,N_695,In_441);
nand U1345 (N_1345,In_716,In_1152);
or U1346 (N_1346,In_2542,In_2817);
xnor U1347 (N_1347,In_2306,In_2972);
and U1348 (N_1348,N_832,N_227);
xnor U1349 (N_1349,In_2031,In_541);
or U1350 (N_1350,In_310,N_1188);
nor U1351 (N_1351,N_950,N_307);
nor U1352 (N_1352,N_1,In_985);
and U1353 (N_1353,N_696,In_2142);
nand U1354 (N_1354,N_875,N_940);
and U1355 (N_1355,N_762,N_1170);
and U1356 (N_1356,In_305,In_2629);
nand U1357 (N_1357,N_37,N_1135);
xnor U1358 (N_1358,In_2101,N_659);
xor U1359 (N_1359,N_571,N_260);
xnor U1360 (N_1360,N_447,N_127);
and U1361 (N_1361,N_444,N_1145);
xnor U1362 (N_1362,In_1338,In_197);
xnor U1363 (N_1363,N_437,In_2215);
nand U1364 (N_1364,In_2457,N_763);
or U1365 (N_1365,N_888,N_642);
nor U1366 (N_1366,N_1104,In_616);
and U1367 (N_1367,N_878,N_625);
or U1368 (N_1368,N_301,In_2265);
or U1369 (N_1369,In_2906,In_2998);
nand U1370 (N_1370,N_737,N_528);
xor U1371 (N_1371,In_13,In_1119);
or U1372 (N_1372,In_1357,In_867);
nand U1373 (N_1373,In_1898,In_1237);
nand U1374 (N_1374,In_2809,N_654);
nand U1375 (N_1375,N_991,In_550);
xor U1376 (N_1376,N_188,N_4);
nand U1377 (N_1377,N_1132,N_980);
and U1378 (N_1378,In_1151,N_1189);
and U1379 (N_1379,N_1120,N_842);
or U1380 (N_1380,N_315,In_1895);
and U1381 (N_1381,N_1127,In_2340);
nand U1382 (N_1382,In_34,N_500);
nand U1383 (N_1383,N_783,In_2026);
xnor U1384 (N_1384,In_1928,In_322);
and U1385 (N_1385,N_30,N_1125);
xnor U1386 (N_1386,In_565,In_2371);
nand U1387 (N_1387,N_254,N_860);
nor U1388 (N_1388,In_1791,In_2294);
nand U1389 (N_1389,N_448,N_843);
xor U1390 (N_1390,N_829,In_1547);
and U1391 (N_1391,N_419,N_665);
and U1392 (N_1392,In_1516,N_338);
xor U1393 (N_1393,N_1029,N_297);
xor U1394 (N_1394,N_1092,N_742);
nand U1395 (N_1395,N_1038,N_884);
and U1396 (N_1396,N_933,In_1604);
xor U1397 (N_1397,N_828,In_1375);
nand U1398 (N_1398,N_774,In_2185);
xnor U1399 (N_1399,In_673,N_960);
xor U1400 (N_1400,N_1065,N_294);
nand U1401 (N_1401,N_947,N_355);
or U1402 (N_1402,In_1788,N_1050);
nand U1403 (N_1403,In_572,In_2647);
nor U1404 (N_1404,In_783,N_648);
or U1405 (N_1405,N_1052,N_822);
and U1406 (N_1406,N_632,In_792);
xnor U1407 (N_1407,N_1163,In_746);
nand U1408 (N_1408,In_603,In_1055);
nor U1409 (N_1409,In_453,In_2691);
nand U1410 (N_1410,In_2487,In_2014);
nand U1411 (N_1411,In_159,In_2401);
or U1412 (N_1412,In_887,N_855);
or U1413 (N_1413,N_680,N_1186);
and U1414 (N_1414,In_1177,In_2671);
and U1415 (N_1415,In_1979,In_1489);
or U1416 (N_1416,In_2524,In_2267);
nor U1417 (N_1417,N_931,N_881);
and U1418 (N_1418,In_1551,N_792);
xnor U1419 (N_1419,In_2640,In_1402);
nor U1420 (N_1420,N_258,In_2659);
nand U1421 (N_1421,In_2580,N_456);
and U1422 (N_1422,In_2556,In_1229);
or U1423 (N_1423,In_2818,N_91);
and U1424 (N_1424,In_1662,In_2067);
nand U1425 (N_1425,N_997,In_2327);
nand U1426 (N_1426,In_267,In_2468);
nor U1427 (N_1427,N_818,N_431);
and U1428 (N_1428,In_522,N_414);
and U1429 (N_1429,In_2925,In_2586);
and U1430 (N_1430,In_1462,N_901);
or U1431 (N_1431,In_2106,In_99);
and U1432 (N_1432,In_7,N_1113);
and U1433 (N_1433,In_1044,N_820);
xor U1434 (N_1434,In_427,In_2119);
nor U1435 (N_1435,In_1002,N_604);
and U1436 (N_1436,N_465,In_2421);
nand U1437 (N_1437,In_1640,In_2152);
nand U1438 (N_1438,N_488,N_1182);
nand U1439 (N_1439,N_752,N_7);
nor U1440 (N_1440,In_2251,N_793);
or U1441 (N_1441,N_821,N_1154);
nand U1442 (N_1442,N_1168,N_894);
xnor U1443 (N_1443,N_1010,In_1538);
or U1444 (N_1444,In_1891,In_1559);
nor U1445 (N_1445,In_2889,N_324);
or U1446 (N_1446,N_797,In_134);
or U1447 (N_1447,N_769,N_135);
and U1448 (N_1448,N_1006,In_480);
or U1449 (N_1449,N_911,N_702);
xor U1450 (N_1450,In_981,N_1160);
nand U1451 (N_1451,In_851,In_703);
or U1452 (N_1452,In_1581,N_948);
or U1453 (N_1453,N_857,N_1042);
and U1454 (N_1454,In_1864,N_1048);
or U1455 (N_1455,N_1021,N_1086);
xnor U1456 (N_1456,In_1473,In_1438);
xor U1457 (N_1457,N_1016,In_2775);
xnor U1458 (N_1458,In_1630,N_660);
nor U1459 (N_1459,N_932,In_2243);
nor U1460 (N_1460,In_1720,N_1077);
nand U1461 (N_1461,In_1583,In_346);
and U1462 (N_1462,N_993,N_1136);
and U1463 (N_1463,In_1567,N_1164);
and U1464 (N_1464,In_2320,N_458);
nand U1465 (N_1465,In_908,In_561);
nand U1466 (N_1466,N_778,N_897);
or U1467 (N_1467,In_2969,N_883);
and U1468 (N_1468,In_1179,In_2893);
nor U1469 (N_1469,In_1396,N_1097);
xnor U1470 (N_1470,In_768,N_977);
or U1471 (N_1471,In_1487,In_1682);
nand U1472 (N_1472,In_20,N_741);
nor U1473 (N_1473,In_776,N_378);
and U1474 (N_1474,N_721,N_617);
xnor U1475 (N_1475,N_552,N_1171);
xnor U1476 (N_1476,N_674,In_2768);
nor U1477 (N_1477,In_1433,In_429);
and U1478 (N_1478,N_917,N_187);
nor U1479 (N_1479,In_1723,In_1764);
nand U1480 (N_1480,In_619,N_47);
or U1481 (N_1481,In_2690,N_88);
or U1482 (N_1482,N_708,N_86);
nand U1483 (N_1483,In_2505,In_245);
or U1484 (N_1484,In_2550,In_662);
or U1485 (N_1485,N_403,In_1550);
and U1486 (N_1486,In_2588,N_163);
nor U1487 (N_1487,In_2892,N_470);
or U1488 (N_1488,N_532,N_417);
nand U1489 (N_1489,In_241,N_641);
or U1490 (N_1490,N_816,N_658);
and U1491 (N_1491,In_1092,In_1185);
nor U1492 (N_1492,In_1093,N_678);
or U1493 (N_1493,In_35,In_1316);
and U1494 (N_1494,N_899,N_1115);
and U1495 (N_1495,N_896,N_777);
and U1496 (N_1496,In_1996,In_880);
xor U1497 (N_1497,N_765,N_1088);
nor U1498 (N_1498,N_1060,In_855);
xnor U1499 (N_1499,In_359,N_802);
xor U1500 (N_1500,N_128,N_1118);
xor U1501 (N_1501,In_249,In_1120);
or U1502 (N_1502,In_1505,In_2239);
nor U1503 (N_1503,N_616,N_968);
nor U1504 (N_1504,In_2160,In_2625);
nor U1505 (N_1505,In_263,N_930);
xor U1506 (N_1506,N_851,In_36);
nor U1507 (N_1507,N_239,N_824);
or U1508 (N_1508,In_2347,N_329);
nand U1509 (N_1509,In_1282,N_634);
nor U1510 (N_1510,N_998,N_840);
xnor U1511 (N_1511,In_1715,N_511);
xor U1512 (N_1512,In_446,In_1056);
nor U1513 (N_1513,N_123,N_874);
or U1514 (N_1514,N_226,N_701);
xor U1515 (N_1515,In_2702,In_2269);
nor U1516 (N_1516,In_2113,In_1743);
nor U1517 (N_1517,N_376,In_456);
nor U1518 (N_1518,N_118,N_937);
nor U1519 (N_1519,N_117,In_1416);
nor U1520 (N_1520,In_2912,N_1133);
nand U1521 (N_1521,N_669,In_527);
nor U1522 (N_1522,In_1327,N_938);
xnor U1523 (N_1523,N_935,In_2293);
nand U1524 (N_1524,In_2959,N_880);
and U1525 (N_1525,In_1187,In_1873);
or U1526 (N_1526,N_1039,In_606);
nor U1527 (N_1527,N_1114,N_1131);
nand U1528 (N_1528,In_2677,N_676);
nor U1529 (N_1529,N_1150,N_895);
or U1530 (N_1530,N_733,In_348);
nand U1531 (N_1531,In_1028,In_2836);
xnor U1532 (N_1532,N_513,In_320);
nand U1533 (N_1533,In_2845,In_924);
xnor U1534 (N_1534,In_2349,N_1165);
xor U1535 (N_1535,N_1055,N_916);
nand U1536 (N_1536,N_69,In_1909);
xor U1537 (N_1537,N_1096,In_948);
nor U1538 (N_1538,N_815,In_2264);
and U1539 (N_1539,In_1533,N_732);
xor U1540 (N_1540,In_1147,In_284);
and U1541 (N_1541,In_534,In_1449);
nand U1542 (N_1542,N_1138,N_49);
xnor U1543 (N_1543,In_2355,N_572);
xor U1544 (N_1544,N_766,In_479);
nor U1545 (N_1545,N_795,In_2284);
nand U1546 (N_1546,N_72,N_18);
and U1547 (N_1547,N_629,N_662);
xnor U1548 (N_1548,In_2755,N_671);
xnor U1549 (N_1549,N_1107,N_740);
and U1550 (N_1550,N_750,N_808);
or U1551 (N_1551,In_2254,In_1713);
nand U1552 (N_1552,N_647,N_814);
nor U1553 (N_1553,In_697,N_611);
xor U1554 (N_1554,In_202,In_2709);
nor U1555 (N_1555,In_417,In_1768);
nand U1556 (N_1556,N_559,In_2303);
nor U1557 (N_1557,N_831,In_2324);
and U1558 (N_1558,N_1106,N_589);
nor U1559 (N_1559,In_2301,In_90);
nand U1560 (N_1560,N_817,N_549);
or U1561 (N_1561,In_504,In_1901);
xnor U1562 (N_1562,N_767,N_946);
xnor U1563 (N_1563,N_557,In_2186);
xnor U1564 (N_1564,N_835,In_1683);
nor U1565 (N_1565,In_1007,In_1548);
nor U1566 (N_1566,In_2918,N_705);
xor U1567 (N_1567,N_958,In_2029);
xor U1568 (N_1568,In_2230,In_319);
nor U1569 (N_1569,In_2953,N_416);
or U1570 (N_1570,N_622,In_1427);
and U1571 (N_1571,In_2812,N_988);
nand U1572 (N_1572,N_1149,N_630);
or U1573 (N_1573,N_1053,N_790);
xnor U1574 (N_1574,N_1130,N_723);
nand U1575 (N_1575,N_636,In_1294);
nand U1576 (N_1576,In_379,In_130);
or U1577 (N_1577,In_2877,N_67);
xor U1578 (N_1578,In_706,N_961);
or U1579 (N_1579,N_628,N_919);
nor U1580 (N_1580,N_1047,In_2132);
or U1581 (N_1581,In_1565,N_627);
or U1582 (N_1582,In_1139,N_344);
nor U1583 (N_1583,In_2332,In_1004);
and U1584 (N_1584,N_801,In_2448);
xor U1585 (N_1585,In_875,N_102);
xnor U1586 (N_1586,N_1193,N_963);
nand U1587 (N_1587,N_587,N_451);
and U1588 (N_1588,N_646,In_1621);
or U1589 (N_1589,In_2277,In_81);
nor U1590 (N_1590,In_2199,In_1074);
nor U1591 (N_1591,N_805,In_440);
nand U1592 (N_1592,In_1678,In_1866);
nand U1593 (N_1593,N_1017,In_857);
and U1594 (N_1594,N_995,N_539);
nor U1595 (N_1595,N_581,In_1336);
nand U1596 (N_1596,In_1990,N_1166);
and U1597 (N_1597,N_927,N_936);
xnor U1598 (N_1598,N_972,In_1381);
xnor U1599 (N_1599,In_378,N_806);
nor U1600 (N_1600,N_60,In_190);
and U1601 (N_1601,N_131,In_189);
or U1602 (N_1602,In_713,In_2729);
and U1603 (N_1603,In_740,In_2200);
nand U1604 (N_1604,In_2107,In_2764);
nor U1605 (N_1605,N_1178,N_220);
or U1606 (N_1606,N_823,In_773);
xor U1607 (N_1607,N_1089,N_601);
and U1608 (N_1608,N_1181,In_2439);
nand U1609 (N_1609,N_1173,In_920);
or U1610 (N_1610,In_1601,In_2679);
nand U1611 (N_1611,N_1035,N_1033);
or U1612 (N_1612,N_1005,N_715);
or U1613 (N_1613,In_2451,N_682);
nand U1614 (N_1614,In_1624,N_781);
xnor U1615 (N_1615,N_858,In_1786);
xnor U1616 (N_1616,In_1805,In_528);
nand U1617 (N_1617,In_2159,N_351);
nor U1618 (N_1618,In_1609,In_1882);
nor U1619 (N_1619,In_490,N_46);
nand U1620 (N_1620,N_1198,N_476);
nand U1621 (N_1621,In_777,N_727);
xnor U1622 (N_1622,In_1872,N_934);
xnor U1623 (N_1623,N_6,In_1441);
nand U1624 (N_1624,In_382,In_710);
or U1625 (N_1625,In_2232,In_2429);
nand U1626 (N_1626,In_1498,N_748);
and U1627 (N_1627,N_1148,N_1174);
nor U1628 (N_1628,N_775,N_1023);
xnor U1629 (N_1629,In_2165,N_56);
nor U1630 (N_1630,N_771,N_904);
nor U1631 (N_1631,N_538,N_130);
nor U1632 (N_1632,N_516,In_2573);
xor U1633 (N_1633,N_108,N_1019);
and U1634 (N_1634,In_2943,In_2073);
or U1635 (N_1635,In_2434,N_1002);
nand U1636 (N_1636,In_2641,In_1920);
and U1637 (N_1637,N_983,In_2571);
nand U1638 (N_1638,In_1905,N_811);
or U1639 (N_1639,In_2733,In_49);
nor U1640 (N_1640,In_2788,N_921);
xor U1641 (N_1641,In_657,In_2008);
nor U1642 (N_1642,In_120,N_640);
and U1643 (N_1643,N_909,In_2415);
nor U1644 (N_1644,N_862,N_749);
or U1645 (N_1645,N_747,In_1880);
nand U1646 (N_1646,N_1187,N_157);
xor U1647 (N_1647,In_923,N_782);
or U1648 (N_1648,In_1530,In_1921);
nor U1649 (N_1649,N_952,N_407);
xnor U1650 (N_1650,N_956,N_753);
xor U1651 (N_1651,In_575,N_892);
nor U1652 (N_1652,N_643,N_27);
and U1653 (N_1653,N_1175,In_2792);
or U1654 (N_1654,In_2634,In_1107);
and U1655 (N_1655,In_1785,In_1495);
or U1656 (N_1656,In_1201,In_1756);
nand U1657 (N_1657,In_652,In_171);
xor U1658 (N_1658,N_420,In_356);
nand U1659 (N_1659,In_2908,N_854);
nor U1660 (N_1660,In_605,N_729);
nand U1661 (N_1661,N_1064,N_1007);
xnor U1662 (N_1662,In_1268,In_1521);
nor U1663 (N_1663,In_1410,In_269);
nor U1664 (N_1664,In_1703,In_2517);
or U1665 (N_1665,N_605,In_1892);
nor U1666 (N_1666,In_32,N_754);
nor U1667 (N_1667,In_2686,In_2162);
xnor U1668 (N_1668,N_595,N_512);
xnor U1669 (N_1669,In_2986,N_798);
nand U1670 (N_1670,In_693,N_1116);
and U1671 (N_1671,In_1385,N_1162);
or U1672 (N_1672,N_1015,In_1456);
and U1673 (N_1673,In_1588,In_2663);
xor U1674 (N_1674,N_1045,N_32);
xor U1675 (N_1675,N_975,In_328);
and U1676 (N_1676,In_256,In_486);
or U1677 (N_1677,N_1062,In_1223);
or U1678 (N_1678,In_1106,N_607);
and U1679 (N_1679,N_834,In_1018);
and U1680 (N_1680,In_1010,In_234);
xor U1681 (N_1681,N_967,N_275);
xor U1682 (N_1682,N_1031,N_1121);
xnor U1683 (N_1683,N_900,In_896);
and U1684 (N_1684,N_1169,In_2662);
nor U1685 (N_1685,In_387,In_138);
nor U1686 (N_1686,N_756,N_725);
nor U1687 (N_1687,In_2786,N_869);
nor U1688 (N_1688,N_540,In_2383);
nand U1689 (N_1689,N_768,In_1746);
nand U1690 (N_1690,N_148,In_2004);
nor U1691 (N_1691,N_1022,N_1095);
xnor U1692 (N_1692,N_308,N_452);
or U1693 (N_1693,N_480,In_2882);
nor U1694 (N_1694,N_850,N_610);
nand U1695 (N_1695,N_716,N_1155);
or U1696 (N_1696,N_664,In_2897);
nand U1697 (N_1697,In_692,N_371);
or U1698 (N_1698,In_1366,In_1694);
or U1699 (N_1699,In_1616,In_1854);
or U1700 (N_1700,In_1954,In_1582);
nand U1701 (N_1701,In_166,In_98);
or U1702 (N_1702,In_2453,N_1003);
or U1703 (N_1703,N_1184,N_357);
xnor U1704 (N_1704,N_255,N_387);
and U1705 (N_1705,N_914,N_978);
or U1706 (N_1706,N_1100,In_1500);
nor U1707 (N_1707,N_939,N_889);
xor U1708 (N_1708,N_143,In_2394);
nand U1709 (N_1709,N_886,In_2801);
or U1710 (N_1710,N_764,In_1);
or U1711 (N_1711,N_602,In_1121);
and U1712 (N_1712,In_1038,In_2784);
nor U1713 (N_1713,N_1140,N_833);
and U1714 (N_1714,In_2583,In_1417);
or U1715 (N_1715,N_666,In_2111);
and U1716 (N_1716,N_1110,N_746);
nor U1717 (N_1717,N_153,N_1194);
or U1718 (N_1718,In_1131,N_567);
nor U1719 (N_1719,In_2087,N_1044);
nand U1720 (N_1720,In_535,In_1998);
and U1721 (N_1721,In_2147,In_471);
nand U1722 (N_1722,N_979,In_464);
nand U1723 (N_1723,In_964,In_238);
nand U1724 (N_1724,N_877,N_1105);
or U1725 (N_1725,N_215,In_1542);
and U1726 (N_1726,N_107,N_1161);
or U1727 (N_1727,N_1069,In_2804);
nor U1728 (N_1728,N_242,In_1902);
nor U1729 (N_1729,N_361,In_408);
nor U1730 (N_1730,In_2005,N_668);
nor U1731 (N_1731,N_1191,N_758);
xnor U1732 (N_1732,In_1907,N_1000);
xor U1733 (N_1733,In_1665,N_974);
xnor U1734 (N_1734,N_761,N_1051);
and U1735 (N_1735,In_2455,N_867);
and U1736 (N_1736,N_249,In_2942);
or U1737 (N_1737,N_677,N_1179);
nand U1738 (N_1738,In_1736,N_698);
nor U1739 (N_1739,In_1951,In_2808);
nor U1740 (N_1740,In_1189,N_827);
nand U1741 (N_1741,In_947,N_724);
nand U1742 (N_1742,In_729,In_833);
nand U1743 (N_1743,N_726,N_1129);
and U1744 (N_1744,N_73,N_1013);
xnor U1745 (N_1745,N_1078,N_1196);
xnor U1746 (N_1746,N_599,N_912);
or U1747 (N_1747,In_1913,In_888);
and U1748 (N_1748,In_46,In_2991);
or U1749 (N_1749,In_53,N_954);
nor U1750 (N_1750,N_274,N_506);
nand U1751 (N_1751,N_1103,In_450);
xnor U1752 (N_1752,N_427,N_84);
or U1753 (N_1753,N_612,In_2385);
or U1754 (N_1754,In_201,In_422);
or U1755 (N_1755,N_1004,In_1352);
nor U1756 (N_1756,In_566,In_27);
or U1757 (N_1757,In_2872,N_309);
and U1758 (N_1758,N_39,In_236);
nand U1759 (N_1759,N_409,In_1968);
or U1760 (N_1760,In_1443,In_1305);
or U1761 (N_1761,In_1273,N_906);
nor U1762 (N_1762,N_325,In_1932);
or U1763 (N_1763,In_1077,In_2040);
nor U1764 (N_1764,N_873,N_1123);
nor U1765 (N_1765,In_1040,N_890);
nor U1766 (N_1766,In_2735,In_2929);
and U1767 (N_1767,N_964,In_1634);
xor U1768 (N_1768,In_810,N_910);
xnor U1769 (N_1769,N_704,In_2392);
or U1770 (N_1770,In_2197,In_336);
nor U1771 (N_1771,In_2880,In_1942);
and U1772 (N_1772,N_365,In_1648);
nor U1773 (N_1773,N_167,N_1056);
and U1774 (N_1774,N_652,In_2372);
nor U1775 (N_1775,In_2514,In_966);
and U1776 (N_1776,N_866,N_399);
or U1777 (N_1777,N_673,N_686);
nor U1778 (N_1778,In_1635,N_929);
nor U1779 (N_1779,In_2482,In_2153);
and U1780 (N_1780,N_168,In_902);
xor U1781 (N_1781,In_1184,N_638);
and U1782 (N_1782,N_352,In_1663);
and U1783 (N_1783,In_128,N_457);
nand U1784 (N_1784,N_1192,N_141);
xnor U1785 (N_1785,In_1155,In_488);
or U1786 (N_1786,N_1063,In_1832);
nor U1787 (N_1787,In_1623,In_2683);
or U1788 (N_1788,In_455,N_561);
and U1789 (N_1789,N_228,In_2464);
xnor U1790 (N_1790,In_872,N_314);
xnor U1791 (N_1791,In_2562,N_521);
xnor U1792 (N_1792,N_323,In_391);
or U1793 (N_1793,N_363,N_1177);
nor U1794 (N_1794,In_1027,N_531);
and U1795 (N_1795,In_483,In_2627);
xor U1796 (N_1796,N_853,N_268);
and U1797 (N_1797,In_2461,N_989);
and U1798 (N_1798,N_263,N_582);
or U1799 (N_1799,N_679,In_2155);
and U1800 (N_1800,N_879,N_1570);
or U1801 (N_1801,In_513,N_1467);
and U1802 (N_1802,N_1153,N_1450);
or U1803 (N_1803,N_1790,N_635);
nor U1804 (N_1804,N_1763,N_1744);
xor U1805 (N_1805,N_29,N_1485);
nand U1806 (N_1806,N_1241,N_1540);
xnor U1807 (N_1807,N_697,N_1754);
or U1808 (N_1808,N_1425,In_714);
nor U1809 (N_1809,N_1779,N_1442);
xnor U1810 (N_1810,In_2738,N_1368);
nor U1811 (N_1811,N_1794,N_1330);
xnor U1812 (N_1812,N_1543,N_1738);
xnor U1813 (N_1813,N_1687,N_1758);
or U1814 (N_1814,N_1317,N_1624);
or U1815 (N_1815,N_1451,N_1632);
xnor U1816 (N_1816,N_1699,N_1698);
nand U1817 (N_1817,In_1195,N_497);
nand U1818 (N_1818,N_626,N_1041);
xnor U1819 (N_1819,N_690,N_1190);
xnor U1820 (N_1820,N_1498,In_118);
xnor U1821 (N_1821,N_1528,N_1567);
xnor U1822 (N_1822,N_1333,N_1487);
and U1823 (N_1823,In_1856,N_786);
nand U1824 (N_1824,In_144,N_1597);
and U1825 (N_1825,In_1837,N_1673);
and U1826 (N_1826,N_1410,In_866);
and U1827 (N_1827,In_1350,N_1761);
nor U1828 (N_1828,N_1374,N_1200);
or U1829 (N_1829,N_1408,N_41);
or U1830 (N_1830,N_1249,N_1008);
nand U1831 (N_1831,N_1709,N_1774);
nand U1832 (N_1832,N_941,In_1479);
nor U1833 (N_1833,N_1367,N_1289);
and U1834 (N_1834,N_1712,In_2403);
xnor U1835 (N_1835,In_2821,N_1586);
and U1836 (N_1836,In_1738,In_663);
xor U1837 (N_1837,N_1310,In_962);
nand U1838 (N_1838,N_426,N_1518);
nand U1839 (N_1839,N_1325,N_159);
nor U1840 (N_1840,N_1716,N_1657);
and U1841 (N_1841,In_789,In_1754);
nand U1842 (N_1842,N_1682,N_1304);
nand U1843 (N_1843,In_2614,In_195);
nand U1844 (N_1844,N_1336,In_1118);
nand U1845 (N_1845,N_1501,N_1395);
and U1846 (N_1846,N_1315,N_1437);
nor U1847 (N_1847,N_1666,In_2751);
xor U1848 (N_1848,N_1380,In_2693);
nor U1849 (N_1849,N_845,N_1722);
xor U1850 (N_1850,N_1458,N_1246);
nor U1851 (N_1851,N_1424,N_547);
xnor U1852 (N_1852,N_1751,N_800);
nor U1853 (N_1853,N_693,N_1211);
and U1854 (N_1854,N_1584,N_1579);
nor U1855 (N_1855,N_990,In_735);
or U1856 (N_1856,N_1678,N_1172);
or U1857 (N_1857,N_1723,In_2868);
xnor U1858 (N_1858,N_1392,N_924);
nor U1859 (N_1859,N_852,In_2842);
or U1860 (N_1860,N_661,N_1688);
nand U1861 (N_1861,N_1219,N_1568);
nor U1862 (N_1862,N_905,In_2011);
and U1863 (N_1863,N_1613,N_1630);
nor U1864 (N_1864,N_913,N_1283);
xor U1865 (N_1865,In_2806,N_574);
and U1866 (N_1866,N_1202,N_1134);
and U1867 (N_1867,N_1775,In_501);
nor U1868 (N_1868,N_1349,N_663);
or U1869 (N_1869,N_1159,N_1476);
nand U1870 (N_1870,In_1890,N_584);
and U1871 (N_1871,N_1555,N_1267);
xnor U1872 (N_1872,N_1468,N_720);
nand U1873 (N_1873,N_1072,N_1411);
xnor U1874 (N_1874,N_1506,N_1469);
or U1875 (N_1875,N_1099,In_2528);
or U1876 (N_1876,N_1252,In_758);
and U1877 (N_1877,N_24,N_1558);
or U1878 (N_1878,N_28,N_606);
and U1879 (N_1879,N_870,N_1565);
nand U1880 (N_1880,In_871,N_1331);
and U1881 (N_1881,N_1282,In_2500);
nand U1882 (N_1882,N_1647,N_1509);
or U1883 (N_1883,In_2143,N_1083);
or U1884 (N_1884,N_1243,In_1883);
xor U1885 (N_1885,N_1535,N_925);
xor U1886 (N_1886,N_728,N_1711);
nand U1887 (N_1887,In_174,N_339);
nor U1888 (N_1888,In_701,In_612);
nor U1889 (N_1889,N_1569,N_631);
xnor U1890 (N_1890,N_1087,N_1554);
and U1891 (N_1891,N_1685,N_1591);
nor U1892 (N_1892,N_1740,N_1212);
nand U1893 (N_1893,In_2947,N_1255);
nor U1894 (N_1894,N_1610,N_1455);
nor U1895 (N_1895,N_1720,N_908);
nand U1896 (N_1896,In_389,N_1596);
xnor U1897 (N_1897,N_1488,N_1585);
or U1898 (N_1898,In_1721,N_1529);
xor U1899 (N_1899,In_2548,N_1435);
xnor U1900 (N_1900,N_1204,N_1332);
nor U1901 (N_1901,N_1542,In_2021);
nand U1902 (N_1902,N_1146,N_1522);
or U1903 (N_1903,N_1385,N_841);
nor U1904 (N_1904,N_1226,N_621);
and U1905 (N_1905,N_551,N_1661);
and U1906 (N_1906,N_201,N_1733);
and U1907 (N_1907,N_1111,In_1629);
nor U1908 (N_1908,N_1718,N_1553);
or U1909 (N_1909,N_1735,In_744);
nand U1910 (N_1910,N_1572,N_1571);
nor U1911 (N_1911,N_1314,N_395);
xor U1912 (N_1912,N_1372,In_785);
or U1913 (N_1913,N_36,N_1510);
nand U1914 (N_1914,N_734,In_2003);
xnor U1915 (N_1915,In_2336,N_1364);
and U1916 (N_1916,N_1564,N_555);
or U1917 (N_1917,In_1641,N_1574);
nand U1918 (N_1918,N_1324,N_1020);
or U1919 (N_1919,N_97,N_1384);
nand U1920 (N_1920,N_1789,N_1616);
nor U1921 (N_1921,N_861,N_757);
or U1922 (N_1922,N_1326,N_1157);
xnor U1923 (N_1923,N_1650,In_520);
nor U1924 (N_1924,N_1335,In_2126);
xnor U1925 (N_1925,N_1386,N_650);
xor U1926 (N_1926,N_1443,N_1223);
xor U1927 (N_1927,In_2247,N_1516);
or U1928 (N_1928,N_703,N_846);
xor U1929 (N_1929,N_404,N_1460);
xnor U1930 (N_1930,N_1358,In_2610);
or U1931 (N_1931,N_508,In_393);
or U1932 (N_1932,N_1538,In_67);
nor U1933 (N_1933,In_1214,N_645);
and U1934 (N_1934,In_254,N_1679);
or U1935 (N_1935,In_1188,In_2952);
nand U1936 (N_1936,N_1195,N_1319);
nor U1937 (N_1937,N_926,N_1413);
nor U1938 (N_1938,N_1672,N_1625);
nor U1939 (N_1939,N_140,N_1313);
nand U1940 (N_1940,In_1207,N_1405);
or U1941 (N_1941,In_1132,N_1258);
nor U1942 (N_1942,In_454,N_459);
nand U1943 (N_1943,N_570,N_1607);
nor U1944 (N_1944,N_976,N_337);
xnor U1945 (N_1945,N_760,N_1623);
or U1946 (N_1946,N_568,N_1222);
nor U1947 (N_1947,N_1480,In_45);
or U1948 (N_1948,In_1015,N_1747);
and U1949 (N_1949,In_2936,N_700);
nand U1950 (N_1950,N_230,In_1977);
and U1951 (N_1951,In_2879,In_465);
nand U1952 (N_1952,In_2353,N_1640);
and U1953 (N_1953,N_1472,In_2432);
nand U1954 (N_1954,In_212,N_620);
nand U1955 (N_1955,N_1416,N_731);
or U1956 (N_1956,N_1406,N_1323);
xor U1957 (N_1957,N_1025,N_197);
nand U1958 (N_1958,In_2613,N_1566);
nand U1959 (N_1959,N_624,In_2103);
xor U1960 (N_1960,N_334,N_1303);
nand U1961 (N_1961,N_1787,N_1749);
nand U1962 (N_1962,N_847,N_1725);
and U1963 (N_1963,In_2289,In_1949);
nor U1964 (N_1964,In_2292,In_686);
xnor U1965 (N_1965,N_1683,N_942);
and U1966 (N_1966,In_938,N_738);
xnor U1967 (N_1967,N_1700,N_1398);
nand U1968 (N_1968,N_1199,In_2658);
nand U1969 (N_1969,N_170,In_708);
nor U1970 (N_1970,N_745,In_2229);
or U1971 (N_1971,In_631,N_1244);
or U1972 (N_1972,N_1644,N_277);
nand U1973 (N_1973,N_1748,N_304);
nand U1974 (N_1974,N_75,N_1415);
and U1975 (N_1975,N_1430,N_706);
xnor U1976 (N_1976,N_1030,In_2493);
nor U1977 (N_1977,In_1105,N_1631);
or U1978 (N_1978,N_1028,In_1128);
xnor U1979 (N_1979,N_856,N_1404);
xnor U1980 (N_1980,In_94,N_1620);
nand U1981 (N_1981,N_1708,N_503);
or U1982 (N_1982,In_2080,N_26);
and U1983 (N_1983,In_2847,N_370);
nor U1984 (N_1984,In_1122,N_1387);
nor U1985 (N_1985,N_1466,In_2302);
nor U1986 (N_1986,In_2205,N_1668);
or U1987 (N_1987,In_2915,N_1339);
and U1988 (N_1988,N_1207,N_1409);
and U1989 (N_1989,N_1221,N_1702);
nor U1990 (N_1990,N_1362,N_813);
or U1991 (N_1991,N_1262,N_1534);
and U1992 (N_1992,In_1680,N_1307);
xnor U1993 (N_1993,In_2574,In_1859);
nor U1994 (N_1994,N_825,N_784);
or U1995 (N_1995,N_744,N_1414);
or U1996 (N_1996,In_2954,N_1598);
xnor U1997 (N_1997,N_1318,N_1124);
nand U1998 (N_1998,N_1057,N_1290);
nor U1999 (N_1999,In_261,N_1704);
or U2000 (N_2000,N_1344,N_1491);
or U2001 (N_2001,N_1767,N_1462);
or U2002 (N_2002,In_1918,In_1974);
and U2003 (N_2003,N_299,N_267);
and U2004 (N_2004,In_181,N_436);
and U2005 (N_2005,N_1743,N_1523);
and U2006 (N_2006,N_1274,N_1357);
nor U2007 (N_2007,N_1772,N_1311);
nand U2008 (N_2008,In_2413,N_603);
nor U2009 (N_2009,In_2665,N_770);
and U2010 (N_2010,N_1287,N_1288);
nand U2011 (N_2011,N_1556,N_1417);
or U2012 (N_2012,N_1795,N_1669);
or U2013 (N_2013,N_1382,In_2958);
nand U2014 (N_2014,N_446,In_37);
and U2015 (N_2015,N_1680,In_481);
nor U2016 (N_2016,N_1503,N_1755);
or U2017 (N_2017,N_1084,N_1375);
or U2018 (N_2018,N_1515,N_1654);
or U2019 (N_2019,In_1673,N_1233);
nor U2020 (N_2020,N_1432,N_1054);
nand U2021 (N_2021,In_579,In_505);
xor U2022 (N_2022,N_1563,N_1773);
or U2023 (N_2023,In_2481,N_614);
nand U2024 (N_2024,N_1507,N_1706);
or U2025 (N_2025,N_1309,N_1611);
or U2026 (N_2026,N_1483,In_2565);
and U2027 (N_2027,N_1511,N_1388);
or U2028 (N_2028,In_1293,N_1697);
xor U2029 (N_2029,N_1302,In_1799);
nand U2030 (N_2030,N_1427,N_1717);
nor U2031 (N_2031,N_1780,N_1225);
nor U2032 (N_2032,N_1454,N_543);
nand U2033 (N_2033,N_1418,N_1627);
nand U2034 (N_2034,N_992,N_1651);
nand U2035 (N_2035,N_16,N_1269);
xor U2036 (N_2036,N_1502,N_1438);
and U2037 (N_2037,N_1238,N_1731);
nor U2038 (N_2038,N_1245,N_62);
nor U2039 (N_2039,N_1732,In_1708);
nand U2040 (N_2040,In_1647,N_623);
xnor U2041 (N_2041,N_1071,N_1272);
and U2042 (N_2042,N_1037,N_281);
nand U2043 (N_2043,N_1628,In_613);
nand U2044 (N_2044,N_1530,N_1692);
nor U2045 (N_2045,N_55,N_1144);
nand U2046 (N_2046,N_1251,In_2964);
nor U2047 (N_2047,N_1421,N_1770);
or U2048 (N_2048,N_283,N_525);
and U2049 (N_2049,N_1517,N_1434);
or U2050 (N_2050,In_123,In_2799);
nand U2051 (N_2051,N_1444,N_1040);
or U2052 (N_2052,N_1765,In_2234);
and U2053 (N_2053,N_1746,In_2687);
nand U2054 (N_2054,In_1173,In_213);
nor U2055 (N_2055,N_1108,N_183);
and U2056 (N_2056,N_1014,N_836);
or U2057 (N_2057,N_1265,N_1422);
nand U2058 (N_2058,N_1508,N_687);
and U2059 (N_2059,In_419,N_1475);
nor U2060 (N_2060,N_271,In_738);
nand U2061 (N_2061,In_298,In_1753);
or U2062 (N_2062,N_1445,N_1715);
and U2063 (N_2063,In_2271,N_1588);
or U2064 (N_2064,In_637,N_1257);
nand U2065 (N_2065,N_1471,N_1286);
xor U2066 (N_2066,In_511,N_1689);
and U2067 (N_2067,N_1359,In_1852);
or U2068 (N_2068,N_1658,N_233);
or U2069 (N_2069,N_1355,N_1228);
xor U2070 (N_2070,N_1297,N_1645);
nand U2071 (N_2071,N_639,In_2779);
nand U2072 (N_2072,N_1280,N_1401);
xor U2073 (N_2073,N_1741,N_1778);
xor U2074 (N_2074,N_1312,N_342);
or U2075 (N_2075,N_327,N_1726);
and U2076 (N_2076,N_1059,N_1684);
nand U2077 (N_2077,In_1001,N_318);
nor U2078 (N_2078,N_943,N_1547);
nand U2079 (N_2079,In_1171,N_1306);
nor U2080 (N_2080,N_969,In_2552);
nand U2081 (N_2081,N_1493,N_586);
xnor U2082 (N_2082,N_887,N_1284);
nand U2083 (N_2083,N_1622,N_644);
xor U2084 (N_2084,N_1490,N_1639);
or U2085 (N_2085,N_1782,N_1407);
or U2086 (N_2086,N_984,N_1484);
nor U2087 (N_2087,N_1268,N_1605);
and U2088 (N_2088,N_1321,In_1176);
and U2089 (N_2089,In_978,In_1078);
nand U2090 (N_2090,In_2226,N_1600);
or U2091 (N_2091,In_1627,In_1378);
xor U2092 (N_2092,N_1348,N_1448);
and U2093 (N_2093,In_2701,N_1520);
and U2094 (N_2094,N_1281,N_1580);
or U2095 (N_2095,In_1755,In_2227);
nand U2096 (N_2096,In_2890,N_1399);
or U2097 (N_2097,N_1066,N_1205);
nor U2098 (N_2098,N_1209,N_1264);
xnor U2099 (N_2099,N_962,N_863);
and U2100 (N_2100,N_1352,N_1082);
xnor U2101 (N_2101,N_1379,In_797);
nor U2102 (N_2102,In_1643,N_1643);
and U2103 (N_2103,N_755,In_1435);
nand U2104 (N_2104,N_1032,N_1609);
and U2105 (N_2105,In_2899,N_1449);
nand U2106 (N_2106,N_1250,In_390);
nor U2107 (N_2107,N_1792,N_1587);
or U2108 (N_2108,N_1714,N_735);
or U2109 (N_2109,In_1940,N_1456);
and U2110 (N_2110,N_1701,N_1426);
nand U2111 (N_2111,N_1316,In_2694);
nor U2112 (N_2112,N_1322,N_1377);
and U2113 (N_2113,N_1637,N_1486);
and U2114 (N_2114,In_2072,N_1576);
nor U2115 (N_2115,N_1351,N_1752);
nor U2116 (N_2116,N_1742,N_1068);
nand U2117 (N_2117,In_971,N_1383);
or U2118 (N_2118,N_1366,N_1695);
or U2119 (N_2119,N_1562,In_1080);
xor U2120 (N_2120,N_1513,N_1514);
nand U2121 (N_2121,N_1730,N_1594);
and U2122 (N_2122,In_1057,N_1389);
and U2123 (N_2123,N_1660,N_1604);
nor U2124 (N_2124,N_1247,N_1236);
xnor U2125 (N_2125,N_672,N_1285);
nand U2126 (N_2126,N_1561,N_1525);
nand U2127 (N_2127,In_1503,N_200);
and U2128 (N_2128,In_1218,N_313);
nand U2129 (N_2129,In_2043,N_1690);
xor U2130 (N_2130,In_1422,N_1603);
or U2131 (N_2131,In_2566,N_311);
nand U2132 (N_2132,N_651,N_1633);
nand U2133 (N_2133,N_1599,In_17);
xor U2134 (N_2134,In_904,N_1231);
xnor U2135 (N_2135,N_54,N_231);
or U2136 (N_2136,N_1391,N_1276);
nor U2137 (N_2137,N_1786,In_437);
nand U2138 (N_2138,N_1781,In_1644);
nor U2139 (N_2139,N_1261,In_1771);
nor U2140 (N_2140,In_176,In_232);
nand U2141 (N_2141,In_2909,N_1796);
nor U2142 (N_2142,N_1360,N_1338);
xor U2143 (N_2143,N_1206,N_1531);
xor U2144 (N_2144,N_1232,N_1655);
nand U2145 (N_2145,In_1897,In_1499);
xor U2146 (N_2146,N_1577,N_1649);
xor U2147 (N_2147,N_199,N_953);
or U2148 (N_2148,In_2361,N_1185);
and U2149 (N_2149,In_2198,N_1703);
or U2150 (N_2150,N_17,N_1278);
nand U2151 (N_2151,In_2206,In_1221);
xnor U2152 (N_2152,N_1431,N_165);
nor U2153 (N_2153,N_1300,N_1769);
xor U2154 (N_2154,N_1641,N_435);
nand U2155 (N_2155,In_1368,N_1473);
nand U2156 (N_2156,N_1667,In_934);
nor U2157 (N_2157,N_279,N_1602);
nand U2158 (N_2158,In_2221,In_458);
xor U2159 (N_2159,N_1396,In_182);
nor U2160 (N_2160,In_386,N_1589);
nand U2161 (N_2161,N_1393,N_1334);
nor U2162 (N_2162,N_1601,In_2329);
xor U2163 (N_2163,N_1527,N_1365);
nor U2164 (N_2164,In_874,N_1612);
or U2165 (N_2165,N_1340,N_1139);
xnor U2166 (N_2166,N_1686,N_1147);
nand U2167 (N_2167,N_1220,N_1737);
nor U2168 (N_2168,N_1126,N_1545);
or U2169 (N_2169,In_1228,In_1697);
and U2170 (N_2170,N_1402,N_1337);
and U2171 (N_2171,N_1012,In_2050);
xor U2172 (N_2172,N_1075,In_1812);
nand U2173 (N_2173,In_2519,N_542);
xor U2174 (N_2174,N_1477,N_1341);
nor U2175 (N_2175,N_1143,In_1964);
nand U2176 (N_2176,In_2853,N_803);
xnor U2177 (N_2177,N_1734,N_1227);
nor U2178 (N_2178,N_1279,N_736);
and U2179 (N_2179,N_1552,N_872);
nand U2180 (N_2180,In_266,N_138);
nand U2181 (N_2181,N_1400,N_42);
nor U2182 (N_2182,N_1370,N_1242);
and U2183 (N_2183,N_1635,N_773);
nand U2184 (N_2184,N_1273,N_1001);
xnor U2185 (N_2185,In_1412,In_626);
and U2186 (N_2186,N_1648,In_763);
and U2187 (N_2187,N_1465,N_609);
or U2188 (N_2188,N_1481,In_687);
and U2189 (N_2189,N_711,In_1843);
or U2190 (N_2190,In_1513,In_2718);
and U2191 (N_2191,N_918,N_1027);
nor U2192 (N_2192,N_1590,N_368);
nand U2193 (N_2193,In_2400,N_1595);
xor U2194 (N_2194,N_1489,In_1425);
or U2195 (N_2195,N_692,In_1163);
nor U2196 (N_2196,N_563,In_1209);
xnor U2197 (N_2197,N_1575,N_1739);
xnor U2198 (N_2198,In_1632,N_1626);
or U2199 (N_2199,In_2156,In_412);
nor U2200 (N_2200,N_1736,N_1634);
or U2201 (N_2201,N_787,N_1759);
or U2202 (N_2202,N_1457,N_174);
nand U2203 (N_2203,N_369,In_2146);
nor U2204 (N_2204,N_1293,N_1216);
or U2205 (N_2205,In_257,In_1198);
nand U2206 (N_2206,N_1524,N_1254);
nor U2207 (N_2207,In_984,N_1046);
or U2208 (N_2208,In_1661,N_1436);
xnor U2209 (N_2209,N_1439,N_1350);
nor U2210 (N_2210,N_667,N_40);
or U2211 (N_2211,N_1674,In_944);
and U2212 (N_2212,N_1533,N_1239);
xor U2213 (N_2213,N_1677,N_1621);
or U2214 (N_2214,N_1428,N_1768);
xnor U2215 (N_2215,In_1215,In_1269);
and U2216 (N_2216,N_657,N_681);
xor U2217 (N_2217,In_2035,N_922);
xor U2218 (N_2218,N_613,N_1294);
nand U2219 (N_2219,In_1862,In_2446);
or U2220 (N_2220,N_1671,In_2257);
nand U2221 (N_2221,In_2878,N_1346);
and U2222 (N_2222,In_1531,N_1259);
or U2223 (N_2223,In_2938,N_1691);
or U2224 (N_2224,N_479,N_709);
and U2225 (N_2225,In_2425,In_2618);
or U2226 (N_2226,N_1557,N_1532);
xnor U2227 (N_2227,N_1447,N_1617);
nor U2228 (N_2228,N_699,N_1369);
nand U2229 (N_2229,In_1611,N_1275);
and U2230 (N_2230,In_1919,N_70);
xnor U2231 (N_2231,N_1670,N_864);
or U2232 (N_2232,N_1343,N_1573);
xnor U2233 (N_2233,N_689,In_2125);
nor U2234 (N_2234,In_1154,N_76);
and U2235 (N_2235,N_1681,In_179);
nand U2236 (N_2236,In_1429,N_1419);
nand U2237 (N_2237,N_1342,N_1423);
nand U2238 (N_2238,N_1710,N_789);
or U2239 (N_2239,In_1937,N_722);
xnor U2240 (N_2240,N_1214,In_1526);
nor U2241 (N_2241,N_987,N_1308);
nand U2242 (N_2242,In_65,In_669);
nand U2243 (N_2243,N_1512,N_1240);
or U2244 (N_2244,N_1329,N_1745);
or U2245 (N_2245,N_475,N_1353);
or U2246 (N_2246,N_359,N_1793);
nand U2247 (N_2247,N_1373,N_1662);
or U2248 (N_2248,In_2098,N_1151);
nand U2249 (N_2249,In_1963,N_554);
xnor U2250 (N_2250,In_332,N_1760);
nor U2251 (N_2251,N_1544,N_83);
or U2252 (N_2252,N_1390,N_1361);
or U2253 (N_2253,N_1581,N_1653);
and U2254 (N_2254,In_58,N_1753);
nand U2255 (N_2255,N_1756,N_1217);
and U2256 (N_2256,N_714,N_1539);
or U2257 (N_2257,N_859,In_2322);
nor U2258 (N_2258,In_2024,N_1606);
xnor U2259 (N_2259,N_1546,In_1916);
and U2260 (N_2260,N_1608,N_1550);
nor U2261 (N_2261,In_2778,N_562);
and U2262 (N_2262,In_1035,In_51);
or U2263 (N_2263,N_1729,N_1256);
and U2264 (N_2264,N_1559,N_1615);
nand U2265 (N_2265,N_1208,In_1800);
nand U2266 (N_2266,N_1420,N_1764);
nand U2267 (N_2267,N_1636,N_1141);
nor U2268 (N_2268,N_1560,N_1079);
or U2269 (N_2269,N_1429,In_903);
nor U2270 (N_2270,N_1646,N_1210);
nor U2271 (N_2271,N_1713,N_285);
and U2272 (N_2272,In_2547,N_1197);
nor U2273 (N_2273,N_951,N_1784);
nand U2274 (N_2274,N_1397,In_1041);
xnor U2275 (N_2275,In_2619,N_1762);
xor U2276 (N_2276,N_1011,N_154);
nor U2277 (N_2277,In_1296,N_970);
nand U2278 (N_2278,N_1320,N_1495);
nor U2279 (N_2279,N_656,N_1665);
nand U2280 (N_2280,N_1201,N_1497);
nor U2281 (N_2281,N_423,In_724);
nor U2282 (N_2282,In_265,N_691);
and U2283 (N_2283,N_1371,N_1705);
and U2284 (N_2284,N_494,N_114);
nor U2285 (N_2285,In_894,N_173);
nor U2286 (N_2286,N_1298,In_442);
nand U2287 (N_2287,N_594,N_1629);
nor U2288 (N_2288,N_1299,N_1504);
nand U2289 (N_2289,In_2081,N_1461);
nand U2290 (N_2290,N_175,N_1788);
nand U2291 (N_2291,In_587,N_1500);
xor U2292 (N_2292,N_585,In_865);
xnor U2293 (N_2293,N_229,In_2133);
and U2294 (N_2294,In_1211,In_1712);
xor U2295 (N_2295,In_1874,In_2078);
and U2296 (N_2296,In_1969,N_1327);
nand U2297 (N_2297,In_946,N_1229);
and U2298 (N_2298,N_1696,N_1328);
nand U2299 (N_2299,N_1693,In_1564);
nor U2300 (N_2300,N_330,In_112);
and U2301 (N_2301,N_1378,N_1356);
and U2302 (N_2302,N_794,In_358);
or U2303 (N_2303,N_1459,N_1536);
or U2304 (N_2304,N_898,N_1235);
nor U2305 (N_2305,N_1776,N_1785);
xor U2306 (N_2306,In_1261,In_2689);
nor U2307 (N_2307,N_1505,N_1496);
or U2308 (N_2308,N_1234,N_713);
or U2309 (N_2309,In_1790,N_1548);
xor U2310 (N_2310,N_1652,N_1541);
xor U2311 (N_2311,N_1619,N_222);
nor U2312 (N_2312,N_608,N_1592);
nand U2313 (N_2313,In_1593,N_77);
or U2314 (N_2314,In_846,In_1610);
or U2315 (N_2315,N_1551,N_1292);
xnor U2316 (N_2316,In_2951,N_1363);
and U2317 (N_2317,N_1642,N_211);
nor U2318 (N_2318,In_2364,N_1345);
and U2319 (N_2319,N_1253,N_1727);
nor U2320 (N_2320,N_1412,N_772);
nand U2321 (N_2321,In_1389,In_1230);
nand U2322 (N_2322,N_1034,N_1799);
nor U2323 (N_2323,N_43,N_1347);
or U2324 (N_2324,N_1403,N_1376);
nand U2325 (N_2325,N_1578,N_1464);
xnor U2326 (N_2326,N_1094,In_757);
or U2327 (N_2327,In_1695,N_812);
nand U2328 (N_2328,N_1521,In_4);
xor U2329 (N_2329,In_2715,In_732);
or U2330 (N_2330,N_1519,In_1692);
nand U2331 (N_2331,In_2150,N_779);
nor U2332 (N_2332,N_1757,N_1080);
xor U2333 (N_2333,N_44,In_2883);
nor U2334 (N_2334,N_1663,In_1250);
or U2335 (N_2335,N_1777,N_1433);
or U2336 (N_2336,N_1659,N_1783);
nand U2337 (N_2337,N_1721,In_1279);
xor U2338 (N_2338,N_871,N_1766);
nand U2339 (N_2339,N_1441,N_1271);
xor U2340 (N_2340,N_1090,N_1203);
nor U2341 (N_2341,N_688,N_1230);
and U2342 (N_2342,N_1656,N_1526);
and U2343 (N_2343,N_1061,N_1492);
xor U2344 (N_2344,N_1463,N_1470);
nand U2345 (N_2345,In_1685,N_1394);
nor U2346 (N_2346,N_1638,In_355);
nand U2347 (N_2347,In_1734,N_1478);
nand U2348 (N_2348,N_1474,N_1277);
nand U2349 (N_2349,N_372,N_1798);
nand U2350 (N_2350,N_1354,N_1618);
nand U2351 (N_2351,In_838,N_1446);
nand U2352 (N_2352,N_1479,N_1301);
nand U2353 (N_2353,In_1062,In_912);
nand U2354 (N_2354,N_1248,In_1829);
xor U2355 (N_2355,In_223,N_1263);
nand U2356 (N_2356,N_1582,N_1675);
nor U2357 (N_2357,N_1583,In_556);
nor U2358 (N_2358,In_2261,N_1270);
and U2359 (N_2359,In_1432,In_974);
and U2360 (N_2360,In_1844,N_1719);
nor U2361 (N_2361,N_1440,N_1676);
or U2362 (N_2362,In_2624,N_1142);
nand U2363 (N_2363,In_653,N_1266);
nor U2364 (N_2364,In_2607,In_2549);
xor U2365 (N_2365,N_34,N_1381);
or U2366 (N_2366,In_2982,N_1291);
nor U2367 (N_2367,N_1224,N_1549);
or U2368 (N_2368,In_791,In_531);
nand U2369 (N_2369,N_1452,N_1237);
or U2370 (N_2370,N_1295,N_973);
and U2371 (N_2371,N_670,N_1724);
nor U2372 (N_2372,N_1494,N_349);
and U2373 (N_2373,N_1614,N_1076);
nor U2374 (N_2374,In_688,N_1073);
xnor U2375 (N_2375,N_1537,In_840);
and U2376 (N_2376,N_1797,N_1024);
and U2377 (N_2377,N_1049,In_1101);
xnor U2378 (N_2378,In_2534,N_1482);
nand U2379 (N_2379,N_1260,N_1707);
xnor U2380 (N_2380,N_785,In_860);
xnor U2381 (N_2381,N_1593,N_707);
or U2382 (N_2382,In_2719,N_354);
nor U2383 (N_2383,N_1453,In_344);
nand U2384 (N_2384,N_1694,In_2489);
nand U2385 (N_2385,In_670,N_1215);
nand U2386 (N_2386,N_156,In_1795);
and U2387 (N_2387,In_289,In_1116);
nand U2388 (N_2388,N_618,N_1791);
and U2389 (N_2389,N_151,N_1296);
xnor U2390 (N_2390,In_2047,In_349);
nand U2391 (N_2391,N_1018,N_1213);
xor U2392 (N_2392,N_393,N_1750);
nor U2393 (N_2393,N_739,N_1664);
or U2394 (N_2394,N_1499,N_791);
nand U2395 (N_2395,N_694,N_1305);
or U2396 (N_2396,N_530,N_1081);
nor U2397 (N_2397,N_205,In_2367);
or U2398 (N_2398,N_1771,In_2888);
nor U2399 (N_2399,N_1218,N_1728);
or U2400 (N_2400,N_2135,N_2377);
xor U2401 (N_2401,N_2257,N_2362);
xor U2402 (N_2402,N_2154,N_1872);
xor U2403 (N_2403,N_1990,N_2124);
and U2404 (N_2404,N_1869,N_2172);
xnor U2405 (N_2405,N_2203,N_2357);
xnor U2406 (N_2406,N_2146,N_2041);
nor U2407 (N_2407,N_2138,N_1934);
xor U2408 (N_2408,N_1976,N_2390);
or U2409 (N_2409,N_1857,N_2057);
or U2410 (N_2410,N_2184,N_2081);
or U2411 (N_2411,N_2358,N_2060);
or U2412 (N_2412,N_1807,N_2248);
and U2413 (N_2413,N_1911,N_1948);
xor U2414 (N_2414,N_2311,N_1979);
nand U2415 (N_2415,N_1825,N_1989);
xor U2416 (N_2416,N_1973,N_2005);
nor U2417 (N_2417,N_2361,N_2394);
nor U2418 (N_2418,N_1884,N_2087);
nor U2419 (N_2419,N_2205,N_2235);
nor U2420 (N_2420,N_1986,N_2156);
xnor U2421 (N_2421,N_2094,N_2313);
or U2422 (N_2422,N_2148,N_2340);
nor U2423 (N_2423,N_1977,N_2030);
or U2424 (N_2424,N_2356,N_2147);
nor U2425 (N_2425,N_1945,N_2003);
xnor U2426 (N_2426,N_1891,N_2028);
nand U2427 (N_2427,N_1912,N_2145);
and U2428 (N_2428,N_2105,N_2023);
or U2429 (N_2429,N_2158,N_1864);
and U2430 (N_2430,N_2083,N_2284);
nand U2431 (N_2431,N_1974,N_1941);
or U2432 (N_2432,N_1987,N_1936);
and U2433 (N_2433,N_1992,N_2366);
nand U2434 (N_2434,N_1985,N_1889);
and U2435 (N_2435,N_2033,N_1914);
nor U2436 (N_2436,N_2183,N_1802);
nand U2437 (N_2437,N_2007,N_2050);
or U2438 (N_2438,N_2144,N_2364);
nand U2439 (N_2439,N_1877,N_1822);
nand U2440 (N_2440,N_2399,N_2268);
nor U2441 (N_2441,N_1996,N_2042);
nor U2442 (N_2442,N_2293,N_2290);
nor U2443 (N_2443,N_2233,N_1844);
and U2444 (N_2444,N_2212,N_2220);
and U2445 (N_2445,N_2376,N_2382);
xor U2446 (N_2446,N_1960,N_2192);
and U2447 (N_2447,N_2274,N_2179);
or U2448 (N_2448,N_2185,N_2052);
nor U2449 (N_2449,N_2092,N_2231);
xor U2450 (N_2450,N_2244,N_1896);
and U2451 (N_2451,N_2353,N_2236);
xnor U2452 (N_2452,N_2080,N_2275);
xor U2453 (N_2453,N_2160,N_1865);
nand U2454 (N_2454,N_1937,N_2139);
and U2455 (N_2455,N_1858,N_1981);
nand U2456 (N_2456,N_2072,N_2064);
nand U2457 (N_2457,N_2354,N_2044);
xnor U2458 (N_2458,N_1863,N_2393);
nor U2459 (N_2459,N_1827,N_2054);
nor U2460 (N_2460,N_1931,N_2206);
nor U2461 (N_2461,N_2073,N_2200);
and U2462 (N_2462,N_1829,N_2306);
or U2463 (N_2463,N_2239,N_2024);
xor U2464 (N_2464,N_2318,N_2036);
nand U2465 (N_2465,N_2258,N_2225);
and U2466 (N_2466,N_1812,N_2343);
and U2467 (N_2467,N_2097,N_1951);
nand U2468 (N_2468,N_1814,N_2093);
nor U2469 (N_2469,N_2101,N_2168);
xnor U2470 (N_2470,N_2304,N_1839);
nor U2471 (N_2471,N_2240,N_2398);
xnor U2472 (N_2472,N_2285,N_2312);
xor U2473 (N_2473,N_2375,N_2056);
xnor U2474 (N_2474,N_1878,N_2230);
xnor U2475 (N_2475,N_2221,N_1848);
and U2476 (N_2476,N_1800,N_2281);
xor U2477 (N_2477,N_2171,N_2242);
xor U2478 (N_2478,N_1843,N_2095);
or U2479 (N_2479,N_2130,N_2226);
nor U2480 (N_2480,N_2025,N_1984);
or U2481 (N_2481,N_2189,N_1925);
nand U2482 (N_2482,N_2218,N_2341);
nand U2483 (N_2483,N_2166,N_2043);
or U2484 (N_2484,N_1815,N_2392);
nor U2485 (N_2485,N_2209,N_1866);
or U2486 (N_2486,N_2061,N_2234);
or U2487 (N_2487,N_1859,N_2053);
xor U2488 (N_2488,N_2252,N_1835);
or U2489 (N_2489,N_2085,N_2336);
and U2490 (N_2490,N_1817,N_1983);
or U2491 (N_2491,N_2090,N_2322);
and U2492 (N_2492,N_2176,N_2165);
nor U2493 (N_2493,N_1968,N_1840);
xnor U2494 (N_2494,N_2187,N_2114);
nand U2495 (N_2495,N_2211,N_2029);
or U2496 (N_2496,N_2153,N_2283);
xnor U2497 (N_2497,N_2262,N_2355);
xnor U2498 (N_2498,N_2074,N_2068);
nor U2499 (N_2499,N_1972,N_2088);
nor U2500 (N_2500,N_2141,N_1927);
xnor U2501 (N_2501,N_2196,N_2113);
or U2502 (N_2502,N_1901,N_2055);
or U2503 (N_2503,N_2129,N_1944);
nand U2504 (N_2504,N_1861,N_2288);
xor U2505 (N_2505,N_2178,N_2110);
or U2506 (N_2506,N_2250,N_1966);
nand U2507 (N_2507,N_2243,N_2259);
xnor U2508 (N_2508,N_1924,N_2107);
nor U2509 (N_2509,N_1913,N_2380);
or U2510 (N_2510,N_2267,N_2102);
and U2511 (N_2511,N_1804,N_1921);
xor U2512 (N_2512,N_2224,N_2098);
nand U2513 (N_2513,N_2278,N_2201);
xor U2514 (N_2514,N_2182,N_2315);
xnor U2515 (N_2515,N_1862,N_1849);
xnor U2516 (N_2516,N_2122,N_2365);
nand U2517 (N_2517,N_1953,N_2379);
nor U2518 (N_2518,N_1845,N_2237);
nand U2519 (N_2519,N_2344,N_1930);
nor U2520 (N_2520,N_2269,N_2077);
xnor U2521 (N_2521,N_1995,N_2381);
nor U2522 (N_2522,N_1853,N_1906);
xor U2523 (N_2523,N_2350,N_2142);
xnor U2524 (N_2524,N_2294,N_1892);
nand U2525 (N_2525,N_2296,N_2099);
xor U2526 (N_2526,N_1824,N_2149);
and U2527 (N_2527,N_1918,N_2317);
nand U2528 (N_2528,N_1886,N_2299);
nand U2529 (N_2529,N_1935,N_2161);
nor U2530 (N_2530,N_2018,N_2048);
xor U2531 (N_2531,N_2216,N_2133);
nand U2532 (N_2532,N_2261,N_1870);
nand U2533 (N_2533,N_2348,N_1938);
xnor U2534 (N_2534,N_2307,N_2316);
nor U2535 (N_2535,N_2324,N_2222);
nor U2536 (N_2536,N_2150,N_1883);
nor U2537 (N_2537,N_2363,N_2241);
or U2538 (N_2538,N_1905,N_2279);
or U2539 (N_2539,N_2163,N_2143);
xor U2540 (N_2540,N_1855,N_2082);
and U2541 (N_2541,N_2345,N_2389);
xnor U2542 (N_2542,N_2188,N_2021);
xnor U2543 (N_2543,N_2228,N_2089);
nor U2544 (N_2544,N_2347,N_2039);
nand U2545 (N_2545,N_1932,N_2351);
and U2546 (N_2546,N_2310,N_2181);
nand U2547 (N_2547,N_2256,N_2286);
and U2548 (N_2548,N_2199,N_2067);
and U2549 (N_2549,N_1809,N_2013);
or U2550 (N_2550,N_2374,N_2096);
or U2551 (N_2551,N_2004,N_2246);
nor U2552 (N_2552,N_1919,N_1908);
xor U2553 (N_2553,N_1888,N_1868);
or U2554 (N_2554,N_2391,N_2397);
or U2555 (N_2555,N_1916,N_2372);
nand U2556 (N_2556,N_1895,N_2308);
nor U2557 (N_2557,N_2155,N_2177);
xor U2558 (N_2558,N_2022,N_2157);
or U2559 (N_2559,N_1851,N_2121);
and U2560 (N_2560,N_2169,N_2352);
nor U2561 (N_2561,N_1920,N_2108);
nand U2562 (N_2562,N_2245,N_1873);
or U2563 (N_2563,N_2213,N_2297);
xnor U2564 (N_2564,N_2333,N_2383);
nor U2565 (N_2565,N_2338,N_2035);
nor U2566 (N_2566,N_1942,N_2008);
and U2567 (N_2567,N_2175,N_2232);
xor U2568 (N_2568,N_2070,N_2049);
nand U2569 (N_2569,N_2038,N_2238);
xor U2570 (N_2570,N_1893,N_2280);
nand U2571 (N_2571,N_2368,N_1867);
nor U2572 (N_2572,N_1847,N_1929);
xor U2573 (N_2573,N_1952,N_2076);
nor U2574 (N_2574,N_1980,N_2020);
and U2575 (N_2575,N_1907,N_2197);
xor U2576 (N_2576,N_2395,N_2136);
xnor U2577 (N_2577,N_2264,N_2137);
and U2578 (N_2578,N_1988,N_1818);
and U2579 (N_2579,N_1882,N_2219);
xnor U2580 (N_2580,N_2120,N_1900);
nand U2581 (N_2581,N_2173,N_1963);
xor U2582 (N_2582,N_1958,N_2058);
and U2583 (N_2583,N_1915,N_1975);
or U2584 (N_2584,N_2190,N_2075);
and U2585 (N_2585,N_1969,N_2263);
or U2586 (N_2586,N_1805,N_1830);
nand U2587 (N_2587,N_2032,N_1831);
nand U2588 (N_2588,N_2112,N_1894);
and U2589 (N_2589,N_2115,N_1806);
xnor U2590 (N_2590,N_2151,N_1950);
and U2591 (N_2591,N_2385,N_2370);
and U2592 (N_2592,N_1993,N_1903);
nor U2593 (N_2593,N_1978,N_2046);
nand U2594 (N_2594,N_1955,N_2027);
or U2595 (N_2595,N_2100,N_1994);
and U2596 (N_2596,N_2387,N_1956);
nor U2597 (N_2597,N_1991,N_2051);
nand U2598 (N_2598,N_2273,N_1816);
xor U2599 (N_2599,N_1833,N_2071);
nor U2600 (N_2600,N_2369,N_2339);
and U2601 (N_2601,N_2065,N_2016);
nor U2602 (N_2602,N_1917,N_2040);
xor U2603 (N_2603,N_2132,N_2265);
xor U2604 (N_2604,N_1887,N_1954);
nand U2605 (N_2605,N_2078,N_2012);
nand U2606 (N_2606,N_2330,N_1998);
nor U2607 (N_2607,N_2002,N_1828);
nor U2608 (N_2608,N_2371,N_2084);
nor U2609 (N_2609,N_2047,N_2069);
xnor U2610 (N_2610,N_2174,N_1964);
and U2611 (N_2611,N_2342,N_2117);
or U2612 (N_2612,N_2277,N_1836);
nand U2613 (N_2613,N_2298,N_2207);
or U2614 (N_2614,N_2119,N_1957);
or U2615 (N_2615,N_1841,N_1810);
xor U2616 (N_2616,N_2170,N_2208);
nand U2617 (N_2617,N_2282,N_2255);
nand U2618 (N_2618,N_2159,N_2204);
and U2619 (N_2619,N_2272,N_1881);
xnor U2620 (N_2620,N_1962,N_2009);
or U2621 (N_2621,N_1943,N_1926);
xnor U2622 (N_2622,N_1904,N_2326);
or U2623 (N_2623,N_2227,N_2223);
nand U2624 (N_2624,N_2271,N_1850);
nor U2625 (N_2625,N_2396,N_2254);
nand U2626 (N_2626,N_1997,N_2063);
and U2627 (N_2627,N_1837,N_2289);
xnor U2628 (N_2628,N_2001,N_1880);
xor U2629 (N_2629,N_2331,N_2266);
xnor U2630 (N_2630,N_2193,N_1821);
xor U2631 (N_2631,N_2152,N_2309);
xor U2632 (N_2632,N_1879,N_1928);
nand U2633 (N_2633,N_2125,N_1939);
and U2634 (N_2634,N_2328,N_2037);
or U2635 (N_2635,N_2337,N_1910);
and U2636 (N_2636,N_2386,N_2126);
nand U2637 (N_2637,N_2010,N_2059);
xnor U2638 (N_2638,N_2118,N_2349);
nand U2639 (N_2639,N_2378,N_1823);
or U2640 (N_2640,N_2217,N_2162);
xnor U2641 (N_2641,N_2314,N_2359);
nor U2642 (N_2642,N_1860,N_2388);
xor U2643 (N_2643,N_2079,N_2164);
xor U2644 (N_2644,N_2017,N_2167);
and U2645 (N_2645,N_1965,N_2031);
and U2646 (N_2646,N_2123,N_2111);
nand U2647 (N_2647,N_1961,N_2015);
xnor U2648 (N_2648,N_1826,N_2116);
and U2649 (N_2649,N_2332,N_2325);
nand U2650 (N_2650,N_1940,N_2360);
nand U2651 (N_2651,N_2215,N_2214);
xor U2652 (N_2652,N_1890,N_1967);
and U2653 (N_2653,N_2091,N_2346);
and U2654 (N_2654,N_2302,N_2253);
nand U2655 (N_2655,N_1856,N_2334);
or U2656 (N_2656,N_2109,N_2367);
nand U2657 (N_2657,N_2045,N_2327);
and U2658 (N_2658,N_1838,N_1834);
and U2659 (N_2659,N_2249,N_2291);
or U2660 (N_2660,N_2198,N_1842);
nand U2661 (N_2661,N_1876,N_2180);
nor U2662 (N_2662,N_1803,N_2301);
nor U2663 (N_2663,N_2335,N_2384);
nand U2664 (N_2664,N_1946,N_2251);
xor U2665 (N_2665,N_1982,N_2006);
nor U2666 (N_2666,N_1902,N_2034);
nor U2667 (N_2667,N_2373,N_2270);
nor U2668 (N_2668,N_2323,N_2295);
or U2669 (N_2669,N_2103,N_1832);
and U2670 (N_2670,N_2191,N_2026);
nor U2671 (N_2671,N_1949,N_1874);
nor U2672 (N_2672,N_2066,N_2106);
xor U2673 (N_2673,N_1846,N_2140);
or U2674 (N_2674,N_2104,N_1875);
or U2675 (N_2675,N_2329,N_1852);
or U2676 (N_2676,N_2247,N_2303);
or U2677 (N_2677,N_2300,N_1959);
or U2678 (N_2678,N_1933,N_2229);
nor U2679 (N_2679,N_1923,N_2320);
nand U2680 (N_2680,N_1999,N_2202);
nand U2681 (N_2681,N_2014,N_1909);
nor U2682 (N_2682,N_2195,N_2210);
nor U2683 (N_2683,N_2186,N_1820);
nand U2684 (N_2684,N_2134,N_2128);
or U2685 (N_2685,N_2062,N_2305);
and U2686 (N_2686,N_2011,N_2131);
and U2687 (N_2687,N_2321,N_1970);
or U2688 (N_2688,N_1897,N_2000);
xnor U2689 (N_2689,N_1947,N_2127);
xor U2690 (N_2690,N_1854,N_2319);
xnor U2691 (N_2691,N_1813,N_2287);
or U2692 (N_2692,N_1801,N_1922);
and U2693 (N_2693,N_1871,N_2292);
xor U2694 (N_2694,N_1811,N_1971);
nand U2695 (N_2695,N_1808,N_1885);
xor U2696 (N_2696,N_2260,N_2194);
and U2697 (N_2697,N_2276,N_1898);
and U2698 (N_2698,N_1819,N_2019);
and U2699 (N_2699,N_1899,N_2086);
or U2700 (N_2700,N_2285,N_1908);
and U2701 (N_2701,N_1825,N_2084);
or U2702 (N_2702,N_2074,N_1965);
and U2703 (N_2703,N_1913,N_2212);
nand U2704 (N_2704,N_2115,N_2319);
nand U2705 (N_2705,N_2085,N_2090);
or U2706 (N_2706,N_2319,N_2157);
and U2707 (N_2707,N_2393,N_2148);
nor U2708 (N_2708,N_2324,N_2190);
nor U2709 (N_2709,N_2224,N_1944);
nor U2710 (N_2710,N_2278,N_1999);
or U2711 (N_2711,N_2038,N_2159);
and U2712 (N_2712,N_2099,N_2271);
nor U2713 (N_2713,N_2098,N_2339);
nor U2714 (N_2714,N_2053,N_2010);
and U2715 (N_2715,N_2209,N_2217);
nor U2716 (N_2716,N_2247,N_2040);
or U2717 (N_2717,N_1815,N_2151);
and U2718 (N_2718,N_1826,N_2043);
or U2719 (N_2719,N_1801,N_1880);
and U2720 (N_2720,N_2242,N_2212);
nand U2721 (N_2721,N_2120,N_2285);
xnor U2722 (N_2722,N_2317,N_1957);
nor U2723 (N_2723,N_1836,N_2328);
or U2724 (N_2724,N_1981,N_2387);
nor U2725 (N_2725,N_2143,N_2089);
and U2726 (N_2726,N_1868,N_2000);
and U2727 (N_2727,N_1882,N_2039);
and U2728 (N_2728,N_1860,N_1874);
xnor U2729 (N_2729,N_1900,N_2316);
or U2730 (N_2730,N_2377,N_2022);
xor U2731 (N_2731,N_1828,N_2299);
and U2732 (N_2732,N_2026,N_2229);
or U2733 (N_2733,N_2256,N_2325);
nor U2734 (N_2734,N_2224,N_1844);
nor U2735 (N_2735,N_1911,N_2167);
nor U2736 (N_2736,N_1940,N_2035);
nor U2737 (N_2737,N_2065,N_2041);
and U2738 (N_2738,N_2016,N_1884);
and U2739 (N_2739,N_2230,N_1931);
xor U2740 (N_2740,N_2297,N_1898);
nand U2741 (N_2741,N_1934,N_2164);
xor U2742 (N_2742,N_2169,N_1912);
nand U2743 (N_2743,N_2185,N_2038);
and U2744 (N_2744,N_2240,N_2018);
or U2745 (N_2745,N_1904,N_2199);
or U2746 (N_2746,N_2217,N_2089);
xor U2747 (N_2747,N_2392,N_1963);
or U2748 (N_2748,N_2080,N_2172);
nand U2749 (N_2749,N_1997,N_2334);
or U2750 (N_2750,N_2230,N_2232);
and U2751 (N_2751,N_2369,N_2308);
and U2752 (N_2752,N_1955,N_2022);
or U2753 (N_2753,N_2155,N_1946);
nand U2754 (N_2754,N_2271,N_2328);
or U2755 (N_2755,N_1950,N_2191);
and U2756 (N_2756,N_2089,N_2321);
nand U2757 (N_2757,N_2352,N_2063);
nor U2758 (N_2758,N_2150,N_2265);
nor U2759 (N_2759,N_2127,N_1923);
or U2760 (N_2760,N_1988,N_1887);
and U2761 (N_2761,N_2096,N_2253);
xor U2762 (N_2762,N_2098,N_2376);
nor U2763 (N_2763,N_2187,N_2354);
xor U2764 (N_2764,N_2189,N_2014);
xor U2765 (N_2765,N_2237,N_2360);
nor U2766 (N_2766,N_2202,N_2010);
xor U2767 (N_2767,N_2251,N_2084);
nor U2768 (N_2768,N_1870,N_2140);
nor U2769 (N_2769,N_2137,N_2281);
or U2770 (N_2770,N_1931,N_2287);
nor U2771 (N_2771,N_2194,N_1889);
or U2772 (N_2772,N_1905,N_2175);
xor U2773 (N_2773,N_1919,N_1849);
nand U2774 (N_2774,N_2291,N_2384);
xnor U2775 (N_2775,N_1959,N_1847);
nor U2776 (N_2776,N_1818,N_1951);
nand U2777 (N_2777,N_2367,N_1957);
and U2778 (N_2778,N_2165,N_2349);
nand U2779 (N_2779,N_2331,N_2272);
or U2780 (N_2780,N_2372,N_1955);
nor U2781 (N_2781,N_2093,N_1811);
and U2782 (N_2782,N_2059,N_1836);
nor U2783 (N_2783,N_2243,N_2167);
xor U2784 (N_2784,N_2333,N_1988);
nor U2785 (N_2785,N_2223,N_2045);
xor U2786 (N_2786,N_1811,N_2084);
xnor U2787 (N_2787,N_1948,N_1951);
or U2788 (N_2788,N_2194,N_1984);
nor U2789 (N_2789,N_1804,N_2221);
and U2790 (N_2790,N_2181,N_2273);
or U2791 (N_2791,N_1812,N_2239);
xor U2792 (N_2792,N_2325,N_2187);
nor U2793 (N_2793,N_1880,N_2233);
and U2794 (N_2794,N_1982,N_2362);
or U2795 (N_2795,N_2392,N_2209);
nand U2796 (N_2796,N_2138,N_2338);
nand U2797 (N_2797,N_2344,N_2114);
nor U2798 (N_2798,N_1804,N_2282);
xor U2799 (N_2799,N_1880,N_2275);
and U2800 (N_2800,N_2272,N_2233);
xnor U2801 (N_2801,N_2266,N_2008);
nor U2802 (N_2802,N_2320,N_2105);
or U2803 (N_2803,N_2129,N_2144);
xnor U2804 (N_2804,N_2047,N_1875);
xor U2805 (N_2805,N_1840,N_2376);
or U2806 (N_2806,N_2231,N_1975);
nand U2807 (N_2807,N_2073,N_2117);
nand U2808 (N_2808,N_2234,N_2130);
or U2809 (N_2809,N_2336,N_2230);
xnor U2810 (N_2810,N_1940,N_2012);
nand U2811 (N_2811,N_2240,N_2006);
and U2812 (N_2812,N_1907,N_1989);
or U2813 (N_2813,N_1919,N_1804);
nor U2814 (N_2814,N_1903,N_1943);
xor U2815 (N_2815,N_2355,N_2060);
nor U2816 (N_2816,N_1951,N_2364);
nand U2817 (N_2817,N_2284,N_2337);
nand U2818 (N_2818,N_1818,N_2219);
and U2819 (N_2819,N_1936,N_2229);
xnor U2820 (N_2820,N_1868,N_2143);
nor U2821 (N_2821,N_1910,N_2059);
and U2822 (N_2822,N_1970,N_2391);
xnor U2823 (N_2823,N_1815,N_2291);
nand U2824 (N_2824,N_2215,N_2202);
nor U2825 (N_2825,N_1902,N_2238);
nor U2826 (N_2826,N_1836,N_2223);
nand U2827 (N_2827,N_1957,N_1827);
and U2828 (N_2828,N_1964,N_2022);
xnor U2829 (N_2829,N_2274,N_2248);
nor U2830 (N_2830,N_2283,N_2136);
and U2831 (N_2831,N_1958,N_1844);
or U2832 (N_2832,N_1842,N_1992);
or U2833 (N_2833,N_1832,N_1860);
or U2834 (N_2834,N_1862,N_2357);
nor U2835 (N_2835,N_1810,N_1813);
or U2836 (N_2836,N_2145,N_1969);
nand U2837 (N_2837,N_1946,N_2206);
xor U2838 (N_2838,N_2213,N_2109);
nor U2839 (N_2839,N_2278,N_1994);
xnor U2840 (N_2840,N_2348,N_1839);
and U2841 (N_2841,N_2153,N_2391);
and U2842 (N_2842,N_2026,N_1852);
nand U2843 (N_2843,N_2228,N_1970);
nor U2844 (N_2844,N_2224,N_2281);
and U2845 (N_2845,N_1914,N_1878);
nand U2846 (N_2846,N_2216,N_2049);
and U2847 (N_2847,N_1895,N_2061);
xor U2848 (N_2848,N_1881,N_1815);
or U2849 (N_2849,N_2079,N_2061);
nor U2850 (N_2850,N_1970,N_2277);
and U2851 (N_2851,N_2335,N_2386);
nand U2852 (N_2852,N_1811,N_2185);
nor U2853 (N_2853,N_2000,N_1855);
or U2854 (N_2854,N_2255,N_1916);
nand U2855 (N_2855,N_1824,N_2137);
xor U2856 (N_2856,N_2322,N_2317);
xor U2857 (N_2857,N_2128,N_1845);
nand U2858 (N_2858,N_2155,N_1845);
nor U2859 (N_2859,N_2006,N_2366);
nand U2860 (N_2860,N_1852,N_2350);
xor U2861 (N_2861,N_2299,N_1944);
nand U2862 (N_2862,N_2229,N_2038);
or U2863 (N_2863,N_2353,N_2266);
nor U2864 (N_2864,N_2218,N_1883);
and U2865 (N_2865,N_2122,N_1998);
or U2866 (N_2866,N_2059,N_2322);
nor U2867 (N_2867,N_2358,N_2227);
and U2868 (N_2868,N_2272,N_2263);
and U2869 (N_2869,N_2152,N_1841);
or U2870 (N_2870,N_2363,N_2299);
or U2871 (N_2871,N_1805,N_2385);
nand U2872 (N_2872,N_2264,N_1837);
xnor U2873 (N_2873,N_2317,N_1884);
nand U2874 (N_2874,N_1898,N_1838);
xor U2875 (N_2875,N_1930,N_2055);
or U2876 (N_2876,N_1890,N_2030);
nand U2877 (N_2877,N_2104,N_2199);
xor U2878 (N_2878,N_2266,N_2100);
or U2879 (N_2879,N_2188,N_1965);
and U2880 (N_2880,N_2227,N_2369);
and U2881 (N_2881,N_1829,N_2301);
nor U2882 (N_2882,N_2349,N_2294);
nand U2883 (N_2883,N_2095,N_2048);
or U2884 (N_2884,N_1807,N_1870);
and U2885 (N_2885,N_1823,N_1923);
nor U2886 (N_2886,N_2175,N_1813);
or U2887 (N_2887,N_2022,N_2161);
and U2888 (N_2888,N_1947,N_1945);
and U2889 (N_2889,N_2019,N_2255);
or U2890 (N_2890,N_1971,N_1881);
and U2891 (N_2891,N_2281,N_2116);
nand U2892 (N_2892,N_2082,N_2189);
and U2893 (N_2893,N_2074,N_1862);
nor U2894 (N_2894,N_1916,N_2132);
nand U2895 (N_2895,N_1858,N_2142);
or U2896 (N_2896,N_2354,N_1975);
or U2897 (N_2897,N_2187,N_1827);
xnor U2898 (N_2898,N_1920,N_2079);
xor U2899 (N_2899,N_2287,N_2165);
or U2900 (N_2900,N_1921,N_2045);
nand U2901 (N_2901,N_2174,N_1894);
nand U2902 (N_2902,N_2376,N_2300);
nor U2903 (N_2903,N_1822,N_1937);
or U2904 (N_2904,N_2207,N_1852);
nand U2905 (N_2905,N_2388,N_2240);
nor U2906 (N_2906,N_1881,N_2057);
or U2907 (N_2907,N_1834,N_2377);
nor U2908 (N_2908,N_1803,N_2216);
or U2909 (N_2909,N_2244,N_2036);
or U2910 (N_2910,N_1905,N_1972);
and U2911 (N_2911,N_2364,N_2188);
or U2912 (N_2912,N_2293,N_1968);
nand U2913 (N_2913,N_1935,N_2334);
xor U2914 (N_2914,N_2002,N_2046);
nand U2915 (N_2915,N_2109,N_2140);
xnor U2916 (N_2916,N_2387,N_2172);
or U2917 (N_2917,N_1947,N_1913);
and U2918 (N_2918,N_2336,N_1988);
and U2919 (N_2919,N_1835,N_1819);
nor U2920 (N_2920,N_1981,N_2352);
or U2921 (N_2921,N_2392,N_1954);
xnor U2922 (N_2922,N_2005,N_2061);
nand U2923 (N_2923,N_2130,N_1864);
or U2924 (N_2924,N_1958,N_2313);
and U2925 (N_2925,N_1895,N_2038);
and U2926 (N_2926,N_2368,N_2229);
nor U2927 (N_2927,N_2200,N_2030);
nand U2928 (N_2928,N_1888,N_1908);
nand U2929 (N_2929,N_1877,N_2392);
or U2930 (N_2930,N_2282,N_2031);
nor U2931 (N_2931,N_1958,N_2013);
and U2932 (N_2932,N_2292,N_2103);
xnor U2933 (N_2933,N_2078,N_2035);
xor U2934 (N_2934,N_1928,N_2277);
nor U2935 (N_2935,N_1951,N_2224);
nand U2936 (N_2936,N_2100,N_2332);
xor U2937 (N_2937,N_2385,N_2347);
nor U2938 (N_2938,N_2002,N_2385);
or U2939 (N_2939,N_2114,N_2103);
xnor U2940 (N_2940,N_1943,N_1855);
xor U2941 (N_2941,N_2399,N_2254);
or U2942 (N_2942,N_2305,N_2342);
or U2943 (N_2943,N_2081,N_1868);
xor U2944 (N_2944,N_2122,N_2001);
nand U2945 (N_2945,N_1959,N_1862);
xor U2946 (N_2946,N_1972,N_2009);
xor U2947 (N_2947,N_2234,N_1914);
nor U2948 (N_2948,N_2043,N_2334);
and U2949 (N_2949,N_2219,N_2212);
and U2950 (N_2950,N_2389,N_1982);
nand U2951 (N_2951,N_1984,N_1821);
xnor U2952 (N_2952,N_2236,N_2142);
nor U2953 (N_2953,N_2146,N_1952);
xnor U2954 (N_2954,N_1882,N_1843);
and U2955 (N_2955,N_2118,N_2243);
or U2956 (N_2956,N_2184,N_2127);
or U2957 (N_2957,N_2336,N_1909);
and U2958 (N_2958,N_2251,N_2064);
and U2959 (N_2959,N_1951,N_2001);
xnor U2960 (N_2960,N_2044,N_2054);
nand U2961 (N_2961,N_2023,N_2050);
xnor U2962 (N_2962,N_2173,N_2258);
and U2963 (N_2963,N_2307,N_1874);
nand U2964 (N_2964,N_1883,N_1959);
nand U2965 (N_2965,N_1819,N_2321);
nor U2966 (N_2966,N_2229,N_1970);
or U2967 (N_2967,N_2172,N_2058);
xor U2968 (N_2968,N_1803,N_1819);
and U2969 (N_2969,N_2032,N_1977);
nor U2970 (N_2970,N_2135,N_1870);
nor U2971 (N_2971,N_1815,N_1907);
nand U2972 (N_2972,N_2226,N_2296);
nor U2973 (N_2973,N_2250,N_1995);
xor U2974 (N_2974,N_2358,N_2305);
or U2975 (N_2975,N_2366,N_2130);
nand U2976 (N_2976,N_1861,N_2205);
xnor U2977 (N_2977,N_1803,N_1942);
or U2978 (N_2978,N_2350,N_2380);
or U2979 (N_2979,N_2332,N_2128);
nor U2980 (N_2980,N_2028,N_1933);
xnor U2981 (N_2981,N_2267,N_2141);
nor U2982 (N_2982,N_2257,N_2116);
and U2983 (N_2983,N_2316,N_1942);
nand U2984 (N_2984,N_2031,N_2106);
nor U2985 (N_2985,N_1844,N_2188);
nor U2986 (N_2986,N_2193,N_1990);
nand U2987 (N_2987,N_2085,N_2126);
and U2988 (N_2988,N_1880,N_2397);
or U2989 (N_2989,N_2246,N_2315);
xnor U2990 (N_2990,N_2205,N_1875);
and U2991 (N_2991,N_1949,N_2077);
or U2992 (N_2992,N_2152,N_2176);
xnor U2993 (N_2993,N_1885,N_2116);
and U2994 (N_2994,N_1926,N_2069);
and U2995 (N_2995,N_1938,N_2218);
nor U2996 (N_2996,N_2226,N_2203);
xor U2997 (N_2997,N_2249,N_1930);
nand U2998 (N_2998,N_2105,N_1903);
or U2999 (N_2999,N_2020,N_2371);
xor U3000 (N_3000,N_2895,N_2767);
and U3001 (N_3001,N_2465,N_2694);
and U3002 (N_3002,N_2860,N_2616);
nand U3003 (N_3003,N_2660,N_2706);
xor U3004 (N_3004,N_2693,N_2984);
nor U3005 (N_3005,N_2586,N_2635);
or U3006 (N_3006,N_2854,N_2549);
nor U3007 (N_3007,N_2638,N_2550);
or U3008 (N_3008,N_2736,N_2732);
xnor U3009 (N_3009,N_2816,N_2653);
nand U3010 (N_3010,N_2527,N_2900);
xnor U3011 (N_3011,N_2750,N_2837);
xor U3012 (N_3012,N_2946,N_2562);
and U3013 (N_3013,N_2713,N_2541);
xnor U3014 (N_3014,N_2899,N_2523);
xnor U3015 (N_3015,N_2494,N_2986);
nor U3016 (N_3016,N_2789,N_2591);
xor U3017 (N_3017,N_2720,N_2651);
nor U3018 (N_3018,N_2463,N_2457);
nand U3019 (N_3019,N_2668,N_2740);
xnor U3020 (N_3020,N_2614,N_2451);
or U3021 (N_3021,N_2864,N_2561);
nand U3022 (N_3022,N_2798,N_2421);
or U3023 (N_3023,N_2546,N_2411);
or U3024 (N_3024,N_2566,N_2771);
nor U3025 (N_3025,N_2743,N_2585);
nand U3026 (N_3026,N_2512,N_2469);
nand U3027 (N_3027,N_2746,N_2803);
nor U3028 (N_3028,N_2593,N_2695);
and U3029 (N_3029,N_2924,N_2447);
or U3030 (N_3030,N_2877,N_2472);
and U3031 (N_3031,N_2827,N_2839);
and U3032 (N_3032,N_2871,N_2489);
xnor U3033 (N_3033,N_2431,N_2733);
or U3034 (N_3034,N_2838,N_2683);
and U3035 (N_3035,N_2701,N_2788);
or U3036 (N_3036,N_2499,N_2406);
or U3037 (N_3037,N_2920,N_2824);
and U3038 (N_3038,N_2475,N_2450);
nand U3039 (N_3039,N_2934,N_2973);
and U3040 (N_3040,N_2907,N_2482);
nor U3041 (N_3041,N_2948,N_2604);
nor U3042 (N_3042,N_2575,N_2843);
and U3043 (N_3043,N_2887,N_2560);
xnor U3044 (N_3044,N_2811,N_2665);
or U3045 (N_3045,N_2744,N_2676);
nand U3046 (N_3046,N_2505,N_2945);
nor U3047 (N_3047,N_2894,N_2699);
nor U3048 (N_3048,N_2805,N_2808);
xnor U3049 (N_3049,N_2800,N_2570);
or U3050 (N_3050,N_2675,N_2865);
or U3051 (N_3051,N_2690,N_2495);
and U3052 (N_3052,N_2987,N_2802);
and U3053 (N_3053,N_2982,N_2405);
and U3054 (N_3054,N_2884,N_2832);
nand U3055 (N_3055,N_2878,N_2914);
xor U3056 (N_3056,N_2939,N_2974);
or U3057 (N_3057,N_2497,N_2813);
nor U3058 (N_3058,N_2415,N_2563);
or U3059 (N_3059,N_2503,N_2420);
or U3060 (N_3060,N_2815,N_2703);
and U3061 (N_3061,N_2967,N_2569);
xnor U3062 (N_3062,N_2810,N_2678);
and U3063 (N_3063,N_2526,N_2904);
xnor U3064 (N_3064,N_2932,N_2613);
xnor U3065 (N_3065,N_2507,N_2674);
or U3066 (N_3066,N_2949,N_2427);
nand U3067 (N_3067,N_2915,N_2756);
xnor U3068 (N_3068,N_2545,N_2990);
and U3069 (N_3069,N_2677,N_2574);
and U3070 (N_3070,N_2705,N_2953);
xnor U3071 (N_3071,N_2539,N_2455);
or U3072 (N_3072,N_2826,N_2985);
or U3073 (N_3073,N_2516,N_2414);
and U3074 (N_3074,N_2589,N_2625);
or U3075 (N_3075,N_2474,N_2478);
or U3076 (N_3076,N_2799,N_2530);
nor U3077 (N_3077,N_2961,N_2938);
xor U3078 (N_3078,N_2761,N_2902);
xor U3079 (N_3079,N_2654,N_2662);
nand U3080 (N_3080,N_2916,N_2568);
nand U3081 (N_3081,N_2922,N_2599);
or U3082 (N_3082,N_2460,N_2734);
or U3083 (N_3083,N_2901,N_2954);
and U3084 (N_3084,N_2712,N_2477);
xor U3085 (N_3085,N_2684,N_2632);
or U3086 (N_3086,N_2708,N_2490);
and U3087 (N_3087,N_2883,N_2829);
xnor U3088 (N_3088,N_2881,N_2951);
nor U3089 (N_3089,N_2640,N_2404);
and U3090 (N_3090,N_2617,N_2501);
and U3091 (N_3091,N_2500,N_2966);
or U3092 (N_3092,N_2791,N_2862);
or U3093 (N_3093,N_2959,N_2778);
nand U3094 (N_3094,N_2487,N_2971);
and U3095 (N_3095,N_2748,N_2646);
and U3096 (N_3096,N_2597,N_2812);
and U3097 (N_3097,N_2786,N_2511);
nand U3098 (N_3098,N_2913,N_2462);
xor U3099 (N_3099,N_2779,N_2538);
nand U3100 (N_3100,N_2680,N_2702);
nor U3101 (N_3101,N_2785,N_2458);
nor U3102 (N_3102,N_2598,N_2970);
xor U3103 (N_3103,N_2547,N_2825);
and U3104 (N_3104,N_2540,N_2636);
xnor U3105 (N_3105,N_2596,N_2848);
and U3106 (N_3106,N_2742,N_2728);
or U3107 (N_3107,N_2822,N_2518);
xnor U3108 (N_3108,N_2754,N_2735);
and U3109 (N_3109,N_2841,N_2558);
or U3110 (N_3110,N_2594,N_2775);
nand U3111 (N_3111,N_2697,N_2814);
nor U3112 (N_3112,N_2506,N_2429);
nand U3113 (N_3113,N_2857,N_2842);
or U3114 (N_3114,N_2739,N_2935);
nand U3115 (N_3115,N_2931,N_2714);
nand U3116 (N_3116,N_2764,N_2757);
or U3117 (N_3117,N_2644,N_2671);
and U3118 (N_3118,N_2473,N_2533);
or U3119 (N_3119,N_2797,N_2804);
and U3120 (N_3120,N_2769,N_2437);
or U3121 (N_3121,N_2760,N_2852);
or U3122 (N_3122,N_2820,N_2872);
or U3123 (N_3123,N_2715,N_2730);
xnor U3124 (N_3124,N_2962,N_2835);
or U3125 (N_3125,N_2433,N_2956);
nand U3126 (N_3126,N_2963,N_2861);
nor U3127 (N_3127,N_2484,N_2611);
nor U3128 (N_3128,N_2584,N_2532);
or U3129 (N_3129,N_2664,N_2819);
nand U3130 (N_3130,N_2576,N_2763);
nor U3131 (N_3131,N_2886,N_2968);
nor U3132 (N_3132,N_2544,N_2426);
nand U3133 (N_3133,N_2719,N_2551);
nor U3134 (N_3134,N_2759,N_2493);
and U3135 (N_3135,N_2737,N_2601);
nand U3136 (N_3136,N_2691,N_2943);
nand U3137 (N_3137,N_2833,N_2818);
xor U3138 (N_3138,N_2400,N_2855);
xnor U3139 (N_3139,N_2806,N_2555);
nor U3140 (N_3140,N_2423,N_2669);
and U3141 (N_3141,N_2731,N_2995);
and U3142 (N_3142,N_2766,N_2988);
or U3143 (N_3143,N_2777,N_2573);
xnor U3144 (N_3144,N_2896,N_2663);
xor U3145 (N_3145,N_2903,N_2793);
nor U3146 (N_3146,N_2911,N_2448);
nor U3147 (N_3147,N_2622,N_2496);
nor U3148 (N_3148,N_2758,N_2588);
nand U3149 (N_3149,N_2483,N_2882);
nor U3150 (N_3150,N_2738,N_2667);
or U3151 (N_3151,N_2722,N_2459);
xnor U3152 (N_3152,N_2942,N_2661);
or U3153 (N_3153,N_2687,N_2930);
nor U3154 (N_3154,N_2401,N_2836);
xor U3155 (N_3155,N_2643,N_2417);
nor U3156 (N_3156,N_2752,N_2554);
and U3157 (N_3157,N_2443,N_2755);
nor U3158 (N_3158,N_2908,N_2817);
or U3159 (N_3159,N_2762,N_2642);
nor U3160 (N_3160,N_2626,N_2940);
or U3161 (N_3161,N_2652,N_2947);
nand U3162 (N_3162,N_2504,N_2408);
xnor U3163 (N_3163,N_2823,N_2592);
xor U3164 (N_3164,N_2543,N_2958);
nor U3165 (N_3165,N_2912,N_2686);
or U3166 (N_3166,N_2941,N_2893);
nand U3167 (N_3167,N_2863,N_2553);
or U3168 (N_3168,N_2422,N_2960);
xor U3169 (N_3169,N_2944,N_2670);
and U3170 (N_3170,N_2655,N_2888);
nand U3171 (N_3171,N_2698,N_2453);
or U3172 (N_3172,N_2828,N_2579);
nand U3173 (N_3173,N_2741,N_2439);
nand U3174 (N_3174,N_2609,N_2726);
nor U3175 (N_3175,N_2851,N_2685);
and U3176 (N_3176,N_2929,N_2783);
nor U3177 (N_3177,N_2464,N_2502);
nand U3178 (N_3178,N_2917,N_2850);
nor U3179 (N_3179,N_2454,N_2991);
or U3180 (N_3180,N_2707,N_2745);
and U3181 (N_3181,N_2787,N_2679);
and U3182 (N_3182,N_2983,N_2795);
nor U3183 (N_3183,N_2476,N_2905);
nor U3184 (N_3184,N_2608,N_2976);
nand U3185 (N_3185,N_2753,N_2510);
or U3186 (N_3186,N_2773,N_2631);
nand U3187 (N_3187,N_2890,N_2909);
nor U3188 (N_3188,N_2681,N_2717);
nor U3189 (N_3189,N_2557,N_2481);
nor U3190 (N_3190,N_2710,N_2989);
nor U3191 (N_3191,N_2981,N_2774);
or U3192 (N_3192,N_2879,N_2898);
nand U3193 (N_3193,N_2416,N_2891);
and U3194 (N_3194,N_2790,N_2950);
or U3195 (N_3195,N_2996,N_2461);
nor U3196 (N_3196,N_2998,N_2537);
xnor U3197 (N_3197,N_2928,N_2784);
nor U3198 (N_3198,N_2466,N_2559);
or U3199 (N_3199,N_2765,N_2979);
xor U3200 (N_3200,N_2910,N_2689);
and U3201 (N_3201,N_2955,N_2456);
nor U3202 (N_3202,N_2615,N_2548);
or U3203 (N_3203,N_2468,N_2656);
xor U3204 (N_3204,N_2542,N_2424);
nor U3205 (N_3205,N_2446,N_2634);
nand U3206 (N_3206,N_2633,N_2925);
nand U3207 (N_3207,N_2868,N_2897);
nor U3208 (N_3208,N_2776,N_2564);
and U3209 (N_3209,N_2639,N_2696);
and U3210 (N_3210,N_2519,N_2610);
nand U3211 (N_3211,N_2418,N_2964);
and U3212 (N_3212,N_2413,N_2556);
nand U3213 (N_3213,N_2700,N_2874);
xnor U3214 (N_3214,N_2580,N_2844);
or U3215 (N_3215,N_2796,N_2866);
or U3216 (N_3216,N_2524,N_2650);
nand U3217 (N_3217,N_2749,N_2567);
xnor U3218 (N_3218,N_2867,N_2520);
nor U3219 (N_3219,N_2936,N_2620);
xnor U3220 (N_3220,N_2830,N_2587);
nor U3221 (N_3221,N_2921,N_2666);
and U3222 (N_3222,N_2618,N_2727);
and U3223 (N_3223,N_2906,N_2847);
xnor U3224 (N_3224,N_2972,N_2999);
xnor U3225 (N_3225,N_2965,N_2794);
xor U3226 (N_3226,N_2870,N_2607);
xnor U3227 (N_3227,N_2629,N_2647);
xor U3228 (N_3228,N_2889,N_2704);
nand U3229 (N_3229,N_2657,N_2412);
or U3230 (N_3230,N_2623,N_2821);
and U3231 (N_3231,N_2438,N_2770);
xor U3232 (N_3232,N_2442,N_2600);
xor U3233 (N_3233,N_2926,N_2581);
nor U3234 (N_3234,N_2430,N_2649);
nand U3235 (N_3235,N_2977,N_2969);
or U3236 (N_3236,N_2612,N_2432);
and U3237 (N_3237,N_2491,N_2792);
and U3238 (N_3238,N_2434,N_2637);
nor U3239 (N_3239,N_2859,N_2853);
and U3240 (N_3240,N_2856,N_2724);
nor U3241 (N_3241,N_2873,N_2403);
and U3242 (N_3242,N_2630,N_2440);
nor U3243 (N_3243,N_2809,N_2711);
nand U3244 (N_3244,N_2428,N_2692);
and U3245 (N_3245,N_2577,N_2845);
or U3246 (N_3246,N_2492,N_2508);
nand U3247 (N_3247,N_2840,N_2552);
nand U3248 (N_3248,N_2768,N_2590);
nand U3249 (N_3249,N_2658,N_2688);
nand U3250 (N_3250,N_2880,N_2565);
and U3251 (N_3251,N_2927,N_2409);
and U3252 (N_3252,N_2498,N_2535);
and U3253 (N_3253,N_2531,N_2673);
and U3254 (N_3254,N_2645,N_2470);
nor U3255 (N_3255,N_2975,N_2725);
nor U3256 (N_3256,N_2751,N_2444);
nor U3257 (N_3257,N_2875,N_2919);
xor U3258 (N_3258,N_2571,N_2407);
xor U3259 (N_3259,N_2488,N_2858);
xor U3260 (N_3260,N_2957,N_2436);
and U3261 (N_3261,N_2606,N_2486);
or U3262 (N_3262,N_2892,N_2595);
nand U3263 (N_3263,N_2513,N_2933);
or U3264 (N_3264,N_2410,N_2509);
and U3265 (N_3265,N_2993,N_2992);
nand U3266 (N_3266,N_2782,N_2718);
and U3267 (N_3267,N_2515,N_2849);
nand U3268 (N_3268,N_2723,N_2521);
and U3269 (N_3269,N_2807,N_2525);
xnor U3270 (N_3270,N_2952,N_2452);
or U3271 (N_3271,N_2831,N_2978);
nor U3272 (N_3272,N_2628,N_2682);
and U3273 (N_3273,N_2846,N_2449);
nand U3274 (N_3274,N_2834,N_2747);
nand U3275 (N_3275,N_2923,N_2534);
and U3276 (N_3276,N_2619,N_2659);
nand U3277 (N_3277,N_2709,N_2721);
or U3278 (N_3278,N_2435,N_2994);
xor U3279 (N_3279,N_2419,N_2578);
and U3280 (N_3280,N_2572,N_2402);
or U3281 (N_3281,N_2514,N_2641);
nand U3282 (N_3282,N_2479,N_2729);
nor U3283 (N_3283,N_2869,N_2624);
nor U3284 (N_3284,N_2937,N_2485);
xor U3285 (N_3285,N_2517,N_2522);
or U3286 (N_3286,N_2536,N_2780);
xnor U3287 (N_3287,N_2602,N_2583);
xnor U3288 (N_3288,N_2441,N_2621);
nor U3289 (N_3289,N_2605,N_2918);
and U3290 (N_3290,N_2425,N_2997);
nor U3291 (N_3291,N_2528,N_2529);
xor U3292 (N_3292,N_2781,N_2648);
nor U3293 (N_3293,N_2876,N_2480);
or U3294 (N_3294,N_2627,N_2467);
and U3295 (N_3295,N_2980,N_2582);
nor U3296 (N_3296,N_2716,N_2885);
nand U3297 (N_3297,N_2445,N_2772);
nor U3298 (N_3298,N_2801,N_2672);
xnor U3299 (N_3299,N_2471,N_2603);
nor U3300 (N_3300,N_2613,N_2562);
xnor U3301 (N_3301,N_2860,N_2438);
nor U3302 (N_3302,N_2626,N_2764);
and U3303 (N_3303,N_2648,N_2634);
nand U3304 (N_3304,N_2802,N_2755);
nor U3305 (N_3305,N_2908,N_2731);
or U3306 (N_3306,N_2965,N_2864);
xor U3307 (N_3307,N_2528,N_2744);
xor U3308 (N_3308,N_2604,N_2906);
nand U3309 (N_3309,N_2739,N_2877);
or U3310 (N_3310,N_2826,N_2591);
nand U3311 (N_3311,N_2943,N_2445);
and U3312 (N_3312,N_2606,N_2774);
xor U3313 (N_3313,N_2588,N_2509);
xor U3314 (N_3314,N_2811,N_2610);
or U3315 (N_3315,N_2884,N_2868);
xor U3316 (N_3316,N_2604,N_2573);
and U3317 (N_3317,N_2778,N_2822);
or U3318 (N_3318,N_2595,N_2526);
xor U3319 (N_3319,N_2526,N_2850);
nor U3320 (N_3320,N_2681,N_2726);
and U3321 (N_3321,N_2499,N_2878);
nand U3322 (N_3322,N_2400,N_2718);
nand U3323 (N_3323,N_2450,N_2455);
or U3324 (N_3324,N_2633,N_2668);
and U3325 (N_3325,N_2507,N_2534);
nand U3326 (N_3326,N_2602,N_2715);
nor U3327 (N_3327,N_2740,N_2955);
or U3328 (N_3328,N_2805,N_2822);
nor U3329 (N_3329,N_2491,N_2760);
or U3330 (N_3330,N_2822,N_2889);
nor U3331 (N_3331,N_2588,N_2717);
and U3332 (N_3332,N_2677,N_2998);
and U3333 (N_3333,N_2513,N_2484);
nand U3334 (N_3334,N_2777,N_2737);
or U3335 (N_3335,N_2479,N_2912);
xor U3336 (N_3336,N_2455,N_2987);
nor U3337 (N_3337,N_2875,N_2885);
or U3338 (N_3338,N_2525,N_2729);
nor U3339 (N_3339,N_2962,N_2415);
and U3340 (N_3340,N_2842,N_2484);
xnor U3341 (N_3341,N_2716,N_2757);
and U3342 (N_3342,N_2920,N_2793);
nor U3343 (N_3343,N_2986,N_2422);
xnor U3344 (N_3344,N_2437,N_2522);
nand U3345 (N_3345,N_2474,N_2465);
nand U3346 (N_3346,N_2981,N_2786);
or U3347 (N_3347,N_2421,N_2922);
nand U3348 (N_3348,N_2812,N_2789);
nor U3349 (N_3349,N_2411,N_2531);
and U3350 (N_3350,N_2727,N_2804);
nor U3351 (N_3351,N_2872,N_2812);
xor U3352 (N_3352,N_2520,N_2573);
nor U3353 (N_3353,N_2705,N_2521);
xor U3354 (N_3354,N_2999,N_2748);
xnor U3355 (N_3355,N_2796,N_2747);
and U3356 (N_3356,N_2857,N_2701);
xnor U3357 (N_3357,N_2544,N_2576);
or U3358 (N_3358,N_2480,N_2715);
nand U3359 (N_3359,N_2775,N_2979);
xor U3360 (N_3360,N_2598,N_2536);
nand U3361 (N_3361,N_2594,N_2975);
nor U3362 (N_3362,N_2636,N_2933);
nand U3363 (N_3363,N_2597,N_2581);
or U3364 (N_3364,N_2794,N_2886);
and U3365 (N_3365,N_2668,N_2656);
nor U3366 (N_3366,N_2488,N_2843);
or U3367 (N_3367,N_2693,N_2646);
and U3368 (N_3368,N_2488,N_2601);
nand U3369 (N_3369,N_2712,N_2434);
nand U3370 (N_3370,N_2616,N_2713);
xnor U3371 (N_3371,N_2969,N_2835);
and U3372 (N_3372,N_2469,N_2823);
or U3373 (N_3373,N_2958,N_2784);
xnor U3374 (N_3374,N_2635,N_2579);
or U3375 (N_3375,N_2462,N_2779);
xnor U3376 (N_3376,N_2497,N_2633);
nand U3377 (N_3377,N_2723,N_2753);
nor U3378 (N_3378,N_2797,N_2936);
xor U3379 (N_3379,N_2444,N_2485);
or U3380 (N_3380,N_2690,N_2998);
xnor U3381 (N_3381,N_2468,N_2644);
nor U3382 (N_3382,N_2975,N_2638);
and U3383 (N_3383,N_2464,N_2713);
xor U3384 (N_3384,N_2748,N_2509);
nand U3385 (N_3385,N_2995,N_2855);
or U3386 (N_3386,N_2531,N_2628);
or U3387 (N_3387,N_2460,N_2676);
nand U3388 (N_3388,N_2611,N_2587);
or U3389 (N_3389,N_2654,N_2957);
nor U3390 (N_3390,N_2435,N_2915);
or U3391 (N_3391,N_2928,N_2821);
xnor U3392 (N_3392,N_2540,N_2477);
xnor U3393 (N_3393,N_2824,N_2687);
or U3394 (N_3394,N_2995,N_2876);
or U3395 (N_3395,N_2821,N_2539);
nor U3396 (N_3396,N_2873,N_2563);
or U3397 (N_3397,N_2751,N_2697);
or U3398 (N_3398,N_2822,N_2952);
and U3399 (N_3399,N_2487,N_2838);
nor U3400 (N_3400,N_2770,N_2409);
and U3401 (N_3401,N_2728,N_2951);
nor U3402 (N_3402,N_2470,N_2440);
or U3403 (N_3403,N_2530,N_2775);
nand U3404 (N_3404,N_2844,N_2620);
nand U3405 (N_3405,N_2774,N_2799);
or U3406 (N_3406,N_2986,N_2939);
or U3407 (N_3407,N_2946,N_2623);
nand U3408 (N_3408,N_2942,N_2502);
xor U3409 (N_3409,N_2888,N_2616);
xnor U3410 (N_3410,N_2588,N_2901);
xnor U3411 (N_3411,N_2953,N_2768);
xnor U3412 (N_3412,N_2425,N_2701);
nor U3413 (N_3413,N_2675,N_2422);
nand U3414 (N_3414,N_2480,N_2457);
xor U3415 (N_3415,N_2993,N_2745);
nor U3416 (N_3416,N_2833,N_2616);
nor U3417 (N_3417,N_2613,N_2624);
nand U3418 (N_3418,N_2805,N_2993);
nor U3419 (N_3419,N_2773,N_2607);
nor U3420 (N_3420,N_2902,N_2651);
nor U3421 (N_3421,N_2777,N_2656);
or U3422 (N_3422,N_2680,N_2571);
or U3423 (N_3423,N_2903,N_2788);
nor U3424 (N_3424,N_2797,N_2694);
and U3425 (N_3425,N_2456,N_2937);
or U3426 (N_3426,N_2505,N_2700);
or U3427 (N_3427,N_2895,N_2702);
and U3428 (N_3428,N_2603,N_2860);
nand U3429 (N_3429,N_2507,N_2422);
nor U3430 (N_3430,N_2572,N_2908);
nor U3431 (N_3431,N_2759,N_2814);
and U3432 (N_3432,N_2536,N_2813);
and U3433 (N_3433,N_2529,N_2729);
xor U3434 (N_3434,N_2587,N_2600);
nand U3435 (N_3435,N_2930,N_2923);
nand U3436 (N_3436,N_2620,N_2654);
nand U3437 (N_3437,N_2595,N_2657);
xor U3438 (N_3438,N_2834,N_2463);
xnor U3439 (N_3439,N_2543,N_2723);
or U3440 (N_3440,N_2738,N_2508);
nand U3441 (N_3441,N_2656,N_2510);
nor U3442 (N_3442,N_2753,N_2817);
nor U3443 (N_3443,N_2695,N_2846);
xnor U3444 (N_3444,N_2944,N_2543);
nand U3445 (N_3445,N_2562,N_2510);
xnor U3446 (N_3446,N_2792,N_2888);
nand U3447 (N_3447,N_2600,N_2983);
and U3448 (N_3448,N_2735,N_2719);
xor U3449 (N_3449,N_2928,N_2831);
and U3450 (N_3450,N_2629,N_2532);
or U3451 (N_3451,N_2682,N_2926);
nand U3452 (N_3452,N_2406,N_2977);
and U3453 (N_3453,N_2779,N_2524);
nor U3454 (N_3454,N_2456,N_2611);
and U3455 (N_3455,N_2592,N_2726);
and U3456 (N_3456,N_2604,N_2871);
nor U3457 (N_3457,N_2966,N_2598);
nor U3458 (N_3458,N_2768,N_2832);
and U3459 (N_3459,N_2882,N_2828);
and U3460 (N_3460,N_2577,N_2675);
or U3461 (N_3461,N_2433,N_2487);
nand U3462 (N_3462,N_2481,N_2712);
xor U3463 (N_3463,N_2769,N_2545);
nor U3464 (N_3464,N_2417,N_2816);
xor U3465 (N_3465,N_2405,N_2703);
and U3466 (N_3466,N_2821,N_2601);
xor U3467 (N_3467,N_2738,N_2476);
nand U3468 (N_3468,N_2437,N_2488);
nand U3469 (N_3469,N_2860,N_2910);
xor U3470 (N_3470,N_2856,N_2536);
or U3471 (N_3471,N_2681,N_2713);
or U3472 (N_3472,N_2685,N_2451);
and U3473 (N_3473,N_2491,N_2988);
or U3474 (N_3474,N_2576,N_2852);
and U3475 (N_3475,N_2698,N_2717);
or U3476 (N_3476,N_2528,N_2983);
xnor U3477 (N_3477,N_2966,N_2730);
and U3478 (N_3478,N_2528,N_2545);
or U3479 (N_3479,N_2620,N_2514);
nor U3480 (N_3480,N_2994,N_2923);
nor U3481 (N_3481,N_2514,N_2728);
xnor U3482 (N_3482,N_2876,N_2801);
or U3483 (N_3483,N_2574,N_2436);
nand U3484 (N_3484,N_2997,N_2922);
or U3485 (N_3485,N_2654,N_2702);
nand U3486 (N_3486,N_2678,N_2898);
and U3487 (N_3487,N_2830,N_2723);
and U3488 (N_3488,N_2456,N_2907);
nor U3489 (N_3489,N_2899,N_2894);
nor U3490 (N_3490,N_2868,N_2883);
nand U3491 (N_3491,N_2548,N_2877);
or U3492 (N_3492,N_2792,N_2590);
xnor U3493 (N_3493,N_2881,N_2814);
nand U3494 (N_3494,N_2688,N_2814);
and U3495 (N_3495,N_2658,N_2520);
nor U3496 (N_3496,N_2829,N_2832);
and U3497 (N_3497,N_2669,N_2927);
nand U3498 (N_3498,N_2529,N_2714);
or U3499 (N_3499,N_2688,N_2520);
or U3500 (N_3500,N_2666,N_2628);
nor U3501 (N_3501,N_2799,N_2592);
nand U3502 (N_3502,N_2893,N_2446);
nand U3503 (N_3503,N_2974,N_2975);
xor U3504 (N_3504,N_2672,N_2693);
nand U3505 (N_3505,N_2808,N_2877);
xor U3506 (N_3506,N_2490,N_2481);
xnor U3507 (N_3507,N_2936,N_2881);
nor U3508 (N_3508,N_2670,N_2614);
or U3509 (N_3509,N_2623,N_2408);
nor U3510 (N_3510,N_2529,N_2748);
or U3511 (N_3511,N_2878,N_2596);
and U3512 (N_3512,N_2791,N_2553);
nor U3513 (N_3513,N_2693,N_2920);
or U3514 (N_3514,N_2989,N_2946);
and U3515 (N_3515,N_2557,N_2791);
nor U3516 (N_3516,N_2825,N_2800);
or U3517 (N_3517,N_2702,N_2871);
or U3518 (N_3518,N_2502,N_2588);
nor U3519 (N_3519,N_2651,N_2938);
xnor U3520 (N_3520,N_2831,N_2879);
nor U3521 (N_3521,N_2639,N_2811);
xor U3522 (N_3522,N_2623,N_2547);
xnor U3523 (N_3523,N_2993,N_2565);
nand U3524 (N_3524,N_2869,N_2770);
and U3525 (N_3525,N_2721,N_2663);
and U3526 (N_3526,N_2701,N_2643);
and U3527 (N_3527,N_2682,N_2592);
xnor U3528 (N_3528,N_2889,N_2695);
and U3529 (N_3529,N_2598,N_2556);
and U3530 (N_3530,N_2776,N_2705);
xor U3531 (N_3531,N_2406,N_2568);
xnor U3532 (N_3532,N_2543,N_2977);
or U3533 (N_3533,N_2820,N_2553);
nor U3534 (N_3534,N_2849,N_2453);
or U3535 (N_3535,N_2900,N_2407);
or U3536 (N_3536,N_2656,N_2930);
xor U3537 (N_3537,N_2732,N_2763);
or U3538 (N_3538,N_2698,N_2832);
or U3539 (N_3539,N_2564,N_2798);
and U3540 (N_3540,N_2551,N_2511);
or U3541 (N_3541,N_2488,N_2482);
or U3542 (N_3542,N_2902,N_2523);
and U3543 (N_3543,N_2559,N_2474);
and U3544 (N_3544,N_2776,N_2888);
and U3545 (N_3545,N_2753,N_2605);
nand U3546 (N_3546,N_2539,N_2840);
nor U3547 (N_3547,N_2464,N_2679);
nand U3548 (N_3548,N_2418,N_2892);
and U3549 (N_3549,N_2942,N_2409);
xnor U3550 (N_3550,N_2425,N_2463);
nor U3551 (N_3551,N_2826,N_2695);
nor U3552 (N_3552,N_2409,N_2725);
or U3553 (N_3553,N_2429,N_2964);
and U3554 (N_3554,N_2595,N_2782);
xor U3555 (N_3555,N_2474,N_2411);
nor U3556 (N_3556,N_2866,N_2783);
or U3557 (N_3557,N_2741,N_2710);
xnor U3558 (N_3558,N_2481,N_2708);
xnor U3559 (N_3559,N_2663,N_2878);
xor U3560 (N_3560,N_2503,N_2977);
or U3561 (N_3561,N_2770,N_2653);
nand U3562 (N_3562,N_2752,N_2715);
or U3563 (N_3563,N_2763,N_2400);
or U3564 (N_3564,N_2732,N_2959);
and U3565 (N_3565,N_2949,N_2917);
or U3566 (N_3566,N_2941,N_2516);
or U3567 (N_3567,N_2521,N_2707);
or U3568 (N_3568,N_2593,N_2411);
xor U3569 (N_3569,N_2786,N_2955);
or U3570 (N_3570,N_2487,N_2794);
nor U3571 (N_3571,N_2808,N_2963);
and U3572 (N_3572,N_2605,N_2744);
nor U3573 (N_3573,N_2703,N_2627);
and U3574 (N_3574,N_2515,N_2977);
xor U3575 (N_3575,N_2911,N_2509);
nor U3576 (N_3576,N_2890,N_2902);
xor U3577 (N_3577,N_2442,N_2676);
and U3578 (N_3578,N_2831,N_2534);
nor U3579 (N_3579,N_2731,N_2912);
or U3580 (N_3580,N_2942,N_2557);
xor U3581 (N_3581,N_2923,N_2595);
and U3582 (N_3582,N_2989,N_2590);
and U3583 (N_3583,N_2621,N_2543);
xnor U3584 (N_3584,N_2892,N_2984);
nand U3585 (N_3585,N_2438,N_2451);
xnor U3586 (N_3586,N_2931,N_2871);
nor U3587 (N_3587,N_2492,N_2418);
nand U3588 (N_3588,N_2413,N_2884);
nor U3589 (N_3589,N_2967,N_2999);
or U3590 (N_3590,N_2775,N_2929);
or U3591 (N_3591,N_2562,N_2631);
or U3592 (N_3592,N_2549,N_2876);
and U3593 (N_3593,N_2514,N_2736);
and U3594 (N_3594,N_2407,N_2576);
xor U3595 (N_3595,N_2996,N_2410);
nor U3596 (N_3596,N_2558,N_2556);
xnor U3597 (N_3597,N_2563,N_2948);
or U3598 (N_3598,N_2688,N_2885);
nand U3599 (N_3599,N_2922,N_2622);
and U3600 (N_3600,N_3397,N_3596);
xnor U3601 (N_3601,N_3402,N_3300);
nand U3602 (N_3602,N_3020,N_3433);
xor U3603 (N_3603,N_3344,N_3113);
nand U3604 (N_3604,N_3352,N_3178);
xor U3605 (N_3605,N_3158,N_3540);
nand U3606 (N_3606,N_3006,N_3516);
xor U3607 (N_3607,N_3170,N_3521);
or U3608 (N_3608,N_3151,N_3353);
or U3609 (N_3609,N_3345,N_3434);
or U3610 (N_3610,N_3590,N_3532);
or U3611 (N_3611,N_3442,N_3138);
nor U3612 (N_3612,N_3340,N_3385);
nor U3613 (N_3613,N_3086,N_3401);
nand U3614 (N_3614,N_3470,N_3507);
and U3615 (N_3615,N_3337,N_3348);
nand U3616 (N_3616,N_3554,N_3363);
nand U3617 (N_3617,N_3387,N_3219);
nor U3618 (N_3618,N_3464,N_3196);
xnor U3619 (N_3619,N_3058,N_3110);
and U3620 (N_3620,N_3189,N_3088);
nand U3621 (N_3621,N_3479,N_3367);
nor U3622 (N_3622,N_3264,N_3114);
nand U3623 (N_3623,N_3395,N_3301);
xor U3624 (N_3624,N_3389,N_3034);
nand U3625 (N_3625,N_3068,N_3234);
nor U3626 (N_3626,N_3202,N_3533);
nor U3627 (N_3627,N_3223,N_3213);
nor U3628 (N_3628,N_3292,N_3326);
and U3629 (N_3629,N_3297,N_3510);
or U3630 (N_3630,N_3026,N_3280);
and U3631 (N_3631,N_3595,N_3023);
or U3632 (N_3632,N_3097,N_3080);
nand U3633 (N_3633,N_3274,N_3412);
nand U3634 (N_3634,N_3041,N_3495);
and U3635 (N_3635,N_3373,N_3181);
and U3636 (N_3636,N_3448,N_3262);
nand U3637 (N_3637,N_3298,N_3523);
or U3638 (N_3638,N_3032,N_3248);
nand U3639 (N_3639,N_3258,N_3406);
nor U3640 (N_3640,N_3116,N_3474);
nand U3641 (N_3641,N_3330,N_3037);
nor U3642 (N_3642,N_3318,N_3064);
nand U3643 (N_3643,N_3375,N_3166);
nor U3644 (N_3644,N_3514,N_3221);
and U3645 (N_3645,N_3529,N_3582);
nor U3646 (N_3646,N_3455,N_3033);
and U3647 (N_3647,N_3316,N_3545);
and U3648 (N_3648,N_3525,N_3293);
nand U3649 (N_3649,N_3518,N_3285);
and U3650 (N_3650,N_3548,N_3253);
or U3651 (N_3651,N_3534,N_3082);
or U3652 (N_3652,N_3208,N_3458);
or U3653 (N_3653,N_3559,N_3429);
xor U3654 (N_3654,N_3451,N_3384);
nand U3655 (N_3655,N_3530,N_3357);
or U3656 (N_3656,N_3200,N_3159);
and U3657 (N_3657,N_3441,N_3081);
or U3658 (N_3658,N_3177,N_3136);
xnor U3659 (N_3659,N_3155,N_3096);
nand U3660 (N_3660,N_3475,N_3594);
xnor U3661 (N_3661,N_3073,N_3065);
xor U3662 (N_3662,N_3564,N_3473);
or U3663 (N_3663,N_3124,N_3439);
nand U3664 (N_3664,N_3319,N_3520);
nor U3665 (N_3665,N_3445,N_3017);
nor U3666 (N_3666,N_3205,N_3162);
xor U3667 (N_3667,N_3211,N_3364);
nor U3668 (N_3668,N_3003,N_3522);
or U3669 (N_3669,N_3209,N_3431);
nor U3670 (N_3670,N_3444,N_3233);
xnor U3671 (N_3671,N_3569,N_3335);
nand U3672 (N_3672,N_3052,N_3583);
nor U3673 (N_3673,N_3598,N_3215);
nand U3674 (N_3674,N_3499,N_3550);
xor U3675 (N_3675,N_3361,N_3541);
nand U3676 (N_3676,N_3098,N_3030);
or U3677 (N_3677,N_3099,N_3180);
nand U3678 (N_3678,N_3415,N_3265);
or U3679 (N_3679,N_3449,N_3339);
and U3680 (N_3680,N_3537,N_3478);
and U3681 (N_3681,N_3046,N_3303);
or U3682 (N_3682,N_3383,N_3506);
or U3683 (N_3683,N_3558,N_3547);
xnor U3684 (N_3684,N_3074,N_3235);
nand U3685 (N_3685,N_3269,N_3167);
nand U3686 (N_3686,N_3149,N_3463);
and U3687 (N_3687,N_3505,N_3152);
and U3688 (N_3688,N_3562,N_3184);
nor U3689 (N_3689,N_3010,N_3408);
xnor U3690 (N_3690,N_3403,N_3242);
or U3691 (N_3691,N_3450,N_3131);
nor U3692 (N_3692,N_3414,N_3480);
nand U3693 (N_3693,N_3460,N_3029);
nor U3694 (N_3694,N_3176,N_3135);
nor U3695 (N_3695,N_3212,N_3091);
nand U3696 (N_3696,N_3296,N_3309);
nand U3697 (N_3697,N_3315,N_3440);
or U3698 (N_3698,N_3137,N_3005);
or U3699 (N_3699,N_3070,N_3536);
or U3700 (N_3700,N_3060,N_3174);
nor U3701 (N_3701,N_3491,N_3025);
and U3702 (N_3702,N_3272,N_3185);
xnor U3703 (N_3703,N_3524,N_3579);
or U3704 (N_3704,N_3063,N_3477);
nand U3705 (N_3705,N_3089,N_3322);
nand U3706 (N_3706,N_3454,N_3483);
nor U3707 (N_3707,N_3571,N_3508);
or U3708 (N_3708,N_3435,N_3061);
nor U3709 (N_3709,N_3323,N_3194);
nand U3710 (N_3710,N_3051,N_3188);
xnor U3711 (N_3711,N_3117,N_3586);
nor U3712 (N_3712,N_3038,N_3278);
xnor U3713 (N_3713,N_3376,N_3103);
xnor U3714 (N_3714,N_3511,N_3472);
xor U3715 (N_3715,N_3245,N_3427);
or U3716 (N_3716,N_3572,N_3009);
xnor U3717 (N_3717,N_3476,N_3372);
and U3718 (N_3718,N_3229,N_3336);
xor U3719 (N_3719,N_3587,N_3142);
nor U3720 (N_3720,N_3349,N_3047);
nor U3721 (N_3721,N_3589,N_3386);
xor U3722 (N_3722,N_3347,N_3066);
nand U3723 (N_3723,N_3462,N_3380);
nand U3724 (N_3724,N_3014,N_3565);
and U3725 (N_3725,N_3538,N_3260);
and U3726 (N_3726,N_3497,N_3365);
and U3727 (N_3727,N_3027,N_3090);
xnor U3728 (N_3728,N_3351,N_3069);
nor U3729 (N_3729,N_3161,N_3379);
xnor U3730 (N_3730,N_3581,N_3574);
and U3731 (N_3731,N_3527,N_3509);
nor U3732 (N_3732,N_3241,N_3231);
xnor U3733 (N_3733,N_3341,N_3216);
or U3734 (N_3734,N_3503,N_3101);
nor U3735 (N_3735,N_3261,N_3405);
or U3736 (N_3736,N_3360,N_3382);
and U3737 (N_3737,N_3201,N_3071);
and U3738 (N_3738,N_3546,N_3561);
and U3739 (N_3739,N_3273,N_3259);
nor U3740 (N_3740,N_3338,N_3588);
nand U3741 (N_3741,N_3053,N_3263);
and U3742 (N_3742,N_3346,N_3502);
or U3743 (N_3743,N_3206,N_3438);
xnor U3744 (N_3744,N_3123,N_3237);
nand U3745 (N_3745,N_3057,N_3542);
nor U3746 (N_3746,N_3410,N_3498);
nand U3747 (N_3747,N_3173,N_3390);
nor U3748 (N_3748,N_3218,N_3432);
xor U3749 (N_3749,N_3157,N_3459);
nor U3750 (N_3750,N_3591,N_3494);
and U3751 (N_3751,N_3004,N_3284);
nand U3752 (N_3752,N_3085,N_3428);
or U3753 (N_3753,N_3129,N_3002);
or U3754 (N_3754,N_3304,N_3560);
and U3755 (N_3755,N_3016,N_3453);
and U3756 (N_3756,N_3400,N_3175);
and U3757 (N_3757,N_3078,N_3493);
and U3758 (N_3758,N_3225,N_3133);
nand U3759 (N_3759,N_3062,N_3040);
or U3760 (N_3760,N_3100,N_3018);
nand U3761 (N_3761,N_3535,N_3250);
or U3762 (N_3762,N_3277,N_3011);
or U3763 (N_3763,N_3093,N_3420);
nor U3764 (N_3764,N_3366,N_3356);
and U3765 (N_3765,N_3371,N_3377);
or U3766 (N_3766,N_3031,N_3172);
xnor U3767 (N_3767,N_3299,N_3430);
and U3768 (N_3768,N_3312,N_3567);
xor U3769 (N_3769,N_3104,N_3224);
and U3770 (N_3770,N_3008,N_3059);
and U3771 (N_3771,N_3198,N_3394);
and U3772 (N_3772,N_3411,N_3313);
xnor U3773 (N_3773,N_3437,N_3199);
xor U3774 (N_3774,N_3305,N_3566);
nor U3775 (N_3775,N_3328,N_3019);
or U3776 (N_3776,N_3120,N_3381);
nand U3777 (N_3777,N_3544,N_3226);
xor U3778 (N_3778,N_3468,N_3079);
xor U3779 (N_3779,N_3324,N_3422);
and U3780 (N_3780,N_3119,N_3368);
nand U3781 (N_3781,N_3543,N_3257);
xor U3782 (N_3782,N_3094,N_3396);
xor U3783 (N_3783,N_3182,N_3236);
nor U3784 (N_3784,N_3306,N_3471);
or U3785 (N_3785,N_3592,N_3416);
xnor U3786 (N_3786,N_3585,N_3072);
xor U3787 (N_3787,N_3391,N_3552);
or U3788 (N_3788,N_3150,N_3148);
or U3789 (N_3789,N_3153,N_3580);
or U3790 (N_3790,N_3276,N_3238);
xor U3791 (N_3791,N_3388,N_3244);
or U3792 (N_3792,N_3426,N_3076);
xnor U3793 (N_3793,N_3147,N_3240);
nand U3794 (N_3794,N_3481,N_3169);
nand U3795 (N_3795,N_3557,N_3271);
nand U3796 (N_3796,N_3399,N_3268);
or U3797 (N_3797,N_3267,N_3279);
nor U3798 (N_3798,N_3597,N_3130);
nor U3799 (N_3799,N_3115,N_3168);
nor U3800 (N_3800,N_3127,N_3232);
nand U3801 (N_3801,N_3109,N_3593);
nor U3802 (N_3802,N_3486,N_3332);
nor U3803 (N_3803,N_3139,N_3049);
nor U3804 (N_3804,N_3055,N_3144);
nor U3805 (N_3805,N_3246,N_3111);
nor U3806 (N_3806,N_3022,N_3393);
nand U3807 (N_3807,N_3563,N_3197);
xor U3808 (N_3808,N_3001,N_3369);
nand U3809 (N_3809,N_3423,N_3482);
and U3810 (N_3810,N_3577,N_3156);
and U3811 (N_3811,N_3203,N_3436);
and U3812 (N_3812,N_3568,N_3140);
nand U3813 (N_3813,N_3256,N_3154);
nor U3814 (N_3814,N_3374,N_3370);
nand U3815 (N_3815,N_3287,N_3355);
xnor U3816 (N_3816,N_3321,N_3112);
nand U3817 (N_3817,N_3539,N_3252);
and U3818 (N_3818,N_3461,N_3465);
or U3819 (N_3819,N_3446,N_3302);
and U3820 (N_3820,N_3578,N_3378);
nand U3821 (N_3821,N_3083,N_3325);
and U3822 (N_3822,N_3492,N_3108);
nor U3823 (N_3823,N_3311,N_3329);
nand U3824 (N_3824,N_3043,N_3186);
xor U3825 (N_3825,N_3599,N_3488);
and U3826 (N_3826,N_3517,N_3171);
nor U3827 (N_3827,N_3500,N_3526);
xnor U3828 (N_3828,N_3036,N_3362);
nor U3829 (N_3829,N_3310,N_3556);
or U3830 (N_3830,N_3334,N_3024);
and U3831 (N_3831,N_3398,N_3570);
and U3832 (N_3832,N_3254,N_3289);
nand U3833 (N_3833,N_3469,N_3183);
nand U3834 (N_3834,N_3095,N_3122);
or U3835 (N_3835,N_3249,N_3295);
and U3836 (N_3836,N_3000,N_3443);
xnor U3837 (N_3837,N_3413,N_3307);
or U3838 (N_3838,N_3075,N_3121);
or U3839 (N_3839,N_3013,N_3584);
or U3840 (N_3840,N_3519,N_3504);
and U3841 (N_3841,N_3489,N_3214);
nor U3842 (N_3842,N_3456,N_3354);
or U3843 (N_3843,N_3195,N_3045);
nand U3844 (N_3844,N_3294,N_3496);
xnor U3845 (N_3845,N_3160,N_3515);
or U3846 (N_3846,N_3331,N_3012);
and U3847 (N_3847,N_3210,N_3359);
and U3848 (N_3848,N_3270,N_3164);
or U3849 (N_3849,N_3457,N_3467);
xnor U3850 (N_3850,N_3204,N_3192);
nand U3851 (N_3851,N_3501,N_3247);
nand U3852 (N_3852,N_3118,N_3409);
or U3853 (N_3853,N_3193,N_3283);
nor U3854 (N_3854,N_3134,N_3191);
nor U3855 (N_3855,N_3132,N_3466);
nand U3856 (N_3856,N_3243,N_3291);
nor U3857 (N_3857,N_3308,N_3054);
nand U3858 (N_3858,N_3419,N_3424);
and U3859 (N_3859,N_3190,N_3290);
nor U3860 (N_3860,N_3048,N_3576);
nor U3861 (N_3861,N_3417,N_3165);
or U3862 (N_3862,N_3230,N_3452);
nand U3863 (N_3863,N_3358,N_3125);
or U3864 (N_3864,N_3145,N_3084);
or U3865 (N_3865,N_3404,N_3421);
and U3866 (N_3866,N_3407,N_3551);
nor U3867 (N_3867,N_3126,N_3228);
nand U3868 (N_3868,N_3220,N_3227);
nor U3869 (N_3869,N_3056,N_3513);
nand U3870 (N_3870,N_3105,N_3392);
xnor U3871 (N_3871,N_3067,N_3050);
and U3872 (N_3872,N_3106,N_3528);
nand U3873 (N_3873,N_3343,N_3487);
nand U3874 (N_3874,N_3553,N_3222);
nor U3875 (N_3875,N_3128,N_3286);
or U3876 (N_3876,N_3207,N_3092);
nor U3877 (N_3877,N_3035,N_3044);
or U3878 (N_3878,N_3317,N_3042);
nand U3879 (N_3879,N_3490,N_3187);
xor U3880 (N_3880,N_3314,N_3087);
or U3881 (N_3881,N_3484,N_3039);
nand U3882 (N_3882,N_3143,N_3447);
xnor U3883 (N_3883,N_3217,N_3251);
or U3884 (N_3884,N_3102,N_3077);
nand U3885 (N_3885,N_3425,N_3327);
and U3886 (N_3886,N_3320,N_3266);
xnor U3887 (N_3887,N_3007,N_3275);
nor U3888 (N_3888,N_3239,N_3028);
xnor U3889 (N_3889,N_3350,N_3575);
or U3890 (N_3890,N_3485,N_3531);
xnor U3891 (N_3891,N_3141,N_3021);
xor U3892 (N_3892,N_3573,N_3418);
xor U3893 (N_3893,N_3179,N_3255);
nor U3894 (N_3894,N_3512,N_3107);
xor U3895 (N_3895,N_3555,N_3288);
or U3896 (N_3896,N_3282,N_3342);
nor U3897 (N_3897,N_3281,N_3333);
nor U3898 (N_3898,N_3549,N_3163);
nand U3899 (N_3899,N_3146,N_3015);
nor U3900 (N_3900,N_3417,N_3509);
nor U3901 (N_3901,N_3120,N_3086);
nand U3902 (N_3902,N_3443,N_3423);
xor U3903 (N_3903,N_3557,N_3066);
nor U3904 (N_3904,N_3308,N_3043);
or U3905 (N_3905,N_3115,N_3278);
xor U3906 (N_3906,N_3531,N_3577);
nor U3907 (N_3907,N_3328,N_3163);
xor U3908 (N_3908,N_3187,N_3457);
nand U3909 (N_3909,N_3401,N_3314);
nand U3910 (N_3910,N_3292,N_3585);
xor U3911 (N_3911,N_3247,N_3274);
xor U3912 (N_3912,N_3097,N_3370);
nand U3913 (N_3913,N_3094,N_3041);
or U3914 (N_3914,N_3372,N_3421);
and U3915 (N_3915,N_3552,N_3273);
and U3916 (N_3916,N_3077,N_3375);
or U3917 (N_3917,N_3328,N_3131);
nand U3918 (N_3918,N_3199,N_3035);
xor U3919 (N_3919,N_3261,N_3199);
and U3920 (N_3920,N_3437,N_3512);
xor U3921 (N_3921,N_3436,N_3424);
or U3922 (N_3922,N_3312,N_3098);
and U3923 (N_3923,N_3524,N_3112);
nand U3924 (N_3924,N_3202,N_3312);
xor U3925 (N_3925,N_3284,N_3384);
and U3926 (N_3926,N_3146,N_3194);
or U3927 (N_3927,N_3302,N_3084);
nand U3928 (N_3928,N_3128,N_3336);
nand U3929 (N_3929,N_3561,N_3127);
and U3930 (N_3930,N_3166,N_3427);
and U3931 (N_3931,N_3455,N_3142);
and U3932 (N_3932,N_3279,N_3544);
nand U3933 (N_3933,N_3120,N_3535);
or U3934 (N_3934,N_3436,N_3485);
nor U3935 (N_3935,N_3347,N_3432);
xor U3936 (N_3936,N_3476,N_3196);
and U3937 (N_3937,N_3218,N_3492);
nor U3938 (N_3938,N_3229,N_3167);
nor U3939 (N_3939,N_3164,N_3521);
xor U3940 (N_3940,N_3005,N_3374);
xor U3941 (N_3941,N_3459,N_3583);
xor U3942 (N_3942,N_3161,N_3367);
nand U3943 (N_3943,N_3122,N_3394);
nand U3944 (N_3944,N_3053,N_3084);
nor U3945 (N_3945,N_3421,N_3478);
or U3946 (N_3946,N_3170,N_3229);
or U3947 (N_3947,N_3226,N_3375);
nand U3948 (N_3948,N_3573,N_3569);
nor U3949 (N_3949,N_3190,N_3486);
and U3950 (N_3950,N_3501,N_3531);
nand U3951 (N_3951,N_3242,N_3591);
nor U3952 (N_3952,N_3242,N_3454);
and U3953 (N_3953,N_3265,N_3131);
and U3954 (N_3954,N_3401,N_3299);
xnor U3955 (N_3955,N_3002,N_3071);
or U3956 (N_3956,N_3560,N_3043);
and U3957 (N_3957,N_3055,N_3494);
nor U3958 (N_3958,N_3169,N_3221);
nand U3959 (N_3959,N_3250,N_3407);
or U3960 (N_3960,N_3272,N_3145);
nand U3961 (N_3961,N_3451,N_3054);
and U3962 (N_3962,N_3586,N_3293);
or U3963 (N_3963,N_3266,N_3191);
nand U3964 (N_3964,N_3030,N_3539);
and U3965 (N_3965,N_3580,N_3502);
xor U3966 (N_3966,N_3234,N_3196);
nand U3967 (N_3967,N_3253,N_3395);
xor U3968 (N_3968,N_3460,N_3560);
nand U3969 (N_3969,N_3115,N_3307);
or U3970 (N_3970,N_3594,N_3063);
xor U3971 (N_3971,N_3002,N_3081);
and U3972 (N_3972,N_3209,N_3428);
xnor U3973 (N_3973,N_3547,N_3332);
xnor U3974 (N_3974,N_3456,N_3327);
or U3975 (N_3975,N_3572,N_3420);
nor U3976 (N_3976,N_3367,N_3256);
nor U3977 (N_3977,N_3252,N_3295);
nor U3978 (N_3978,N_3201,N_3057);
xnor U3979 (N_3979,N_3078,N_3122);
xor U3980 (N_3980,N_3381,N_3339);
or U3981 (N_3981,N_3560,N_3371);
nor U3982 (N_3982,N_3266,N_3175);
or U3983 (N_3983,N_3155,N_3208);
or U3984 (N_3984,N_3470,N_3421);
nor U3985 (N_3985,N_3190,N_3053);
xor U3986 (N_3986,N_3498,N_3508);
or U3987 (N_3987,N_3369,N_3261);
xor U3988 (N_3988,N_3148,N_3272);
xor U3989 (N_3989,N_3084,N_3409);
xor U3990 (N_3990,N_3143,N_3151);
nor U3991 (N_3991,N_3205,N_3457);
nand U3992 (N_3992,N_3099,N_3298);
and U3993 (N_3993,N_3505,N_3120);
and U3994 (N_3994,N_3249,N_3206);
nor U3995 (N_3995,N_3081,N_3596);
xnor U3996 (N_3996,N_3147,N_3334);
nand U3997 (N_3997,N_3515,N_3460);
xor U3998 (N_3998,N_3269,N_3546);
nand U3999 (N_3999,N_3485,N_3433);
xor U4000 (N_4000,N_3282,N_3321);
nand U4001 (N_4001,N_3345,N_3387);
or U4002 (N_4002,N_3153,N_3348);
or U4003 (N_4003,N_3032,N_3279);
nand U4004 (N_4004,N_3304,N_3046);
xor U4005 (N_4005,N_3542,N_3297);
xnor U4006 (N_4006,N_3478,N_3312);
nor U4007 (N_4007,N_3321,N_3063);
xnor U4008 (N_4008,N_3060,N_3026);
nor U4009 (N_4009,N_3560,N_3378);
or U4010 (N_4010,N_3537,N_3455);
nor U4011 (N_4011,N_3052,N_3286);
or U4012 (N_4012,N_3452,N_3058);
or U4013 (N_4013,N_3102,N_3522);
xor U4014 (N_4014,N_3546,N_3531);
nor U4015 (N_4015,N_3064,N_3307);
nor U4016 (N_4016,N_3046,N_3160);
nand U4017 (N_4017,N_3433,N_3325);
and U4018 (N_4018,N_3437,N_3170);
or U4019 (N_4019,N_3091,N_3412);
nor U4020 (N_4020,N_3333,N_3585);
and U4021 (N_4021,N_3539,N_3226);
and U4022 (N_4022,N_3007,N_3598);
nand U4023 (N_4023,N_3266,N_3429);
or U4024 (N_4024,N_3445,N_3563);
nand U4025 (N_4025,N_3287,N_3140);
xor U4026 (N_4026,N_3446,N_3438);
nand U4027 (N_4027,N_3458,N_3380);
or U4028 (N_4028,N_3379,N_3382);
nor U4029 (N_4029,N_3403,N_3396);
xnor U4030 (N_4030,N_3458,N_3254);
or U4031 (N_4031,N_3597,N_3435);
or U4032 (N_4032,N_3202,N_3479);
and U4033 (N_4033,N_3317,N_3505);
xor U4034 (N_4034,N_3312,N_3402);
nor U4035 (N_4035,N_3594,N_3500);
xnor U4036 (N_4036,N_3464,N_3208);
and U4037 (N_4037,N_3515,N_3054);
xnor U4038 (N_4038,N_3226,N_3289);
nand U4039 (N_4039,N_3009,N_3263);
and U4040 (N_4040,N_3044,N_3338);
nand U4041 (N_4041,N_3268,N_3201);
and U4042 (N_4042,N_3226,N_3407);
xnor U4043 (N_4043,N_3437,N_3103);
nand U4044 (N_4044,N_3123,N_3103);
and U4045 (N_4045,N_3199,N_3027);
nor U4046 (N_4046,N_3273,N_3537);
nor U4047 (N_4047,N_3059,N_3413);
or U4048 (N_4048,N_3301,N_3114);
and U4049 (N_4049,N_3512,N_3483);
or U4050 (N_4050,N_3041,N_3454);
or U4051 (N_4051,N_3262,N_3564);
nand U4052 (N_4052,N_3563,N_3553);
xor U4053 (N_4053,N_3187,N_3038);
or U4054 (N_4054,N_3205,N_3035);
or U4055 (N_4055,N_3136,N_3070);
or U4056 (N_4056,N_3224,N_3069);
and U4057 (N_4057,N_3596,N_3499);
nor U4058 (N_4058,N_3225,N_3237);
nand U4059 (N_4059,N_3383,N_3589);
nand U4060 (N_4060,N_3472,N_3321);
nand U4061 (N_4061,N_3402,N_3537);
nor U4062 (N_4062,N_3243,N_3237);
or U4063 (N_4063,N_3283,N_3007);
xor U4064 (N_4064,N_3109,N_3579);
nand U4065 (N_4065,N_3049,N_3016);
xor U4066 (N_4066,N_3444,N_3075);
and U4067 (N_4067,N_3179,N_3256);
nor U4068 (N_4068,N_3085,N_3400);
or U4069 (N_4069,N_3317,N_3406);
nor U4070 (N_4070,N_3301,N_3451);
and U4071 (N_4071,N_3367,N_3239);
xnor U4072 (N_4072,N_3317,N_3192);
nand U4073 (N_4073,N_3133,N_3315);
nand U4074 (N_4074,N_3050,N_3344);
and U4075 (N_4075,N_3223,N_3309);
and U4076 (N_4076,N_3359,N_3568);
and U4077 (N_4077,N_3260,N_3522);
nand U4078 (N_4078,N_3499,N_3132);
or U4079 (N_4079,N_3491,N_3196);
xor U4080 (N_4080,N_3337,N_3308);
nand U4081 (N_4081,N_3438,N_3532);
xnor U4082 (N_4082,N_3330,N_3583);
nor U4083 (N_4083,N_3137,N_3058);
xnor U4084 (N_4084,N_3265,N_3325);
nor U4085 (N_4085,N_3249,N_3208);
xnor U4086 (N_4086,N_3199,N_3398);
nor U4087 (N_4087,N_3563,N_3236);
nand U4088 (N_4088,N_3286,N_3555);
xnor U4089 (N_4089,N_3354,N_3004);
nor U4090 (N_4090,N_3015,N_3000);
and U4091 (N_4091,N_3278,N_3149);
xor U4092 (N_4092,N_3156,N_3360);
xor U4093 (N_4093,N_3052,N_3144);
and U4094 (N_4094,N_3150,N_3145);
nor U4095 (N_4095,N_3401,N_3408);
nand U4096 (N_4096,N_3414,N_3076);
nor U4097 (N_4097,N_3094,N_3130);
and U4098 (N_4098,N_3295,N_3293);
and U4099 (N_4099,N_3216,N_3050);
and U4100 (N_4100,N_3267,N_3184);
nor U4101 (N_4101,N_3582,N_3138);
or U4102 (N_4102,N_3204,N_3261);
nand U4103 (N_4103,N_3182,N_3327);
and U4104 (N_4104,N_3081,N_3007);
or U4105 (N_4105,N_3303,N_3392);
and U4106 (N_4106,N_3334,N_3393);
or U4107 (N_4107,N_3514,N_3305);
xor U4108 (N_4108,N_3389,N_3013);
xnor U4109 (N_4109,N_3091,N_3414);
xor U4110 (N_4110,N_3570,N_3550);
and U4111 (N_4111,N_3273,N_3282);
or U4112 (N_4112,N_3088,N_3261);
nand U4113 (N_4113,N_3213,N_3406);
or U4114 (N_4114,N_3373,N_3133);
xnor U4115 (N_4115,N_3293,N_3246);
nand U4116 (N_4116,N_3304,N_3029);
nand U4117 (N_4117,N_3255,N_3076);
and U4118 (N_4118,N_3128,N_3595);
nand U4119 (N_4119,N_3243,N_3357);
and U4120 (N_4120,N_3528,N_3382);
xnor U4121 (N_4121,N_3393,N_3318);
and U4122 (N_4122,N_3239,N_3424);
nand U4123 (N_4123,N_3238,N_3043);
or U4124 (N_4124,N_3472,N_3126);
or U4125 (N_4125,N_3170,N_3118);
or U4126 (N_4126,N_3540,N_3510);
xor U4127 (N_4127,N_3572,N_3460);
nor U4128 (N_4128,N_3250,N_3360);
nor U4129 (N_4129,N_3283,N_3434);
nor U4130 (N_4130,N_3292,N_3331);
xnor U4131 (N_4131,N_3133,N_3208);
nor U4132 (N_4132,N_3251,N_3258);
and U4133 (N_4133,N_3196,N_3034);
and U4134 (N_4134,N_3405,N_3196);
and U4135 (N_4135,N_3311,N_3564);
or U4136 (N_4136,N_3542,N_3557);
or U4137 (N_4137,N_3366,N_3348);
xor U4138 (N_4138,N_3168,N_3486);
nand U4139 (N_4139,N_3422,N_3266);
nor U4140 (N_4140,N_3211,N_3537);
xor U4141 (N_4141,N_3177,N_3475);
nor U4142 (N_4142,N_3258,N_3104);
and U4143 (N_4143,N_3358,N_3466);
nand U4144 (N_4144,N_3046,N_3578);
nand U4145 (N_4145,N_3138,N_3380);
xnor U4146 (N_4146,N_3403,N_3287);
and U4147 (N_4147,N_3547,N_3367);
nor U4148 (N_4148,N_3285,N_3571);
xor U4149 (N_4149,N_3091,N_3388);
xnor U4150 (N_4150,N_3471,N_3273);
or U4151 (N_4151,N_3480,N_3252);
or U4152 (N_4152,N_3010,N_3069);
nand U4153 (N_4153,N_3068,N_3319);
and U4154 (N_4154,N_3479,N_3595);
and U4155 (N_4155,N_3218,N_3344);
nand U4156 (N_4156,N_3545,N_3131);
nor U4157 (N_4157,N_3449,N_3147);
and U4158 (N_4158,N_3048,N_3363);
and U4159 (N_4159,N_3198,N_3520);
xor U4160 (N_4160,N_3116,N_3200);
nor U4161 (N_4161,N_3521,N_3575);
nand U4162 (N_4162,N_3351,N_3349);
nor U4163 (N_4163,N_3457,N_3209);
or U4164 (N_4164,N_3075,N_3429);
or U4165 (N_4165,N_3084,N_3016);
or U4166 (N_4166,N_3034,N_3435);
and U4167 (N_4167,N_3490,N_3499);
or U4168 (N_4168,N_3431,N_3158);
xnor U4169 (N_4169,N_3150,N_3023);
xor U4170 (N_4170,N_3229,N_3356);
or U4171 (N_4171,N_3539,N_3437);
and U4172 (N_4172,N_3156,N_3578);
nand U4173 (N_4173,N_3135,N_3496);
nand U4174 (N_4174,N_3211,N_3171);
and U4175 (N_4175,N_3237,N_3041);
nor U4176 (N_4176,N_3512,N_3480);
or U4177 (N_4177,N_3095,N_3395);
or U4178 (N_4178,N_3475,N_3541);
xor U4179 (N_4179,N_3525,N_3557);
nor U4180 (N_4180,N_3407,N_3146);
or U4181 (N_4181,N_3335,N_3336);
or U4182 (N_4182,N_3546,N_3398);
and U4183 (N_4183,N_3439,N_3350);
and U4184 (N_4184,N_3547,N_3128);
or U4185 (N_4185,N_3555,N_3598);
nor U4186 (N_4186,N_3373,N_3357);
nand U4187 (N_4187,N_3271,N_3218);
nand U4188 (N_4188,N_3522,N_3439);
nand U4189 (N_4189,N_3488,N_3456);
xnor U4190 (N_4190,N_3052,N_3174);
or U4191 (N_4191,N_3174,N_3209);
nand U4192 (N_4192,N_3535,N_3500);
nand U4193 (N_4193,N_3322,N_3442);
and U4194 (N_4194,N_3462,N_3513);
xnor U4195 (N_4195,N_3448,N_3516);
or U4196 (N_4196,N_3440,N_3230);
and U4197 (N_4197,N_3189,N_3404);
and U4198 (N_4198,N_3117,N_3070);
and U4199 (N_4199,N_3466,N_3442);
and U4200 (N_4200,N_3711,N_4042);
nor U4201 (N_4201,N_4020,N_3852);
xor U4202 (N_4202,N_4064,N_3961);
nand U4203 (N_4203,N_3949,N_3725);
or U4204 (N_4204,N_3873,N_3703);
xor U4205 (N_4205,N_4045,N_3997);
nor U4206 (N_4206,N_3792,N_3821);
nor U4207 (N_4207,N_3657,N_4044);
and U4208 (N_4208,N_3698,N_3655);
xor U4209 (N_4209,N_3764,N_4016);
nand U4210 (N_4210,N_3660,N_3983);
xor U4211 (N_4211,N_3752,N_3883);
nor U4212 (N_4212,N_3683,N_3771);
or U4213 (N_4213,N_3663,N_3741);
xor U4214 (N_4214,N_4123,N_3819);
nand U4215 (N_4215,N_3673,N_4147);
xnor U4216 (N_4216,N_4056,N_3775);
nand U4217 (N_4217,N_3788,N_3796);
or U4218 (N_4218,N_3602,N_3837);
or U4219 (N_4219,N_3692,N_4178);
xor U4220 (N_4220,N_4017,N_3789);
xnor U4221 (N_4221,N_4050,N_3760);
nor U4222 (N_4222,N_4192,N_4019);
xnor U4223 (N_4223,N_4115,N_3665);
nor U4224 (N_4224,N_3649,N_3936);
or U4225 (N_4225,N_3981,N_3704);
xnor U4226 (N_4226,N_3661,N_3705);
nor U4227 (N_4227,N_4104,N_3800);
nand U4228 (N_4228,N_4150,N_3613);
or U4229 (N_4229,N_3892,N_3757);
xor U4230 (N_4230,N_4021,N_3847);
xnor U4231 (N_4231,N_3749,N_3957);
nor U4232 (N_4232,N_3753,N_3923);
nand U4233 (N_4233,N_3820,N_3674);
and U4234 (N_4234,N_4060,N_3933);
nand U4235 (N_4235,N_3601,N_3992);
nand U4236 (N_4236,N_3710,N_4069);
nand U4237 (N_4237,N_3851,N_4040);
or U4238 (N_4238,N_3776,N_3728);
and U4239 (N_4239,N_3912,N_3893);
and U4240 (N_4240,N_3624,N_3989);
nor U4241 (N_4241,N_3790,N_3805);
nor U4242 (N_4242,N_3785,N_3614);
xor U4243 (N_4243,N_3914,N_3802);
nor U4244 (N_4244,N_4151,N_4059);
or U4245 (N_4245,N_3921,N_4096);
or U4246 (N_4246,N_3600,N_3818);
nor U4247 (N_4247,N_4043,N_3736);
and U4248 (N_4248,N_3784,N_3787);
xor U4249 (N_4249,N_4125,N_3621);
nor U4250 (N_4250,N_3849,N_3814);
xor U4251 (N_4251,N_3694,N_3833);
and U4252 (N_4252,N_4072,N_3908);
or U4253 (N_4253,N_3695,N_3778);
and U4254 (N_4254,N_3666,N_4141);
and U4255 (N_4255,N_4006,N_3877);
and U4256 (N_4256,N_4095,N_3606);
or U4257 (N_4257,N_3740,N_3935);
nor U4258 (N_4258,N_4098,N_3843);
nor U4259 (N_4259,N_3795,N_3638);
nand U4260 (N_4260,N_4127,N_3697);
xor U4261 (N_4261,N_3756,N_3642);
xnor U4262 (N_4262,N_4008,N_3662);
nor U4263 (N_4263,N_3720,N_3995);
or U4264 (N_4264,N_4145,N_4120);
or U4265 (N_4265,N_3941,N_4077);
or U4266 (N_4266,N_3920,N_4185);
nand U4267 (N_4267,N_3617,N_4167);
or U4268 (N_4268,N_4011,N_3744);
nand U4269 (N_4269,N_4058,N_4085);
nor U4270 (N_4270,N_3632,N_3682);
and U4271 (N_4271,N_3654,N_4015);
or U4272 (N_4272,N_4074,N_3659);
and U4273 (N_4273,N_4087,N_4129);
nor U4274 (N_4274,N_3605,N_3706);
or U4275 (N_4275,N_4100,N_4156);
nand U4276 (N_4276,N_4162,N_4140);
or U4277 (N_4277,N_3607,N_3629);
nor U4278 (N_4278,N_3636,N_3643);
or U4279 (N_4279,N_3906,N_4121);
xor U4280 (N_4280,N_3754,N_4119);
nand U4281 (N_4281,N_4078,N_3747);
nor U4282 (N_4282,N_3731,N_3766);
nand U4283 (N_4283,N_3804,N_3715);
or U4284 (N_4284,N_4184,N_4190);
nand U4285 (N_4285,N_3664,N_3631);
nand U4286 (N_4286,N_3887,N_4089);
nor U4287 (N_4287,N_3960,N_3729);
nor U4288 (N_4288,N_3721,N_3679);
and U4289 (N_4289,N_4028,N_3990);
or U4290 (N_4290,N_4038,N_3954);
nor U4291 (N_4291,N_4024,N_4079);
and U4292 (N_4292,N_3658,N_3878);
and U4293 (N_4293,N_4143,N_3689);
or U4294 (N_4294,N_4102,N_3816);
or U4295 (N_4295,N_3611,N_3862);
nand U4296 (N_4296,N_3861,N_3942);
nor U4297 (N_4297,N_4065,N_3651);
and U4298 (N_4298,N_3952,N_3925);
and U4299 (N_4299,N_3890,N_4084);
xor U4300 (N_4300,N_3964,N_3737);
and U4301 (N_4301,N_4128,N_3670);
nor U4302 (N_4302,N_4114,N_3948);
and U4303 (N_4303,N_4073,N_4090);
and U4304 (N_4304,N_3966,N_3889);
nor U4305 (N_4305,N_3916,N_4035);
or U4306 (N_4306,N_3653,N_3722);
nand U4307 (N_4307,N_3848,N_3962);
and U4308 (N_4308,N_3931,N_3973);
nand U4309 (N_4309,N_4000,N_4148);
nand U4310 (N_4310,N_3869,N_4003);
or U4311 (N_4311,N_4166,N_4130);
xnor U4312 (N_4312,N_3884,N_3678);
xor U4313 (N_4313,N_4110,N_3770);
or U4314 (N_4314,N_3668,N_3841);
nand U4315 (N_4315,N_4014,N_3812);
or U4316 (N_4316,N_3856,N_3610);
xor U4317 (N_4317,N_3732,N_3797);
nor U4318 (N_4318,N_3693,N_3699);
nor U4319 (N_4319,N_3686,N_4194);
nor U4320 (N_4320,N_3768,N_3707);
nor U4321 (N_4321,N_3926,N_3615);
nor U4322 (N_4322,N_4152,N_3874);
xnor U4323 (N_4323,N_4107,N_3772);
or U4324 (N_4324,N_4149,N_4196);
nand U4325 (N_4325,N_3898,N_3751);
nand U4326 (N_4326,N_4174,N_3999);
xor U4327 (N_4327,N_3619,N_4132);
or U4328 (N_4328,N_4076,N_3635);
and U4329 (N_4329,N_3652,N_4183);
nand U4330 (N_4330,N_4198,N_3761);
or U4331 (N_4331,N_3738,N_4004);
or U4332 (N_4332,N_4091,N_3876);
xor U4333 (N_4333,N_3813,N_3958);
xor U4334 (N_4334,N_3627,N_3680);
and U4335 (N_4335,N_4188,N_3781);
or U4336 (N_4336,N_3971,N_3904);
nor U4337 (N_4337,N_3899,N_4010);
nor U4338 (N_4338,N_4112,N_3701);
xnor U4339 (N_4339,N_3894,N_3886);
nand U4340 (N_4340,N_4159,N_3854);
or U4341 (N_4341,N_3640,N_3690);
nand U4342 (N_4342,N_3903,N_3969);
xnor U4343 (N_4343,N_4146,N_3970);
nor U4344 (N_4344,N_3647,N_3972);
or U4345 (N_4345,N_3824,N_3986);
and U4346 (N_4346,N_3672,N_4142);
nand U4347 (N_4347,N_4134,N_4086);
and U4348 (N_4348,N_3864,N_3859);
or U4349 (N_4349,N_3719,N_3924);
nor U4350 (N_4350,N_4182,N_4082);
nand U4351 (N_4351,N_4081,N_3700);
xor U4352 (N_4352,N_3675,N_3860);
and U4353 (N_4353,N_3763,N_3947);
or U4354 (N_4354,N_3681,N_3801);
xnor U4355 (N_4355,N_4111,N_4037);
xnor U4356 (N_4356,N_4018,N_4007);
nor U4357 (N_4357,N_3743,N_4113);
xor U4358 (N_4358,N_4048,N_3733);
nor U4359 (N_4359,N_3810,N_3677);
nand U4360 (N_4360,N_3730,N_4136);
or U4361 (N_4361,N_4034,N_3950);
nand U4362 (N_4362,N_4153,N_3855);
nor U4363 (N_4363,N_3857,N_4195);
and U4364 (N_4364,N_3782,N_3807);
nand U4365 (N_4365,N_4181,N_3965);
and U4366 (N_4366,N_3832,N_4173);
and U4367 (N_4367,N_4108,N_4179);
nor U4368 (N_4368,N_4168,N_3793);
xor U4369 (N_4369,N_3691,N_3838);
xnor U4370 (N_4370,N_3939,N_3932);
nor U4371 (N_4371,N_3900,N_3646);
nor U4372 (N_4372,N_3979,N_4116);
nand U4373 (N_4373,N_4067,N_3853);
nor U4374 (N_4374,N_3687,N_3863);
or U4375 (N_4375,N_4169,N_3718);
xor U4376 (N_4376,N_3896,N_3656);
nand U4377 (N_4377,N_4180,N_3727);
xor U4378 (N_4378,N_3987,N_3917);
xnor U4379 (N_4379,N_4062,N_3604);
nand U4380 (N_4380,N_3623,N_3823);
nor U4381 (N_4381,N_3955,N_3844);
nand U4382 (N_4382,N_3645,N_4131);
or U4383 (N_4383,N_4002,N_3735);
nand U4384 (N_4384,N_4118,N_4103);
and U4385 (N_4385,N_3734,N_3723);
xnor U4386 (N_4386,N_3967,N_4063);
and U4387 (N_4387,N_4071,N_4061);
or U4388 (N_4388,N_4177,N_4083);
or U4389 (N_4389,N_4070,N_3993);
or U4390 (N_4390,N_3938,N_3842);
nand U4391 (N_4391,N_3834,N_3830);
xor U4392 (N_4392,N_3786,N_3836);
or U4393 (N_4393,N_3959,N_4158);
nor U4394 (N_4394,N_3907,N_3928);
nor U4395 (N_4395,N_4036,N_3829);
or U4396 (N_4396,N_3835,N_3676);
nand U4397 (N_4397,N_3745,N_3976);
nor U4398 (N_4398,N_3991,N_3822);
or U4399 (N_4399,N_3905,N_3762);
or U4400 (N_4400,N_4097,N_3750);
nand U4401 (N_4401,N_4139,N_4001);
and U4402 (N_4402,N_3902,N_3978);
xor U4403 (N_4403,N_4068,N_4005);
xor U4404 (N_4404,N_3620,N_3910);
xnor U4405 (N_4405,N_4175,N_3980);
xnor U4406 (N_4406,N_3875,N_3669);
and U4407 (N_4407,N_3911,N_3944);
and U4408 (N_4408,N_4033,N_4088);
xor U4409 (N_4409,N_3612,N_4094);
and U4410 (N_4410,N_4049,N_3616);
nand U4411 (N_4411,N_3934,N_4054);
and U4412 (N_4412,N_4199,N_3891);
nand U4413 (N_4413,N_3783,N_4046);
or U4414 (N_4414,N_3865,N_3609);
nor U4415 (N_4415,N_3702,N_3885);
and U4416 (N_4416,N_3953,N_3739);
xnor U4417 (N_4417,N_4161,N_3811);
or U4418 (N_4418,N_3714,N_3839);
and U4419 (N_4419,N_3872,N_3858);
nand U4420 (N_4420,N_4124,N_3994);
xor U4421 (N_4421,N_3827,N_4026);
xor U4422 (N_4422,N_3746,N_4176);
xor U4423 (N_4423,N_3968,N_3650);
nor U4424 (N_4424,N_4075,N_3634);
xnor U4425 (N_4425,N_3633,N_3828);
xnor U4426 (N_4426,N_3696,N_4165);
xnor U4427 (N_4427,N_3671,N_4157);
nand U4428 (N_4428,N_3626,N_3882);
or U4429 (N_4429,N_3982,N_3825);
xor U4430 (N_4430,N_4154,N_4027);
and U4431 (N_4431,N_3826,N_3798);
xnor U4432 (N_4432,N_4171,N_3806);
and U4433 (N_4433,N_3791,N_3867);
and U4434 (N_4434,N_3881,N_4093);
nor U4435 (N_4435,N_3773,N_3913);
xor U4436 (N_4436,N_3915,N_3644);
xor U4437 (N_4437,N_3943,N_4051);
and U4438 (N_4438,N_3769,N_4197);
xor U4439 (N_4439,N_4032,N_3708);
nand U4440 (N_4440,N_3625,N_4155);
nor U4441 (N_4441,N_3779,N_3716);
and U4442 (N_4442,N_4193,N_3850);
and U4443 (N_4443,N_3685,N_4187);
nor U4444 (N_4444,N_4066,N_3755);
or U4445 (N_4445,N_4029,N_3963);
nand U4446 (N_4446,N_3603,N_4164);
and U4447 (N_4447,N_3777,N_3622);
nand U4448 (N_4448,N_3975,N_4106);
and U4449 (N_4449,N_4039,N_3871);
nor U4450 (N_4450,N_3929,N_3759);
xnor U4451 (N_4451,N_4137,N_3717);
and U4452 (N_4452,N_3919,N_4138);
or U4453 (N_4453,N_3951,N_3840);
and U4454 (N_4454,N_3726,N_3767);
nor U4455 (N_4455,N_3713,N_3808);
and U4456 (N_4456,N_4117,N_3809);
nor U4457 (N_4457,N_4009,N_4189);
or U4458 (N_4458,N_3868,N_4170);
nor U4459 (N_4459,N_3984,N_3774);
nand U4460 (N_4460,N_3940,N_4105);
and U4461 (N_4461,N_3977,N_3815);
nor U4462 (N_4462,N_4186,N_3918);
nand U4463 (N_4463,N_4052,N_3895);
or U4464 (N_4464,N_3996,N_3641);
nand U4465 (N_4465,N_4191,N_3927);
xnor U4466 (N_4466,N_3803,N_3937);
nor U4467 (N_4467,N_3985,N_4013);
or U4468 (N_4468,N_4031,N_3780);
or U4469 (N_4469,N_4144,N_3748);
nor U4470 (N_4470,N_3724,N_4025);
nand U4471 (N_4471,N_3930,N_4133);
nor U4472 (N_4472,N_3988,N_3922);
and U4473 (N_4473,N_3712,N_3879);
and U4474 (N_4474,N_4135,N_3870);
xnor U4475 (N_4475,N_4126,N_3888);
or U4476 (N_4476,N_3846,N_3765);
or U4477 (N_4477,N_4022,N_4057);
or U4478 (N_4478,N_3608,N_4030);
and U4479 (N_4479,N_3956,N_4012);
nand U4480 (N_4480,N_3639,N_3742);
or U4481 (N_4481,N_3974,N_4160);
xnor U4482 (N_4482,N_3909,N_4055);
nor U4483 (N_4483,N_3667,N_3758);
and U4484 (N_4484,N_4092,N_3880);
nor U4485 (N_4485,N_3901,N_3945);
or U4486 (N_4486,N_3831,N_4041);
nor U4487 (N_4487,N_3817,N_3866);
xnor U4488 (N_4488,N_3897,N_3630);
nor U4489 (N_4489,N_4122,N_4053);
nand U4490 (N_4490,N_3794,N_4023);
nor U4491 (N_4491,N_4109,N_4101);
or U4492 (N_4492,N_4047,N_3628);
nand U4493 (N_4493,N_4163,N_3618);
and U4494 (N_4494,N_3799,N_4099);
or U4495 (N_4495,N_3709,N_4080);
and U4496 (N_4496,N_3648,N_3684);
or U4497 (N_4497,N_3998,N_3946);
xnor U4498 (N_4498,N_3845,N_3688);
and U4499 (N_4499,N_4172,N_3637);
nor U4500 (N_4500,N_3610,N_3694);
and U4501 (N_4501,N_4155,N_3707);
nand U4502 (N_4502,N_3723,N_3787);
or U4503 (N_4503,N_3988,N_4069);
and U4504 (N_4504,N_3769,N_4136);
nor U4505 (N_4505,N_3804,N_4068);
or U4506 (N_4506,N_3766,N_3643);
and U4507 (N_4507,N_4034,N_3903);
or U4508 (N_4508,N_4046,N_3674);
xnor U4509 (N_4509,N_3886,N_3710);
and U4510 (N_4510,N_3833,N_3969);
xor U4511 (N_4511,N_3698,N_4004);
or U4512 (N_4512,N_3920,N_3874);
or U4513 (N_4513,N_3785,N_3752);
and U4514 (N_4514,N_3681,N_3750);
xor U4515 (N_4515,N_4025,N_4026);
and U4516 (N_4516,N_3861,N_4087);
nand U4517 (N_4517,N_3978,N_4075);
and U4518 (N_4518,N_3991,N_4040);
or U4519 (N_4519,N_3734,N_3993);
or U4520 (N_4520,N_3651,N_4136);
and U4521 (N_4521,N_3958,N_3940);
nand U4522 (N_4522,N_3793,N_4087);
nor U4523 (N_4523,N_3698,N_4023);
nand U4524 (N_4524,N_3880,N_4160);
xnor U4525 (N_4525,N_4034,N_3897);
or U4526 (N_4526,N_4096,N_4152);
or U4527 (N_4527,N_3615,N_3679);
nor U4528 (N_4528,N_4171,N_4015);
and U4529 (N_4529,N_3722,N_3947);
nand U4530 (N_4530,N_3889,N_3702);
or U4531 (N_4531,N_4073,N_4105);
xor U4532 (N_4532,N_3800,N_3855);
nor U4533 (N_4533,N_4087,N_4077);
nand U4534 (N_4534,N_3885,N_3973);
nor U4535 (N_4535,N_4110,N_3753);
or U4536 (N_4536,N_3623,N_4116);
or U4537 (N_4537,N_4082,N_3679);
xor U4538 (N_4538,N_3802,N_3942);
and U4539 (N_4539,N_4128,N_3647);
nand U4540 (N_4540,N_3881,N_4150);
nand U4541 (N_4541,N_3918,N_4138);
or U4542 (N_4542,N_4184,N_4047);
nand U4543 (N_4543,N_3884,N_3807);
nand U4544 (N_4544,N_3843,N_3795);
nor U4545 (N_4545,N_3966,N_4012);
nor U4546 (N_4546,N_3607,N_3798);
or U4547 (N_4547,N_3746,N_3790);
xnor U4548 (N_4548,N_3935,N_3908);
xnor U4549 (N_4549,N_3793,N_3835);
xor U4550 (N_4550,N_3985,N_3753);
and U4551 (N_4551,N_4044,N_3917);
nand U4552 (N_4552,N_3658,N_3837);
xor U4553 (N_4553,N_3985,N_4137);
or U4554 (N_4554,N_3991,N_4019);
nand U4555 (N_4555,N_3703,N_4187);
and U4556 (N_4556,N_3775,N_4064);
nand U4557 (N_4557,N_4184,N_4123);
xor U4558 (N_4558,N_3984,N_3781);
nor U4559 (N_4559,N_3959,N_3770);
and U4560 (N_4560,N_4064,N_3989);
or U4561 (N_4561,N_4067,N_3933);
nand U4562 (N_4562,N_3956,N_4096);
xnor U4563 (N_4563,N_4081,N_3724);
xnor U4564 (N_4564,N_3853,N_4014);
nand U4565 (N_4565,N_3740,N_3967);
xor U4566 (N_4566,N_3845,N_4143);
xnor U4567 (N_4567,N_3773,N_3783);
nor U4568 (N_4568,N_4076,N_4159);
xnor U4569 (N_4569,N_4014,N_3731);
or U4570 (N_4570,N_3784,N_3704);
and U4571 (N_4571,N_3690,N_4043);
nand U4572 (N_4572,N_3915,N_4039);
nor U4573 (N_4573,N_3883,N_4132);
nor U4574 (N_4574,N_4136,N_4073);
xnor U4575 (N_4575,N_4164,N_4137);
nor U4576 (N_4576,N_4011,N_4167);
xnor U4577 (N_4577,N_4098,N_3624);
and U4578 (N_4578,N_3915,N_4073);
and U4579 (N_4579,N_3663,N_4140);
nand U4580 (N_4580,N_3899,N_3802);
or U4581 (N_4581,N_3810,N_3852);
and U4582 (N_4582,N_3805,N_4104);
and U4583 (N_4583,N_3783,N_4178);
or U4584 (N_4584,N_3802,N_3931);
and U4585 (N_4585,N_4036,N_3747);
nand U4586 (N_4586,N_3620,N_4018);
and U4587 (N_4587,N_4054,N_3618);
and U4588 (N_4588,N_3622,N_3761);
and U4589 (N_4589,N_4127,N_3716);
nand U4590 (N_4590,N_4004,N_3761);
nor U4591 (N_4591,N_3820,N_3654);
and U4592 (N_4592,N_4113,N_3917);
or U4593 (N_4593,N_4079,N_4174);
nand U4594 (N_4594,N_3694,N_3989);
nand U4595 (N_4595,N_3672,N_3668);
nor U4596 (N_4596,N_4053,N_3920);
and U4597 (N_4597,N_3682,N_4104);
nand U4598 (N_4598,N_3852,N_3647);
and U4599 (N_4599,N_4199,N_4185);
nor U4600 (N_4600,N_3624,N_4003);
and U4601 (N_4601,N_3671,N_3953);
nor U4602 (N_4602,N_3893,N_4140);
nand U4603 (N_4603,N_3926,N_3694);
or U4604 (N_4604,N_3868,N_3761);
and U4605 (N_4605,N_3730,N_4050);
nand U4606 (N_4606,N_3616,N_4073);
xor U4607 (N_4607,N_3925,N_4036);
nand U4608 (N_4608,N_4134,N_3948);
xnor U4609 (N_4609,N_3976,N_4099);
and U4610 (N_4610,N_4009,N_3662);
nand U4611 (N_4611,N_3819,N_4043);
nor U4612 (N_4612,N_4119,N_4158);
nor U4613 (N_4613,N_3942,N_3800);
or U4614 (N_4614,N_3613,N_4049);
nand U4615 (N_4615,N_4062,N_3735);
nor U4616 (N_4616,N_4127,N_3642);
nand U4617 (N_4617,N_3820,N_3677);
nor U4618 (N_4618,N_3907,N_3639);
and U4619 (N_4619,N_4026,N_3972);
or U4620 (N_4620,N_3807,N_3957);
nand U4621 (N_4621,N_3891,N_3602);
nor U4622 (N_4622,N_3812,N_3804);
nand U4623 (N_4623,N_4146,N_4105);
or U4624 (N_4624,N_3984,N_3760);
nand U4625 (N_4625,N_4064,N_3829);
or U4626 (N_4626,N_4137,N_3866);
nand U4627 (N_4627,N_4166,N_3975);
nand U4628 (N_4628,N_3980,N_3975);
xor U4629 (N_4629,N_3696,N_3815);
and U4630 (N_4630,N_4023,N_3898);
nand U4631 (N_4631,N_3718,N_3875);
nor U4632 (N_4632,N_3733,N_3649);
or U4633 (N_4633,N_4121,N_4150);
xnor U4634 (N_4634,N_3679,N_3687);
xor U4635 (N_4635,N_4167,N_3683);
nand U4636 (N_4636,N_3886,N_3878);
or U4637 (N_4637,N_3902,N_3695);
and U4638 (N_4638,N_3657,N_3638);
or U4639 (N_4639,N_4155,N_3961);
and U4640 (N_4640,N_4096,N_3627);
nor U4641 (N_4641,N_3861,N_3611);
nor U4642 (N_4642,N_4152,N_3899);
or U4643 (N_4643,N_3811,N_3943);
and U4644 (N_4644,N_4024,N_3888);
xor U4645 (N_4645,N_3801,N_4120);
nand U4646 (N_4646,N_3695,N_4083);
nand U4647 (N_4647,N_3801,N_4035);
nor U4648 (N_4648,N_3708,N_3759);
or U4649 (N_4649,N_4190,N_4115);
nand U4650 (N_4650,N_4026,N_4182);
xnor U4651 (N_4651,N_4188,N_3631);
and U4652 (N_4652,N_3834,N_4196);
xor U4653 (N_4653,N_3610,N_3699);
nor U4654 (N_4654,N_3856,N_3785);
nand U4655 (N_4655,N_3930,N_4142);
and U4656 (N_4656,N_3827,N_4196);
xnor U4657 (N_4657,N_4096,N_4139);
nor U4658 (N_4658,N_3977,N_4146);
xor U4659 (N_4659,N_4020,N_4000);
nand U4660 (N_4660,N_3851,N_3909);
and U4661 (N_4661,N_3947,N_3997);
nor U4662 (N_4662,N_3955,N_3899);
or U4663 (N_4663,N_3960,N_3850);
or U4664 (N_4664,N_4119,N_3846);
or U4665 (N_4665,N_4044,N_3606);
nor U4666 (N_4666,N_3982,N_3756);
nand U4667 (N_4667,N_4182,N_3748);
nand U4668 (N_4668,N_3658,N_3739);
nand U4669 (N_4669,N_3778,N_3697);
and U4670 (N_4670,N_3827,N_4101);
nor U4671 (N_4671,N_3988,N_4094);
and U4672 (N_4672,N_3713,N_3730);
or U4673 (N_4673,N_3812,N_3772);
and U4674 (N_4674,N_4189,N_3650);
and U4675 (N_4675,N_3848,N_4092);
and U4676 (N_4676,N_3731,N_4159);
nand U4677 (N_4677,N_3630,N_3870);
nor U4678 (N_4678,N_3686,N_3687);
xor U4679 (N_4679,N_3609,N_3868);
xor U4680 (N_4680,N_3923,N_4099);
nor U4681 (N_4681,N_3726,N_4066);
xor U4682 (N_4682,N_3875,N_3762);
or U4683 (N_4683,N_4011,N_4188);
nand U4684 (N_4684,N_4160,N_3875);
and U4685 (N_4685,N_3864,N_4185);
or U4686 (N_4686,N_4193,N_3732);
nor U4687 (N_4687,N_3997,N_4162);
and U4688 (N_4688,N_3602,N_4050);
or U4689 (N_4689,N_3958,N_3816);
and U4690 (N_4690,N_4163,N_4161);
nand U4691 (N_4691,N_3699,N_3620);
and U4692 (N_4692,N_3949,N_3662);
and U4693 (N_4693,N_4013,N_3622);
nand U4694 (N_4694,N_3929,N_3900);
nand U4695 (N_4695,N_4079,N_4120);
nand U4696 (N_4696,N_3885,N_4151);
or U4697 (N_4697,N_3894,N_3915);
nand U4698 (N_4698,N_3979,N_4113);
or U4699 (N_4699,N_3885,N_3977);
nor U4700 (N_4700,N_3664,N_3875);
xnor U4701 (N_4701,N_4142,N_3694);
nor U4702 (N_4702,N_4054,N_3974);
or U4703 (N_4703,N_4158,N_3718);
xnor U4704 (N_4704,N_3626,N_4025);
and U4705 (N_4705,N_4179,N_4190);
nor U4706 (N_4706,N_4174,N_4074);
and U4707 (N_4707,N_3827,N_4181);
xor U4708 (N_4708,N_4191,N_4046);
xor U4709 (N_4709,N_3625,N_3643);
nand U4710 (N_4710,N_4076,N_3995);
xor U4711 (N_4711,N_4177,N_3972);
nor U4712 (N_4712,N_3942,N_4027);
nand U4713 (N_4713,N_4196,N_4111);
nand U4714 (N_4714,N_3893,N_3935);
nor U4715 (N_4715,N_4101,N_4015);
xnor U4716 (N_4716,N_4199,N_4132);
nor U4717 (N_4717,N_3863,N_4055);
and U4718 (N_4718,N_4005,N_4198);
or U4719 (N_4719,N_3867,N_3655);
nand U4720 (N_4720,N_3904,N_4012);
or U4721 (N_4721,N_3964,N_3715);
nand U4722 (N_4722,N_3656,N_3678);
nand U4723 (N_4723,N_3748,N_3675);
or U4724 (N_4724,N_4088,N_3845);
xor U4725 (N_4725,N_4098,N_3916);
nand U4726 (N_4726,N_3869,N_3753);
or U4727 (N_4727,N_3688,N_3664);
or U4728 (N_4728,N_4120,N_3788);
nand U4729 (N_4729,N_4150,N_3936);
xor U4730 (N_4730,N_3799,N_3902);
xnor U4731 (N_4731,N_3859,N_3969);
nand U4732 (N_4732,N_4066,N_3781);
and U4733 (N_4733,N_3972,N_3732);
xor U4734 (N_4734,N_4118,N_3908);
nor U4735 (N_4735,N_3691,N_4056);
or U4736 (N_4736,N_3862,N_3765);
nor U4737 (N_4737,N_3677,N_4185);
xor U4738 (N_4738,N_4062,N_3762);
and U4739 (N_4739,N_4097,N_3959);
nand U4740 (N_4740,N_4029,N_3757);
or U4741 (N_4741,N_3790,N_3696);
nand U4742 (N_4742,N_3630,N_3830);
nand U4743 (N_4743,N_3857,N_3912);
and U4744 (N_4744,N_4092,N_4179);
or U4745 (N_4745,N_4068,N_3899);
and U4746 (N_4746,N_4105,N_3759);
and U4747 (N_4747,N_3742,N_4138);
xor U4748 (N_4748,N_4005,N_4007);
or U4749 (N_4749,N_4061,N_4182);
nor U4750 (N_4750,N_3726,N_4035);
nor U4751 (N_4751,N_4016,N_3772);
nand U4752 (N_4752,N_3891,N_3658);
nand U4753 (N_4753,N_3893,N_3864);
xor U4754 (N_4754,N_4042,N_4005);
nor U4755 (N_4755,N_3880,N_3754);
nor U4756 (N_4756,N_3692,N_3742);
nor U4757 (N_4757,N_4044,N_3888);
xnor U4758 (N_4758,N_3806,N_3679);
nor U4759 (N_4759,N_3896,N_4000);
and U4760 (N_4760,N_3864,N_3655);
nor U4761 (N_4761,N_3837,N_4082);
nor U4762 (N_4762,N_3666,N_3674);
and U4763 (N_4763,N_3752,N_3903);
nand U4764 (N_4764,N_3740,N_3930);
or U4765 (N_4765,N_3968,N_3673);
or U4766 (N_4766,N_4106,N_3957);
or U4767 (N_4767,N_3616,N_4083);
or U4768 (N_4768,N_4145,N_4105);
and U4769 (N_4769,N_4040,N_4066);
or U4770 (N_4770,N_3855,N_4159);
xor U4771 (N_4771,N_3664,N_3662);
xnor U4772 (N_4772,N_3860,N_4089);
and U4773 (N_4773,N_3772,N_3824);
or U4774 (N_4774,N_3911,N_3752);
nand U4775 (N_4775,N_4104,N_4187);
or U4776 (N_4776,N_3960,N_4053);
and U4777 (N_4777,N_3764,N_3883);
or U4778 (N_4778,N_3627,N_3850);
nor U4779 (N_4779,N_4031,N_4118);
nand U4780 (N_4780,N_3977,N_3666);
nand U4781 (N_4781,N_3804,N_3907);
nor U4782 (N_4782,N_3704,N_3925);
nor U4783 (N_4783,N_4043,N_3862);
or U4784 (N_4784,N_3882,N_4096);
nor U4785 (N_4785,N_4165,N_3920);
or U4786 (N_4786,N_3827,N_4068);
or U4787 (N_4787,N_3633,N_4008);
or U4788 (N_4788,N_4094,N_4078);
and U4789 (N_4789,N_3913,N_4032);
nor U4790 (N_4790,N_4121,N_3769);
nor U4791 (N_4791,N_4195,N_3803);
nor U4792 (N_4792,N_4150,N_3982);
nand U4793 (N_4793,N_4199,N_4139);
or U4794 (N_4794,N_3772,N_4014);
nand U4795 (N_4795,N_4145,N_3881);
and U4796 (N_4796,N_3681,N_4185);
nor U4797 (N_4797,N_3909,N_3616);
or U4798 (N_4798,N_3743,N_4021);
nand U4799 (N_4799,N_3990,N_3784);
or U4800 (N_4800,N_4726,N_4289);
or U4801 (N_4801,N_4234,N_4264);
nor U4802 (N_4802,N_4374,N_4243);
nor U4803 (N_4803,N_4200,N_4716);
and U4804 (N_4804,N_4571,N_4325);
nand U4805 (N_4805,N_4398,N_4501);
nand U4806 (N_4806,N_4293,N_4504);
or U4807 (N_4807,N_4259,N_4590);
nand U4808 (N_4808,N_4321,N_4759);
nand U4809 (N_4809,N_4793,N_4579);
or U4810 (N_4810,N_4225,N_4328);
nor U4811 (N_4811,N_4787,N_4622);
xnor U4812 (N_4812,N_4657,N_4639);
or U4813 (N_4813,N_4449,N_4311);
xor U4814 (N_4814,N_4732,N_4468);
and U4815 (N_4815,N_4296,N_4313);
nand U4816 (N_4816,N_4209,N_4424);
and U4817 (N_4817,N_4361,N_4530);
and U4818 (N_4818,N_4621,N_4618);
xor U4819 (N_4819,N_4485,N_4436);
and U4820 (N_4820,N_4244,N_4546);
nand U4821 (N_4821,N_4344,N_4735);
xnor U4822 (N_4822,N_4399,N_4454);
xor U4823 (N_4823,N_4228,N_4393);
nor U4824 (N_4824,N_4332,N_4747);
xor U4825 (N_4825,N_4533,N_4473);
and U4826 (N_4826,N_4655,N_4300);
nand U4827 (N_4827,N_4592,N_4547);
xor U4828 (N_4828,N_4373,N_4308);
or U4829 (N_4829,N_4681,N_4691);
nand U4830 (N_4830,N_4320,N_4771);
xnor U4831 (N_4831,N_4617,N_4528);
and U4832 (N_4832,N_4426,N_4438);
nand U4833 (N_4833,N_4260,N_4394);
nand U4834 (N_4834,N_4381,N_4347);
nor U4835 (N_4835,N_4380,N_4428);
or U4836 (N_4836,N_4589,N_4695);
xnor U4837 (N_4837,N_4582,N_4684);
xor U4838 (N_4838,N_4378,N_4524);
and U4839 (N_4839,N_4369,N_4372);
and U4840 (N_4840,N_4465,N_4673);
or U4841 (N_4841,N_4627,N_4511);
nor U4842 (N_4842,N_4593,N_4569);
and U4843 (N_4843,N_4461,N_4672);
and U4844 (N_4844,N_4407,N_4435);
and U4845 (N_4845,N_4391,N_4202);
nand U4846 (N_4846,N_4699,N_4696);
nand U4847 (N_4847,N_4542,N_4301);
nor U4848 (N_4848,N_4409,N_4437);
or U4849 (N_4849,N_4580,N_4703);
or U4850 (N_4850,N_4595,N_4367);
and U4851 (N_4851,N_4737,N_4233);
nand U4852 (N_4852,N_4348,N_4223);
nor U4853 (N_4853,N_4448,N_4493);
nor U4854 (N_4854,N_4641,N_4548);
and U4855 (N_4855,N_4470,N_4701);
or U4856 (N_4856,N_4322,N_4575);
or U4857 (N_4857,N_4566,N_4292);
or U4858 (N_4858,N_4739,N_4420);
xnor U4859 (N_4859,N_4362,N_4215);
or U4860 (N_4860,N_4752,N_4230);
and U4861 (N_4861,N_4784,N_4294);
xnor U4862 (N_4862,N_4298,N_4240);
xor U4863 (N_4863,N_4457,N_4483);
and U4864 (N_4864,N_4423,N_4785);
xor U4865 (N_4865,N_4711,N_4773);
and U4866 (N_4866,N_4763,N_4272);
xnor U4867 (N_4867,N_4366,N_4368);
or U4868 (N_4868,N_4708,N_4724);
or U4869 (N_4869,N_4730,N_4219);
nor U4870 (N_4870,N_4421,N_4505);
nor U4871 (N_4871,N_4634,N_4265);
xnor U4872 (N_4872,N_4517,N_4690);
nor U4873 (N_4873,N_4309,N_4757);
xor U4874 (N_4874,N_4597,N_4565);
nor U4875 (N_4875,N_4714,N_4594);
or U4876 (N_4876,N_4256,N_4476);
and U4877 (N_4877,N_4644,N_4652);
and U4878 (N_4878,N_4255,N_4648);
nor U4879 (N_4879,N_4799,N_4527);
or U4880 (N_4880,N_4487,N_4236);
xnor U4881 (N_4881,N_4683,N_4610);
and U4882 (N_4882,N_4318,N_4798);
nor U4883 (N_4883,N_4682,N_4231);
nor U4884 (N_4884,N_4466,N_4499);
and U4885 (N_4885,N_4553,N_4664);
and U4886 (N_4886,N_4611,N_4523);
or U4887 (N_4887,N_4520,N_4535);
xor U4888 (N_4888,N_4375,N_4556);
and U4889 (N_4889,N_4494,N_4662);
and U4890 (N_4890,N_4522,N_4371);
or U4891 (N_4891,N_4563,N_4349);
xnor U4892 (N_4892,N_4603,N_4728);
xnor U4893 (N_4893,N_4356,N_4395);
or U4894 (N_4894,N_4679,N_4458);
nor U4895 (N_4895,N_4615,N_4498);
and U4896 (N_4896,N_4463,N_4509);
nand U4897 (N_4897,N_4512,N_4317);
nand U4898 (N_4898,N_4790,N_4386);
nor U4899 (N_4899,N_4382,N_4620);
and U4900 (N_4900,N_4341,N_4766);
nor U4901 (N_4901,N_4433,N_4379);
nand U4902 (N_4902,N_4729,N_4649);
and U4903 (N_4903,N_4208,N_4585);
xor U4904 (N_4904,N_4447,N_4334);
and U4905 (N_4905,N_4507,N_4775);
and U4906 (N_4906,N_4459,N_4632);
nor U4907 (N_4907,N_4554,N_4377);
or U4908 (N_4908,N_4707,N_4354);
and U4909 (N_4909,N_4794,N_4624);
and U4910 (N_4910,N_4671,N_4774);
nand U4911 (N_4911,N_4414,N_4640);
xnor U4912 (N_4912,N_4541,N_4510);
nor U4913 (N_4913,N_4647,N_4797);
or U4914 (N_4914,N_4670,N_4286);
nor U4915 (N_4915,N_4452,N_4568);
and U4916 (N_4916,N_4283,N_4278);
or U4917 (N_4917,N_4754,N_4429);
xor U4918 (N_4918,N_4385,N_4257);
xnor U4919 (N_4919,N_4719,N_4412);
or U4920 (N_4920,N_4227,N_4205);
nand U4921 (N_4921,N_4674,N_4273);
xnor U4922 (N_4922,N_4702,N_4760);
nand U4923 (N_4923,N_4705,N_4596);
xnor U4924 (N_4924,N_4567,N_4742);
nor U4925 (N_4925,N_4629,N_4680);
nand U4926 (N_4926,N_4731,N_4287);
nand U4927 (N_4927,N_4704,N_4478);
nand U4928 (N_4928,N_4676,N_4425);
or U4929 (N_4929,N_4578,N_4345);
xor U4930 (N_4930,N_4350,N_4335);
or U4931 (N_4931,N_4687,N_4303);
and U4932 (N_4932,N_4637,N_4538);
and U4933 (N_4933,N_4753,N_4472);
nand U4934 (N_4934,N_4623,N_4544);
xor U4935 (N_4935,N_4446,N_4583);
nor U4936 (N_4936,N_4275,N_4779);
nor U4937 (N_4937,N_4792,N_4207);
nor U4938 (N_4938,N_4307,N_4586);
xnor U4939 (N_4939,N_4451,N_4489);
xor U4940 (N_4940,N_4268,N_4645);
xor U4941 (N_4941,N_4722,N_4306);
and U4942 (N_4942,N_4484,N_4216);
xor U4943 (N_4943,N_4503,N_4288);
and U4944 (N_4944,N_4279,N_4351);
xor U4945 (N_4945,N_4295,N_4337);
or U4946 (N_4946,N_4340,N_4781);
nor U4947 (N_4947,N_4692,N_4249);
xor U4948 (N_4948,N_4689,N_4235);
xnor U4949 (N_4949,N_4712,N_4756);
or U4950 (N_4950,N_4762,N_4282);
and U4951 (N_4951,N_4749,N_4650);
and U4952 (N_4952,N_4357,N_4531);
nor U4953 (N_4953,N_4625,N_4738);
or U4954 (N_4954,N_4333,N_4270);
or U4955 (N_4955,N_4666,N_4297);
nor U4956 (N_4956,N_4392,N_4561);
nand U4957 (N_4957,N_4364,N_4427);
xnor U4958 (N_4958,N_4750,N_4405);
or U4959 (N_4959,N_4352,N_4677);
nand U4960 (N_4960,N_4387,N_4727);
xnor U4961 (N_4961,N_4400,N_4444);
or U4962 (N_4962,N_4768,N_4401);
xor U4963 (N_4963,N_4269,N_4570);
or U4964 (N_4964,N_4612,N_4471);
and U4965 (N_4965,N_4229,N_4607);
nand U4966 (N_4966,N_4519,N_4430);
nand U4967 (N_4967,N_4602,N_4564);
xor U4968 (N_4968,N_4660,N_4488);
or U4969 (N_4969,N_4330,N_4734);
xnor U4970 (N_4970,N_4276,N_4685);
or U4971 (N_4971,N_4305,N_4479);
nor U4972 (N_4972,N_4667,N_4253);
and U4973 (N_4973,N_4363,N_4482);
and U4974 (N_4974,N_4778,N_4434);
nor U4975 (N_4975,N_4245,N_4700);
and U4976 (N_4976,N_4559,N_4481);
or U4977 (N_4977,N_4456,N_4764);
nand U4978 (N_4978,N_4339,N_4525);
or U4979 (N_4979,N_4213,N_4659);
or U4980 (N_4980,N_4480,N_4406);
or U4981 (N_4981,N_4521,N_4608);
or U4982 (N_4982,N_4646,N_4748);
or U4983 (N_4983,N_4740,N_4271);
nor U4984 (N_4984,N_4761,N_4751);
and U4985 (N_4985,N_4694,N_4628);
nor U4986 (N_4986,N_4221,N_4767);
xnor U4987 (N_4987,N_4715,N_4324);
nand U4988 (N_4988,N_4658,N_4247);
nor U4989 (N_4989,N_4299,N_4788);
nand U4990 (N_4990,N_4495,N_4419);
nand U4991 (N_4991,N_4258,N_4442);
xor U4992 (N_4992,N_4581,N_4720);
or U4993 (N_4993,N_4529,N_4262);
nor U4994 (N_4994,N_4591,N_4226);
and U4995 (N_4995,N_4777,N_4314);
and U4996 (N_4996,N_4693,N_4417);
xor U4997 (N_4997,N_4631,N_4327);
and U4998 (N_4998,N_4477,N_4601);
nor U4999 (N_4999,N_4573,N_4360);
and U5000 (N_5000,N_4532,N_4252);
nor U5001 (N_5001,N_4789,N_4403);
nor U5002 (N_5002,N_4284,N_4274);
or U5003 (N_5003,N_4201,N_4323);
or U5004 (N_5004,N_4540,N_4224);
xor U5005 (N_5005,N_4706,N_4678);
xnor U5006 (N_5006,N_4238,N_4642);
or U5007 (N_5007,N_4331,N_4217);
xor U5008 (N_5008,N_4518,N_4786);
nand U5009 (N_5009,N_4254,N_4576);
and U5010 (N_5010,N_4772,N_4263);
xnor U5011 (N_5011,N_4630,N_4765);
nor U5012 (N_5012,N_4638,N_4326);
xnor U5013 (N_5013,N_4709,N_4242);
nor U5014 (N_5014,N_4599,N_4422);
nor U5015 (N_5015,N_4598,N_4758);
nand U5016 (N_5016,N_4551,N_4474);
xnor U5017 (N_5017,N_4462,N_4543);
nand U5018 (N_5018,N_4633,N_4450);
nand U5019 (N_5019,N_4411,N_4302);
or U5020 (N_5020,N_4241,N_4497);
xnor U5021 (N_5021,N_4534,N_4232);
nor U5022 (N_5022,N_4467,N_4508);
and U5023 (N_5023,N_4281,N_4310);
xnor U5024 (N_5024,N_4537,N_4211);
xor U5025 (N_5025,N_4744,N_4415);
or U5026 (N_5026,N_4440,N_4619);
nand U5027 (N_5027,N_4698,N_4514);
nand U5028 (N_5028,N_4552,N_4669);
nand U5029 (N_5029,N_4746,N_4237);
and U5030 (N_5030,N_4741,N_4769);
and U5031 (N_5031,N_4432,N_4315);
or U5032 (N_5032,N_4656,N_4725);
and U5033 (N_5033,N_4783,N_4600);
or U5034 (N_5034,N_4416,N_4469);
or U5035 (N_5035,N_4574,N_4572);
xor U5036 (N_5036,N_4250,N_4261);
xnor U5037 (N_5037,N_4587,N_4343);
xnor U5038 (N_5038,N_4550,N_4404);
nor U5039 (N_5039,N_4782,N_4614);
or U5040 (N_5040,N_4291,N_4588);
xnor U5041 (N_5041,N_4791,N_4312);
nand U5042 (N_5042,N_4445,N_4486);
nand U5043 (N_5043,N_4717,N_4316);
or U5044 (N_5044,N_4285,N_4246);
or U5045 (N_5045,N_4408,N_4439);
and U5046 (N_5046,N_4277,N_4376);
xnor U5047 (N_5047,N_4780,N_4496);
xor U5048 (N_5048,N_4549,N_4358);
or U5049 (N_5049,N_4500,N_4526);
or U5050 (N_5050,N_4370,N_4513);
nor U5051 (N_5051,N_4220,N_4663);
nor U5052 (N_5052,N_4441,N_4795);
nand U5053 (N_5053,N_4336,N_4460);
or U5054 (N_5054,N_4609,N_4267);
xor U5055 (N_5055,N_4651,N_4346);
nor U5056 (N_5056,N_4654,N_4353);
and U5057 (N_5057,N_4502,N_4584);
and U5058 (N_5058,N_4604,N_4776);
or U5059 (N_5059,N_4418,N_4723);
xor U5060 (N_5060,N_4492,N_4248);
nor U5061 (N_5061,N_4755,N_4606);
nand U5062 (N_5062,N_4506,N_4710);
and U5063 (N_5063,N_4397,N_4222);
xnor U5064 (N_5064,N_4733,N_4796);
xor U5065 (N_5065,N_4713,N_4455);
or U5066 (N_5066,N_4410,N_4668);
or U5067 (N_5067,N_4539,N_4204);
nor U5068 (N_5068,N_4383,N_4515);
nor U5069 (N_5069,N_4210,N_4688);
or U5070 (N_5070,N_4251,N_4697);
xnor U5071 (N_5071,N_4214,N_4365);
nand U5072 (N_5072,N_4389,N_4218);
xor U5073 (N_5073,N_4721,N_4743);
or U5074 (N_5074,N_4736,N_4636);
xor U5075 (N_5075,N_4388,N_4661);
xnor U5076 (N_5076,N_4464,N_4304);
xor U5077 (N_5077,N_4557,N_4616);
or U5078 (N_5078,N_4212,N_4613);
nand U5079 (N_5079,N_4718,N_4562);
nand U5080 (N_5080,N_4558,N_4431);
and U5081 (N_5081,N_4516,N_4203);
nand U5082 (N_5082,N_4355,N_4675);
nand U5083 (N_5083,N_4605,N_4560);
nand U5084 (N_5084,N_4545,N_4390);
or U5085 (N_5085,N_4491,N_4206);
xor U5086 (N_5086,N_4626,N_4643);
nor U5087 (N_5087,N_4635,N_4745);
xnor U5088 (N_5088,N_4329,N_4396);
and U5089 (N_5089,N_4239,N_4577);
and U5090 (N_5090,N_4475,N_4555);
xnor U5091 (N_5091,N_4443,N_4266);
or U5092 (N_5092,N_4490,N_4342);
nand U5093 (N_5093,N_4453,N_4686);
or U5094 (N_5094,N_4665,N_4536);
nand U5095 (N_5095,N_4280,N_4359);
xnor U5096 (N_5096,N_4770,N_4290);
and U5097 (N_5097,N_4413,N_4338);
and U5098 (N_5098,N_4384,N_4319);
or U5099 (N_5099,N_4402,N_4653);
nor U5100 (N_5100,N_4553,N_4546);
and U5101 (N_5101,N_4462,N_4634);
or U5102 (N_5102,N_4508,N_4293);
and U5103 (N_5103,N_4673,N_4518);
xor U5104 (N_5104,N_4487,N_4785);
nor U5105 (N_5105,N_4243,N_4782);
xnor U5106 (N_5106,N_4244,N_4727);
or U5107 (N_5107,N_4428,N_4596);
nand U5108 (N_5108,N_4411,N_4629);
and U5109 (N_5109,N_4741,N_4323);
nor U5110 (N_5110,N_4316,N_4329);
nor U5111 (N_5111,N_4220,N_4495);
nand U5112 (N_5112,N_4300,N_4576);
xnor U5113 (N_5113,N_4680,N_4399);
and U5114 (N_5114,N_4215,N_4315);
nor U5115 (N_5115,N_4723,N_4279);
nor U5116 (N_5116,N_4315,N_4522);
nor U5117 (N_5117,N_4560,N_4334);
nor U5118 (N_5118,N_4748,N_4449);
nor U5119 (N_5119,N_4428,N_4416);
and U5120 (N_5120,N_4280,N_4723);
and U5121 (N_5121,N_4265,N_4748);
nand U5122 (N_5122,N_4219,N_4641);
xnor U5123 (N_5123,N_4377,N_4784);
nand U5124 (N_5124,N_4635,N_4612);
nor U5125 (N_5125,N_4615,N_4385);
and U5126 (N_5126,N_4299,N_4319);
nor U5127 (N_5127,N_4707,N_4795);
nand U5128 (N_5128,N_4467,N_4793);
nor U5129 (N_5129,N_4598,N_4585);
xnor U5130 (N_5130,N_4733,N_4226);
xnor U5131 (N_5131,N_4605,N_4686);
or U5132 (N_5132,N_4732,N_4539);
xor U5133 (N_5133,N_4587,N_4592);
and U5134 (N_5134,N_4278,N_4777);
xnor U5135 (N_5135,N_4562,N_4531);
nor U5136 (N_5136,N_4489,N_4240);
or U5137 (N_5137,N_4752,N_4741);
nor U5138 (N_5138,N_4429,N_4424);
nand U5139 (N_5139,N_4211,N_4478);
or U5140 (N_5140,N_4440,N_4369);
nor U5141 (N_5141,N_4731,N_4659);
or U5142 (N_5142,N_4613,N_4633);
and U5143 (N_5143,N_4581,N_4467);
or U5144 (N_5144,N_4364,N_4206);
nand U5145 (N_5145,N_4582,N_4351);
and U5146 (N_5146,N_4331,N_4656);
nor U5147 (N_5147,N_4231,N_4392);
nor U5148 (N_5148,N_4655,N_4535);
xor U5149 (N_5149,N_4207,N_4762);
and U5150 (N_5150,N_4549,N_4367);
or U5151 (N_5151,N_4519,N_4727);
nor U5152 (N_5152,N_4241,N_4703);
and U5153 (N_5153,N_4617,N_4348);
nor U5154 (N_5154,N_4634,N_4745);
nor U5155 (N_5155,N_4229,N_4493);
and U5156 (N_5156,N_4200,N_4319);
nand U5157 (N_5157,N_4565,N_4780);
or U5158 (N_5158,N_4537,N_4523);
and U5159 (N_5159,N_4491,N_4384);
or U5160 (N_5160,N_4608,N_4452);
xor U5161 (N_5161,N_4536,N_4634);
nand U5162 (N_5162,N_4640,N_4681);
and U5163 (N_5163,N_4259,N_4403);
and U5164 (N_5164,N_4267,N_4357);
nand U5165 (N_5165,N_4352,N_4683);
nand U5166 (N_5166,N_4703,N_4386);
or U5167 (N_5167,N_4784,N_4693);
and U5168 (N_5168,N_4237,N_4202);
nand U5169 (N_5169,N_4395,N_4282);
and U5170 (N_5170,N_4697,N_4749);
and U5171 (N_5171,N_4516,N_4452);
nand U5172 (N_5172,N_4477,N_4228);
nor U5173 (N_5173,N_4276,N_4272);
nor U5174 (N_5174,N_4600,N_4529);
nor U5175 (N_5175,N_4413,N_4491);
and U5176 (N_5176,N_4754,N_4779);
xnor U5177 (N_5177,N_4466,N_4592);
xor U5178 (N_5178,N_4589,N_4677);
nor U5179 (N_5179,N_4784,N_4542);
xnor U5180 (N_5180,N_4414,N_4784);
and U5181 (N_5181,N_4761,N_4246);
and U5182 (N_5182,N_4573,N_4227);
and U5183 (N_5183,N_4370,N_4778);
xor U5184 (N_5184,N_4217,N_4270);
or U5185 (N_5185,N_4348,N_4239);
nand U5186 (N_5186,N_4329,N_4451);
nand U5187 (N_5187,N_4248,N_4402);
and U5188 (N_5188,N_4419,N_4415);
xnor U5189 (N_5189,N_4774,N_4610);
or U5190 (N_5190,N_4504,N_4561);
nand U5191 (N_5191,N_4375,N_4210);
or U5192 (N_5192,N_4778,N_4278);
nand U5193 (N_5193,N_4446,N_4338);
nor U5194 (N_5194,N_4249,N_4649);
nor U5195 (N_5195,N_4493,N_4577);
nand U5196 (N_5196,N_4490,N_4658);
xnor U5197 (N_5197,N_4547,N_4232);
and U5198 (N_5198,N_4620,N_4560);
nand U5199 (N_5199,N_4268,N_4285);
or U5200 (N_5200,N_4315,N_4470);
xor U5201 (N_5201,N_4334,N_4482);
nand U5202 (N_5202,N_4712,N_4584);
and U5203 (N_5203,N_4304,N_4603);
and U5204 (N_5204,N_4243,N_4350);
xnor U5205 (N_5205,N_4485,N_4749);
nand U5206 (N_5206,N_4250,N_4450);
xnor U5207 (N_5207,N_4241,N_4570);
nor U5208 (N_5208,N_4349,N_4242);
and U5209 (N_5209,N_4356,N_4309);
or U5210 (N_5210,N_4708,N_4390);
and U5211 (N_5211,N_4624,N_4458);
nand U5212 (N_5212,N_4456,N_4396);
or U5213 (N_5213,N_4592,N_4631);
and U5214 (N_5214,N_4736,N_4567);
or U5215 (N_5215,N_4407,N_4666);
nor U5216 (N_5216,N_4396,N_4740);
nand U5217 (N_5217,N_4397,N_4354);
or U5218 (N_5218,N_4425,N_4773);
nor U5219 (N_5219,N_4568,N_4316);
nor U5220 (N_5220,N_4798,N_4577);
nor U5221 (N_5221,N_4669,N_4777);
and U5222 (N_5222,N_4525,N_4459);
xor U5223 (N_5223,N_4552,N_4284);
xor U5224 (N_5224,N_4470,N_4565);
xnor U5225 (N_5225,N_4471,N_4792);
or U5226 (N_5226,N_4430,N_4444);
nor U5227 (N_5227,N_4603,N_4521);
xnor U5228 (N_5228,N_4548,N_4496);
nand U5229 (N_5229,N_4201,N_4674);
nand U5230 (N_5230,N_4363,N_4551);
nor U5231 (N_5231,N_4632,N_4462);
xor U5232 (N_5232,N_4227,N_4271);
or U5233 (N_5233,N_4561,N_4468);
xor U5234 (N_5234,N_4357,N_4259);
xnor U5235 (N_5235,N_4772,N_4520);
and U5236 (N_5236,N_4534,N_4696);
nand U5237 (N_5237,N_4737,N_4223);
or U5238 (N_5238,N_4540,N_4269);
xor U5239 (N_5239,N_4779,N_4310);
nand U5240 (N_5240,N_4519,N_4629);
nor U5241 (N_5241,N_4769,N_4293);
nor U5242 (N_5242,N_4435,N_4733);
nand U5243 (N_5243,N_4316,N_4264);
nand U5244 (N_5244,N_4694,N_4542);
nand U5245 (N_5245,N_4689,N_4405);
xor U5246 (N_5246,N_4722,N_4658);
or U5247 (N_5247,N_4426,N_4239);
and U5248 (N_5248,N_4594,N_4618);
xor U5249 (N_5249,N_4287,N_4695);
nor U5250 (N_5250,N_4422,N_4378);
and U5251 (N_5251,N_4750,N_4280);
nor U5252 (N_5252,N_4795,N_4628);
nand U5253 (N_5253,N_4638,N_4697);
xnor U5254 (N_5254,N_4411,N_4253);
nand U5255 (N_5255,N_4699,N_4670);
and U5256 (N_5256,N_4220,N_4216);
or U5257 (N_5257,N_4310,N_4302);
nor U5258 (N_5258,N_4519,N_4759);
nand U5259 (N_5259,N_4570,N_4362);
xor U5260 (N_5260,N_4566,N_4513);
xnor U5261 (N_5261,N_4468,N_4721);
xnor U5262 (N_5262,N_4328,N_4722);
xor U5263 (N_5263,N_4645,N_4208);
or U5264 (N_5264,N_4428,N_4353);
and U5265 (N_5265,N_4773,N_4204);
nor U5266 (N_5266,N_4604,N_4365);
nand U5267 (N_5267,N_4272,N_4444);
xor U5268 (N_5268,N_4423,N_4315);
and U5269 (N_5269,N_4376,N_4282);
and U5270 (N_5270,N_4570,N_4691);
nand U5271 (N_5271,N_4314,N_4707);
xnor U5272 (N_5272,N_4622,N_4555);
or U5273 (N_5273,N_4472,N_4305);
xnor U5274 (N_5274,N_4670,N_4628);
nand U5275 (N_5275,N_4669,N_4717);
and U5276 (N_5276,N_4397,N_4506);
nor U5277 (N_5277,N_4424,N_4203);
or U5278 (N_5278,N_4759,N_4674);
xnor U5279 (N_5279,N_4600,N_4662);
and U5280 (N_5280,N_4730,N_4322);
nor U5281 (N_5281,N_4265,N_4611);
nor U5282 (N_5282,N_4699,N_4389);
xnor U5283 (N_5283,N_4701,N_4709);
nor U5284 (N_5284,N_4373,N_4683);
nor U5285 (N_5285,N_4621,N_4750);
or U5286 (N_5286,N_4337,N_4523);
nor U5287 (N_5287,N_4723,N_4295);
xor U5288 (N_5288,N_4707,N_4607);
xor U5289 (N_5289,N_4662,N_4752);
nand U5290 (N_5290,N_4201,N_4504);
and U5291 (N_5291,N_4666,N_4329);
nand U5292 (N_5292,N_4320,N_4406);
and U5293 (N_5293,N_4613,N_4561);
nand U5294 (N_5294,N_4410,N_4667);
nand U5295 (N_5295,N_4585,N_4237);
or U5296 (N_5296,N_4585,N_4548);
and U5297 (N_5297,N_4717,N_4359);
and U5298 (N_5298,N_4722,N_4397);
xnor U5299 (N_5299,N_4777,N_4246);
xor U5300 (N_5300,N_4629,N_4710);
nor U5301 (N_5301,N_4410,N_4324);
nor U5302 (N_5302,N_4785,N_4604);
nand U5303 (N_5303,N_4436,N_4361);
nor U5304 (N_5304,N_4492,N_4309);
nor U5305 (N_5305,N_4475,N_4487);
and U5306 (N_5306,N_4316,N_4373);
nand U5307 (N_5307,N_4288,N_4633);
or U5308 (N_5308,N_4499,N_4404);
or U5309 (N_5309,N_4328,N_4728);
or U5310 (N_5310,N_4286,N_4776);
nand U5311 (N_5311,N_4634,N_4598);
xnor U5312 (N_5312,N_4417,N_4333);
or U5313 (N_5313,N_4450,N_4389);
nand U5314 (N_5314,N_4515,N_4574);
xor U5315 (N_5315,N_4730,N_4432);
or U5316 (N_5316,N_4217,N_4409);
or U5317 (N_5317,N_4623,N_4214);
nand U5318 (N_5318,N_4457,N_4506);
or U5319 (N_5319,N_4785,N_4271);
or U5320 (N_5320,N_4279,N_4731);
nand U5321 (N_5321,N_4583,N_4667);
nor U5322 (N_5322,N_4244,N_4507);
or U5323 (N_5323,N_4398,N_4302);
xnor U5324 (N_5324,N_4211,N_4493);
or U5325 (N_5325,N_4290,N_4482);
or U5326 (N_5326,N_4385,N_4619);
and U5327 (N_5327,N_4585,N_4340);
xnor U5328 (N_5328,N_4334,N_4450);
xor U5329 (N_5329,N_4300,N_4764);
and U5330 (N_5330,N_4618,N_4692);
nand U5331 (N_5331,N_4395,N_4238);
nand U5332 (N_5332,N_4791,N_4380);
nor U5333 (N_5333,N_4274,N_4375);
or U5334 (N_5334,N_4547,N_4273);
and U5335 (N_5335,N_4708,N_4686);
and U5336 (N_5336,N_4224,N_4699);
nand U5337 (N_5337,N_4317,N_4629);
or U5338 (N_5338,N_4388,N_4233);
nor U5339 (N_5339,N_4708,N_4527);
and U5340 (N_5340,N_4419,N_4580);
xor U5341 (N_5341,N_4606,N_4741);
or U5342 (N_5342,N_4475,N_4270);
and U5343 (N_5343,N_4219,N_4649);
nand U5344 (N_5344,N_4703,N_4371);
or U5345 (N_5345,N_4475,N_4533);
xnor U5346 (N_5346,N_4581,N_4532);
nor U5347 (N_5347,N_4307,N_4624);
nand U5348 (N_5348,N_4715,N_4604);
xor U5349 (N_5349,N_4634,N_4645);
nor U5350 (N_5350,N_4259,N_4750);
or U5351 (N_5351,N_4557,N_4506);
or U5352 (N_5352,N_4572,N_4311);
nand U5353 (N_5353,N_4640,N_4331);
nand U5354 (N_5354,N_4562,N_4737);
and U5355 (N_5355,N_4392,N_4540);
nor U5356 (N_5356,N_4363,N_4787);
nor U5357 (N_5357,N_4659,N_4681);
nand U5358 (N_5358,N_4210,N_4495);
or U5359 (N_5359,N_4477,N_4578);
nor U5360 (N_5360,N_4470,N_4342);
xnor U5361 (N_5361,N_4216,N_4563);
nand U5362 (N_5362,N_4355,N_4415);
or U5363 (N_5363,N_4488,N_4288);
nor U5364 (N_5364,N_4421,N_4686);
and U5365 (N_5365,N_4649,N_4358);
nand U5366 (N_5366,N_4654,N_4496);
xnor U5367 (N_5367,N_4451,N_4265);
or U5368 (N_5368,N_4302,N_4689);
nor U5369 (N_5369,N_4418,N_4449);
nor U5370 (N_5370,N_4586,N_4724);
or U5371 (N_5371,N_4665,N_4761);
or U5372 (N_5372,N_4620,N_4739);
nand U5373 (N_5373,N_4239,N_4428);
nand U5374 (N_5374,N_4744,N_4433);
xnor U5375 (N_5375,N_4476,N_4606);
xnor U5376 (N_5376,N_4239,N_4324);
nand U5377 (N_5377,N_4474,N_4303);
and U5378 (N_5378,N_4466,N_4559);
or U5379 (N_5379,N_4559,N_4378);
and U5380 (N_5380,N_4266,N_4242);
and U5381 (N_5381,N_4590,N_4799);
and U5382 (N_5382,N_4466,N_4313);
and U5383 (N_5383,N_4514,N_4275);
or U5384 (N_5384,N_4631,N_4449);
xor U5385 (N_5385,N_4623,N_4794);
nor U5386 (N_5386,N_4287,N_4616);
and U5387 (N_5387,N_4566,N_4308);
and U5388 (N_5388,N_4653,N_4287);
nor U5389 (N_5389,N_4630,N_4607);
xor U5390 (N_5390,N_4577,N_4738);
nand U5391 (N_5391,N_4654,N_4326);
and U5392 (N_5392,N_4728,N_4584);
nand U5393 (N_5393,N_4772,N_4465);
and U5394 (N_5394,N_4586,N_4674);
nand U5395 (N_5395,N_4393,N_4713);
nand U5396 (N_5396,N_4550,N_4361);
nand U5397 (N_5397,N_4656,N_4237);
nand U5398 (N_5398,N_4773,N_4211);
xor U5399 (N_5399,N_4526,N_4401);
nor U5400 (N_5400,N_4961,N_5028);
or U5401 (N_5401,N_5017,N_5105);
and U5402 (N_5402,N_4911,N_4842);
nor U5403 (N_5403,N_5221,N_4947);
or U5404 (N_5404,N_4995,N_5037);
nand U5405 (N_5405,N_4991,N_4993);
nor U5406 (N_5406,N_5324,N_5067);
nand U5407 (N_5407,N_4808,N_5129);
xor U5408 (N_5408,N_4968,N_5008);
and U5409 (N_5409,N_4813,N_5298);
and U5410 (N_5410,N_4800,N_5378);
nand U5411 (N_5411,N_5228,N_5155);
nand U5412 (N_5412,N_5262,N_5281);
or U5413 (N_5413,N_5388,N_5394);
nor U5414 (N_5414,N_5166,N_5000);
nor U5415 (N_5415,N_5391,N_5360);
and U5416 (N_5416,N_5106,N_5347);
xor U5417 (N_5417,N_4985,N_5261);
nand U5418 (N_5418,N_4957,N_4871);
xnor U5419 (N_5419,N_5119,N_4830);
nand U5420 (N_5420,N_4989,N_5098);
nor U5421 (N_5421,N_4858,N_5024);
and U5422 (N_5422,N_4884,N_5030);
or U5423 (N_5423,N_4918,N_5237);
xnor U5424 (N_5424,N_5308,N_5303);
nand U5425 (N_5425,N_5134,N_5160);
nor U5426 (N_5426,N_5173,N_4907);
nor U5427 (N_5427,N_5276,N_5260);
xnor U5428 (N_5428,N_5003,N_5123);
xnor U5429 (N_5429,N_5014,N_4945);
and U5430 (N_5430,N_5361,N_4988);
nor U5431 (N_5431,N_5265,N_5257);
nor U5432 (N_5432,N_4978,N_5002);
xor U5433 (N_5433,N_5384,N_4937);
nor U5434 (N_5434,N_5127,N_5194);
or U5435 (N_5435,N_5269,N_4929);
or U5436 (N_5436,N_4867,N_5035);
and U5437 (N_5437,N_5337,N_4891);
and U5438 (N_5438,N_5329,N_4893);
xor U5439 (N_5439,N_5353,N_4981);
and U5440 (N_5440,N_5079,N_5357);
and U5441 (N_5441,N_5182,N_5006);
nor U5442 (N_5442,N_4831,N_5231);
xnor U5443 (N_5443,N_4987,N_5332);
and U5444 (N_5444,N_5310,N_4827);
nor U5445 (N_5445,N_5007,N_4982);
or U5446 (N_5446,N_5158,N_5051);
nor U5447 (N_5447,N_4976,N_4856);
or U5448 (N_5448,N_5043,N_5187);
nand U5449 (N_5449,N_5009,N_5235);
nand U5450 (N_5450,N_5141,N_4874);
xnor U5451 (N_5451,N_5382,N_5033);
xor U5452 (N_5452,N_4977,N_5131);
and U5453 (N_5453,N_4924,N_5052);
xor U5454 (N_5454,N_4927,N_4926);
or U5455 (N_5455,N_5071,N_5075);
nor U5456 (N_5456,N_4885,N_4857);
nand U5457 (N_5457,N_4928,N_5211);
nand U5458 (N_5458,N_5209,N_5338);
nor U5459 (N_5459,N_4906,N_4805);
or U5460 (N_5460,N_5188,N_5143);
xor U5461 (N_5461,N_5295,N_5316);
nand U5462 (N_5462,N_5090,N_4815);
or U5463 (N_5463,N_4963,N_4921);
or U5464 (N_5464,N_4868,N_5056);
xor U5465 (N_5465,N_5251,N_5040);
nor U5466 (N_5466,N_4994,N_5393);
nand U5467 (N_5467,N_5199,N_5088);
and U5468 (N_5468,N_4999,N_5038);
or U5469 (N_5469,N_4912,N_4922);
nor U5470 (N_5470,N_5138,N_5020);
or U5471 (N_5471,N_5306,N_5004);
or U5472 (N_5472,N_5381,N_5026);
nor U5473 (N_5473,N_5241,N_5159);
nand U5474 (N_5474,N_5317,N_5059);
xor U5475 (N_5475,N_4853,N_5366);
nor U5476 (N_5476,N_5321,N_5350);
nand U5477 (N_5477,N_5248,N_5323);
or U5478 (N_5478,N_4939,N_4938);
or U5479 (N_5479,N_5046,N_4872);
or U5480 (N_5480,N_5149,N_5358);
or U5481 (N_5481,N_4930,N_5132);
nand U5482 (N_5482,N_5266,N_5197);
and U5483 (N_5483,N_5163,N_5085);
nand U5484 (N_5484,N_4886,N_5124);
xnor U5485 (N_5485,N_5282,N_5230);
or U5486 (N_5486,N_5270,N_4946);
xnor U5487 (N_5487,N_5117,N_5354);
nor U5488 (N_5488,N_5076,N_5184);
nor U5489 (N_5489,N_4895,N_5325);
nor U5490 (N_5490,N_5355,N_5278);
nor U5491 (N_5491,N_5299,N_5379);
xnor U5492 (N_5492,N_5147,N_5082);
and U5493 (N_5493,N_4866,N_5128);
nand U5494 (N_5494,N_5320,N_5144);
nor U5495 (N_5495,N_4801,N_5212);
or U5496 (N_5496,N_5207,N_5178);
and U5497 (N_5497,N_5372,N_4960);
or U5498 (N_5498,N_4920,N_5240);
nand U5499 (N_5499,N_4948,N_5263);
nor U5500 (N_5500,N_5239,N_4950);
and U5501 (N_5501,N_4863,N_4917);
nor U5502 (N_5502,N_5191,N_5068);
or U5503 (N_5503,N_5198,N_5275);
or U5504 (N_5504,N_5005,N_5179);
xor U5505 (N_5505,N_4969,N_5218);
or U5506 (N_5506,N_5034,N_4826);
nor U5507 (N_5507,N_5335,N_5377);
xnor U5508 (N_5508,N_5204,N_5150);
nand U5509 (N_5509,N_4971,N_4965);
or U5510 (N_5510,N_4802,N_5193);
xnor U5511 (N_5511,N_5313,N_5322);
nand U5512 (N_5512,N_5219,N_5208);
nor U5513 (N_5513,N_4975,N_4835);
xnor U5514 (N_5514,N_4958,N_5289);
xnor U5515 (N_5515,N_5121,N_4925);
or U5516 (N_5516,N_5063,N_5195);
xnor U5517 (N_5517,N_5114,N_5293);
and U5518 (N_5518,N_5380,N_5081);
xnor U5519 (N_5519,N_5302,N_4845);
xnor U5520 (N_5520,N_4878,N_5069);
and U5521 (N_5521,N_4889,N_5120);
and U5522 (N_5522,N_5162,N_5365);
nor U5523 (N_5523,N_5174,N_5042);
nand U5524 (N_5524,N_4953,N_4941);
and U5525 (N_5525,N_5074,N_5255);
xnor U5526 (N_5526,N_4823,N_5236);
nor U5527 (N_5527,N_4903,N_5001);
nand U5528 (N_5528,N_5374,N_5122);
or U5529 (N_5529,N_5012,N_5053);
and U5530 (N_5530,N_5383,N_4850);
nand U5531 (N_5531,N_5154,N_4942);
xnor U5532 (N_5532,N_5346,N_5238);
nand U5533 (N_5533,N_4964,N_5078);
xor U5534 (N_5534,N_5362,N_4905);
xor U5535 (N_5535,N_5061,N_5058);
or U5536 (N_5536,N_4869,N_5330);
nor U5537 (N_5537,N_5140,N_5274);
or U5538 (N_5538,N_5151,N_4882);
nor U5539 (N_5539,N_4908,N_5213);
or U5540 (N_5540,N_5291,N_5279);
xnor U5541 (N_5541,N_5364,N_5334);
or U5542 (N_5542,N_4998,N_5258);
nand U5543 (N_5543,N_5373,N_5234);
xnor U5544 (N_5544,N_5185,N_5227);
nor U5545 (N_5545,N_5080,N_5169);
nand U5546 (N_5546,N_5328,N_5153);
xnor U5547 (N_5547,N_5290,N_5060);
or U5548 (N_5548,N_4973,N_5376);
or U5549 (N_5549,N_5062,N_5267);
xor U5550 (N_5550,N_5152,N_5319);
and U5551 (N_5551,N_5342,N_4898);
xnor U5552 (N_5552,N_5250,N_5139);
or U5553 (N_5553,N_5047,N_4862);
nand U5554 (N_5554,N_5101,N_4833);
and U5555 (N_5555,N_5205,N_5215);
xnor U5556 (N_5556,N_5351,N_4841);
nand U5557 (N_5557,N_4851,N_5089);
nor U5558 (N_5558,N_5224,N_5167);
xnor U5559 (N_5559,N_5156,N_5126);
nand U5560 (N_5560,N_5148,N_4811);
and U5561 (N_5561,N_4967,N_4966);
xor U5562 (N_5562,N_5375,N_4897);
and U5563 (N_5563,N_5192,N_5259);
xor U5564 (N_5564,N_5170,N_5200);
xor U5565 (N_5565,N_4980,N_4996);
nor U5566 (N_5566,N_5217,N_5064);
nand U5567 (N_5567,N_5049,N_5084);
or U5568 (N_5568,N_5116,N_4888);
xor U5569 (N_5569,N_5369,N_4847);
or U5570 (N_5570,N_5363,N_5368);
xnor U5571 (N_5571,N_5157,N_4936);
and U5572 (N_5572,N_5183,N_5109);
nand U5573 (N_5573,N_4865,N_4812);
and U5574 (N_5574,N_5091,N_4859);
or U5575 (N_5575,N_5386,N_5083);
and U5576 (N_5576,N_5339,N_4970);
or U5577 (N_5577,N_5304,N_4954);
nand U5578 (N_5578,N_4890,N_5271);
or U5579 (N_5579,N_4875,N_4949);
xor U5580 (N_5580,N_5093,N_5073);
nand U5581 (N_5581,N_5284,N_5253);
or U5582 (N_5582,N_4984,N_4913);
or U5583 (N_5583,N_5110,N_4959);
xor U5584 (N_5584,N_5107,N_5130);
nand U5585 (N_5585,N_5301,N_5390);
nor U5586 (N_5586,N_5318,N_4838);
nor U5587 (N_5587,N_4931,N_4894);
and U5588 (N_5588,N_5296,N_4849);
nor U5589 (N_5589,N_4990,N_5222);
and U5590 (N_5590,N_5327,N_5243);
and U5591 (N_5591,N_4951,N_5272);
and U5592 (N_5592,N_5086,N_4879);
xnor U5593 (N_5593,N_5055,N_5387);
nor U5594 (N_5594,N_5229,N_4877);
and U5595 (N_5595,N_5181,N_5010);
xnor U5596 (N_5596,N_5018,N_4914);
and U5597 (N_5597,N_5349,N_5118);
nor U5598 (N_5598,N_5196,N_5135);
or U5599 (N_5599,N_5095,N_5226);
or U5600 (N_5600,N_4979,N_5142);
xor U5601 (N_5601,N_4821,N_4820);
or U5602 (N_5602,N_4870,N_5113);
nor U5603 (N_5603,N_5343,N_4825);
nor U5604 (N_5604,N_4846,N_5168);
nor U5605 (N_5605,N_4818,N_4901);
nand U5606 (N_5606,N_5125,N_5264);
nand U5607 (N_5607,N_5044,N_5172);
nand U5608 (N_5608,N_4814,N_5385);
nand U5609 (N_5609,N_5203,N_4983);
or U5610 (N_5610,N_4956,N_4940);
nor U5611 (N_5611,N_4915,N_4997);
or U5612 (N_5612,N_4902,N_4974);
xor U5613 (N_5613,N_4840,N_5225);
nor U5614 (N_5614,N_4803,N_5025);
xnor U5615 (N_5615,N_5331,N_4828);
and U5616 (N_5616,N_4900,N_5297);
nand U5617 (N_5617,N_5161,N_5341);
xnor U5618 (N_5618,N_5016,N_5104);
nand U5619 (N_5619,N_4962,N_5097);
nand U5620 (N_5620,N_5392,N_5108);
nand U5621 (N_5621,N_4839,N_4873);
nor U5622 (N_5622,N_5345,N_4881);
and U5623 (N_5623,N_5036,N_5111);
nor U5624 (N_5624,N_5072,N_4880);
nor U5625 (N_5625,N_4916,N_5244);
nor U5626 (N_5626,N_5309,N_5359);
nand U5627 (N_5627,N_5054,N_4919);
nand U5628 (N_5628,N_5277,N_5395);
xor U5629 (N_5629,N_5136,N_5344);
or U5630 (N_5630,N_5232,N_4829);
nand U5631 (N_5631,N_4934,N_4822);
nor U5632 (N_5632,N_5397,N_5077);
or U5633 (N_5633,N_5396,N_4816);
xor U5634 (N_5634,N_5210,N_5294);
and U5635 (N_5635,N_5050,N_5112);
or U5636 (N_5636,N_5186,N_5177);
nand U5637 (N_5637,N_5307,N_4836);
nand U5638 (N_5638,N_4807,N_4844);
or U5639 (N_5639,N_4923,N_4876);
xor U5640 (N_5640,N_4933,N_5220);
nor U5641 (N_5641,N_5065,N_4809);
xor U5642 (N_5642,N_5146,N_5249);
or U5643 (N_5643,N_5340,N_5286);
nand U5644 (N_5644,N_4944,N_5094);
and U5645 (N_5645,N_5022,N_5145);
or U5646 (N_5646,N_5370,N_5326);
xnor U5647 (N_5647,N_5070,N_4932);
nor U5648 (N_5648,N_5314,N_5133);
nand U5649 (N_5649,N_5245,N_5015);
or U5650 (N_5650,N_4864,N_4909);
and U5651 (N_5651,N_4832,N_5312);
xnor U5652 (N_5652,N_5287,N_5292);
nand U5653 (N_5653,N_5216,N_5288);
and U5654 (N_5654,N_5039,N_5206);
nor U5655 (N_5655,N_5171,N_5180);
or U5656 (N_5656,N_5398,N_5164);
nor U5657 (N_5657,N_4837,N_5189);
nor U5658 (N_5658,N_5202,N_5214);
nand U5659 (N_5659,N_5019,N_5256);
nand U5660 (N_5660,N_4972,N_4910);
xor U5661 (N_5661,N_5103,N_5201);
and U5662 (N_5662,N_5367,N_4804);
nand U5663 (N_5663,N_4817,N_5285);
nor U5664 (N_5664,N_4883,N_5048);
nor U5665 (N_5665,N_4819,N_5371);
xor U5666 (N_5666,N_5092,N_5096);
nor U5667 (N_5667,N_5031,N_5246);
nand U5668 (N_5668,N_4834,N_4904);
xor U5669 (N_5669,N_5315,N_5102);
nor U5670 (N_5670,N_5252,N_5057);
nand U5671 (N_5671,N_5352,N_4892);
nor U5672 (N_5672,N_5280,N_5041);
nand U5673 (N_5673,N_4860,N_4986);
or U5674 (N_5674,N_5099,N_4952);
xor U5675 (N_5675,N_4843,N_5087);
or U5676 (N_5676,N_5023,N_5190);
and U5677 (N_5677,N_5242,N_5254);
nand U5678 (N_5678,N_4896,N_4806);
nand U5679 (N_5679,N_5045,N_5032);
xor U5680 (N_5680,N_4935,N_5348);
nor U5681 (N_5681,N_4854,N_5175);
xnor U5682 (N_5682,N_4899,N_5273);
nand U5683 (N_5683,N_4848,N_5399);
and U5684 (N_5684,N_5029,N_5305);
nand U5685 (N_5685,N_4824,N_5223);
and U5686 (N_5686,N_4861,N_4943);
or U5687 (N_5687,N_5011,N_5066);
xor U5688 (N_5688,N_5165,N_5356);
xor U5689 (N_5689,N_5021,N_5283);
or U5690 (N_5690,N_5115,N_5333);
and U5691 (N_5691,N_4852,N_5027);
and U5692 (N_5692,N_4955,N_5311);
nor U5693 (N_5693,N_5336,N_5137);
xnor U5694 (N_5694,N_4810,N_5389);
xnor U5695 (N_5695,N_5176,N_5233);
nor U5696 (N_5696,N_5013,N_5300);
and U5697 (N_5697,N_4887,N_5247);
or U5698 (N_5698,N_5100,N_4855);
nor U5699 (N_5699,N_4992,N_5268);
and U5700 (N_5700,N_4816,N_5301);
or U5701 (N_5701,N_4816,N_4928);
or U5702 (N_5702,N_5033,N_5296);
and U5703 (N_5703,N_4871,N_5025);
nor U5704 (N_5704,N_5113,N_5287);
xor U5705 (N_5705,N_5153,N_5072);
nand U5706 (N_5706,N_5294,N_4874);
and U5707 (N_5707,N_4841,N_5283);
or U5708 (N_5708,N_4881,N_5195);
nand U5709 (N_5709,N_5075,N_4980);
nor U5710 (N_5710,N_5330,N_5289);
xor U5711 (N_5711,N_5286,N_5068);
nand U5712 (N_5712,N_5267,N_4828);
nor U5713 (N_5713,N_4828,N_4935);
nor U5714 (N_5714,N_5330,N_5098);
nor U5715 (N_5715,N_4826,N_4884);
xor U5716 (N_5716,N_5345,N_5204);
or U5717 (N_5717,N_5238,N_5322);
and U5718 (N_5718,N_5091,N_5209);
or U5719 (N_5719,N_4971,N_5366);
and U5720 (N_5720,N_5340,N_5139);
and U5721 (N_5721,N_5216,N_4992);
nor U5722 (N_5722,N_5030,N_5283);
nor U5723 (N_5723,N_5212,N_5210);
nor U5724 (N_5724,N_4972,N_5164);
nor U5725 (N_5725,N_4854,N_5163);
nor U5726 (N_5726,N_4947,N_5382);
nor U5727 (N_5727,N_4859,N_4898);
xnor U5728 (N_5728,N_5270,N_5119);
xnor U5729 (N_5729,N_4986,N_5213);
nand U5730 (N_5730,N_5352,N_5219);
nand U5731 (N_5731,N_4824,N_4811);
nand U5732 (N_5732,N_4923,N_5203);
or U5733 (N_5733,N_4966,N_5217);
nor U5734 (N_5734,N_4976,N_4932);
nor U5735 (N_5735,N_5362,N_5209);
nand U5736 (N_5736,N_5268,N_5158);
xnor U5737 (N_5737,N_4848,N_4869);
xor U5738 (N_5738,N_4897,N_5247);
or U5739 (N_5739,N_4829,N_5231);
and U5740 (N_5740,N_5377,N_5387);
or U5741 (N_5741,N_4904,N_5153);
nand U5742 (N_5742,N_4940,N_4825);
xnor U5743 (N_5743,N_4866,N_5379);
nor U5744 (N_5744,N_4926,N_4946);
and U5745 (N_5745,N_5177,N_4806);
nand U5746 (N_5746,N_5267,N_5103);
xor U5747 (N_5747,N_5151,N_4847);
or U5748 (N_5748,N_4981,N_5380);
nor U5749 (N_5749,N_5109,N_5225);
nor U5750 (N_5750,N_5392,N_4998);
nor U5751 (N_5751,N_5113,N_5257);
and U5752 (N_5752,N_5152,N_4978);
nor U5753 (N_5753,N_5175,N_4937);
and U5754 (N_5754,N_5055,N_5138);
or U5755 (N_5755,N_5250,N_5280);
nor U5756 (N_5756,N_5084,N_4989);
or U5757 (N_5757,N_5094,N_5295);
xnor U5758 (N_5758,N_4818,N_5244);
and U5759 (N_5759,N_5113,N_5032);
and U5760 (N_5760,N_5073,N_5075);
nor U5761 (N_5761,N_5207,N_5126);
or U5762 (N_5762,N_5237,N_5017);
and U5763 (N_5763,N_4833,N_4852);
or U5764 (N_5764,N_5174,N_4855);
and U5765 (N_5765,N_4959,N_5186);
xnor U5766 (N_5766,N_5093,N_5214);
nand U5767 (N_5767,N_5035,N_4842);
or U5768 (N_5768,N_5345,N_5281);
or U5769 (N_5769,N_4934,N_4907);
xor U5770 (N_5770,N_4862,N_4849);
nand U5771 (N_5771,N_5150,N_5026);
xor U5772 (N_5772,N_5229,N_5045);
and U5773 (N_5773,N_5311,N_4839);
and U5774 (N_5774,N_5119,N_4895);
nand U5775 (N_5775,N_4872,N_5098);
nand U5776 (N_5776,N_4924,N_5158);
or U5777 (N_5777,N_5369,N_5330);
and U5778 (N_5778,N_5380,N_4984);
xor U5779 (N_5779,N_5358,N_5085);
nand U5780 (N_5780,N_4885,N_4802);
or U5781 (N_5781,N_5374,N_4899);
or U5782 (N_5782,N_5385,N_4972);
nor U5783 (N_5783,N_4971,N_4902);
and U5784 (N_5784,N_5333,N_4868);
xor U5785 (N_5785,N_4893,N_5038);
nand U5786 (N_5786,N_4914,N_5332);
nand U5787 (N_5787,N_5086,N_5393);
and U5788 (N_5788,N_5192,N_5234);
or U5789 (N_5789,N_5121,N_5323);
or U5790 (N_5790,N_5120,N_4944);
xor U5791 (N_5791,N_4839,N_5268);
nand U5792 (N_5792,N_5291,N_5247);
or U5793 (N_5793,N_5012,N_5332);
nor U5794 (N_5794,N_4846,N_4869);
and U5795 (N_5795,N_5030,N_5203);
nor U5796 (N_5796,N_5328,N_5368);
xnor U5797 (N_5797,N_5261,N_5198);
or U5798 (N_5798,N_5001,N_5048);
or U5799 (N_5799,N_5250,N_4824);
nand U5800 (N_5800,N_4869,N_5242);
and U5801 (N_5801,N_5002,N_5011);
nand U5802 (N_5802,N_4827,N_5025);
nor U5803 (N_5803,N_5360,N_5091);
or U5804 (N_5804,N_5279,N_5275);
and U5805 (N_5805,N_5235,N_5228);
xor U5806 (N_5806,N_4924,N_5221);
nor U5807 (N_5807,N_5366,N_5035);
and U5808 (N_5808,N_5199,N_5363);
nand U5809 (N_5809,N_5249,N_5151);
nor U5810 (N_5810,N_5081,N_4912);
nand U5811 (N_5811,N_5335,N_5275);
or U5812 (N_5812,N_5081,N_5230);
or U5813 (N_5813,N_5020,N_5220);
nand U5814 (N_5814,N_5297,N_5179);
nor U5815 (N_5815,N_5022,N_5051);
xor U5816 (N_5816,N_5240,N_5067);
xnor U5817 (N_5817,N_5131,N_4926);
nor U5818 (N_5818,N_4809,N_5132);
nor U5819 (N_5819,N_5320,N_4915);
xnor U5820 (N_5820,N_4965,N_5013);
xnor U5821 (N_5821,N_4919,N_5008);
xnor U5822 (N_5822,N_5217,N_4959);
nor U5823 (N_5823,N_5288,N_4995);
nor U5824 (N_5824,N_5359,N_5136);
nand U5825 (N_5825,N_4885,N_5305);
or U5826 (N_5826,N_4909,N_5125);
nor U5827 (N_5827,N_4892,N_4857);
and U5828 (N_5828,N_4895,N_4855);
and U5829 (N_5829,N_5213,N_5385);
and U5830 (N_5830,N_5033,N_5221);
nand U5831 (N_5831,N_4833,N_5084);
nor U5832 (N_5832,N_4917,N_5256);
xor U5833 (N_5833,N_5191,N_5130);
or U5834 (N_5834,N_4805,N_5118);
nand U5835 (N_5835,N_5366,N_5270);
nand U5836 (N_5836,N_5046,N_4989);
and U5837 (N_5837,N_5343,N_5367);
or U5838 (N_5838,N_4994,N_5128);
and U5839 (N_5839,N_5264,N_4837);
and U5840 (N_5840,N_4974,N_5261);
or U5841 (N_5841,N_4881,N_5391);
or U5842 (N_5842,N_5104,N_5132);
and U5843 (N_5843,N_5064,N_4830);
and U5844 (N_5844,N_4983,N_4987);
nor U5845 (N_5845,N_5270,N_5314);
nand U5846 (N_5846,N_5342,N_5123);
or U5847 (N_5847,N_4943,N_5194);
nand U5848 (N_5848,N_4861,N_4907);
and U5849 (N_5849,N_5023,N_5325);
nor U5850 (N_5850,N_4809,N_4891);
or U5851 (N_5851,N_5265,N_4817);
or U5852 (N_5852,N_5316,N_5119);
or U5853 (N_5853,N_5226,N_4875);
or U5854 (N_5854,N_5315,N_4934);
or U5855 (N_5855,N_5314,N_5172);
nor U5856 (N_5856,N_5128,N_4850);
nand U5857 (N_5857,N_5293,N_4858);
nor U5858 (N_5858,N_5354,N_5216);
and U5859 (N_5859,N_5145,N_5265);
or U5860 (N_5860,N_4878,N_5267);
nor U5861 (N_5861,N_5344,N_5358);
nor U5862 (N_5862,N_5284,N_5190);
nand U5863 (N_5863,N_5232,N_5068);
or U5864 (N_5864,N_5006,N_5160);
and U5865 (N_5865,N_4826,N_5113);
nand U5866 (N_5866,N_4867,N_5340);
nand U5867 (N_5867,N_5052,N_5372);
and U5868 (N_5868,N_4870,N_5349);
nor U5869 (N_5869,N_5384,N_4898);
nor U5870 (N_5870,N_5243,N_4964);
or U5871 (N_5871,N_4868,N_5046);
nand U5872 (N_5872,N_4901,N_5028);
nor U5873 (N_5873,N_5301,N_5334);
nand U5874 (N_5874,N_5027,N_5387);
nor U5875 (N_5875,N_5324,N_5378);
xor U5876 (N_5876,N_5259,N_4836);
nand U5877 (N_5877,N_5185,N_5203);
xor U5878 (N_5878,N_5026,N_5105);
nand U5879 (N_5879,N_5346,N_5188);
nand U5880 (N_5880,N_4907,N_4967);
nand U5881 (N_5881,N_5392,N_5337);
xor U5882 (N_5882,N_4851,N_5074);
xor U5883 (N_5883,N_5255,N_5017);
xnor U5884 (N_5884,N_5342,N_5285);
nand U5885 (N_5885,N_5240,N_5063);
or U5886 (N_5886,N_5298,N_5381);
nor U5887 (N_5887,N_4925,N_5189);
nand U5888 (N_5888,N_5032,N_4982);
nor U5889 (N_5889,N_4857,N_4830);
xor U5890 (N_5890,N_4945,N_5197);
nor U5891 (N_5891,N_5367,N_5200);
xnor U5892 (N_5892,N_5143,N_5281);
nand U5893 (N_5893,N_5009,N_4907);
nor U5894 (N_5894,N_4852,N_5166);
and U5895 (N_5895,N_5013,N_5136);
or U5896 (N_5896,N_5275,N_4833);
nor U5897 (N_5897,N_5092,N_4924);
nand U5898 (N_5898,N_4917,N_5187);
xnor U5899 (N_5899,N_4901,N_5021);
xnor U5900 (N_5900,N_5379,N_5057);
or U5901 (N_5901,N_4930,N_5242);
and U5902 (N_5902,N_5264,N_5082);
or U5903 (N_5903,N_5093,N_5008);
nand U5904 (N_5904,N_5096,N_4856);
xor U5905 (N_5905,N_5162,N_5062);
nand U5906 (N_5906,N_4834,N_5214);
or U5907 (N_5907,N_4878,N_4946);
or U5908 (N_5908,N_5209,N_4873);
nor U5909 (N_5909,N_5104,N_5095);
nor U5910 (N_5910,N_4968,N_5139);
nor U5911 (N_5911,N_5383,N_5279);
and U5912 (N_5912,N_5078,N_5336);
and U5913 (N_5913,N_4941,N_4896);
nor U5914 (N_5914,N_5075,N_5088);
or U5915 (N_5915,N_5046,N_5266);
xnor U5916 (N_5916,N_5116,N_4936);
and U5917 (N_5917,N_5236,N_5156);
xor U5918 (N_5918,N_5155,N_4877);
xnor U5919 (N_5919,N_5374,N_5265);
or U5920 (N_5920,N_4967,N_4848);
or U5921 (N_5921,N_4835,N_4950);
nor U5922 (N_5922,N_5345,N_5354);
or U5923 (N_5923,N_4808,N_5284);
xor U5924 (N_5924,N_5205,N_5379);
or U5925 (N_5925,N_5332,N_5148);
nor U5926 (N_5926,N_5312,N_5118);
or U5927 (N_5927,N_5018,N_5397);
and U5928 (N_5928,N_5092,N_4867);
xor U5929 (N_5929,N_5150,N_5341);
nand U5930 (N_5930,N_5024,N_4982);
or U5931 (N_5931,N_5089,N_4872);
or U5932 (N_5932,N_5295,N_5221);
xor U5933 (N_5933,N_5040,N_4948);
nor U5934 (N_5934,N_5214,N_5013);
xnor U5935 (N_5935,N_5395,N_4992);
nor U5936 (N_5936,N_5004,N_5034);
xor U5937 (N_5937,N_5347,N_4934);
or U5938 (N_5938,N_5308,N_4955);
and U5939 (N_5939,N_4864,N_5312);
nor U5940 (N_5940,N_5196,N_5236);
nand U5941 (N_5941,N_5120,N_5243);
nand U5942 (N_5942,N_5107,N_5365);
xor U5943 (N_5943,N_5266,N_5145);
xnor U5944 (N_5944,N_5020,N_4961);
or U5945 (N_5945,N_5046,N_5206);
nand U5946 (N_5946,N_5243,N_5258);
xnor U5947 (N_5947,N_4844,N_4833);
and U5948 (N_5948,N_4840,N_4907);
and U5949 (N_5949,N_4967,N_4889);
nor U5950 (N_5950,N_5046,N_5388);
and U5951 (N_5951,N_5084,N_5275);
xor U5952 (N_5952,N_4916,N_5316);
xor U5953 (N_5953,N_5259,N_4831);
nor U5954 (N_5954,N_5144,N_4866);
or U5955 (N_5955,N_5014,N_5323);
or U5956 (N_5956,N_5054,N_5172);
xnor U5957 (N_5957,N_5026,N_5217);
nor U5958 (N_5958,N_5351,N_5035);
or U5959 (N_5959,N_5228,N_4814);
or U5960 (N_5960,N_4848,N_5202);
nand U5961 (N_5961,N_5161,N_4826);
and U5962 (N_5962,N_5067,N_4892);
nor U5963 (N_5963,N_5136,N_5262);
and U5964 (N_5964,N_5360,N_5163);
nor U5965 (N_5965,N_5045,N_4971);
or U5966 (N_5966,N_5177,N_5383);
xnor U5967 (N_5967,N_5202,N_5138);
and U5968 (N_5968,N_4815,N_4914);
and U5969 (N_5969,N_5262,N_5035);
nand U5970 (N_5970,N_4898,N_4884);
nor U5971 (N_5971,N_5324,N_4899);
xor U5972 (N_5972,N_5262,N_5141);
nand U5973 (N_5973,N_5000,N_4961);
xnor U5974 (N_5974,N_4968,N_5037);
nor U5975 (N_5975,N_5162,N_5002);
and U5976 (N_5976,N_5308,N_5061);
nand U5977 (N_5977,N_5003,N_5113);
nand U5978 (N_5978,N_5074,N_4818);
nor U5979 (N_5979,N_5104,N_5255);
or U5980 (N_5980,N_5076,N_5167);
xor U5981 (N_5981,N_5246,N_4987);
xnor U5982 (N_5982,N_4893,N_4897);
nor U5983 (N_5983,N_5217,N_5223);
and U5984 (N_5984,N_5247,N_5278);
xnor U5985 (N_5985,N_5363,N_4881);
xor U5986 (N_5986,N_4890,N_5113);
or U5987 (N_5987,N_5103,N_4928);
nand U5988 (N_5988,N_4995,N_5098);
nor U5989 (N_5989,N_5392,N_5153);
nor U5990 (N_5990,N_4961,N_4957);
xnor U5991 (N_5991,N_5395,N_5266);
nor U5992 (N_5992,N_5360,N_4803);
nand U5993 (N_5993,N_5334,N_5297);
nand U5994 (N_5994,N_5389,N_4980);
nor U5995 (N_5995,N_4834,N_5266);
xor U5996 (N_5996,N_4985,N_5340);
or U5997 (N_5997,N_5068,N_5093);
nand U5998 (N_5998,N_5264,N_5308);
or U5999 (N_5999,N_5379,N_4944);
and U6000 (N_6000,N_5660,N_5912);
or U6001 (N_6001,N_5434,N_5498);
or U6002 (N_6002,N_5693,N_5549);
and U6003 (N_6003,N_5403,N_5503);
or U6004 (N_6004,N_5993,N_5541);
xnor U6005 (N_6005,N_5510,N_5746);
xnor U6006 (N_6006,N_5910,N_5475);
or U6007 (N_6007,N_5633,N_5548);
nor U6008 (N_6008,N_5531,N_5720);
or U6009 (N_6009,N_5597,N_5563);
or U6010 (N_6010,N_5680,N_5905);
and U6011 (N_6011,N_5655,N_5412);
nand U6012 (N_6012,N_5555,N_5585);
and U6013 (N_6013,N_5729,N_5463);
nand U6014 (N_6014,N_5952,N_5895);
and U6015 (N_6015,N_5805,N_5406);
and U6016 (N_6016,N_5817,N_5410);
and U6017 (N_6017,N_5842,N_5962);
or U6018 (N_6018,N_5702,N_5416);
and U6019 (N_6019,N_5981,N_5437);
nand U6020 (N_6020,N_5456,N_5978);
or U6021 (N_6021,N_5886,N_5681);
nand U6022 (N_6022,N_5689,N_5831);
and U6023 (N_6023,N_5879,N_5966);
and U6024 (N_6024,N_5683,N_5770);
nor U6025 (N_6025,N_5652,N_5760);
nand U6026 (N_6026,N_5898,N_5838);
or U6027 (N_6027,N_5989,N_5419);
or U6028 (N_6028,N_5618,N_5421);
nor U6029 (N_6029,N_5947,N_5853);
and U6030 (N_6030,N_5866,N_5765);
and U6031 (N_6031,N_5488,N_5430);
or U6032 (N_6032,N_5581,N_5833);
and U6033 (N_6033,N_5494,N_5502);
xnor U6034 (N_6034,N_5478,N_5659);
xor U6035 (N_6035,N_5967,N_5462);
and U6036 (N_6036,N_5644,N_5663);
and U6037 (N_6037,N_5707,N_5642);
and U6038 (N_6038,N_5742,N_5848);
nor U6039 (N_6039,N_5771,N_5880);
or U6040 (N_6040,N_5767,N_5856);
or U6041 (N_6041,N_5487,N_5933);
xor U6042 (N_6042,N_5684,N_5453);
nand U6043 (N_6043,N_5575,N_5861);
nand U6044 (N_6044,N_5552,N_5534);
and U6045 (N_6045,N_5649,N_5505);
or U6046 (N_6046,N_5669,N_5537);
xnor U6047 (N_6047,N_5839,N_5712);
and U6048 (N_6048,N_5825,N_5677);
nor U6049 (N_6049,N_5553,N_5664);
nor U6050 (N_6050,N_5759,N_5578);
or U6051 (N_6051,N_5977,N_5855);
xnor U6052 (N_6052,N_5885,N_5559);
and U6053 (N_6053,N_5479,N_5927);
xor U6054 (N_6054,N_5971,N_5704);
nand U6055 (N_6055,N_5763,N_5506);
xnor U6056 (N_6056,N_5917,N_5471);
xnor U6057 (N_6057,N_5526,N_5590);
nand U6058 (N_6058,N_5946,N_5938);
nand U6059 (N_6059,N_5661,N_5811);
xnor U6060 (N_6060,N_5774,N_5455);
nand U6061 (N_6061,N_5944,N_5916);
nor U6062 (N_6062,N_5779,N_5647);
xor U6063 (N_6063,N_5605,N_5705);
nor U6064 (N_6064,N_5643,N_5999);
and U6065 (N_6065,N_5539,N_5405);
or U6066 (N_6066,N_5620,N_5940);
xnor U6067 (N_6067,N_5924,N_5925);
or U6068 (N_6068,N_5998,N_5452);
or U6069 (N_6069,N_5586,N_5588);
or U6070 (N_6070,N_5599,N_5903);
xor U6071 (N_6071,N_5454,N_5509);
or U6072 (N_6072,N_5567,N_5963);
nand U6073 (N_6073,N_5570,N_5816);
nor U6074 (N_6074,N_5934,N_5894);
xor U6075 (N_6075,N_5727,N_5573);
or U6076 (N_6076,N_5635,N_5859);
nor U6077 (N_6077,N_5666,N_5854);
nor U6078 (N_6078,N_5422,N_5914);
and U6079 (N_6079,N_5891,N_5769);
and U6080 (N_6080,N_5748,N_5814);
nor U6081 (N_6081,N_5409,N_5810);
nand U6082 (N_6082,N_5423,N_5948);
nor U6083 (N_6083,N_5432,N_5547);
or U6084 (N_6084,N_5992,N_5464);
nor U6085 (N_6085,N_5899,N_5524);
xor U6086 (N_6086,N_5958,N_5561);
nor U6087 (N_6087,N_5577,N_5565);
xor U6088 (N_6088,N_5497,N_5744);
nand U6089 (N_6089,N_5909,N_5717);
or U6090 (N_6090,N_5755,N_5554);
nand U6091 (N_6091,N_5665,N_5809);
or U6092 (N_6092,N_5691,N_5592);
nand U6093 (N_6093,N_5785,N_5844);
nand U6094 (N_6094,N_5822,N_5613);
xor U6095 (N_6095,N_5863,N_5583);
nor U6096 (N_6096,N_5697,N_5733);
or U6097 (N_6097,N_5737,N_5974);
or U6098 (N_6098,N_5686,N_5623);
nor U6099 (N_6099,N_5685,N_5892);
nor U6100 (N_6100,N_5741,N_5429);
and U6101 (N_6101,N_5931,N_5530);
nand U6102 (N_6102,N_5443,N_5657);
or U6103 (N_6103,N_5874,N_5991);
and U6104 (N_6104,N_5493,N_5724);
nor U6105 (N_6105,N_5404,N_5614);
or U6106 (N_6106,N_5504,N_5499);
xnor U6107 (N_6107,N_5602,N_5923);
nor U6108 (N_6108,N_5436,N_5922);
xnor U6109 (N_6109,N_5786,N_5593);
nor U6110 (N_6110,N_5616,N_5511);
and U6111 (N_6111,N_5709,N_5507);
or U6112 (N_6112,N_5641,N_5699);
nand U6113 (N_6113,N_5517,N_5907);
nand U6114 (N_6114,N_5850,N_5735);
nand U6115 (N_6115,N_5569,N_5582);
or U6116 (N_6116,N_5900,N_5890);
nor U6117 (N_6117,N_5734,N_5716);
or U6118 (N_6118,N_5761,N_5519);
xnor U6119 (N_6119,N_5417,N_5965);
and U6120 (N_6120,N_5433,N_5953);
or U6121 (N_6121,N_5489,N_5461);
nor U6122 (N_6122,N_5738,N_5612);
or U6123 (N_6123,N_5609,N_5957);
nor U6124 (N_6124,N_5420,N_5913);
or U6125 (N_6125,N_5472,N_5536);
or U6126 (N_6126,N_5674,N_5596);
or U6127 (N_6127,N_5711,N_5701);
xnor U6128 (N_6128,N_5961,N_5911);
or U6129 (N_6129,N_5440,N_5513);
xor U6130 (N_6130,N_5622,N_5846);
and U6131 (N_6131,N_5402,N_5745);
nor U6132 (N_6132,N_5688,N_5692);
nor U6133 (N_6133,N_5682,N_5673);
nor U6134 (N_6134,N_5869,N_5932);
or U6135 (N_6135,N_5935,N_5439);
or U6136 (N_6136,N_5964,N_5546);
and U6137 (N_6137,N_5544,N_5865);
nor U6138 (N_6138,N_5607,N_5926);
xnor U6139 (N_6139,N_5799,N_5988);
nand U6140 (N_6140,N_5970,N_5984);
and U6141 (N_6141,N_5939,N_5518);
and U6142 (N_6142,N_5749,N_5784);
nand U6143 (N_6143,N_5543,N_5975);
nand U6144 (N_6144,N_5773,N_5972);
nand U6145 (N_6145,N_5813,N_5918);
xor U6146 (N_6146,N_5820,N_5973);
or U6147 (N_6147,N_5696,N_5783);
or U6148 (N_6148,N_5798,N_5941);
and U6149 (N_6149,N_5662,N_5610);
nand U6150 (N_6150,N_5551,N_5654);
xnor U6151 (N_6151,N_5427,N_5750);
xor U6152 (N_6152,N_5426,N_5790);
or U6153 (N_6153,N_5864,N_5802);
and U6154 (N_6154,N_5458,N_5762);
and U6155 (N_6155,N_5851,N_5920);
xor U6156 (N_6156,N_5540,N_5512);
nor U6157 (N_6157,N_5640,N_5449);
nor U6158 (N_6158,N_5778,N_5852);
nor U6159 (N_6159,N_5730,N_5772);
or U6160 (N_6160,N_5606,N_5834);
and U6161 (N_6161,N_5757,N_5447);
xnor U6162 (N_6162,N_5728,N_5884);
or U6163 (N_6163,N_5545,N_5515);
or U6164 (N_6164,N_5603,N_5626);
nor U6165 (N_6165,N_5435,N_5732);
nor U6166 (N_6166,N_5782,N_5400);
or U6167 (N_6167,N_5470,N_5979);
xor U6168 (N_6168,N_5698,N_5801);
xor U6169 (N_6169,N_5803,N_5994);
xnor U6170 (N_6170,N_5928,N_5739);
or U6171 (N_6171,N_5492,N_5841);
and U6172 (N_6172,N_5424,N_5906);
nor U6173 (N_6173,N_5690,N_5714);
or U6174 (N_6174,N_5921,N_5843);
and U6175 (N_6175,N_5983,N_5558);
or U6176 (N_6176,N_5679,N_5904);
nor U6177 (N_6177,N_5639,N_5937);
nand U6178 (N_6178,N_5710,N_5789);
or U6179 (N_6179,N_5700,N_5636);
nor U6180 (N_6180,N_5721,N_5576);
and U6181 (N_6181,N_5878,N_5584);
nor U6182 (N_6182,N_5650,N_5827);
nor U6183 (N_6183,N_5408,N_5457);
or U6184 (N_6184,N_5797,N_5672);
nand U6185 (N_6185,N_5625,N_5431);
xnor U6186 (N_6186,N_5837,N_5791);
xnor U6187 (N_6187,N_5425,N_5758);
or U6188 (N_6188,N_5477,N_5556);
and U6189 (N_6189,N_5560,N_5826);
xnor U6190 (N_6190,N_5413,N_5522);
xor U6191 (N_6191,N_5997,N_5883);
and U6192 (N_6192,N_5954,N_5525);
nand U6193 (N_6193,N_5428,N_5538);
nor U6194 (N_6194,N_5829,N_5753);
nand U6195 (N_6195,N_5571,N_5671);
nand U6196 (N_6196,N_5819,N_5594);
xor U6197 (N_6197,N_5466,N_5959);
and U6198 (N_6198,N_5637,N_5646);
xor U6199 (N_6199,N_5823,N_5670);
nand U6200 (N_6200,N_5668,N_5467);
or U6201 (N_6201,N_5448,N_5960);
or U6202 (N_6202,N_5482,N_5776);
nor U6203 (N_6203,N_5736,N_5870);
and U6204 (N_6204,N_5812,N_5876);
nor U6205 (N_6205,N_5486,N_5821);
and U6206 (N_6206,N_5579,N_5747);
nand U6207 (N_6207,N_5630,N_5523);
nor U6208 (N_6208,N_5562,N_5469);
and U6209 (N_6209,N_5580,N_5754);
xor U6210 (N_6210,N_5777,N_5535);
nand U6211 (N_6211,N_5514,N_5807);
or U6212 (N_6212,N_5788,N_5632);
or U6213 (N_6213,N_5678,N_5676);
and U6214 (N_6214,N_5627,N_5550);
and U6215 (N_6215,N_5990,N_5756);
xor U6216 (N_6216,N_5713,N_5780);
or U6217 (N_6217,N_5490,N_5631);
and U6218 (N_6218,N_5945,N_5715);
nor U6219 (N_6219,N_5653,N_5695);
nand U6220 (N_6220,N_5694,N_5615);
and U6221 (N_6221,N_5868,N_5706);
nand U6222 (N_6222,N_5996,N_5459);
or U6223 (N_6223,N_5484,N_5589);
nor U6224 (N_6224,N_5687,N_5415);
nand U6225 (N_6225,N_5942,N_5896);
nand U6226 (N_6226,N_5815,N_5985);
nand U6227 (N_6227,N_5617,N_5845);
nand U6228 (N_6228,N_5450,N_5474);
xnor U6229 (N_6229,N_5438,N_5766);
nand U6230 (N_6230,N_5483,N_5619);
and U6231 (N_6231,N_5794,N_5658);
nor U6232 (N_6232,N_5743,N_5800);
nand U6233 (N_6233,N_5862,N_5595);
nor U6234 (N_6234,N_5611,N_5723);
or U6235 (N_6235,N_5407,N_5930);
and U6236 (N_6236,N_5476,N_5516);
and U6237 (N_6237,N_5726,N_5951);
nor U6238 (N_6238,N_5792,N_5528);
xnor U6239 (N_6239,N_5598,N_5496);
or U6240 (N_6240,N_5529,N_5401);
nor U6241 (N_6241,N_5835,N_5468);
or U6242 (N_6242,N_5882,N_5969);
nor U6243 (N_6243,N_5987,N_5830);
xor U6244 (N_6244,N_5929,N_5719);
and U6245 (N_6245,N_5446,N_5849);
xnor U6246 (N_6246,N_5718,N_5955);
nor U6247 (N_6247,N_5956,N_5441);
or U6248 (N_6248,N_5444,N_5840);
nor U6249 (N_6249,N_5520,N_5638);
nor U6250 (N_6250,N_5949,N_5731);
nand U6251 (N_6251,N_5950,N_5936);
nor U6252 (N_6252,N_5445,N_5465);
or U6253 (N_6253,N_5752,N_5703);
nand U6254 (N_6254,N_5836,N_5473);
nor U6255 (N_6255,N_5451,N_5889);
or U6256 (N_6256,N_5624,N_5600);
or U6257 (N_6257,N_5793,N_5656);
xnor U6258 (N_6258,N_5873,N_5881);
xnor U6259 (N_6259,N_5872,N_5982);
xnor U6260 (N_6260,N_5867,N_5976);
nand U6261 (N_6261,N_5485,N_5574);
xnor U6262 (N_6262,N_5414,N_5521);
nand U6263 (N_6263,N_5564,N_5858);
or U6264 (N_6264,N_5888,N_5568);
xor U6265 (N_6265,N_5501,N_5943);
xnor U6266 (N_6266,N_5725,N_5919);
nand U6267 (N_6267,N_5787,N_5557);
or U6268 (N_6268,N_5628,N_5795);
or U6269 (N_6269,N_5897,N_5818);
nor U6270 (N_6270,N_5418,N_5781);
or U6271 (N_6271,N_5481,N_5480);
nor U6272 (N_6272,N_5740,N_5621);
nor U6273 (N_6273,N_5495,N_5893);
nand U6274 (N_6274,N_5645,N_5591);
nor U6275 (N_6275,N_5722,N_5491);
nand U6276 (N_6276,N_5648,N_5608);
and U6277 (N_6277,N_5601,N_5877);
or U6278 (N_6278,N_5667,N_5871);
and U6279 (N_6279,N_5986,N_5411);
nand U6280 (N_6280,N_5908,N_5804);
nand U6281 (N_6281,N_5968,N_5572);
nand U6282 (N_6282,N_5651,N_5542);
and U6283 (N_6283,N_5847,N_5824);
or U6284 (N_6284,N_5533,N_5751);
or U6285 (N_6285,N_5566,N_5675);
nor U6286 (N_6286,N_5527,N_5860);
nand U6287 (N_6287,N_5901,N_5460);
nand U6288 (N_6288,N_5980,N_5764);
nand U6289 (N_6289,N_5587,N_5708);
nand U6290 (N_6290,N_5500,N_5796);
or U6291 (N_6291,N_5768,N_5806);
nor U6292 (N_6292,N_5775,N_5857);
xor U6293 (N_6293,N_5532,N_5604);
nor U6294 (N_6294,N_5887,N_5875);
nand U6295 (N_6295,N_5995,N_5634);
nand U6296 (N_6296,N_5629,N_5902);
or U6297 (N_6297,N_5832,N_5442);
nand U6298 (N_6298,N_5808,N_5915);
or U6299 (N_6299,N_5508,N_5828);
nor U6300 (N_6300,N_5710,N_5411);
nand U6301 (N_6301,N_5517,N_5928);
and U6302 (N_6302,N_5931,N_5978);
nor U6303 (N_6303,N_5959,N_5560);
nand U6304 (N_6304,N_5481,N_5694);
xnor U6305 (N_6305,N_5618,N_5499);
or U6306 (N_6306,N_5896,N_5826);
xor U6307 (N_6307,N_5865,N_5870);
or U6308 (N_6308,N_5916,N_5536);
xor U6309 (N_6309,N_5655,N_5939);
nor U6310 (N_6310,N_5822,N_5785);
and U6311 (N_6311,N_5781,N_5434);
and U6312 (N_6312,N_5968,N_5481);
and U6313 (N_6313,N_5916,N_5572);
and U6314 (N_6314,N_5564,N_5631);
nand U6315 (N_6315,N_5965,N_5501);
and U6316 (N_6316,N_5429,N_5742);
nand U6317 (N_6317,N_5841,N_5461);
nand U6318 (N_6318,N_5406,N_5861);
nand U6319 (N_6319,N_5628,N_5983);
nor U6320 (N_6320,N_5914,N_5424);
nor U6321 (N_6321,N_5414,N_5547);
xor U6322 (N_6322,N_5543,N_5951);
xor U6323 (N_6323,N_5680,N_5431);
nand U6324 (N_6324,N_5545,N_5479);
xor U6325 (N_6325,N_5873,N_5898);
nor U6326 (N_6326,N_5594,N_5530);
nand U6327 (N_6327,N_5634,N_5818);
or U6328 (N_6328,N_5909,N_5498);
nor U6329 (N_6329,N_5908,N_5521);
nor U6330 (N_6330,N_5892,N_5565);
nand U6331 (N_6331,N_5507,N_5856);
nand U6332 (N_6332,N_5612,N_5865);
xor U6333 (N_6333,N_5503,N_5890);
or U6334 (N_6334,N_5636,N_5821);
nand U6335 (N_6335,N_5882,N_5998);
nor U6336 (N_6336,N_5610,N_5812);
or U6337 (N_6337,N_5721,N_5583);
and U6338 (N_6338,N_5779,N_5943);
and U6339 (N_6339,N_5797,N_5537);
or U6340 (N_6340,N_5738,N_5770);
and U6341 (N_6341,N_5913,N_5523);
or U6342 (N_6342,N_5905,N_5778);
nand U6343 (N_6343,N_5749,N_5954);
nor U6344 (N_6344,N_5911,N_5663);
or U6345 (N_6345,N_5736,N_5430);
xor U6346 (N_6346,N_5423,N_5700);
nand U6347 (N_6347,N_5770,N_5784);
xor U6348 (N_6348,N_5489,N_5965);
or U6349 (N_6349,N_5831,N_5497);
xnor U6350 (N_6350,N_5813,N_5929);
xnor U6351 (N_6351,N_5987,N_5562);
xnor U6352 (N_6352,N_5681,N_5571);
xor U6353 (N_6353,N_5704,N_5465);
or U6354 (N_6354,N_5996,N_5488);
and U6355 (N_6355,N_5449,N_5731);
nand U6356 (N_6356,N_5526,N_5681);
and U6357 (N_6357,N_5783,N_5416);
and U6358 (N_6358,N_5599,N_5944);
and U6359 (N_6359,N_5606,N_5465);
nor U6360 (N_6360,N_5826,N_5773);
nand U6361 (N_6361,N_5898,N_5673);
nor U6362 (N_6362,N_5747,N_5651);
nor U6363 (N_6363,N_5608,N_5944);
or U6364 (N_6364,N_5628,N_5954);
and U6365 (N_6365,N_5507,N_5590);
or U6366 (N_6366,N_5925,N_5652);
nand U6367 (N_6367,N_5594,N_5983);
nand U6368 (N_6368,N_5796,N_5719);
nor U6369 (N_6369,N_5651,N_5870);
nand U6370 (N_6370,N_5749,N_5593);
and U6371 (N_6371,N_5707,N_5812);
nor U6372 (N_6372,N_5556,N_5882);
and U6373 (N_6373,N_5878,N_5583);
and U6374 (N_6374,N_5528,N_5771);
xor U6375 (N_6375,N_5462,N_5789);
nand U6376 (N_6376,N_5952,N_5433);
and U6377 (N_6377,N_5601,N_5438);
and U6378 (N_6378,N_5770,N_5736);
and U6379 (N_6379,N_5537,N_5874);
and U6380 (N_6380,N_5418,N_5463);
or U6381 (N_6381,N_5564,N_5957);
or U6382 (N_6382,N_5401,N_5839);
or U6383 (N_6383,N_5788,N_5533);
xnor U6384 (N_6384,N_5851,N_5957);
nor U6385 (N_6385,N_5982,N_5874);
or U6386 (N_6386,N_5834,N_5740);
and U6387 (N_6387,N_5797,N_5470);
nand U6388 (N_6388,N_5931,N_5944);
or U6389 (N_6389,N_5883,N_5956);
xor U6390 (N_6390,N_5851,N_5600);
xnor U6391 (N_6391,N_5824,N_5584);
or U6392 (N_6392,N_5681,N_5486);
or U6393 (N_6393,N_5825,N_5799);
and U6394 (N_6394,N_5665,N_5534);
nand U6395 (N_6395,N_5842,N_5520);
or U6396 (N_6396,N_5709,N_5894);
nor U6397 (N_6397,N_5472,N_5473);
nor U6398 (N_6398,N_5686,N_5672);
and U6399 (N_6399,N_5642,N_5687);
nand U6400 (N_6400,N_5753,N_5552);
or U6401 (N_6401,N_5754,N_5922);
xnor U6402 (N_6402,N_5450,N_5637);
and U6403 (N_6403,N_5405,N_5802);
or U6404 (N_6404,N_5405,N_5860);
nor U6405 (N_6405,N_5684,N_5558);
or U6406 (N_6406,N_5487,N_5881);
nand U6407 (N_6407,N_5403,N_5690);
nand U6408 (N_6408,N_5892,N_5590);
and U6409 (N_6409,N_5429,N_5521);
nor U6410 (N_6410,N_5519,N_5825);
nor U6411 (N_6411,N_5997,N_5977);
xor U6412 (N_6412,N_5650,N_5627);
nor U6413 (N_6413,N_5728,N_5708);
and U6414 (N_6414,N_5600,N_5651);
xor U6415 (N_6415,N_5735,N_5793);
nor U6416 (N_6416,N_5463,N_5976);
xnor U6417 (N_6417,N_5847,N_5535);
nor U6418 (N_6418,N_5603,N_5414);
xnor U6419 (N_6419,N_5478,N_5972);
nor U6420 (N_6420,N_5405,N_5799);
or U6421 (N_6421,N_5999,N_5405);
xnor U6422 (N_6422,N_5910,N_5999);
nor U6423 (N_6423,N_5751,N_5604);
and U6424 (N_6424,N_5578,N_5440);
nor U6425 (N_6425,N_5916,N_5810);
nor U6426 (N_6426,N_5448,N_5548);
nand U6427 (N_6427,N_5974,N_5758);
nand U6428 (N_6428,N_5848,N_5403);
or U6429 (N_6429,N_5805,N_5563);
nor U6430 (N_6430,N_5818,N_5433);
xnor U6431 (N_6431,N_5425,N_5619);
nand U6432 (N_6432,N_5863,N_5758);
nand U6433 (N_6433,N_5957,N_5427);
nand U6434 (N_6434,N_5618,N_5446);
xnor U6435 (N_6435,N_5523,N_5841);
nor U6436 (N_6436,N_5958,N_5606);
xor U6437 (N_6437,N_5994,N_5622);
and U6438 (N_6438,N_5413,N_5868);
xor U6439 (N_6439,N_5502,N_5436);
nand U6440 (N_6440,N_5621,N_5696);
nand U6441 (N_6441,N_5966,N_5932);
nand U6442 (N_6442,N_5554,N_5542);
nor U6443 (N_6443,N_5995,N_5815);
nor U6444 (N_6444,N_5637,N_5869);
nor U6445 (N_6445,N_5644,N_5600);
nand U6446 (N_6446,N_5968,N_5551);
nand U6447 (N_6447,N_5555,N_5536);
and U6448 (N_6448,N_5585,N_5441);
and U6449 (N_6449,N_5660,N_5656);
and U6450 (N_6450,N_5424,N_5504);
xnor U6451 (N_6451,N_5774,N_5867);
and U6452 (N_6452,N_5828,N_5553);
nor U6453 (N_6453,N_5452,N_5885);
and U6454 (N_6454,N_5623,N_5809);
and U6455 (N_6455,N_5805,N_5870);
or U6456 (N_6456,N_5668,N_5772);
xor U6457 (N_6457,N_5988,N_5648);
nand U6458 (N_6458,N_5911,N_5493);
and U6459 (N_6459,N_5700,N_5877);
nor U6460 (N_6460,N_5481,N_5451);
nor U6461 (N_6461,N_5432,N_5441);
and U6462 (N_6462,N_5747,N_5813);
xnor U6463 (N_6463,N_5588,N_5844);
xor U6464 (N_6464,N_5988,N_5907);
and U6465 (N_6465,N_5999,N_5922);
xor U6466 (N_6466,N_5783,N_5550);
nand U6467 (N_6467,N_5886,N_5704);
nand U6468 (N_6468,N_5414,N_5435);
nor U6469 (N_6469,N_5668,N_5538);
nand U6470 (N_6470,N_5602,N_5927);
xnor U6471 (N_6471,N_5803,N_5556);
nor U6472 (N_6472,N_5612,N_5773);
nor U6473 (N_6473,N_5629,N_5863);
xor U6474 (N_6474,N_5662,N_5904);
nand U6475 (N_6475,N_5728,N_5477);
and U6476 (N_6476,N_5646,N_5870);
or U6477 (N_6477,N_5653,N_5412);
nand U6478 (N_6478,N_5423,N_5882);
nand U6479 (N_6479,N_5790,N_5887);
nand U6480 (N_6480,N_5949,N_5606);
or U6481 (N_6481,N_5668,N_5440);
nand U6482 (N_6482,N_5572,N_5664);
xor U6483 (N_6483,N_5804,N_5727);
nor U6484 (N_6484,N_5582,N_5520);
or U6485 (N_6485,N_5591,N_5793);
or U6486 (N_6486,N_5787,N_5494);
and U6487 (N_6487,N_5952,N_5458);
nand U6488 (N_6488,N_5759,N_5508);
nor U6489 (N_6489,N_5552,N_5471);
and U6490 (N_6490,N_5985,N_5770);
nand U6491 (N_6491,N_5739,N_5943);
nor U6492 (N_6492,N_5401,N_5547);
and U6493 (N_6493,N_5592,N_5913);
nand U6494 (N_6494,N_5984,N_5640);
nor U6495 (N_6495,N_5437,N_5936);
and U6496 (N_6496,N_5926,N_5752);
nor U6497 (N_6497,N_5935,N_5487);
nand U6498 (N_6498,N_5985,N_5786);
or U6499 (N_6499,N_5652,N_5771);
or U6500 (N_6500,N_5715,N_5813);
nor U6501 (N_6501,N_5649,N_5906);
nor U6502 (N_6502,N_5802,N_5460);
nand U6503 (N_6503,N_5731,N_5846);
xnor U6504 (N_6504,N_5827,N_5746);
nand U6505 (N_6505,N_5555,N_5609);
nor U6506 (N_6506,N_5491,N_5555);
and U6507 (N_6507,N_5842,N_5408);
nand U6508 (N_6508,N_5676,N_5992);
or U6509 (N_6509,N_5762,N_5989);
or U6510 (N_6510,N_5668,N_5963);
xnor U6511 (N_6511,N_5855,N_5416);
nand U6512 (N_6512,N_5480,N_5802);
or U6513 (N_6513,N_5619,N_5781);
and U6514 (N_6514,N_5618,N_5969);
or U6515 (N_6515,N_5415,N_5681);
xor U6516 (N_6516,N_5611,N_5963);
nor U6517 (N_6517,N_5482,N_5680);
nor U6518 (N_6518,N_5852,N_5424);
and U6519 (N_6519,N_5425,N_5801);
xnor U6520 (N_6520,N_5431,N_5726);
nor U6521 (N_6521,N_5754,N_5623);
nor U6522 (N_6522,N_5579,N_5569);
xor U6523 (N_6523,N_5912,N_5798);
nor U6524 (N_6524,N_5679,N_5515);
nand U6525 (N_6525,N_5427,N_5888);
or U6526 (N_6526,N_5902,N_5503);
nand U6527 (N_6527,N_5695,N_5801);
nand U6528 (N_6528,N_5509,N_5812);
and U6529 (N_6529,N_5996,N_5833);
nor U6530 (N_6530,N_5792,N_5978);
or U6531 (N_6531,N_5779,N_5841);
xnor U6532 (N_6532,N_5588,N_5830);
and U6533 (N_6533,N_5586,N_5904);
and U6534 (N_6534,N_5718,N_5934);
xnor U6535 (N_6535,N_5606,N_5513);
nand U6536 (N_6536,N_5446,N_5761);
and U6537 (N_6537,N_5549,N_5556);
nor U6538 (N_6538,N_5810,N_5992);
or U6539 (N_6539,N_5650,N_5978);
or U6540 (N_6540,N_5849,N_5905);
and U6541 (N_6541,N_5456,N_5804);
or U6542 (N_6542,N_5685,N_5806);
and U6543 (N_6543,N_5406,N_5602);
xnor U6544 (N_6544,N_5627,N_5871);
nor U6545 (N_6545,N_5796,N_5861);
nand U6546 (N_6546,N_5663,N_5650);
xor U6547 (N_6547,N_5458,N_5935);
xnor U6548 (N_6548,N_5745,N_5486);
and U6549 (N_6549,N_5627,N_5534);
nand U6550 (N_6550,N_5987,N_5938);
nor U6551 (N_6551,N_5922,N_5847);
nor U6552 (N_6552,N_5919,N_5743);
or U6553 (N_6553,N_5847,N_5756);
and U6554 (N_6554,N_5655,N_5468);
xnor U6555 (N_6555,N_5500,N_5942);
or U6556 (N_6556,N_5941,N_5502);
nor U6557 (N_6557,N_5733,N_5584);
nor U6558 (N_6558,N_5936,N_5843);
or U6559 (N_6559,N_5482,N_5892);
xnor U6560 (N_6560,N_5454,N_5491);
xnor U6561 (N_6561,N_5737,N_5812);
xor U6562 (N_6562,N_5498,N_5700);
nor U6563 (N_6563,N_5501,N_5782);
and U6564 (N_6564,N_5848,N_5729);
xor U6565 (N_6565,N_5546,N_5857);
and U6566 (N_6566,N_5607,N_5747);
nand U6567 (N_6567,N_5470,N_5929);
nand U6568 (N_6568,N_5894,N_5441);
nor U6569 (N_6569,N_5921,N_5419);
and U6570 (N_6570,N_5995,N_5861);
or U6571 (N_6571,N_5907,N_5755);
and U6572 (N_6572,N_5529,N_5776);
and U6573 (N_6573,N_5775,N_5446);
xnor U6574 (N_6574,N_5498,N_5787);
or U6575 (N_6575,N_5948,N_5426);
nor U6576 (N_6576,N_5860,N_5809);
and U6577 (N_6577,N_5496,N_5476);
or U6578 (N_6578,N_5511,N_5932);
nand U6579 (N_6579,N_5499,N_5434);
xnor U6580 (N_6580,N_5558,N_5799);
or U6581 (N_6581,N_5529,N_5819);
or U6582 (N_6582,N_5532,N_5971);
or U6583 (N_6583,N_5402,N_5852);
xnor U6584 (N_6584,N_5566,N_5694);
nand U6585 (N_6585,N_5796,N_5476);
xnor U6586 (N_6586,N_5961,N_5898);
xor U6587 (N_6587,N_5535,N_5812);
and U6588 (N_6588,N_5809,N_5821);
nor U6589 (N_6589,N_5640,N_5646);
or U6590 (N_6590,N_5929,N_5915);
and U6591 (N_6591,N_5697,N_5589);
nor U6592 (N_6592,N_5441,N_5733);
nand U6593 (N_6593,N_5563,N_5915);
xor U6594 (N_6594,N_5788,N_5733);
and U6595 (N_6595,N_5517,N_5778);
and U6596 (N_6596,N_5802,N_5926);
nor U6597 (N_6597,N_5405,N_5655);
nand U6598 (N_6598,N_5535,N_5576);
or U6599 (N_6599,N_5944,N_5871);
and U6600 (N_6600,N_6076,N_6400);
or U6601 (N_6601,N_6377,N_6468);
xor U6602 (N_6602,N_6219,N_6385);
xnor U6603 (N_6603,N_6574,N_6101);
xnor U6604 (N_6604,N_6397,N_6163);
nand U6605 (N_6605,N_6159,N_6124);
and U6606 (N_6606,N_6207,N_6316);
nand U6607 (N_6607,N_6596,N_6266);
nor U6608 (N_6608,N_6452,N_6012);
or U6609 (N_6609,N_6195,N_6418);
xor U6610 (N_6610,N_6017,N_6551);
nor U6611 (N_6611,N_6188,N_6431);
nand U6612 (N_6612,N_6319,N_6057);
and U6613 (N_6613,N_6194,N_6429);
nor U6614 (N_6614,N_6486,N_6090);
nand U6615 (N_6615,N_6364,N_6407);
nor U6616 (N_6616,N_6306,N_6558);
or U6617 (N_6617,N_6153,N_6465);
or U6618 (N_6618,N_6568,N_6318);
and U6619 (N_6619,N_6544,N_6144);
or U6620 (N_6620,N_6487,N_6136);
and U6621 (N_6621,N_6506,N_6478);
xor U6622 (N_6622,N_6118,N_6193);
nand U6623 (N_6623,N_6001,N_6222);
or U6624 (N_6624,N_6126,N_6489);
nor U6625 (N_6625,N_6029,N_6360);
xnor U6626 (N_6626,N_6192,N_6132);
or U6627 (N_6627,N_6223,N_6511);
and U6628 (N_6628,N_6184,N_6295);
nand U6629 (N_6629,N_6236,N_6448);
xor U6630 (N_6630,N_6515,N_6432);
and U6631 (N_6631,N_6592,N_6462);
or U6632 (N_6632,N_6459,N_6538);
nor U6633 (N_6633,N_6066,N_6503);
nand U6634 (N_6634,N_6567,N_6243);
or U6635 (N_6635,N_6372,N_6393);
xnor U6636 (N_6636,N_6036,N_6447);
or U6637 (N_6637,N_6548,N_6082);
nand U6638 (N_6638,N_6226,N_6518);
and U6639 (N_6639,N_6024,N_6004);
or U6640 (N_6640,N_6209,N_6214);
and U6641 (N_6641,N_6181,N_6552);
and U6642 (N_6642,N_6414,N_6026);
nand U6643 (N_6643,N_6191,N_6321);
xnor U6644 (N_6644,N_6399,N_6485);
or U6645 (N_6645,N_6002,N_6178);
nand U6646 (N_6646,N_6204,N_6235);
or U6647 (N_6647,N_6030,N_6573);
or U6648 (N_6648,N_6111,N_6237);
or U6649 (N_6649,N_6115,N_6028);
nand U6650 (N_6650,N_6096,N_6304);
nand U6651 (N_6651,N_6249,N_6562);
or U6652 (N_6652,N_6083,N_6412);
and U6653 (N_6653,N_6559,N_6196);
and U6654 (N_6654,N_6234,N_6541);
and U6655 (N_6655,N_6311,N_6247);
nor U6656 (N_6656,N_6441,N_6182);
or U6657 (N_6657,N_6152,N_6477);
or U6658 (N_6658,N_6370,N_6583);
nand U6659 (N_6659,N_6167,N_6157);
and U6660 (N_6660,N_6492,N_6406);
xor U6661 (N_6661,N_6109,N_6077);
xor U6662 (N_6662,N_6050,N_6164);
nor U6663 (N_6663,N_6320,N_6451);
nand U6664 (N_6664,N_6179,N_6035);
xnor U6665 (N_6665,N_6070,N_6476);
nand U6666 (N_6666,N_6245,N_6392);
or U6667 (N_6667,N_6206,N_6225);
nand U6668 (N_6668,N_6282,N_6174);
nor U6669 (N_6669,N_6381,N_6241);
nand U6670 (N_6670,N_6228,N_6430);
nor U6671 (N_6671,N_6527,N_6122);
and U6672 (N_6672,N_6327,N_6287);
nand U6673 (N_6673,N_6442,N_6127);
nor U6674 (N_6674,N_6580,N_6051);
or U6675 (N_6675,N_6339,N_6540);
nor U6676 (N_6676,N_6497,N_6061);
or U6677 (N_6677,N_6239,N_6461);
or U6678 (N_6678,N_6481,N_6526);
and U6679 (N_6679,N_6524,N_6137);
nand U6680 (N_6680,N_6274,N_6114);
and U6681 (N_6681,N_6064,N_6175);
nor U6682 (N_6682,N_6123,N_6220);
and U6683 (N_6683,N_6217,N_6269);
or U6684 (N_6684,N_6043,N_6420);
nor U6685 (N_6685,N_6322,N_6224);
xnor U6686 (N_6686,N_6308,N_6215);
nor U6687 (N_6687,N_6480,N_6584);
xnor U6688 (N_6688,N_6532,N_6590);
nor U6689 (N_6689,N_6436,N_6065);
nor U6690 (N_6690,N_6367,N_6099);
and U6691 (N_6691,N_6404,N_6071);
xor U6692 (N_6692,N_6398,N_6208);
and U6693 (N_6693,N_6309,N_6464);
or U6694 (N_6694,N_6593,N_6265);
and U6695 (N_6695,N_6203,N_6286);
xor U6696 (N_6696,N_6354,N_6294);
and U6697 (N_6697,N_6351,N_6120);
or U6698 (N_6698,N_6458,N_6263);
or U6699 (N_6699,N_6095,N_6353);
and U6700 (N_6700,N_6015,N_6113);
nand U6701 (N_6701,N_6105,N_6554);
and U6702 (N_6702,N_6572,N_6210);
or U6703 (N_6703,N_6500,N_6453);
or U6704 (N_6704,N_6484,N_6068);
nand U6705 (N_6705,N_6373,N_6074);
nand U6706 (N_6706,N_6110,N_6508);
and U6707 (N_6707,N_6359,N_6437);
and U6708 (N_6708,N_6557,N_6097);
or U6709 (N_6709,N_6504,N_6314);
or U6710 (N_6710,N_6063,N_6374);
nor U6711 (N_6711,N_6577,N_6255);
and U6712 (N_6712,N_6421,N_6289);
or U6713 (N_6713,N_6342,N_6084);
nand U6714 (N_6714,N_6450,N_6575);
nor U6715 (N_6715,N_6387,N_6542);
or U6716 (N_6716,N_6034,N_6537);
or U6717 (N_6717,N_6280,N_6176);
nand U6718 (N_6718,N_6394,N_6025);
nand U6719 (N_6719,N_6530,N_6042);
nand U6720 (N_6720,N_6325,N_6018);
and U6721 (N_6721,N_6116,N_6067);
nand U6722 (N_6722,N_6037,N_6102);
and U6723 (N_6723,N_6128,N_6479);
nor U6724 (N_6724,N_6131,N_6368);
nor U6725 (N_6725,N_6470,N_6356);
nand U6726 (N_6726,N_6343,N_6324);
nand U6727 (N_6727,N_6014,N_6560);
and U6728 (N_6728,N_6300,N_6233);
or U6729 (N_6729,N_6160,N_6463);
or U6730 (N_6730,N_6089,N_6005);
nand U6731 (N_6731,N_6579,N_6296);
nand U6732 (N_6732,N_6338,N_6553);
or U6733 (N_6733,N_6080,N_6169);
and U6734 (N_6734,N_6232,N_6361);
and U6735 (N_6735,N_6516,N_6410);
xor U6736 (N_6736,N_6121,N_6041);
nor U6737 (N_6737,N_6297,N_6349);
nor U6738 (N_6738,N_6509,N_6049);
nand U6739 (N_6739,N_6257,N_6594);
and U6740 (N_6740,N_6020,N_6161);
xor U6741 (N_6741,N_6514,N_6039);
xnor U6742 (N_6742,N_6048,N_6307);
nor U6743 (N_6743,N_6455,N_6352);
or U6744 (N_6744,N_6107,N_6130);
nor U6745 (N_6745,N_6268,N_6411);
and U6746 (N_6746,N_6366,N_6202);
nor U6747 (N_6747,N_6299,N_6386);
and U6748 (N_6748,N_6000,N_6417);
xor U6749 (N_6749,N_6317,N_6438);
xnor U6750 (N_6750,N_6329,N_6185);
and U6751 (N_6751,N_6402,N_6545);
and U6752 (N_6752,N_6469,N_6434);
or U6753 (N_6753,N_6326,N_6413);
and U6754 (N_6754,N_6170,N_6578);
nand U6755 (N_6755,N_6473,N_6143);
nand U6756 (N_6756,N_6347,N_6081);
and U6757 (N_6757,N_6059,N_6357);
and U6758 (N_6758,N_6595,N_6403);
or U6759 (N_6759,N_6507,N_6079);
nor U6760 (N_6760,N_6426,N_6363);
or U6761 (N_6761,N_6145,N_6288);
nor U6762 (N_6762,N_6585,N_6382);
nor U6763 (N_6763,N_6493,N_6301);
or U6764 (N_6764,N_6396,N_6173);
and U6765 (N_6765,N_6358,N_6279);
xor U6766 (N_6766,N_6488,N_6046);
and U6767 (N_6767,N_6419,N_6284);
or U6768 (N_6768,N_6088,N_6180);
and U6769 (N_6769,N_6154,N_6103);
xnor U6770 (N_6770,N_6440,N_6531);
nand U6771 (N_6771,N_6401,N_6369);
nand U6772 (N_6772,N_6533,N_6589);
and U6773 (N_6773,N_6148,N_6058);
and U6774 (N_6774,N_6547,N_6543);
or U6775 (N_6775,N_6264,N_6038);
nor U6776 (N_6776,N_6275,N_6561);
xnor U6777 (N_6777,N_6555,N_6460);
xor U6778 (N_6778,N_6529,N_6104);
and U6779 (N_6779,N_6528,N_6588);
nand U6780 (N_6780,N_6213,N_6494);
and U6781 (N_6781,N_6045,N_6201);
or U6782 (N_6782,N_6582,N_6383);
and U6783 (N_6783,N_6415,N_6505);
xnor U6784 (N_6784,N_6525,N_6456);
or U6785 (N_6785,N_6272,N_6569);
and U6786 (N_6786,N_6108,N_6491);
nor U6787 (N_6787,N_6521,N_6564);
nand U6788 (N_6788,N_6337,N_6200);
and U6789 (N_6789,N_6599,N_6230);
xnor U6790 (N_6790,N_6252,N_6134);
nor U6791 (N_6791,N_6032,N_6549);
nor U6792 (N_6792,N_6502,N_6416);
xor U6793 (N_6793,N_6365,N_6053);
or U6794 (N_6794,N_6348,N_6454);
xor U6795 (N_6795,N_6016,N_6187);
xor U6796 (N_6796,N_6172,N_6119);
and U6797 (N_6797,N_6586,N_6250);
nand U6798 (N_6798,N_6011,N_6427);
nor U6799 (N_6799,N_6008,N_6085);
nor U6800 (N_6800,N_6443,N_6146);
nand U6801 (N_6801,N_6267,N_6093);
nor U6802 (N_6802,N_6242,N_6536);
nand U6803 (N_6803,N_6092,N_6023);
nor U6804 (N_6804,N_6422,N_6168);
and U6805 (N_6805,N_6598,N_6229);
xor U6806 (N_6806,N_6581,N_6186);
xor U6807 (N_6807,N_6190,N_6331);
xnor U6808 (N_6808,N_6371,N_6444);
nand U6809 (N_6809,N_6133,N_6240);
xor U6810 (N_6810,N_6138,N_6490);
nand U6811 (N_6811,N_6376,N_6091);
and U6812 (N_6812,N_6171,N_6117);
nor U6813 (N_6813,N_6409,N_6060);
and U6814 (N_6814,N_6312,N_6062);
nor U6815 (N_6815,N_6391,N_6519);
and U6816 (N_6816,N_6587,N_6424);
nor U6817 (N_6817,N_6405,N_6248);
nand U6818 (N_6818,N_6052,N_6199);
or U6819 (N_6819,N_6475,N_6147);
nand U6820 (N_6820,N_6205,N_6135);
xnor U6821 (N_6821,N_6256,N_6495);
xor U6822 (N_6822,N_6498,N_6428);
nand U6823 (N_6823,N_6010,N_6198);
or U6824 (N_6824,N_6512,N_6474);
or U6825 (N_6825,N_6335,N_6260);
and U6826 (N_6826,N_6216,N_6534);
and U6827 (N_6827,N_6140,N_6466);
and U6828 (N_6828,N_6341,N_6069);
nor U6829 (N_6829,N_6566,N_6094);
nand U6830 (N_6830,N_6022,N_6246);
and U6831 (N_6831,N_6496,N_6162);
and U6832 (N_6832,N_6482,N_6183);
or U6833 (N_6833,N_6330,N_6323);
nor U6834 (N_6834,N_6513,N_6254);
xor U6835 (N_6835,N_6375,N_6563);
or U6836 (N_6836,N_6336,N_6379);
or U6837 (N_6837,N_6021,N_6253);
or U6838 (N_6838,N_6238,N_6395);
or U6839 (N_6839,N_6100,N_6449);
nor U6840 (N_6840,N_6259,N_6125);
nand U6841 (N_6841,N_6078,N_6003);
nand U6842 (N_6842,N_6425,N_6344);
or U6843 (N_6843,N_6106,N_6310);
and U6844 (N_6844,N_6539,N_6556);
nand U6845 (N_6845,N_6546,N_6087);
or U6846 (N_6846,N_6522,N_6298);
or U6847 (N_6847,N_6273,N_6047);
nand U6848 (N_6848,N_6292,N_6283);
or U6849 (N_6849,N_6340,N_6073);
nor U6850 (N_6850,N_6328,N_6510);
nor U6851 (N_6851,N_6333,N_6390);
or U6852 (N_6852,N_6345,N_6293);
or U6853 (N_6853,N_6197,N_6520);
and U6854 (N_6854,N_6027,N_6302);
nor U6855 (N_6855,N_6378,N_6211);
nand U6856 (N_6856,N_6007,N_6278);
nand U6857 (N_6857,N_6501,N_6571);
xnor U6858 (N_6858,N_6231,N_6218);
xnor U6859 (N_6859,N_6550,N_6389);
nor U6860 (N_6860,N_6086,N_6156);
and U6861 (N_6861,N_6150,N_6221);
nand U6862 (N_6862,N_6006,N_6499);
nor U6863 (N_6863,N_6346,N_6570);
or U6864 (N_6864,N_6313,N_6472);
nand U6865 (N_6865,N_6408,N_6139);
xor U6866 (N_6866,N_6446,N_6565);
xnor U6867 (N_6867,N_6433,N_6129);
nor U6868 (N_6868,N_6388,N_6523);
nand U6869 (N_6869,N_6166,N_6155);
and U6870 (N_6870,N_6165,N_6467);
and U6871 (N_6871,N_6350,N_6013);
xnor U6872 (N_6872,N_6056,N_6270);
and U6873 (N_6873,N_6141,N_6040);
nand U6874 (N_6874,N_6142,N_6044);
or U6875 (N_6875,N_6576,N_6291);
or U6876 (N_6876,N_6303,N_6019);
xnor U6877 (N_6877,N_6535,N_6212);
nand U6878 (N_6878,N_6031,N_6277);
xor U6879 (N_6879,N_6072,N_6597);
and U6880 (N_6880,N_6380,N_6075);
xor U6881 (N_6881,N_6362,N_6457);
nand U6882 (N_6882,N_6244,N_6009);
or U6883 (N_6883,N_6276,N_6334);
nor U6884 (N_6884,N_6251,N_6384);
nand U6885 (N_6885,N_6517,N_6055);
nor U6886 (N_6886,N_6112,N_6355);
nand U6887 (N_6887,N_6262,N_6290);
or U6888 (N_6888,N_6158,N_6591);
and U6889 (N_6889,N_6471,N_6423);
nor U6890 (N_6890,N_6177,N_6305);
nand U6891 (N_6891,N_6151,N_6227);
and U6892 (N_6892,N_6258,N_6098);
xnor U6893 (N_6893,N_6261,N_6332);
nand U6894 (N_6894,N_6315,N_6189);
and U6895 (N_6895,N_6033,N_6445);
nor U6896 (N_6896,N_6054,N_6271);
xnor U6897 (N_6897,N_6483,N_6439);
nand U6898 (N_6898,N_6285,N_6435);
xnor U6899 (N_6899,N_6281,N_6149);
nor U6900 (N_6900,N_6401,N_6127);
nor U6901 (N_6901,N_6509,N_6212);
xnor U6902 (N_6902,N_6413,N_6429);
or U6903 (N_6903,N_6202,N_6443);
or U6904 (N_6904,N_6333,N_6187);
nand U6905 (N_6905,N_6448,N_6578);
nand U6906 (N_6906,N_6462,N_6439);
or U6907 (N_6907,N_6189,N_6105);
nor U6908 (N_6908,N_6173,N_6453);
and U6909 (N_6909,N_6396,N_6121);
nor U6910 (N_6910,N_6378,N_6222);
or U6911 (N_6911,N_6021,N_6529);
or U6912 (N_6912,N_6187,N_6426);
or U6913 (N_6913,N_6323,N_6244);
nand U6914 (N_6914,N_6227,N_6394);
and U6915 (N_6915,N_6572,N_6313);
xor U6916 (N_6916,N_6367,N_6481);
or U6917 (N_6917,N_6461,N_6458);
or U6918 (N_6918,N_6391,N_6427);
nand U6919 (N_6919,N_6047,N_6414);
nor U6920 (N_6920,N_6447,N_6456);
or U6921 (N_6921,N_6198,N_6513);
and U6922 (N_6922,N_6363,N_6130);
nand U6923 (N_6923,N_6373,N_6156);
xnor U6924 (N_6924,N_6389,N_6295);
xnor U6925 (N_6925,N_6441,N_6069);
and U6926 (N_6926,N_6339,N_6233);
nor U6927 (N_6927,N_6155,N_6456);
or U6928 (N_6928,N_6048,N_6380);
or U6929 (N_6929,N_6588,N_6182);
xnor U6930 (N_6930,N_6581,N_6245);
nor U6931 (N_6931,N_6058,N_6313);
nor U6932 (N_6932,N_6474,N_6149);
xor U6933 (N_6933,N_6374,N_6290);
nand U6934 (N_6934,N_6072,N_6215);
nor U6935 (N_6935,N_6006,N_6093);
or U6936 (N_6936,N_6245,N_6282);
nand U6937 (N_6937,N_6079,N_6549);
xor U6938 (N_6938,N_6393,N_6155);
nor U6939 (N_6939,N_6112,N_6268);
and U6940 (N_6940,N_6134,N_6510);
xor U6941 (N_6941,N_6190,N_6178);
and U6942 (N_6942,N_6347,N_6256);
and U6943 (N_6943,N_6240,N_6588);
nor U6944 (N_6944,N_6492,N_6099);
nand U6945 (N_6945,N_6491,N_6583);
nand U6946 (N_6946,N_6540,N_6338);
nor U6947 (N_6947,N_6078,N_6255);
xor U6948 (N_6948,N_6044,N_6522);
nor U6949 (N_6949,N_6173,N_6121);
or U6950 (N_6950,N_6196,N_6297);
nor U6951 (N_6951,N_6062,N_6292);
nor U6952 (N_6952,N_6028,N_6490);
or U6953 (N_6953,N_6239,N_6448);
and U6954 (N_6954,N_6298,N_6161);
or U6955 (N_6955,N_6438,N_6363);
or U6956 (N_6956,N_6233,N_6271);
or U6957 (N_6957,N_6347,N_6072);
or U6958 (N_6958,N_6546,N_6218);
nor U6959 (N_6959,N_6209,N_6161);
or U6960 (N_6960,N_6044,N_6473);
nand U6961 (N_6961,N_6255,N_6591);
xnor U6962 (N_6962,N_6053,N_6229);
xor U6963 (N_6963,N_6517,N_6301);
or U6964 (N_6964,N_6289,N_6197);
nand U6965 (N_6965,N_6105,N_6426);
and U6966 (N_6966,N_6492,N_6169);
nor U6967 (N_6967,N_6576,N_6240);
nand U6968 (N_6968,N_6154,N_6342);
nor U6969 (N_6969,N_6239,N_6531);
nor U6970 (N_6970,N_6099,N_6383);
or U6971 (N_6971,N_6467,N_6474);
nand U6972 (N_6972,N_6457,N_6570);
or U6973 (N_6973,N_6332,N_6354);
and U6974 (N_6974,N_6325,N_6234);
xnor U6975 (N_6975,N_6020,N_6287);
or U6976 (N_6976,N_6357,N_6485);
or U6977 (N_6977,N_6112,N_6044);
and U6978 (N_6978,N_6447,N_6302);
xnor U6979 (N_6979,N_6315,N_6346);
nor U6980 (N_6980,N_6084,N_6216);
or U6981 (N_6981,N_6536,N_6581);
nand U6982 (N_6982,N_6348,N_6439);
and U6983 (N_6983,N_6217,N_6172);
xor U6984 (N_6984,N_6284,N_6306);
nor U6985 (N_6985,N_6143,N_6550);
or U6986 (N_6986,N_6407,N_6451);
and U6987 (N_6987,N_6206,N_6168);
nand U6988 (N_6988,N_6032,N_6317);
and U6989 (N_6989,N_6129,N_6477);
or U6990 (N_6990,N_6170,N_6430);
and U6991 (N_6991,N_6237,N_6087);
xnor U6992 (N_6992,N_6137,N_6383);
or U6993 (N_6993,N_6027,N_6213);
nor U6994 (N_6994,N_6577,N_6480);
or U6995 (N_6995,N_6478,N_6569);
and U6996 (N_6996,N_6031,N_6263);
nand U6997 (N_6997,N_6030,N_6295);
and U6998 (N_6998,N_6070,N_6023);
nor U6999 (N_6999,N_6451,N_6327);
and U7000 (N_7000,N_6588,N_6373);
or U7001 (N_7001,N_6137,N_6473);
or U7002 (N_7002,N_6288,N_6249);
xnor U7003 (N_7003,N_6390,N_6498);
nand U7004 (N_7004,N_6291,N_6400);
nand U7005 (N_7005,N_6118,N_6394);
xor U7006 (N_7006,N_6374,N_6182);
nand U7007 (N_7007,N_6078,N_6122);
or U7008 (N_7008,N_6130,N_6531);
and U7009 (N_7009,N_6136,N_6171);
nor U7010 (N_7010,N_6156,N_6299);
nor U7011 (N_7011,N_6470,N_6155);
nor U7012 (N_7012,N_6001,N_6506);
xor U7013 (N_7013,N_6512,N_6224);
and U7014 (N_7014,N_6582,N_6355);
xnor U7015 (N_7015,N_6426,N_6299);
or U7016 (N_7016,N_6492,N_6268);
nor U7017 (N_7017,N_6192,N_6372);
nor U7018 (N_7018,N_6515,N_6297);
or U7019 (N_7019,N_6037,N_6518);
nand U7020 (N_7020,N_6479,N_6180);
or U7021 (N_7021,N_6241,N_6196);
nor U7022 (N_7022,N_6506,N_6483);
or U7023 (N_7023,N_6479,N_6053);
nand U7024 (N_7024,N_6376,N_6101);
xnor U7025 (N_7025,N_6320,N_6010);
and U7026 (N_7026,N_6219,N_6001);
xnor U7027 (N_7027,N_6086,N_6176);
and U7028 (N_7028,N_6230,N_6552);
xnor U7029 (N_7029,N_6154,N_6129);
nand U7030 (N_7030,N_6497,N_6379);
and U7031 (N_7031,N_6202,N_6291);
xor U7032 (N_7032,N_6229,N_6558);
xnor U7033 (N_7033,N_6067,N_6278);
or U7034 (N_7034,N_6234,N_6475);
or U7035 (N_7035,N_6457,N_6150);
or U7036 (N_7036,N_6260,N_6097);
and U7037 (N_7037,N_6305,N_6269);
xnor U7038 (N_7038,N_6580,N_6040);
xnor U7039 (N_7039,N_6162,N_6285);
and U7040 (N_7040,N_6110,N_6055);
xor U7041 (N_7041,N_6083,N_6155);
nand U7042 (N_7042,N_6515,N_6442);
nand U7043 (N_7043,N_6358,N_6251);
nor U7044 (N_7044,N_6411,N_6153);
and U7045 (N_7045,N_6596,N_6171);
nand U7046 (N_7046,N_6025,N_6456);
nor U7047 (N_7047,N_6054,N_6246);
xor U7048 (N_7048,N_6454,N_6367);
and U7049 (N_7049,N_6281,N_6224);
nand U7050 (N_7050,N_6335,N_6217);
nor U7051 (N_7051,N_6135,N_6070);
or U7052 (N_7052,N_6278,N_6398);
and U7053 (N_7053,N_6540,N_6413);
nand U7054 (N_7054,N_6536,N_6584);
nor U7055 (N_7055,N_6313,N_6148);
nor U7056 (N_7056,N_6400,N_6381);
or U7057 (N_7057,N_6269,N_6135);
and U7058 (N_7058,N_6208,N_6046);
nor U7059 (N_7059,N_6113,N_6452);
nand U7060 (N_7060,N_6547,N_6421);
or U7061 (N_7061,N_6471,N_6434);
xnor U7062 (N_7062,N_6432,N_6570);
or U7063 (N_7063,N_6099,N_6014);
nor U7064 (N_7064,N_6594,N_6270);
xor U7065 (N_7065,N_6337,N_6466);
xor U7066 (N_7066,N_6142,N_6118);
nor U7067 (N_7067,N_6550,N_6004);
nand U7068 (N_7068,N_6439,N_6181);
nor U7069 (N_7069,N_6558,N_6108);
or U7070 (N_7070,N_6230,N_6133);
nand U7071 (N_7071,N_6347,N_6134);
nor U7072 (N_7072,N_6499,N_6240);
nor U7073 (N_7073,N_6262,N_6339);
nor U7074 (N_7074,N_6260,N_6298);
xor U7075 (N_7075,N_6306,N_6272);
xnor U7076 (N_7076,N_6390,N_6185);
nor U7077 (N_7077,N_6583,N_6390);
and U7078 (N_7078,N_6587,N_6348);
nor U7079 (N_7079,N_6521,N_6191);
or U7080 (N_7080,N_6001,N_6365);
xnor U7081 (N_7081,N_6129,N_6227);
nor U7082 (N_7082,N_6207,N_6557);
or U7083 (N_7083,N_6472,N_6325);
nand U7084 (N_7084,N_6471,N_6087);
xor U7085 (N_7085,N_6467,N_6432);
nor U7086 (N_7086,N_6101,N_6598);
and U7087 (N_7087,N_6038,N_6257);
xnor U7088 (N_7088,N_6074,N_6198);
and U7089 (N_7089,N_6065,N_6261);
nand U7090 (N_7090,N_6340,N_6049);
or U7091 (N_7091,N_6083,N_6538);
or U7092 (N_7092,N_6039,N_6136);
and U7093 (N_7093,N_6280,N_6043);
or U7094 (N_7094,N_6548,N_6083);
nand U7095 (N_7095,N_6497,N_6467);
xor U7096 (N_7096,N_6393,N_6206);
and U7097 (N_7097,N_6300,N_6216);
and U7098 (N_7098,N_6488,N_6400);
or U7099 (N_7099,N_6573,N_6207);
nand U7100 (N_7100,N_6561,N_6472);
and U7101 (N_7101,N_6011,N_6208);
nand U7102 (N_7102,N_6134,N_6569);
or U7103 (N_7103,N_6196,N_6400);
xnor U7104 (N_7104,N_6022,N_6515);
xnor U7105 (N_7105,N_6336,N_6122);
xor U7106 (N_7106,N_6592,N_6342);
nor U7107 (N_7107,N_6346,N_6214);
nor U7108 (N_7108,N_6582,N_6344);
nor U7109 (N_7109,N_6439,N_6415);
nand U7110 (N_7110,N_6597,N_6461);
and U7111 (N_7111,N_6307,N_6323);
nor U7112 (N_7112,N_6417,N_6234);
xor U7113 (N_7113,N_6526,N_6222);
nand U7114 (N_7114,N_6123,N_6447);
nand U7115 (N_7115,N_6351,N_6092);
xnor U7116 (N_7116,N_6483,N_6410);
and U7117 (N_7117,N_6013,N_6232);
nor U7118 (N_7118,N_6021,N_6519);
nor U7119 (N_7119,N_6399,N_6499);
and U7120 (N_7120,N_6389,N_6424);
nor U7121 (N_7121,N_6183,N_6359);
or U7122 (N_7122,N_6022,N_6206);
and U7123 (N_7123,N_6260,N_6523);
and U7124 (N_7124,N_6312,N_6471);
and U7125 (N_7125,N_6065,N_6384);
or U7126 (N_7126,N_6101,N_6441);
nand U7127 (N_7127,N_6051,N_6561);
and U7128 (N_7128,N_6115,N_6037);
and U7129 (N_7129,N_6380,N_6451);
and U7130 (N_7130,N_6232,N_6213);
or U7131 (N_7131,N_6094,N_6109);
or U7132 (N_7132,N_6099,N_6430);
nor U7133 (N_7133,N_6301,N_6319);
or U7134 (N_7134,N_6264,N_6341);
or U7135 (N_7135,N_6169,N_6194);
nand U7136 (N_7136,N_6317,N_6366);
nor U7137 (N_7137,N_6242,N_6552);
or U7138 (N_7138,N_6495,N_6238);
xor U7139 (N_7139,N_6003,N_6318);
xnor U7140 (N_7140,N_6525,N_6099);
nor U7141 (N_7141,N_6578,N_6560);
nor U7142 (N_7142,N_6406,N_6325);
or U7143 (N_7143,N_6442,N_6261);
and U7144 (N_7144,N_6407,N_6514);
nor U7145 (N_7145,N_6019,N_6317);
xor U7146 (N_7146,N_6503,N_6436);
nor U7147 (N_7147,N_6503,N_6012);
and U7148 (N_7148,N_6162,N_6508);
xnor U7149 (N_7149,N_6197,N_6082);
nor U7150 (N_7150,N_6154,N_6341);
and U7151 (N_7151,N_6215,N_6008);
nand U7152 (N_7152,N_6356,N_6200);
or U7153 (N_7153,N_6176,N_6266);
or U7154 (N_7154,N_6487,N_6546);
nor U7155 (N_7155,N_6376,N_6473);
and U7156 (N_7156,N_6252,N_6068);
or U7157 (N_7157,N_6077,N_6088);
or U7158 (N_7158,N_6476,N_6018);
or U7159 (N_7159,N_6590,N_6498);
xor U7160 (N_7160,N_6003,N_6335);
nor U7161 (N_7161,N_6496,N_6534);
nand U7162 (N_7162,N_6436,N_6045);
xor U7163 (N_7163,N_6266,N_6022);
nor U7164 (N_7164,N_6416,N_6153);
nand U7165 (N_7165,N_6290,N_6264);
and U7166 (N_7166,N_6559,N_6581);
or U7167 (N_7167,N_6198,N_6116);
nor U7168 (N_7168,N_6350,N_6406);
nor U7169 (N_7169,N_6454,N_6564);
and U7170 (N_7170,N_6083,N_6305);
and U7171 (N_7171,N_6434,N_6132);
xor U7172 (N_7172,N_6325,N_6097);
and U7173 (N_7173,N_6367,N_6188);
and U7174 (N_7174,N_6003,N_6035);
xnor U7175 (N_7175,N_6337,N_6015);
or U7176 (N_7176,N_6525,N_6551);
xor U7177 (N_7177,N_6496,N_6011);
nor U7178 (N_7178,N_6378,N_6546);
xor U7179 (N_7179,N_6145,N_6532);
nor U7180 (N_7180,N_6175,N_6313);
and U7181 (N_7181,N_6452,N_6235);
nand U7182 (N_7182,N_6169,N_6568);
or U7183 (N_7183,N_6476,N_6324);
and U7184 (N_7184,N_6568,N_6148);
or U7185 (N_7185,N_6410,N_6407);
xor U7186 (N_7186,N_6359,N_6424);
nand U7187 (N_7187,N_6387,N_6313);
xor U7188 (N_7188,N_6114,N_6346);
nor U7189 (N_7189,N_6564,N_6072);
and U7190 (N_7190,N_6157,N_6099);
xnor U7191 (N_7191,N_6031,N_6236);
and U7192 (N_7192,N_6542,N_6263);
or U7193 (N_7193,N_6076,N_6509);
nand U7194 (N_7194,N_6079,N_6045);
and U7195 (N_7195,N_6412,N_6368);
or U7196 (N_7196,N_6072,N_6235);
and U7197 (N_7197,N_6498,N_6289);
or U7198 (N_7198,N_6329,N_6187);
and U7199 (N_7199,N_6076,N_6045);
xnor U7200 (N_7200,N_6768,N_6991);
xnor U7201 (N_7201,N_6814,N_6981);
or U7202 (N_7202,N_6792,N_6916);
nor U7203 (N_7203,N_7020,N_7155);
nand U7204 (N_7204,N_6834,N_6955);
and U7205 (N_7205,N_6801,N_7162);
xor U7206 (N_7206,N_7026,N_6890);
xor U7207 (N_7207,N_6965,N_6812);
xnor U7208 (N_7208,N_6788,N_6951);
or U7209 (N_7209,N_6789,N_6726);
and U7210 (N_7210,N_6840,N_7051);
xnor U7211 (N_7211,N_7046,N_6849);
nand U7212 (N_7212,N_6641,N_6624);
xor U7213 (N_7213,N_7062,N_6912);
xnor U7214 (N_7214,N_6645,N_6870);
and U7215 (N_7215,N_6715,N_6829);
xor U7216 (N_7216,N_6717,N_6983);
and U7217 (N_7217,N_7097,N_7085);
or U7218 (N_7218,N_7102,N_6659);
and U7219 (N_7219,N_7004,N_7030);
and U7220 (N_7220,N_6640,N_7093);
xor U7221 (N_7221,N_6978,N_6701);
and U7222 (N_7222,N_7158,N_6727);
and U7223 (N_7223,N_6618,N_7188);
nand U7224 (N_7224,N_6879,N_6620);
xnor U7225 (N_7225,N_6841,N_6807);
nor U7226 (N_7226,N_6649,N_6854);
nand U7227 (N_7227,N_6658,N_7041);
nor U7228 (N_7228,N_7134,N_7048);
nor U7229 (N_7229,N_6853,N_6730);
nand U7230 (N_7230,N_6937,N_6868);
nor U7231 (N_7231,N_6838,N_7074);
or U7232 (N_7232,N_6857,N_6652);
or U7233 (N_7233,N_7038,N_6986);
nor U7234 (N_7234,N_7112,N_7068);
nand U7235 (N_7235,N_7096,N_6646);
nor U7236 (N_7236,N_6610,N_7057);
or U7237 (N_7237,N_6785,N_7084);
nand U7238 (N_7238,N_6704,N_6975);
and U7239 (N_7239,N_7125,N_6990);
nor U7240 (N_7240,N_6636,N_6821);
xnor U7241 (N_7241,N_6989,N_6667);
nand U7242 (N_7242,N_7178,N_6781);
nor U7243 (N_7243,N_7056,N_6804);
xor U7244 (N_7244,N_6777,N_6631);
or U7245 (N_7245,N_7145,N_7010);
and U7246 (N_7246,N_6694,N_7121);
nand U7247 (N_7247,N_6628,N_6762);
nand U7248 (N_7248,N_6939,N_6712);
nand U7249 (N_7249,N_7189,N_6839);
and U7250 (N_7250,N_7065,N_6865);
or U7251 (N_7251,N_7027,N_6705);
nand U7252 (N_7252,N_7042,N_6711);
xnor U7253 (N_7253,N_6710,N_6832);
nor U7254 (N_7254,N_7153,N_6621);
nor U7255 (N_7255,N_6703,N_7183);
nor U7256 (N_7256,N_6896,N_7031);
nand U7257 (N_7257,N_7163,N_6984);
xnor U7258 (N_7258,N_7135,N_6752);
or U7259 (N_7259,N_7156,N_6793);
and U7260 (N_7260,N_6976,N_7137);
nor U7261 (N_7261,N_6889,N_6842);
xor U7262 (N_7262,N_6791,N_6906);
nand U7263 (N_7263,N_6784,N_6681);
nand U7264 (N_7264,N_6707,N_6608);
nand U7265 (N_7265,N_6815,N_6958);
and U7266 (N_7266,N_6682,N_6880);
or U7267 (N_7267,N_6696,N_6940);
nand U7268 (N_7268,N_6823,N_6771);
and U7269 (N_7269,N_6739,N_6790);
or U7270 (N_7270,N_6905,N_6898);
nor U7271 (N_7271,N_7117,N_6936);
nand U7272 (N_7272,N_6846,N_6946);
nor U7273 (N_7273,N_7069,N_7127);
and U7274 (N_7274,N_7089,N_6613);
xnor U7275 (N_7275,N_7076,N_6921);
and U7276 (N_7276,N_6918,N_6885);
nand U7277 (N_7277,N_6883,N_6616);
and U7278 (N_7278,N_6670,N_6735);
or U7279 (N_7279,N_7071,N_7081);
or U7280 (N_7280,N_6714,N_6644);
or U7281 (N_7281,N_7035,N_7072);
xor U7282 (N_7282,N_7091,N_6909);
nor U7283 (N_7283,N_6766,N_7122);
nand U7284 (N_7284,N_7021,N_7019);
xnor U7285 (N_7285,N_6723,N_7025);
or U7286 (N_7286,N_6973,N_6678);
xor U7287 (N_7287,N_6760,N_7087);
or U7288 (N_7288,N_6943,N_7083);
and U7289 (N_7289,N_6622,N_7172);
xor U7290 (N_7290,N_7040,N_7133);
nor U7291 (N_7291,N_7186,N_6996);
nand U7292 (N_7292,N_7118,N_6875);
nand U7293 (N_7293,N_6850,N_6968);
and U7294 (N_7294,N_6695,N_7138);
nor U7295 (N_7295,N_6873,N_7104);
nand U7296 (N_7296,N_7070,N_7168);
xnor U7297 (N_7297,N_6864,N_7124);
nor U7298 (N_7298,N_7011,N_6774);
or U7299 (N_7299,N_6716,N_6617);
or U7300 (N_7300,N_6897,N_7106);
and U7301 (N_7301,N_6605,N_7060);
nand U7302 (N_7302,N_6919,N_6692);
and U7303 (N_7303,N_6686,N_6928);
and U7304 (N_7304,N_6929,N_7181);
or U7305 (N_7305,N_6706,N_6950);
and U7306 (N_7306,N_6655,N_6687);
or U7307 (N_7307,N_6754,N_6871);
nand U7308 (N_7308,N_6887,N_6900);
nand U7309 (N_7309,N_6600,N_6825);
nand U7310 (N_7310,N_7128,N_7002);
nand U7311 (N_7311,N_7029,N_6925);
nor U7312 (N_7312,N_7080,N_6718);
xor U7313 (N_7313,N_6819,N_7184);
or U7314 (N_7314,N_6786,N_7018);
nand U7315 (N_7315,N_6901,N_6720);
and U7316 (N_7316,N_7054,N_6988);
xor U7317 (N_7317,N_6748,N_6851);
nor U7318 (N_7318,N_7176,N_6810);
xnor U7319 (N_7319,N_6660,N_6765);
or U7320 (N_7320,N_6953,N_7034);
and U7321 (N_7321,N_7157,N_6957);
nand U7322 (N_7322,N_6809,N_6904);
and U7323 (N_7323,N_6627,N_7006);
and U7324 (N_7324,N_6891,N_6917);
and U7325 (N_7325,N_7101,N_6893);
and U7326 (N_7326,N_6878,N_7141);
nor U7327 (N_7327,N_6997,N_7009);
nor U7328 (N_7328,N_6626,N_7197);
nor U7329 (N_7329,N_6759,N_6673);
and U7330 (N_7330,N_6648,N_7115);
xor U7331 (N_7331,N_6866,N_7024);
and U7332 (N_7332,N_6833,N_6637);
nand U7333 (N_7333,N_7014,N_6818);
nor U7334 (N_7334,N_6732,N_6799);
nor U7335 (N_7335,N_6972,N_6805);
xnor U7336 (N_7336,N_7045,N_7103);
or U7337 (N_7337,N_7159,N_6861);
nand U7338 (N_7338,N_6734,N_6954);
xnor U7339 (N_7339,N_6782,N_6974);
or U7340 (N_7340,N_7196,N_6941);
nor U7341 (N_7341,N_6822,N_6606);
nor U7342 (N_7342,N_7150,N_6926);
nor U7343 (N_7343,N_7092,N_7039);
nand U7344 (N_7344,N_7180,N_6743);
and U7345 (N_7345,N_6657,N_7140);
xor U7346 (N_7346,N_6930,N_6740);
or U7347 (N_7347,N_6862,N_6664);
nor U7348 (N_7348,N_6653,N_6876);
nand U7349 (N_7349,N_6836,N_7095);
nand U7350 (N_7350,N_6947,N_6647);
and U7351 (N_7351,N_6945,N_6858);
or U7352 (N_7352,N_7160,N_6757);
and U7353 (N_7353,N_6787,N_6676);
nand U7354 (N_7354,N_6744,N_7049);
and U7355 (N_7355,N_6629,N_6601);
or U7356 (N_7356,N_6859,N_6722);
nor U7357 (N_7357,N_7146,N_7000);
and U7358 (N_7358,N_6775,N_7037);
or U7359 (N_7359,N_6602,N_7116);
or U7360 (N_7360,N_6699,N_6827);
xor U7361 (N_7361,N_6662,N_6728);
nand U7362 (N_7362,N_7098,N_6632);
xor U7363 (N_7363,N_6902,N_6778);
xnor U7364 (N_7364,N_6999,N_7131);
xnor U7365 (N_7365,N_6994,N_7055);
or U7366 (N_7366,N_6964,N_6679);
and U7367 (N_7367,N_6808,N_7050);
or U7368 (N_7368,N_7142,N_6835);
nand U7369 (N_7369,N_6713,N_7110);
and U7370 (N_7370,N_6960,N_6654);
xor U7371 (N_7371,N_6907,N_6803);
xnor U7372 (N_7372,N_6860,N_7123);
or U7373 (N_7373,N_7136,N_7171);
and U7374 (N_7374,N_7017,N_6745);
or U7375 (N_7375,N_6719,N_6697);
nand U7376 (N_7376,N_6747,N_6761);
and U7377 (N_7377,N_7194,N_6817);
or U7378 (N_7378,N_6733,N_7170);
or U7379 (N_7379,N_7052,N_7044);
nor U7380 (N_7380,N_7167,N_7152);
and U7381 (N_7381,N_6795,N_7120);
nand U7382 (N_7382,N_7198,N_6603);
and U7383 (N_7383,N_6746,N_6800);
nand U7384 (N_7384,N_6985,N_7099);
and U7385 (N_7385,N_6663,N_6680);
or U7386 (N_7386,N_6852,N_6806);
nand U7387 (N_7387,N_6993,N_6635);
and U7388 (N_7388,N_6668,N_6843);
or U7389 (N_7389,N_7023,N_6867);
and U7390 (N_7390,N_6779,N_6982);
xnor U7391 (N_7391,N_6837,N_6855);
nor U7392 (N_7392,N_6820,N_7195);
nor U7393 (N_7393,N_6656,N_6758);
xnor U7394 (N_7394,N_6738,N_6625);
nor U7395 (N_7395,N_6903,N_6816);
xnor U7396 (N_7396,N_6750,N_7173);
xor U7397 (N_7397,N_6773,N_6729);
nand U7398 (N_7398,N_7139,N_6931);
nor U7399 (N_7399,N_7013,N_6736);
nor U7400 (N_7400,N_6970,N_6721);
xnor U7401 (N_7401,N_6708,N_7066);
nor U7402 (N_7402,N_6642,N_7126);
xnor U7403 (N_7403,N_7130,N_6848);
and U7404 (N_7404,N_6948,N_7105);
xnor U7405 (N_7405,N_6922,N_6796);
nand U7406 (N_7406,N_6998,N_6770);
or U7407 (N_7407,N_7005,N_6908);
xor U7408 (N_7408,N_7036,N_6798);
or U7409 (N_7409,N_6856,N_6671);
nor U7410 (N_7410,N_6888,N_7192);
xnor U7411 (N_7411,N_6693,N_6623);
xor U7412 (N_7412,N_6741,N_6828);
nor U7413 (N_7413,N_6685,N_6844);
and U7414 (N_7414,N_7182,N_6971);
and U7415 (N_7415,N_6604,N_7090);
xor U7416 (N_7416,N_6892,N_7107);
xnor U7417 (N_7417,N_7193,N_6731);
or U7418 (N_7418,N_6612,N_7111);
xnor U7419 (N_7419,N_6675,N_6932);
or U7420 (N_7420,N_7094,N_6992);
or U7421 (N_7421,N_7077,N_6987);
or U7422 (N_7422,N_7082,N_7064);
or U7423 (N_7423,N_7012,N_6755);
xnor U7424 (N_7424,N_6672,N_6977);
and U7425 (N_7425,N_6884,N_7185);
and U7426 (N_7426,N_6944,N_6933);
nand U7427 (N_7427,N_6935,N_7149);
and U7428 (N_7428,N_7148,N_6927);
or U7429 (N_7429,N_6920,N_6633);
or U7430 (N_7430,N_6961,N_6874);
nand U7431 (N_7431,N_6639,N_6689);
nor U7432 (N_7432,N_6702,N_6756);
nand U7433 (N_7433,N_6698,N_6630);
and U7434 (N_7434,N_6959,N_6763);
xnor U7435 (N_7435,N_7022,N_7151);
or U7436 (N_7436,N_7129,N_7086);
or U7437 (N_7437,N_6826,N_6938);
xnor U7438 (N_7438,N_7119,N_7001);
or U7439 (N_7439,N_7187,N_7166);
nor U7440 (N_7440,N_6742,N_6845);
and U7441 (N_7441,N_7109,N_7063);
nor U7442 (N_7442,N_6709,N_6877);
nand U7443 (N_7443,N_6615,N_7191);
nand U7444 (N_7444,N_7075,N_6751);
or U7445 (N_7445,N_7008,N_6683);
nand U7446 (N_7446,N_6651,N_7073);
nor U7447 (N_7447,N_6952,N_6776);
nor U7448 (N_7448,N_6737,N_6811);
xor U7449 (N_7449,N_6609,N_6638);
or U7450 (N_7450,N_6963,N_7190);
nor U7451 (N_7451,N_6611,N_6881);
xnor U7452 (N_7452,N_6666,N_6783);
and U7453 (N_7453,N_6688,N_7015);
nor U7454 (N_7454,N_7033,N_6914);
nand U7455 (N_7455,N_6753,N_6749);
nand U7456 (N_7456,N_6772,N_6665);
nor U7457 (N_7457,N_7047,N_7061);
nor U7458 (N_7458,N_7164,N_6980);
xor U7459 (N_7459,N_6831,N_6942);
nor U7460 (N_7460,N_6797,N_7199);
or U7461 (N_7461,N_6910,N_7043);
nor U7462 (N_7462,N_7059,N_6924);
and U7463 (N_7463,N_7174,N_6824);
or U7464 (N_7464,N_7016,N_6830);
nor U7465 (N_7465,N_7100,N_6895);
xor U7466 (N_7466,N_6725,N_6995);
xnor U7467 (N_7467,N_7161,N_6724);
nand U7468 (N_7468,N_6691,N_6962);
xnor U7469 (N_7469,N_7007,N_6872);
xor U7470 (N_7470,N_7078,N_6802);
nand U7471 (N_7471,N_6847,N_6634);
or U7472 (N_7472,N_7169,N_7154);
nand U7473 (N_7473,N_7132,N_6767);
and U7474 (N_7474,N_7165,N_6869);
nand U7475 (N_7475,N_6794,N_7088);
nand U7476 (N_7476,N_6684,N_6934);
and U7477 (N_7477,N_6967,N_6886);
xnor U7478 (N_7478,N_7053,N_7114);
or U7479 (N_7479,N_6607,N_7113);
or U7480 (N_7480,N_6911,N_7144);
nor U7481 (N_7481,N_6863,N_6614);
nor U7482 (N_7482,N_6949,N_6966);
xnor U7483 (N_7483,N_6661,N_6915);
nor U7484 (N_7484,N_6894,N_6769);
and U7485 (N_7485,N_6956,N_7147);
nor U7486 (N_7486,N_6923,N_6690);
and U7487 (N_7487,N_7143,N_7079);
xor U7488 (N_7488,N_6899,N_7058);
and U7489 (N_7489,N_7108,N_6619);
or U7490 (N_7490,N_6643,N_7032);
nor U7491 (N_7491,N_6969,N_7177);
or U7492 (N_7492,N_6700,N_7175);
and U7493 (N_7493,N_7179,N_6650);
nor U7494 (N_7494,N_7028,N_6674);
and U7495 (N_7495,N_7067,N_6764);
nor U7496 (N_7496,N_6913,N_6780);
nor U7497 (N_7497,N_6813,N_6669);
xor U7498 (N_7498,N_6677,N_6882);
nor U7499 (N_7499,N_6979,N_7003);
or U7500 (N_7500,N_6729,N_6885);
and U7501 (N_7501,N_6767,N_6647);
nor U7502 (N_7502,N_6628,N_6851);
nor U7503 (N_7503,N_6999,N_6706);
and U7504 (N_7504,N_7192,N_6635);
nor U7505 (N_7505,N_6880,N_6965);
and U7506 (N_7506,N_6983,N_6971);
and U7507 (N_7507,N_6833,N_6643);
nor U7508 (N_7508,N_6873,N_6729);
nand U7509 (N_7509,N_7076,N_6998);
nor U7510 (N_7510,N_6792,N_6646);
nor U7511 (N_7511,N_6848,N_6947);
xor U7512 (N_7512,N_6775,N_6636);
and U7513 (N_7513,N_6931,N_6690);
nand U7514 (N_7514,N_6960,N_6606);
nor U7515 (N_7515,N_7186,N_7136);
nand U7516 (N_7516,N_7016,N_6747);
or U7517 (N_7517,N_6815,N_7193);
or U7518 (N_7518,N_6605,N_7158);
or U7519 (N_7519,N_7120,N_6785);
xor U7520 (N_7520,N_7158,N_6877);
nor U7521 (N_7521,N_6649,N_7151);
xor U7522 (N_7522,N_7166,N_7174);
xor U7523 (N_7523,N_7003,N_6955);
and U7524 (N_7524,N_7062,N_7170);
and U7525 (N_7525,N_6655,N_6863);
nor U7526 (N_7526,N_7120,N_6881);
nor U7527 (N_7527,N_6825,N_7077);
or U7528 (N_7528,N_6666,N_7165);
nand U7529 (N_7529,N_6742,N_7186);
or U7530 (N_7530,N_6703,N_7158);
and U7531 (N_7531,N_7093,N_6763);
and U7532 (N_7532,N_6951,N_6975);
or U7533 (N_7533,N_6665,N_6825);
nand U7534 (N_7534,N_6606,N_7198);
nand U7535 (N_7535,N_7124,N_6970);
and U7536 (N_7536,N_7167,N_6649);
nand U7537 (N_7537,N_6838,N_6682);
and U7538 (N_7538,N_6936,N_6897);
xnor U7539 (N_7539,N_7193,N_7015);
nand U7540 (N_7540,N_6712,N_7005);
xor U7541 (N_7541,N_7012,N_6981);
nand U7542 (N_7542,N_6654,N_6962);
or U7543 (N_7543,N_7002,N_6708);
and U7544 (N_7544,N_6720,N_7131);
nand U7545 (N_7545,N_7111,N_6887);
and U7546 (N_7546,N_6860,N_6987);
nand U7547 (N_7547,N_6632,N_7053);
nor U7548 (N_7548,N_6663,N_6900);
xor U7549 (N_7549,N_6990,N_6629);
or U7550 (N_7550,N_6806,N_6761);
or U7551 (N_7551,N_7146,N_7194);
nand U7552 (N_7552,N_6655,N_6815);
or U7553 (N_7553,N_6606,N_7146);
nor U7554 (N_7554,N_6723,N_7118);
xnor U7555 (N_7555,N_7058,N_6781);
nor U7556 (N_7556,N_7140,N_6817);
nor U7557 (N_7557,N_6743,N_6602);
or U7558 (N_7558,N_7135,N_6716);
xor U7559 (N_7559,N_7137,N_6658);
or U7560 (N_7560,N_6671,N_7112);
nor U7561 (N_7561,N_7008,N_6630);
nand U7562 (N_7562,N_6773,N_7030);
xor U7563 (N_7563,N_6927,N_6718);
nand U7564 (N_7564,N_6868,N_7153);
xnor U7565 (N_7565,N_7156,N_6938);
nor U7566 (N_7566,N_6801,N_7192);
nand U7567 (N_7567,N_6752,N_6893);
or U7568 (N_7568,N_6750,N_6962);
and U7569 (N_7569,N_6976,N_6746);
nand U7570 (N_7570,N_6609,N_6765);
and U7571 (N_7571,N_7135,N_7091);
xor U7572 (N_7572,N_6981,N_7193);
nand U7573 (N_7573,N_6615,N_6658);
or U7574 (N_7574,N_6655,N_6758);
nor U7575 (N_7575,N_7195,N_6919);
nor U7576 (N_7576,N_7108,N_6784);
nand U7577 (N_7577,N_6658,N_6742);
xor U7578 (N_7578,N_6759,N_7037);
and U7579 (N_7579,N_7048,N_6806);
xor U7580 (N_7580,N_7104,N_7102);
or U7581 (N_7581,N_6638,N_6838);
and U7582 (N_7582,N_6870,N_7197);
or U7583 (N_7583,N_6900,N_6755);
nand U7584 (N_7584,N_6609,N_6844);
nor U7585 (N_7585,N_7025,N_7031);
and U7586 (N_7586,N_6619,N_6939);
xnor U7587 (N_7587,N_6982,N_6754);
xnor U7588 (N_7588,N_7005,N_7059);
nand U7589 (N_7589,N_6973,N_6958);
and U7590 (N_7590,N_6646,N_6748);
nand U7591 (N_7591,N_7077,N_6880);
xor U7592 (N_7592,N_6762,N_6706);
or U7593 (N_7593,N_7177,N_7188);
xor U7594 (N_7594,N_6672,N_6984);
and U7595 (N_7595,N_6911,N_7135);
xnor U7596 (N_7596,N_7075,N_6703);
xnor U7597 (N_7597,N_7128,N_6837);
and U7598 (N_7598,N_6657,N_6998);
xnor U7599 (N_7599,N_6703,N_6958);
or U7600 (N_7600,N_6778,N_6996);
nand U7601 (N_7601,N_6736,N_6656);
nand U7602 (N_7602,N_7175,N_6749);
and U7603 (N_7603,N_6827,N_6987);
nor U7604 (N_7604,N_6716,N_7024);
nor U7605 (N_7605,N_7041,N_7186);
or U7606 (N_7606,N_7192,N_6982);
and U7607 (N_7607,N_7164,N_6634);
nor U7608 (N_7608,N_7120,N_7102);
xor U7609 (N_7609,N_7056,N_7071);
nor U7610 (N_7610,N_7195,N_7061);
and U7611 (N_7611,N_6611,N_6705);
nor U7612 (N_7612,N_6914,N_6911);
and U7613 (N_7613,N_6619,N_7189);
or U7614 (N_7614,N_6652,N_7133);
xor U7615 (N_7615,N_7102,N_6943);
xor U7616 (N_7616,N_6804,N_6662);
nand U7617 (N_7617,N_7182,N_6792);
and U7618 (N_7618,N_6713,N_6729);
and U7619 (N_7619,N_6696,N_6828);
xor U7620 (N_7620,N_6984,N_6756);
xor U7621 (N_7621,N_6683,N_6950);
nor U7622 (N_7622,N_7081,N_6654);
or U7623 (N_7623,N_7004,N_6702);
or U7624 (N_7624,N_6997,N_6775);
or U7625 (N_7625,N_6885,N_7181);
nor U7626 (N_7626,N_6708,N_7178);
xor U7627 (N_7627,N_7078,N_7143);
and U7628 (N_7628,N_7179,N_6719);
and U7629 (N_7629,N_7072,N_6925);
nor U7630 (N_7630,N_7152,N_7140);
nor U7631 (N_7631,N_7195,N_6696);
and U7632 (N_7632,N_6681,N_7018);
xor U7633 (N_7633,N_6950,N_6867);
nor U7634 (N_7634,N_6628,N_6759);
nor U7635 (N_7635,N_6770,N_6971);
and U7636 (N_7636,N_7165,N_7055);
or U7637 (N_7637,N_7026,N_6937);
xnor U7638 (N_7638,N_6940,N_7055);
nand U7639 (N_7639,N_6683,N_6625);
nand U7640 (N_7640,N_6999,N_7143);
and U7641 (N_7641,N_7050,N_7042);
nor U7642 (N_7642,N_7140,N_7128);
or U7643 (N_7643,N_6870,N_6702);
xnor U7644 (N_7644,N_7125,N_6887);
xnor U7645 (N_7645,N_7091,N_6898);
nor U7646 (N_7646,N_6747,N_6898);
nor U7647 (N_7647,N_7175,N_6937);
or U7648 (N_7648,N_6813,N_7145);
and U7649 (N_7649,N_6915,N_6689);
xnor U7650 (N_7650,N_6782,N_7055);
or U7651 (N_7651,N_7149,N_7078);
nor U7652 (N_7652,N_7053,N_7065);
xnor U7653 (N_7653,N_7084,N_7135);
xor U7654 (N_7654,N_7024,N_6657);
and U7655 (N_7655,N_6866,N_7079);
and U7656 (N_7656,N_6908,N_7113);
xor U7657 (N_7657,N_7004,N_6967);
or U7658 (N_7658,N_6886,N_6639);
or U7659 (N_7659,N_6624,N_7124);
nor U7660 (N_7660,N_6741,N_6647);
nor U7661 (N_7661,N_7026,N_7033);
nor U7662 (N_7662,N_7175,N_6629);
nand U7663 (N_7663,N_7123,N_6784);
nand U7664 (N_7664,N_6695,N_6604);
xor U7665 (N_7665,N_7084,N_6955);
nor U7666 (N_7666,N_6704,N_6850);
or U7667 (N_7667,N_6800,N_6727);
xor U7668 (N_7668,N_7108,N_6767);
and U7669 (N_7669,N_7073,N_7003);
and U7670 (N_7670,N_7150,N_6845);
nor U7671 (N_7671,N_7124,N_6716);
nor U7672 (N_7672,N_7075,N_7185);
and U7673 (N_7673,N_6746,N_7117);
nand U7674 (N_7674,N_6726,N_6834);
nor U7675 (N_7675,N_7129,N_7153);
nand U7676 (N_7676,N_6829,N_6762);
nor U7677 (N_7677,N_6807,N_6720);
nand U7678 (N_7678,N_6847,N_6779);
and U7679 (N_7679,N_7040,N_6642);
or U7680 (N_7680,N_6872,N_7106);
nand U7681 (N_7681,N_7158,N_6989);
or U7682 (N_7682,N_6676,N_6947);
xor U7683 (N_7683,N_6766,N_7091);
or U7684 (N_7684,N_7171,N_6633);
nand U7685 (N_7685,N_6818,N_6894);
xor U7686 (N_7686,N_6876,N_6746);
nor U7687 (N_7687,N_6698,N_7082);
xnor U7688 (N_7688,N_6965,N_6777);
and U7689 (N_7689,N_6955,N_6728);
nand U7690 (N_7690,N_6753,N_6754);
and U7691 (N_7691,N_6653,N_7059);
nand U7692 (N_7692,N_7127,N_6947);
xor U7693 (N_7693,N_7048,N_6782);
and U7694 (N_7694,N_6942,N_6784);
or U7695 (N_7695,N_6868,N_6744);
nand U7696 (N_7696,N_7182,N_6824);
nor U7697 (N_7697,N_6649,N_6762);
nor U7698 (N_7698,N_6914,N_7029);
xor U7699 (N_7699,N_6666,N_6910);
nor U7700 (N_7700,N_7137,N_6702);
xnor U7701 (N_7701,N_6660,N_6701);
nor U7702 (N_7702,N_7186,N_7183);
and U7703 (N_7703,N_6784,N_7181);
or U7704 (N_7704,N_6770,N_6964);
nor U7705 (N_7705,N_6965,N_6867);
and U7706 (N_7706,N_6955,N_6703);
nand U7707 (N_7707,N_6791,N_7197);
or U7708 (N_7708,N_7023,N_7015);
nor U7709 (N_7709,N_7072,N_7041);
and U7710 (N_7710,N_6756,N_7180);
or U7711 (N_7711,N_6915,N_6638);
or U7712 (N_7712,N_7019,N_7144);
xnor U7713 (N_7713,N_6891,N_7033);
nand U7714 (N_7714,N_6863,N_6838);
nand U7715 (N_7715,N_6611,N_7006);
nor U7716 (N_7716,N_6851,N_7053);
and U7717 (N_7717,N_6657,N_7186);
and U7718 (N_7718,N_6820,N_6723);
xor U7719 (N_7719,N_6686,N_6993);
nor U7720 (N_7720,N_7076,N_7039);
xor U7721 (N_7721,N_6647,N_6894);
nand U7722 (N_7722,N_6609,N_6651);
nor U7723 (N_7723,N_6792,N_6955);
xnor U7724 (N_7724,N_7106,N_6935);
and U7725 (N_7725,N_6808,N_6616);
nand U7726 (N_7726,N_7128,N_6921);
nand U7727 (N_7727,N_6870,N_6601);
and U7728 (N_7728,N_6662,N_6870);
nor U7729 (N_7729,N_6785,N_6689);
or U7730 (N_7730,N_7041,N_6862);
and U7731 (N_7731,N_7101,N_6870);
and U7732 (N_7732,N_7152,N_6959);
nor U7733 (N_7733,N_6835,N_6842);
nand U7734 (N_7734,N_6620,N_7160);
and U7735 (N_7735,N_7008,N_6928);
nor U7736 (N_7736,N_6884,N_6809);
nor U7737 (N_7737,N_7176,N_6728);
xnor U7738 (N_7738,N_7092,N_6974);
nor U7739 (N_7739,N_6752,N_6835);
and U7740 (N_7740,N_6639,N_7099);
and U7741 (N_7741,N_6834,N_7043);
and U7742 (N_7742,N_6905,N_6619);
and U7743 (N_7743,N_6791,N_6650);
or U7744 (N_7744,N_7010,N_7175);
nand U7745 (N_7745,N_7011,N_6716);
xnor U7746 (N_7746,N_7104,N_6999);
nor U7747 (N_7747,N_6639,N_6825);
nor U7748 (N_7748,N_6865,N_6891);
nor U7749 (N_7749,N_6814,N_6699);
and U7750 (N_7750,N_6758,N_7138);
xor U7751 (N_7751,N_6625,N_6726);
nand U7752 (N_7752,N_6742,N_6857);
and U7753 (N_7753,N_7018,N_6818);
nand U7754 (N_7754,N_7041,N_6641);
nor U7755 (N_7755,N_6804,N_6960);
nand U7756 (N_7756,N_6856,N_6714);
nand U7757 (N_7757,N_7094,N_7131);
and U7758 (N_7758,N_6760,N_6844);
nor U7759 (N_7759,N_6935,N_7019);
and U7760 (N_7760,N_7095,N_6752);
xor U7761 (N_7761,N_6960,N_6931);
nand U7762 (N_7762,N_6918,N_6603);
or U7763 (N_7763,N_6639,N_7067);
and U7764 (N_7764,N_6933,N_7160);
nor U7765 (N_7765,N_7071,N_6630);
nor U7766 (N_7766,N_6902,N_6705);
nor U7767 (N_7767,N_6863,N_7117);
and U7768 (N_7768,N_6642,N_6993);
xor U7769 (N_7769,N_6654,N_7138);
nand U7770 (N_7770,N_7072,N_6996);
or U7771 (N_7771,N_6883,N_6901);
xor U7772 (N_7772,N_6617,N_6879);
or U7773 (N_7773,N_7125,N_6648);
xor U7774 (N_7774,N_6846,N_6944);
xor U7775 (N_7775,N_7110,N_6693);
xnor U7776 (N_7776,N_6706,N_6834);
nand U7777 (N_7777,N_7094,N_6637);
xnor U7778 (N_7778,N_6674,N_6842);
or U7779 (N_7779,N_6662,N_6680);
xnor U7780 (N_7780,N_7053,N_6615);
xnor U7781 (N_7781,N_7122,N_6850);
nor U7782 (N_7782,N_6723,N_7144);
xor U7783 (N_7783,N_7185,N_6968);
nand U7784 (N_7784,N_6615,N_7136);
nand U7785 (N_7785,N_6802,N_6729);
and U7786 (N_7786,N_6754,N_6797);
nor U7787 (N_7787,N_7078,N_6811);
nand U7788 (N_7788,N_7015,N_7094);
or U7789 (N_7789,N_6680,N_6618);
and U7790 (N_7790,N_6714,N_6793);
nor U7791 (N_7791,N_6774,N_6876);
nand U7792 (N_7792,N_7198,N_7103);
and U7793 (N_7793,N_6741,N_6654);
nand U7794 (N_7794,N_6805,N_6863);
xor U7795 (N_7795,N_6665,N_6888);
nor U7796 (N_7796,N_6863,N_6884);
or U7797 (N_7797,N_7107,N_6983);
xor U7798 (N_7798,N_6883,N_7194);
nand U7799 (N_7799,N_6700,N_6834);
xnor U7800 (N_7800,N_7425,N_7764);
xnor U7801 (N_7801,N_7725,N_7218);
xor U7802 (N_7802,N_7549,N_7414);
nor U7803 (N_7803,N_7701,N_7594);
or U7804 (N_7804,N_7598,N_7780);
nand U7805 (N_7805,N_7299,N_7774);
or U7806 (N_7806,N_7451,N_7672);
nand U7807 (N_7807,N_7342,N_7271);
nand U7808 (N_7808,N_7267,N_7762);
or U7809 (N_7809,N_7423,N_7263);
or U7810 (N_7810,N_7250,N_7562);
xor U7811 (N_7811,N_7752,N_7782);
xnor U7812 (N_7812,N_7678,N_7772);
nor U7813 (N_7813,N_7795,N_7429);
and U7814 (N_7814,N_7748,N_7335);
nor U7815 (N_7815,N_7475,N_7473);
or U7816 (N_7816,N_7515,N_7502);
or U7817 (N_7817,N_7791,N_7213);
xnor U7818 (N_7818,N_7489,N_7239);
nand U7819 (N_7819,N_7685,N_7212);
and U7820 (N_7820,N_7571,N_7629);
and U7821 (N_7821,N_7529,N_7301);
nor U7822 (N_7822,N_7447,N_7362);
xnor U7823 (N_7823,N_7757,N_7613);
nand U7824 (N_7824,N_7655,N_7368);
nor U7825 (N_7825,N_7719,N_7611);
or U7826 (N_7826,N_7215,N_7624);
nand U7827 (N_7827,N_7330,N_7394);
nand U7828 (N_7828,N_7426,N_7274);
nor U7829 (N_7829,N_7480,N_7221);
nand U7830 (N_7830,N_7641,N_7694);
xor U7831 (N_7831,N_7588,N_7495);
and U7832 (N_7832,N_7496,N_7441);
xnor U7833 (N_7833,N_7726,N_7770);
or U7834 (N_7834,N_7525,N_7751);
xnor U7835 (N_7835,N_7716,N_7548);
and U7836 (N_7836,N_7769,N_7667);
xor U7837 (N_7837,N_7679,N_7659);
xnor U7838 (N_7838,N_7688,N_7352);
nand U7839 (N_7839,N_7379,N_7369);
nor U7840 (N_7840,N_7241,N_7375);
and U7841 (N_7841,N_7732,N_7333);
xor U7842 (N_7842,N_7510,N_7508);
xnor U7843 (N_7843,N_7443,N_7437);
and U7844 (N_7844,N_7298,N_7457);
nor U7845 (N_7845,N_7645,N_7491);
nand U7846 (N_7846,N_7202,N_7662);
nor U7847 (N_7847,N_7327,N_7490);
nand U7848 (N_7848,N_7654,N_7567);
xnor U7849 (N_7849,N_7663,N_7756);
nand U7850 (N_7850,N_7294,N_7350);
nor U7851 (N_7851,N_7755,N_7455);
or U7852 (N_7852,N_7300,N_7612);
and U7853 (N_7853,N_7763,N_7317);
and U7854 (N_7854,N_7297,N_7517);
xor U7855 (N_7855,N_7699,N_7675);
xor U7856 (N_7856,N_7599,N_7210);
nor U7857 (N_7857,N_7403,N_7436);
or U7858 (N_7858,N_7246,N_7776);
xnor U7859 (N_7859,N_7545,N_7650);
nor U7860 (N_7860,N_7319,N_7523);
nand U7861 (N_7861,N_7636,N_7606);
or U7862 (N_7862,N_7604,N_7378);
nor U7863 (N_7863,N_7551,N_7334);
nand U7864 (N_7864,N_7575,N_7530);
and U7865 (N_7865,N_7313,N_7345);
and U7866 (N_7866,N_7228,N_7402);
xnor U7867 (N_7867,N_7398,N_7367);
nand U7868 (N_7868,N_7463,N_7391);
nor U7869 (N_7869,N_7503,N_7631);
nand U7870 (N_7870,N_7279,N_7435);
nand U7871 (N_7871,N_7323,N_7200);
xor U7872 (N_7872,N_7702,N_7661);
or U7873 (N_7873,N_7256,N_7261);
or U7874 (N_7874,N_7698,N_7784);
and U7875 (N_7875,N_7620,N_7539);
nor U7876 (N_7876,N_7460,N_7617);
and U7877 (N_7877,N_7277,N_7265);
xor U7878 (N_7878,N_7434,N_7586);
or U7879 (N_7879,N_7208,N_7603);
nor U7880 (N_7880,N_7534,N_7303);
or U7881 (N_7881,N_7407,N_7642);
or U7882 (N_7882,N_7427,N_7306);
or U7883 (N_7883,N_7392,N_7458);
nand U7884 (N_7884,N_7236,N_7209);
and U7885 (N_7885,N_7563,N_7415);
nand U7886 (N_7886,N_7582,N_7374);
or U7887 (N_7887,N_7632,N_7615);
or U7888 (N_7888,N_7793,N_7536);
nor U7889 (N_7889,N_7467,N_7505);
and U7890 (N_7890,N_7608,N_7640);
xnor U7891 (N_7891,N_7431,N_7232);
and U7892 (N_7892,N_7387,N_7477);
and U7893 (N_7893,N_7204,N_7358);
nand U7894 (N_7894,N_7580,N_7343);
or U7895 (N_7895,N_7328,N_7281);
and U7896 (N_7896,N_7715,N_7733);
and U7897 (N_7897,N_7238,N_7373);
nand U7898 (N_7898,N_7581,N_7653);
nor U7899 (N_7899,N_7227,N_7749);
nor U7900 (N_7900,N_7583,N_7771);
xnor U7901 (N_7901,N_7380,N_7635);
xor U7902 (N_7902,N_7600,N_7648);
nor U7903 (N_7903,N_7665,N_7476);
and U7904 (N_7904,N_7553,N_7225);
xnor U7905 (N_7905,N_7388,N_7484);
xnor U7906 (N_7906,N_7664,N_7633);
or U7907 (N_7907,N_7417,N_7518);
nor U7908 (N_7908,N_7356,N_7428);
or U7909 (N_7909,N_7201,N_7399);
and U7910 (N_7910,N_7370,N_7766);
or U7911 (N_7911,N_7721,N_7628);
and U7912 (N_7912,N_7276,N_7727);
nor U7913 (N_7913,N_7657,N_7643);
xor U7914 (N_7914,N_7322,N_7700);
or U7915 (N_7915,N_7761,N_7729);
and U7916 (N_7916,N_7479,N_7759);
xor U7917 (N_7917,N_7359,N_7789);
or U7918 (N_7918,N_7214,N_7506);
nor U7919 (N_7919,N_7411,N_7704);
and U7920 (N_7920,N_7619,N_7669);
or U7921 (N_7921,N_7708,N_7783);
and U7922 (N_7922,N_7446,N_7507);
xor U7923 (N_7923,N_7248,N_7235);
xnor U7924 (N_7924,N_7282,N_7741);
or U7925 (N_7925,N_7296,N_7357);
nand U7926 (N_7926,N_7605,N_7418);
or U7927 (N_7927,N_7532,N_7785);
xor U7928 (N_7928,N_7377,N_7709);
or U7929 (N_7929,N_7538,N_7237);
nand U7930 (N_7930,N_7487,N_7778);
nand U7931 (N_7931,N_7408,N_7651);
and U7932 (N_7932,N_7670,N_7231);
nand U7933 (N_7933,N_7430,N_7302);
nor U7934 (N_7934,N_7483,N_7469);
xor U7935 (N_7935,N_7372,N_7644);
or U7936 (N_7936,N_7737,N_7680);
and U7937 (N_7937,N_7295,N_7336);
nand U7938 (N_7938,N_7541,N_7395);
and U7939 (N_7939,N_7245,N_7416);
nor U7940 (N_7940,N_7597,N_7331);
nand U7941 (N_7941,N_7365,N_7318);
nand U7942 (N_7942,N_7254,N_7222);
or U7943 (N_7943,N_7444,N_7382);
nor U7944 (N_7944,N_7341,N_7521);
and U7945 (N_7945,N_7647,N_7462);
xnor U7946 (N_7946,N_7361,N_7572);
and U7947 (N_7947,N_7668,N_7354);
nor U7948 (N_7948,N_7305,N_7682);
nor U7949 (N_7949,N_7555,N_7316);
or U7950 (N_7950,N_7767,N_7440);
nor U7951 (N_7951,N_7747,N_7260);
nor U7952 (N_7952,N_7409,N_7384);
nor U7953 (N_7953,N_7206,N_7292);
xnor U7954 (N_7954,N_7758,N_7442);
nand U7955 (N_7955,N_7243,N_7714);
or U7956 (N_7956,N_7681,N_7230);
and U7957 (N_7957,N_7697,N_7692);
or U7958 (N_7958,N_7329,N_7742);
nand U7959 (N_7959,N_7285,N_7283);
or U7960 (N_7960,N_7393,N_7673);
nand U7961 (N_7961,N_7513,N_7671);
or U7962 (N_7962,N_7637,N_7421);
or U7963 (N_7963,N_7481,N_7516);
and U7964 (N_7964,N_7486,N_7660);
and U7965 (N_7965,N_7717,N_7270);
nand U7966 (N_7966,N_7251,N_7351);
nor U7967 (N_7967,N_7710,N_7565);
and U7968 (N_7968,N_7312,N_7683);
nand U7969 (N_7969,N_7573,N_7564);
nand U7970 (N_7970,N_7514,N_7207);
nor U7971 (N_7971,N_7610,N_7713);
or U7972 (N_7972,N_7556,N_7658);
or U7973 (N_7973,N_7788,N_7569);
nand U7974 (N_7974,N_7711,N_7579);
nand U7975 (N_7975,N_7269,N_7307);
and U7976 (N_7976,N_7730,N_7790);
or U7977 (N_7977,N_7400,N_7258);
or U7978 (N_7978,N_7638,N_7304);
nand U7979 (N_7979,N_7478,N_7308);
nor U7980 (N_7980,N_7259,N_7286);
xor U7981 (N_7981,N_7554,N_7205);
nor U7982 (N_7982,N_7578,N_7736);
and U7983 (N_7983,N_7590,N_7546);
and U7984 (N_7984,N_7796,N_7381);
or U7985 (N_7985,N_7450,N_7280);
or U7986 (N_7986,N_7346,N_7405);
nand U7987 (N_7987,N_7607,N_7371);
nor U7988 (N_7988,N_7453,N_7459);
or U7989 (N_7989,N_7456,N_7739);
xnor U7990 (N_7990,N_7275,N_7284);
or U7991 (N_7991,N_7574,N_7524);
or U7992 (N_7992,N_7509,N_7470);
nand U7993 (N_7993,N_7233,N_7649);
nand U7994 (N_7994,N_7389,N_7511);
and U7995 (N_7995,N_7433,N_7745);
and U7996 (N_7996,N_7686,N_7461);
xnor U7997 (N_7997,N_7325,N_7500);
and U7998 (N_7998,N_7482,N_7324);
xnor U7999 (N_7999,N_7311,N_7364);
and U8000 (N_8000,N_7519,N_7492);
nor U8001 (N_8001,N_7677,N_7626);
and U8002 (N_8002,N_7242,N_7687);
xor U8003 (N_8003,N_7587,N_7656);
nor U8004 (N_8004,N_7268,N_7779);
nor U8005 (N_8005,N_7754,N_7314);
nand U8006 (N_8006,N_7353,N_7255);
nor U8007 (N_8007,N_7396,N_7249);
and U8008 (N_8008,N_7684,N_7712);
and U8009 (N_8009,N_7595,N_7464);
nand U8010 (N_8010,N_7410,N_7760);
or U8011 (N_8011,N_7445,N_7383);
or U8012 (N_8012,N_7310,N_7630);
and U8013 (N_8013,N_7738,N_7768);
and U8014 (N_8014,N_7332,N_7591);
nand U8015 (N_8015,N_7439,N_7340);
xor U8016 (N_8016,N_7797,N_7531);
nor U8017 (N_8017,N_7253,N_7257);
nand U8018 (N_8018,N_7560,N_7625);
xnor U8019 (N_8019,N_7498,N_7705);
and U8020 (N_8020,N_7485,N_7674);
and U8021 (N_8021,N_7217,N_7544);
nand U8022 (N_8022,N_7547,N_7224);
and U8023 (N_8023,N_7420,N_7568);
xnor U8024 (N_8024,N_7349,N_7493);
and U8025 (N_8025,N_7321,N_7406);
and U8026 (N_8026,N_7244,N_7424);
nand U8027 (N_8027,N_7723,N_7614);
and U8028 (N_8028,N_7291,N_7229);
or U8029 (N_8029,N_7593,N_7616);
nand U8030 (N_8030,N_7691,N_7618);
and U8031 (N_8031,N_7622,N_7792);
nor U8032 (N_8032,N_7468,N_7602);
nor U8033 (N_8033,N_7753,N_7707);
nand U8034 (N_8034,N_7273,N_7360);
or U8035 (N_8035,N_7397,N_7731);
or U8036 (N_8036,N_7216,N_7474);
xor U8037 (N_8037,N_7315,N_7432);
and U8038 (N_8038,N_7786,N_7522);
xor U8039 (N_8039,N_7559,N_7696);
xor U8040 (N_8040,N_7211,N_7693);
and U8041 (N_8041,N_7278,N_7386);
or U8042 (N_8042,N_7488,N_7466);
nor U8043 (N_8043,N_7592,N_7234);
and U8044 (N_8044,N_7497,N_7471);
xnor U8045 (N_8045,N_7596,N_7777);
nand U8046 (N_8046,N_7526,N_7540);
nand U8047 (N_8047,N_7203,N_7765);
and U8048 (N_8048,N_7537,N_7775);
and U8049 (N_8049,N_7533,N_7535);
nand U8050 (N_8050,N_7390,N_7623);
xor U8051 (N_8051,N_7787,N_7743);
nand U8052 (N_8052,N_7557,N_7288);
nand U8053 (N_8053,N_7609,N_7589);
nor U8054 (N_8054,N_7355,N_7454);
xor U8055 (N_8055,N_7676,N_7448);
or U8056 (N_8056,N_7724,N_7347);
or U8057 (N_8057,N_7652,N_7264);
nor U8058 (N_8058,N_7695,N_7344);
nand U8059 (N_8059,N_7320,N_7706);
and U8060 (N_8060,N_7337,N_7746);
and U8061 (N_8061,N_7419,N_7601);
nor U8062 (N_8062,N_7561,N_7252);
or U8063 (N_8063,N_7223,N_7520);
xnor U8064 (N_8064,N_7501,N_7240);
and U8065 (N_8065,N_7781,N_7744);
xnor U8066 (N_8066,N_7499,N_7718);
xor U8067 (N_8067,N_7585,N_7465);
and U8068 (N_8068,N_7634,N_7438);
xnor U8069 (N_8069,N_7627,N_7494);
or U8070 (N_8070,N_7799,N_7740);
or U8071 (N_8071,N_7689,N_7542);
xor U8072 (N_8072,N_7734,N_7363);
nand U8073 (N_8073,N_7452,N_7690);
or U8074 (N_8074,N_7728,N_7449);
nand U8075 (N_8075,N_7226,N_7412);
nand U8076 (N_8076,N_7290,N_7576);
or U8077 (N_8077,N_7376,N_7794);
xor U8078 (N_8078,N_7512,N_7504);
and U8079 (N_8079,N_7348,N_7385);
nor U8080 (N_8080,N_7798,N_7735);
and U8081 (N_8081,N_7287,N_7266);
or U8082 (N_8082,N_7366,N_7309);
and U8083 (N_8083,N_7338,N_7326);
and U8084 (N_8084,N_7404,N_7621);
or U8085 (N_8085,N_7584,N_7720);
and U8086 (N_8086,N_7422,N_7570);
nor U8087 (N_8087,N_7558,N_7550);
or U8088 (N_8088,N_7527,N_7339);
and U8089 (N_8089,N_7773,N_7289);
nand U8090 (N_8090,N_7219,N_7262);
nor U8091 (N_8091,N_7247,N_7413);
nand U8092 (N_8092,N_7666,N_7543);
or U8093 (N_8093,N_7577,N_7566);
xor U8094 (N_8094,N_7220,N_7646);
and U8095 (N_8095,N_7722,N_7401);
xnor U8096 (N_8096,N_7703,N_7750);
nand U8097 (N_8097,N_7472,N_7293);
or U8098 (N_8098,N_7272,N_7639);
and U8099 (N_8099,N_7552,N_7528);
xnor U8100 (N_8100,N_7426,N_7711);
nand U8101 (N_8101,N_7411,N_7536);
nor U8102 (N_8102,N_7211,N_7538);
and U8103 (N_8103,N_7322,N_7684);
nand U8104 (N_8104,N_7589,N_7637);
or U8105 (N_8105,N_7240,N_7275);
and U8106 (N_8106,N_7360,N_7354);
nor U8107 (N_8107,N_7677,N_7405);
nor U8108 (N_8108,N_7795,N_7352);
or U8109 (N_8109,N_7273,N_7593);
or U8110 (N_8110,N_7322,N_7338);
nor U8111 (N_8111,N_7781,N_7389);
xor U8112 (N_8112,N_7399,N_7695);
xnor U8113 (N_8113,N_7204,N_7766);
nand U8114 (N_8114,N_7696,N_7724);
nand U8115 (N_8115,N_7297,N_7798);
nor U8116 (N_8116,N_7349,N_7602);
and U8117 (N_8117,N_7402,N_7702);
nor U8118 (N_8118,N_7576,N_7241);
nor U8119 (N_8119,N_7656,N_7705);
nor U8120 (N_8120,N_7386,N_7328);
and U8121 (N_8121,N_7758,N_7645);
nand U8122 (N_8122,N_7546,N_7222);
or U8123 (N_8123,N_7506,N_7494);
nor U8124 (N_8124,N_7238,N_7209);
xor U8125 (N_8125,N_7487,N_7692);
nand U8126 (N_8126,N_7545,N_7608);
or U8127 (N_8127,N_7736,N_7714);
nor U8128 (N_8128,N_7297,N_7291);
nor U8129 (N_8129,N_7226,N_7231);
nor U8130 (N_8130,N_7512,N_7311);
xor U8131 (N_8131,N_7532,N_7268);
nor U8132 (N_8132,N_7581,N_7434);
xnor U8133 (N_8133,N_7651,N_7392);
and U8134 (N_8134,N_7485,N_7668);
nand U8135 (N_8135,N_7740,N_7396);
xnor U8136 (N_8136,N_7691,N_7729);
xor U8137 (N_8137,N_7211,N_7705);
nor U8138 (N_8138,N_7633,N_7223);
or U8139 (N_8139,N_7710,N_7465);
or U8140 (N_8140,N_7271,N_7394);
xnor U8141 (N_8141,N_7287,N_7558);
nor U8142 (N_8142,N_7231,N_7413);
nand U8143 (N_8143,N_7258,N_7756);
nor U8144 (N_8144,N_7607,N_7402);
nor U8145 (N_8145,N_7584,N_7621);
nor U8146 (N_8146,N_7560,N_7304);
nor U8147 (N_8147,N_7784,N_7395);
xor U8148 (N_8148,N_7211,N_7323);
nand U8149 (N_8149,N_7349,N_7325);
and U8150 (N_8150,N_7688,N_7570);
nand U8151 (N_8151,N_7548,N_7255);
xor U8152 (N_8152,N_7646,N_7328);
and U8153 (N_8153,N_7619,N_7497);
nor U8154 (N_8154,N_7479,N_7400);
nor U8155 (N_8155,N_7272,N_7631);
or U8156 (N_8156,N_7724,N_7577);
xnor U8157 (N_8157,N_7752,N_7565);
nor U8158 (N_8158,N_7410,N_7275);
nor U8159 (N_8159,N_7447,N_7721);
xnor U8160 (N_8160,N_7542,N_7577);
xor U8161 (N_8161,N_7452,N_7588);
or U8162 (N_8162,N_7260,N_7336);
nor U8163 (N_8163,N_7497,N_7360);
and U8164 (N_8164,N_7627,N_7379);
and U8165 (N_8165,N_7356,N_7460);
or U8166 (N_8166,N_7253,N_7421);
xor U8167 (N_8167,N_7231,N_7463);
or U8168 (N_8168,N_7333,N_7237);
or U8169 (N_8169,N_7744,N_7727);
nand U8170 (N_8170,N_7418,N_7593);
nand U8171 (N_8171,N_7268,N_7607);
or U8172 (N_8172,N_7733,N_7709);
xor U8173 (N_8173,N_7736,N_7459);
nor U8174 (N_8174,N_7442,N_7680);
nand U8175 (N_8175,N_7306,N_7729);
nor U8176 (N_8176,N_7255,N_7400);
nor U8177 (N_8177,N_7312,N_7450);
xor U8178 (N_8178,N_7349,N_7643);
and U8179 (N_8179,N_7244,N_7228);
and U8180 (N_8180,N_7213,N_7625);
nor U8181 (N_8181,N_7432,N_7770);
xor U8182 (N_8182,N_7772,N_7454);
xnor U8183 (N_8183,N_7773,N_7713);
nand U8184 (N_8184,N_7311,N_7471);
xnor U8185 (N_8185,N_7459,N_7577);
nor U8186 (N_8186,N_7487,N_7252);
xor U8187 (N_8187,N_7236,N_7538);
or U8188 (N_8188,N_7532,N_7295);
nor U8189 (N_8189,N_7394,N_7223);
nand U8190 (N_8190,N_7493,N_7339);
nand U8191 (N_8191,N_7734,N_7563);
or U8192 (N_8192,N_7589,N_7400);
xnor U8193 (N_8193,N_7596,N_7239);
and U8194 (N_8194,N_7733,N_7253);
nor U8195 (N_8195,N_7481,N_7750);
nand U8196 (N_8196,N_7301,N_7290);
xor U8197 (N_8197,N_7562,N_7776);
nor U8198 (N_8198,N_7258,N_7302);
nor U8199 (N_8199,N_7255,N_7275);
nor U8200 (N_8200,N_7356,N_7506);
or U8201 (N_8201,N_7705,N_7228);
or U8202 (N_8202,N_7255,N_7323);
and U8203 (N_8203,N_7448,N_7738);
nor U8204 (N_8204,N_7533,N_7334);
xnor U8205 (N_8205,N_7431,N_7620);
nor U8206 (N_8206,N_7558,N_7632);
nor U8207 (N_8207,N_7512,N_7565);
or U8208 (N_8208,N_7662,N_7567);
or U8209 (N_8209,N_7213,N_7398);
or U8210 (N_8210,N_7300,N_7769);
xnor U8211 (N_8211,N_7414,N_7343);
nand U8212 (N_8212,N_7315,N_7702);
or U8213 (N_8213,N_7347,N_7509);
xnor U8214 (N_8214,N_7506,N_7332);
nand U8215 (N_8215,N_7375,N_7510);
or U8216 (N_8216,N_7788,N_7716);
xnor U8217 (N_8217,N_7562,N_7657);
and U8218 (N_8218,N_7707,N_7393);
nor U8219 (N_8219,N_7506,N_7777);
nand U8220 (N_8220,N_7253,N_7435);
nand U8221 (N_8221,N_7396,N_7509);
or U8222 (N_8222,N_7213,N_7673);
or U8223 (N_8223,N_7551,N_7577);
and U8224 (N_8224,N_7642,N_7587);
xor U8225 (N_8225,N_7455,N_7241);
or U8226 (N_8226,N_7668,N_7392);
or U8227 (N_8227,N_7453,N_7404);
xor U8228 (N_8228,N_7368,N_7208);
nand U8229 (N_8229,N_7770,N_7458);
xor U8230 (N_8230,N_7493,N_7645);
and U8231 (N_8231,N_7383,N_7479);
xor U8232 (N_8232,N_7772,N_7394);
or U8233 (N_8233,N_7548,N_7315);
or U8234 (N_8234,N_7360,N_7448);
nor U8235 (N_8235,N_7215,N_7225);
or U8236 (N_8236,N_7642,N_7557);
nor U8237 (N_8237,N_7322,N_7657);
or U8238 (N_8238,N_7479,N_7239);
nor U8239 (N_8239,N_7706,N_7764);
and U8240 (N_8240,N_7281,N_7796);
or U8241 (N_8241,N_7655,N_7506);
nor U8242 (N_8242,N_7419,N_7481);
xnor U8243 (N_8243,N_7566,N_7313);
and U8244 (N_8244,N_7716,N_7609);
nor U8245 (N_8245,N_7734,N_7489);
nor U8246 (N_8246,N_7431,N_7365);
xnor U8247 (N_8247,N_7410,N_7422);
and U8248 (N_8248,N_7679,N_7721);
or U8249 (N_8249,N_7637,N_7742);
nand U8250 (N_8250,N_7314,N_7480);
xor U8251 (N_8251,N_7793,N_7417);
nand U8252 (N_8252,N_7367,N_7401);
and U8253 (N_8253,N_7787,N_7350);
and U8254 (N_8254,N_7797,N_7689);
nand U8255 (N_8255,N_7388,N_7596);
and U8256 (N_8256,N_7524,N_7532);
and U8257 (N_8257,N_7797,N_7590);
xor U8258 (N_8258,N_7329,N_7455);
nor U8259 (N_8259,N_7414,N_7606);
nor U8260 (N_8260,N_7706,N_7399);
and U8261 (N_8261,N_7330,N_7268);
or U8262 (N_8262,N_7352,N_7644);
and U8263 (N_8263,N_7420,N_7330);
or U8264 (N_8264,N_7298,N_7631);
and U8265 (N_8265,N_7232,N_7360);
and U8266 (N_8266,N_7481,N_7435);
or U8267 (N_8267,N_7278,N_7328);
and U8268 (N_8268,N_7366,N_7704);
and U8269 (N_8269,N_7254,N_7546);
and U8270 (N_8270,N_7506,N_7778);
or U8271 (N_8271,N_7487,N_7249);
and U8272 (N_8272,N_7702,N_7289);
xor U8273 (N_8273,N_7443,N_7341);
xor U8274 (N_8274,N_7600,N_7434);
nor U8275 (N_8275,N_7527,N_7705);
xnor U8276 (N_8276,N_7531,N_7459);
or U8277 (N_8277,N_7324,N_7425);
nor U8278 (N_8278,N_7501,N_7703);
or U8279 (N_8279,N_7504,N_7418);
xor U8280 (N_8280,N_7211,N_7459);
and U8281 (N_8281,N_7728,N_7747);
xor U8282 (N_8282,N_7665,N_7525);
or U8283 (N_8283,N_7496,N_7483);
and U8284 (N_8284,N_7616,N_7548);
and U8285 (N_8285,N_7527,N_7748);
xnor U8286 (N_8286,N_7206,N_7267);
xnor U8287 (N_8287,N_7504,N_7443);
nor U8288 (N_8288,N_7684,N_7222);
nor U8289 (N_8289,N_7761,N_7684);
or U8290 (N_8290,N_7355,N_7788);
and U8291 (N_8291,N_7252,N_7670);
nor U8292 (N_8292,N_7358,N_7374);
xnor U8293 (N_8293,N_7626,N_7573);
nor U8294 (N_8294,N_7589,N_7518);
nand U8295 (N_8295,N_7564,N_7221);
xnor U8296 (N_8296,N_7649,N_7370);
nand U8297 (N_8297,N_7235,N_7433);
nand U8298 (N_8298,N_7342,N_7202);
xor U8299 (N_8299,N_7393,N_7289);
or U8300 (N_8300,N_7528,N_7677);
or U8301 (N_8301,N_7411,N_7507);
nor U8302 (N_8302,N_7338,N_7227);
and U8303 (N_8303,N_7568,N_7632);
nor U8304 (N_8304,N_7238,N_7671);
and U8305 (N_8305,N_7390,N_7315);
xor U8306 (N_8306,N_7308,N_7782);
xor U8307 (N_8307,N_7380,N_7704);
xor U8308 (N_8308,N_7570,N_7621);
or U8309 (N_8309,N_7332,N_7737);
nor U8310 (N_8310,N_7360,N_7511);
nand U8311 (N_8311,N_7565,N_7774);
xnor U8312 (N_8312,N_7406,N_7249);
nand U8313 (N_8313,N_7434,N_7369);
or U8314 (N_8314,N_7352,N_7284);
xor U8315 (N_8315,N_7479,N_7531);
xnor U8316 (N_8316,N_7483,N_7603);
and U8317 (N_8317,N_7408,N_7757);
nor U8318 (N_8318,N_7762,N_7716);
and U8319 (N_8319,N_7348,N_7417);
or U8320 (N_8320,N_7386,N_7257);
and U8321 (N_8321,N_7323,N_7389);
nor U8322 (N_8322,N_7314,N_7669);
or U8323 (N_8323,N_7410,N_7597);
nor U8324 (N_8324,N_7788,N_7677);
nand U8325 (N_8325,N_7430,N_7272);
nand U8326 (N_8326,N_7416,N_7696);
and U8327 (N_8327,N_7608,N_7590);
or U8328 (N_8328,N_7356,N_7410);
or U8329 (N_8329,N_7477,N_7397);
or U8330 (N_8330,N_7452,N_7782);
or U8331 (N_8331,N_7311,N_7501);
xnor U8332 (N_8332,N_7290,N_7420);
or U8333 (N_8333,N_7513,N_7432);
and U8334 (N_8334,N_7385,N_7245);
nor U8335 (N_8335,N_7583,N_7426);
xnor U8336 (N_8336,N_7559,N_7783);
nand U8337 (N_8337,N_7278,N_7634);
nor U8338 (N_8338,N_7266,N_7375);
xor U8339 (N_8339,N_7572,N_7320);
or U8340 (N_8340,N_7549,N_7400);
and U8341 (N_8341,N_7221,N_7239);
xnor U8342 (N_8342,N_7465,N_7562);
nand U8343 (N_8343,N_7301,N_7355);
nor U8344 (N_8344,N_7485,N_7790);
nor U8345 (N_8345,N_7657,N_7210);
or U8346 (N_8346,N_7513,N_7209);
nand U8347 (N_8347,N_7738,N_7555);
xor U8348 (N_8348,N_7584,N_7676);
nor U8349 (N_8349,N_7417,N_7495);
xor U8350 (N_8350,N_7729,N_7474);
or U8351 (N_8351,N_7766,N_7244);
or U8352 (N_8352,N_7546,N_7370);
and U8353 (N_8353,N_7609,N_7297);
and U8354 (N_8354,N_7585,N_7706);
xor U8355 (N_8355,N_7467,N_7644);
nor U8356 (N_8356,N_7659,N_7504);
and U8357 (N_8357,N_7338,N_7479);
or U8358 (N_8358,N_7793,N_7702);
nor U8359 (N_8359,N_7581,N_7681);
and U8360 (N_8360,N_7373,N_7590);
nor U8361 (N_8361,N_7238,N_7686);
or U8362 (N_8362,N_7720,N_7315);
nand U8363 (N_8363,N_7631,N_7553);
or U8364 (N_8364,N_7202,N_7639);
and U8365 (N_8365,N_7282,N_7568);
xor U8366 (N_8366,N_7510,N_7750);
or U8367 (N_8367,N_7582,N_7342);
or U8368 (N_8368,N_7590,N_7593);
xnor U8369 (N_8369,N_7459,N_7792);
nand U8370 (N_8370,N_7451,N_7264);
nand U8371 (N_8371,N_7204,N_7342);
or U8372 (N_8372,N_7766,N_7358);
or U8373 (N_8373,N_7596,N_7693);
and U8374 (N_8374,N_7293,N_7584);
xnor U8375 (N_8375,N_7340,N_7715);
nand U8376 (N_8376,N_7726,N_7571);
nor U8377 (N_8377,N_7402,N_7731);
nor U8378 (N_8378,N_7660,N_7434);
and U8379 (N_8379,N_7772,N_7584);
xnor U8380 (N_8380,N_7757,N_7279);
xor U8381 (N_8381,N_7213,N_7390);
nor U8382 (N_8382,N_7359,N_7699);
xor U8383 (N_8383,N_7283,N_7571);
nor U8384 (N_8384,N_7445,N_7391);
nand U8385 (N_8385,N_7686,N_7571);
nand U8386 (N_8386,N_7616,N_7572);
and U8387 (N_8387,N_7341,N_7618);
xor U8388 (N_8388,N_7543,N_7729);
xor U8389 (N_8389,N_7739,N_7453);
nor U8390 (N_8390,N_7460,N_7201);
and U8391 (N_8391,N_7624,N_7437);
nor U8392 (N_8392,N_7692,N_7397);
nand U8393 (N_8393,N_7629,N_7785);
xnor U8394 (N_8394,N_7390,N_7245);
or U8395 (N_8395,N_7507,N_7513);
xnor U8396 (N_8396,N_7623,N_7342);
xnor U8397 (N_8397,N_7294,N_7415);
or U8398 (N_8398,N_7700,N_7308);
or U8399 (N_8399,N_7490,N_7628);
nor U8400 (N_8400,N_8065,N_8333);
xnor U8401 (N_8401,N_8165,N_8372);
or U8402 (N_8402,N_8131,N_7855);
or U8403 (N_8403,N_7825,N_8335);
xnor U8404 (N_8404,N_7984,N_8338);
and U8405 (N_8405,N_7918,N_8116);
or U8406 (N_8406,N_8339,N_7800);
or U8407 (N_8407,N_8028,N_7922);
nor U8408 (N_8408,N_8197,N_7866);
nand U8409 (N_8409,N_8375,N_8385);
nand U8410 (N_8410,N_7864,N_7996);
or U8411 (N_8411,N_8107,N_7870);
nand U8412 (N_8412,N_8268,N_7896);
nand U8413 (N_8413,N_8363,N_8256);
nor U8414 (N_8414,N_8094,N_8216);
xnor U8415 (N_8415,N_8003,N_7813);
and U8416 (N_8416,N_8193,N_8234);
nor U8417 (N_8417,N_8013,N_7971);
and U8418 (N_8418,N_7807,N_8031);
xnor U8419 (N_8419,N_8232,N_8161);
and U8420 (N_8420,N_8045,N_8024);
nor U8421 (N_8421,N_7903,N_8389);
xor U8422 (N_8422,N_8042,N_8320);
nand U8423 (N_8423,N_8077,N_7880);
or U8424 (N_8424,N_7814,N_8285);
or U8425 (N_8425,N_8266,N_8344);
nor U8426 (N_8426,N_8006,N_8377);
and U8427 (N_8427,N_8322,N_8262);
nand U8428 (N_8428,N_8225,N_7835);
nand U8429 (N_8429,N_8257,N_7879);
and U8430 (N_8430,N_7958,N_7832);
xor U8431 (N_8431,N_7848,N_8251);
or U8432 (N_8432,N_7889,N_8088);
nor U8433 (N_8433,N_7955,N_8070);
nand U8434 (N_8434,N_8394,N_7947);
or U8435 (N_8435,N_7977,N_7821);
nor U8436 (N_8436,N_7989,N_8382);
nand U8437 (N_8437,N_8168,N_8245);
or U8438 (N_8438,N_8307,N_8215);
nor U8439 (N_8439,N_8075,N_8171);
nor U8440 (N_8440,N_8114,N_8179);
or U8441 (N_8441,N_7854,N_8093);
nor U8442 (N_8442,N_8063,N_7941);
nand U8443 (N_8443,N_8046,N_8252);
nand U8444 (N_8444,N_7904,N_8356);
and U8445 (N_8445,N_8166,N_8291);
and U8446 (N_8446,N_7925,N_8314);
nor U8447 (N_8447,N_8121,N_7822);
nand U8448 (N_8448,N_8090,N_8255);
and U8449 (N_8449,N_8352,N_8249);
nand U8450 (N_8450,N_8302,N_8124);
nand U8451 (N_8451,N_8383,N_8106);
or U8452 (N_8452,N_8250,N_8240);
and U8453 (N_8453,N_8361,N_8128);
or U8454 (N_8454,N_8136,N_8187);
xnor U8455 (N_8455,N_7956,N_8272);
nor U8456 (N_8456,N_7998,N_8364);
nand U8457 (N_8457,N_8007,N_7926);
nand U8458 (N_8458,N_8380,N_7846);
or U8459 (N_8459,N_7933,N_7884);
or U8460 (N_8460,N_7859,N_8016);
nor U8461 (N_8461,N_8032,N_7905);
nor U8462 (N_8462,N_8083,N_8157);
nand U8463 (N_8463,N_8164,N_8154);
or U8464 (N_8464,N_8306,N_8048);
nand U8465 (N_8465,N_8205,N_8125);
nand U8466 (N_8466,N_8012,N_8146);
nor U8467 (N_8467,N_8043,N_8130);
and U8468 (N_8468,N_8260,N_8297);
nand U8469 (N_8469,N_8067,N_7838);
and U8470 (N_8470,N_8156,N_7827);
nand U8471 (N_8471,N_8310,N_8284);
nand U8472 (N_8472,N_8160,N_7843);
xor U8473 (N_8473,N_8348,N_8243);
nand U8474 (N_8474,N_7873,N_8336);
and U8475 (N_8475,N_7954,N_7869);
nand U8476 (N_8476,N_8362,N_7908);
nor U8477 (N_8477,N_7802,N_8044);
and U8478 (N_8478,N_8235,N_8017);
or U8479 (N_8479,N_8064,N_8059);
nand U8480 (N_8480,N_7811,N_8370);
or U8481 (N_8481,N_7945,N_8393);
xor U8482 (N_8482,N_8230,N_8174);
nand U8483 (N_8483,N_7915,N_7979);
and U8484 (N_8484,N_7963,N_8137);
xor U8485 (N_8485,N_7853,N_8289);
xnor U8486 (N_8486,N_8217,N_7997);
or U8487 (N_8487,N_7886,N_8294);
nand U8488 (N_8488,N_7897,N_7868);
nand U8489 (N_8489,N_8169,N_8329);
nand U8490 (N_8490,N_8265,N_8060);
xnor U8491 (N_8491,N_8184,N_8180);
nor U8492 (N_8492,N_8095,N_8087);
xor U8493 (N_8493,N_8309,N_8072);
nor U8494 (N_8494,N_8143,N_8023);
nand U8495 (N_8495,N_8221,N_8145);
xor U8496 (N_8496,N_8010,N_7883);
or U8497 (N_8497,N_8376,N_8034);
nand U8498 (N_8498,N_7959,N_8279);
or U8499 (N_8499,N_8267,N_8152);
nand U8500 (N_8500,N_7965,N_8037);
or U8501 (N_8501,N_7881,N_8325);
nor U8502 (N_8502,N_8319,N_8276);
nand U8503 (N_8503,N_8055,N_7867);
or U8504 (N_8504,N_8392,N_8286);
and U8505 (N_8505,N_8273,N_8304);
nand U8506 (N_8506,N_8219,N_8354);
and U8507 (N_8507,N_8246,N_8203);
xor U8508 (N_8508,N_7919,N_8270);
or U8509 (N_8509,N_8229,N_8386);
or U8510 (N_8510,N_8355,N_7944);
and U8511 (N_8511,N_7893,N_7992);
and U8512 (N_8512,N_7983,N_7875);
or U8513 (N_8513,N_8318,N_7948);
nand U8514 (N_8514,N_8073,N_8119);
xor U8515 (N_8515,N_8275,N_8259);
or U8516 (N_8516,N_8308,N_7967);
nor U8517 (N_8517,N_8379,N_7931);
nand U8518 (N_8518,N_8122,N_7845);
xor U8519 (N_8519,N_8288,N_8258);
xnor U8520 (N_8520,N_8208,N_8030);
nand U8521 (N_8521,N_7874,N_7877);
or U8522 (N_8522,N_7999,N_7934);
and U8523 (N_8523,N_8244,N_7985);
nor U8524 (N_8524,N_8239,N_8305);
or U8525 (N_8525,N_8231,N_7840);
nand U8526 (N_8526,N_8082,N_8378);
and U8527 (N_8527,N_8212,N_8347);
xnor U8528 (N_8528,N_8029,N_8008);
and U8529 (N_8529,N_8185,N_7901);
and U8530 (N_8530,N_8141,N_8254);
xnor U8531 (N_8531,N_7966,N_8149);
and U8532 (N_8532,N_8020,N_8295);
and U8533 (N_8533,N_8147,N_8371);
or U8534 (N_8534,N_8326,N_8269);
nand U8535 (N_8535,N_7841,N_7882);
or U8536 (N_8536,N_8248,N_7852);
and U8537 (N_8537,N_7953,N_8117);
nor U8538 (N_8538,N_7913,N_7943);
nor U8539 (N_8539,N_8188,N_8102);
or U8540 (N_8540,N_7910,N_7935);
nand U8541 (N_8541,N_8190,N_8351);
xor U8542 (N_8542,N_7930,N_7824);
nor U8543 (N_8543,N_7924,N_7981);
and U8544 (N_8544,N_7842,N_8022);
or U8545 (N_8545,N_7860,N_8109);
xor U8546 (N_8546,N_8140,N_8182);
nand U8547 (N_8547,N_7892,N_7899);
xor U8548 (N_8548,N_8050,N_8224);
or U8549 (N_8549,N_8346,N_7823);
xor U8550 (N_8550,N_7865,N_8388);
nand U8551 (N_8551,N_8366,N_7833);
xor U8552 (N_8552,N_8345,N_8150);
nor U8553 (N_8553,N_8253,N_8058);
or U8554 (N_8554,N_8051,N_8177);
xnor U8555 (N_8555,N_8196,N_8039);
nor U8556 (N_8556,N_7806,N_8342);
xor U8557 (N_8557,N_8242,N_8155);
and U8558 (N_8558,N_7949,N_8237);
nand U8559 (N_8559,N_8186,N_7888);
nor U8560 (N_8560,N_7952,N_8033);
and U8561 (N_8561,N_8103,N_8298);
nor U8562 (N_8562,N_8014,N_8315);
or U8563 (N_8563,N_8038,N_8151);
or U8564 (N_8564,N_8214,N_8384);
nor U8565 (N_8565,N_7872,N_7849);
nor U8566 (N_8566,N_8066,N_8009);
nand U8567 (N_8567,N_7862,N_8391);
nand U8568 (N_8568,N_8011,N_7812);
nand U8569 (N_8569,N_8303,N_7826);
or U8570 (N_8570,N_7836,N_7885);
nor U8571 (N_8571,N_8118,N_8211);
nor U8572 (N_8572,N_8158,N_7839);
or U8573 (N_8573,N_8399,N_8316);
and U8574 (N_8574,N_7988,N_7801);
or U8575 (N_8575,N_8062,N_7817);
nand U8576 (N_8576,N_8162,N_8127);
or U8577 (N_8577,N_7891,N_8005);
xor U8578 (N_8578,N_8049,N_7994);
nand U8579 (N_8579,N_8293,N_7895);
nand U8580 (N_8580,N_8198,N_8280);
nor U8581 (N_8581,N_8281,N_7830);
nand U8582 (N_8582,N_7834,N_8101);
and U8583 (N_8583,N_8334,N_8337);
or U8584 (N_8584,N_8263,N_7973);
nor U8585 (N_8585,N_8057,N_8027);
xnor U8586 (N_8586,N_8163,N_8176);
xor U8587 (N_8587,N_8015,N_8359);
or U8588 (N_8588,N_8287,N_8173);
nor U8589 (N_8589,N_8159,N_8092);
nand U8590 (N_8590,N_8282,N_7923);
nor U8591 (N_8591,N_7847,N_8115);
and U8592 (N_8592,N_7968,N_8052);
nor U8593 (N_8593,N_7819,N_8192);
xnor U8594 (N_8594,N_7995,N_8367);
or U8595 (N_8595,N_7928,N_8021);
nor U8596 (N_8596,N_7932,N_8181);
or U8597 (N_8597,N_8189,N_7871);
and U8598 (N_8598,N_8331,N_7831);
and U8599 (N_8599,N_8387,N_8290);
and U8600 (N_8600,N_7829,N_8317);
nor U8601 (N_8601,N_8191,N_8080);
or U8602 (N_8602,N_8123,N_8133);
or U8603 (N_8603,N_8089,N_7929);
nor U8604 (N_8604,N_8278,N_8144);
xor U8605 (N_8605,N_8026,N_7916);
nand U8606 (N_8606,N_8078,N_8327);
nand U8607 (N_8607,N_7921,N_8132);
xor U8608 (N_8608,N_8202,N_7898);
nand U8609 (N_8609,N_8368,N_8301);
nor U8610 (N_8610,N_8357,N_8349);
xor U8611 (N_8611,N_8330,N_7837);
nand U8612 (N_8612,N_8068,N_7912);
nand U8613 (N_8613,N_7974,N_8096);
nor U8614 (N_8614,N_8398,N_7844);
or U8615 (N_8615,N_7951,N_8126);
and U8616 (N_8616,N_8148,N_7911);
or U8617 (N_8617,N_7818,N_8247);
xor U8618 (N_8618,N_8264,N_8227);
xor U8619 (N_8619,N_8210,N_8079);
nand U8620 (N_8620,N_8172,N_8313);
or U8621 (N_8621,N_8120,N_7856);
xor U8622 (N_8622,N_8271,N_8358);
nand U8623 (N_8623,N_8300,N_8153);
or U8624 (N_8624,N_7851,N_8274);
nand U8625 (N_8625,N_7828,N_8134);
or U8626 (N_8626,N_8194,N_7991);
nand U8627 (N_8627,N_7803,N_7815);
xor U8628 (N_8628,N_8111,N_7960);
nor U8629 (N_8629,N_7957,N_8396);
nand U8630 (N_8630,N_7976,N_7894);
nand U8631 (N_8631,N_7920,N_8129);
or U8632 (N_8632,N_8299,N_7861);
nand U8633 (N_8633,N_8110,N_8311);
nor U8634 (N_8634,N_7993,N_7964);
nand U8635 (N_8635,N_8236,N_8277);
and U8636 (N_8636,N_8204,N_8340);
nor U8637 (N_8637,N_8142,N_8195);
nor U8638 (N_8638,N_8369,N_8312);
and U8639 (N_8639,N_8040,N_7857);
xnor U8640 (N_8640,N_7902,N_8081);
or U8641 (N_8641,N_8084,N_8019);
nand U8642 (N_8642,N_8035,N_7907);
nand U8643 (N_8643,N_8213,N_7982);
nand U8644 (N_8644,N_7978,N_7878);
and U8645 (N_8645,N_7810,N_8397);
and U8646 (N_8646,N_7809,N_8332);
xnor U8647 (N_8647,N_7804,N_8098);
nor U8648 (N_8648,N_7986,N_8209);
nor U8649 (N_8649,N_8071,N_8000);
or U8650 (N_8650,N_8341,N_8199);
xnor U8651 (N_8651,N_8360,N_8086);
or U8652 (N_8652,N_8390,N_8138);
nand U8653 (N_8653,N_7942,N_8381);
or U8654 (N_8654,N_7972,N_8343);
or U8655 (N_8655,N_8324,N_7970);
nor U8656 (N_8656,N_7917,N_8222);
or U8657 (N_8657,N_7962,N_8076);
or U8658 (N_8658,N_7987,N_8167);
or U8659 (N_8659,N_8170,N_7990);
xor U8660 (N_8660,N_8292,N_7950);
xnor U8661 (N_8661,N_8074,N_8175);
and U8662 (N_8662,N_8113,N_8135);
or U8663 (N_8663,N_8099,N_8395);
or U8664 (N_8664,N_7808,N_8001);
xnor U8665 (N_8665,N_8054,N_8241);
nor U8666 (N_8666,N_8047,N_7927);
and U8667 (N_8667,N_8085,N_8061);
and U8668 (N_8668,N_8365,N_8041);
and U8669 (N_8669,N_8233,N_7940);
nor U8670 (N_8670,N_8100,N_7900);
or U8671 (N_8671,N_7939,N_7936);
or U8672 (N_8672,N_8105,N_7969);
or U8673 (N_8673,N_8200,N_8004);
xnor U8674 (N_8674,N_7820,N_8206);
or U8675 (N_8675,N_8112,N_8069);
nor U8676 (N_8676,N_8296,N_8283);
and U8677 (N_8677,N_8104,N_8036);
and U8678 (N_8678,N_8373,N_8091);
nand U8679 (N_8679,N_8056,N_8374);
nor U8680 (N_8680,N_7946,N_7906);
or U8681 (N_8681,N_8350,N_7805);
nand U8682 (N_8682,N_8328,N_7863);
nor U8683 (N_8683,N_8353,N_8097);
nor U8684 (N_8684,N_8178,N_7937);
and U8685 (N_8685,N_8139,N_8261);
xnor U8686 (N_8686,N_8223,N_8053);
nand U8687 (N_8687,N_8321,N_8218);
xnor U8688 (N_8688,N_8183,N_8323);
nor U8689 (N_8689,N_8108,N_8002);
or U8690 (N_8690,N_8228,N_7858);
xor U8691 (N_8691,N_7975,N_7938);
and U8692 (N_8692,N_8207,N_7816);
and U8693 (N_8693,N_8238,N_7876);
and U8694 (N_8694,N_7914,N_7980);
and U8695 (N_8695,N_7909,N_8201);
and U8696 (N_8696,N_8226,N_8220);
nor U8697 (N_8697,N_7961,N_7887);
nand U8698 (N_8698,N_8025,N_7850);
and U8699 (N_8699,N_8018,N_7890);
or U8700 (N_8700,N_7829,N_7941);
nor U8701 (N_8701,N_8034,N_8087);
nand U8702 (N_8702,N_7984,N_8121);
nand U8703 (N_8703,N_7896,N_8033);
and U8704 (N_8704,N_8255,N_8098);
and U8705 (N_8705,N_8074,N_7879);
or U8706 (N_8706,N_7948,N_8061);
xor U8707 (N_8707,N_8031,N_8345);
or U8708 (N_8708,N_8323,N_8262);
xor U8709 (N_8709,N_7878,N_8254);
nand U8710 (N_8710,N_7994,N_8240);
or U8711 (N_8711,N_8112,N_7899);
or U8712 (N_8712,N_8338,N_8085);
nor U8713 (N_8713,N_8373,N_8151);
nand U8714 (N_8714,N_8315,N_8017);
nor U8715 (N_8715,N_7939,N_8139);
xor U8716 (N_8716,N_7809,N_7979);
nand U8717 (N_8717,N_7843,N_8191);
and U8718 (N_8718,N_8350,N_8266);
nand U8719 (N_8719,N_7856,N_7884);
nor U8720 (N_8720,N_8330,N_8190);
or U8721 (N_8721,N_7936,N_7834);
or U8722 (N_8722,N_7979,N_7918);
and U8723 (N_8723,N_8314,N_8173);
nor U8724 (N_8724,N_8300,N_8111);
or U8725 (N_8725,N_7984,N_8000);
or U8726 (N_8726,N_8186,N_8119);
and U8727 (N_8727,N_7894,N_8070);
and U8728 (N_8728,N_8096,N_8366);
nor U8729 (N_8729,N_7914,N_7899);
nor U8730 (N_8730,N_8030,N_7801);
nor U8731 (N_8731,N_7889,N_8157);
or U8732 (N_8732,N_8348,N_8375);
nor U8733 (N_8733,N_8325,N_7867);
or U8734 (N_8734,N_8359,N_8215);
xnor U8735 (N_8735,N_8139,N_7854);
and U8736 (N_8736,N_7925,N_8062);
nand U8737 (N_8737,N_8228,N_7929);
or U8738 (N_8738,N_7899,N_7928);
and U8739 (N_8739,N_8102,N_7937);
xor U8740 (N_8740,N_8276,N_8153);
nand U8741 (N_8741,N_8163,N_8263);
or U8742 (N_8742,N_7853,N_7896);
or U8743 (N_8743,N_8245,N_8040);
nor U8744 (N_8744,N_7941,N_8142);
nand U8745 (N_8745,N_7908,N_7954);
or U8746 (N_8746,N_8240,N_8040);
and U8747 (N_8747,N_8328,N_8107);
or U8748 (N_8748,N_8328,N_7822);
nor U8749 (N_8749,N_8109,N_7986);
and U8750 (N_8750,N_8211,N_7856);
and U8751 (N_8751,N_8182,N_8167);
nand U8752 (N_8752,N_8366,N_8047);
or U8753 (N_8753,N_8399,N_8386);
nand U8754 (N_8754,N_8121,N_8221);
nand U8755 (N_8755,N_7870,N_8231);
nand U8756 (N_8756,N_8253,N_7930);
nand U8757 (N_8757,N_8309,N_7869);
nor U8758 (N_8758,N_7928,N_8339);
or U8759 (N_8759,N_8044,N_8165);
xnor U8760 (N_8760,N_8007,N_8156);
nand U8761 (N_8761,N_7964,N_8314);
nand U8762 (N_8762,N_7839,N_8115);
nand U8763 (N_8763,N_8321,N_8081);
and U8764 (N_8764,N_8064,N_7917);
and U8765 (N_8765,N_8230,N_8227);
or U8766 (N_8766,N_8063,N_7832);
and U8767 (N_8767,N_7830,N_7875);
or U8768 (N_8768,N_8125,N_7923);
or U8769 (N_8769,N_8245,N_8204);
xor U8770 (N_8770,N_8344,N_7836);
or U8771 (N_8771,N_7954,N_8077);
nand U8772 (N_8772,N_7870,N_8183);
nor U8773 (N_8773,N_8114,N_7989);
xor U8774 (N_8774,N_8356,N_7826);
nand U8775 (N_8775,N_8269,N_8129);
nor U8776 (N_8776,N_7850,N_7907);
nor U8777 (N_8777,N_7937,N_8254);
xnor U8778 (N_8778,N_8178,N_8192);
and U8779 (N_8779,N_7935,N_7862);
xnor U8780 (N_8780,N_8001,N_7918);
nand U8781 (N_8781,N_8114,N_7852);
or U8782 (N_8782,N_8158,N_8159);
xnor U8783 (N_8783,N_8329,N_8074);
or U8784 (N_8784,N_8199,N_7815);
xor U8785 (N_8785,N_8077,N_7832);
xnor U8786 (N_8786,N_8283,N_8314);
and U8787 (N_8787,N_8349,N_8306);
or U8788 (N_8788,N_8290,N_8384);
and U8789 (N_8789,N_8344,N_7933);
nand U8790 (N_8790,N_8175,N_8307);
and U8791 (N_8791,N_8296,N_7822);
nor U8792 (N_8792,N_8175,N_7986);
nand U8793 (N_8793,N_7922,N_7951);
or U8794 (N_8794,N_7988,N_8296);
or U8795 (N_8795,N_8080,N_7967);
xor U8796 (N_8796,N_8068,N_8281);
and U8797 (N_8797,N_7961,N_7938);
or U8798 (N_8798,N_7917,N_8309);
nor U8799 (N_8799,N_7859,N_7978);
or U8800 (N_8800,N_8237,N_8185);
and U8801 (N_8801,N_8261,N_7934);
nor U8802 (N_8802,N_7874,N_7837);
xor U8803 (N_8803,N_8018,N_7803);
or U8804 (N_8804,N_7950,N_8239);
xor U8805 (N_8805,N_8135,N_8024);
nand U8806 (N_8806,N_8236,N_8361);
or U8807 (N_8807,N_8010,N_8127);
nor U8808 (N_8808,N_7872,N_8317);
nor U8809 (N_8809,N_7984,N_7834);
xor U8810 (N_8810,N_8381,N_7893);
nand U8811 (N_8811,N_8396,N_8127);
nor U8812 (N_8812,N_8375,N_8043);
and U8813 (N_8813,N_8306,N_7912);
nor U8814 (N_8814,N_8045,N_8233);
xnor U8815 (N_8815,N_8326,N_7847);
nor U8816 (N_8816,N_8233,N_7861);
or U8817 (N_8817,N_8314,N_7851);
xor U8818 (N_8818,N_7859,N_8386);
nor U8819 (N_8819,N_8225,N_8293);
xnor U8820 (N_8820,N_8209,N_8340);
nand U8821 (N_8821,N_8007,N_8049);
or U8822 (N_8822,N_8244,N_7906);
nor U8823 (N_8823,N_8047,N_7891);
nor U8824 (N_8824,N_7887,N_7901);
xor U8825 (N_8825,N_8353,N_8120);
or U8826 (N_8826,N_8335,N_8227);
xnor U8827 (N_8827,N_8374,N_8394);
xor U8828 (N_8828,N_8053,N_8068);
and U8829 (N_8829,N_8343,N_8120);
nand U8830 (N_8830,N_8195,N_8085);
nor U8831 (N_8831,N_8292,N_7982);
or U8832 (N_8832,N_7834,N_7934);
nor U8833 (N_8833,N_8259,N_8095);
nand U8834 (N_8834,N_7998,N_7959);
nor U8835 (N_8835,N_8389,N_8211);
or U8836 (N_8836,N_7936,N_8292);
or U8837 (N_8837,N_7811,N_7958);
and U8838 (N_8838,N_7990,N_7828);
xor U8839 (N_8839,N_8264,N_8105);
nand U8840 (N_8840,N_8363,N_8382);
nor U8841 (N_8841,N_7971,N_7986);
xnor U8842 (N_8842,N_7847,N_8022);
and U8843 (N_8843,N_8069,N_8120);
xnor U8844 (N_8844,N_7960,N_8009);
nor U8845 (N_8845,N_8192,N_8343);
and U8846 (N_8846,N_7879,N_7804);
and U8847 (N_8847,N_8149,N_8271);
or U8848 (N_8848,N_7803,N_7850);
xor U8849 (N_8849,N_8315,N_8306);
xnor U8850 (N_8850,N_8365,N_8222);
nand U8851 (N_8851,N_8084,N_8169);
and U8852 (N_8852,N_8271,N_7845);
nand U8853 (N_8853,N_8273,N_8130);
nand U8854 (N_8854,N_8353,N_7959);
and U8855 (N_8855,N_8285,N_7815);
xnor U8856 (N_8856,N_7993,N_8084);
or U8857 (N_8857,N_8392,N_8264);
nor U8858 (N_8858,N_8339,N_7950);
or U8859 (N_8859,N_8387,N_8164);
and U8860 (N_8860,N_8105,N_7802);
xnor U8861 (N_8861,N_7891,N_8174);
or U8862 (N_8862,N_7980,N_7951);
nor U8863 (N_8863,N_7894,N_7965);
nor U8864 (N_8864,N_7855,N_8207);
xor U8865 (N_8865,N_7982,N_7831);
xor U8866 (N_8866,N_8177,N_8231);
xnor U8867 (N_8867,N_7862,N_8215);
xnor U8868 (N_8868,N_7917,N_8120);
nor U8869 (N_8869,N_7957,N_7981);
and U8870 (N_8870,N_8100,N_8222);
nand U8871 (N_8871,N_8168,N_8196);
nand U8872 (N_8872,N_7905,N_8282);
or U8873 (N_8873,N_8082,N_8193);
xor U8874 (N_8874,N_8068,N_8255);
nor U8875 (N_8875,N_8314,N_8197);
and U8876 (N_8876,N_8245,N_8311);
or U8877 (N_8877,N_7991,N_8302);
xor U8878 (N_8878,N_7949,N_7847);
xor U8879 (N_8879,N_7834,N_8074);
and U8880 (N_8880,N_8232,N_8194);
xor U8881 (N_8881,N_7876,N_8154);
nor U8882 (N_8882,N_8183,N_8372);
xor U8883 (N_8883,N_8131,N_7925);
or U8884 (N_8884,N_7953,N_7832);
or U8885 (N_8885,N_8307,N_8373);
xnor U8886 (N_8886,N_8158,N_8177);
or U8887 (N_8887,N_7969,N_7820);
and U8888 (N_8888,N_7825,N_7852);
nand U8889 (N_8889,N_8366,N_8046);
nor U8890 (N_8890,N_8241,N_8388);
or U8891 (N_8891,N_7865,N_8151);
xor U8892 (N_8892,N_8159,N_8304);
xnor U8893 (N_8893,N_8302,N_8016);
and U8894 (N_8894,N_8000,N_7850);
nor U8895 (N_8895,N_7979,N_8087);
or U8896 (N_8896,N_8181,N_7897);
and U8897 (N_8897,N_7998,N_8261);
xor U8898 (N_8898,N_7963,N_8201);
xor U8899 (N_8899,N_8045,N_8170);
or U8900 (N_8900,N_7977,N_8198);
xnor U8901 (N_8901,N_7859,N_8234);
xor U8902 (N_8902,N_8051,N_8072);
or U8903 (N_8903,N_7815,N_8195);
nand U8904 (N_8904,N_8286,N_7853);
xor U8905 (N_8905,N_7810,N_7827);
xnor U8906 (N_8906,N_8307,N_7975);
and U8907 (N_8907,N_7928,N_8277);
nor U8908 (N_8908,N_8330,N_8065);
and U8909 (N_8909,N_8180,N_8043);
nor U8910 (N_8910,N_8397,N_8188);
nor U8911 (N_8911,N_8103,N_8343);
xnor U8912 (N_8912,N_7846,N_7924);
and U8913 (N_8913,N_8077,N_8341);
or U8914 (N_8914,N_8242,N_7992);
or U8915 (N_8915,N_8169,N_7859);
nand U8916 (N_8916,N_8045,N_8112);
or U8917 (N_8917,N_7869,N_8386);
or U8918 (N_8918,N_7899,N_7871);
and U8919 (N_8919,N_7898,N_8132);
or U8920 (N_8920,N_7803,N_8115);
xor U8921 (N_8921,N_7973,N_7972);
and U8922 (N_8922,N_7982,N_8391);
or U8923 (N_8923,N_8083,N_8345);
nor U8924 (N_8924,N_7808,N_8338);
nor U8925 (N_8925,N_8185,N_8027);
nor U8926 (N_8926,N_7978,N_7820);
xor U8927 (N_8927,N_8062,N_8281);
or U8928 (N_8928,N_8183,N_7955);
xor U8929 (N_8929,N_8347,N_7861);
nor U8930 (N_8930,N_8134,N_7971);
xor U8931 (N_8931,N_8127,N_8160);
xnor U8932 (N_8932,N_8118,N_8166);
or U8933 (N_8933,N_8310,N_8015);
nor U8934 (N_8934,N_8369,N_8066);
and U8935 (N_8935,N_7885,N_8265);
nor U8936 (N_8936,N_7837,N_7904);
nand U8937 (N_8937,N_8007,N_7823);
or U8938 (N_8938,N_8278,N_8348);
and U8939 (N_8939,N_8246,N_8098);
nand U8940 (N_8940,N_7984,N_7963);
xor U8941 (N_8941,N_8352,N_7954);
nand U8942 (N_8942,N_8272,N_8270);
nand U8943 (N_8943,N_8137,N_8195);
nand U8944 (N_8944,N_8010,N_7846);
xor U8945 (N_8945,N_8048,N_8076);
nand U8946 (N_8946,N_8377,N_8310);
xnor U8947 (N_8947,N_8334,N_8379);
xor U8948 (N_8948,N_8245,N_8387);
nand U8949 (N_8949,N_7871,N_8238);
and U8950 (N_8950,N_7958,N_8203);
and U8951 (N_8951,N_8194,N_7975);
xor U8952 (N_8952,N_7930,N_7848);
nand U8953 (N_8953,N_7923,N_8259);
and U8954 (N_8954,N_7960,N_8344);
or U8955 (N_8955,N_8155,N_7913);
nor U8956 (N_8956,N_8324,N_8278);
nand U8957 (N_8957,N_8151,N_8336);
xor U8958 (N_8958,N_8381,N_7999);
and U8959 (N_8959,N_7859,N_8125);
and U8960 (N_8960,N_7997,N_8381);
nor U8961 (N_8961,N_8238,N_7917);
nand U8962 (N_8962,N_8219,N_8355);
nor U8963 (N_8963,N_7942,N_8322);
xnor U8964 (N_8964,N_8013,N_8374);
nand U8965 (N_8965,N_8186,N_8321);
or U8966 (N_8966,N_8019,N_8022);
and U8967 (N_8967,N_8129,N_8378);
nor U8968 (N_8968,N_7947,N_7992);
xor U8969 (N_8969,N_8016,N_7881);
nand U8970 (N_8970,N_7858,N_7805);
xor U8971 (N_8971,N_8148,N_8275);
and U8972 (N_8972,N_8197,N_8037);
or U8973 (N_8973,N_8241,N_8266);
nand U8974 (N_8974,N_7873,N_8366);
and U8975 (N_8975,N_8321,N_7885);
and U8976 (N_8976,N_8162,N_8051);
or U8977 (N_8977,N_8057,N_8096);
xnor U8978 (N_8978,N_8383,N_7882);
xnor U8979 (N_8979,N_7860,N_8032);
and U8980 (N_8980,N_8167,N_8232);
nand U8981 (N_8981,N_7808,N_8130);
nor U8982 (N_8982,N_7853,N_8121);
xor U8983 (N_8983,N_8177,N_8243);
xnor U8984 (N_8984,N_7823,N_8177);
and U8985 (N_8985,N_8129,N_7930);
nor U8986 (N_8986,N_7965,N_8069);
nand U8987 (N_8987,N_7970,N_8054);
nand U8988 (N_8988,N_8269,N_8085);
xnor U8989 (N_8989,N_7849,N_8381);
or U8990 (N_8990,N_8366,N_7999);
xor U8991 (N_8991,N_8183,N_8235);
xnor U8992 (N_8992,N_8299,N_8130);
and U8993 (N_8993,N_8022,N_7865);
or U8994 (N_8994,N_7818,N_8126);
and U8995 (N_8995,N_7843,N_7810);
and U8996 (N_8996,N_8025,N_8041);
xnor U8997 (N_8997,N_8341,N_7858);
and U8998 (N_8998,N_7931,N_8030);
xor U8999 (N_8999,N_7933,N_8155);
and U9000 (N_9000,N_8919,N_8638);
nand U9001 (N_9001,N_8460,N_8504);
and U9002 (N_9002,N_8535,N_8511);
or U9003 (N_9003,N_8680,N_8846);
and U9004 (N_9004,N_8952,N_8814);
and U9005 (N_9005,N_8906,N_8736);
nor U9006 (N_9006,N_8608,N_8982);
and U9007 (N_9007,N_8577,N_8762);
xnor U9008 (N_9008,N_8611,N_8921);
nor U9009 (N_9009,N_8813,N_8594);
nor U9010 (N_9010,N_8918,N_8439);
nand U9011 (N_9011,N_8849,N_8667);
xor U9012 (N_9012,N_8576,N_8865);
nor U9013 (N_9013,N_8668,N_8490);
nand U9014 (N_9014,N_8602,N_8796);
and U9015 (N_9015,N_8695,N_8420);
and U9016 (N_9016,N_8791,N_8761);
xor U9017 (N_9017,N_8842,N_8401);
or U9018 (N_9018,N_8689,N_8558);
and U9019 (N_9019,N_8973,N_8896);
xnor U9020 (N_9020,N_8400,N_8655);
nand U9021 (N_9021,N_8531,N_8549);
and U9022 (N_9022,N_8542,N_8769);
nand U9023 (N_9023,N_8752,N_8725);
nor U9024 (N_9024,N_8671,N_8845);
or U9025 (N_9025,N_8673,N_8800);
and U9026 (N_9026,N_8884,N_8651);
xnor U9027 (N_9027,N_8749,N_8471);
xnor U9028 (N_9028,N_8678,N_8719);
nor U9029 (N_9029,N_8585,N_8710);
nor U9030 (N_9030,N_8767,N_8771);
xor U9031 (N_9031,N_8459,N_8751);
nor U9032 (N_9032,N_8830,N_8886);
nor U9033 (N_9033,N_8766,N_8850);
xor U9034 (N_9034,N_8709,N_8554);
and U9035 (N_9035,N_8835,N_8499);
xor U9036 (N_9036,N_8449,N_8496);
or U9037 (N_9037,N_8652,N_8661);
xor U9038 (N_9038,N_8534,N_8741);
or U9039 (N_9039,N_8819,N_8505);
nor U9040 (N_9040,N_8684,N_8702);
xor U9041 (N_9041,N_8546,N_8917);
and U9042 (N_9042,N_8979,N_8737);
or U9043 (N_9043,N_8625,N_8959);
xor U9044 (N_9044,N_8871,N_8698);
nand U9045 (N_9045,N_8786,N_8616);
and U9046 (N_9046,N_8501,N_8561);
nand U9047 (N_9047,N_8488,N_8507);
nor U9048 (N_9048,N_8448,N_8636);
or U9049 (N_9049,N_8923,N_8729);
nor U9050 (N_9050,N_8432,N_8985);
nor U9051 (N_9051,N_8408,N_8980);
and U9052 (N_9052,N_8885,N_8949);
or U9053 (N_9053,N_8634,N_8453);
xnor U9054 (N_9054,N_8848,N_8747);
and U9055 (N_9055,N_8628,N_8415);
and U9056 (N_9056,N_8669,N_8722);
or U9057 (N_9057,N_8847,N_8508);
and U9058 (N_9058,N_8656,N_8431);
nand U9059 (N_9059,N_8553,N_8863);
or U9060 (N_9060,N_8828,N_8640);
and U9061 (N_9061,N_8824,N_8476);
nand U9062 (N_9062,N_8509,N_8545);
xor U9063 (N_9063,N_8880,N_8853);
xnor U9064 (N_9064,N_8468,N_8579);
and U9065 (N_9065,N_8475,N_8569);
and U9066 (N_9066,N_8570,N_8650);
or U9067 (N_9067,N_8797,N_8765);
or U9068 (N_9068,N_8404,N_8861);
or U9069 (N_9069,N_8962,N_8993);
nor U9070 (N_9070,N_8944,N_8816);
or U9071 (N_9071,N_8890,N_8901);
nor U9072 (N_9072,N_8532,N_8900);
nor U9073 (N_9073,N_8739,N_8954);
and U9074 (N_9074,N_8455,N_8812);
nand U9075 (N_9075,N_8473,N_8615);
nor U9076 (N_9076,N_8539,N_8868);
nand U9077 (N_9077,N_8986,N_8688);
or U9078 (N_9078,N_8726,N_8551);
nor U9079 (N_9079,N_8687,N_8773);
nor U9080 (N_9080,N_8493,N_8412);
nand U9081 (N_9081,N_8984,N_8734);
xnor U9082 (N_9082,N_8754,N_8596);
and U9083 (N_9083,N_8435,N_8706);
xor U9084 (N_9084,N_8823,N_8945);
and U9085 (N_9085,N_8785,N_8595);
and U9086 (N_9086,N_8555,N_8593);
xnor U9087 (N_9087,N_8931,N_8907);
xor U9088 (N_9088,N_8426,N_8443);
xor U9089 (N_9089,N_8755,N_8604);
or U9090 (N_9090,N_8676,N_8990);
and U9091 (N_9091,N_8597,N_8793);
and U9092 (N_9092,N_8855,N_8735);
or U9093 (N_9093,N_8416,N_8694);
nor U9094 (N_9094,N_8920,N_8815);
nor U9095 (N_9095,N_8529,N_8905);
nor U9096 (N_9096,N_8712,N_8502);
nor U9097 (N_9097,N_8701,N_8929);
and U9098 (N_9098,N_8926,N_8746);
and U9099 (N_9099,N_8480,N_8789);
and U9100 (N_9100,N_8512,N_8924);
xnor U9101 (N_9101,N_8631,N_8756);
xor U9102 (N_9102,N_8575,N_8707);
or U9103 (N_9103,N_8744,N_8866);
or U9104 (N_9104,N_8753,N_8467);
and U9105 (N_9105,N_8682,N_8566);
or U9106 (N_9106,N_8792,N_8444);
or U9107 (N_9107,N_8913,N_8544);
nor U9108 (N_9108,N_8413,N_8659);
nor U9109 (N_9109,N_8647,N_8437);
xnor U9110 (N_9110,N_8888,N_8700);
xor U9111 (N_9111,N_8732,N_8728);
and U9112 (N_9112,N_8515,N_8718);
nor U9113 (N_9113,N_8930,N_8599);
or U9114 (N_9114,N_8434,N_8521);
nor U9115 (N_9115,N_8881,N_8810);
xor U9116 (N_9116,N_8510,N_8469);
xnor U9117 (N_9117,N_8564,N_8450);
nor U9118 (N_9118,N_8821,N_8967);
xor U9119 (N_9119,N_8902,N_8981);
or U9120 (N_9120,N_8870,N_8768);
nor U9121 (N_9121,N_8742,N_8581);
nor U9122 (N_9122,N_8914,N_8430);
or U9123 (N_9123,N_8548,N_8658);
nor U9124 (N_9124,N_8903,N_8626);
nor U9125 (N_9125,N_8939,N_8983);
nand U9126 (N_9126,N_8692,N_8715);
xor U9127 (N_9127,N_8748,N_8573);
and U9128 (N_9128,N_8567,N_8988);
nand U9129 (N_9129,N_8470,N_8418);
xnor U9130 (N_9130,N_8780,N_8965);
or U9131 (N_9131,N_8811,N_8464);
nor U9132 (N_9132,N_8612,N_8831);
and U9133 (N_9133,N_8481,N_8740);
nor U9134 (N_9134,N_8825,N_8927);
and U9135 (N_9135,N_8803,N_8759);
nand U9136 (N_9136,N_8911,N_8966);
and U9137 (N_9137,N_8491,N_8827);
nand U9138 (N_9138,N_8937,N_8820);
and U9139 (N_9139,N_8424,N_8497);
xnor U9140 (N_9140,N_8971,N_8910);
nand U9141 (N_9141,N_8590,N_8589);
or U9142 (N_9142,N_8660,N_8841);
and U9143 (N_9143,N_8518,N_8969);
or U9144 (N_9144,N_8843,N_8889);
or U9145 (N_9145,N_8869,N_8500);
or U9146 (N_9146,N_8711,N_8898);
nor U9147 (N_9147,N_8445,N_8644);
xnor U9148 (N_9148,N_8617,N_8807);
and U9149 (N_9149,N_8557,N_8957);
or U9150 (N_9150,N_8801,N_8428);
nand U9151 (N_9151,N_8516,N_8991);
xor U9152 (N_9152,N_8723,N_8601);
nor U9153 (N_9153,N_8458,N_8614);
nor U9154 (N_9154,N_8419,N_8600);
and U9155 (N_9155,N_8916,N_8536);
nand U9156 (N_9156,N_8730,N_8506);
nor U9157 (N_9157,N_8696,N_8943);
nor U9158 (N_9158,N_8887,N_8685);
and U9159 (N_9159,N_8528,N_8764);
or U9160 (N_9160,N_8717,N_8583);
nor U9161 (N_9161,N_8461,N_8524);
and U9162 (N_9162,N_8859,N_8837);
or U9163 (N_9163,N_8895,N_8790);
and U9164 (N_9164,N_8619,N_8621);
or U9165 (N_9165,N_8877,N_8513);
nand U9166 (N_9166,N_8520,N_8477);
or U9167 (N_9167,N_8699,N_8844);
or U9168 (N_9168,N_8787,N_8757);
nand U9169 (N_9169,N_8484,N_8955);
and U9170 (N_9170,N_8964,N_8677);
xor U9171 (N_9171,N_8750,N_8832);
nand U9172 (N_9172,N_8494,N_8587);
or U9173 (N_9173,N_8873,N_8975);
and U9174 (N_9174,N_8995,N_8406);
and U9175 (N_9175,N_8833,N_8864);
and U9176 (N_9176,N_8879,N_8703);
nor U9177 (N_9177,N_8654,N_8635);
nor U9178 (N_9178,N_8568,N_8526);
nand U9179 (N_9179,N_8578,N_8904);
xnor U9180 (N_9180,N_8433,N_8463);
nand U9181 (N_9181,N_8643,N_8618);
xnor U9182 (N_9182,N_8666,N_8860);
nor U9183 (N_9183,N_8998,N_8857);
xnor U9184 (N_9184,N_8407,N_8795);
nor U9185 (N_9185,N_8485,N_8425);
and U9186 (N_9186,N_8999,N_8645);
nor U9187 (N_9187,N_8519,N_8486);
nand U9188 (N_9188,N_8641,N_8883);
nor U9189 (N_9189,N_8708,N_8851);
and U9190 (N_9190,N_8478,N_8947);
or U9191 (N_9191,N_8716,N_8705);
xor U9192 (N_9192,N_8552,N_8514);
nor U9193 (N_9193,N_8987,N_8953);
nand U9194 (N_9194,N_8540,N_8670);
xnor U9195 (N_9195,N_8452,N_8745);
and U9196 (N_9196,N_8892,N_8472);
xor U9197 (N_9197,N_8648,N_8805);
nand U9198 (N_9198,N_8775,N_8778);
nand U9199 (N_9199,N_8958,N_8598);
nand U9200 (N_9200,N_8838,N_8405);
nand U9201 (N_9201,N_8456,N_8808);
or U9202 (N_9202,N_8622,N_8961);
nand U9203 (N_9203,N_8427,N_8487);
xor U9204 (N_9204,N_8411,N_8674);
or U9205 (N_9205,N_8779,N_8683);
xor U9206 (N_9206,N_8731,N_8530);
nand U9207 (N_9207,N_8799,N_8776);
and U9208 (N_9208,N_8533,N_8642);
nand U9209 (N_9209,N_8922,N_8421);
nand U9210 (N_9210,N_8690,N_8956);
or U9211 (N_9211,N_8950,N_8894);
and U9212 (N_9212,N_8479,N_8629);
nand U9213 (N_9213,N_8992,N_8550);
nand U9214 (N_9214,N_8720,N_8454);
nand U9215 (N_9215,N_8727,N_8862);
or U9216 (N_9216,N_8942,N_8940);
or U9217 (N_9217,N_8525,N_8681);
xor U9218 (N_9218,N_8936,N_8760);
nor U9219 (N_9219,N_8482,N_8704);
and U9220 (N_9220,N_8462,N_8733);
xor U9221 (N_9221,N_8657,N_8743);
nand U9222 (N_9222,N_8409,N_8951);
nand U9223 (N_9223,N_8562,N_8977);
and U9224 (N_9224,N_8996,N_8770);
xnor U9225 (N_9225,N_8442,N_8414);
or U9226 (N_9226,N_8788,N_8909);
and U9227 (N_9227,N_8836,N_8686);
nand U9228 (N_9228,N_8802,N_8782);
nor U9229 (N_9229,N_8438,N_8772);
or U9230 (N_9230,N_8466,N_8817);
or U9231 (N_9231,N_8968,N_8784);
nor U9232 (N_9232,N_8517,N_8932);
nand U9233 (N_9233,N_8875,N_8403);
nand U9234 (N_9234,N_8609,N_8649);
xnor U9235 (N_9235,N_8697,N_8465);
nand U9236 (N_9236,N_8798,N_8925);
nand U9237 (N_9237,N_8429,N_8829);
or U9238 (N_9238,N_8826,N_8994);
or U9239 (N_9239,N_8970,N_8627);
nand U9240 (N_9240,N_8665,N_8447);
or U9241 (N_9241,N_8582,N_8989);
nand U9242 (N_9242,N_8915,N_8624);
nand U9243 (N_9243,N_8560,N_8498);
or U9244 (N_9244,N_8818,N_8897);
xnor U9245 (N_9245,N_8809,N_8457);
xnor U9246 (N_9246,N_8781,N_8653);
nand U9247 (N_9247,N_8423,N_8928);
nand U9248 (N_9248,N_8783,N_8948);
xnor U9249 (N_9249,N_8483,N_8446);
nor U9250 (N_9250,N_8410,N_8946);
nor U9251 (N_9251,N_8672,N_8876);
and U9252 (N_9252,N_8559,N_8899);
nor U9253 (N_9253,N_8632,N_8933);
nor U9254 (N_9254,N_8997,N_8503);
and U9255 (N_9255,N_8592,N_8417);
or U9256 (N_9256,N_8547,N_8572);
or U9257 (N_9257,N_8588,N_8663);
xnor U9258 (N_9258,N_8804,N_8522);
xor U9259 (N_9259,N_8440,N_8607);
or U9260 (N_9260,N_8623,N_8978);
xor U9261 (N_9261,N_8637,N_8822);
nand U9262 (N_9262,N_8495,N_8774);
and U9263 (N_9263,N_8664,N_8758);
nor U9264 (N_9264,N_8935,N_8858);
nand U9265 (N_9265,N_8537,N_8834);
nand U9266 (N_9266,N_8941,N_8639);
or U9267 (N_9267,N_8840,N_8794);
nand U9268 (N_9268,N_8527,N_8839);
nor U9269 (N_9269,N_8620,N_8972);
or U9270 (N_9270,N_8422,N_8960);
nand U9271 (N_9271,N_8724,N_8974);
nor U9272 (N_9272,N_8586,N_8714);
nor U9273 (N_9273,N_8436,N_8854);
nor U9274 (N_9274,N_8451,N_8713);
or U9275 (N_9275,N_8523,N_8606);
nand U9276 (N_9276,N_8610,N_8402);
nor U9277 (N_9277,N_8675,N_8912);
nand U9278 (N_9278,N_8691,N_8679);
and U9279 (N_9279,N_8882,N_8878);
nor U9280 (N_9280,N_8806,N_8693);
and U9281 (N_9281,N_8605,N_8613);
or U9282 (N_9282,N_8538,N_8630);
xnor U9283 (N_9283,N_8556,N_8721);
nor U9284 (N_9284,N_8646,N_8867);
and U9285 (N_9285,N_8738,N_8893);
nand U9286 (N_9286,N_8633,N_8584);
xnor U9287 (N_9287,N_8489,N_8934);
nand U9288 (N_9288,N_8563,N_8763);
nand U9289 (N_9289,N_8852,N_8441);
and U9290 (N_9290,N_8591,N_8908);
nor U9291 (N_9291,N_8777,N_8938);
nor U9292 (N_9292,N_8580,N_8603);
nand U9293 (N_9293,N_8565,N_8874);
xor U9294 (N_9294,N_8474,N_8571);
or U9295 (N_9295,N_8963,N_8662);
nor U9296 (N_9296,N_8492,N_8574);
or U9297 (N_9297,N_8891,N_8543);
nor U9298 (N_9298,N_8976,N_8856);
nor U9299 (N_9299,N_8541,N_8872);
or U9300 (N_9300,N_8799,N_8791);
or U9301 (N_9301,N_8709,N_8520);
xnor U9302 (N_9302,N_8853,N_8839);
xor U9303 (N_9303,N_8985,N_8553);
xor U9304 (N_9304,N_8939,N_8810);
and U9305 (N_9305,N_8668,N_8752);
nand U9306 (N_9306,N_8684,N_8655);
and U9307 (N_9307,N_8536,N_8782);
or U9308 (N_9308,N_8439,N_8472);
nand U9309 (N_9309,N_8506,N_8902);
or U9310 (N_9310,N_8587,N_8408);
nand U9311 (N_9311,N_8946,N_8856);
nand U9312 (N_9312,N_8519,N_8692);
nand U9313 (N_9313,N_8996,N_8861);
or U9314 (N_9314,N_8968,N_8403);
nand U9315 (N_9315,N_8944,N_8474);
xor U9316 (N_9316,N_8515,N_8756);
or U9317 (N_9317,N_8701,N_8472);
nor U9318 (N_9318,N_8825,N_8705);
or U9319 (N_9319,N_8905,N_8640);
nand U9320 (N_9320,N_8662,N_8938);
and U9321 (N_9321,N_8423,N_8501);
nor U9322 (N_9322,N_8451,N_8411);
or U9323 (N_9323,N_8824,N_8996);
nand U9324 (N_9324,N_8811,N_8829);
or U9325 (N_9325,N_8965,N_8726);
or U9326 (N_9326,N_8835,N_8874);
xnor U9327 (N_9327,N_8820,N_8428);
xor U9328 (N_9328,N_8637,N_8839);
nor U9329 (N_9329,N_8815,N_8886);
or U9330 (N_9330,N_8492,N_8469);
xor U9331 (N_9331,N_8631,N_8809);
or U9332 (N_9332,N_8513,N_8935);
or U9333 (N_9333,N_8926,N_8692);
nand U9334 (N_9334,N_8835,N_8921);
nand U9335 (N_9335,N_8789,N_8525);
and U9336 (N_9336,N_8580,N_8855);
or U9337 (N_9337,N_8660,N_8790);
or U9338 (N_9338,N_8511,N_8714);
nor U9339 (N_9339,N_8918,N_8722);
and U9340 (N_9340,N_8997,N_8597);
nor U9341 (N_9341,N_8626,N_8740);
or U9342 (N_9342,N_8412,N_8415);
or U9343 (N_9343,N_8590,N_8910);
nand U9344 (N_9344,N_8912,N_8608);
or U9345 (N_9345,N_8444,N_8505);
nand U9346 (N_9346,N_8843,N_8466);
nor U9347 (N_9347,N_8717,N_8837);
nor U9348 (N_9348,N_8501,N_8877);
xor U9349 (N_9349,N_8492,N_8579);
and U9350 (N_9350,N_8757,N_8675);
nand U9351 (N_9351,N_8953,N_8472);
or U9352 (N_9352,N_8430,N_8805);
nand U9353 (N_9353,N_8576,N_8668);
and U9354 (N_9354,N_8621,N_8921);
or U9355 (N_9355,N_8648,N_8692);
xnor U9356 (N_9356,N_8418,N_8548);
nand U9357 (N_9357,N_8601,N_8569);
xnor U9358 (N_9358,N_8556,N_8643);
or U9359 (N_9359,N_8417,N_8678);
and U9360 (N_9360,N_8540,N_8501);
and U9361 (N_9361,N_8502,N_8919);
and U9362 (N_9362,N_8759,N_8873);
xor U9363 (N_9363,N_8872,N_8581);
nand U9364 (N_9364,N_8597,N_8411);
and U9365 (N_9365,N_8765,N_8888);
xor U9366 (N_9366,N_8685,N_8412);
xnor U9367 (N_9367,N_8744,N_8425);
nor U9368 (N_9368,N_8696,N_8794);
or U9369 (N_9369,N_8730,N_8603);
xnor U9370 (N_9370,N_8437,N_8788);
xor U9371 (N_9371,N_8471,N_8689);
and U9372 (N_9372,N_8942,N_8614);
or U9373 (N_9373,N_8611,N_8577);
nand U9374 (N_9374,N_8879,N_8814);
and U9375 (N_9375,N_8674,N_8963);
or U9376 (N_9376,N_8602,N_8888);
nand U9377 (N_9377,N_8743,N_8481);
nand U9378 (N_9378,N_8889,N_8696);
nor U9379 (N_9379,N_8795,N_8522);
nand U9380 (N_9380,N_8755,N_8853);
and U9381 (N_9381,N_8584,N_8759);
nor U9382 (N_9382,N_8647,N_8616);
nand U9383 (N_9383,N_8553,N_8851);
xnor U9384 (N_9384,N_8894,N_8743);
xor U9385 (N_9385,N_8559,N_8608);
or U9386 (N_9386,N_8867,N_8753);
xor U9387 (N_9387,N_8966,N_8671);
xnor U9388 (N_9388,N_8845,N_8922);
nand U9389 (N_9389,N_8982,N_8841);
and U9390 (N_9390,N_8896,N_8603);
nand U9391 (N_9391,N_8882,N_8648);
and U9392 (N_9392,N_8552,N_8729);
nand U9393 (N_9393,N_8694,N_8706);
nor U9394 (N_9394,N_8570,N_8461);
and U9395 (N_9395,N_8847,N_8811);
or U9396 (N_9396,N_8871,N_8485);
and U9397 (N_9397,N_8948,N_8561);
nand U9398 (N_9398,N_8400,N_8610);
and U9399 (N_9399,N_8768,N_8767);
or U9400 (N_9400,N_8463,N_8796);
nor U9401 (N_9401,N_8420,N_8453);
nor U9402 (N_9402,N_8618,N_8657);
nor U9403 (N_9403,N_8844,N_8541);
or U9404 (N_9404,N_8494,N_8746);
xnor U9405 (N_9405,N_8475,N_8831);
nor U9406 (N_9406,N_8814,N_8701);
and U9407 (N_9407,N_8789,N_8786);
xnor U9408 (N_9408,N_8511,N_8939);
nor U9409 (N_9409,N_8767,N_8427);
and U9410 (N_9410,N_8851,N_8967);
nand U9411 (N_9411,N_8876,N_8547);
or U9412 (N_9412,N_8434,N_8653);
nor U9413 (N_9413,N_8719,N_8454);
xnor U9414 (N_9414,N_8580,N_8492);
or U9415 (N_9415,N_8439,N_8535);
nor U9416 (N_9416,N_8429,N_8537);
nand U9417 (N_9417,N_8787,N_8747);
nand U9418 (N_9418,N_8958,N_8445);
or U9419 (N_9419,N_8775,N_8636);
or U9420 (N_9420,N_8940,N_8505);
nand U9421 (N_9421,N_8714,N_8472);
and U9422 (N_9422,N_8628,N_8990);
xnor U9423 (N_9423,N_8701,N_8768);
xnor U9424 (N_9424,N_8851,N_8837);
or U9425 (N_9425,N_8620,N_8697);
and U9426 (N_9426,N_8816,N_8929);
nand U9427 (N_9427,N_8455,N_8692);
nand U9428 (N_9428,N_8776,N_8678);
nand U9429 (N_9429,N_8895,N_8743);
nand U9430 (N_9430,N_8901,N_8932);
nand U9431 (N_9431,N_8415,N_8986);
nand U9432 (N_9432,N_8632,N_8735);
xor U9433 (N_9433,N_8704,N_8977);
nor U9434 (N_9434,N_8774,N_8699);
nand U9435 (N_9435,N_8532,N_8590);
nand U9436 (N_9436,N_8516,N_8575);
nand U9437 (N_9437,N_8539,N_8442);
and U9438 (N_9438,N_8964,N_8822);
nor U9439 (N_9439,N_8664,N_8683);
nand U9440 (N_9440,N_8771,N_8765);
nor U9441 (N_9441,N_8818,N_8822);
and U9442 (N_9442,N_8998,N_8599);
xor U9443 (N_9443,N_8930,N_8909);
nor U9444 (N_9444,N_8699,N_8967);
nand U9445 (N_9445,N_8871,N_8639);
nor U9446 (N_9446,N_8692,N_8587);
nand U9447 (N_9447,N_8635,N_8804);
xor U9448 (N_9448,N_8563,N_8529);
nor U9449 (N_9449,N_8772,N_8419);
nand U9450 (N_9450,N_8679,N_8566);
xnor U9451 (N_9451,N_8886,N_8509);
nor U9452 (N_9452,N_8923,N_8678);
and U9453 (N_9453,N_8589,N_8594);
nor U9454 (N_9454,N_8567,N_8899);
nand U9455 (N_9455,N_8846,N_8405);
nor U9456 (N_9456,N_8993,N_8849);
xor U9457 (N_9457,N_8456,N_8560);
nor U9458 (N_9458,N_8850,N_8564);
nand U9459 (N_9459,N_8724,N_8950);
or U9460 (N_9460,N_8452,N_8449);
nand U9461 (N_9461,N_8520,N_8766);
or U9462 (N_9462,N_8931,N_8795);
and U9463 (N_9463,N_8936,N_8521);
nand U9464 (N_9464,N_8634,N_8652);
and U9465 (N_9465,N_8990,N_8962);
or U9466 (N_9466,N_8647,N_8506);
nand U9467 (N_9467,N_8837,N_8875);
nor U9468 (N_9468,N_8603,N_8970);
nor U9469 (N_9469,N_8629,N_8494);
nand U9470 (N_9470,N_8973,N_8796);
nand U9471 (N_9471,N_8626,N_8698);
nor U9472 (N_9472,N_8589,N_8729);
or U9473 (N_9473,N_8662,N_8481);
and U9474 (N_9474,N_8712,N_8998);
and U9475 (N_9475,N_8733,N_8907);
xnor U9476 (N_9476,N_8728,N_8941);
xor U9477 (N_9477,N_8606,N_8966);
or U9478 (N_9478,N_8408,N_8681);
nand U9479 (N_9479,N_8869,N_8677);
xor U9480 (N_9480,N_8596,N_8864);
nor U9481 (N_9481,N_8484,N_8535);
or U9482 (N_9482,N_8756,N_8814);
and U9483 (N_9483,N_8463,N_8591);
xnor U9484 (N_9484,N_8893,N_8682);
nand U9485 (N_9485,N_8518,N_8938);
nand U9486 (N_9486,N_8829,N_8806);
nand U9487 (N_9487,N_8698,N_8473);
or U9488 (N_9488,N_8670,N_8443);
nor U9489 (N_9489,N_8667,N_8924);
xnor U9490 (N_9490,N_8570,N_8859);
or U9491 (N_9491,N_8935,N_8690);
nor U9492 (N_9492,N_8491,N_8801);
nor U9493 (N_9493,N_8825,N_8856);
and U9494 (N_9494,N_8983,N_8660);
nand U9495 (N_9495,N_8425,N_8790);
and U9496 (N_9496,N_8444,N_8916);
nor U9497 (N_9497,N_8783,N_8819);
and U9498 (N_9498,N_8560,N_8959);
xnor U9499 (N_9499,N_8494,N_8787);
or U9500 (N_9500,N_8466,N_8540);
xor U9501 (N_9501,N_8413,N_8809);
or U9502 (N_9502,N_8591,N_8824);
nand U9503 (N_9503,N_8779,N_8518);
or U9504 (N_9504,N_8808,N_8620);
and U9505 (N_9505,N_8552,N_8428);
or U9506 (N_9506,N_8659,N_8815);
and U9507 (N_9507,N_8693,N_8846);
nor U9508 (N_9508,N_8519,N_8881);
xnor U9509 (N_9509,N_8886,N_8640);
or U9510 (N_9510,N_8827,N_8546);
nor U9511 (N_9511,N_8813,N_8566);
or U9512 (N_9512,N_8993,N_8545);
or U9513 (N_9513,N_8857,N_8958);
or U9514 (N_9514,N_8865,N_8735);
nand U9515 (N_9515,N_8483,N_8688);
nor U9516 (N_9516,N_8731,N_8527);
and U9517 (N_9517,N_8766,N_8904);
or U9518 (N_9518,N_8771,N_8504);
or U9519 (N_9519,N_8801,N_8634);
nand U9520 (N_9520,N_8668,N_8545);
nor U9521 (N_9521,N_8419,N_8515);
nand U9522 (N_9522,N_8986,N_8997);
xor U9523 (N_9523,N_8903,N_8896);
xnor U9524 (N_9524,N_8566,N_8907);
nand U9525 (N_9525,N_8543,N_8754);
or U9526 (N_9526,N_8738,N_8805);
and U9527 (N_9527,N_8571,N_8623);
or U9528 (N_9528,N_8795,N_8404);
and U9529 (N_9529,N_8508,N_8580);
xnor U9530 (N_9530,N_8557,N_8882);
nor U9531 (N_9531,N_8728,N_8821);
xnor U9532 (N_9532,N_8993,N_8637);
and U9533 (N_9533,N_8564,N_8523);
and U9534 (N_9534,N_8610,N_8935);
xor U9535 (N_9535,N_8675,N_8846);
nor U9536 (N_9536,N_8768,N_8505);
nor U9537 (N_9537,N_8829,N_8730);
nor U9538 (N_9538,N_8449,N_8534);
or U9539 (N_9539,N_8947,N_8488);
nand U9540 (N_9540,N_8737,N_8560);
and U9541 (N_9541,N_8783,N_8926);
nor U9542 (N_9542,N_8627,N_8573);
and U9543 (N_9543,N_8677,N_8955);
or U9544 (N_9544,N_8602,N_8692);
or U9545 (N_9545,N_8989,N_8969);
xnor U9546 (N_9546,N_8644,N_8427);
xnor U9547 (N_9547,N_8809,N_8872);
or U9548 (N_9548,N_8468,N_8964);
nor U9549 (N_9549,N_8595,N_8604);
and U9550 (N_9550,N_8649,N_8419);
nor U9551 (N_9551,N_8841,N_8624);
or U9552 (N_9552,N_8656,N_8991);
nor U9553 (N_9553,N_8459,N_8555);
xnor U9554 (N_9554,N_8592,N_8759);
nor U9555 (N_9555,N_8418,N_8591);
or U9556 (N_9556,N_8677,N_8512);
or U9557 (N_9557,N_8662,N_8865);
and U9558 (N_9558,N_8513,N_8711);
or U9559 (N_9559,N_8941,N_8818);
nor U9560 (N_9560,N_8862,N_8696);
xnor U9561 (N_9561,N_8410,N_8983);
nor U9562 (N_9562,N_8723,N_8777);
xor U9563 (N_9563,N_8488,N_8857);
and U9564 (N_9564,N_8562,N_8624);
nor U9565 (N_9565,N_8770,N_8640);
nand U9566 (N_9566,N_8698,N_8995);
and U9567 (N_9567,N_8527,N_8583);
nor U9568 (N_9568,N_8770,N_8537);
nand U9569 (N_9569,N_8828,N_8876);
and U9570 (N_9570,N_8768,N_8446);
xnor U9571 (N_9571,N_8607,N_8405);
xnor U9572 (N_9572,N_8800,N_8655);
nand U9573 (N_9573,N_8648,N_8893);
nand U9574 (N_9574,N_8802,N_8778);
nand U9575 (N_9575,N_8592,N_8715);
nand U9576 (N_9576,N_8670,N_8750);
and U9577 (N_9577,N_8916,N_8682);
nand U9578 (N_9578,N_8879,N_8782);
nand U9579 (N_9579,N_8910,N_8985);
nor U9580 (N_9580,N_8903,N_8640);
xor U9581 (N_9581,N_8504,N_8474);
xnor U9582 (N_9582,N_8655,N_8584);
nand U9583 (N_9583,N_8480,N_8989);
xor U9584 (N_9584,N_8538,N_8650);
nor U9585 (N_9585,N_8543,N_8799);
xor U9586 (N_9586,N_8880,N_8533);
nor U9587 (N_9587,N_8662,N_8467);
xnor U9588 (N_9588,N_8931,N_8743);
xor U9589 (N_9589,N_8726,N_8449);
nor U9590 (N_9590,N_8428,N_8609);
xnor U9591 (N_9591,N_8692,N_8606);
and U9592 (N_9592,N_8621,N_8640);
nand U9593 (N_9593,N_8827,N_8886);
nor U9594 (N_9594,N_8453,N_8611);
xor U9595 (N_9595,N_8708,N_8731);
nor U9596 (N_9596,N_8515,N_8508);
nor U9597 (N_9597,N_8710,N_8794);
and U9598 (N_9598,N_8602,N_8986);
nand U9599 (N_9599,N_8966,N_8417);
nor U9600 (N_9600,N_9460,N_9534);
nor U9601 (N_9601,N_9312,N_9155);
or U9602 (N_9602,N_9220,N_9005);
xnor U9603 (N_9603,N_9316,N_9486);
and U9604 (N_9604,N_9524,N_9371);
xor U9605 (N_9605,N_9161,N_9348);
xor U9606 (N_9606,N_9477,N_9326);
nor U9607 (N_9607,N_9124,N_9301);
nor U9608 (N_9608,N_9347,N_9239);
nor U9609 (N_9609,N_9284,N_9015);
xor U9610 (N_9610,N_9075,N_9370);
and U9611 (N_9611,N_9364,N_9232);
nor U9612 (N_9612,N_9212,N_9331);
xor U9613 (N_9613,N_9508,N_9247);
and U9614 (N_9614,N_9057,N_9048);
or U9615 (N_9615,N_9596,N_9406);
and U9616 (N_9616,N_9039,N_9554);
nor U9617 (N_9617,N_9384,N_9575);
nand U9618 (N_9618,N_9393,N_9139);
nor U9619 (N_9619,N_9398,N_9181);
and U9620 (N_9620,N_9550,N_9471);
and U9621 (N_9621,N_9569,N_9073);
nand U9622 (N_9622,N_9016,N_9046);
or U9623 (N_9623,N_9437,N_9149);
nor U9624 (N_9624,N_9590,N_9008);
nand U9625 (N_9625,N_9093,N_9339);
nor U9626 (N_9626,N_9188,N_9307);
xnor U9627 (N_9627,N_9333,N_9510);
nor U9628 (N_9628,N_9147,N_9434);
or U9629 (N_9629,N_9376,N_9017);
nor U9630 (N_9630,N_9221,N_9055);
or U9631 (N_9631,N_9352,N_9226);
nor U9632 (N_9632,N_9213,N_9243);
nand U9633 (N_9633,N_9513,N_9063);
and U9634 (N_9634,N_9553,N_9447);
and U9635 (N_9635,N_9336,N_9077);
xor U9636 (N_9636,N_9323,N_9234);
nor U9637 (N_9637,N_9196,N_9351);
xnor U9638 (N_9638,N_9580,N_9094);
and U9639 (N_9639,N_9570,N_9224);
nor U9640 (N_9640,N_9388,N_9480);
nor U9641 (N_9641,N_9318,N_9303);
or U9642 (N_9642,N_9292,N_9296);
xnor U9643 (N_9643,N_9254,N_9202);
nand U9644 (N_9644,N_9571,N_9069);
xor U9645 (N_9645,N_9379,N_9459);
nand U9646 (N_9646,N_9125,N_9193);
xnor U9647 (N_9647,N_9419,N_9417);
and U9648 (N_9648,N_9389,N_9546);
xnor U9649 (N_9649,N_9442,N_9011);
and U9650 (N_9650,N_9478,N_9558);
or U9651 (N_9651,N_9573,N_9006);
and U9652 (N_9652,N_9222,N_9429);
or U9653 (N_9653,N_9367,N_9433);
nor U9654 (N_9654,N_9516,N_9404);
nor U9655 (N_9655,N_9241,N_9283);
or U9656 (N_9656,N_9564,N_9185);
nor U9657 (N_9657,N_9047,N_9171);
or U9658 (N_9658,N_9211,N_9131);
or U9659 (N_9659,N_9054,N_9096);
and U9660 (N_9660,N_9383,N_9200);
nor U9661 (N_9661,N_9018,N_9444);
and U9662 (N_9662,N_9128,N_9523);
nor U9663 (N_9663,N_9502,N_9158);
nor U9664 (N_9664,N_9293,N_9214);
and U9665 (N_9665,N_9026,N_9002);
or U9666 (N_9666,N_9207,N_9204);
nand U9667 (N_9667,N_9427,N_9540);
or U9668 (N_9668,N_9410,N_9541);
nand U9669 (N_9669,N_9304,N_9042);
nor U9670 (N_9670,N_9458,N_9085);
nand U9671 (N_9671,N_9407,N_9566);
nor U9672 (N_9672,N_9431,N_9137);
or U9673 (N_9673,N_9386,N_9079);
xnor U9674 (N_9674,N_9595,N_9394);
nand U9675 (N_9675,N_9010,N_9556);
nand U9676 (N_9676,N_9416,N_9350);
and U9677 (N_9677,N_9536,N_9468);
and U9678 (N_9678,N_9559,N_9080);
or U9679 (N_9679,N_9259,N_9387);
xnor U9680 (N_9680,N_9062,N_9356);
xnor U9681 (N_9681,N_9560,N_9519);
xnor U9682 (N_9682,N_9110,N_9365);
nand U9683 (N_9683,N_9172,N_9027);
xnor U9684 (N_9684,N_9157,N_9402);
nand U9685 (N_9685,N_9390,N_9432);
nor U9686 (N_9686,N_9142,N_9512);
nor U9687 (N_9687,N_9266,N_9197);
and U9688 (N_9688,N_9330,N_9428);
nor U9689 (N_9689,N_9176,N_9021);
nor U9690 (N_9690,N_9036,N_9170);
nand U9691 (N_9691,N_9260,N_9229);
and U9692 (N_9692,N_9332,N_9092);
and U9693 (N_9693,N_9245,N_9578);
nor U9694 (N_9694,N_9114,N_9533);
or U9695 (N_9695,N_9454,N_9599);
nor U9696 (N_9696,N_9579,N_9014);
nor U9697 (N_9697,N_9572,N_9525);
nand U9698 (N_9698,N_9342,N_9515);
nand U9699 (N_9699,N_9413,N_9242);
nand U9700 (N_9700,N_9050,N_9089);
or U9701 (N_9701,N_9289,N_9252);
nand U9702 (N_9702,N_9520,N_9194);
xnor U9703 (N_9703,N_9225,N_9377);
or U9704 (N_9704,N_9076,N_9236);
nor U9705 (N_9705,N_9363,N_9127);
or U9706 (N_9706,N_9380,N_9274);
nor U9707 (N_9707,N_9581,N_9217);
nor U9708 (N_9708,N_9315,N_9163);
xor U9709 (N_9709,N_9280,N_9216);
nand U9710 (N_9710,N_9425,N_9111);
and U9711 (N_9711,N_9396,N_9150);
xnor U9712 (N_9712,N_9215,N_9522);
nor U9713 (N_9713,N_9038,N_9058);
nand U9714 (N_9714,N_9494,N_9001);
and U9715 (N_9715,N_9208,N_9133);
nand U9716 (N_9716,N_9244,N_9409);
nand U9717 (N_9717,N_9251,N_9209);
xnor U9718 (N_9718,N_9308,N_9070);
nand U9719 (N_9719,N_9141,N_9190);
and U9720 (N_9720,N_9030,N_9210);
xnor U9721 (N_9721,N_9526,N_9025);
or U9722 (N_9722,N_9311,N_9445);
or U9723 (N_9723,N_9143,N_9594);
and U9724 (N_9724,N_9426,N_9148);
nand U9725 (N_9725,N_9116,N_9343);
or U9726 (N_9726,N_9009,N_9360);
or U9727 (N_9727,N_9294,N_9305);
nor U9728 (N_9728,N_9175,N_9324);
or U9729 (N_9729,N_9506,N_9322);
and U9730 (N_9730,N_9366,N_9435);
nor U9731 (N_9731,N_9189,N_9498);
xor U9732 (N_9732,N_9145,N_9473);
xnor U9733 (N_9733,N_9557,N_9320);
nand U9734 (N_9734,N_9112,N_9481);
and U9735 (N_9735,N_9562,N_9123);
xor U9736 (N_9736,N_9532,N_9321);
xor U9737 (N_9737,N_9195,N_9357);
and U9738 (N_9738,N_9151,N_9577);
nor U9739 (N_9739,N_9449,N_9338);
or U9740 (N_9740,N_9275,N_9415);
xor U9741 (N_9741,N_9485,N_9452);
or U9742 (N_9742,N_9592,N_9253);
nand U9743 (N_9743,N_9088,N_9490);
nor U9744 (N_9744,N_9263,N_9180);
nand U9745 (N_9745,N_9474,N_9037);
or U9746 (N_9746,N_9401,N_9574);
nor U9747 (N_9747,N_9053,N_9103);
xnor U9748 (N_9748,N_9507,N_9593);
or U9749 (N_9749,N_9531,N_9511);
or U9750 (N_9750,N_9529,N_9344);
nand U9751 (N_9751,N_9166,N_9064);
and U9752 (N_9752,N_9203,N_9081);
xnor U9753 (N_9753,N_9505,N_9464);
xnor U9754 (N_9754,N_9403,N_9132);
nor U9755 (N_9755,N_9378,N_9543);
xor U9756 (N_9756,N_9013,N_9306);
and U9757 (N_9757,N_9493,N_9418);
nor U9758 (N_9758,N_9405,N_9456);
nor U9759 (N_9759,N_9597,N_9091);
nand U9760 (N_9760,N_9567,N_9290);
nor U9761 (N_9761,N_9327,N_9061);
xor U9762 (N_9762,N_9340,N_9022);
xor U9763 (N_9763,N_9530,N_9273);
nor U9764 (N_9764,N_9095,N_9272);
nor U9765 (N_9765,N_9514,N_9361);
xor U9766 (N_9766,N_9129,N_9153);
xor U9767 (N_9767,N_9049,N_9487);
or U9768 (N_9768,N_9463,N_9362);
nand U9769 (N_9769,N_9443,N_9119);
or U9770 (N_9770,N_9467,N_9205);
xor U9771 (N_9771,N_9334,N_9246);
nor U9772 (N_9772,N_9173,N_9035);
and U9773 (N_9773,N_9358,N_9504);
and U9774 (N_9774,N_9023,N_9184);
nand U9775 (N_9775,N_9261,N_9489);
and U9776 (N_9776,N_9101,N_9302);
nor U9777 (N_9777,N_9551,N_9067);
nor U9778 (N_9778,N_9300,N_9255);
and U9779 (N_9779,N_9517,N_9500);
nor U9780 (N_9780,N_9098,N_9281);
nand U9781 (N_9781,N_9156,N_9033);
and U9782 (N_9782,N_9084,N_9482);
or U9783 (N_9783,N_9430,N_9000);
or U9784 (N_9784,N_9100,N_9159);
nand U9785 (N_9785,N_9382,N_9450);
or U9786 (N_9786,N_9107,N_9040);
nor U9787 (N_9787,N_9421,N_9183);
or U9788 (N_9788,N_9448,N_9012);
or U9789 (N_9789,N_9154,N_9328);
nand U9790 (N_9790,N_9034,N_9568);
nand U9791 (N_9791,N_9056,N_9105);
xor U9792 (N_9792,N_9346,N_9024);
nand U9793 (N_9793,N_9231,N_9545);
xnor U9794 (N_9794,N_9375,N_9438);
nor U9795 (N_9795,N_9257,N_9068);
nand U9796 (N_9796,N_9121,N_9270);
nand U9797 (N_9797,N_9065,N_9399);
xor U9798 (N_9798,N_9267,N_9457);
and U9799 (N_9799,N_9249,N_9535);
or U9800 (N_9800,N_9537,N_9099);
or U9801 (N_9801,N_9019,N_9223);
xor U9802 (N_9802,N_9341,N_9262);
or U9803 (N_9803,N_9074,N_9583);
or U9804 (N_9804,N_9174,N_9495);
xor U9805 (N_9805,N_9233,N_9130);
nand U9806 (N_9806,N_9598,N_9455);
nand U9807 (N_9807,N_9059,N_9527);
and U9808 (N_9808,N_9186,N_9288);
nor U9809 (N_9809,N_9397,N_9104);
and U9810 (N_9810,N_9400,N_9256);
xor U9811 (N_9811,N_9408,N_9167);
and U9812 (N_9812,N_9368,N_9240);
nor U9813 (N_9813,N_9521,N_9492);
and U9814 (N_9814,N_9317,N_9491);
or U9815 (N_9815,N_9271,N_9276);
xnor U9816 (N_9816,N_9483,N_9538);
or U9817 (N_9817,N_9299,N_9469);
or U9818 (N_9818,N_9325,N_9446);
and U9819 (N_9819,N_9286,N_9138);
xor U9820 (N_9820,N_9354,N_9282);
nor U9821 (N_9821,N_9392,N_9497);
and U9822 (N_9822,N_9582,N_9087);
or U9823 (N_9823,N_9265,N_9160);
nor U9824 (N_9824,N_9206,N_9359);
nand U9825 (N_9825,N_9178,N_9250);
xnor U9826 (N_9826,N_9140,N_9279);
or U9827 (N_9827,N_9120,N_9144);
nor U9828 (N_9828,N_9182,N_9539);
xor U9829 (N_9829,N_9462,N_9470);
xor U9830 (N_9830,N_9310,N_9043);
nor U9831 (N_9831,N_9227,N_9349);
or U9832 (N_9832,N_9484,N_9051);
nand U9833 (N_9833,N_9385,N_9264);
and U9834 (N_9834,N_9028,N_9277);
nor U9835 (N_9835,N_9238,N_9235);
nor U9836 (N_9836,N_9373,N_9004);
and U9837 (N_9837,N_9335,N_9177);
or U9838 (N_9838,N_9549,N_9258);
xor U9839 (N_9839,N_9411,N_9298);
nor U9840 (N_9840,N_9218,N_9576);
or U9841 (N_9841,N_9441,N_9309);
nor U9842 (N_9842,N_9285,N_9071);
nor U9843 (N_9843,N_9122,N_9108);
nand U9844 (N_9844,N_9007,N_9548);
and U9845 (N_9845,N_9314,N_9381);
or U9846 (N_9846,N_9372,N_9423);
xor U9847 (N_9847,N_9501,N_9453);
and U9848 (N_9848,N_9106,N_9329);
xor U9849 (N_9849,N_9586,N_9134);
nand U9850 (N_9850,N_9422,N_9563);
and U9851 (N_9851,N_9589,N_9496);
and U9852 (N_9852,N_9374,N_9109);
or U9853 (N_9853,N_9518,N_9391);
and U9854 (N_9854,N_9345,N_9192);
and U9855 (N_9855,N_9117,N_9083);
nand U9856 (N_9856,N_9461,N_9420);
nand U9857 (N_9857,N_9113,N_9169);
nand U9858 (N_9858,N_9542,N_9297);
nor U9859 (N_9859,N_9509,N_9097);
nand U9860 (N_9860,N_9369,N_9488);
nand U9861 (N_9861,N_9066,N_9465);
nand U9862 (N_9862,N_9278,N_9191);
xnor U9863 (N_9863,N_9565,N_9136);
nand U9864 (N_9864,N_9135,N_9146);
and U9865 (N_9865,N_9078,N_9499);
xnor U9866 (N_9866,N_9319,N_9591);
and U9867 (N_9867,N_9198,N_9060);
and U9868 (N_9868,N_9269,N_9475);
or U9869 (N_9869,N_9451,N_9126);
nand U9870 (N_9870,N_9152,N_9228);
or U9871 (N_9871,N_9031,N_9395);
xnor U9872 (N_9872,N_9584,N_9295);
and U9873 (N_9873,N_9086,N_9199);
or U9874 (N_9874,N_9187,N_9472);
and U9875 (N_9875,N_9291,N_9164);
or U9876 (N_9876,N_9412,N_9237);
nand U9877 (N_9877,N_9072,N_9424);
or U9878 (N_9878,N_9479,N_9547);
or U9879 (N_9879,N_9503,N_9248);
xnor U9880 (N_9880,N_9439,N_9003);
nand U9881 (N_9881,N_9476,N_9561);
xor U9882 (N_9882,N_9165,N_9020);
xor U9883 (N_9883,N_9588,N_9044);
and U9884 (N_9884,N_9587,N_9440);
and U9885 (N_9885,N_9337,N_9082);
and U9886 (N_9886,N_9045,N_9168);
nand U9887 (N_9887,N_9585,N_9115);
and U9888 (N_9888,N_9029,N_9179);
xor U9889 (N_9889,N_9219,N_9555);
or U9890 (N_9890,N_9090,N_9052);
or U9891 (N_9891,N_9544,N_9102);
xor U9892 (N_9892,N_9268,N_9552);
nor U9893 (N_9893,N_9201,N_9032);
nand U9894 (N_9894,N_9041,N_9230);
nand U9895 (N_9895,N_9287,N_9414);
nor U9896 (N_9896,N_9528,N_9162);
and U9897 (N_9897,N_9118,N_9466);
nand U9898 (N_9898,N_9313,N_9355);
nand U9899 (N_9899,N_9353,N_9436);
or U9900 (N_9900,N_9059,N_9123);
xor U9901 (N_9901,N_9441,N_9053);
and U9902 (N_9902,N_9306,N_9397);
nor U9903 (N_9903,N_9562,N_9552);
nor U9904 (N_9904,N_9542,N_9447);
nor U9905 (N_9905,N_9066,N_9421);
nand U9906 (N_9906,N_9452,N_9253);
and U9907 (N_9907,N_9107,N_9003);
or U9908 (N_9908,N_9329,N_9523);
or U9909 (N_9909,N_9572,N_9170);
or U9910 (N_9910,N_9194,N_9364);
and U9911 (N_9911,N_9558,N_9472);
and U9912 (N_9912,N_9377,N_9011);
nor U9913 (N_9913,N_9539,N_9353);
or U9914 (N_9914,N_9164,N_9144);
xnor U9915 (N_9915,N_9563,N_9032);
xnor U9916 (N_9916,N_9463,N_9037);
xor U9917 (N_9917,N_9313,N_9437);
and U9918 (N_9918,N_9336,N_9166);
or U9919 (N_9919,N_9306,N_9373);
or U9920 (N_9920,N_9554,N_9456);
and U9921 (N_9921,N_9124,N_9357);
and U9922 (N_9922,N_9330,N_9183);
nand U9923 (N_9923,N_9008,N_9282);
nand U9924 (N_9924,N_9143,N_9278);
xnor U9925 (N_9925,N_9283,N_9538);
xnor U9926 (N_9926,N_9324,N_9403);
nand U9927 (N_9927,N_9039,N_9279);
and U9928 (N_9928,N_9111,N_9534);
nor U9929 (N_9929,N_9323,N_9198);
or U9930 (N_9930,N_9363,N_9262);
xor U9931 (N_9931,N_9531,N_9452);
or U9932 (N_9932,N_9051,N_9431);
nor U9933 (N_9933,N_9595,N_9500);
or U9934 (N_9934,N_9250,N_9211);
nor U9935 (N_9935,N_9560,N_9255);
nand U9936 (N_9936,N_9222,N_9113);
xnor U9937 (N_9937,N_9239,N_9379);
nand U9938 (N_9938,N_9196,N_9583);
or U9939 (N_9939,N_9318,N_9107);
nand U9940 (N_9940,N_9356,N_9304);
xor U9941 (N_9941,N_9374,N_9274);
xnor U9942 (N_9942,N_9162,N_9125);
nand U9943 (N_9943,N_9462,N_9256);
or U9944 (N_9944,N_9189,N_9507);
nor U9945 (N_9945,N_9581,N_9161);
nor U9946 (N_9946,N_9042,N_9511);
nand U9947 (N_9947,N_9058,N_9391);
nand U9948 (N_9948,N_9480,N_9393);
or U9949 (N_9949,N_9474,N_9251);
nand U9950 (N_9950,N_9290,N_9376);
nand U9951 (N_9951,N_9190,N_9336);
nand U9952 (N_9952,N_9147,N_9233);
xor U9953 (N_9953,N_9075,N_9565);
nand U9954 (N_9954,N_9159,N_9460);
and U9955 (N_9955,N_9060,N_9254);
nand U9956 (N_9956,N_9540,N_9203);
nand U9957 (N_9957,N_9109,N_9177);
nor U9958 (N_9958,N_9439,N_9422);
nor U9959 (N_9959,N_9117,N_9549);
nor U9960 (N_9960,N_9330,N_9253);
or U9961 (N_9961,N_9548,N_9439);
nor U9962 (N_9962,N_9521,N_9174);
nor U9963 (N_9963,N_9101,N_9033);
nor U9964 (N_9964,N_9057,N_9064);
or U9965 (N_9965,N_9591,N_9367);
nand U9966 (N_9966,N_9340,N_9173);
nand U9967 (N_9967,N_9232,N_9060);
nor U9968 (N_9968,N_9037,N_9009);
nor U9969 (N_9969,N_9375,N_9403);
and U9970 (N_9970,N_9318,N_9124);
or U9971 (N_9971,N_9451,N_9147);
nor U9972 (N_9972,N_9572,N_9281);
xnor U9973 (N_9973,N_9158,N_9086);
nor U9974 (N_9974,N_9130,N_9046);
and U9975 (N_9975,N_9061,N_9459);
nor U9976 (N_9976,N_9252,N_9592);
and U9977 (N_9977,N_9055,N_9558);
or U9978 (N_9978,N_9589,N_9253);
and U9979 (N_9979,N_9461,N_9090);
xor U9980 (N_9980,N_9433,N_9530);
and U9981 (N_9981,N_9590,N_9226);
or U9982 (N_9982,N_9532,N_9529);
nor U9983 (N_9983,N_9210,N_9173);
xor U9984 (N_9984,N_9536,N_9247);
or U9985 (N_9985,N_9397,N_9355);
or U9986 (N_9986,N_9304,N_9270);
and U9987 (N_9987,N_9393,N_9175);
nand U9988 (N_9988,N_9353,N_9355);
nand U9989 (N_9989,N_9491,N_9199);
xnor U9990 (N_9990,N_9535,N_9267);
xnor U9991 (N_9991,N_9599,N_9054);
xnor U9992 (N_9992,N_9065,N_9125);
and U9993 (N_9993,N_9583,N_9187);
and U9994 (N_9994,N_9475,N_9083);
and U9995 (N_9995,N_9440,N_9023);
xor U9996 (N_9996,N_9392,N_9156);
and U9997 (N_9997,N_9223,N_9430);
and U9998 (N_9998,N_9194,N_9347);
or U9999 (N_9999,N_9312,N_9412);
or U10000 (N_10000,N_9197,N_9274);
nand U10001 (N_10001,N_9589,N_9407);
and U10002 (N_10002,N_9041,N_9286);
nand U10003 (N_10003,N_9170,N_9319);
xor U10004 (N_10004,N_9010,N_9322);
or U10005 (N_10005,N_9321,N_9513);
or U10006 (N_10006,N_9108,N_9562);
and U10007 (N_10007,N_9457,N_9046);
xor U10008 (N_10008,N_9166,N_9357);
and U10009 (N_10009,N_9537,N_9398);
nand U10010 (N_10010,N_9098,N_9113);
nand U10011 (N_10011,N_9419,N_9312);
and U10012 (N_10012,N_9107,N_9192);
xnor U10013 (N_10013,N_9286,N_9441);
or U10014 (N_10014,N_9205,N_9030);
nand U10015 (N_10015,N_9324,N_9541);
or U10016 (N_10016,N_9500,N_9116);
xor U10017 (N_10017,N_9527,N_9407);
nand U10018 (N_10018,N_9202,N_9286);
and U10019 (N_10019,N_9412,N_9277);
nand U10020 (N_10020,N_9082,N_9495);
nor U10021 (N_10021,N_9380,N_9188);
nand U10022 (N_10022,N_9554,N_9286);
or U10023 (N_10023,N_9049,N_9424);
xnor U10024 (N_10024,N_9434,N_9168);
and U10025 (N_10025,N_9098,N_9118);
xor U10026 (N_10026,N_9438,N_9145);
xor U10027 (N_10027,N_9433,N_9554);
and U10028 (N_10028,N_9045,N_9232);
nand U10029 (N_10029,N_9094,N_9534);
or U10030 (N_10030,N_9176,N_9333);
nand U10031 (N_10031,N_9478,N_9396);
and U10032 (N_10032,N_9353,N_9260);
nand U10033 (N_10033,N_9444,N_9236);
and U10034 (N_10034,N_9416,N_9289);
nor U10035 (N_10035,N_9305,N_9435);
nor U10036 (N_10036,N_9128,N_9036);
nor U10037 (N_10037,N_9588,N_9308);
or U10038 (N_10038,N_9072,N_9431);
or U10039 (N_10039,N_9259,N_9325);
nand U10040 (N_10040,N_9249,N_9394);
nor U10041 (N_10041,N_9590,N_9139);
or U10042 (N_10042,N_9551,N_9384);
nor U10043 (N_10043,N_9370,N_9095);
nand U10044 (N_10044,N_9567,N_9139);
nor U10045 (N_10045,N_9187,N_9382);
xor U10046 (N_10046,N_9384,N_9300);
and U10047 (N_10047,N_9053,N_9197);
or U10048 (N_10048,N_9084,N_9357);
and U10049 (N_10049,N_9341,N_9585);
nand U10050 (N_10050,N_9307,N_9393);
xor U10051 (N_10051,N_9223,N_9129);
nand U10052 (N_10052,N_9128,N_9486);
xor U10053 (N_10053,N_9572,N_9117);
nor U10054 (N_10054,N_9088,N_9169);
xnor U10055 (N_10055,N_9097,N_9385);
nor U10056 (N_10056,N_9208,N_9123);
xor U10057 (N_10057,N_9056,N_9106);
or U10058 (N_10058,N_9512,N_9120);
nor U10059 (N_10059,N_9224,N_9409);
or U10060 (N_10060,N_9542,N_9327);
xor U10061 (N_10061,N_9032,N_9188);
nand U10062 (N_10062,N_9441,N_9166);
and U10063 (N_10063,N_9076,N_9096);
or U10064 (N_10064,N_9213,N_9520);
xnor U10065 (N_10065,N_9025,N_9102);
xor U10066 (N_10066,N_9021,N_9093);
or U10067 (N_10067,N_9410,N_9279);
or U10068 (N_10068,N_9246,N_9400);
and U10069 (N_10069,N_9461,N_9488);
and U10070 (N_10070,N_9577,N_9186);
xor U10071 (N_10071,N_9410,N_9519);
or U10072 (N_10072,N_9328,N_9399);
and U10073 (N_10073,N_9406,N_9324);
and U10074 (N_10074,N_9550,N_9106);
and U10075 (N_10075,N_9189,N_9559);
nand U10076 (N_10076,N_9302,N_9342);
nor U10077 (N_10077,N_9429,N_9388);
nor U10078 (N_10078,N_9275,N_9372);
and U10079 (N_10079,N_9008,N_9192);
xor U10080 (N_10080,N_9076,N_9050);
or U10081 (N_10081,N_9418,N_9143);
xor U10082 (N_10082,N_9176,N_9520);
or U10083 (N_10083,N_9379,N_9345);
nand U10084 (N_10084,N_9239,N_9290);
nand U10085 (N_10085,N_9327,N_9507);
and U10086 (N_10086,N_9249,N_9369);
nor U10087 (N_10087,N_9565,N_9021);
nor U10088 (N_10088,N_9235,N_9250);
and U10089 (N_10089,N_9024,N_9113);
and U10090 (N_10090,N_9364,N_9184);
and U10091 (N_10091,N_9302,N_9241);
and U10092 (N_10092,N_9363,N_9459);
or U10093 (N_10093,N_9024,N_9198);
and U10094 (N_10094,N_9213,N_9041);
or U10095 (N_10095,N_9457,N_9569);
nand U10096 (N_10096,N_9148,N_9191);
or U10097 (N_10097,N_9283,N_9197);
and U10098 (N_10098,N_9490,N_9000);
nand U10099 (N_10099,N_9016,N_9569);
or U10100 (N_10100,N_9463,N_9192);
or U10101 (N_10101,N_9296,N_9065);
and U10102 (N_10102,N_9342,N_9100);
or U10103 (N_10103,N_9229,N_9397);
or U10104 (N_10104,N_9483,N_9513);
nor U10105 (N_10105,N_9564,N_9485);
and U10106 (N_10106,N_9566,N_9029);
nand U10107 (N_10107,N_9421,N_9487);
or U10108 (N_10108,N_9205,N_9028);
nor U10109 (N_10109,N_9146,N_9157);
xnor U10110 (N_10110,N_9171,N_9449);
xor U10111 (N_10111,N_9087,N_9299);
nand U10112 (N_10112,N_9513,N_9564);
xor U10113 (N_10113,N_9331,N_9166);
and U10114 (N_10114,N_9493,N_9468);
xor U10115 (N_10115,N_9377,N_9413);
nor U10116 (N_10116,N_9018,N_9283);
nand U10117 (N_10117,N_9423,N_9518);
nand U10118 (N_10118,N_9316,N_9348);
nand U10119 (N_10119,N_9370,N_9226);
or U10120 (N_10120,N_9123,N_9287);
nand U10121 (N_10121,N_9383,N_9190);
or U10122 (N_10122,N_9247,N_9370);
or U10123 (N_10123,N_9122,N_9562);
or U10124 (N_10124,N_9497,N_9034);
nand U10125 (N_10125,N_9183,N_9283);
nand U10126 (N_10126,N_9167,N_9549);
nor U10127 (N_10127,N_9283,N_9501);
xor U10128 (N_10128,N_9570,N_9459);
nor U10129 (N_10129,N_9491,N_9450);
xnor U10130 (N_10130,N_9170,N_9075);
nand U10131 (N_10131,N_9397,N_9111);
nor U10132 (N_10132,N_9200,N_9585);
xnor U10133 (N_10133,N_9227,N_9044);
and U10134 (N_10134,N_9399,N_9565);
and U10135 (N_10135,N_9018,N_9316);
nand U10136 (N_10136,N_9313,N_9021);
nor U10137 (N_10137,N_9533,N_9031);
nand U10138 (N_10138,N_9517,N_9199);
or U10139 (N_10139,N_9109,N_9087);
or U10140 (N_10140,N_9219,N_9256);
or U10141 (N_10141,N_9277,N_9392);
and U10142 (N_10142,N_9427,N_9163);
xnor U10143 (N_10143,N_9238,N_9417);
and U10144 (N_10144,N_9485,N_9042);
nor U10145 (N_10145,N_9006,N_9173);
or U10146 (N_10146,N_9513,N_9091);
and U10147 (N_10147,N_9335,N_9383);
nand U10148 (N_10148,N_9589,N_9392);
xnor U10149 (N_10149,N_9317,N_9231);
xor U10150 (N_10150,N_9507,N_9396);
or U10151 (N_10151,N_9208,N_9212);
and U10152 (N_10152,N_9473,N_9048);
or U10153 (N_10153,N_9302,N_9435);
and U10154 (N_10154,N_9150,N_9446);
xor U10155 (N_10155,N_9083,N_9397);
and U10156 (N_10156,N_9395,N_9445);
nor U10157 (N_10157,N_9358,N_9006);
nor U10158 (N_10158,N_9250,N_9076);
and U10159 (N_10159,N_9238,N_9427);
and U10160 (N_10160,N_9453,N_9353);
or U10161 (N_10161,N_9402,N_9015);
and U10162 (N_10162,N_9134,N_9282);
nand U10163 (N_10163,N_9081,N_9064);
xnor U10164 (N_10164,N_9471,N_9245);
or U10165 (N_10165,N_9408,N_9015);
or U10166 (N_10166,N_9017,N_9460);
or U10167 (N_10167,N_9405,N_9003);
nor U10168 (N_10168,N_9592,N_9594);
or U10169 (N_10169,N_9098,N_9535);
nand U10170 (N_10170,N_9435,N_9029);
nor U10171 (N_10171,N_9570,N_9028);
nand U10172 (N_10172,N_9511,N_9134);
nand U10173 (N_10173,N_9485,N_9291);
nor U10174 (N_10174,N_9414,N_9207);
and U10175 (N_10175,N_9533,N_9254);
or U10176 (N_10176,N_9229,N_9287);
or U10177 (N_10177,N_9553,N_9127);
nand U10178 (N_10178,N_9378,N_9593);
nor U10179 (N_10179,N_9208,N_9458);
xnor U10180 (N_10180,N_9034,N_9060);
nand U10181 (N_10181,N_9573,N_9069);
nand U10182 (N_10182,N_9239,N_9163);
nor U10183 (N_10183,N_9311,N_9226);
and U10184 (N_10184,N_9325,N_9027);
nor U10185 (N_10185,N_9120,N_9255);
xor U10186 (N_10186,N_9365,N_9310);
or U10187 (N_10187,N_9464,N_9530);
or U10188 (N_10188,N_9144,N_9208);
xor U10189 (N_10189,N_9374,N_9549);
nand U10190 (N_10190,N_9400,N_9512);
nand U10191 (N_10191,N_9256,N_9084);
or U10192 (N_10192,N_9154,N_9511);
nand U10193 (N_10193,N_9525,N_9090);
nand U10194 (N_10194,N_9527,N_9348);
nand U10195 (N_10195,N_9229,N_9275);
xor U10196 (N_10196,N_9028,N_9599);
nand U10197 (N_10197,N_9267,N_9408);
nand U10198 (N_10198,N_9105,N_9578);
and U10199 (N_10199,N_9376,N_9038);
nor U10200 (N_10200,N_10188,N_10146);
nand U10201 (N_10201,N_10079,N_9912);
or U10202 (N_10202,N_10141,N_9718);
or U10203 (N_10203,N_9725,N_9868);
or U10204 (N_10204,N_10170,N_9984);
nor U10205 (N_10205,N_10097,N_9849);
nor U10206 (N_10206,N_9885,N_9715);
and U10207 (N_10207,N_9829,N_9982);
or U10208 (N_10208,N_9993,N_9756);
nor U10209 (N_10209,N_9850,N_10154);
and U10210 (N_10210,N_9954,N_9866);
and U10211 (N_10211,N_10047,N_10031);
nor U10212 (N_10212,N_9925,N_10044);
and U10213 (N_10213,N_10169,N_10106);
or U10214 (N_10214,N_9729,N_9830);
nand U10215 (N_10215,N_9975,N_9844);
and U10216 (N_10216,N_9669,N_9940);
xor U10217 (N_10217,N_9709,N_9748);
and U10218 (N_10218,N_10160,N_9825);
xnor U10219 (N_10219,N_9661,N_9839);
nand U10220 (N_10220,N_9968,N_9969);
nor U10221 (N_10221,N_9600,N_9651);
xnor U10222 (N_10222,N_9989,N_10016);
and U10223 (N_10223,N_9689,N_9738);
and U10224 (N_10224,N_10005,N_10042);
nor U10225 (N_10225,N_9906,N_9821);
nor U10226 (N_10226,N_10165,N_9619);
or U10227 (N_10227,N_10043,N_9869);
xor U10228 (N_10228,N_10093,N_9743);
and U10229 (N_10229,N_9774,N_9882);
xnor U10230 (N_10230,N_10197,N_9811);
or U10231 (N_10231,N_9935,N_9727);
nand U10232 (N_10232,N_9790,N_10134);
nand U10233 (N_10233,N_9795,N_10184);
xor U10234 (N_10234,N_10173,N_9806);
nand U10235 (N_10235,N_10088,N_9653);
or U10236 (N_10236,N_9636,N_10126);
nand U10237 (N_10237,N_9688,N_9734);
and U10238 (N_10238,N_9919,N_9623);
nor U10239 (N_10239,N_9958,N_9762);
and U10240 (N_10240,N_9916,N_9941);
xnor U10241 (N_10241,N_9854,N_9780);
nor U10242 (N_10242,N_9652,N_9786);
or U10243 (N_10243,N_9787,N_9929);
xor U10244 (N_10244,N_9713,N_9741);
and U10245 (N_10245,N_9892,N_9603);
nor U10246 (N_10246,N_9633,N_9660);
or U10247 (N_10247,N_9957,N_10183);
nand U10248 (N_10248,N_9986,N_9634);
and U10249 (N_10249,N_10178,N_10102);
nand U10250 (N_10250,N_9802,N_9717);
or U10251 (N_10251,N_9883,N_10096);
and U10252 (N_10252,N_9755,N_9744);
or U10253 (N_10253,N_9629,N_9617);
or U10254 (N_10254,N_9827,N_9675);
or U10255 (N_10255,N_9997,N_9668);
or U10256 (N_10256,N_9648,N_10071);
and U10257 (N_10257,N_10123,N_10137);
nand U10258 (N_10258,N_10019,N_9698);
and U10259 (N_10259,N_10060,N_9974);
nand U10260 (N_10260,N_9872,N_10013);
nand U10261 (N_10261,N_10116,N_9608);
and U10262 (N_10262,N_9628,N_10176);
and U10263 (N_10263,N_9764,N_10131);
nor U10264 (N_10264,N_9807,N_9895);
and U10265 (N_10265,N_9938,N_9604);
xnor U10266 (N_10266,N_9972,N_9931);
and U10267 (N_10267,N_9799,N_9739);
xnor U10268 (N_10268,N_10034,N_10084);
and U10269 (N_10269,N_10006,N_10192);
or U10270 (N_10270,N_9772,N_9837);
nand U10271 (N_10271,N_9881,N_9967);
or U10272 (N_10272,N_9947,N_10129);
xor U10273 (N_10273,N_10189,N_9971);
xor U10274 (N_10274,N_10166,N_9991);
and U10275 (N_10275,N_9711,N_10077);
or U10276 (N_10276,N_10098,N_9845);
nand U10277 (N_10277,N_9720,N_10048);
nor U10278 (N_10278,N_9871,N_9961);
nand U10279 (N_10279,N_9949,N_9813);
or U10280 (N_10280,N_9656,N_9682);
or U10281 (N_10281,N_10151,N_10063);
xor U10282 (N_10282,N_9952,N_9988);
nand U10283 (N_10283,N_9831,N_9922);
xor U10284 (N_10284,N_9768,N_9693);
nand U10285 (N_10285,N_9887,N_9897);
xor U10286 (N_10286,N_9612,N_10074);
nor U10287 (N_10287,N_9822,N_9726);
nand U10288 (N_10288,N_9722,N_9773);
nand U10289 (N_10289,N_9970,N_9816);
xnor U10290 (N_10290,N_9955,N_9678);
and U10291 (N_10291,N_10128,N_9686);
or U10292 (N_10292,N_9804,N_9640);
nand U10293 (N_10293,N_9785,N_9817);
xor U10294 (N_10294,N_9815,N_9769);
xnor U10295 (N_10295,N_9611,N_9848);
or U10296 (N_10296,N_10112,N_10091);
or U10297 (N_10297,N_9724,N_10114);
and U10298 (N_10298,N_10145,N_9927);
nor U10299 (N_10299,N_9907,N_9679);
nand U10300 (N_10300,N_9903,N_9708);
nand U10301 (N_10301,N_10025,N_9823);
nand U10302 (N_10302,N_9856,N_10039);
and U10303 (N_10303,N_9891,N_9663);
and U10304 (N_10304,N_9719,N_9980);
or U10305 (N_10305,N_9613,N_9728);
nand U10306 (N_10306,N_9605,N_10046);
and U10307 (N_10307,N_10167,N_9767);
nand U10308 (N_10308,N_9878,N_9702);
and U10309 (N_10309,N_9805,N_10018);
xor U10310 (N_10310,N_9789,N_9911);
nand U10311 (N_10311,N_10092,N_9915);
nor U10312 (N_10312,N_9776,N_9737);
nor U10313 (N_10313,N_9664,N_10163);
nor U10314 (N_10314,N_9690,N_9812);
nand U10315 (N_10315,N_9828,N_10158);
nor U10316 (N_10316,N_10120,N_9614);
nand U10317 (N_10317,N_9631,N_9880);
or U10318 (N_10318,N_9865,N_9654);
xnor U10319 (N_10319,N_10179,N_9998);
and U10320 (N_10320,N_10058,N_9921);
nor U10321 (N_10321,N_9758,N_10159);
and U10322 (N_10322,N_9707,N_10132);
nand U10323 (N_10323,N_10127,N_10100);
xor U10324 (N_10324,N_10105,N_9879);
nor U10325 (N_10325,N_10078,N_10182);
nor U10326 (N_10326,N_9870,N_10143);
and U10327 (N_10327,N_9705,N_9966);
and U10328 (N_10328,N_10064,N_10156);
or U10329 (N_10329,N_10081,N_10144);
nor U10330 (N_10330,N_10045,N_9778);
or U10331 (N_10331,N_9981,N_10161);
or U10332 (N_10332,N_9913,N_10136);
or U10333 (N_10333,N_9853,N_10130);
and U10334 (N_10334,N_9959,N_9681);
nand U10335 (N_10335,N_9863,N_9751);
and U10336 (N_10336,N_9917,N_9641);
nor U10337 (N_10337,N_9930,N_9723);
or U10338 (N_10338,N_10087,N_9624);
xor U10339 (N_10339,N_9884,N_9920);
xnor U10340 (N_10340,N_9939,N_9609);
and U10341 (N_10341,N_9834,N_9635);
nand U10342 (N_10342,N_10014,N_9944);
xnor U10343 (N_10343,N_9747,N_9838);
xnor U10344 (N_10344,N_9783,N_10065);
and U10345 (N_10345,N_9937,N_9857);
xnor U10346 (N_10346,N_9618,N_10038);
xnor U10347 (N_10347,N_10172,N_9800);
xnor U10348 (N_10348,N_9736,N_9820);
nor U10349 (N_10349,N_10061,N_9852);
nor U10350 (N_10350,N_9962,N_9902);
or U10351 (N_10351,N_10059,N_9985);
nand U10352 (N_10352,N_9630,N_9900);
or U10353 (N_10353,N_9753,N_9840);
or U10354 (N_10354,N_10012,N_10086);
and U10355 (N_10355,N_10193,N_9752);
nor U10356 (N_10356,N_9735,N_9687);
or U10357 (N_10357,N_10015,N_10023);
or U10358 (N_10358,N_9796,N_9683);
or U10359 (N_10359,N_9810,N_10009);
nor U10360 (N_10360,N_9625,N_9616);
or U10361 (N_10361,N_9740,N_10111);
and U10362 (N_10362,N_9627,N_10196);
nor U10363 (N_10363,N_9964,N_10011);
and U10364 (N_10364,N_10149,N_9639);
nand U10365 (N_10365,N_10153,N_9775);
nor U10366 (N_10366,N_9846,N_10041);
nand U10367 (N_10367,N_9643,N_9847);
nand U10368 (N_10368,N_10032,N_9650);
or U10369 (N_10369,N_10186,N_9889);
or U10370 (N_10370,N_9781,N_9696);
xnor U10371 (N_10371,N_9754,N_9996);
or U10372 (N_10372,N_9910,N_9667);
nand U10373 (N_10373,N_9714,N_9901);
and U10374 (N_10374,N_10085,N_10008);
or U10375 (N_10375,N_9615,N_9923);
or U10376 (N_10376,N_9750,N_9607);
nor U10377 (N_10377,N_9859,N_10140);
nor U10378 (N_10378,N_9951,N_9914);
or U10379 (N_10379,N_9973,N_9864);
or U10380 (N_10380,N_10017,N_10024);
nand U10381 (N_10381,N_10083,N_9861);
nand U10382 (N_10382,N_10198,N_9770);
or U10383 (N_10383,N_9842,N_9908);
and U10384 (N_10384,N_9983,N_10035);
nor U10385 (N_10385,N_9746,N_9798);
nor U10386 (N_10386,N_9894,N_10053);
xnor U10387 (N_10387,N_9620,N_10108);
nor U10388 (N_10388,N_10168,N_10033);
nor U10389 (N_10389,N_10199,N_9803);
nand U10390 (N_10390,N_9995,N_9784);
nor U10391 (N_10391,N_9704,N_9953);
nand U10392 (N_10392,N_9695,N_10051);
nand U10393 (N_10393,N_9703,N_9670);
nor U10394 (N_10394,N_10150,N_9948);
and U10395 (N_10395,N_9987,N_9877);
or U10396 (N_10396,N_9644,N_9950);
nand U10397 (N_10397,N_9874,N_9875);
nand U10398 (N_10398,N_9858,N_9936);
xnor U10399 (N_10399,N_9888,N_10164);
xnor U10400 (N_10400,N_9946,N_10073);
xor U10401 (N_10401,N_9909,N_9779);
and U10402 (N_10402,N_9763,N_9963);
nor U10403 (N_10403,N_10115,N_9833);
or U10404 (N_10404,N_9677,N_9645);
or U10405 (N_10405,N_10101,N_9626);
and U10406 (N_10406,N_10110,N_9824);
nand U10407 (N_10407,N_9818,N_9791);
or U10408 (N_10408,N_9855,N_10142);
xor U10409 (N_10409,N_10062,N_10147);
and U10410 (N_10410,N_9646,N_9692);
and U10411 (N_10411,N_9965,N_10089);
and U10412 (N_10412,N_9706,N_9918);
xor U10413 (N_10413,N_9749,N_9826);
and U10414 (N_10414,N_9760,N_9979);
nand U10415 (N_10415,N_10066,N_10094);
or U10416 (N_10416,N_9956,N_10117);
xor U10417 (N_10417,N_10118,N_9701);
and U10418 (N_10418,N_9610,N_10056);
and U10419 (N_10419,N_9851,N_9899);
or U10420 (N_10420,N_10185,N_9876);
xnor U10421 (N_10421,N_10028,N_10162);
and U10422 (N_10422,N_10095,N_10026);
or U10423 (N_10423,N_10122,N_9647);
xnor U10424 (N_10424,N_10075,N_9924);
nand U10425 (N_10425,N_10054,N_10195);
and U10426 (N_10426,N_9674,N_9662);
nand U10427 (N_10427,N_10181,N_9777);
nor U10428 (N_10428,N_9676,N_9694);
or U10429 (N_10429,N_10190,N_9638);
nand U10430 (N_10430,N_9797,N_10194);
nor U10431 (N_10431,N_9928,N_9836);
nor U10432 (N_10432,N_10072,N_9978);
nor U10433 (N_10433,N_9782,N_9699);
nor U10434 (N_10434,N_10000,N_9637);
and U10435 (N_10435,N_10113,N_9771);
nand U10436 (N_10436,N_9697,N_10124);
nand U10437 (N_10437,N_9657,N_10004);
xnor U10438 (N_10438,N_10125,N_9673);
nor U10439 (N_10439,N_9757,N_10027);
nand U10440 (N_10440,N_9886,N_10037);
nor U10441 (N_10441,N_9671,N_10067);
nor U10442 (N_10442,N_10138,N_9642);
nand U10443 (N_10443,N_9765,N_9860);
and U10444 (N_10444,N_10121,N_9666);
or U10445 (N_10445,N_9808,N_9934);
or U10446 (N_10446,N_10068,N_10157);
and U10447 (N_10447,N_10001,N_10029);
nor U10448 (N_10448,N_10174,N_10040);
xnor U10449 (N_10449,N_10191,N_9621);
xor U10450 (N_10450,N_9658,N_9793);
nand U10451 (N_10451,N_10187,N_10175);
nor U10452 (N_10452,N_9942,N_10052);
and U10453 (N_10453,N_9731,N_9684);
nand U10454 (N_10454,N_9710,N_9685);
and U10455 (N_10455,N_9926,N_9742);
and U10456 (N_10456,N_10082,N_10036);
and U10457 (N_10457,N_9898,N_10076);
nor U10458 (N_10458,N_9992,N_10148);
and U10459 (N_10459,N_10069,N_9994);
or U10460 (N_10460,N_9943,N_10007);
nor U10461 (N_10461,N_9814,N_9606);
or U10462 (N_10462,N_10177,N_9896);
xnor U10463 (N_10463,N_9832,N_10133);
and U10464 (N_10464,N_9905,N_10119);
or U10465 (N_10465,N_9843,N_9999);
or U10466 (N_10466,N_9841,N_10020);
and U10467 (N_10467,N_9960,N_9761);
nor U10468 (N_10468,N_9665,N_9904);
or U10469 (N_10469,N_10109,N_9794);
and U10470 (N_10470,N_9712,N_10152);
or U10471 (N_10471,N_9801,N_9977);
xnor U10472 (N_10472,N_10090,N_9733);
nor U10473 (N_10473,N_10171,N_9716);
nor U10474 (N_10474,N_9788,N_10155);
nor U10475 (N_10475,N_10104,N_9976);
nor U10476 (N_10476,N_9672,N_9732);
xnor U10477 (N_10477,N_9835,N_10139);
xnor U10478 (N_10478,N_9893,N_9655);
and U10479 (N_10479,N_9622,N_9792);
nand U10480 (N_10480,N_10070,N_10022);
xnor U10481 (N_10481,N_9890,N_9721);
or U10482 (N_10482,N_10080,N_9766);
xor U10483 (N_10483,N_9649,N_9632);
nor U10484 (N_10484,N_10030,N_9867);
xor U10485 (N_10485,N_10057,N_9990);
or U10486 (N_10486,N_9602,N_10099);
nor U10487 (N_10487,N_10135,N_10021);
nand U10488 (N_10488,N_9945,N_10103);
or U10489 (N_10489,N_9819,N_10010);
and U10490 (N_10490,N_9809,N_9601);
and U10491 (N_10491,N_9745,N_9759);
or U10492 (N_10492,N_9680,N_10003);
nand U10493 (N_10493,N_9862,N_9691);
nor U10494 (N_10494,N_10055,N_9932);
xor U10495 (N_10495,N_10049,N_9659);
xnor U10496 (N_10496,N_9873,N_10002);
or U10497 (N_10497,N_9933,N_9700);
xnor U10498 (N_10498,N_10107,N_9730);
nand U10499 (N_10499,N_10180,N_10050);
or U10500 (N_10500,N_9652,N_9678);
nor U10501 (N_10501,N_9748,N_10035);
or U10502 (N_10502,N_10048,N_9867);
and U10503 (N_10503,N_9705,N_9836);
nor U10504 (N_10504,N_9623,N_9620);
nor U10505 (N_10505,N_9636,N_10149);
nand U10506 (N_10506,N_10042,N_10107);
or U10507 (N_10507,N_10157,N_9652);
or U10508 (N_10508,N_9820,N_10070);
or U10509 (N_10509,N_9616,N_10071);
nor U10510 (N_10510,N_10131,N_10127);
or U10511 (N_10511,N_9653,N_9650);
or U10512 (N_10512,N_10156,N_9787);
nor U10513 (N_10513,N_9938,N_10131);
or U10514 (N_10514,N_9669,N_9740);
nor U10515 (N_10515,N_9937,N_9806);
xor U10516 (N_10516,N_10092,N_10022);
nor U10517 (N_10517,N_9751,N_9930);
and U10518 (N_10518,N_10197,N_9607);
xor U10519 (N_10519,N_9913,N_9711);
nand U10520 (N_10520,N_9628,N_9776);
xor U10521 (N_10521,N_9811,N_9693);
xnor U10522 (N_10522,N_9622,N_10181);
or U10523 (N_10523,N_9685,N_9840);
nor U10524 (N_10524,N_9953,N_10156);
nand U10525 (N_10525,N_9742,N_9961);
xor U10526 (N_10526,N_9925,N_9865);
or U10527 (N_10527,N_9677,N_9713);
or U10528 (N_10528,N_10129,N_10049);
and U10529 (N_10529,N_10107,N_9778);
or U10530 (N_10530,N_10172,N_9708);
nor U10531 (N_10531,N_9976,N_10119);
xor U10532 (N_10532,N_10073,N_10172);
xnor U10533 (N_10533,N_10035,N_9757);
xnor U10534 (N_10534,N_9718,N_9707);
xor U10535 (N_10535,N_9874,N_9622);
nand U10536 (N_10536,N_10095,N_10088);
or U10537 (N_10537,N_9995,N_9782);
nand U10538 (N_10538,N_10169,N_9905);
and U10539 (N_10539,N_10096,N_10088);
xor U10540 (N_10540,N_9648,N_9836);
xor U10541 (N_10541,N_9631,N_9622);
nor U10542 (N_10542,N_9628,N_9694);
nor U10543 (N_10543,N_10121,N_10177);
and U10544 (N_10544,N_10011,N_9661);
nand U10545 (N_10545,N_10147,N_9940);
or U10546 (N_10546,N_10009,N_9719);
or U10547 (N_10547,N_10100,N_9837);
nor U10548 (N_10548,N_9994,N_9891);
nand U10549 (N_10549,N_9898,N_9607);
nand U10550 (N_10550,N_9824,N_9843);
or U10551 (N_10551,N_10012,N_9832);
nand U10552 (N_10552,N_9766,N_10188);
nand U10553 (N_10553,N_9853,N_9872);
and U10554 (N_10554,N_10081,N_9620);
nand U10555 (N_10555,N_9764,N_9846);
nor U10556 (N_10556,N_9762,N_10076);
xnor U10557 (N_10557,N_9805,N_10127);
nand U10558 (N_10558,N_9673,N_9931);
xor U10559 (N_10559,N_9800,N_10023);
xnor U10560 (N_10560,N_9703,N_9632);
xor U10561 (N_10561,N_10022,N_10148);
xor U10562 (N_10562,N_9611,N_10160);
or U10563 (N_10563,N_10174,N_9976);
nand U10564 (N_10564,N_9943,N_9926);
nand U10565 (N_10565,N_9729,N_9774);
nor U10566 (N_10566,N_9961,N_9896);
and U10567 (N_10567,N_9993,N_9692);
xnor U10568 (N_10568,N_9692,N_9961);
and U10569 (N_10569,N_9959,N_10178);
and U10570 (N_10570,N_9645,N_9972);
nand U10571 (N_10571,N_10161,N_10014);
nor U10572 (N_10572,N_9948,N_10177);
and U10573 (N_10573,N_10034,N_9605);
and U10574 (N_10574,N_9710,N_10171);
nand U10575 (N_10575,N_10089,N_10007);
nor U10576 (N_10576,N_9846,N_9835);
nand U10577 (N_10577,N_9978,N_10191);
nor U10578 (N_10578,N_9909,N_9876);
nand U10579 (N_10579,N_9755,N_9655);
nor U10580 (N_10580,N_9709,N_9873);
xor U10581 (N_10581,N_10051,N_9788);
nand U10582 (N_10582,N_9762,N_9849);
nand U10583 (N_10583,N_10094,N_9600);
and U10584 (N_10584,N_9649,N_9637);
xor U10585 (N_10585,N_9949,N_9737);
and U10586 (N_10586,N_9788,N_10180);
and U10587 (N_10587,N_10175,N_9739);
xnor U10588 (N_10588,N_10130,N_10019);
nor U10589 (N_10589,N_9846,N_10172);
or U10590 (N_10590,N_10170,N_9887);
nand U10591 (N_10591,N_9938,N_9953);
xor U10592 (N_10592,N_9763,N_9823);
xnor U10593 (N_10593,N_10187,N_10139);
nand U10594 (N_10594,N_9794,N_9714);
xor U10595 (N_10595,N_9699,N_9717);
xor U10596 (N_10596,N_9929,N_9820);
nand U10597 (N_10597,N_10001,N_10016);
nor U10598 (N_10598,N_10025,N_9901);
xnor U10599 (N_10599,N_9712,N_10059);
and U10600 (N_10600,N_9653,N_9859);
nor U10601 (N_10601,N_9791,N_10035);
nand U10602 (N_10602,N_9744,N_10165);
and U10603 (N_10603,N_10177,N_9831);
nor U10604 (N_10604,N_10167,N_10150);
nor U10605 (N_10605,N_9861,N_10100);
and U10606 (N_10606,N_9765,N_10195);
nor U10607 (N_10607,N_10145,N_9947);
nand U10608 (N_10608,N_10184,N_9699);
nor U10609 (N_10609,N_9635,N_10164);
nand U10610 (N_10610,N_10157,N_9991);
or U10611 (N_10611,N_10168,N_10171);
xnor U10612 (N_10612,N_9682,N_9797);
and U10613 (N_10613,N_10182,N_10136);
and U10614 (N_10614,N_9646,N_9752);
nor U10615 (N_10615,N_9876,N_9703);
xnor U10616 (N_10616,N_9647,N_9776);
nand U10617 (N_10617,N_9751,N_9653);
nor U10618 (N_10618,N_10048,N_10080);
xor U10619 (N_10619,N_9955,N_9837);
nand U10620 (N_10620,N_9981,N_10157);
and U10621 (N_10621,N_9613,N_9662);
xor U10622 (N_10622,N_9806,N_9755);
nand U10623 (N_10623,N_9972,N_9981);
and U10624 (N_10624,N_9772,N_9869);
xnor U10625 (N_10625,N_10116,N_9828);
xnor U10626 (N_10626,N_10020,N_9772);
xor U10627 (N_10627,N_9923,N_9643);
or U10628 (N_10628,N_10058,N_9843);
nand U10629 (N_10629,N_9661,N_10155);
and U10630 (N_10630,N_9664,N_9885);
and U10631 (N_10631,N_9907,N_9993);
and U10632 (N_10632,N_9884,N_9893);
or U10633 (N_10633,N_10108,N_9837);
nand U10634 (N_10634,N_10121,N_9794);
or U10635 (N_10635,N_9799,N_10094);
nor U10636 (N_10636,N_10059,N_9612);
and U10637 (N_10637,N_9742,N_9806);
and U10638 (N_10638,N_10103,N_10010);
nand U10639 (N_10639,N_9994,N_9917);
and U10640 (N_10640,N_10170,N_9846);
xnor U10641 (N_10641,N_10061,N_10074);
nand U10642 (N_10642,N_9623,N_10068);
nand U10643 (N_10643,N_10006,N_9690);
or U10644 (N_10644,N_9613,N_9950);
or U10645 (N_10645,N_10000,N_9662);
or U10646 (N_10646,N_10031,N_9632);
or U10647 (N_10647,N_10175,N_10143);
and U10648 (N_10648,N_9896,N_10069);
nor U10649 (N_10649,N_10154,N_9816);
nor U10650 (N_10650,N_9726,N_9832);
and U10651 (N_10651,N_9866,N_9845);
nand U10652 (N_10652,N_9880,N_10067);
or U10653 (N_10653,N_10119,N_9603);
nor U10654 (N_10654,N_9918,N_10092);
xnor U10655 (N_10655,N_9693,N_9711);
and U10656 (N_10656,N_10026,N_9761);
xor U10657 (N_10657,N_10022,N_10155);
nand U10658 (N_10658,N_9811,N_10133);
nand U10659 (N_10659,N_9858,N_9625);
or U10660 (N_10660,N_9792,N_9623);
nand U10661 (N_10661,N_10038,N_9601);
xnor U10662 (N_10662,N_9749,N_10080);
xnor U10663 (N_10663,N_10163,N_9901);
xnor U10664 (N_10664,N_9961,N_9960);
and U10665 (N_10665,N_9951,N_9703);
nor U10666 (N_10666,N_9981,N_10067);
nor U10667 (N_10667,N_10147,N_9926);
nor U10668 (N_10668,N_9613,N_9637);
nor U10669 (N_10669,N_9996,N_9917);
or U10670 (N_10670,N_9794,N_9640);
nand U10671 (N_10671,N_9993,N_10103);
xor U10672 (N_10672,N_10140,N_9709);
or U10673 (N_10673,N_9839,N_9672);
nand U10674 (N_10674,N_10153,N_9661);
nand U10675 (N_10675,N_10098,N_10136);
and U10676 (N_10676,N_10062,N_10125);
nand U10677 (N_10677,N_9693,N_9947);
nor U10678 (N_10678,N_9854,N_9973);
nand U10679 (N_10679,N_9817,N_9713);
and U10680 (N_10680,N_10003,N_10038);
xor U10681 (N_10681,N_9861,N_9817);
nor U10682 (N_10682,N_10015,N_10082);
and U10683 (N_10683,N_10157,N_9787);
xor U10684 (N_10684,N_9936,N_9623);
nor U10685 (N_10685,N_9969,N_9716);
nand U10686 (N_10686,N_10184,N_10029);
and U10687 (N_10687,N_9776,N_10066);
nor U10688 (N_10688,N_9724,N_10144);
xor U10689 (N_10689,N_10079,N_9962);
nor U10690 (N_10690,N_10178,N_10013);
and U10691 (N_10691,N_9737,N_10020);
or U10692 (N_10692,N_10069,N_10136);
nor U10693 (N_10693,N_9628,N_10020);
nand U10694 (N_10694,N_9863,N_9995);
nor U10695 (N_10695,N_10075,N_9826);
nand U10696 (N_10696,N_9888,N_9755);
nand U10697 (N_10697,N_10084,N_10089);
xor U10698 (N_10698,N_10127,N_10196);
xor U10699 (N_10699,N_9984,N_9825);
and U10700 (N_10700,N_9759,N_9832);
nand U10701 (N_10701,N_9711,N_9626);
and U10702 (N_10702,N_9977,N_9616);
xor U10703 (N_10703,N_9817,N_9932);
or U10704 (N_10704,N_9723,N_10051);
and U10705 (N_10705,N_10189,N_9739);
and U10706 (N_10706,N_9629,N_10109);
xor U10707 (N_10707,N_9773,N_9920);
nand U10708 (N_10708,N_10181,N_9941);
and U10709 (N_10709,N_9886,N_9818);
or U10710 (N_10710,N_9604,N_10155);
xnor U10711 (N_10711,N_9847,N_9893);
and U10712 (N_10712,N_10107,N_9604);
xor U10713 (N_10713,N_9737,N_9755);
and U10714 (N_10714,N_9951,N_10180);
xnor U10715 (N_10715,N_10049,N_9923);
xor U10716 (N_10716,N_9884,N_10130);
nor U10717 (N_10717,N_10178,N_9824);
nor U10718 (N_10718,N_9653,N_10006);
and U10719 (N_10719,N_9944,N_9964);
xor U10720 (N_10720,N_9918,N_9814);
nor U10721 (N_10721,N_9625,N_10148);
xor U10722 (N_10722,N_10069,N_10053);
and U10723 (N_10723,N_9757,N_10172);
or U10724 (N_10724,N_9980,N_9899);
nor U10725 (N_10725,N_9618,N_9945);
nor U10726 (N_10726,N_9965,N_9970);
and U10727 (N_10727,N_10127,N_10040);
nor U10728 (N_10728,N_10070,N_10040);
xnor U10729 (N_10729,N_9857,N_9633);
xor U10730 (N_10730,N_9634,N_9613);
nand U10731 (N_10731,N_10182,N_10165);
xnor U10732 (N_10732,N_10104,N_9769);
and U10733 (N_10733,N_10120,N_10092);
and U10734 (N_10734,N_10124,N_9699);
or U10735 (N_10735,N_9930,N_9767);
nor U10736 (N_10736,N_9699,N_9799);
or U10737 (N_10737,N_9719,N_10059);
nand U10738 (N_10738,N_9824,N_9842);
or U10739 (N_10739,N_9804,N_9647);
nand U10740 (N_10740,N_9692,N_10149);
xor U10741 (N_10741,N_9822,N_10072);
nor U10742 (N_10742,N_9782,N_9921);
nand U10743 (N_10743,N_9878,N_9900);
and U10744 (N_10744,N_10042,N_9736);
nand U10745 (N_10745,N_9721,N_10028);
nor U10746 (N_10746,N_10021,N_9671);
xnor U10747 (N_10747,N_9675,N_9986);
nand U10748 (N_10748,N_9625,N_10041);
nand U10749 (N_10749,N_9847,N_10040);
nor U10750 (N_10750,N_10063,N_10179);
or U10751 (N_10751,N_9650,N_10117);
or U10752 (N_10752,N_9855,N_10093);
xor U10753 (N_10753,N_10025,N_9716);
and U10754 (N_10754,N_9865,N_9617);
nor U10755 (N_10755,N_9924,N_9618);
and U10756 (N_10756,N_10014,N_9785);
xor U10757 (N_10757,N_9872,N_9795);
nand U10758 (N_10758,N_9656,N_9625);
nor U10759 (N_10759,N_9861,N_9724);
nand U10760 (N_10760,N_10062,N_9814);
xor U10761 (N_10761,N_10000,N_10066);
nor U10762 (N_10762,N_9991,N_9800);
nand U10763 (N_10763,N_9851,N_9794);
nor U10764 (N_10764,N_9991,N_9618);
nor U10765 (N_10765,N_10101,N_9965);
or U10766 (N_10766,N_9821,N_9740);
nor U10767 (N_10767,N_9904,N_9640);
and U10768 (N_10768,N_10178,N_10076);
or U10769 (N_10769,N_10107,N_9632);
xnor U10770 (N_10770,N_9659,N_9939);
nor U10771 (N_10771,N_9870,N_9875);
nand U10772 (N_10772,N_9868,N_10160);
nor U10773 (N_10773,N_9941,N_9983);
or U10774 (N_10774,N_9692,N_9974);
nor U10775 (N_10775,N_9814,N_9888);
nor U10776 (N_10776,N_10030,N_10038);
nand U10777 (N_10777,N_9627,N_10054);
nand U10778 (N_10778,N_9674,N_9978);
and U10779 (N_10779,N_10069,N_9652);
and U10780 (N_10780,N_9911,N_9694);
nand U10781 (N_10781,N_9954,N_9817);
or U10782 (N_10782,N_10007,N_9637);
xor U10783 (N_10783,N_9736,N_10124);
or U10784 (N_10784,N_9838,N_9982);
and U10785 (N_10785,N_9669,N_9698);
xor U10786 (N_10786,N_9631,N_9817);
nor U10787 (N_10787,N_10154,N_9774);
nand U10788 (N_10788,N_9654,N_9722);
or U10789 (N_10789,N_10124,N_9682);
nor U10790 (N_10790,N_10114,N_9629);
and U10791 (N_10791,N_9838,N_9874);
and U10792 (N_10792,N_9984,N_10045);
xor U10793 (N_10793,N_9704,N_9827);
xor U10794 (N_10794,N_10117,N_9813);
and U10795 (N_10795,N_9897,N_9673);
or U10796 (N_10796,N_9968,N_10060);
or U10797 (N_10797,N_10108,N_10024);
and U10798 (N_10798,N_9999,N_9766);
nor U10799 (N_10799,N_10117,N_9938);
nand U10800 (N_10800,N_10520,N_10560);
and U10801 (N_10801,N_10705,N_10353);
nand U10802 (N_10802,N_10262,N_10258);
and U10803 (N_10803,N_10625,N_10530);
nand U10804 (N_10804,N_10278,N_10314);
xnor U10805 (N_10805,N_10698,N_10539);
nand U10806 (N_10806,N_10462,N_10292);
and U10807 (N_10807,N_10207,N_10521);
nor U10808 (N_10808,N_10431,N_10397);
nand U10809 (N_10809,N_10382,N_10685);
xor U10810 (N_10810,N_10387,N_10799);
nor U10811 (N_10811,N_10457,N_10343);
xor U10812 (N_10812,N_10384,N_10205);
xor U10813 (N_10813,N_10246,N_10307);
nand U10814 (N_10814,N_10360,N_10671);
nor U10815 (N_10815,N_10612,N_10613);
nor U10816 (N_10816,N_10363,N_10789);
or U10817 (N_10817,N_10794,N_10589);
nand U10818 (N_10818,N_10726,N_10237);
and U10819 (N_10819,N_10713,N_10779);
xnor U10820 (N_10820,N_10433,N_10471);
nor U10821 (N_10821,N_10432,N_10646);
nor U10822 (N_10822,N_10504,N_10531);
nor U10823 (N_10823,N_10308,N_10265);
and U10824 (N_10824,N_10655,N_10489);
and U10825 (N_10825,N_10320,N_10275);
and U10826 (N_10826,N_10649,N_10730);
and U10827 (N_10827,N_10456,N_10700);
nand U10828 (N_10828,N_10426,N_10510);
and U10829 (N_10829,N_10774,N_10249);
and U10830 (N_10830,N_10399,N_10715);
nor U10831 (N_10831,N_10256,N_10621);
and U10832 (N_10832,N_10543,N_10230);
and U10833 (N_10833,N_10264,N_10326);
nand U10834 (N_10834,N_10344,N_10466);
and U10835 (N_10835,N_10744,N_10712);
and U10836 (N_10836,N_10672,N_10358);
nand U10837 (N_10837,N_10518,N_10409);
or U10838 (N_10838,N_10599,N_10651);
xnor U10839 (N_10839,N_10381,N_10354);
nor U10840 (N_10840,N_10757,N_10351);
or U10841 (N_10841,N_10272,N_10291);
xnor U10842 (N_10842,N_10626,N_10514);
and U10843 (N_10843,N_10670,N_10372);
xnor U10844 (N_10844,N_10238,N_10405);
or U10845 (N_10845,N_10785,N_10214);
or U10846 (N_10846,N_10577,N_10483);
or U10847 (N_10847,N_10711,N_10355);
and U10848 (N_10848,N_10380,N_10622);
nand U10849 (N_10849,N_10460,N_10224);
nor U10850 (N_10850,N_10547,N_10250);
xnor U10851 (N_10851,N_10459,N_10290);
xnor U10852 (N_10852,N_10691,N_10487);
xnor U10853 (N_10853,N_10748,N_10758);
xor U10854 (N_10854,N_10346,N_10368);
or U10855 (N_10855,N_10310,N_10442);
and U10856 (N_10856,N_10552,N_10282);
nand U10857 (N_10857,N_10745,N_10479);
nor U10858 (N_10858,N_10413,N_10777);
xor U10859 (N_10859,N_10367,N_10721);
xnor U10860 (N_10860,N_10752,N_10274);
xor U10861 (N_10861,N_10443,N_10753);
nor U10862 (N_10862,N_10534,N_10614);
and U10863 (N_10863,N_10775,N_10682);
and U10864 (N_10864,N_10505,N_10760);
or U10865 (N_10865,N_10338,N_10780);
nand U10866 (N_10866,N_10349,N_10475);
nand U10867 (N_10867,N_10664,N_10464);
xnor U10868 (N_10868,N_10203,N_10316);
and U10869 (N_10869,N_10683,N_10782);
nand U10870 (N_10870,N_10647,N_10605);
or U10871 (N_10871,N_10241,N_10554);
xor U10872 (N_10872,N_10796,N_10564);
nor U10873 (N_10873,N_10473,N_10635);
xnor U10874 (N_10874,N_10490,N_10301);
and U10875 (N_10875,N_10669,N_10379);
xor U10876 (N_10876,N_10707,N_10731);
xnor U10877 (N_10877,N_10798,N_10773);
and U10878 (N_10878,N_10394,N_10425);
nand U10879 (N_10879,N_10364,N_10660);
nand U10880 (N_10880,N_10632,N_10766);
or U10881 (N_10881,N_10268,N_10716);
nand U10882 (N_10882,N_10797,N_10681);
or U10883 (N_10883,N_10347,N_10763);
and U10884 (N_10884,N_10677,N_10269);
xnor U10885 (N_10885,N_10486,N_10735);
nor U10886 (N_10886,N_10550,N_10508);
nor U10887 (N_10887,N_10759,N_10689);
xnor U10888 (N_10888,N_10311,N_10279);
xor U10889 (N_10889,N_10704,N_10319);
nand U10890 (N_10890,N_10538,N_10200);
xnor U10891 (N_10891,N_10213,N_10401);
nand U10892 (N_10892,N_10450,N_10255);
or U10893 (N_10893,N_10580,N_10586);
and U10894 (N_10894,N_10556,N_10416);
and U10895 (N_10895,N_10678,N_10693);
xnor U10896 (N_10896,N_10666,N_10574);
and U10897 (N_10897,N_10403,N_10225);
nand U10898 (N_10898,N_10545,N_10616);
xnor U10899 (N_10899,N_10417,N_10506);
nor U10900 (N_10900,N_10211,N_10484);
nand U10901 (N_10901,N_10708,N_10451);
nand U10902 (N_10902,N_10595,N_10388);
and U10903 (N_10903,N_10219,N_10458);
xnor U10904 (N_10904,N_10212,N_10369);
and U10905 (N_10905,N_10667,N_10428);
or U10906 (N_10906,N_10267,N_10640);
or U10907 (N_10907,N_10260,N_10566);
or U10908 (N_10908,N_10551,N_10688);
xnor U10909 (N_10909,N_10648,N_10598);
and U10910 (N_10910,N_10631,N_10216);
and U10911 (N_10911,N_10680,N_10630);
nand U10912 (N_10912,N_10289,N_10546);
and U10913 (N_10913,N_10657,N_10247);
nor U10914 (N_10914,N_10732,N_10366);
xor U10915 (N_10915,N_10350,N_10561);
or U10916 (N_10916,N_10668,N_10422);
nand U10917 (N_10917,N_10628,N_10209);
nor U10918 (N_10918,N_10576,N_10529);
nand U10919 (N_10919,N_10424,N_10714);
xnor U10920 (N_10920,N_10581,N_10513);
nand U10921 (N_10921,N_10468,N_10607);
and U10922 (N_10922,N_10788,N_10270);
xor U10923 (N_10923,N_10597,N_10341);
xor U10924 (N_10924,N_10340,N_10724);
nand U10925 (N_10925,N_10309,N_10563);
xnor U10926 (N_10926,N_10567,N_10378);
nor U10927 (N_10927,N_10624,N_10485);
nor U10928 (N_10928,N_10588,N_10527);
and U10929 (N_10929,N_10562,N_10786);
nor U10930 (N_10930,N_10277,N_10604);
nor U10931 (N_10931,N_10488,N_10697);
xor U10932 (N_10932,N_10575,N_10661);
nor U10933 (N_10933,N_10359,N_10374);
or U10934 (N_10934,N_10227,N_10734);
and U10935 (N_10935,N_10480,N_10755);
and U10936 (N_10936,N_10396,N_10283);
and U10937 (N_10937,N_10694,N_10411);
and U10938 (N_10938,N_10402,N_10421);
or U10939 (N_10939,N_10315,N_10699);
and U10940 (N_10940,N_10727,N_10645);
and U10941 (N_10941,N_10717,N_10204);
or U10942 (N_10942,N_10474,N_10537);
nand U10943 (N_10943,N_10558,N_10373);
nand U10944 (N_10944,N_10617,N_10463);
and U10945 (N_10945,N_10702,N_10342);
nor U10946 (N_10946,N_10516,N_10610);
nor U10947 (N_10947,N_10582,N_10541);
nand U10948 (N_10948,N_10511,N_10594);
nor U10949 (N_10949,N_10438,N_10492);
nand U10950 (N_10950,N_10754,N_10454);
and U10951 (N_10951,N_10477,N_10536);
nand U10952 (N_10952,N_10410,N_10592);
nand U10953 (N_10953,N_10749,N_10601);
nand U10954 (N_10954,N_10352,N_10776);
or U10955 (N_10955,N_10494,N_10792);
or U10956 (N_10956,N_10679,N_10652);
nand U10957 (N_10957,N_10495,N_10642);
nand U10958 (N_10958,N_10201,N_10619);
xor U10959 (N_10959,N_10781,N_10294);
and U10960 (N_10960,N_10312,N_10331);
nor U10961 (N_10961,N_10623,N_10345);
nand U10962 (N_10962,N_10427,N_10254);
nand U10963 (N_10963,N_10235,N_10447);
nand U10964 (N_10964,N_10287,N_10523);
nand U10965 (N_10965,N_10362,N_10765);
or U10966 (N_10966,N_10634,N_10728);
and U10967 (N_10967,N_10687,N_10305);
or U10968 (N_10968,N_10606,N_10418);
nor U10969 (N_10969,N_10787,N_10257);
nand U10970 (N_10970,N_10240,N_10673);
or U10971 (N_10971,N_10318,N_10503);
or U10972 (N_10972,N_10482,N_10528);
or U10973 (N_10973,N_10720,N_10676);
and U10974 (N_10974,N_10220,N_10361);
nor U10975 (N_10975,N_10709,N_10633);
nand U10976 (N_10976,N_10502,N_10453);
or U10977 (N_10977,N_10217,N_10740);
nand U10978 (N_10978,N_10725,N_10579);
and U10979 (N_10979,N_10747,N_10519);
nor U10980 (N_10980,N_10750,N_10448);
xnor U10981 (N_10981,N_10242,N_10334);
nor U10982 (N_10982,N_10446,N_10583);
and U10983 (N_10983,N_10659,N_10286);
xnor U10984 (N_10984,N_10674,N_10557);
nor U10985 (N_10985,N_10584,N_10650);
xor U10986 (N_10986,N_10578,N_10791);
xnor U10987 (N_10987,N_10415,N_10498);
nand U10988 (N_10988,N_10703,N_10441);
xnor U10989 (N_10989,N_10232,N_10675);
nand U10990 (N_10990,N_10357,N_10636);
and U10991 (N_10991,N_10701,N_10284);
xor U10992 (N_10992,N_10222,N_10496);
xnor U10993 (N_10993,N_10706,N_10321);
xnor U10994 (N_10994,N_10404,N_10293);
nand U10995 (N_10995,N_10215,N_10365);
nand U10996 (N_10996,N_10393,N_10768);
or U10997 (N_10997,N_10228,N_10332);
nand U10998 (N_10998,N_10435,N_10452);
and U10999 (N_10999,N_10542,N_10375);
nor U11000 (N_11000,N_10386,N_10243);
xor U11001 (N_11001,N_10298,N_10271);
xnor U11002 (N_11002,N_10525,N_10322);
and U11003 (N_11003,N_10692,N_10587);
and U11004 (N_11004,N_10437,N_10790);
xnor U11005 (N_11005,N_10276,N_10762);
and U11006 (N_11006,N_10377,N_10221);
or U11007 (N_11007,N_10273,N_10608);
nor U11008 (N_11008,N_10500,N_10414);
nand U11009 (N_11009,N_10723,N_10304);
nand U11010 (N_11010,N_10390,N_10684);
nor U11011 (N_11011,N_10718,N_10729);
xnor U11012 (N_11012,N_10327,N_10783);
nor U11013 (N_11013,N_10423,N_10202);
or U11014 (N_11014,N_10767,N_10398);
nand U11015 (N_11015,N_10261,N_10370);
nand U11016 (N_11016,N_10507,N_10371);
nor U11017 (N_11017,N_10236,N_10764);
nor U11018 (N_11018,N_10515,N_10653);
nor U11019 (N_11019,N_10407,N_10430);
xnor U11020 (N_11020,N_10266,N_10549);
or U11021 (N_11021,N_10299,N_10348);
and U11022 (N_11022,N_10336,N_10231);
or U11023 (N_11023,N_10532,N_10429);
nor U11024 (N_11024,N_10313,N_10793);
nor U11025 (N_11025,N_10497,N_10555);
nand U11026 (N_11026,N_10253,N_10590);
nor U11027 (N_11027,N_10408,N_10695);
nand U11028 (N_11028,N_10644,N_10654);
nor U11029 (N_11029,N_10395,N_10339);
and U11030 (N_11030,N_10263,N_10565);
or U11031 (N_11031,N_10335,N_10470);
xnor U11032 (N_11032,N_10795,N_10559);
nor U11033 (N_11033,N_10285,N_10639);
nand U11034 (N_11034,N_10244,N_10696);
nand U11035 (N_11035,N_10376,N_10784);
or U11036 (N_11036,N_10736,N_10738);
xnor U11037 (N_11037,N_10722,N_10761);
or U11038 (N_11038,N_10481,N_10383);
nand U11039 (N_11039,N_10603,N_10569);
nand U11040 (N_11040,N_10434,N_10306);
nand U11041 (N_11041,N_10751,N_10288);
nand U11042 (N_11042,N_10517,N_10665);
nor U11043 (N_11043,N_10658,N_10300);
or U11044 (N_11044,N_10719,N_10280);
nor U11045 (N_11045,N_10419,N_10618);
xor U11046 (N_11046,N_10218,N_10445);
nand U11047 (N_11047,N_10449,N_10248);
nand U11048 (N_11048,N_10686,N_10444);
and U11049 (N_11049,N_10323,N_10239);
nand U11050 (N_11050,N_10302,N_10467);
and U11051 (N_11051,N_10535,N_10245);
xor U11052 (N_11052,N_10499,N_10333);
nand U11053 (N_11053,N_10206,N_10771);
xor U11054 (N_11054,N_10629,N_10406);
and U11055 (N_11055,N_10226,N_10526);
or U11056 (N_11056,N_10743,N_10328);
nor U11057 (N_11057,N_10662,N_10615);
xor U11058 (N_11058,N_10251,N_10593);
nor U11059 (N_11059,N_10472,N_10690);
xnor U11060 (N_11060,N_10746,N_10317);
and U11061 (N_11061,N_10356,N_10609);
xor U11062 (N_11062,N_10210,N_10741);
nand U11063 (N_11063,N_10572,N_10739);
or U11064 (N_11064,N_10533,N_10602);
nand U11065 (N_11065,N_10259,N_10234);
and U11066 (N_11066,N_10476,N_10436);
nor U11067 (N_11067,N_10325,N_10600);
nand U11068 (N_11068,N_10570,N_10522);
or U11069 (N_11069,N_10737,N_10420);
nor U11070 (N_11070,N_10553,N_10656);
nand U11071 (N_11071,N_10392,N_10233);
and U11072 (N_11072,N_10295,N_10573);
nand U11073 (N_11073,N_10641,N_10524);
nand U11074 (N_11074,N_10512,N_10491);
or U11075 (N_11075,N_10385,N_10337);
or U11076 (N_11076,N_10439,N_10769);
or U11077 (N_11077,N_10568,N_10548);
and U11078 (N_11078,N_10540,N_10770);
and U11079 (N_11079,N_10742,N_10229);
nand U11080 (N_11080,N_10465,N_10389);
nor U11081 (N_11081,N_10509,N_10778);
or U11082 (N_11082,N_10400,N_10281);
xnor U11083 (N_11083,N_10627,N_10663);
or U11084 (N_11084,N_10591,N_10296);
xor U11085 (N_11085,N_10493,N_10772);
xnor U11086 (N_11086,N_10611,N_10297);
and U11087 (N_11087,N_10596,N_10620);
nor U11088 (N_11088,N_10469,N_10585);
nand U11089 (N_11089,N_10710,N_10208);
and U11090 (N_11090,N_10330,N_10637);
xor U11091 (N_11091,N_10324,N_10455);
nand U11092 (N_11092,N_10571,N_10643);
nand U11093 (N_11093,N_10440,N_10303);
nand U11094 (N_11094,N_10329,N_10461);
and U11095 (N_11095,N_10756,N_10223);
or U11096 (N_11096,N_10501,N_10252);
and U11097 (N_11097,N_10544,N_10638);
nand U11098 (N_11098,N_10412,N_10391);
or U11099 (N_11099,N_10733,N_10478);
and U11100 (N_11100,N_10416,N_10310);
or U11101 (N_11101,N_10743,N_10419);
nor U11102 (N_11102,N_10752,N_10412);
nand U11103 (N_11103,N_10514,N_10458);
nand U11104 (N_11104,N_10392,N_10753);
nand U11105 (N_11105,N_10393,N_10717);
and U11106 (N_11106,N_10285,N_10682);
nor U11107 (N_11107,N_10551,N_10454);
and U11108 (N_11108,N_10273,N_10200);
and U11109 (N_11109,N_10242,N_10534);
and U11110 (N_11110,N_10704,N_10680);
nand U11111 (N_11111,N_10388,N_10454);
nor U11112 (N_11112,N_10644,N_10251);
nor U11113 (N_11113,N_10717,N_10363);
nor U11114 (N_11114,N_10289,N_10487);
or U11115 (N_11115,N_10647,N_10297);
xor U11116 (N_11116,N_10289,N_10426);
and U11117 (N_11117,N_10349,N_10240);
nor U11118 (N_11118,N_10764,N_10507);
or U11119 (N_11119,N_10293,N_10642);
nor U11120 (N_11120,N_10622,N_10575);
or U11121 (N_11121,N_10746,N_10304);
nand U11122 (N_11122,N_10341,N_10675);
nand U11123 (N_11123,N_10325,N_10577);
or U11124 (N_11124,N_10438,N_10298);
and U11125 (N_11125,N_10436,N_10344);
nand U11126 (N_11126,N_10449,N_10240);
or U11127 (N_11127,N_10345,N_10237);
nor U11128 (N_11128,N_10544,N_10569);
nor U11129 (N_11129,N_10324,N_10462);
nand U11130 (N_11130,N_10724,N_10625);
xor U11131 (N_11131,N_10204,N_10635);
or U11132 (N_11132,N_10484,N_10436);
nand U11133 (N_11133,N_10676,N_10678);
nor U11134 (N_11134,N_10680,N_10281);
nor U11135 (N_11135,N_10767,N_10513);
nor U11136 (N_11136,N_10671,N_10380);
or U11137 (N_11137,N_10489,N_10466);
xor U11138 (N_11138,N_10514,N_10290);
and U11139 (N_11139,N_10512,N_10233);
or U11140 (N_11140,N_10262,N_10284);
xnor U11141 (N_11141,N_10442,N_10784);
nor U11142 (N_11142,N_10259,N_10445);
nor U11143 (N_11143,N_10239,N_10798);
or U11144 (N_11144,N_10745,N_10580);
and U11145 (N_11145,N_10254,N_10211);
nor U11146 (N_11146,N_10215,N_10633);
and U11147 (N_11147,N_10752,N_10669);
nand U11148 (N_11148,N_10298,N_10367);
and U11149 (N_11149,N_10486,N_10309);
nand U11150 (N_11150,N_10731,N_10558);
nand U11151 (N_11151,N_10474,N_10271);
or U11152 (N_11152,N_10537,N_10200);
and U11153 (N_11153,N_10419,N_10341);
nor U11154 (N_11154,N_10509,N_10773);
xor U11155 (N_11155,N_10260,N_10471);
nand U11156 (N_11156,N_10766,N_10586);
nand U11157 (N_11157,N_10536,N_10529);
nor U11158 (N_11158,N_10626,N_10536);
and U11159 (N_11159,N_10314,N_10698);
xor U11160 (N_11160,N_10303,N_10434);
or U11161 (N_11161,N_10540,N_10695);
nor U11162 (N_11162,N_10464,N_10712);
xnor U11163 (N_11163,N_10241,N_10411);
and U11164 (N_11164,N_10358,N_10637);
nand U11165 (N_11165,N_10451,N_10525);
xor U11166 (N_11166,N_10308,N_10346);
or U11167 (N_11167,N_10205,N_10211);
xnor U11168 (N_11168,N_10454,N_10206);
or U11169 (N_11169,N_10369,N_10326);
and U11170 (N_11170,N_10243,N_10567);
xor U11171 (N_11171,N_10610,N_10514);
nor U11172 (N_11172,N_10485,N_10518);
nand U11173 (N_11173,N_10479,N_10655);
nand U11174 (N_11174,N_10250,N_10513);
xor U11175 (N_11175,N_10400,N_10749);
xor U11176 (N_11176,N_10547,N_10379);
nor U11177 (N_11177,N_10473,N_10661);
or U11178 (N_11178,N_10684,N_10443);
and U11179 (N_11179,N_10730,N_10395);
and U11180 (N_11180,N_10215,N_10521);
or U11181 (N_11181,N_10645,N_10666);
nor U11182 (N_11182,N_10350,N_10370);
nor U11183 (N_11183,N_10461,N_10437);
and U11184 (N_11184,N_10730,N_10538);
and U11185 (N_11185,N_10468,N_10354);
nor U11186 (N_11186,N_10303,N_10787);
and U11187 (N_11187,N_10401,N_10755);
or U11188 (N_11188,N_10446,N_10576);
xnor U11189 (N_11189,N_10698,N_10449);
nor U11190 (N_11190,N_10329,N_10260);
and U11191 (N_11191,N_10767,N_10234);
and U11192 (N_11192,N_10463,N_10380);
xor U11193 (N_11193,N_10598,N_10448);
nor U11194 (N_11194,N_10330,N_10488);
or U11195 (N_11195,N_10271,N_10411);
nor U11196 (N_11196,N_10607,N_10305);
and U11197 (N_11197,N_10549,N_10250);
or U11198 (N_11198,N_10695,N_10704);
or U11199 (N_11199,N_10552,N_10214);
or U11200 (N_11200,N_10603,N_10293);
nor U11201 (N_11201,N_10700,N_10489);
nor U11202 (N_11202,N_10479,N_10546);
or U11203 (N_11203,N_10750,N_10366);
nand U11204 (N_11204,N_10766,N_10692);
xor U11205 (N_11205,N_10590,N_10763);
nor U11206 (N_11206,N_10780,N_10371);
or U11207 (N_11207,N_10735,N_10642);
xnor U11208 (N_11208,N_10574,N_10767);
nor U11209 (N_11209,N_10583,N_10640);
and U11210 (N_11210,N_10331,N_10239);
nand U11211 (N_11211,N_10229,N_10499);
nand U11212 (N_11212,N_10568,N_10420);
and U11213 (N_11213,N_10212,N_10705);
nand U11214 (N_11214,N_10236,N_10670);
or U11215 (N_11215,N_10613,N_10677);
nand U11216 (N_11216,N_10324,N_10237);
and U11217 (N_11217,N_10310,N_10698);
nand U11218 (N_11218,N_10580,N_10267);
nand U11219 (N_11219,N_10546,N_10742);
xnor U11220 (N_11220,N_10387,N_10501);
nand U11221 (N_11221,N_10739,N_10232);
xnor U11222 (N_11222,N_10490,N_10476);
xor U11223 (N_11223,N_10672,N_10403);
xnor U11224 (N_11224,N_10542,N_10405);
xor U11225 (N_11225,N_10210,N_10554);
nor U11226 (N_11226,N_10527,N_10754);
nor U11227 (N_11227,N_10574,N_10472);
xor U11228 (N_11228,N_10320,N_10449);
and U11229 (N_11229,N_10346,N_10405);
or U11230 (N_11230,N_10454,N_10549);
and U11231 (N_11231,N_10705,N_10510);
nor U11232 (N_11232,N_10546,N_10797);
xor U11233 (N_11233,N_10619,N_10485);
nand U11234 (N_11234,N_10752,N_10252);
and U11235 (N_11235,N_10670,N_10331);
and U11236 (N_11236,N_10765,N_10573);
nand U11237 (N_11237,N_10365,N_10701);
and U11238 (N_11238,N_10445,N_10495);
and U11239 (N_11239,N_10739,N_10484);
xnor U11240 (N_11240,N_10665,N_10720);
nand U11241 (N_11241,N_10659,N_10425);
or U11242 (N_11242,N_10226,N_10304);
nand U11243 (N_11243,N_10216,N_10753);
nand U11244 (N_11244,N_10647,N_10395);
and U11245 (N_11245,N_10307,N_10699);
and U11246 (N_11246,N_10436,N_10363);
xnor U11247 (N_11247,N_10568,N_10390);
nor U11248 (N_11248,N_10780,N_10588);
nor U11249 (N_11249,N_10489,N_10568);
nand U11250 (N_11250,N_10318,N_10295);
nand U11251 (N_11251,N_10418,N_10339);
xor U11252 (N_11252,N_10370,N_10541);
nor U11253 (N_11253,N_10225,N_10210);
and U11254 (N_11254,N_10546,N_10454);
and U11255 (N_11255,N_10744,N_10359);
nand U11256 (N_11256,N_10332,N_10759);
and U11257 (N_11257,N_10235,N_10606);
nand U11258 (N_11258,N_10455,N_10553);
xor U11259 (N_11259,N_10316,N_10301);
nor U11260 (N_11260,N_10463,N_10404);
xor U11261 (N_11261,N_10329,N_10315);
xor U11262 (N_11262,N_10456,N_10382);
or U11263 (N_11263,N_10748,N_10438);
or U11264 (N_11264,N_10555,N_10232);
nor U11265 (N_11265,N_10511,N_10670);
nand U11266 (N_11266,N_10294,N_10677);
xor U11267 (N_11267,N_10234,N_10773);
and U11268 (N_11268,N_10758,N_10331);
and U11269 (N_11269,N_10517,N_10630);
and U11270 (N_11270,N_10264,N_10726);
xor U11271 (N_11271,N_10394,N_10727);
xor U11272 (N_11272,N_10770,N_10492);
or U11273 (N_11273,N_10408,N_10433);
nor U11274 (N_11274,N_10516,N_10606);
and U11275 (N_11275,N_10267,N_10352);
nor U11276 (N_11276,N_10658,N_10346);
xor U11277 (N_11277,N_10629,N_10522);
nand U11278 (N_11278,N_10582,N_10347);
or U11279 (N_11279,N_10386,N_10249);
or U11280 (N_11280,N_10374,N_10604);
nor U11281 (N_11281,N_10408,N_10341);
nand U11282 (N_11282,N_10333,N_10611);
or U11283 (N_11283,N_10730,N_10312);
xor U11284 (N_11284,N_10750,N_10687);
nor U11285 (N_11285,N_10525,N_10344);
nor U11286 (N_11286,N_10518,N_10205);
xor U11287 (N_11287,N_10216,N_10355);
nor U11288 (N_11288,N_10345,N_10460);
xnor U11289 (N_11289,N_10782,N_10321);
nand U11290 (N_11290,N_10414,N_10787);
and U11291 (N_11291,N_10373,N_10256);
or U11292 (N_11292,N_10766,N_10603);
xor U11293 (N_11293,N_10375,N_10661);
and U11294 (N_11294,N_10679,N_10554);
nor U11295 (N_11295,N_10241,N_10678);
and U11296 (N_11296,N_10369,N_10500);
nor U11297 (N_11297,N_10415,N_10218);
and U11298 (N_11298,N_10538,N_10314);
nand U11299 (N_11299,N_10400,N_10690);
nand U11300 (N_11300,N_10658,N_10642);
nand U11301 (N_11301,N_10395,N_10716);
nor U11302 (N_11302,N_10266,N_10390);
xor U11303 (N_11303,N_10527,N_10275);
nand U11304 (N_11304,N_10375,N_10366);
and U11305 (N_11305,N_10489,N_10633);
nand U11306 (N_11306,N_10454,N_10590);
nor U11307 (N_11307,N_10449,N_10437);
and U11308 (N_11308,N_10320,N_10376);
or U11309 (N_11309,N_10448,N_10440);
and U11310 (N_11310,N_10664,N_10638);
or U11311 (N_11311,N_10475,N_10255);
nand U11312 (N_11312,N_10610,N_10220);
and U11313 (N_11313,N_10759,N_10281);
xor U11314 (N_11314,N_10686,N_10573);
or U11315 (N_11315,N_10487,N_10661);
or U11316 (N_11316,N_10473,N_10287);
xnor U11317 (N_11317,N_10332,N_10251);
or U11318 (N_11318,N_10331,N_10334);
xnor U11319 (N_11319,N_10341,N_10285);
and U11320 (N_11320,N_10585,N_10695);
nand U11321 (N_11321,N_10531,N_10770);
nand U11322 (N_11322,N_10378,N_10397);
nand U11323 (N_11323,N_10710,N_10282);
and U11324 (N_11324,N_10444,N_10302);
or U11325 (N_11325,N_10302,N_10579);
xnor U11326 (N_11326,N_10461,N_10495);
nand U11327 (N_11327,N_10707,N_10313);
xnor U11328 (N_11328,N_10529,N_10651);
nor U11329 (N_11329,N_10440,N_10371);
xnor U11330 (N_11330,N_10647,N_10778);
nand U11331 (N_11331,N_10644,N_10226);
and U11332 (N_11332,N_10358,N_10750);
and U11333 (N_11333,N_10730,N_10729);
nor U11334 (N_11334,N_10704,N_10329);
xor U11335 (N_11335,N_10635,N_10461);
nor U11336 (N_11336,N_10572,N_10714);
xor U11337 (N_11337,N_10295,N_10680);
nand U11338 (N_11338,N_10315,N_10472);
or U11339 (N_11339,N_10657,N_10785);
or U11340 (N_11340,N_10288,N_10241);
xor U11341 (N_11341,N_10222,N_10487);
nand U11342 (N_11342,N_10758,N_10689);
and U11343 (N_11343,N_10312,N_10610);
nor U11344 (N_11344,N_10335,N_10276);
or U11345 (N_11345,N_10492,N_10520);
or U11346 (N_11346,N_10229,N_10551);
xor U11347 (N_11347,N_10585,N_10509);
nor U11348 (N_11348,N_10374,N_10630);
and U11349 (N_11349,N_10239,N_10638);
nand U11350 (N_11350,N_10724,N_10277);
and U11351 (N_11351,N_10557,N_10776);
xnor U11352 (N_11352,N_10635,N_10457);
nor U11353 (N_11353,N_10753,N_10388);
nand U11354 (N_11354,N_10795,N_10308);
and U11355 (N_11355,N_10419,N_10374);
nor U11356 (N_11356,N_10640,N_10452);
and U11357 (N_11357,N_10383,N_10355);
xor U11358 (N_11358,N_10501,N_10777);
and U11359 (N_11359,N_10797,N_10447);
nand U11360 (N_11360,N_10566,N_10338);
or U11361 (N_11361,N_10331,N_10243);
nand U11362 (N_11362,N_10627,N_10563);
and U11363 (N_11363,N_10645,N_10596);
nand U11364 (N_11364,N_10653,N_10518);
or U11365 (N_11365,N_10767,N_10324);
nor U11366 (N_11366,N_10521,N_10779);
and U11367 (N_11367,N_10474,N_10418);
nand U11368 (N_11368,N_10272,N_10377);
nor U11369 (N_11369,N_10252,N_10556);
or U11370 (N_11370,N_10400,N_10367);
nor U11371 (N_11371,N_10530,N_10251);
xnor U11372 (N_11372,N_10359,N_10396);
or U11373 (N_11373,N_10692,N_10249);
nand U11374 (N_11374,N_10248,N_10266);
and U11375 (N_11375,N_10794,N_10458);
nor U11376 (N_11376,N_10499,N_10636);
nand U11377 (N_11377,N_10506,N_10336);
or U11378 (N_11378,N_10705,N_10300);
nor U11379 (N_11379,N_10356,N_10576);
and U11380 (N_11380,N_10237,N_10646);
or U11381 (N_11381,N_10425,N_10520);
nor U11382 (N_11382,N_10233,N_10493);
nor U11383 (N_11383,N_10675,N_10295);
and U11384 (N_11384,N_10501,N_10661);
and U11385 (N_11385,N_10486,N_10336);
or U11386 (N_11386,N_10506,N_10700);
xor U11387 (N_11387,N_10253,N_10469);
nor U11388 (N_11388,N_10259,N_10451);
nand U11389 (N_11389,N_10568,N_10665);
nand U11390 (N_11390,N_10255,N_10548);
xor U11391 (N_11391,N_10543,N_10507);
or U11392 (N_11392,N_10381,N_10630);
and U11393 (N_11393,N_10656,N_10751);
and U11394 (N_11394,N_10275,N_10263);
or U11395 (N_11395,N_10215,N_10205);
and U11396 (N_11396,N_10403,N_10704);
nand U11397 (N_11397,N_10492,N_10740);
nor U11398 (N_11398,N_10294,N_10229);
and U11399 (N_11399,N_10773,N_10404);
nand U11400 (N_11400,N_11089,N_11102);
nand U11401 (N_11401,N_10951,N_11210);
xnor U11402 (N_11402,N_10949,N_11318);
and U11403 (N_11403,N_11206,N_11162);
xnor U11404 (N_11404,N_10865,N_10909);
xnor U11405 (N_11405,N_10976,N_11031);
or U11406 (N_11406,N_11025,N_10875);
and U11407 (N_11407,N_10966,N_10916);
or U11408 (N_11408,N_10946,N_11218);
nor U11409 (N_11409,N_11095,N_10867);
nor U11410 (N_11410,N_11118,N_11198);
and U11411 (N_11411,N_11081,N_11141);
or U11412 (N_11412,N_11125,N_11295);
xor U11413 (N_11413,N_11035,N_10806);
and U11414 (N_11414,N_11147,N_11201);
xor U11415 (N_11415,N_11258,N_11010);
nor U11416 (N_11416,N_11268,N_11070);
and U11417 (N_11417,N_10918,N_11055);
xnor U11418 (N_11418,N_11034,N_11378);
xor U11419 (N_11419,N_11273,N_11282);
nand U11420 (N_11420,N_11220,N_10826);
and U11421 (N_11421,N_11324,N_11233);
nor U11422 (N_11422,N_10886,N_11001);
nand U11423 (N_11423,N_11300,N_11367);
xor U11424 (N_11424,N_11397,N_11345);
nand U11425 (N_11425,N_10996,N_11167);
xor U11426 (N_11426,N_11382,N_11006);
and U11427 (N_11427,N_11068,N_10900);
nand U11428 (N_11428,N_11338,N_10919);
xnor U11429 (N_11429,N_10964,N_11003);
xnor U11430 (N_11430,N_10862,N_11110);
or U11431 (N_11431,N_11204,N_11082);
nand U11432 (N_11432,N_11163,N_10864);
nor U11433 (N_11433,N_11079,N_10913);
and U11434 (N_11434,N_11265,N_11049);
and U11435 (N_11435,N_11175,N_11094);
nor U11436 (N_11436,N_11045,N_11359);
nor U11437 (N_11437,N_11191,N_11388);
xor U11438 (N_11438,N_10992,N_10963);
and U11439 (N_11439,N_11289,N_11277);
nor U11440 (N_11440,N_11296,N_11224);
or U11441 (N_11441,N_11309,N_11169);
or U11442 (N_11442,N_10915,N_10857);
nand U11443 (N_11443,N_11390,N_11087);
nand U11444 (N_11444,N_10827,N_10930);
xor U11445 (N_11445,N_10820,N_11287);
nand U11446 (N_11446,N_11337,N_10863);
xor U11447 (N_11447,N_11033,N_11291);
nor U11448 (N_11448,N_11246,N_11393);
nor U11449 (N_11449,N_11336,N_10914);
xnor U11450 (N_11450,N_11263,N_11293);
nand U11451 (N_11451,N_11040,N_11152);
nor U11452 (N_11452,N_11354,N_10835);
nand U11453 (N_11453,N_11202,N_11155);
and U11454 (N_11454,N_11271,N_11389);
nand U11455 (N_11455,N_10877,N_11103);
and U11456 (N_11456,N_11015,N_11348);
and U11457 (N_11457,N_11022,N_10885);
and U11458 (N_11458,N_10809,N_11355);
nand U11459 (N_11459,N_11294,N_10852);
xor U11460 (N_11460,N_11161,N_10961);
nand U11461 (N_11461,N_11126,N_11267);
xnor U11462 (N_11462,N_11283,N_10939);
nand U11463 (N_11463,N_11187,N_11078);
xor U11464 (N_11464,N_11226,N_10831);
xor U11465 (N_11465,N_11330,N_10926);
nand U11466 (N_11466,N_11188,N_11120);
xor U11467 (N_11467,N_11362,N_10829);
nor U11468 (N_11468,N_11060,N_10962);
and U11469 (N_11469,N_11377,N_10837);
and U11470 (N_11470,N_10997,N_11099);
nand U11471 (N_11471,N_11156,N_10944);
xor U11472 (N_11472,N_11140,N_11366);
xor U11473 (N_11473,N_11153,N_11225);
xor U11474 (N_11474,N_11000,N_11379);
nand U11475 (N_11475,N_10948,N_11058);
nand U11476 (N_11476,N_11086,N_10856);
xnor U11477 (N_11477,N_10908,N_11349);
nor U11478 (N_11478,N_11303,N_11384);
nand U11479 (N_11479,N_10878,N_11116);
xor U11480 (N_11480,N_11052,N_11251);
or U11481 (N_11481,N_10813,N_11158);
nor U11482 (N_11482,N_10925,N_10984);
nand U11483 (N_11483,N_11173,N_11036);
nand U11484 (N_11484,N_11215,N_11193);
and U11485 (N_11485,N_11278,N_11091);
and U11486 (N_11486,N_11128,N_11316);
and U11487 (N_11487,N_11012,N_10824);
nor U11488 (N_11488,N_10933,N_11171);
and U11489 (N_11489,N_10975,N_11321);
xor U11490 (N_11490,N_11335,N_10912);
or U11491 (N_11491,N_10884,N_10855);
or U11492 (N_11492,N_11149,N_11160);
and U11493 (N_11493,N_10868,N_11229);
nor U11494 (N_11494,N_10982,N_11257);
xor U11495 (N_11495,N_11264,N_11299);
nor U11496 (N_11496,N_11199,N_10905);
xnor U11497 (N_11497,N_11370,N_10987);
and U11498 (N_11498,N_10986,N_10853);
nand U11499 (N_11499,N_11106,N_10805);
nand U11500 (N_11500,N_10811,N_11298);
or U11501 (N_11501,N_10989,N_10931);
or U11502 (N_11502,N_11333,N_11307);
or U11503 (N_11503,N_11253,N_10812);
or U11504 (N_11504,N_11157,N_11395);
and U11505 (N_11505,N_11067,N_11143);
and U11506 (N_11506,N_11329,N_11088);
xor U11507 (N_11507,N_11242,N_10906);
or U11508 (N_11508,N_10840,N_10881);
xor U11509 (N_11509,N_11097,N_11261);
and U11510 (N_11510,N_11374,N_11028);
and U11511 (N_11511,N_11074,N_10988);
and U11512 (N_11512,N_11044,N_11248);
nor U11513 (N_11513,N_11208,N_11274);
nand U11514 (N_11514,N_11363,N_11130);
xor U11515 (N_11515,N_10947,N_11376);
nor U11516 (N_11516,N_11305,N_11138);
nand U11517 (N_11517,N_10954,N_10817);
or U11518 (N_11518,N_10983,N_11350);
nand U11519 (N_11519,N_11083,N_11260);
xor U11520 (N_11520,N_11018,N_11325);
nor U11521 (N_11521,N_10993,N_11071);
nand U11522 (N_11522,N_10843,N_11178);
and U11523 (N_11523,N_11315,N_10911);
or U11524 (N_11524,N_10956,N_11284);
xor U11525 (N_11525,N_11281,N_11240);
and U11526 (N_11526,N_11117,N_11269);
and U11527 (N_11527,N_10800,N_11219);
nor U11528 (N_11528,N_10816,N_11129);
nor U11529 (N_11529,N_10935,N_10825);
and U11530 (N_11530,N_11230,N_11327);
nand U11531 (N_11531,N_11017,N_10943);
or U11532 (N_11532,N_11174,N_11013);
xnor U11533 (N_11533,N_11019,N_11214);
xnor U11534 (N_11534,N_11054,N_11093);
nor U11535 (N_11535,N_10971,N_11323);
xor U11536 (N_11536,N_11255,N_11047);
and U11537 (N_11537,N_11101,N_10861);
or U11538 (N_11538,N_10883,N_11061);
nand U11539 (N_11539,N_10860,N_10891);
nand U11540 (N_11540,N_10985,N_10953);
nor U11541 (N_11541,N_11286,N_11351);
xor U11542 (N_11542,N_11011,N_11146);
and U11543 (N_11543,N_11008,N_10848);
xor U11544 (N_11544,N_11181,N_10940);
nand U11545 (N_11545,N_10998,N_10854);
nand U11546 (N_11546,N_11150,N_10810);
nand U11547 (N_11547,N_10801,N_11347);
and U11548 (N_11548,N_10836,N_11112);
and U11549 (N_11549,N_11275,N_10960);
or U11550 (N_11550,N_11029,N_11096);
and U11551 (N_11551,N_10942,N_11197);
nand U11552 (N_11552,N_10879,N_11238);
xor U11553 (N_11553,N_10904,N_11084);
nand U11554 (N_11554,N_11236,N_11075);
nor U11555 (N_11555,N_11005,N_10959);
or U11556 (N_11556,N_10974,N_10818);
and U11557 (N_11557,N_11057,N_10934);
nand U11558 (N_11558,N_10957,N_11072);
and U11559 (N_11559,N_10822,N_10873);
nand U11560 (N_11560,N_11334,N_10832);
and U11561 (N_11561,N_10844,N_11109);
or U11562 (N_11562,N_10802,N_10928);
xnor U11563 (N_11563,N_11123,N_11050);
and U11564 (N_11564,N_11203,N_11217);
and U11565 (N_11565,N_11317,N_11342);
xor U11566 (N_11566,N_10950,N_10927);
nor U11567 (N_11567,N_11232,N_10849);
or U11568 (N_11568,N_11166,N_11245);
xor U11569 (N_11569,N_11062,N_11186);
or U11570 (N_11570,N_11032,N_10823);
xnor U11571 (N_11571,N_10907,N_10894);
nor U11572 (N_11572,N_10970,N_10921);
xnor U11573 (N_11573,N_11212,N_11209);
and U11574 (N_11574,N_10924,N_11185);
or U11575 (N_11575,N_11127,N_10977);
or U11576 (N_11576,N_11249,N_11092);
xor U11577 (N_11577,N_10859,N_11319);
and U11578 (N_11578,N_11151,N_11383);
nor U11579 (N_11579,N_11256,N_11159);
or U11580 (N_11580,N_10880,N_11237);
nand U11581 (N_11581,N_11285,N_10808);
nor U11582 (N_11582,N_11252,N_11235);
or U11583 (N_11583,N_11241,N_11373);
or U11584 (N_11584,N_11134,N_11247);
and U11585 (N_11585,N_10902,N_11365);
nor U11586 (N_11586,N_11399,N_11385);
or U11587 (N_11587,N_10819,N_10807);
nand U11588 (N_11588,N_10833,N_10952);
or U11589 (N_11589,N_11310,N_11020);
xor U11590 (N_11590,N_11262,N_11090);
xor U11591 (N_11591,N_11180,N_11254);
or U11592 (N_11592,N_10929,N_11023);
nand U11593 (N_11593,N_10932,N_11014);
xor U11594 (N_11594,N_11165,N_10847);
nor U11595 (N_11595,N_11176,N_11195);
nand U11596 (N_11596,N_11297,N_10999);
and U11597 (N_11597,N_11056,N_11002);
nand U11598 (N_11598,N_10979,N_11392);
nand U11599 (N_11599,N_10972,N_11266);
nor U11600 (N_11600,N_11372,N_11302);
nand U11601 (N_11601,N_10920,N_11039);
nor U11602 (N_11602,N_10839,N_10901);
nand U11603 (N_11603,N_11381,N_11168);
nand U11604 (N_11604,N_10893,N_11007);
and U11605 (N_11605,N_11364,N_11121);
and U11606 (N_11606,N_11085,N_11114);
nand U11607 (N_11607,N_11142,N_11353);
nand U11608 (N_11608,N_11065,N_11053);
nor U11609 (N_11609,N_11113,N_11177);
and U11610 (N_11610,N_11190,N_11250);
xor U11611 (N_11611,N_10981,N_11328);
or U11612 (N_11612,N_11346,N_11243);
nand U11613 (N_11613,N_11205,N_11038);
nor U11614 (N_11614,N_11341,N_11132);
xnor U11615 (N_11615,N_10814,N_11391);
or U11616 (N_11616,N_10828,N_11108);
nor U11617 (N_11617,N_11073,N_11228);
xor U11618 (N_11618,N_11343,N_11396);
xnor U11619 (N_11619,N_11037,N_11292);
or U11620 (N_11620,N_11320,N_11148);
or U11621 (N_11621,N_11344,N_10871);
xnor U11622 (N_11622,N_11306,N_11313);
nand U11623 (N_11623,N_11192,N_11358);
nand U11624 (N_11624,N_10830,N_10973);
and U11625 (N_11625,N_11100,N_10850);
and U11626 (N_11626,N_11222,N_11207);
nor U11627 (N_11627,N_11213,N_11122);
nand U11628 (N_11628,N_11398,N_11137);
xnor U11629 (N_11629,N_11290,N_11308);
and U11630 (N_11630,N_10967,N_11189);
or U11631 (N_11631,N_11144,N_11133);
and U11632 (N_11632,N_10882,N_10841);
and U11633 (N_11633,N_10958,N_11145);
nand U11634 (N_11634,N_11386,N_10910);
and U11635 (N_11635,N_11288,N_10991);
nand U11636 (N_11636,N_11154,N_11164);
and U11637 (N_11637,N_10866,N_11009);
nand U11638 (N_11638,N_10870,N_10874);
nor U11639 (N_11639,N_11024,N_10994);
nand U11640 (N_11640,N_11194,N_11076);
and U11641 (N_11641,N_11200,N_11021);
nor U11642 (N_11642,N_10838,N_10980);
nor U11643 (N_11643,N_10990,N_11360);
and U11644 (N_11644,N_10941,N_10842);
or U11645 (N_11645,N_10834,N_11394);
xnor U11646 (N_11646,N_11311,N_10869);
and U11647 (N_11647,N_11332,N_11059);
xnor U11648 (N_11648,N_11280,N_11041);
and U11649 (N_11649,N_11183,N_10872);
and U11650 (N_11650,N_10804,N_11239);
and U11651 (N_11651,N_11371,N_11276);
nand U11652 (N_11652,N_11098,N_11111);
nand U11653 (N_11653,N_11304,N_11115);
and U11654 (N_11654,N_11211,N_11339);
nor U11655 (N_11655,N_11119,N_11107);
xnor U11656 (N_11656,N_10821,N_10897);
or U11657 (N_11657,N_11124,N_10858);
xor U11658 (N_11658,N_11048,N_10815);
xor U11659 (N_11659,N_11380,N_10845);
or U11660 (N_11660,N_11234,N_10995);
xnor U11661 (N_11661,N_11131,N_10896);
nand U11662 (N_11662,N_10922,N_11004);
nor U11663 (N_11663,N_11135,N_11368);
xnor U11664 (N_11664,N_10846,N_11063);
xnor U11665 (N_11665,N_10936,N_11026);
or U11666 (N_11666,N_10903,N_11027);
xnor U11667 (N_11667,N_11196,N_11069);
nand U11668 (N_11668,N_11080,N_11314);
or U11669 (N_11669,N_10887,N_11182);
or U11670 (N_11670,N_10965,N_11139);
xnor U11671 (N_11671,N_10945,N_10969);
nand U11672 (N_11672,N_11375,N_11301);
and U11673 (N_11673,N_10803,N_10968);
or U11674 (N_11674,N_11357,N_11326);
nand U11675 (N_11675,N_10938,N_11331);
or U11676 (N_11676,N_11270,N_11279);
nor U11677 (N_11677,N_11184,N_10889);
and U11678 (N_11678,N_11042,N_10923);
and U11679 (N_11679,N_11104,N_11172);
nor U11680 (N_11680,N_11030,N_10917);
nor U11681 (N_11681,N_11361,N_10892);
nor U11682 (N_11682,N_11179,N_11227);
and U11683 (N_11683,N_11231,N_11369);
or U11684 (N_11684,N_11016,N_11352);
xnor U11685 (N_11685,N_11312,N_11066);
nand U11686 (N_11686,N_10898,N_11046);
and U11687 (N_11687,N_10888,N_11221);
nor U11688 (N_11688,N_11272,N_11387);
or U11689 (N_11689,N_11064,N_11170);
nor U11690 (N_11690,N_11043,N_10876);
or U11691 (N_11691,N_11259,N_10937);
nor U11692 (N_11692,N_10895,N_11322);
nor U11693 (N_11693,N_11340,N_11077);
and U11694 (N_11694,N_11223,N_11136);
nand U11695 (N_11695,N_11356,N_10978);
or U11696 (N_11696,N_10851,N_10899);
nand U11697 (N_11697,N_11051,N_10955);
or U11698 (N_11698,N_10890,N_11216);
xor U11699 (N_11699,N_11105,N_11244);
nand U11700 (N_11700,N_11318,N_11102);
or U11701 (N_11701,N_10858,N_10913);
or U11702 (N_11702,N_11263,N_10923);
nand U11703 (N_11703,N_11130,N_11061);
or U11704 (N_11704,N_11145,N_11029);
or U11705 (N_11705,N_11220,N_11095);
xnor U11706 (N_11706,N_11059,N_10939);
or U11707 (N_11707,N_11178,N_10851);
nand U11708 (N_11708,N_10821,N_10880);
nand U11709 (N_11709,N_10859,N_11207);
and U11710 (N_11710,N_10862,N_11370);
or U11711 (N_11711,N_11153,N_11169);
nand U11712 (N_11712,N_10980,N_11075);
or U11713 (N_11713,N_11148,N_11274);
xor U11714 (N_11714,N_11163,N_10927);
xor U11715 (N_11715,N_11267,N_10800);
or U11716 (N_11716,N_10913,N_11169);
and U11717 (N_11717,N_10918,N_11172);
nand U11718 (N_11718,N_11157,N_10843);
nand U11719 (N_11719,N_10967,N_10830);
nor U11720 (N_11720,N_11246,N_10990);
nor U11721 (N_11721,N_11126,N_10863);
xor U11722 (N_11722,N_10821,N_11313);
nor U11723 (N_11723,N_11012,N_11354);
xnor U11724 (N_11724,N_11095,N_10840);
nand U11725 (N_11725,N_10868,N_11055);
xor U11726 (N_11726,N_10897,N_10802);
and U11727 (N_11727,N_11327,N_11342);
nor U11728 (N_11728,N_10854,N_11190);
and U11729 (N_11729,N_11250,N_11346);
or U11730 (N_11730,N_11163,N_11014);
nand U11731 (N_11731,N_11029,N_11193);
nor U11732 (N_11732,N_10802,N_11382);
or U11733 (N_11733,N_11192,N_11098);
or U11734 (N_11734,N_10915,N_10822);
nand U11735 (N_11735,N_11281,N_11243);
nand U11736 (N_11736,N_11340,N_10874);
or U11737 (N_11737,N_11000,N_11315);
and U11738 (N_11738,N_11055,N_11052);
nand U11739 (N_11739,N_11273,N_11326);
xnor U11740 (N_11740,N_11363,N_10908);
nor U11741 (N_11741,N_11130,N_10888);
nor U11742 (N_11742,N_11175,N_10889);
xor U11743 (N_11743,N_10920,N_11072);
and U11744 (N_11744,N_11144,N_11082);
nand U11745 (N_11745,N_10951,N_11190);
or U11746 (N_11746,N_11397,N_11074);
nand U11747 (N_11747,N_10925,N_11133);
xor U11748 (N_11748,N_11082,N_10917);
nor U11749 (N_11749,N_10974,N_11107);
nor U11750 (N_11750,N_11357,N_10924);
nand U11751 (N_11751,N_10827,N_11199);
or U11752 (N_11752,N_10934,N_10895);
nor U11753 (N_11753,N_11305,N_11253);
and U11754 (N_11754,N_11159,N_10903);
or U11755 (N_11755,N_11098,N_10912);
or U11756 (N_11756,N_11340,N_11325);
nor U11757 (N_11757,N_11128,N_11371);
or U11758 (N_11758,N_10976,N_10900);
xnor U11759 (N_11759,N_11140,N_11139);
and U11760 (N_11760,N_11279,N_11009);
nand U11761 (N_11761,N_11060,N_11169);
xnor U11762 (N_11762,N_11366,N_11142);
xor U11763 (N_11763,N_10842,N_10806);
nor U11764 (N_11764,N_10966,N_11211);
or U11765 (N_11765,N_11305,N_11042);
nor U11766 (N_11766,N_11066,N_11266);
nand U11767 (N_11767,N_11061,N_11249);
nand U11768 (N_11768,N_11317,N_11389);
nand U11769 (N_11769,N_10903,N_10873);
nor U11770 (N_11770,N_11144,N_11284);
or U11771 (N_11771,N_10941,N_11363);
or U11772 (N_11772,N_11185,N_11075);
nor U11773 (N_11773,N_10990,N_11131);
and U11774 (N_11774,N_10940,N_11316);
xnor U11775 (N_11775,N_11093,N_10892);
nand U11776 (N_11776,N_11307,N_10917);
or U11777 (N_11777,N_11132,N_11304);
or U11778 (N_11778,N_11173,N_11310);
xnor U11779 (N_11779,N_11104,N_10854);
nand U11780 (N_11780,N_11068,N_10925);
nor U11781 (N_11781,N_11027,N_11076);
xor U11782 (N_11782,N_11068,N_10935);
and U11783 (N_11783,N_10808,N_11307);
nand U11784 (N_11784,N_11115,N_10885);
nand U11785 (N_11785,N_11189,N_11245);
and U11786 (N_11786,N_11099,N_11178);
xor U11787 (N_11787,N_11130,N_11086);
nand U11788 (N_11788,N_10860,N_10827);
nand U11789 (N_11789,N_11141,N_10972);
nor U11790 (N_11790,N_10833,N_10962);
nand U11791 (N_11791,N_11097,N_11190);
xnor U11792 (N_11792,N_10870,N_11032);
nor U11793 (N_11793,N_11150,N_10805);
and U11794 (N_11794,N_10945,N_10955);
and U11795 (N_11795,N_11272,N_11083);
and U11796 (N_11796,N_11284,N_10833);
xnor U11797 (N_11797,N_11119,N_10810);
xnor U11798 (N_11798,N_11349,N_10881);
xnor U11799 (N_11799,N_11130,N_11292);
nand U11800 (N_11800,N_10920,N_11190);
nor U11801 (N_11801,N_11363,N_11242);
or U11802 (N_11802,N_11129,N_11063);
or U11803 (N_11803,N_11027,N_10969);
and U11804 (N_11804,N_11244,N_11109);
or U11805 (N_11805,N_11057,N_11302);
or U11806 (N_11806,N_10887,N_11024);
or U11807 (N_11807,N_11030,N_10934);
nor U11808 (N_11808,N_11086,N_10809);
xnor U11809 (N_11809,N_11135,N_11286);
or U11810 (N_11810,N_11386,N_11180);
nand U11811 (N_11811,N_11056,N_10804);
nor U11812 (N_11812,N_11367,N_10938);
nor U11813 (N_11813,N_11033,N_10931);
nand U11814 (N_11814,N_11243,N_11123);
xnor U11815 (N_11815,N_11049,N_11123);
xnor U11816 (N_11816,N_10939,N_11312);
nor U11817 (N_11817,N_11309,N_11024);
or U11818 (N_11818,N_11308,N_10862);
nand U11819 (N_11819,N_10885,N_11178);
or U11820 (N_11820,N_11045,N_11054);
nand U11821 (N_11821,N_11248,N_10854);
or U11822 (N_11822,N_11354,N_11043);
and U11823 (N_11823,N_11349,N_10977);
and U11824 (N_11824,N_11385,N_10810);
or U11825 (N_11825,N_11043,N_11149);
or U11826 (N_11826,N_11360,N_10827);
nand U11827 (N_11827,N_11127,N_11065);
and U11828 (N_11828,N_11292,N_10889);
xnor U11829 (N_11829,N_11168,N_10893);
nand U11830 (N_11830,N_10931,N_11169);
or U11831 (N_11831,N_11300,N_10852);
xnor U11832 (N_11832,N_10836,N_11370);
or U11833 (N_11833,N_11163,N_10938);
and U11834 (N_11834,N_11175,N_10933);
nand U11835 (N_11835,N_10888,N_10890);
xnor U11836 (N_11836,N_11052,N_11116);
or U11837 (N_11837,N_11084,N_10864);
nor U11838 (N_11838,N_10854,N_11090);
or U11839 (N_11839,N_11235,N_11292);
or U11840 (N_11840,N_10917,N_10934);
nand U11841 (N_11841,N_11106,N_11394);
and U11842 (N_11842,N_10951,N_11021);
xor U11843 (N_11843,N_11244,N_11287);
and U11844 (N_11844,N_10949,N_10948);
nand U11845 (N_11845,N_11178,N_10989);
nor U11846 (N_11846,N_11022,N_11236);
xnor U11847 (N_11847,N_11129,N_11216);
nand U11848 (N_11848,N_11000,N_10929);
nor U11849 (N_11849,N_11295,N_10987);
or U11850 (N_11850,N_11003,N_11270);
xnor U11851 (N_11851,N_11356,N_11164);
nor U11852 (N_11852,N_11141,N_11316);
xnor U11853 (N_11853,N_10820,N_11125);
nand U11854 (N_11854,N_10818,N_10840);
nor U11855 (N_11855,N_11238,N_11107);
xnor U11856 (N_11856,N_11187,N_11006);
or U11857 (N_11857,N_11391,N_11267);
nand U11858 (N_11858,N_11323,N_11190);
xnor U11859 (N_11859,N_11231,N_11348);
nor U11860 (N_11860,N_11094,N_11039);
xor U11861 (N_11861,N_10935,N_10947);
nor U11862 (N_11862,N_11202,N_11102);
or U11863 (N_11863,N_10938,N_11144);
and U11864 (N_11864,N_11216,N_11092);
or U11865 (N_11865,N_11050,N_11297);
and U11866 (N_11866,N_11279,N_11269);
or U11867 (N_11867,N_11084,N_10806);
nand U11868 (N_11868,N_11075,N_11338);
nor U11869 (N_11869,N_11003,N_11240);
xnor U11870 (N_11870,N_11084,N_11279);
nor U11871 (N_11871,N_10909,N_11011);
or U11872 (N_11872,N_10876,N_11325);
and U11873 (N_11873,N_11151,N_10834);
nor U11874 (N_11874,N_11398,N_11028);
xnor U11875 (N_11875,N_11311,N_11035);
nand U11876 (N_11876,N_10873,N_11053);
or U11877 (N_11877,N_11016,N_11103);
xnor U11878 (N_11878,N_11069,N_11355);
or U11879 (N_11879,N_11350,N_10995);
xor U11880 (N_11880,N_11246,N_10802);
xor U11881 (N_11881,N_11124,N_10959);
xnor U11882 (N_11882,N_11186,N_11277);
xor U11883 (N_11883,N_11311,N_10966);
nor U11884 (N_11884,N_11070,N_11396);
nor U11885 (N_11885,N_11116,N_11130);
xor U11886 (N_11886,N_11311,N_10912);
and U11887 (N_11887,N_11239,N_11228);
nor U11888 (N_11888,N_11033,N_11055);
xnor U11889 (N_11889,N_11193,N_11083);
xnor U11890 (N_11890,N_11304,N_10845);
or U11891 (N_11891,N_11029,N_10857);
and U11892 (N_11892,N_10862,N_11368);
nor U11893 (N_11893,N_11185,N_10925);
nand U11894 (N_11894,N_11147,N_11111);
and U11895 (N_11895,N_11137,N_10851);
or U11896 (N_11896,N_11224,N_11076);
and U11897 (N_11897,N_11166,N_10977);
xnor U11898 (N_11898,N_11361,N_10810);
nand U11899 (N_11899,N_11170,N_11229);
nand U11900 (N_11900,N_11357,N_11338);
and U11901 (N_11901,N_10989,N_10958);
xor U11902 (N_11902,N_11376,N_10983);
and U11903 (N_11903,N_11010,N_11084);
or U11904 (N_11904,N_10926,N_11024);
or U11905 (N_11905,N_11303,N_10938);
or U11906 (N_11906,N_11251,N_11381);
nor U11907 (N_11907,N_11168,N_11215);
and U11908 (N_11908,N_11010,N_10889);
xnor U11909 (N_11909,N_11067,N_10996);
nand U11910 (N_11910,N_11118,N_11390);
xor U11911 (N_11911,N_11378,N_10836);
xnor U11912 (N_11912,N_10995,N_11386);
xor U11913 (N_11913,N_10955,N_10939);
nor U11914 (N_11914,N_10926,N_11044);
nor U11915 (N_11915,N_11098,N_11213);
nand U11916 (N_11916,N_10941,N_11045);
nor U11917 (N_11917,N_11221,N_11309);
nand U11918 (N_11918,N_10817,N_10854);
or U11919 (N_11919,N_10985,N_11057);
and U11920 (N_11920,N_11290,N_11345);
xor U11921 (N_11921,N_11271,N_11125);
or U11922 (N_11922,N_11393,N_10997);
or U11923 (N_11923,N_11015,N_11165);
nand U11924 (N_11924,N_10869,N_11295);
and U11925 (N_11925,N_10916,N_10913);
or U11926 (N_11926,N_11371,N_11296);
nor U11927 (N_11927,N_10925,N_10811);
and U11928 (N_11928,N_11038,N_11270);
and U11929 (N_11929,N_10850,N_10956);
nor U11930 (N_11930,N_10857,N_10878);
and U11931 (N_11931,N_11085,N_11097);
nand U11932 (N_11932,N_11128,N_11132);
nand U11933 (N_11933,N_10974,N_11036);
xor U11934 (N_11934,N_10930,N_10990);
nor U11935 (N_11935,N_11073,N_11315);
and U11936 (N_11936,N_11054,N_10924);
nand U11937 (N_11937,N_11084,N_10885);
or U11938 (N_11938,N_11283,N_11252);
xnor U11939 (N_11939,N_11326,N_10956);
or U11940 (N_11940,N_10807,N_11238);
or U11941 (N_11941,N_11220,N_11122);
xnor U11942 (N_11942,N_11315,N_11257);
xor U11943 (N_11943,N_11254,N_11139);
or U11944 (N_11944,N_11189,N_11341);
and U11945 (N_11945,N_11132,N_10831);
and U11946 (N_11946,N_11099,N_10817);
nor U11947 (N_11947,N_11194,N_11059);
nand U11948 (N_11948,N_11043,N_11355);
xnor U11949 (N_11949,N_10970,N_11130);
and U11950 (N_11950,N_11051,N_11242);
nor U11951 (N_11951,N_11395,N_10809);
or U11952 (N_11952,N_11089,N_10997);
nor U11953 (N_11953,N_11180,N_10820);
nor U11954 (N_11954,N_11384,N_10892);
xor U11955 (N_11955,N_11136,N_11159);
and U11956 (N_11956,N_10977,N_11297);
or U11957 (N_11957,N_11284,N_11058);
and U11958 (N_11958,N_11234,N_11312);
and U11959 (N_11959,N_11125,N_11006);
or U11960 (N_11960,N_10994,N_10803);
nand U11961 (N_11961,N_11039,N_10806);
and U11962 (N_11962,N_10967,N_11392);
nor U11963 (N_11963,N_10930,N_11191);
and U11964 (N_11964,N_11159,N_11247);
xor U11965 (N_11965,N_11260,N_11108);
nand U11966 (N_11966,N_10848,N_11332);
or U11967 (N_11967,N_11263,N_11371);
nor U11968 (N_11968,N_11107,N_10905);
nor U11969 (N_11969,N_11242,N_11180);
or U11970 (N_11970,N_11119,N_11165);
and U11971 (N_11971,N_11078,N_11339);
nand U11972 (N_11972,N_11381,N_11063);
nand U11973 (N_11973,N_10892,N_10959);
nor U11974 (N_11974,N_10981,N_11253);
and U11975 (N_11975,N_11052,N_11111);
nor U11976 (N_11976,N_11038,N_11219);
xor U11977 (N_11977,N_11177,N_10847);
and U11978 (N_11978,N_11019,N_11095);
and U11979 (N_11979,N_10883,N_10961);
nor U11980 (N_11980,N_11273,N_11209);
nand U11981 (N_11981,N_10909,N_10829);
or U11982 (N_11982,N_11160,N_11069);
or U11983 (N_11983,N_11131,N_11098);
xor U11984 (N_11984,N_10989,N_10917);
nor U11985 (N_11985,N_11029,N_10995);
nor U11986 (N_11986,N_11026,N_10967);
nor U11987 (N_11987,N_10891,N_10975);
or U11988 (N_11988,N_11184,N_11004);
and U11989 (N_11989,N_11322,N_11251);
nor U11990 (N_11990,N_11145,N_10876);
xnor U11991 (N_11991,N_11323,N_10867);
or U11992 (N_11992,N_11326,N_11032);
nand U11993 (N_11993,N_11191,N_11021);
nand U11994 (N_11994,N_10919,N_11327);
nor U11995 (N_11995,N_10836,N_11033);
or U11996 (N_11996,N_11340,N_10968);
nor U11997 (N_11997,N_11141,N_11088);
and U11998 (N_11998,N_10908,N_10824);
nor U11999 (N_11999,N_11005,N_10963);
xor U12000 (N_12000,N_11964,N_11679);
xor U12001 (N_12001,N_11888,N_11510);
xnor U12002 (N_12002,N_11752,N_11419);
nor U12003 (N_12003,N_11639,N_11803);
or U12004 (N_12004,N_11598,N_11766);
and U12005 (N_12005,N_11885,N_11946);
nand U12006 (N_12006,N_11859,N_11996);
nand U12007 (N_12007,N_11978,N_11729);
and U12008 (N_12008,N_11967,N_11809);
nand U12009 (N_12009,N_11602,N_11477);
nand U12010 (N_12010,N_11654,N_11658);
and U12011 (N_12011,N_11599,N_11693);
xor U12012 (N_12012,N_11895,N_11966);
xor U12013 (N_12013,N_11512,N_11673);
xnor U12014 (N_12014,N_11807,N_11619);
xnor U12015 (N_12015,N_11539,N_11605);
nand U12016 (N_12016,N_11706,N_11798);
or U12017 (N_12017,N_11681,N_11454);
or U12018 (N_12018,N_11561,N_11692);
xor U12019 (N_12019,N_11969,N_11956);
xnor U12020 (N_12020,N_11879,N_11995);
nor U12021 (N_12021,N_11558,N_11814);
or U12022 (N_12022,N_11850,N_11436);
or U12023 (N_12023,N_11636,N_11970);
nand U12024 (N_12024,N_11638,N_11427);
xnor U12025 (N_12025,N_11723,N_11755);
nor U12026 (N_12026,N_11630,N_11670);
xnor U12027 (N_12027,N_11715,N_11853);
xor U12028 (N_12028,N_11551,N_11781);
xor U12029 (N_12029,N_11604,N_11981);
nand U12030 (N_12030,N_11666,N_11833);
or U12031 (N_12031,N_11898,N_11515);
and U12032 (N_12032,N_11963,N_11446);
nand U12033 (N_12033,N_11408,N_11851);
xor U12034 (N_12034,N_11533,N_11699);
nand U12035 (N_12035,N_11453,N_11908);
nor U12036 (N_12036,N_11431,N_11503);
or U12037 (N_12037,N_11549,N_11911);
nand U12038 (N_12038,N_11507,N_11548);
and U12039 (N_12039,N_11501,N_11663);
or U12040 (N_12040,N_11499,N_11938);
xnor U12041 (N_12041,N_11661,N_11952);
nor U12042 (N_12042,N_11754,N_11472);
xor U12043 (N_12043,N_11433,N_11674);
and U12044 (N_12044,N_11724,N_11883);
nand U12045 (N_12045,N_11659,N_11535);
nand U12046 (N_12046,N_11768,N_11793);
nor U12047 (N_12047,N_11517,N_11703);
nand U12048 (N_12048,N_11606,N_11450);
nand U12049 (N_12049,N_11442,N_11465);
nand U12050 (N_12050,N_11451,N_11610);
or U12051 (N_12051,N_11702,N_11652);
nor U12052 (N_12052,N_11439,N_11470);
nor U12053 (N_12053,N_11444,N_11878);
xnor U12054 (N_12054,N_11756,N_11530);
xor U12055 (N_12055,N_11521,N_11730);
and U12056 (N_12056,N_11601,N_11954);
xnor U12057 (N_12057,N_11513,N_11740);
nor U12058 (N_12058,N_11986,N_11993);
nand U12059 (N_12059,N_11965,N_11891);
nor U12060 (N_12060,N_11957,N_11790);
and U12061 (N_12061,N_11866,N_11443);
xnor U12062 (N_12062,N_11989,N_11417);
and U12063 (N_12063,N_11595,N_11627);
or U12064 (N_12064,N_11900,N_11626);
and U12065 (N_12065,N_11894,N_11678);
nand U12066 (N_12066,N_11422,N_11532);
nand U12067 (N_12067,N_11929,N_11916);
xnor U12068 (N_12068,N_11893,N_11460);
or U12069 (N_12069,N_11493,N_11880);
nand U12070 (N_12070,N_11941,N_11557);
or U12071 (N_12071,N_11823,N_11409);
and U12072 (N_12072,N_11990,N_11924);
xnor U12073 (N_12073,N_11852,N_11538);
or U12074 (N_12074,N_11700,N_11556);
and U12075 (N_12075,N_11907,N_11788);
xor U12076 (N_12076,N_11482,N_11719);
or U12077 (N_12077,N_11633,N_11994);
nand U12078 (N_12078,N_11708,N_11704);
and U12079 (N_12079,N_11922,N_11779);
xor U12080 (N_12080,N_11890,N_11757);
xnor U12081 (N_12081,N_11920,N_11608);
or U12082 (N_12082,N_11865,N_11410);
nand U12083 (N_12083,N_11589,N_11563);
or U12084 (N_12084,N_11497,N_11792);
or U12085 (N_12085,N_11484,N_11928);
or U12086 (N_12086,N_11874,N_11435);
nor U12087 (N_12087,N_11985,N_11582);
or U12088 (N_12088,N_11694,N_11821);
nor U12089 (N_12089,N_11889,N_11615);
nand U12090 (N_12090,N_11849,N_11411);
or U12091 (N_12091,N_11457,N_11945);
and U12092 (N_12092,N_11747,N_11571);
or U12093 (N_12093,N_11437,N_11463);
and U12094 (N_12094,N_11816,N_11618);
and U12095 (N_12095,N_11919,N_11725);
xnor U12096 (N_12096,N_11732,N_11867);
and U12097 (N_12097,N_11820,N_11488);
and U12098 (N_12098,N_11675,N_11910);
xnor U12099 (N_12099,N_11462,N_11544);
nor U12100 (N_12100,N_11759,N_11461);
or U12101 (N_12101,N_11817,N_11741);
nor U12102 (N_12102,N_11742,N_11855);
xnor U12103 (N_12103,N_11944,N_11511);
and U12104 (N_12104,N_11813,N_11498);
nor U12105 (N_12105,N_11677,N_11858);
or U12106 (N_12106,N_11690,N_11974);
nor U12107 (N_12107,N_11592,N_11429);
and U12108 (N_12108,N_11651,N_11543);
and U12109 (N_12109,N_11918,N_11418);
or U12110 (N_12110,N_11585,N_11887);
and U12111 (N_12111,N_11426,N_11791);
nand U12112 (N_12112,N_11689,N_11844);
xnor U12113 (N_12113,N_11830,N_11467);
or U12114 (N_12114,N_11466,N_11913);
and U12115 (N_12115,N_11886,N_11490);
and U12116 (N_12116,N_11516,N_11770);
xnor U12117 (N_12117,N_11537,N_11669);
xor U12118 (N_12118,N_11728,N_11933);
nand U12119 (N_12119,N_11400,N_11837);
nand U12120 (N_12120,N_11458,N_11709);
nand U12121 (N_12121,N_11713,N_11802);
nor U12122 (N_12122,N_11485,N_11459);
or U12123 (N_12123,N_11877,N_11831);
and U12124 (N_12124,N_11832,N_11936);
xor U12125 (N_12125,N_11575,N_11438);
and U12126 (N_12126,N_11940,N_11523);
nor U12127 (N_12127,N_11785,N_11800);
nand U12128 (N_12128,N_11407,N_11553);
or U12129 (N_12129,N_11518,N_11761);
xnor U12130 (N_12130,N_11819,N_11641);
or U12131 (N_12131,N_11780,N_11600);
and U12132 (N_12132,N_11483,N_11705);
nand U12133 (N_12133,N_11491,N_11420);
nand U12134 (N_12134,N_11687,N_11495);
nand U12135 (N_12135,N_11447,N_11711);
or U12136 (N_12136,N_11672,N_11617);
nand U12137 (N_12137,N_11810,N_11801);
and U12138 (N_12138,N_11881,N_11455);
nor U12139 (N_12139,N_11547,N_11577);
nand U12140 (N_12140,N_11991,N_11736);
xnor U12141 (N_12141,N_11710,N_11901);
or U12142 (N_12142,N_11988,N_11869);
xor U12143 (N_12143,N_11489,N_11951);
nor U12144 (N_12144,N_11861,N_11603);
or U12145 (N_12145,N_11947,N_11842);
nand U12146 (N_12146,N_11960,N_11469);
or U12147 (N_12147,N_11856,N_11860);
or U12148 (N_12148,N_11441,N_11931);
and U12149 (N_12149,N_11829,N_11591);
and U12150 (N_12150,N_11424,N_11581);
or U12151 (N_12151,N_11587,N_11906);
or U12152 (N_12152,N_11789,N_11475);
and U12153 (N_12153,N_11746,N_11722);
and U12154 (N_12154,N_11769,N_11733);
xor U12155 (N_12155,N_11653,N_11403);
and U12156 (N_12156,N_11632,N_11806);
nor U12157 (N_12157,N_11644,N_11767);
and U12158 (N_12158,N_11734,N_11784);
and U12159 (N_12159,N_11502,N_11686);
nand U12160 (N_12160,N_11479,N_11868);
nor U12161 (N_12161,N_11846,N_11540);
xor U12162 (N_12162,N_11811,N_11760);
xnor U12163 (N_12163,N_11872,N_11775);
and U12164 (N_12164,N_11440,N_11508);
or U12165 (N_12165,N_11925,N_11930);
nand U12166 (N_12166,N_11721,N_11808);
xor U12167 (N_12167,N_11795,N_11764);
and U12168 (N_12168,N_11487,N_11468);
or U12169 (N_12169,N_11425,N_11959);
or U12170 (N_12170,N_11701,N_11423);
and U12171 (N_12171,N_11797,N_11642);
xnor U12172 (N_12172,N_11939,N_11805);
xnor U12173 (N_12173,N_11902,N_11528);
and U12174 (N_12174,N_11613,N_11737);
or U12175 (N_12175,N_11696,N_11594);
xor U12176 (N_12176,N_11452,N_11405);
and U12177 (N_12177,N_11862,N_11771);
nor U12178 (N_12178,N_11683,N_11609);
nor U12179 (N_12179,N_11682,N_11648);
and U12180 (N_12180,N_11876,N_11979);
nor U12181 (N_12181,N_11778,N_11905);
or U12182 (N_12182,N_11597,N_11656);
xor U12183 (N_12183,N_11949,N_11854);
or U12184 (N_12184,N_11564,N_11509);
nor U12185 (N_12185,N_11568,N_11909);
and U12186 (N_12186,N_11912,N_11815);
nand U12187 (N_12187,N_11657,N_11845);
xor U12188 (N_12188,N_11720,N_11695);
and U12189 (N_12189,N_11735,N_11524);
and U12190 (N_12190,N_11456,N_11975);
nand U12191 (N_12191,N_11545,N_11496);
nor U12192 (N_12192,N_11635,N_11968);
nor U12193 (N_12193,N_11492,N_11932);
nor U12194 (N_12194,N_11934,N_11588);
and U12195 (N_12195,N_11473,N_11903);
xnor U12196 (N_12196,N_11818,N_11471);
or U12197 (N_12197,N_11526,N_11566);
xor U12198 (N_12198,N_11958,N_11825);
nand U12199 (N_12199,N_11448,N_11999);
and U12200 (N_12200,N_11474,N_11998);
nand U12201 (N_12201,N_11796,N_11971);
or U12202 (N_12202,N_11923,N_11662);
xor U12203 (N_12203,N_11536,N_11621);
nand U12204 (N_12204,N_11576,N_11973);
and U12205 (N_12205,N_11584,N_11804);
xnor U12206 (N_12206,N_11643,N_11667);
nand U12207 (N_12207,N_11717,N_11750);
nor U12208 (N_12208,N_11840,N_11432);
or U12209 (N_12209,N_11915,N_11743);
nand U12210 (N_12210,N_11664,N_11712);
nand U12211 (N_12211,N_11421,N_11622);
or U12212 (N_12212,N_11783,N_11841);
and U12213 (N_12213,N_11870,N_11892);
xnor U12214 (N_12214,N_11884,N_11406);
and U12215 (N_12215,N_11625,N_11727);
nor U12216 (N_12216,N_11647,N_11554);
or U12217 (N_12217,N_11917,N_11478);
nand U12218 (N_12218,N_11772,N_11763);
nor U12219 (N_12219,N_11623,N_11765);
and U12220 (N_12220,N_11871,N_11476);
and U12221 (N_12221,N_11749,N_11449);
and U12222 (N_12222,N_11751,N_11745);
xnor U12223 (N_12223,N_11646,N_11718);
nor U12224 (N_12224,N_11620,N_11977);
and U12225 (N_12225,N_11527,N_11707);
and U12226 (N_12226,N_11583,N_11612);
or U12227 (N_12227,N_11428,N_11731);
and U12228 (N_12228,N_11776,N_11739);
nand U12229 (N_12229,N_11836,N_11787);
or U12230 (N_12230,N_11607,N_11640);
or U12231 (N_12231,N_11481,N_11414);
nand U12232 (N_12232,N_11777,N_11572);
nand U12233 (N_12233,N_11586,N_11982);
nor U12234 (N_12234,N_11569,N_11857);
or U12235 (N_12235,N_11637,N_11698);
or U12236 (N_12236,N_11688,N_11774);
xnor U12237 (N_12237,N_11826,N_11504);
or U12238 (N_12238,N_11786,N_11943);
xor U12239 (N_12239,N_11559,N_11691);
and U12240 (N_12240,N_11838,N_11983);
nor U12241 (N_12241,N_11697,N_11505);
or U12242 (N_12242,N_11794,N_11834);
and U12243 (N_12243,N_11843,N_11955);
and U12244 (N_12244,N_11645,N_11748);
or U12245 (N_12245,N_11997,N_11629);
or U12246 (N_12246,N_11628,N_11534);
xnor U12247 (N_12247,N_11514,N_11671);
xor U12248 (N_12248,N_11828,N_11542);
and U12249 (N_12249,N_11914,N_11839);
and U12250 (N_12250,N_11744,N_11953);
nand U12251 (N_12251,N_11948,N_11896);
or U12252 (N_12252,N_11579,N_11402);
and U12253 (N_12253,N_11873,N_11899);
xor U12254 (N_12254,N_11655,N_11950);
and U12255 (N_12255,N_11555,N_11416);
xor U12256 (N_12256,N_11520,N_11897);
nand U12257 (N_12257,N_11992,N_11684);
xor U12258 (N_12258,N_11773,N_11624);
nand U12259 (N_12259,N_11616,N_11926);
nand U12260 (N_12260,N_11570,N_11961);
nor U12261 (N_12261,N_11593,N_11714);
or U12262 (N_12262,N_11590,N_11580);
nand U12263 (N_12263,N_11987,N_11882);
xnor U12264 (N_12264,N_11976,N_11480);
nand U12265 (N_12265,N_11634,N_11812);
and U12266 (N_12266,N_11578,N_11753);
xor U12267 (N_12267,N_11413,N_11412);
and U12268 (N_12268,N_11762,N_11430);
nand U12269 (N_12269,N_11847,N_11676);
xnor U12270 (N_12270,N_11782,N_11935);
nor U12271 (N_12271,N_11921,N_11962);
xnor U12272 (N_12272,N_11552,N_11614);
xor U12273 (N_12273,N_11500,N_11863);
nor U12274 (N_12274,N_11560,N_11550);
or U12275 (N_12275,N_11529,N_11927);
nand U12276 (N_12276,N_11680,N_11401);
nor U12277 (N_12277,N_11665,N_11631);
nor U12278 (N_12278,N_11486,N_11726);
xor U12279 (N_12279,N_11685,N_11522);
nand U12280 (N_12280,N_11660,N_11596);
and U12281 (N_12281,N_11415,N_11464);
nand U12282 (N_12282,N_11835,N_11531);
and U12283 (N_12283,N_11404,N_11758);
xnor U12284 (N_12284,N_11567,N_11525);
nor U12285 (N_12285,N_11562,N_11980);
xor U12286 (N_12286,N_11848,N_11864);
or U12287 (N_12287,N_11565,N_11904);
xor U12288 (N_12288,N_11445,N_11824);
or U12289 (N_12289,N_11984,N_11434);
and U12290 (N_12290,N_11822,N_11506);
xnor U12291 (N_12291,N_11494,N_11972);
or U12292 (N_12292,N_11942,N_11668);
or U12293 (N_12293,N_11573,N_11519);
xnor U12294 (N_12294,N_11827,N_11650);
or U12295 (N_12295,N_11716,N_11649);
nand U12296 (N_12296,N_11611,N_11574);
nand U12297 (N_12297,N_11875,N_11738);
or U12298 (N_12298,N_11799,N_11541);
xor U12299 (N_12299,N_11546,N_11937);
nor U12300 (N_12300,N_11889,N_11964);
nand U12301 (N_12301,N_11742,N_11751);
nand U12302 (N_12302,N_11504,N_11694);
nor U12303 (N_12303,N_11840,N_11959);
nand U12304 (N_12304,N_11711,N_11886);
and U12305 (N_12305,N_11917,N_11774);
nor U12306 (N_12306,N_11838,N_11440);
nor U12307 (N_12307,N_11690,N_11831);
and U12308 (N_12308,N_11619,N_11892);
nor U12309 (N_12309,N_11779,N_11660);
nand U12310 (N_12310,N_11840,N_11543);
or U12311 (N_12311,N_11483,N_11509);
xnor U12312 (N_12312,N_11536,N_11910);
nor U12313 (N_12313,N_11899,N_11672);
nand U12314 (N_12314,N_11846,N_11828);
nand U12315 (N_12315,N_11560,N_11477);
or U12316 (N_12316,N_11779,N_11993);
nand U12317 (N_12317,N_11560,N_11885);
and U12318 (N_12318,N_11561,N_11432);
xor U12319 (N_12319,N_11705,N_11710);
xor U12320 (N_12320,N_11440,N_11876);
and U12321 (N_12321,N_11569,N_11683);
nand U12322 (N_12322,N_11985,N_11798);
and U12323 (N_12323,N_11732,N_11642);
nand U12324 (N_12324,N_11592,N_11625);
or U12325 (N_12325,N_11564,N_11664);
nor U12326 (N_12326,N_11861,N_11986);
or U12327 (N_12327,N_11658,N_11557);
and U12328 (N_12328,N_11934,N_11514);
nor U12329 (N_12329,N_11677,N_11745);
nand U12330 (N_12330,N_11921,N_11619);
nand U12331 (N_12331,N_11995,N_11809);
nand U12332 (N_12332,N_11638,N_11729);
nor U12333 (N_12333,N_11755,N_11987);
or U12334 (N_12334,N_11630,N_11435);
xor U12335 (N_12335,N_11585,N_11704);
and U12336 (N_12336,N_11504,N_11788);
and U12337 (N_12337,N_11748,N_11447);
nand U12338 (N_12338,N_11947,N_11794);
or U12339 (N_12339,N_11574,N_11610);
nand U12340 (N_12340,N_11761,N_11844);
xnor U12341 (N_12341,N_11997,N_11673);
nand U12342 (N_12342,N_11483,N_11809);
and U12343 (N_12343,N_11407,N_11902);
xor U12344 (N_12344,N_11883,N_11537);
nand U12345 (N_12345,N_11485,N_11422);
or U12346 (N_12346,N_11625,N_11885);
nand U12347 (N_12347,N_11668,N_11426);
xor U12348 (N_12348,N_11793,N_11817);
nand U12349 (N_12349,N_11664,N_11863);
xor U12350 (N_12350,N_11602,N_11619);
nand U12351 (N_12351,N_11772,N_11724);
nor U12352 (N_12352,N_11976,N_11686);
xor U12353 (N_12353,N_11701,N_11457);
nand U12354 (N_12354,N_11606,N_11593);
or U12355 (N_12355,N_11533,N_11733);
nor U12356 (N_12356,N_11621,N_11711);
nand U12357 (N_12357,N_11764,N_11975);
nand U12358 (N_12358,N_11446,N_11876);
nor U12359 (N_12359,N_11916,N_11652);
and U12360 (N_12360,N_11741,N_11625);
xnor U12361 (N_12361,N_11800,N_11781);
xnor U12362 (N_12362,N_11521,N_11735);
nor U12363 (N_12363,N_11757,N_11873);
nor U12364 (N_12364,N_11844,N_11497);
or U12365 (N_12365,N_11566,N_11459);
and U12366 (N_12366,N_11434,N_11765);
and U12367 (N_12367,N_11985,N_11859);
nand U12368 (N_12368,N_11475,N_11958);
xor U12369 (N_12369,N_11914,N_11945);
and U12370 (N_12370,N_11922,N_11830);
or U12371 (N_12371,N_11553,N_11878);
xnor U12372 (N_12372,N_11830,N_11663);
nand U12373 (N_12373,N_11990,N_11684);
nor U12374 (N_12374,N_11614,N_11636);
nand U12375 (N_12375,N_11879,N_11878);
nand U12376 (N_12376,N_11553,N_11921);
nand U12377 (N_12377,N_11890,N_11650);
xor U12378 (N_12378,N_11639,N_11600);
nor U12379 (N_12379,N_11928,N_11764);
or U12380 (N_12380,N_11680,N_11738);
nand U12381 (N_12381,N_11576,N_11916);
xor U12382 (N_12382,N_11949,N_11425);
nand U12383 (N_12383,N_11948,N_11955);
nor U12384 (N_12384,N_11655,N_11986);
nand U12385 (N_12385,N_11806,N_11986);
or U12386 (N_12386,N_11829,N_11710);
and U12387 (N_12387,N_11838,N_11575);
or U12388 (N_12388,N_11709,N_11794);
or U12389 (N_12389,N_11670,N_11826);
xnor U12390 (N_12390,N_11972,N_11843);
nor U12391 (N_12391,N_11603,N_11767);
nand U12392 (N_12392,N_11642,N_11490);
xor U12393 (N_12393,N_11705,N_11753);
and U12394 (N_12394,N_11929,N_11977);
nor U12395 (N_12395,N_11627,N_11490);
xor U12396 (N_12396,N_11603,N_11402);
and U12397 (N_12397,N_11462,N_11618);
nor U12398 (N_12398,N_11991,N_11458);
and U12399 (N_12399,N_11750,N_11856);
or U12400 (N_12400,N_11401,N_11443);
and U12401 (N_12401,N_11788,N_11600);
nor U12402 (N_12402,N_11400,N_11621);
and U12403 (N_12403,N_11462,N_11759);
xor U12404 (N_12404,N_11429,N_11499);
nand U12405 (N_12405,N_11686,N_11437);
nor U12406 (N_12406,N_11707,N_11993);
nor U12407 (N_12407,N_11569,N_11696);
nor U12408 (N_12408,N_11412,N_11932);
or U12409 (N_12409,N_11678,N_11895);
xor U12410 (N_12410,N_11487,N_11593);
nand U12411 (N_12411,N_11656,N_11802);
nand U12412 (N_12412,N_11522,N_11950);
or U12413 (N_12413,N_11740,N_11730);
or U12414 (N_12414,N_11938,N_11780);
or U12415 (N_12415,N_11631,N_11598);
xnor U12416 (N_12416,N_11691,N_11839);
or U12417 (N_12417,N_11841,N_11636);
or U12418 (N_12418,N_11890,N_11473);
and U12419 (N_12419,N_11590,N_11780);
nor U12420 (N_12420,N_11403,N_11936);
or U12421 (N_12421,N_11725,N_11975);
and U12422 (N_12422,N_11524,N_11788);
xor U12423 (N_12423,N_11995,N_11403);
and U12424 (N_12424,N_11531,N_11903);
and U12425 (N_12425,N_11607,N_11545);
xnor U12426 (N_12426,N_11925,N_11516);
and U12427 (N_12427,N_11716,N_11947);
nor U12428 (N_12428,N_11778,N_11801);
nor U12429 (N_12429,N_11810,N_11506);
or U12430 (N_12430,N_11951,N_11593);
xnor U12431 (N_12431,N_11801,N_11643);
xnor U12432 (N_12432,N_11625,N_11980);
xnor U12433 (N_12433,N_11407,N_11601);
or U12434 (N_12434,N_11609,N_11867);
or U12435 (N_12435,N_11451,N_11449);
nand U12436 (N_12436,N_11528,N_11411);
nand U12437 (N_12437,N_11573,N_11522);
and U12438 (N_12438,N_11849,N_11520);
nor U12439 (N_12439,N_11555,N_11961);
nand U12440 (N_12440,N_11453,N_11917);
nand U12441 (N_12441,N_11966,N_11739);
or U12442 (N_12442,N_11584,N_11799);
nor U12443 (N_12443,N_11636,N_11671);
xnor U12444 (N_12444,N_11787,N_11862);
and U12445 (N_12445,N_11442,N_11825);
nand U12446 (N_12446,N_11585,N_11506);
xnor U12447 (N_12447,N_11659,N_11409);
nand U12448 (N_12448,N_11850,N_11456);
xor U12449 (N_12449,N_11861,N_11613);
or U12450 (N_12450,N_11731,N_11821);
and U12451 (N_12451,N_11733,N_11814);
and U12452 (N_12452,N_11777,N_11675);
nand U12453 (N_12453,N_11562,N_11740);
nand U12454 (N_12454,N_11534,N_11541);
nand U12455 (N_12455,N_11734,N_11891);
xor U12456 (N_12456,N_11949,N_11675);
xnor U12457 (N_12457,N_11942,N_11971);
nor U12458 (N_12458,N_11686,N_11595);
or U12459 (N_12459,N_11521,N_11813);
nor U12460 (N_12460,N_11718,N_11735);
and U12461 (N_12461,N_11673,N_11560);
nor U12462 (N_12462,N_11765,N_11420);
xnor U12463 (N_12463,N_11620,N_11543);
xor U12464 (N_12464,N_11791,N_11868);
xnor U12465 (N_12465,N_11899,N_11493);
nand U12466 (N_12466,N_11515,N_11860);
or U12467 (N_12467,N_11847,N_11660);
nand U12468 (N_12468,N_11457,N_11975);
nor U12469 (N_12469,N_11728,N_11563);
xnor U12470 (N_12470,N_11523,N_11891);
and U12471 (N_12471,N_11498,N_11782);
nand U12472 (N_12472,N_11536,N_11608);
nand U12473 (N_12473,N_11672,N_11678);
nor U12474 (N_12474,N_11645,N_11933);
and U12475 (N_12475,N_11504,N_11725);
nor U12476 (N_12476,N_11868,N_11810);
nor U12477 (N_12477,N_11798,N_11708);
nand U12478 (N_12478,N_11618,N_11713);
nand U12479 (N_12479,N_11673,N_11713);
nand U12480 (N_12480,N_11788,N_11996);
xnor U12481 (N_12481,N_11417,N_11421);
nand U12482 (N_12482,N_11609,N_11599);
and U12483 (N_12483,N_11552,N_11543);
nand U12484 (N_12484,N_11803,N_11645);
and U12485 (N_12485,N_11519,N_11860);
xnor U12486 (N_12486,N_11758,N_11464);
nor U12487 (N_12487,N_11509,N_11925);
xor U12488 (N_12488,N_11838,N_11674);
nor U12489 (N_12489,N_11950,N_11846);
xor U12490 (N_12490,N_11863,N_11616);
xor U12491 (N_12491,N_11664,N_11447);
nand U12492 (N_12492,N_11543,N_11764);
nand U12493 (N_12493,N_11529,N_11632);
nor U12494 (N_12494,N_11787,N_11718);
nand U12495 (N_12495,N_11904,N_11802);
and U12496 (N_12496,N_11935,N_11520);
and U12497 (N_12497,N_11597,N_11971);
or U12498 (N_12498,N_11671,N_11577);
xnor U12499 (N_12499,N_11509,N_11648);
nor U12500 (N_12500,N_11530,N_11538);
nand U12501 (N_12501,N_11456,N_11688);
nand U12502 (N_12502,N_11999,N_11609);
or U12503 (N_12503,N_11930,N_11756);
or U12504 (N_12504,N_11676,N_11642);
and U12505 (N_12505,N_11418,N_11929);
nor U12506 (N_12506,N_11808,N_11487);
nand U12507 (N_12507,N_11590,N_11833);
nor U12508 (N_12508,N_11430,N_11663);
nor U12509 (N_12509,N_11810,N_11861);
nand U12510 (N_12510,N_11625,N_11559);
or U12511 (N_12511,N_11469,N_11524);
or U12512 (N_12512,N_11535,N_11523);
nor U12513 (N_12513,N_11414,N_11798);
nor U12514 (N_12514,N_11930,N_11824);
and U12515 (N_12515,N_11539,N_11477);
nor U12516 (N_12516,N_11785,N_11557);
nand U12517 (N_12517,N_11402,N_11759);
and U12518 (N_12518,N_11477,N_11860);
and U12519 (N_12519,N_11985,N_11475);
or U12520 (N_12520,N_11641,N_11625);
nand U12521 (N_12521,N_11847,N_11806);
nor U12522 (N_12522,N_11587,N_11876);
nor U12523 (N_12523,N_11450,N_11639);
nand U12524 (N_12524,N_11518,N_11662);
or U12525 (N_12525,N_11638,N_11515);
nand U12526 (N_12526,N_11975,N_11604);
nand U12527 (N_12527,N_11681,N_11492);
xor U12528 (N_12528,N_11938,N_11461);
nor U12529 (N_12529,N_11715,N_11974);
and U12530 (N_12530,N_11687,N_11500);
nand U12531 (N_12531,N_11507,N_11714);
xor U12532 (N_12532,N_11689,N_11995);
nand U12533 (N_12533,N_11897,N_11859);
nand U12534 (N_12534,N_11630,N_11572);
nor U12535 (N_12535,N_11928,N_11625);
xor U12536 (N_12536,N_11634,N_11514);
and U12537 (N_12537,N_11477,N_11940);
or U12538 (N_12538,N_11454,N_11517);
nand U12539 (N_12539,N_11823,N_11697);
xor U12540 (N_12540,N_11636,N_11417);
xnor U12541 (N_12541,N_11511,N_11862);
nor U12542 (N_12542,N_11988,N_11999);
or U12543 (N_12543,N_11786,N_11845);
and U12544 (N_12544,N_11882,N_11907);
nand U12545 (N_12545,N_11622,N_11851);
and U12546 (N_12546,N_11826,N_11682);
nand U12547 (N_12547,N_11730,N_11520);
xnor U12548 (N_12548,N_11950,N_11812);
or U12549 (N_12549,N_11966,N_11912);
nand U12550 (N_12550,N_11513,N_11923);
and U12551 (N_12551,N_11881,N_11642);
or U12552 (N_12552,N_11461,N_11743);
nand U12553 (N_12553,N_11728,N_11825);
or U12554 (N_12554,N_11775,N_11627);
nor U12555 (N_12555,N_11747,N_11827);
nand U12556 (N_12556,N_11803,N_11697);
or U12557 (N_12557,N_11615,N_11718);
nand U12558 (N_12558,N_11591,N_11409);
nor U12559 (N_12559,N_11455,N_11408);
nor U12560 (N_12560,N_11816,N_11933);
xnor U12561 (N_12561,N_11863,N_11966);
nand U12562 (N_12562,N_11859,N_11419);
xor U12563 (N_12563,N_11620,N_11479);
xor U12564 (N_12564,N_11744,N_11743);
nand U12565 (N_12565,N_11746,N_11980);
and U12566 (N_12566,N_11718,N_11878);
nor U12567 (N_12567,N_11657,N_11706);
and U12568 (N_12568,N_11951,N_11955);
or U12569 (N_12569,N_11449,N_11637);
and U12570 (N_12570,N_11846,N_11785);
and U12571 (N_12571,N_11757,N_11654);
nand U12572 (N_12572,N_11692,N_11839);
and U12573 (N_12573,N_11911,N_11448);
or U12574 (N_12574,N_11427,N_11774);
and U12575 (N_12575,N_11923,N_11779);
and U12576 (N_12576,N_11826,N_11840);
nand U12577 (N_12577,N_11714,N_11855);
or U12578 (N_12578,N_11730,N_11425);
xnor U12579 (N_12579,N_11447,N_11863);
nor U12580 (N_12580,N_11792,N_11674);
or U12581 (N_12581,N_11770,N_11998);
nand U12582 (N_12582,N_11520,N_11732);
nand U12583 (N_12583,N_11646,N_11422);
or U12584 (N_12584,N_11527,N_11763);
or U12585 (N_12585,N_11778,N_11828);
nor U12586 (N_12586,N_11915,N_11644);
or U12587 (N_12587,N_11517,N_11964);
or U12588 (N_12588,N_11777,N_11408);
nand U12589 (N_12589,N_11838,N_11984);
nand U12590 (N_12590,N_11482,N_11848);
nand U12591 (N_12591,N_11730,N_11798);
and U12592 (N_12592,N_11425,N_11534);
xor U12593 (N_12593,N_11495,N_11586);
and U12594 (N_12594,N_11462,N_11905);
and U12595 (N_12595,N_11504,N_11880);
xor U12596 (N_12596,N_11880,N_11792);
or U12597 (N_12597,N_11401,N_11616);
and U12598 (N_12598,N_11931,N_11771);
and U12599 (N_12599,N_11614,N_11658);
xor U12600 (N_12600,N_12204,N_12024);
nand U12601 (N_12601,N_12583,N_12334);
nor U12602 (N_12602,N_12070,N_12187);
nand U12603 (N_12603,N_12549,N_12189);
or U12604 (N_12604,N_12474,N_12177);
and U12605 (N_12605,N_12476,N_12430);
xor U12606 (N_12606,N_12292,N_12069);
nor U12607 (N_12607,N_12079,N_12023);
and U12608 (N_12608,N_12447,N_12271);
and U12609 (N_12609,N_12360,N_12379);
and U12610 (N_12610,N_12308,N_12550);
nor U12611 (N_12611,N_12105,N_12016);
nor U12612 (N_12612,N_12585,N_12009);
and U12613 (N_12613,N_12061,N_12504);
nand U12614 (N_12614,N_12175,N_12561);
nor U12615 (N_12615,N_12290,N_12176);
nor U12616 (N_12616,N_12399,N_12555);
or U12617 (N_12617,N_12587,N_12395);
nor U12618 (N_12618,N_12309,N_12442);
and U12619 (N_12619,N_12378,N_12118);
and U12620 (N_12620,N_12059,N_12331);
nor U12621 (N_12621,N_12517,N_12147);
or U12622 (N_12622,N_12344,N_12169);
and U12623 (N_12623,N_12201,N_12060);
nand U12624 (N_12624,N_12015,N_12164);
nor U12625 (N_12625,N_12248,N_12314);
and U12626 (N_12626,N_12302,N_12250);
or U12627 (N_12627,N_12514,N_12579);
nor U12628 (N_12628,N_12325,N_12202);
nor U12629 (N_12629,N_12380,N_12184);
nor U12630 (N_12630,N_12007,N_12212);
xnor U12631 (N_12631,N_12149,N_12244);
xor U12632 (N_12632,N_12075,N_12027);
xnor U12633 (N_12633,N_12017,N_12095);
xor U12634 (N_12634,N_12339,N_12558);
xnor U12635 (N_12635,N_12537,N_12246);
or U12636 (N_12636,N_12590,N_12192);
xor U12637 (N_12637,N_12569,N_12371);
xor U12638 (N_12638,N_12127,N_12006);
xnor U12639 (N_12639,N_12531,N_12272);
or U12640 (N_12640,N_12256,N_12274);
nor U12641 (N_12641,N_12416,N_12042);
and U12642 (N_12642,N_12479,N_12444);
or U12643 (N_12643,N_12289,N_12566);
and U12644 (N_12644,N_12459,N_12520);
and U12645 (N_12645,N_12232,N_12300);
xnor U12646 (N_12646,N_12054,N_12093);
and U12647 (N_12647,N_12159,N_12172);
nor U12648 (N_12648,N_12564,N_12056);
or U12649 (N_12649,N_12083,N_12515);
nand U12650 (N_12650,N_12461,N_12032);
nor U12651 (N_12651,N_12073,N_12365);
and U12652 (N_12652,N_12264,N_12364);
nand U12653 (N_12653,N_12422,N_12151);
and U12654 (N_12654,N_12110,N_12130);
or U12655 (N_12655,N_12091,N_12100);
nand U12656 (N_12656,N_12280,N_12522);
xnor U12657 (N_12657,N_12484,N_12320);
nand U12658 (N_12658,N_12472,N_12085);
or U12659 (N_12659,N_12008,N_12021);
or U12660 (N_12660,N_12262,N_12082);
xor U12661 (N_12661,N_12124,N_12431);
and U12662 (N_12662,N_12166,N_12539);
or U12663 (N_12663,N_12065,N_12045);
xnor U12664 (N_12664,N_12327,N_12552);
or U12665 (N_12665,N_12198,N_12038);
and U12666 (N_12666,N_12348,N_12078);
xnor U12667 (N_12667,N_12146,N_12443);
and U12668 (N_12668,N_12374,N_12414);
nand U12669 (N_12669,N_12421,N_12532);
nand U12670 (N_12670,N_12261,N_12129);
nand U12671 (N_12671,N_12133,N_12286);
nor U12672 (N_12672,N_12209,N_12115);
nand U12673 (N_12673,N_12597,N_12516);
xnor U12674 (N_12674,N_12557,N_12301);
nand U12675 (N_12675,N_12171,N_12234);
or U12676 (N_12676,N_12071,N_12485);
nand U12677 (N_12677,N_12230,N_12036);
or U12678 (N_12678,N_12375,N_12362);
or U12679 (N_12679,N_12551,N_12575);
nand U12680 (N_12680,N_12162,N_12340);
and U12681 (N_12681,N_12063,N_12119);
nand U12682 (N_12682,N_12150,N_12584);
xnor U12683 (N_12683,N_12132,N_12243);
nor U12684 (N_12684,N_12004,N_12306);
xor U12685 (N_12685,N_12505,N_12452);
nor U12686 (N_12686,N_12295,N_12219);
and U12687 (N_12687,N_12346,N_12384);
or U12688 (N_12688,N_12040,N_12237);
nor U12689 (N_12689,N_12102,N_12324);
or U12690 (N_12690,N_12586,N_12254);
nor U12691 (N_12691,N_12429,N_12594);
nand U12692 (N_12692,N_12012,N_12253);
or U12693 (N_12693,N_12477,N_12310);
xor U12694 (N_12694,N_12456,N_12455);
and U12695 (N_12695,N_12178,N_12353);
xor U12696 (N_12696,N_12490,N_12086);
nor U12697 (N_12697,N_12229,N_12396);
nand U12698 (N_12698,N_12596,N_12037);
xor U12699 (N_12699,N_12376,N_12231);
or U12700 (N_12700,N_12465,N_12134);
nor U12701 (N_12701,N_12293,N_12047);
and U12702 (N_12702,N_12556,N_12480);
xor U12703 (N_12703,N_12413,N_12260);
xor U12704 (N_12704,N_12528,N_12043);
or U12705 (N_12705,N_12001,N_12299);
nor U12706 (N_12706,N_12251,N_12407);
nand U12707 (N_12707,N_12279,N_12161);
nand U12708 (N_12708,N_12473,N_12225);
xor U12709 (N_12709,N_12464,N_12410);
nand U12710 (N_12710,N_12144,N_12155);
nor U12711 (N_12711,N_12185,N_12457);
nor U12712 (N_12712,N_12002,N_12533);
and U12713 (N_12713,N_12143,N_12215);
nand U12714 (N_12714,N_12049,N_12417);
nor U12715 (N_12715,N_12165,N_12578);
or U12716 (N_12716,N_12535,N_12233);
nor U12717 (N_12717,N_12336,N_12525);
or U12718 (N_12718,N_12534,N_12350);
and U12719 (N_12719,N_12568,N_12033);
and U12720 (N_12720,N_12529,N_12275);
nor U12721 (N_12721,N_12546,N_12018);
and U12722 (N_12722,N_12333,N_12548);
xnor U12723 (N_12723,N_12194,N_12536);
nand U12724 (N_12724,N_12258,N_12291);
xor U12725 (N_12725,N_12276,N_12022);
or U12726 (N_12726,N_12257,N_12141);
nand U12727 (N_12727,N_12326,N_12341);
nor U12728 (N_12728,N_12495,N_12449);
nor U12729 (N_12729,N_12530,N_12298);
nand U12730 (N_12730,N_12335,N_12186);
and U12731 (N_12731,N_12524,N_12170);
xnor U12732 (N_12732,N_12440,N_12598);
nor U12733 (N_12733,N_12542,N_12218);
nor U12734 (N_12734,N_12211,N_12462);
nand U12735 (N_12735,N_12565,N_12241);
and U12736 (N_12736,N_12481,N_12106);
nand U12737 (N_12737,N_12328,N_12160);
and U12738 (N_12738,N_12377,N_12190);
xor U12739 (N_12739,N_12200,N_12148);
xnor U12740 (N_12740,N_12540,N_12010);
xnor U12741 (N_12741,N_12304,N_12057);
and U12742 (N_12742,N_12098,N_12562);
and U12743 (N_12743,N_12424,N_12064);
and U12744 (N_12744,N_12103,N_12471);
and U12745 (N_12745,N_12511,N_12181);
xnor U12746 (N_12746,N_12080,N_12434);
nor U12747 (N_12747,N_12437,N_12307);
or U12748 (N_12748,N_12268,N_12446);
nand U12749 (N_12749,N_12277,N_12389);
nor U12750 (N_12750,N_12356,N_12125);
and U12751 (N_12751,N_12199,N_12519);
nor U12752 (N_12752,N_12120,N_12267);
or U12753 (N_12753,N_12497,N_12242);
nor U12754 (N_12754,N_12428,N_12383);
nor U12755 (N_12755,N_12385,N_12288);
nor U12756 (N_12756,N_12297,N_12468);
xor U12757 (N_12757,N_12094,N_12240);
nand U12758 (N_12758,N_12122,N_12030);
xor U12759 (N_12759,N_12580,N_12508);
xnor U12760 (N_12760,N_12588,N_12401);
or U12761 (N_12761,N_12195,N_12019);
nor U12762 (N_12762,N_12197,N_12259);
nor U12763 (N_12763,N_12581,N_12466);
xnor U12764 (N_12764,N_12174,N_12591);
nor U12765 (N_12765,N_12107,N_12527);
nand U12766 (N_12766,N_12116,N_12453);
and U12767 (N_12767,N_12338,N_12403);
nor U12768 (N_12768,N_12330,N_12084);
or U12769 (N_12769,N_12285,N_12035);
and U12770 (N_12770,N_12478,N_12337);
or U12771 (N_12771,N_12411,N_12111);
or U12772 (N_12772,N_12191,N_12205);
or U12773 (N_12773,N_12117,N_12108);
and U12774 (N_12774,N_12226,N_12312);
and U12775 (N_12775,N_12034,N_12589);
and U12776 (N_12776,N_12222,N_12510);
nor U12777 (N_12777,N_12076,N_12553);
or U12778 (N_12778,N_12090,N_12196);
nor U12779 (N_12779,N_12432,N_12089);
or U12780 (N_12780,N_12157,N_12025);
and U12781 (N_12781,N_12492,N_12168);
or U12782 (N_12782,N_12224,N_12349);
nand U12783 (N_12783,N_12450,N_12386);
and U12784 (N_12784,N_12577,N_12303);
nor U12785 (N_12785,N_12426,N_12592);
nor U12786 (N_12786,N_12438,N_12255);
or U12787 (N_12787,N_12567,N_12572);
xor U12788 (N_12788,N_12239,N_12097);
and U12789 (N_12789,N_12563,N_12315);
nand U12790 (N_12790,N_12322,N_12469);
nor U12791 (N_12791,N_12112,N_12113);
or U12792 (N_12792,N_12390,N_12460);
nor U12793 (N_12793,N_12087,N_12415);
nand U12794 (N_12794,N_12368,N_12372);
and U12795 (N_12795,N_12152,N_12354);
and U12796 (N_12796,N_12313,N_12343);
nor U12797 (N_12797,N_12412,N_12278);
and U12798 (N_12798,N_12544,N_12055);
xor U12799 (N_12799,N_12281,N_12284);
nor U12800 (N_12800,N_12142,N_12236);
nor U12801 (N_12801,N_12109,N_12046);
nor U12802 (N_12802,N_12131,N_12135);
xnor U12803 (N_12803,N_12294,N_12296);
nand U12804 (N_12804,N_12217,N_12066);
xnor U12805 (N_12805,N_12099,N_12573);
or U12806 (N_12806,N_12595,N_12506);
or U12807 (N_12807,N_12269,N_12221);
or U12808 (N_12808,N_12538,N_12039);
nand U12809 (N_12809,N_12488,N_12287);
nor U12810 (N_12810,N_12053,N_12096);
or U12811 (N_12811,N_12458,N_12467);
or U12812 (N_12812,N_12487,N_12247);
or U12813 (N_12813,N_12020,N_12074);
xor U12814 (N_12814,N_12387,N_12173);
or U12815 (N_12815,N_12501,N_12351);
or U12816 (N_12816,N_12409,N_12317);
nor U12817 (N_12817,N_12570,N_12448);
nor U12818 (N_12818,N_12203,N_12154);
xor U12819 (N_12819,N_12183,N_12547);
nand U12820 (N_12820,N_12439,N_12206);
nor U12821 (N_12821,N_12593,N_12266);
nand U12822 (N_12822,N_12463,N_12398);
xor U12823 (N_12823,N_12545,N_12050);
nor U12824 (N_12824,N_12345,N_12483);
and U12825 (N_12825,N_12482,N_12321);
or U12826 (N_12826,N_12332,N_12139);
and U12827 (N_12827,N_12153,N_12238);
and U12828 (N_12828,N_12235,N_12489);
or U12829 (N_12829,N_12392,N_12088);
nor U12830 (N_12830,N_12114,N_12418);
nor U12831 (N_12831,N_12493,N_12503);
xor U12832 (N_12832,N_12005,N_12445);
xor U12833 (N_12833,N_12397,N_12180);
nand U12834 (N_12834,N_12560,N_12044);
nor U12835 (N_12835,N_12509,N_12491);
or U12836 (N_12836,N_12028,N_12104);
nand U12837 (N_12837,N_12423,N_12179);
nand U12838 (N_12838,N_12029,N_12311);
or U12839 (N_12839,N_12433,N_12513);
xnor U12840 (N_12840,N_12370,N_12427);
xnor U12841 (N_12841,N_12543,N_12216);
or U12842 (N_12842,N_12026,N_12145);
xnor U12843 (N_12843,N_12355,N_12394);
nand U12844 (N_12844,N_12316,N_12526);
nand U12845 (N_12845,N_12011,N_12051);
nor U12846 (N_12846,N_12363,N_12470);
and U12847 (N_12847,N_12245,N_12062);
nor U12848 (N_12848,N_12014,N_12193);
and U12849 (N_12849,N_12512,N_12419);
and U12850 (N_12850,N_12270,N_12158);
and U12851 (N_12851,N_12072,N_12381);
nand U12852 (N_12852,N_12359,N_12329);
nor U12853 (N_12853,N_12388,N_12400);
xnor U12854 (N_12854,N_12352,N_12502);
or U12855 (N_12855,N_12357,N_12496);
nand U12856 (N_12856,N_12123,N_12220);
xor U12857 (N_12857,N_12101,N_12369);
and U12858 (N_12858,N_12435,N_12052);
and U12859 (N_12859,N_12518,N_12420);
nand U12860 (N_12860,N_12582,N_12571);
or U12861 (N_12861,N_12366,N_12402);
nor U12862 (N_12862,N_12121,N_12541);
nand U12863 (N_12863,N_12265,N_12404);
and U12864 (N_12864,N_12323,N_12128);
nor U12865 (N_12865,N_12425,N_12003);
nor U12866 (N_12866,N_12406,N_12599);
xnor U12867 (N_12867,N_12227,N_12058);
nor U12868 (N_12868,N_12393,N_12136);
nand U12869 (N_12869,N_12182,N_12361);
and U12870 (N_12870,N_12000,N_12283);
xnor U12871 (N_12871,N_12405,N_12214);
nor U12872 (N_12872,N_12373,N_12041);
or U12873 (N_12873,N_12475,N_12454);
or U12874 (N_12874,N_12263,N_12521);
nand U12875 (N_12875,N_12137,N_12067);
or U12876 (N_12876,N_12282,N_12167);
or U12877 (N_12877,N_12319,N_12126);
nand U12878 (N_12878,N_12391,N_12507);
or U12879 (N_12879,N_12249,N_12081);
xor U12880 (N_12880,N_12092,N_12252);
nand U12881 (N_12881,N_12494,N_12559);
or U12882 (N_12882,N_12013,N_12031);
and U12883 (N_12883,N_12382,N_12500);
and U12884 (N_12884,N_12523,N_12367);
or U12885 (N_12885,N_12436,N_12140);
xnor U12886 (N_12886,N_12499,N_12441);
nand U12887 (N_12887,N_12498,N_12486);
and U12888 (N_12888,N_12068,N_12048);
nand U12889 (N_12889,N_12210,N_12273);
xor U12890 (N_12890,N_12208,N_12223);
nor U12891 (N_12891,N_12207,N_12347);
nand U12892 (N_12892,N_12188,N_12576);
or U12893 (N_12893,N_12077,N_12213);
nand U12894 (N_12894,N_12138,N_12342);
or U12895 (N_12895,N_12554,N_12451);
xor U12896 (N_12896,N_12318,N_12156);
and U12897 (N_12897,N_12574,N_12408);
and U12898 (N_12898,N_12305,N_12358);
nand U12899 (N_12899,N_12228,N_12163);
or U12900 (N_12900,N_12343,N_12558);
xnor U12901 (N_12901,N_12598,N_12069);
nor U12902 (N_12902,N_12162,N_12342);
nand U12903 (N_12903,N_12376,N_12132);
or U12904 (N_12904,N_12548,N_12582);
xnor U12905 (N_12905,N_12156,N_12533);
nor U12906 (N_12906,N_12254,N_12521);
nand U12907 (N_12907,N_12501,N_12170);
nor U12908 (N_12908,N_12436,N_12354);
and U12909 (N_12909,N_12316,N_12521);
xor U12910 (N_12910,N_12348,N_12445);
and U12911 (N_12911,N_12114,N_12595);
or U12912 (N_12912,N_12331,N_12391);
or U12913 (N_12913,N_12056,N_12213);
or U12914 (N_12914,N_12333,N_12512);
nor U12915 (N_12915,N_12319,N_12501);
xnor U12916 (N_12916,N_12474,N_12244);
or U12917 (N_12917,N_12231,N_12190);
and U12918 (N_12918,N_12128,N_12026);
and U12919 (N_12919,N_12004,N_12353);
or U12920 (N_12920,N_12366,N_12060);
nand U12921 (N_12921,N_12213,N_12511);
and U12922 (N_12922,N_12319,N_12176);
and U12923 (N_12923,N_12403,N_12324);
or U12924 (N_12924,N_12351,N_12038);
or U12925 (N_12925,N_12212,N_12483);
or U12926 (N_12926,N_12055,N_12541);
nand U12927 (N_12927,N_12182,N_12370);
nand U12928 (N_12928,N_12251,N_12269);
nand U12929 (N_12929,N_12443,N_12054);
nand U12930 (N_12930,N_12107,N_12176);
or U12931 (N_12931,N_12368,N_12395);
xor U12932 (N_12932,N_12592,N_12533);
or U12933 (N_12933,N_12275,N_12172);
nand U12934 (N_12934,N_12384,N_12019);
or U12935 (N_12935,N_12364,N_12431);
xnor U12936 (N_12936,N_12449,N_12216);
nor U12937 (N_12937,N_12259,N_12193);
xor U12938 (N_12938,N_12533,N_12336);
nand U12939 (N_12939,N_12305,N_12194);
xor U12940 (N_12940,N_12297,N_12438);
nor U12941 (N_12941,N_12218,N_12151);
nor U12942 (N_12942,N_12523,N_12148);
nand U12943 (N_12943,N_12073,N_12376);
or U12944 (N_12944,N_12483,N_12126);
xor U12945 (N_12945,N_12257,N_12219);
and U12946 (N_12946,N_12269,N_12259);
xnor U12947 (N_12947,N_12450,N_12115);
and U12948 (N_12948,N_12462,N_12012);
or U12949 (N_12949,N_12033,N_12362);
and U12950 (N_12950,N_12008,N_12313);
xnor U12951 (N_12951,N_12503,N_12556);
nor U12952 (N_12952,N_12596,N_12074);
xnor U12953 (N_12953,N_12521,N_12030);
nor U12954 (N_12954,N_12550,N_12502);
or U12955 (N_12955,N_12424,N_12570);
nor U12956 (N_12956,N_12167,N_12450);
nor U12957 (N_12957,N_12034,N_12567);
xnor U12958 (N_12958,N_12319,N_12512);
or U12959 (N_12959,N_12332,N_12599);
xnor U12960 (N_12960,N_12421,N_12482);
nand U12961 (N_12961,N_12500,N_12439);
nand U12962 (N_12962,N_12102,N_12240);
or U12963 (N_12963,N_12391,N_12473);
nor U12964 (N_12964,N_12478,N_12112);
nor U12965 (N_12965,N_12031,N_12209);
or U12966 (N_12966,N_12292,N_12090);
nand U12967 (N_12967,N_12434,N_12348);
and U12968 (N_12968,N_12286,N_12059);
and U12969 (N_12969,N_12377,N_12325);
nor U12970 (N_12970,N_12306,N_12459);
or U12971 (N_12971,N_12060,N_12539);
xnor U12972 (N_12972,N_12436,N_12408);
nor U12973 (N_12973,N_12536,N_12567);
nor U12974 (N_12974,N_12570,N_12413);
nand U12975 (N_12975,N_12005,N_12458);
nor U12976 (N_12976,N_12406,N_12341);
or U12977 (N_12977,N_12585,N_12296);
nor U12978 (N_12978,N_12304,N_12463);
nand U12979 (N_12979,N_12433,N_12041);
or U12980 (N_12980,N_12580,N_12250);
and U12981 (N_12981,N_12509,N_12356);
xnor U12982 (N_12982,N_12009,N_12070);
or U12983 (N_12983,N_12399,N_12240);
xor U12984 (N_12984,N_12317,N_12080);
nand U12985 (N_12985,N_12005,N_12346);
xnor U12986 (N_12986,N_12129,N_12505);
nor U12987 (N_12987,N_12295,N_12166);
xnor U12988 (N_12988,N_12378,N_12247);
and U12989 (N_12989,N_12116,N_12505);
and U12990 (N_12990,N_12510,N_12072);
xor U12991 (N_12991,N_12080,N_12476);
xnor U12992 (N_12992,N_12222,N_12145);
and U12993 (N_12993,N_12283,N_12577);
xnor U12994 (N_12994,N_12113,N_12430);
and U12995 (N_12995,N_12597,N_12591);
nor U12996 (N_12996,N_12153,N_12436);
xor U12997 (N_12997,N_12044,N_12305);
nor U12998 (N_12998,N_12491,N_12314);
nor U12999 (N_12999,N_12033,N_12001);
or U13000 (N_13000,N_12589,N_12592);
and U13001 (N_13001,N_12547,N_12435);
or U13002 (N_13002,N_12298,N_12125);
nand U13003 (N_13003,N_12114,N_12340);
and U13004 (N_13004,N_12446,N_12164);
and U13005 (N_13005,N_12544,N_12426);
xor U13006 (N_13006,N_12185,N_12064);
nand U13007 (N_13007,N_12021,N_12156);
and U13008 (N_13008,N_12010,N_12480);
or U13009 (N_13009,N_12483,N_12573);
nor U13010 (N_13010,N_12334,N_12091);
nor U13011 (N_13011,N_12350,N_12011);
nand U13012 (N_13012,N_12228,N_12482);
or U13013 (N_13013,N_12591,N_12074);
or U13014 (N_13014,N_12431,N_12476);
xnor U13015 (N_13015,N_12155,N_12025);
or U13016 (N_13016,N_12397,N_12517);
and U13017 (N_13017,N_12499,N_12274);
nor U13018 (N_13018,N_12499,N_12222);
xor U13019 (N_13019,N_12269,N_12580);
nor U13020 (N_13020,N_12352,N_12236);
xnor U13021 (N_13021,N_12088,N_12523);
nand U13022 (N_13022,N_12171,N_12247);
xor U13023 (N_13023,N_12048,N_12137);
nand U13024 (N_13024,N_12240,N_12485);
nor U13025 (N_13025,N_12236,N_12416);
or U13026 (N_13026,N_12118,N_12438);
nand U13027 (N_13027,N_12440,N_12479);
and U13028 (N_13028,N_12398,N_12147);
nand U13029 (N_13029,N_12590,N_12279);
xnor U13030 (N_13030,N_12286,N_12126);
xor U13031 (N_13031,N_12323,N_12386);
xnor U13032 (N_13032,N_12357,N_12012);
xor U13033 (N_13033,N_12320,N_12523);
xnor U13034 (N_13034,N_12359,N_12492);
nor U13035 (N_13035,N_12595,N_12499);
nor U13036 (N_13036,N_12240,N_12460);
and U13037 (N_13037,N_12233,N_12594);
nand U13038 (N_13038,N_12383,N_12016);
and U13039 (N_13039,N_12205,N_12424);
xor U13040 (N_13040,N_12588,N_12504);
or U13041 (N_13041,N_12435,N_12146);
nor U13042 (N_13042,N_12387,N_12151);
xnor U13043 (N_13043,N_12325,N_12380);
nand U13044 (N_13044,N_12102,N_12177);
or U13045 (N_13045,N_12595,N_12361);
nand U13046 (N_13046,N_12433,N_12119);
nand U13047 (N_13047,N_12191,N_12136);
and U13048 (N_13048,N_12171,N_12118);
and U13049 (N_13049,N_12432,N_12477);
or U13050 (N_13050,N_12411,N_12232);
or U13051 (N_13051,N_12549,N_12059);
or U13052 (N_13052,N_12502,N_12198);
nor U13053 (N_13053,N_12521,N_12223);
nand U13054 (N_13054,N_12321,N_12218);
and U13055 (N_13055,N_12069,N_12371);
nor U13056 (N_13056,N_12080,N_12200);
or U13057 (N_13057,N_12149,N_12181);
xor U13058 (N_13058,N_12300,N_12171);
nand U13059 (N_13059,N_12093,N_12263);
and U13060 (N_13060,N_12407,N_12324);
and U13061 (N_13061,N_12545,N_12348);
and U13062 (N_13062,N_12384,N_12028);
or U13063 (N_13063,N_12305,N_12240);
and U13064 (N_13064,N_12494,N_12263);
xor U13065 (N_13065,N_12253,N_12140);
and U13066 (N_13066,N_12282,N_12517);
nand U13067 (N_13067,N_12249,N_12143);
and U13068 (N_13068,N_12485,N_12409);
nand U13069 (N_13069,N_12006,N_12049);
and U13070 (N_13070,N_12168,N_12151);
xnor U13071 (N_13071,N_12227,N_12052);
nor U13072 (N_13072,N_12152,N_12449);
xnor U13073 (N_13073,N_12001,N_12011);
xnor U13074 (N_13074,N_12068,N_12371);
and U13075 (N_13075,N_12056,N_12308);
nor U13076 (N_13076,N_12067,N_12493);
or U13077 (N_13077,N_12048,N_12355);
nand U13078 (N_13078,N_12443,N_12063);
nor U13079 (N_13079,N_12175,N_12358);
and U13080 (N_13080,N_12172,N_12500);
xnor U13081 (N_13081,N_12549,N_12437);
and U13082 (N_13082,N_12331,N_12554);
nand U13083 (N_13083,N_12297,N_12483);
nand U13084 (N_13084,N_12094,N_12275);
or U13085 (N_13085,N_12587,N_12537);
or U13086 (N_13086,N_12345,N_12224);
nor U13087 (N_13087,N_12068,N_12144);
and U13088 (N_13088,N_12470,N_12001);
and U13089 (N_13089,N_12596,N_12498);
or U13090 (N_13090,N_12543,N_12071);
nand U13091 (N_13091,N_12441,N_12381);
nor U13092 (N_13092,N_12382,N_12330);
nand U13093 (N_13093,N_12082,N_12363);
nand U13094 (N_13094,N_12442,N_12456);
nand U13095 (N_13095,N_12462,N_12229);
nand U13096 (N_13096,N_12124,N_12265);
or U13097 (N_13097,N_12113,N_12147);
and U13098 (N_13098,N_12547,N_12420);
nor U13099 (N_13099,N_12152,N_12405);
xor U13100 (N_13100,N_12502,N_12348);
or U13101 (N_13101,N_12122,N_12047);
nor U13102 (N_13102,N_12592,N_12309);
nand U13103 (N_13103,N_12497,N_12107);
nor U13104 (N_13104,N_12280,N_12227);
nand U13105 (N_13105,N_12161,N_12082);
or U13106 (N_13106,N_12574,N_12320);
nor U13107 (N_13107,N_12196,N_12563);
and U13108 (N_13108,N_12139,N_12504);
nand U13109 (N_13109,N_12504,N_12549);
and U13110 (N_13110,N_12580,N_12502);
nor U13111 (N_13111,N_12533,N_12132);
and U13112 (N_13112,N_12369,N_12590);
and U13113 (N_13113,N_12395,N_12123);
nor U13114 (N_13114,N_12084,N_12465);
nor U13115 (N_13115,N_12486,N_12013);
nand U13116 (N_13116,N_12541,N_12064);
nor U13117 (N_13117,N_12301,N_12453);
or U13118 (N_13118,N_12425,N_12335);
nand U13119 (N_13119,N_12464,N_12217);
xnor U13120 (N_13120,N_12150,N_12196);
nand U13121 (N_13121,N_12395,N_12124);
nor U13122 (N_13122,N_12288,N_12574);
or U13123 (N_13123,N_12385,N_12152);
xnor U13124 (N_13124,N_12480,N_12445);
xor U13125 (N_13125,N_12227,N_12101);
nor U13126 (N_13126,N_12570,N_12139);
and U13127 (N_13127,N_12298,N_12504);
or U13128 (N_13128,N_12445,N_12481);
nor U13129 (N_13129,N_12552,N_12078);
nand U13130 (N_13130,N_12560,N_12045);
xor U13131 (N_13131,N_12302,N_12138);
and U13132 (N_13132,N_12007,N_12036);
and U13133 (N_13133,N_12505,N_12391);
nor U13134 (N_13134,N_12427,N_12177);
or U13135 (N_13135,N_12436,N_12562);
or U13136 (N_13136,N_12263,N_12097);
xor U13137 (N_13137,N_12443,N_12394);
xor U13138 (N_13138,N_12333,N_12499);
or U13139 (N_13139,N_12369,N_12217);
or U13140 (N_13140,N_12002,N_12432);
nand U13141 (N_13141,N_12261,N_12232);
xnor U13142 (N_13142,N_12046,N_12130);
or U13143 (N_13143,N_12387,N_12272);
and U13144 (N_13144,N_12341,N_12146);
and U13145 (N_13145,N_12163,N_12507);
nor U13146 (N_13146,N_12169,N_12420);
and U13147 (N_13147,N_12169,N_12343);
or U13148 (N_13148,N_12340,N_12535);
nand U13149 (N_13149,N_12377,N_12337);
xor U13150 (N_13150,N_12538,N_12196);
xnor U13151 (N_13151,N_12551,N_12562);
or U13152 (N_13152,N_12597,N_12497);
nor U13153 (N_13153,N_12292,N_12589);
nand U13154 (N_13154,N_12477,N_12157);
xnor U13155 (N_13155,N_12046,N_12592);
nand U13156 (N_13156,N_12192,N_12463);
nor U13157 (N_13157,N_12006,N_12418);
nand U13158 (N_13158,N_12361,N_12091);
nand U13159 (N_13159,N_12032,N_12108);
xnor U13160 (N_13160,N_12579,N_12079);
and U13161 (N_13161,N_12206,N_12344);
xor U13162 (N_13162,N_12268,N_12441);
nand U13163 (N_13163,N_12265,N_12391);
nor U13164 (N_13164,N_12068,N_12533);
and U13165 (N_13165,N_12598,N_12160);
nor U13166 (N_13166,N_12231,N_12252);
or U13167 (N_13167,N_12400,N_12353);
nand U13168 (N_13168,N_12417,N_12571);
nor U13169 (N_13169,N_12361,N_12567);
or U13170 (N_13170,N_12285,N_12367);
nor U13171 (N_13171,N_12590,N_12462);
or U13172 (N_13172,N_12341,N_12561);
nor U13173 (N_13173,N_12364,N_12237);
or U13174 (N_13174,N_12204,N_12528);
and U13175 (N_13175,N_12318,N_12270);
nor U13176 (N_13176,N_12149,N_12313);
and U13177 (N_13177,N_12465,N_12423);
and U13178 (N_13178,N_12298,N_12574);
and U13179 (N_13179,N_12423,N_12526);
xnor U13180 (N_13180,N_12418,N_12122);
nor U13181 (N_13181,N_12044,N_12541);
xor U13182 (N_13182,N_12184,N_12593);
or U13183 (N_13183,N_12295,N_12023);
or U13184 (N_13184,N_12528,N_12549);
or U13185 (N_13185,N_12553,N_12060);
xor U13186 (N_13186,N_12088,N_12474);
and U13187 (N_13187,N_12461,N_12014);
or U13188 (N_13188,N_12295,N_12341);
or U13189 (N_13189,N_12362,N_12495);
nor U13190 (N_13190,N_12102,N_12052);
nand U13191 (N_13191,N_12546,N_12285);
or U13192 (N_13192,N_12140,N_12366);
xor U13193 (N_13193,N_12126,N_12029);
xor U13194 (N_13194,N_12381,N_12453);
or U13195 (N_13195,N_12597,N_12575);
nand U13196 (N_13196,N_12213,N_12568);
xor U13197 (N_13197,N_12566,N_12551);
or U13198 (N_13198,N_12538,N_12170);
nor U13199 (N_13199,N_12348,N_12087);
nor U13200 (N_13200,N_13053,N_12633);
and U13201 (N_13201,N_12654,N_13194);
xnor U13202 (N_13202,N_13083,N_13060);
nand U13203 (N_13203,N_13070,N_12849);
xnor U13204 (N_13204,N_12947,N_12876);
or U13205 (N_13205,N_13190,N_13109);
nor U13206 (N_13206,N_13038,N_12870);
or U13207 (N_13207,N_13013,N_12943);
and U13208 (N_13208,N_12722,N_13097);
or U13209 (N_13209,N_12887,N_12999);
or U13210 (N_13210,N_13191,N_12745);
nor U13211 (N_13211,N_12914,N_12704);
nor U13212 (N_13212,N_12702,N_12858);
nand U13213 (N_13213,N_12924,N_13029);
nand U13214 (N_13214,N_12683,N_12687);
nand U13215 (N_13215,N_13164,N_13188);
xnor U13216 (N_13216,N_12988,N_12853);
nand U13217 (N_13217,N_12651,N_13000);
or U13218 (N_13218,N_13193,N_13110);
and U13219 (N_13219,N_12779,N_12739);
xnor U13220 (N_13220,N_12711,N_12882);
nor U13221 (N_13221,N_13098,N_12823);
nor U13222 (N_13222,N_12819,N_13156);
nand U13223 (N_13223,N_13159,N_13167);
and U13224 (N_13224,N_13199,N_12606);
or U13225 (N_13225,N_12657,N_12861);
nor U13226 (N_13226,N_12623,N_13006);
or U13227 (N_13227,N_12954,N_13130);
xnor U13228 (N_13228,N_13106,N_13135);
xor U13229 (N_13229,N_13021,N_12996);
nor U13230 (N_13230,N_12743,N_12729);
nor U13231 (N_13231,N_12768,N_13059);
nor U13232 (N_13232,N_13198,N_12670);
and U13233 (N_13233,N_12799,N_12913);
nor U13234 (N_13234,N_12886,N_12697);
nand U13235 (N_13235,N_12964,N_12970);
and U13236 (N_13236,N_13004,N_12663);
nand U13237 (N_13237,N_12820,N_12762);
nor U13238 (N_13238,N_12808,N_12863);
nor U13239 (N_13239,N_12978,N_12881);
xnor U13240 (N_13240,N_13008,N_12727);
and U13241 (N_13241,N_12967,N_12987);
xor U13242 (N_13242,N_13080,N_12754);
xor U13243 (N_13243,N_13035,N_12952);
xnor U13244 (N_13244,N_12777,N_13129);
nand U13245 (N_13245,N_12681,N_12844);
nor U13246 (N_13246,N_13161,N_13108);
nor U13247 (N_13247,N_12880,N_12939);
nand U13248 (N_13248,N_12766,N_12950);
nor U13249 (N_13249,N_13003,N_12692);
nand U13250 (N_13250,N_12634,N_13066);
and U13251 (N_13251,N_12982,N_13015);
nand U13252 (N_13252,N_12991,N_12966);
and U13253 (N_13253,N_13174,N_12802);
nand U13254 (N_13254,N_13044,N_13065);
xor U13255 (N_13255,N_13033,N_12610);
or U13256 (N_13256,N_12728,N_12751);
nor U13257 (N_13257,N_13137,N_12708);
nand U13258 (N_13258,N_13165,N_12804);
xnor U13259 (N_13259,N_12911,N_13048);
or U13260 (N_13260,N_12721,N_13152);
and U13261 (N_13261,N_12669,N_12738);
and U13262 (N_13262,N_12749,N_12953);
nor U13263 (N_13263,N_12998,N_13122);
or U13264 (N_13264,N_12829,N_13128);
nor U13265 (N_13265,N_13145,N_13075);
and U13266 (N_13266,N_12753,N_13104);
nand U13267 (N_13267,N_12747,N_13117);
nand U13268 (N_13268,N_13195,N_12645);
nor U13269 (N_13269,N_12686,N_12788);
xnor U13270 (N_13270,N_12856,N_12928);
and U13271 (N_13271,N_12699,N_12627);
nand U13272 (N_13272,N_12841,N_13037);
nor U13273 (N_13273,N_12984,N_12885);
xnor U13274 (N_13274,N_12850,N_12895);
nor U13275 (N_13275,N_13045,N_13031);
nor U13276 (N_13276,N_13185,N_13125);
xor U13277 (N_13277,N_13092,N_13077);
and U13278 (N_13278,N_12701,N_12626);
or U13279 (N_13279,N_12741,N_12960);
xnor U13280 (N_13280,N_12905,N_12646);
nor U13281 (N_13281,N_12784,N_13018);
xnor U13282 (N_13282,N_12857,N_12616);
and U13283 (N_13283,N_12983,N_12825);
xnor U13284 (N_13284,N_13168,N_13134);
nor U13285 (N_13285,N_12782,N_12761);
nand U13286 (N_13286,N_13192,N_12839);
nand U13287 (N_13287,N_12718,N_12621);
nor U13288 (N_13288,N_13126,N_12973);
xnor U13289 (N_13289,N_13173,N_12682);
and U13290 (N_13290,N_12814,N_12958);
xnor U13291 (N_13291,N_13020,N_13172);
and U13292 (N_13292,N_12672,N_13149);
and U13293 (N_13293,N_12688,N_12707);
nand U13294 (N_13294,N_12684,N_12828);
or U13295 (N_13295,N_13076,N_12842);
nand U13296 (N_13296,N_12740,N_12714);
and U13297 (N_13297,N_12717,N_12851);
and U13298 (N_13298,N_12685,N_13081);
nor U13299 (N_13299,N_13176,N_12665);
and U13300 (N_13300,N_12733,N_12852);
or U13301 (N_13301,N_13071,N_13099);
xor U13302 (N_13302,N_12946,N_12748);
nand U13303 (N_13303,N_13072,N_13118);
and U13304 (N_13304,N_13163,N_13111);
or U13305 (N_13305,N_12730,N_12860);
nand U13306 (N_13306,N_12894,N_12787);
and U13307 (N_13307,N_12824,N_13002);
and U13308 (N_13308,N_12703,N_13041);
xor U13309 (N_13309,N_12872,N_12818);
nand U13310 (N_13310,N_12690,N_12752);
nor U13311 (N_13311,N_12827,N_13057);
nor U13312 (N_13312,N_12866,N_12930);
and U13313 (N_13313,N_12974,N_13181);
xor U13314 (N_13314,N_12840,N_12603);
xnor U13315 (N_13315,N_13042,N_13032);
xor U13316 (N_13316,N_12622,N_13155);
nor U13317 (N_13317,N_13114,N_12644);
xor U13318 (N_13318,N_12647,N_12661);
or U13319 (N_13319,N_12656,N_13170);
nand U13320 (N_13320,N_12618,N_12901);
nand U13321 (N_13321,N_12759,N_12720);
nand U13322 (N_13322,N_13142,N_12658);
and U13323 (N_13323,N_12698,N_12710);
nor U13324 (N_13324,N_12831,N_13138);
nor U13325 (N_13325,N_13052,N_12628);
nand U13326 (N_13326,N_12900,N_13196);
and U13327 (N_13327,N_13051,N_13007);
nand U13328 (N_13328,N_12909,N_12744);
or U13329 (N_13329,N_12813,N_13025);
xor U13330 (N_13330,N_12796,N_12934);
xor U13331 (N_13331,N_12674,N_13014);
nand U13332 (N_13332,N_12920,N_12636);
and U13333 (N_13333,N_12625,N_12667);
and U13334 (N_13334,N_13093,N_12847);
or U13335 (N_13335,N_12875,N_13011);
or U13336 (N_13336,N_12812,N_13096);
xnor U13337 (N_13337,N_12919,N_12933);
and U13338 (N_13338,N_13089,N_12868);
nand U13339 (N_13339,N_12780,N_12968);
and U13340 (N_13340,N_12927,N_12836);
and U13341 (N_13341,N_12854,N_12929);
nand U13342 (N_13342,N_13091,N_12758);
or U13343 (N_13343,N_13132,N_12791);
xnor U13344 (N_13344,N_12865,N_13115);
and U13345 (N_13345,N_13180,N_12944);
xor U13346 (N_13346,N_12737,N_13189);
nand U13347 (N_13347,N_12877,N_12971);
or U13348 (N_13348,N_12725,N_12993);
nor U13349 (N_13349,N_12835,N_12951);
nand U13350 (N_13350,N_13055,N_12889);
or U13351 (N_13351,N_12602,N_12926);
nand U13352 (N_13352,N_12807,N_12871);
nor U13353 (N_13353,N_12941,N_12811);
and U13354 (N_13354,N_12679,N_12666);
nand U13355 (N_13355,N_13169,N_12936);
and U13356 (N_13356,N_12873,N_12726);
xor U13357 (N_13357,N_12822,N_13073);
nor U13358 (N_13358,N_12611,N_13088);
or U13359 (N_13359,N_12648,N_12972);
xor U13360 (N_13360,N_12785,N_12869);
nand U13361 (N_13361,N_12965,N_13078);
xnor U13362 (N_13362,N_12907,N_13123);
nor U13363 (N_13363,N_12884,N_12629);
nor U13364 (N_13364,N_12843,N_13095);
nand U13365 (N_13365,N_13184,N_13056);
xor U13366 (N_13366,N_12899,N_12801);
nand U13367 (N_13367,N_13105,N_13121);
xor U13368 (N_13368,N_12961,N_12997);
xnor U13369 (N_13369,N_12915,N_13166);
or U13370 (N_13370,N_12767,N_12662);
and U13371 (N_13371,N_12689,N_12832);
or U13372 (N_13372,N_12723,N_13197);
nand U13373 (N_13373,N_12677,N_13124);
or U13374 (N_13374,N_12792,N_12923);
xnor U13375 (N_13375,N_12653,N_13141);
nor U13376 (N_13376,N_12879,N_13119);
nor U13377 (N_13377,N_12680,N_12945);
nor U13378 (N_13378,N_12992,N_13040);
nand U13379 (N_13379,N_12770,N_12937);
and U13380 (N_13380,N_12632,N_12691);
and U13381 (N_13381,N_12922,N_13147);
nand U13382 (N_13382,N_12990,N_12916);
xor U13383 (N_13383,N_12794,N_12659);
and U13384 (N_13384,N_12910,N_12673);
or U13385 (N_13385,N_12675,N_12620);
xnor U13386 (N_13386,N_12678,N_12630);
or U13387 (N_13387,N_13046,N_12609);
nor U13388 (N_13388,N_12918,N_13094);
xnor U13389 (N_13389,N_12908,N_13064);
or U13390 (N_13390,N_12848,N_12601);
xor U13391 (N_13391,N_13027,N_13133);
or U13392 (N_13392,N_13107,N_12912);
and U13393 (N_13393,N_12898,N_13102);
nand U13394 (N_13394,N_12883,N_12734);
nand U13395 (N_13395,N_13101,N_13116);
nor U13396 (N_13396,N_12994,N_12709);
xor U13397 (N_13397,N_13017,N_12715);
xnor U13398 (N_13398,N_12816,N_13079);
or U13399 (N_13399,N_12962,N_12649);
xor U13400 (N_13400,N_12642,N_12846);
xor U13401 (N_13401,N_12817,N_12763);
xnor U13402 (N_13402,N_13085,N_12896);
nand U13403 (N_13403,N_12948,N_12890);
xor U13404 (N_13404,N_12830,N_13074);
and U13405 (N_13405,N_12652,N_12774);
nor U13406 (N_13406,N_12949,N_13019);
and U13407 (N_13407,N_12955,N_12862);
nor U13408 (N_13408,N_12985,N_12724);
or U13409 (N_13409,N_13010,N_12891);
nand U13410 (N_13410,N_13162,N_13039);
xor U13411 (N_13411,N_13036,N_13030);
nor U13412 (N_13412,N_13049,N_12719);
and U13413 (N_13413,N_12980,N_12775);
nor U13414 (N_13414,N_13150,N_12638);
nor U13415 (N_13415,N_13069,N_12750);
and U13416 (N_13416,N_13175,N_13144);
nand U13417 (N_13417,N_12809,N_13054);
nand U13418 (N_13418,N_13154,N_13131);
nor U13419 (N_13419,N_12641,N_12765);
nor U13420 (N_13420,N_13143,N_12859);
xor U13421 (N_13421,N_12706,N_13086);
xor U13422 (N_13422,N_13016,N_12639);
and U13423 (N_13423,N_12878,N_12668);
nor U13424 (N_13424,N_12778,N_12833);
and U13425 (N_13425,N_12742,N_13084);
nand U13426 (N_13426,N_13012,N_12906);
xnor U13427 (N_13427,N_12771,N_12693);
xnor U13428 (N_13428,N_12746,N_12643);
or U13429 (N_13429,N_12855,N_12925);
and U13430 (N_13430,N_13140,N_13179);
or U13431 (N_13431,N_12904,N_13160);
and U13432 (N_13432,N_12783,N_12821);
nand U13433 (N_13433,N_12938,N_12864);
or U13434 (N_13434,N_12612,N_12977);
nand U13435 (N_13435,N_12769,N_13047);
xnor U13436 (N_13436,N_12772,N_13087);
nor U13437 (N_13437,N_13001,N_13058);
xor U13438 (N_13438,N_12607,N_12764);
nand U13439 (N_13439,N_13148,N_13171);
or U13440 (N_13440,N_13061,N_13034);
and U13441 (N_13441,N_12845,N_12986);
or U13442 (N_13442,N_13063,N_12874);
and U13443 (N_13443,N_12838,N_12795);
nor U13444 (N_13444,N_13139,N_13136);
nand U13445 (N_13445,N_12614,N_12805);
and U13446 (N_13446,N_12963,N_12732);
or U13447 (N_13447,N_12940,N_13023);
xnor U13448 (N_13448,N_13100,N_13028);
xnor U13449 (N_13449,N_13043,N_13153);
nor U13450 (N_13450,N_12650,N_12776);
and U13451 (N_13451,N_12893,N_13050);
and U13452 (N_13452,N_12989,N_13068);
xor U13453 (N_13453,N_13187,N_12615);
or U13454 (N_13454,N_12773,N_13113);
or U13455 (N_13455,N_12716,N_12760);
nor U13456 (N_13456,N_13112,N_12789);
nor U13457 (N_13457,N_12637,N_12935);
nand U13458 (N_13458,N_13146,N_13009);
and U13459 (N_13459,N_12903,N_12837);
or U13460 (N_13460,N_13090,N_12735);
and U13461 (N_13461,N_12608,N_12731);
or U13462 (N_13462,N_12696,N_12640);
xor U13463 (N_13463,N_12867,N_12655);
nor U13464 (N_13464,N_12613,N_12959);
or U13465 (N_13465,N_13067,N_12736);
and U13466 (N_13466,N_12712,N_12676);
nand U13467 (N_13467,N_12981,N_12921);
and U13468 (N_13468,N_12781,N_12790);
nand U13469 (N_13469,N_12619,N_12635);
nor U13470 (N_13470,N_12756,N_12956);
nand U13471 (N_13471,N_12834,N_12713);
or U13472 (N_13472,N_13158,N_13103);
xor U13473 (N_13473,N_12975,N_13026);
nor U13474 (N_13474,N_12604,N_13186);
and U13475 (N_13475,N_13157,N_13178);
xnor U13476 (N_13476,N_12969,N_13151);
nor U13477 (N_13477,N_12892,N_13022);
xor U13478 (N_13478,N_12797,N_12806);
xor U13479 (N_13479,N_13177,N_12979);
nand U13480 (N_13480,N_12694,N_12793);
nand U13481 (N_13481,N_13183,N_12931);
or U13482 (N_13482,N_12695,N_12803);
nor U13483 (N_13483,N_12786,N_12700);
nand U13484 (N_13484,N_12888,N_12705);
nor U13485 (N_13485,N_12798,N_12810);
nand U13486 (N_13486,N_12976,N_12757);
nor U13487 (N_13487,N_12800,N_12942);
and U13488 (N_13488,N_12932,N_12664);
and U13489 (N_13489,N_13005,N_13062);
nor U13490 (N_13490,N_12957,N_12917);
or U13491 (N_13491,N_13024,N_12897);
and U13492 (N_13492,N_12600,N_12631);
and U13493 (N_13493,N_13182,N_12617);
and U13494 (N_13494,N_12995,N_12671);
nand U13495 (N_13495,N_12902,N_12624);
nand U13496 (N_13496,N_13082,N_12826);
nand U13497 (N_13497,N_13120,N_12605);
and U13498 (N_13498,N_12815,N_13127);
or U13499 (N_13499,N_12660,N_12755);
xor U13500 (N_13500,N_13137,N_12655);
nand U13501 (N_13501,N_12644,N_12827);
nor U13502 (N_13502,N_13011,N_12858);
or U13503 (N_13503,N_12877,N_12923);
and U13504 (N_13504,N_12741,N_12944);
and U13505 (N_13505,N_12744,N_12819);
or U13506 (N_13506,N_12743,N_12718);
and U13507 (N_13507,N_12693,N_12788);
nor U13508 (N_13508,N_13185,N_13180);
or U13509 (N_13509,N_12768,N_12708);
xnor U13510 (N_13510,N_13176,N_12757);
xor U13511 (N_13511,N_13015,N_12744);
nand U13512 (N_13512,N_12683,N_12680);
nand U13513 (N_13513,N_12633,N_13115);
xnor U13514 (N_13514,N_12805,N_12760);
xnor U13515 (N_13515,N_12975,N_12754);
xnor U13516 (N_13516,N_12604,N_12769);
nor U13517 (N_13517,N_13071,N_12841);
nor U13518 (N_13518,N_12721,N_13078);
or U13519 (N_13519,N_12761,N_12929);
nor U13520 (N_13520,N_12986,N_12852);
and U13521 (N_13521,N_13042,N_12763);
or U13522 (N_13522,N_12778,N_12724);
nand U13523 (N_13523,N_12724,N_12933);
or U13524 (N_13524,N_12780,N_13041);
or U13525 (N_13525,N_12858,N_12784);
xnor U13526 (N_13526,N_12815,N_12975);
or U13527 (N_13527,N_12625,N_12982);
nor U13528 (N_13528,N_12668,N_12848);
or U13529 (N_13529,N_12819,N_13180);
and U13530 (N_13530,N_13094,N_12907);
xnor U13531 (N_13531,N_13033,N_13062);
nand U13532 (N_13532,N_12957,N_12648);
or U13533 (N_13533,N_12763,N_12994);
or U13534 (N_13534,N_12916,N_12946);
nand U13535 (N_13535,N_13199,N_12729);
nor U13536 (N_13536,N_12845,N_12782);
or U13537 (N_13537,N_12865,N_12702);
and U13538 (N_13538,N_12817,N_12843);
xor U13539 (N_13539,N_13152,N_13095);
or U13540 (N_13540,N_12901,N_13093);
or U13541 (N_13541,N_12640,N_12967);
and U13542 (N_13542,N_12601,N_12824);
or U13543 (N_13543,N_12627,N_13006);
xor U13544 (N_13544,N_13099,N_12939);
nand U13545 (N_13545,N_12947,N_12822);
nor U13546 (N_13546,N_13144,N_13034);
or U13547 (N_13547,N_12692,N_13169);
and U13548 (N_13548,N_12874,N_13095);
xor U13549 (N_13549,N_13001,N_12704);
nor U13550 (N_13550,N_13089,N_12964);
or U13551 (N_13551,N_12641,N_13083);
or U13552 (N_13552,N_12965,N_13023);
or U13553 (N_13553,N_12785,N_12867);
nand U13554 (N_13554,N_13081,N_12619);
and U13555 (N_13555,N_12753,N_12742);
or U13556 (N_13556,N_12618,N_13177);
nor U13557 (N_13557,N_12876,N_12666);
xnor U13558 (N_13558,N_12932,N_12845);
and U13559 (N_13559,N_13015,N_13170);
nor U13560 (N_13560,N_12903,N_12842);
nand U13561 (N_13561,N_12758,N_12819);
nor U13562 (N_13562,N_12940,N_13032);
xor U13563 (N_13563,N_13002,N_12727);
nand U13564 (N_13564,N_12937,N_12885);
nand U13565 (N_13565,N_12705,N_12667);
and U13566 (N_13566,N_13188,N_12801);
and U13567 (N_13567,N_12811,N_13063);
xnor U13568 (N_13568,N_12876,N_13164);
xnor U13569 (N_13569,N_12646,N_12865);
nor U13570 (N_13570,N_12908,N_13005);
and U13571 (N_13571,N_13065,N_12876);
or U13572 (N_13572,N_12746,N_13132);
nand U13573 (N_13573,N_13026,N_13196);
and U13574 (N_13574,N_12811,N_12972);
and U13575 (N_13575,N_12907,N_12820);
nand U13576 (N_13576,N_12749,N_13170);
nand U13577 (N_13577,N_12823,N_12965);
nand U13578 (N_13578,N_12605,N_12816);
or U13579 (N_13579,N_12778,N_13174);
nand U13580 (N_13580,N_12909,N_12939);
xnor U13581 (N_13581,N_12962,N_13117);
nand U13582 (N_13582,N_12989,N_13102);
nor U13583 (N_13583,N_13154,N_13143);
xor U13584 (N_13584,N_12888,N_12783);
xnor U13585 (N_13585,N_13062,N_12921);
and U13586 (N_13586,N_12609,N_12725);
xor U13587 (N_13587,N_12986,N_12756);
nor U13588 (N_13588,N_12943,N_13025);
or U13589 (N_13589,N_12740,N_12733);
or U13590 (N_13590,N_12828,N_13029);
nand U13591 (N_13591,N_12722,N_12846);
xor U13592 (N_13592,N_13031,N_12824);
and U13593 (N_13593,N_12872,N_13105);
nand U13594 (N_13594,N_12718,N_13053);
xnor U13595 (N_13595,N_13115,N_13118);
nand U13596 (N_13596,N_13034,N_13107);
nand U13597 (N_13597,N_12841,N_13042);
or U13598 (N_13598,N_13169,N_12742);
and U13599 (N_13599,N_12859,N_13163);
and U13600 (N_13600,N_12726,N_12787);
xor U13601 (N_13601,N_12882,N_13122);
nand U13602 (N_13602,N_12858,N_12861);
and U13603 (N_13603,N_12769,N_13194);
nand U13604 (N_13604,N_12731,N_13163);
or U13605 (N_13605,N_13029,N_12648);
xor U13606 (N_13606,N_12803,N_12749);
and U13607 (N_13607,N_13196,N_12808);
xnor U13608 (N_13608,N_12960,N_13168);
nor U13609 (N_13609,N_12898,N_13046);
nand U13610 (N_13610,N_12949,N_12659);
or U13611 (N_13611,N_12734,N_12699);
nand U13612 (N_13612,N_12749,N_13185);
nand U13613 (N_13613,N_13048,N_12870);
nand U13614 (N_13614,N_12805,N_13179);
and U13615 (N_13615,N_12616,N_12750);
nand U13616 (N_13616,N_12999,N_12972);
nand U13617 (N_13617,N_12762,N_13037);
nand U13618 (N_13618,N_13143,N_12775);
nor U13619 (N_13619,N_12912,N_13157);
nand U13620 (N_13620,N_12616,N_12672);
and U13621 (N_13621,N_12892,N_12718);
xor U13622 (N_13622,N_12984,N_13027);
xor U13623 (N_13623,N_12974,N_13089);
and U13624 (N_13624,N_12661,N_12969);
and U13625 (N_13625,N_12619,N_12610);
nor U13626 (N_13626,N_13156,N_12617);
nand U13627 (N_13627,N_12688,N_12949);
or U13628 (N_13628,N_12938,N_12793);
nor U13629 (N_13629,N_12878,N_12980);
xnor U13630 (N_13630,N_12891,N_12614);
and U13631 (N_13631,N_12669,N_13133);
nand U13632 (N_13632,N_12626,N_12639);
nor U13633 (N_13633,N_12783,N_13132);
nor U13634 (N_13634,N_12784,N_12880);
or U13635 (N_13635,N_12881,N_13077);
and U13636 (N_13636,N_12831,N_12885);
or U13637 (N_13637,N_13138,N_13111);
or U13638 (N_13638,N_13049,N_13127);
nand U13639 (N_13639,N_12664,N_12799);
nand U13640 (N_13640,N_12831,N_12882);
nand U13641 (N_13641,N_12628,N_13119);
nor U13642 (N_13642,N_12851,N_12711);
nor U13643 (N_13643,N_12612,N_12978);
and U13644 (N_13644,N_12888,N_12676);
or U13645 (N_13645,N_12795,N_13077);
or U13646 (N_13646,N_12905,N_13060);
xnor U13647 (N_13647,N_13060,N_12622);
and U13648 (N_13648,N_12687,N_12700);
and U13649 (N_13649,N_13085,N_13141);
and U13650 (N_13650,N_12967,N_12994);
nand U13651 (N_13651,N_13070,N_12628);
and U13652 (N_13652,N_12672,N_12692);
and U13653 (N_13653,N_13124,N_12785);
xor U13654 (N_13654,N_12824,N_13162);
and U13655 (N_13655,N_12955,N_12924);
nor U13656 (N_13656,N_12853,N_12813);
nor U13657 (N_13657,N_12839,N_13156);
xor U13658 (N_13658,N_12827,N_12972);
and U13659 (N_13659,N_13142,N_12927);
or U13660 (N_13660,N_12850,N_12962);
nand U13661 (N_13661,N_12853,N_12602);
xnor U13662 (N_13662,N_12928,N_12853);
nor U13663 (N_13663,N_13037,N_12812);
xor U13664 (N_13664,N_12767,N_12865);
xnor U13665 (N_13665,N_12788,N_12759);
or U13666 (N_13666,N_12742,N_13114);
nand U13667 (N_13667,N_12974,N_12724);
and U13668 (N_13668,N_13161,N_13039);
nand U13669 (N_13669,N_13035,N_13031);
or U13670 (N_13670,N_13051,N_13197);
nand U13671 (N_13671,N_12877,N_12852);
xor U13672 (N_13672,N_13014,N_12728);
nand U13673 (N_13673,N_12743,N_12672);
nand U13674 (N_13674,N_12654,N_12866);
nor U13675 (N_13675,N_12678,N_12694);
or U13676 (N_13676,N_12788,N_12993);
and U13677 (N_13677,N_12943,N_12817);
or U13678 (N_13678,N_12892,N_13103);
or U13679 (N_13679,N_12745,N_13167);
or U13680 (N_13680,N_12623,N_12702);
or U13681 (N_13681,N_13088,N_12905);
nand U13682 (N_13682,N_13196,N_13184);
or U13683 (N_13683,N_13194,N_12658);
or U13684 (N_13684,N_12600,N_12759);
nor U13685 (N_13685,N_12611,N_12994);
and U13686 (N_13686,N_13084,N_12973);
or U13687 (N_13687,N_13080,N_13053);
nor U13688 (N_13688,N_12614,N_12929);
nor U13689 (N_13689,N_12621,N_13151);
or U13690 (N_13690,N_12818,N_12736);
or U13691 (N_13691,N_12941,N_13177);
nor U13692 (N_13692,N_12906,N_12975);
xor U13693 (N_13693,N_13084,N_12647);
nand U13694 (N_13694,N_12695,N_12992);
or U13695 (N_13695,N_13026,N_12646);
nor U13696 (N_13696,N_12661,N_12760);
or U13697 (N_13697,N_12969,N_13140);
nor U13698 (N_13698,N_12807,N_12844);
nand U13699 (N_13699,N_13104,N_12848);
nor U13700 (N_13700,N_13031,N_12691);
nand U13701 (N_13701,N_12961,N_12999);
nor U13702 (N_13702,N_13077,N_13019);
nand U13703 (N_13703,N_13159,N_12703);
nand U13704 (N_13704,N_13081,N_13096);
xor U13705 (N_13705,N_12998,N_12726);
and U13706 (N_13706,N_12638,N_12641);
nand U13707 (N_13707,N_13071,N_12730);
nand U13708 (N_13708,N_12615,N_12882);
or U13709 (N_13709,N_13044,N_12957);
xor U13710 (N_13710,N_12829,N_12774);
xor U13711 (N_13711,N_13190,N_12950);
nand U13712 (N_13712,N_12939,N_12648);
and U13713 (N_13713,N_12911,N_12698);
or U13714 (N_13714,N_13171,N_12765);
nor U13715 (N_13715,N_12870,N_12991);
nor U13716 (N_13716,N_12968,N_13170);
or U13717 (N_13717,N_12762,N_12613);
or U13718 (N_13718,N_13038,N_13127);
nand U13719 (N_13719,N_12855,N_12739);
and U13720 (N_13720,N_13007,N_12958);
or U13721 (N_13721,N_13136,N_12942);
nor U13722 (N_13722,N_12956,N_12675);
or U13723 (N_13723,N_12984,N_12647);
nor U13724 (N_13724,N_12838,N_12625);
and U13725 (N_13725,N_13046,N_12743);
xnor U13726 (N_13726,N_12789,N_12995);
or U13727 (N_13727,N_12719,N_12722);
xor U13728 (N_13728,N_13164,N_13096);
xnor U13729 (N_13729,N_13091,N_12634);
or U13730 (N_13730,N_12681,N_12911);
nand U13731 (N_13731,N_12858,N_12695);
or U13732 (N_13732,N_13197,N_12648);
nand U13733 (N_13733,N_12679,N_12630);
nor U13734 (N_13734,N_12626,N_13167);
nand U13735 (N_13735,N_13096,N_13070);
nand U13736 (N_13736,N_12845,N_12901);
nand U13737 (N_13737,N_12851,N_12650);
nand U13738 (N_13738,N_13088,N_13087);
and U13739 (N_13739,N_12842,N_12791);
nor U13740 (N_13740,N_12615,N_12774);
and U13741 (N_13741,N_12954,N_13142);
xor U13742 (N_13742,N_12608,N_12777);
xnor U13743 (N_13743,N_12841,N_12806);
and U13744 (N_13744,N_12713,N_13196);
and U13745 (N_13745,N_12895,N_13048);
or U13746 (N_13746,N_12993,N_12705);
nand U13747 (N_13747,N_12795,N_12682);
xor U13748 (N_13748,N_13001,N_13190);
xnor U13749 (N_13749,N_13122,N_12700);
and U13750 (N_13750,N_12792,N_12863);
nor U13751 (N_13751,N_12622,N_12760);
nor U13752 (N_13752,N_12650,N_12857);
nand U13753 (N_13753,N_12787,N_12682);
and U13754 (N_13754,N_13155,N_12908);
and U13755 (N_13755,N_13020,N_12702);
and U13756 (N_13756,N_12842,N_12702);
nand U13757 (N_13757,N_13072,N_12853);
xnor U13758 (N_13758,N_12877,N_13062);
and U13759 (N_13759,N_13126,N_12656);
nand U13760 (N_13760,N_12635,N_12880);
or U13761 (N_13761,N_13145,N_13032);
xor U13762 (N_13762,N_12702,N_12604);
xnor U13763 (N_13763,N_12960,N_12911);
nor U13764 (N_13764,N_12748,N_12827);
nand U13765 (N_13765,N_12643,N_13155);
nor U13766 (N_13766,N_13107,N_13052);
nand U13767 (N_13767,N_13091,N_12997);
xnor U13768 (N_13768,N_13172,N_13122);
or U13769 (N_13769,N_12977,N_12966);
nand U13770 (N_13770,N_12774,N_13077);
xor U13771 (N_13771,N_13153,N_13137);
nand U13772 (N_13772,N_12826,N_12621);
nand U13773 (N_13773,N_13115,N_12816);
and U13774 (N_13774,N_13051,N_12825);
xnor U13775 (N_13775,N_13121,N_12852);
nand U13776 (N_13776,N_13112,N_13169);
and U13777 (N_13777,N_12926,N_13014);
and U13778 (N_13778,N_12857,N_13033);
and U13779 (N_13779,N_12923,N_12648);
nor U13780 (N_13780,N_12906,N_13124);
and U13781 (N_13781,N_13042,N_12894);
nor U13782 (N_13782,N_12797,N_12792);
nor U13783 (N_13783,N_12871,N_12747);
xor U13784 (N_13784,N_12993,N_12782);
xor U13785 (N_13785,N_12908,N_13097);
and U13786 (N_13786,N_12869,N_13108);
or U13787 (N_13787,N_12800,N_12668);
nor U13788 (N_13788,N_13142,N_12741);
and U13789 (N_13789,N_13127,N_12936);
nand U13790 (N_13790,N_13052,N_12730);
or U13791 (N_13791,N_13199,N_13041);
and U13792 (N_13792,N_12802,N_13025);
nor U13793 (N_13793,N_12943,N_12908);
nand U13794 (N_13794,N_12905,N_12634);
xor U13795 (N_13795,N_12761,N_13168);
nand U13796 (N_13796,N_12673,N_12761);
nand U13797 (N_13797,N_12980,N_12608);
or U13798 (N_13798,N_12925,N_12630);
or U13799 (N_13799,N_12828,N_13144);
nor U13800 (N_13800,N_13233,N_13739);
nor U13801 (N_13801,N_13644,N_13356);
nand U13802 (N_13802,N_13314,N_13380);
and U13803 (N_13803,N_13389,N_13401);
nand U13804 (N_13804,N_13561,N_13336);
nand U13805 (N_13805,N_13683,N_13236);
xor U13806 (N_13806,N_13681,N_13661);
and U13807 (N_13807,N_13604,N_13284);
nand U13808 (N_13808,N_13541,N_13768);
or U13809 (N_13809,N_13760,N_13369);
nor U13810 (N_13810,N_13776,N_13650);
and U13811 (N_13811,N_13657,N_13419);
nand U13812 (N_13812,N_13576,N_13432);
and U13813 (N_13813,N_13772,N_13213);
and U13814 (N_13814,N_13619,N_13782);
xor U13815 (N_13815,N_13711,N_13338);
nor U13816 (N_13816,N_13734,N_13365);
nand U13817 (N_13817,N_13246,N_13430);
or U13818 (N_13818,N_13224,N_13656);
nand U13819 (N_13819,N_13308,N_13633);
xnor U13820 (N_13820,N_13203,N_13746);
or U13821 (N_13821,N_13567,N_13266);
or U13822 (N_13822,N_13674,N_13736);
xor U13823 (N_13823,N_13513,N_13453);
nand U13824 (N_13824,N_13276,N_13570);
xnor U13825 (N_13825,N_13415,N_13395);
or U13826 (N_13826,N_13384,N_13434);
or U13827 (N_13827,N_13406,N_13322);
xor U13828 (N_13828,N_13602,N_13547);
nor U13829 (N_13829,N_13737,N_13254);
and U13830 (N_13830,N_13536,N_13719);
and U13831 (N_13831,N_13708,N_13582);
and U13832 (N_13832,N_13222,N_13712);
nor U13833 (N_13833,N_13361,N_13529);
xor U13834 (N_13834,N_13366,N_13269);
xor U13835 (N_13835,N_13367,N_13793);
nand U13836 (N_13836,N_13429,N_13554);
and U13837 (N_13837,N_13480,N_13206);
nor U13838 (N_13838,N_13362,N_13786);
nor U13839 (N_13839,N_13634,N_13723);
or U13840 (N_13840,N_13540,N_13449);
or U13841 (N_13841,N_13718,N_13294);
and U13842 (N_13842,N_13679,N_13493);
and U13843 (N_13843,N_13358,N_13397);
nor U13844 (N_13844,N_13289,N_13629);
nand U13845 (N_13845,N_13459,N_13328);
or U13846 (N_13846,N_13474,N_13682);
nor U13847 (N_13847,N_13249,N_13744);
and U13848 (N_13848,N_13589,N_13798);
xnor U13849 (N_13849,N_13423,N_13235);
xnor U13850 (N_13850,N_13710,N_13371);
and U13851 (N_13851,N_13765,N_13225);
or U13852 (N_13852,N_13797,N_13667);
nand U13853 (N_13853,N_13329,N_13616);
and U13854 (N_13854,N_13748,N_13278);
and U13855 (N_13855,N_13640,N_13566);
and U13856 (N_13856,N_13487,N_13373);
and U13857 (N_13857,N_13594,N_13240);
nand U13858 (N_13858,N_13439,N_13307);
and U13859 (N_13859,N_13202,N_13524);
nand U13860 (N_13860,N_13789,N_13283);
or U13861 (N_13861,N_13648,N_13315);
xor U13862 (N_13862,N_13761,N_13752);
xnor U13863 (N_13863,N_13579,N_13715);
xnor U13864 (N_13864,N_13291,N_13749);
or U13865 (N_13865,N_13611,N_13591);
and U13866 (N_13866,N_13649,N_13669);
or U13867 (N_13867,N_13303,N_13298);
nor U13868 (N_13868,N_13754,N_13517);
xor U13869 (N_13869,N_13720,N_13345);
nand U13870 (N_13870,N_13295,N_13446);
or U13871 (N_13871,N_13774,N_13645);
xnor U13872 (N_13872,N_13721,N_13275);
nand U13873 (N_13873,N_13458,N_13217);
nand U13874 (N_13874,N_13334,N_13730);
nor U13875 (N_13875,N_13523,N_13701);
and U13876 (N_13876,N_13526,N_13273);
nand U13877 (N_13877,N_13515,N_13753);
nand U13878 (N_13878,N_13638,N_13301);
or U13879 (N_13879,N_13646,N_13532);
and U13880 (N_13880,N_13585,N_13799);
xor U13881 (N_13881,N_13673,N_13431);
or U13882 (N_13882,N_13660,N_13537);
xor U13883 (N_13883,N_13758,N_13218);
nor U13884 (N_13884,N_13781,N_13595);
xnor U13885 (N_13885,N_13605,N_13316);
xor U13886 (N_13886,N_13299,N_13704);
nor U13887 (N_13887,N_13507,N_13238);
nand U13888 (N_13888,N_13386,N_13435);
and U13889 (N_13889,N_13339,N_13466);
and U13890 (N_13890,N_13557,N_13492);
nand U13891 (N_13891,N_13684,N_13639);
xor U13892 (N_13892,N_13571,N_13499);
nand U13893 (N_13893,N_13775,N_13784);
nand U13894 (N_13894,N_13689,N_13508);
or U13895 (N_13895,N_13450,N_13313);
nor U13896 (N_13896,N_13272,N_13501);
nand U13897 (N_13897,N_13709,N_13751);
and U13898 (N_13898,N_13205,N_13405);
nor U13899 (N_13899,N_13569,N_13747);
and U13900 (N_13900,N_13424,N_13548);
nor U13901 (N_13901,N_13256,N_13552);
nand U13902 (N_13902,N_13764,N_13471);
nand U13903 (N_13903,N_13229,N_13766);
nand U13904 (N_13904,N_13464,N_13521);
nand U13905 (N_13905,N_13743,N_13592);
xor U13906 (N_13906,N_13539,N_13637);
or U13907 (N_13907,N_13641,N_13227);
nand U13908 (N_13908,N_13323,N_13534);
and U13909 (N_13909,N_13705,N_13578);
and U13910 (N_13910,N_13232,N_13707);
xnor U13911 (N_13911,N_13263,N_13378);
xor U13912 (N_13912,N_13491,N_13628);
nand U13913 (N_13913,N_13488,N_13538);
nand U13914 (N_13914,N_13281,N_13399);
nor U13915 (N_13915,N_13770,N_13265);
xor U13916 (N_13916,N_13456,N_13382);
or U13917 (N_13917,N_13654,N_13426);
and U13918 (N_13918,N_13652,N_13357);
nor U13919 (N_13919,N_13259,N_13261);
and U13920 (N_13920,N_13237,N_13727);
nor U13921 (N_13921,N_13580,N_13411);
nand U13922 (N_13922,N_13732,N_13433);
and U13923 (N_13923,N_13516,N_13664);
nor U13924 (N_13924,N_13783,N_13676);
nand U13925 (N_13925,N_13497,N_13713);
and U13926 (N_13926,N_13465,N_13416);
xnor U13927 (N_13927,N_13742,N_13477);
nand U13928 (N_13928,N_13476,N_13584);
xnor U13929 (N_13929,N_13531,N_13420);
nand U13930 (N_13930,N_13342,N_13494);
nor U13931 (N_13931,N_13262,N_13651);
nor U13932 (N_13932,N_13672,N_13771);
or U13933 (N_13933,N_13250,N_13398);
and U13934 (N_13934,N_13428,N_13658);
nor U13935 (N_13935,N_13258,N_13596);
nor U13936 (N_13936,N_13502,N_13642);
or U13937 (N_13937,N_13247,N_13740);
and U13938 (N_13938,N_13773,N_13485);
nor U13939 (N_13939,N_13230,N_13305);
or U13940 (N_13940,N_13274,N_13452);
nand U13941 (N_13941,N_13410,N_13777);
xnor U13942 (N_13942,N_13455,N_13483);
or U13943 (N_13943,N_13436,N_13304);
and U13944 (N_13944,N_13785,N_13677);
nand U13945 (N_13945,N_13687,N_13757);
xnor U13946 (N_13946,N_13372,N_13680);
and U13947 (N_13947,N_13542,N_13255);
and U13948 (N_13948,N_13312,N_13422);
nand U13949 (N_13949,N_13208,N_13468);
or U13950 (N_13950,N_13500,N_13735);
nor U13951 (N_13951,N_13581,N_13791);
or U13952 (N_13952,N_13327,N_13769);
nor U13953 (N_13953,N_13319,N_13630);
nand U13954 (N_13954,N_13467,N_13267);
xnor U13955 (N_13955,N_13318,N_13354);
xnor U13956 (N_13956,N_13478,N_13564);
xnor U13957 (N_13957,N_13506,N_13383);
nand U13958 (N_13958,N_13599,N_13454);
nor U13959 (N_13959,N_13795,N_13527);
nor U13960 (N_13960,N_13414,N_13320);
nand U13961 (N_13961,N_13490,N_13724);
or U13962 (N_13962,N_13586,N_13310);
nand U13963 (N_13963,N_13583,N_13700);
or U13964 (N_13964,N_13463,N_13608);
or U13965 (N_13965,N_13214,N_13385);
nand U13966 (N_13966,N_13543,N_13519);
and U13967 (N_13967,N_13694,N_13317);
nor U13968 (N_13968,N_13553,N_13504);
xnor U13969 (N_13969,N_13448,N_13377);
nor U13970 (N_13970,N_13438,N_13341);
and U13971 (N_13971,N_13200,N_13201);
and U13972 (N_13972,N_13550,N_13413);
or U13973 (N_13973,N_13796,N_13400);
xnor U13974 (N_13974,N_13577,N_13535);
xor U13975 (N_13975,N_13615,N_13391);
xor U13976 (N_13976,N_13551,N_13302);
or U13977 (N_13977,N_13509,N_13620);
and U13978 (N_13978,N_13792,N_13244);
nor U13979 (N_13979,N_13659,N_13560);
nand U13980 (N_13980,N_13325,N_13279);
xor U13981 (N_13981,N_13559,N_13292);
nor U13982 (N_13982,N_13359,N_13212);
or U13983 (N_13983,N_13696,N_13788);
and U13984 (N_13984,N_13418,N_13290);
nand U13985 (N_13985,N_13253,N_13215);
or U13986 (N_13986,N_13239,N_13606);
xnor U13987 (N_13987,N_13368,N_13482);
or U13988 (N_13988,N_13350,N_13525);
nor U13989 (N_13989,N_13496,N_13486);
or U13990 (N_13990,N_13442,N_13461);
nand U13991 (N_13991,N_13759,N_13309);
and U13992 (N_13992,N_13662,N_13376);
or U13993 (N_13993,N_13293,N_13697);
nor U13994 (N_13994,N_13437,N_13495);
xor U13995 (N_13995,N_13333,N_13216);
nor U13996 (N_13996,N_13306,N_13600);
nand U13997 (N_13997,N_13663,N_13364);
nor U13998 (N_13998,N_13481,N_13503);
xor U13999 (N_13999,N_13282,N_13425);
nor U14000 (N_14000,N_13546,N_13794);
nand U14001 (N_14001,N_13219,N_13270);
or U14002 (N_14002,N_13344,N_13349);
or U14003 (N_14003,N_13441,N_13587);
nand U14004 (N_14004,N_13598,N_13204);
nand U14005 (N_14005,N_13653,N_13631);
or U14006 (N_14006,N_13451,N_13343);
or U14007 (N_14007,N_13346,N_13311);
or U14008 (N_14008,N_13716,N_13280);
xnor U14009 (N_14009,N_13593,N_13409);
xor U14010 (N_14010,N_13324,N_13787);
or U14011 (N_14011,N_13228,N_13636);
and U14012 (N_14012,N_13288,N_13417);
nor U14013 (N_14013,N_13489,N_13755);
xnor U14014 (N_14014,N_13655,N_13207);
xor U14015 (N_14015,N_13260,N_13220);
xor U14016 (N_14016,N_13574,N_13241);
or U14017 (N_14017,N_13609,N_13528);
or U14018 (N_14018,N_13702,N_13624);
nor U14019 (N_14019,N_13470,N_13522);
xor U14020 (N_14020,N_13264,N_13612);
or U14021 (N_14021,N_13686,N_13518);
xor U14022 (N_14022,N_13403,N_13392);
or U14023 (N_14023,N_13603,N_13665);
and U14024 (N_14024,N_13297,N_13374);
xor U14025 (N_14025,N_13778,N_13443);
nor U14026 (N_14026,N_13271,N_13296);
and U14027 (N_14027,N_13394,N_13625);
xnor U14028 (N_14028,N_13390,N_13530);
xor U14029 (N_14029,N_13698,N_13321);
nor U14030 (N_14030,N_13555,N_13678);
nor U14031 (N_14031,N_13243,N_13268);
or U14032 (N_14032,N_13556,N_13381);
nor U14033 (N_14033,N_13445,N_13726);
xnor U14034 (N_14034,N_13286,N_13375);
or U14035 (N_14035,N_13562,N_13627);
nand U14036 (N_14036,N_13252,N_13331);
or U14037 (N_14037,N_13337,N_13643);
nand U14038 (N_14038,N_13573,N_13635);
and U14039 (N_14039,N_13352,N_13460);
nor U14040 (N_14040,N_13691,N_13209);
xnor U14041 (N_14041,N_13335,N_13607);
nor U14042 (N_14042,N_13447,N_13565);
nor U14043 (N_14043,N_13725,N_13472);
and U14044 (N_14044,N_13457,N_13326);
nand U14045 (N_14045,N_13479,N_13340);
xor U14046 (N_14046,N_13622,N_13484);
and U14047 (N_14047,N_13613,N_13412);
xor U14048 (N_14048,N_13407,N_13693);
nand U14049 (N_14049,N_13671,N_13427);
nor U14050 (N_14050,N_13351,N_13421);
nor U14051 (N_14051,N_13514,N_13388);
xnor U14052 (N_14052,N_13277,N_13440);
or U14053 (N_14053,N_13762,N_13714);
xor U14054 (N_14054,N_13750,N_13670);
nand U14055 (N_14055,N_13610,N_13379);
nor U14056 (N_14056,N_13210,N_13473);
nand U14057 (N_14057,N_13614,N_13545);
and U14058 (N_14058,N_13287,N_13763);
or U14059 (N_14059,N_13731,N_13475);
xnor U14060 (N_14060,N_13402,N_13688);
nor U14061 (N_14061,N_13520,N_13717);
xnor U14062 (N_14062,N_13647,N_13568);
nor U14063 (N_14063,N_13257,N_13563);
xnor U14064 (N_14064,N_13692,N_13728);
and U14065 (N_14065,N_13575,N_13444);
or U14066 (N_14066,N_13251,N_13511);
and U14067 (N_14067,N_13211,N_13408);
nor U14068 (N_14068,N_13733,N_13544);
and U14069 (N_14069,N_13512,N_13767);
nor U14070 (N_14070,N_13623,N_13355);
or U14071 (N_14071,N_13588,N_13745);
nor U14072 (N_14072,N_13780,N_13706);
nor U14073 (N_14073,N_13234,N_13404);
or U14074 (N_14074,N_13695,N_13363);
or U14075 (N_14075,N_13248,N_13505);
nor U14076 (N_14076,N_13245,N_13396);
nor U14077 (N_14077,N_13738,N_13231);
or U14078 (N_14078,N_13223,N_13685);
or U14079 (N_14079,N_13572,N_13498);
and U14080 (N_14080,N_13330,N_13347);
xor U14081 (N_14081,N_13675,N_13549);
xnor U14082 (N_14082,N_13242,N_13756);
nand U14083 (N_14083,N_13332,N_13393);
or U14084 (N_14084,N_13632,N_13790);
and U14085 (N_14085,N_13601,N_13285);
nand U14086 (N_14086,N_13221,N_13370);
and U14087 (N_14087,N_13510,N_13469);
or U14088 (N_14088,N_13741,N_13533);
nand U14089 (N_14089,N_13666,N_13779);
nand U14090 (N_14090,N_13729,N_13353);
nand U14091 (N_14091,N_13618,N_13722);
or U14092 (N_14092,N_13558,N_13462);
or U14093 (N_14093,N_13703,N_13617);
or U14094 (N_14094,N_13626,N_13300);
xor U14095 (N_14095,N_13360,N_13226);
xnor U14096 (N_14096,N_13590,N_13699);
or U14097 (N_14097,N_13621,N_13387);
or U14098 (N_14098,N_13668,N_13690);
or U14099 (N_14099,N_13348,N_13597);
nand U14100 (N_14100,N_13750,N_13710);
and U14101 (N_14101,N_13234,N_13212);
or U14102 (N_14102,N_13490,N_13756);
nand U14103 (N_14103,N_13246,N_13310);
nand U14104 (N_14104,N_13489,N_13798);
xnor U14105 (N_14105,N_13492,N_13420);
nor U14106 (N_14106,N_13259,N_13415);
xnor U14107 (N_14107,N_13463,N_13358);
nor U14108 (N_14108,N_13553,N_13478);
or U14109 (N_14109,N_13433,N_13527);
or U14110 (N_14110,N_13593,N_13402);
nor U14111 (N_14111,N_13363,N_13248);
nand U14112 (N_14112,N_13483,N_13670);
or U14113 (N_14113,N_13424,N_13642);
and U14114 (N_14114,N_13797,N_13663);
nand U14115 (N_14115,N_13763,N_13638);
nor U14116 (N_14116,N_13200,N_13536);
nand U14117 (N_14117,N_13610,N_13210);
nand U14118 (N_14118,N_13610,N_13565);
xor U14119 (N_14119,N_13686,N_13788);
and U14120 (N_14120,N_13739,N_13371);
xnor U14121 (N_14121,N_13282,N_13447);
xnor U14122 (N_14122,N_13683,N_13630);
nor U14123 (N_14123,N_13306,N_13244);
nor U14124 (N_14124,N_13454,N_13340);
xor U14125 (N_14125,N_13694,N_13682);
nor U14126 (N_14126,N_13757,N_13243);
nand U14127 (N_14127,N_13261,N_13599);
xnor U14128 (N_14128,N_13246,N_13550);
nor U14129 (N_14129,N_13433,N_13712);
or U14130 (N_14130,N_13640,N_13646);
or U14131 (N_14131,N_13558,N_13699);
or U14132 (N_14132,N_13597,N_13314);
and U14133 (N_14133,N_13352,N_13316);
xor U14134 (N_14134,N_13645,N_13407);
nand U14135 (N_14135,N_13336,N_13421);
nor U14136 (N_14136,N_13714,N_13570);
nand U14137 (N_14137,N_13779,N_13394);
nor U14138 (N_14138,N_13248,N_13244);
nor U14139 (N_14139,N_13323,N_13672);
or U14140 (N_14140,N_13599,N_13587);
nor U14141 (N_14141,N_13218,N_13383);
nand U14142 (N_14142,N_13275,N_13621);
and U14143 (N_14143,N_13653,N_13323);
xnor U14144 (N_14144,N_13629,N_13438);
and U14145 (N_14145,N_13350,N_13497);
nand U14146 (N_14146,N_13563,N_13360);
or U14147 (N_14147,N_13334,N_13515);
nand U14148 (N_14148,N_13279,N_13433);
and U14149 (N_14149,N_13635,N_13600);
and U14150 (N_14150,N_13607,N_13263);
nor U14151 (N_14151,N_13706,N_13592);
nor U14152 (N_14152,N_13344,N_13497);
xnor U14153 (N_14153,N_13695,N_13252);
xnor U14154 (N_14154,N_13247,N_13616);
or U14155 (N_14155,N_13414,N_13309);
or U14156 (N_14156,N_13246,N_13230);
nand U14157 (N_14157,N_13225,N_13376);
and U14158 (N_14158,N_13282,N_13305);
nand U14159 (N_14159,N_13382,N_13395);
and U14160 (N_14160,N_13488,N_13285);
or U14161 (N_14161,N_13744,N_13518);
xnor U14162 (N_14162,N_13701,N_13789);
or U14163 (N_14163,N_13607,N_13344);
and U14164 (N_14164,N_13389,N_13695);
and U14165 (N_14165,N_13576,N_13617);
nand U14166 (N_14166,N_13624,N_13254);
nor U14167 (N_14167,N_13551,N_13614);
xor U14168 (N_14168,N_13318,N_13733);
nor U14169 (N_14169,N_13313,N_13293);
nand U14170 (N_14170,N_13261,N_13653);
nand U14171 (N_14171,N_13453,N_13254);
or U14172 (N_14172,N_13784,N_13674);
nor U14173 (N_14173,N_13405,N_13353);
or U14174 (N_14174,N_13321,N_13348);
or U14175 (N_14175,N_13493,N_13738);
nand U14176 (N_14176,N_13209,N_13392);
nor U14177 (N_14177,N_13273,N_13551);
and U14178 (N_14178,N_13215,N_13582);
and U14179 (N_14179,N_13496,N_13612);
xnor U14180 (N_14180,N_13546,N_13368);
nor U14181 (N_14181,N_13606,N_13774);
nand U14182 (N_14182,N_13367,N_13747);
nand U14183 (N_14183,N_13612,N_13747);
nor U14184 (N_14184,N_13254,N_13431);
and U14185 (N_14185,N_13775,N_13647);
and U14186 (N_14186,N_13353,N_13385);
nor U14187 (N_14187,N_13275,N_13447);
xnor U14188 (N_14188,N_13629,N_13634);
and U14189 (N_14189,N_13791,N_13482);
nor U14190 (N_14190,N_13512,N_13295);
or U14191 (N_14191,N_13293,N_13786);
and U14192 (N_14192,N_13776,N_13304);
and U14193 (N_14193,N_13711,N_13489);
nand U14194 (N_14194,N_13220,N_13695);
nor U14195 (N_14195,N_13757,N_13525);
and U14196 (N_14196,N_13410,N_13589);
nand U14197 (N_14197,N_13479,N_13360);
xnor U14198 (N_14198,N_13576,N_13218);
nor U14199 (N_14199,N_13355,N_13394);
and U14200 (N_14200,N_13499,N_13784);
nor U14201 (N_14201,N_13658,N_13213);
and U14202 (N_14202,N_13277,N_13597);
or U14203 (N_14203,N_13752,N_13452);
xor U14204 (N_14204,N_13762,N_13499);
nor U14205 (N_14205,N_13621,N_13749);
nor U14206 (N_14206,N_13685,N_13222);
and U14207 (N_14207,N_13539,N_13735);
and U14208 (N_14208,N_13714,N_13300);
or U14209 (N_14209,N_13266,N_13760);
xnor U14210 (N_14210,N_13646,N_13748);
and U14211 (N_14211,N_13442,N_13575);
and U14212 (N_14212,N_13252,N_13780);
xor U14213 (N_14213,N_13484,N_13676);
or U14214 (N_14214,N_13543,N_13362);
and U14215 (N_14215,N_13746,N_13556);
and U14216 (N_14216,N_13706,N_13356);
or U14217 (N_14217,N_13483,N_13423);
nand U14218 (N_14218,N_13628,N_13221);
nand U14219 (N_14219,N_13768,N_13361);
xor U14220 (N_14220,N_13472,N_13712);
nor U14221 (N_14221,N_13750,N_13693);
and U14222 (N_14222,N_13334,N_13202);
nand U14223 (N_14223,N_13670,N_13225);
and U14224 (N_14224,N_13790,N_13513);
or U14225 (N_14225,N_13326,N_13597);
or U14226 (N_14226,N_13641,N_13519);
xor U14227 (N_14227,N_13260,N_13709);
and U14228 (N_14228,N_13585,N_13546);
or U14229 (N_14229,N_13428,N_13557);
or U14230 (N_14230,N_13214,N_13663);
nor U14231 (N_14231,N_13342,N_13408);
or U14232 (N_14232,N_13475,N_13386);
xor U14233 (N_14233,N_13237,N_13574);
or U14234 (N_14234,N_13740,N_13298);
and U14235 (N_14235,N_13316,N_13493);
nand U14236 (N_14236,N_13522,N_13666);
nand U14237 (N_14237,N_13654,N_13667);
and U14238 (N_14238,N_13688,N_13745);
xor U14239 (N_14239,N_13486,N_13674);
and U14240 (N_14240,N_13279,N_13683);
and U14241 (N_14241,N_13635,N_13507);
nand U14242 (N_14242,N_13402,N_13796);
or U14243 (N_14243,N_13270,N_13793);
xnor U14244 (N_14244,N_13537,N_13386);
xor U14245 (N_14245,N_13482,N_13715);
xor U14246 (N_14246,N_13315,N_13530);
nand U14247 (N_14247,N_13262,N_13590);
or U14248 (N_14248,N_13670,N_13788);
xnor U14249 (N_14249,N_13539,N_13760);
and U14250 (N_14250,N_13399,N_13361);
nand U14251 (N_14251,N_13514,N_13233);
and U14252 (N_14252,N_13712,N_13721);
nand U14253 (N_14253,N_13612,N_13379);
or U14254 (N_14254,N_13483,N_13565);
nand U14255 (N_14255,N_13367,N_13534);
and U14256 (N_14256,N_13509,N_13534);
xnor U14257 (N_14257,N_13421,N_13696);
nor U14258 (N_14258,N_13404,N_13659);
xor U14259 (N_14259,N_13644,N_13284);
or U14260 (N_14260,N_13773,N_13396);
nor U14261 (N_14261,N_13250,N_13617);
nand U14262 (N_14262,N_13306,N_13259);
nand U14263 (N_14263,N_13608,N_13390);
and U14264 (N_14264,N_13713,N_13299);
or U14265 (N_14265,N_13747,N_13289);
xnor U14266 (N_14266,N_13330,N_13621);
or U14267 (N_14267,N_13750,N_13339);
nor U14268 (N_14268,N_13539,N_13442);
nand U14269 (N_14269,N_13661,N_13731);
nand U14270 (N_14270,N_13400,N_13629);
nand U14271 (N_14271,N_13787,N_13724);
nand U14272 (N_14272,N_13607,N_13546);
and U14273 (N_14273,N_13356,N_13777);
and U14274 (N_14274,N_13262,N_13648);
nand U14275 (N_14275,N_13594,N_13203);
nand U14276 (N_14276,N_13687,N_13357);
nand U14277 (N_14277,N_13271,N_13407);
nor U14278 (N_14278,N_13444,N_13351);
nor U14279 (N_14279,N_13421,N_13238);
xor U14280 (N_14280,N_13710,N_13358);
nand U14281 (N_14281,N_13327,N_13628);
nand U14282 (N_14282,N_13627,N_13488);
xnor U14283 (N_14283,N_13688,N_13682);
nor U14284 (N_14284,N_13294,N_13675);
xnor U14285 (N_14285,N_13763,N_13561);
and U14286 (N_14286,N_13356,N_13600);
xnor U14287 (N_14287,N_13433,N_13285);
nor U14288 (N_14288,N_13392,N_13510);
nor U14289 (N_14289,N_13359,N_13392);
and U14290 (N_14290,N_13514,N_13236);
nand U14291 (N_14291,N_13416,N_13256);
or U14292 (N_14292,N_13394,N_13685);
nand U14293 (N_14293,N_13221,N_13737);
and U14294 (N_14294,N_13466,N_13494);
nor U14295 (N_14295,N_13225,N_13464);
or U14296 (N_14296,N_13633,N_13318);
and U14297 (N_14297,N_13203,N_13316);
xor U14298 (N_14298,N_13751,N_13785);
nor U14299 (N_14299,N_13562,N_13386);
nor U14300 (N_14300,N_13592,N_13544);
nor U14301 (N_14301,N_13742,N_13495);
xnor U14302 (N_14302,N_13797,N_13580);
nor U14303 (N_14303,N_13379,N_13750);
nor U14304 (N_14304,N_13348,N_13583);
nor U14305 (N_14305,N_13738,N_13716);
or U14306 (N_14306,N_13582,N_13471);
and U14307 (N_14307,N_13641,N_13767);
xnor U14308 (N_14308,N_13615,N_13209);
xor U14309 (N_14309,N_13779,N_13744);
and U14310 (N_14310,N_13583,N_13449);
or U14311 (N_14311,N_13337,N_13640);
nor U14312 (N_14312,N_13651,N_13477);
nand U14313 (N_14313,N_13555,N_13449);
nor U14314 (N_14314,N_13373,N_13412);
xor U14315 (N_14315,N_13726,N_13330);
or U14316 (N_14316,N_13399,N_13690);
nand U14317 (N_14317,N_13703,N_13286);
xnor U14318 (N_14318,N_13397,N_13243);
and U14319 (N_14319,N_13678,N_13794);
or U14320 (N_14320,N_13281,N_13250);
and U14321 (N_14321,N_13598,N_13435);
nand U14322 (N_14322,N_13410,N_13441);
nand U14323 (N_14323,N_13505,N_13652);
or U14324 (N_14324,N_13457,N_13412);
nand U14325 (N_14325,N_13583,N_13487);
xnor U14326 (N_14326,N_13240,N_13499);
xor U14327 (N_14327,N_13404,N_13623);
nand U14328 (N_14328,N_13319,N_13206);
xor U14329 (N_14329,N_13753,N_13780);
nor U14330 (N_14330,N_13438,N_13713);
and U14331 (N_14331,N_13241,N_13566);
nand U14332 (N_14332,N_13590,N_13311);
nor U14333 (N_14333,N_13507,N_13418);
or U14334 (N_14334,N_13778,N_13525);
or U14335 (N_14335,N_13645,N_13643);
nand U14336 (N_14336,N_13609,N_13217);
or U14337 (N_14337,N_13436,N_13698);
or U14338 (N_14338,N_13356,N_13647);
or U14339 (N_14339,N_13679,N_13486);
or U14340 (N_14340,N_13487,N_13469);
or U14341 (N_14341,N_13409,N_13392);
and U14342 (N_14342,N_13453,N_13293);
nand U14343 (N_14343,N_13679,N_13248);
xor U14344 (N_14344,N_13206,N_13507);
nand U14345 (N_14345,N_13480,N_13318);
or U14346 (N_14346,N_13410,N_13432);
or U14347 (N_14347,N_13406,N_13347);
nand U14348 (N_14348,N_13724,N_13451);
nor U14349 (N_14349,N_13271,N_13324);
nand U14350 (N_14350,N_13594,N_13275);
xnor U14351 (N_14351,N_13484,N_13502);
nor U14352 (N_14352,N_13753,N_13200);
nor U14353 (N_14353,N_13418,N_13753);
and U14354 (N_14354,N_13293,N_13306);
and U14355 (N_14355,N_13378,N_13623);
and U14356 (N_14356,N_13649,N_13430);
nor U14357 (N_14357,N_13466,N_13236);
nand U14358 (N_14358,N_13319,N_13628);
nor U14359 (N_14359,N_13417,N_13658);
xor U14360 (N_14360,N_13284,N_13790);
xnor U14361 (N_14361,N_13598,N_13555);
and U14362 (N_14362,N_13721,N_13422);
or U14363 (N_14363,N_13343,N_13402);
nand U14364 (N_14364,N_13751,N_13584);
xor U14365 (N_14365,N_13499,N_13620);
xor U14366 (N_14366,N_13326,N_13689);
xor U14367 (N_14367,N_13421,N_13744);
xnor U14368 (N_14368,N_13360,N_13675);
and U14369 (N_14369,N_13585,N_13619);
nor U14370 (N_14370,N_13626,N_13290);
and U14371 (N_14371,N_13511,N_13269);
nor U14372 (N_14372,N_13383,N_13582);
nor U14373 (N_14373,N_13291,N_13590);
nor U14374 (N_14374,N_13635,N_13603);
nor U14375 (N_14375,N_13489,N_13695);
xor U14376 (N_14376,N_13355,N_13201);
and U14377 (N_14377,N_13428,N_13265);
nor U14378 (N_14378,N_13365,N_13374);
and U14379 (N_14379,N_13738,N_13487);
or U14380 (N_14380,N_13491,N_13773);
nor U14381 (N_14381,N_13774,N_13649);
and U14382 (N_14382,N_13330,N_13624);
or U14383 (N_14383,N_13632,N_13512);
xor U14384 (N_14384,N_13739,N_13594);
and U14385 (N_14385,N_13449,N_13715);
and U14386 (N_14386,N_13512,N_13348);
xor U14387 (N_14387,N_13324,N_13653);
nor U14388 (N_14388,N_13432,N_13527);
and U14389 (N_14389,N_13429,N_13423);
or U14390 (N_14390,N_13326,N_13453);
xor U14391 (N_14391,N_13217,N_13259);
xor U14392 (N_14392,N_13465,N_13760);
nand U14393 (N_14393,N_13319,N_13512);
xnor U14394 (N_14394,N_13366,N_13568);
or U14395 (N_14395,N_13412,N_13238);
nor U14396 (N_14396,N_13620,N_13782);
nor U14397 (N_14397,N_13632,N_13534);
and U14398 (N_14398,N_13200,N_13575);
and U14399 (N_14399,N_13383,N_13394);
xnor U14400 (N_14400,N_13854,N_14275);
xnor U14401 (N_14401,N_14272,N_14266);
or U14402 (N_14402,N_13839,N_13843);
nand U14403 (N_14403,N_14299,N_14186);
nand U14404 (N_14404,N_14352,N_14317);
xor U14405 (N_14405,N_13960,N_14035);
nor U14406 (N_14406,N_13978,N_13982);
and U14407 (N_14407,N_13884,N_13812);
nor U14408 (N_14408,N_14367,N_13935);
xor U14409 (N_14409,N_13836,N_13904);
or U14410 (N_14410,N_14364,N_14348);
xnor U14411 (N_14411,N_14302,N_13976);
nor U14412 (N_14412,N_14255,N_13828);
xor U14413 (N_14413,N_13965,N_14044);
nand U14414 (N_14414,N_14286,N_14237);
or U14415 (N_14415,N_13838,N_14223);
and U14416 (N_14416,N_14268,N_14087);
nor U14417 (N_14417,N_14165,N_14333);
xor U14418 (N_14418,N_14310,N_14305);
xor U14419 (N_14419,N_13971,N_13847);
or U14420 (N_14420,N_13860,N_14030);
nand U14421 (N_14421,N_14289,N_14207);
and U14422 (N_14422,N_14105,N_13887);
and U14423 (N_14423,N_13820,N_14011);
or U14424 (N_14424,N_13996,N_13888);
and U14425 (N_14425,N_13802,N_13808);
nor U14426 (N_14426,N_14171,N_14216);
or U14427 (N_14427,N_14218,N_14159);
xnor U14428 (N_14428,N_13878,N_13925);
and U14429 (N_14429,N_14196,N_14101);
nand U14430 (N_14430,N_14325,N_13941);
nor U14431 (N_14431,N_14270,N_14227);
xor U14432 (N_14432,N_14148,N_14076);
and U14433 (N_14433,N_14180,N_14215);
xor U14434 (N_14434,N_14194,N_14341);
nor U14435 (N_14435,N_14066,N_14259);
xnor U14436 (N_14436,N_14345,N_14031);
and U14437 (N_14437,N_14205,N_14059);
and U14438 (N_14438,N_13892,N_14058);
nor U14439 (N_14439,N_14130,N_14175);
nor U14440 (N_14440,N_14151,N_14383);
nand U14441 (N_14441,N_13988,N_13898);
or U14442 (N_14442,N_14269,N_14250);
and U14443 (N_14443,N_13848,N_14306);
or U14444 (N_14444,N_14154,N_14274);
or U14445 (N_14445,N_14106,N_14176);
or U14446 (N_14446,N_14129,N_14354);
xnor U14447 (N_14447,N_14150,N_14397);
xor U14448 (N_14448,N_13818,N_14075);
and U14449 (N_14449,N_13910,N_14070);
nand U14450 (N_14450,N_14022,N_14096);
or U14451 (N_14451,N_14251,N_14208);
nand U14452 (N_14452,N_13852,N_14220);
and U14453 (N_14453,N_13856,N_14261);
nand U14454 (N_14454,N_14100,N_14376);
or U14455 (N_14455,N_13939,N_13950);
xor U14456 (N_14456,N_13855,N_14026);
nand U14457 (N_14457,N_13929,N_14012);
or U14458 (N_14458,N_14265,N_14188);
nand U14459 (N_14459,N_13918,N_13803);
nor U14460 (N_14460,N_14143,N_14173);
or U14461 (N_14461,N_14245,N_13917);
nor U14462 (N_14462,N_14353,N_14189);
nor U14463 (N_14463,N_14170,N_13926);
nor U14464 (N_14464,N_14371,N_14000);
nor U14465 (N_14465,N_13846,N_14002);
nor U14466 (N_14466,N_14363,N_13851);
xnor U14467 (N_14467,N_14224,N_14343);
nor U14468 (N_14468,N_14004,N_13810);
nor U14469 (N_14469,N_14377,N_14280);
and U14470 (N_14470,N_14273,N_14051);
nor U14471 (N_14471,N_13825,N_14036);
nand U14472 (N_14472,N_14077,N_14115);
and U14473 (N_14473,N_14267,N_14212);
and U14474 (N_14474,N_14217,N_14158);
or U14475 (N_14475,N_14140,N_13930);
nor U14476 (N_14476,N_14128,N_14144);
and U14477 (N_14477,N_14249,N_14321);
or U14478 (N_14478,N_14332,N_14262);
and U14479 (N_14479,N_14329,N_13977);
nor U14480 (N_14480,N_13850,N_14193);
xor U14481 (N_14481,N_14136,N_14055);
and U14482 (N_14482,N_13864,N_14240);
and U14483 (N_14483,N_14396,N_14389);
and U14484 (N_14484,N_14198,N_13893);
nor U14485 (N_14485,N_14213,N_14290);
nor U14486 (N_14486,N_13897,N_14112);
or U14487 (N_14487,N_14349,N_14256);
nor U14488 (N_14488,N_14013,N_14358);
nand U14489 (N_14489,N_14088,N_13924);
xor U14490 (N_14490,N_14393,N_14362);
xor U14491 (N_14491,N_14038,N_14132);
xor U14492 (N_14492,N_14162,N_14357);
nor U14493 (N_14493,N_13829,N_14247);
nor U14494 (N_14494,N_13958,N_14328);
nand U14495 (N_14495,N_14190,N_14001);
or U14496 (N_14496,N_13841,N_14387);
xor U14497 (N_14497,N_14327,N_13895);
nand U14498 (N_14498,N_14334,N_14123);
or U14499 (N_14499,N_14338,N_14201);
nand U14500 (N_14500,N_13991,N_13814);
or U14501 (N_14501,N_14127,N_14174);
nand U14502 (N_14502,N_13928,N_14009);
and U14503 (N_14503,N_13949,N_14307);
or U14504 (N_14504,N_14164,N_13948);
and U14505 (N_14505,N_14089,N_14177);
nand U14506 (N_14506,N_14301,N_13819);
or U14507 (N_14507,N_14390,N_14394);
nor U14508 (N_14508,N_13908,N_14119);
xnor U14509 (N_14509,N_13936,N_14337);
nand U14510 (N_14510,N_13900,N_13877);
or U14511 (N_14511,N_14388,N_13832);
and U14512 (N_14512,N_14392,N_14064);
nor U14513 (N_14513,N_14108,N_14039);
or U14514 (N_14514,N_14222,N_14258);
nor U14515 (N_14515,N_14054,N_14257);
or U14516 (N_14516,N_13845,N_13871);
or U14517 (N_14517,N_14169,N_14024);
or U14518 (N_14518,N_14368,N_14326);
or U14519 (N_14519,N_14010,N_14291);
or U14520 (N_14520,N_14241,N_14008);
nor U14521 (N_14521,N_14084,N_13883);
or U14522 (N_14522,N_14060,N_14080);
nand U14523 (N_14523,N_14082,N_14003);
nor U14524 (N_14524,N_13914,N_14342);
nor U14525 (N_14525,N_14116,N_14202);
or U14526 (N_14526,N_13987,N_13901);
nand U14527 (N_14527,N_14356,N_13959);
and U14528 (N_14528,N_14372,N_13955);
nor U14529 (N_14529,N_14233,N_14293);
nand U14530 (N_14530,N_13946,N_13970);
or U14531 (N_14531,N_13980,N_14139);
xor U14532 (N_14532,N_14335,N_14316);
or U14533 (N_14533,N_13986,N_13922);
nand U14534 (N_14534,N_14191,N_14228);
nor U14535 (N_14535,N_14146,N_13801);
xor U14536 (N_14536,N_14179,N_13992);
or U14537 (N_14537,N_14133,N_14381);
nand U14538 (N_14538,N_13826,N_13875);
xor U14539 (N_14539,N_14067,N_14157);
and U14540 (N_14540,N_14141,N_14163);
xor U14541 (N_14541,N_14303,N_14199);
nor U14542 (N_14542,N_14029,N_14018);
xnor U14543 (N_14543,N_14056,N_14073);
xor U14544 (N_14544,N_14373,N_13861);
nand U14545 (N_14545,N_14086,N_13902);
nor U14546 (N_14546,N_14279,N_14244);
and U14547 (N_14547,N_14017,N_14184);
nand U14548 (N_14548,N_14187,N_13868);
or U14549 (N_14549,N_13984,N_14296);
xor U14550 (N_14550,N_14043,N_14072);
xnor U14551 (N_14551,N_14308,N_14069);
nand U14552 (N_14552,N_13966,N_13805);
nand U14553 (N_14553,N_14045,N_14049);
or U14554 (N_14554,N_14344,N_13994);
nand U14555 (N_14555,N_14048,N_13804);
xor U14556 (N_14556,N_14324,N_14318);
nand U14557 (N_14557,N_14297,N_13811);
and U14558 (N_14558,N_14350,N_13870);
or U14559 (N_14559,N_13969,N_14203);
and U14560 (N_14560,N_14160,N_14037);
or U14561 (N_14561,N_13867,N_13920);
and U14562 (N_14562,N_13889,N_14107);
and U14563 (N_14563,N_14135,N_14330);
nand U14564 (N_14564,N_14221,N_13858);
nand U14565 (N_14565,N_13849,N_13822);
xnor U14566 (N_14566,N_13940,N_14091);
nand U14567 (N_14567,N_13815,N_14040);
xor U14568 (N_14568,N_13831,N_14379);
nand U14569 (N_14569,N_14053,N_14346);
nand U14570 (N_14570,N_14034,N_14032);
and U14571 (N_14571,N_14102,N_13899);
or U14572 (N_14572,N_13943,N_14355);
and U14573 (N_14573,N_14278,N_14230);
nor U14574 (N_14574,N_14068,N_13800);
nand U14575 (N_14575,N_14282,N_13891);
or U14576 (N_14576,N_13830,N_14122);
and U14577 (N_14577,N_13905,N_13954);
or U14578 (N_14578,N_14020,N_13885);
nor U14579 (N_14579,N_13972,N_13913);
nand U14580 (N_14580,N_14145,N_14090);
or U14581 (N_14581,N_13859,N_14021);
nor U14582 (N_14582,N_14281,N_13981);
nand U14583 (N_14583,N_13821,N_14097);
xnor U14584 (N_14584,N_14178,N_14260);
nor U14585 (N_14585,N_14161,N_13834);
and U14586 (N_14586,N_13837,N_13915);
nor U14587 (N_14587,N_13813,N_13863);
or U14588 (N_14588,N_14225,N_13906);
nand U14589 (N_14589,N_14340,N_14313);
nand U14590 (N_14590,N_14041,N_13975);
or U14591 (N_14591,N_14033,N_13909);
xnor U14592 (N_14592,N_14284,N_14300);
nand U14593 (N_14593,N_13894,N_14374);
and U14594 (N_14594,N_13953,N_14312);
and U14595 (N_14595,N_14085,N_14172);
and U14596 (N_14596,N_14320,N_14098);
nand U14597 (N_14597,N_13962,N_14311);
or U14598 (N_14598,N_14263,N_14126);
nand U14599 (N_14599,N_14071,N_14276);
xor U14600 (N_14600,N_13923,N_14209);
nor U14601 (N_14601,N_14182,N_14234);
xor U14602 (N_14602,N_14147,N_13961);
xnor U14603 (N_14603,N_14375,N_14192);
nor U14604 (N_14604,N_13817,N_13872);
nor U14605 (N_14605,N_13932,N_13934);
nand U14606 (N_14606,N_14398,N_14025);
and U14607 (N_14607,N_14361,N_14226);
xnor U14608 (N_14608,N_14065,N_13879);
or U14609 (N_14609,N_14109,N_14028);
or U14610 (N_14610,N_14314,N_13983);
xor U14611 (N_14611,N_13890,N_14131);
nand U14612 (N_14612,N_14378,N_14219);
or U14613 (N_14613,N_13957,N_14138);
nand U14614 (N_14614,N_13874,N_14078);
nand U14615 (N_14615,N_14246,N_14264);
nor U14616 (N_14616,N_14370,N_13873);
nand U14617 (N_14617,N_14236,N_14210);
nor U14618 (N_14618,N_14079,N_14283);
and U14619 (N_14619,N_14391,N_14351);
xor U14620 (N_14620,N_13945,N_13989);
xor U14621 (N_14621,N_13857,N_14023);
nand U14622 (N_14622,N_14093,N_14197);
and U14623 (N_14623,N_13807,N_13985);
nor U14624 (N_14624,N_14253,N_14235);
xor U14625 (N_14625,N_13880,N_14385);
nor U14626 (N_14626,N_14057,N_13853);
and U14627 (N_14627,N_14063,N_14254);
and U14628 (N_14628,N_14042,N_13921);
or U14629 (N_14629,N_14099,N_14195);
nand U14630 (N_14630,N_13842,N_14319);
nand U14631 (N_14631,N_14395,N_14103);
or U14632 (N_14632,N_13835,N_13881);
xor U14633 (N_14633,N_13916,N_14016);
and U14634 (N_14634,N_14095,N_14366);
xor U14635 (N_14635,N_14336,N_13809);
and U14636 (N_14636,N_13956,N_13806);
xor U14637 (N_14637,N_13907,N_14185);
nor U14638 (N_14638,N_13896,N_13995);
and U14639 (N_14639,N_14114,N_14027);
nor U14640 (N_14640,N_14294,N_13973);
nand U14641 (N_14641,N_13993,N_14200);
and U14642 (N_14642,N_14304,N_13944);
xor U14643 (N_14643,N_13968,N_13974);
nor U14644 (N_14644,N_14214,N_13951);
nand U14645 (N_14645,N_14052,N_14295);
nand U14646 (N_14646,N_14094,N_13903);
nand U14647 (N_14647,N_14238,N_14110);
and U14648 (N_14648,N_14181,N_13979);
and U14649 (N_14649,N_14137,N_13997);
xor U14650 (N_14650,N_13927,N_14322);
xor U14651 (N_14651,N_13827,N_14050);
xor U14652 (N_14652,N_14331,N_14062);
nand U14653 (N_14653,N_13823,N_13947);
xnor U14654 (N_14654,N_13886,N_13866);
xor U14655 (N_14655,N_14339,N_14149);
nor U14656 (N_14656,N_13840,N_14061);
nand U14657 (N_14657,N_14323,N_13869);
nor U14658 (N_14658,N_13816,N_14231);
nor U14659 (N_14659,N_14156,N_14074);
nand U14660 (N_14660,N_13844,N_14229);
nor U14661 (N_14661,N_14285,N_14113);
xnor U14662 (N_14662,N_14347,N_14232);
and U14663 (N_14663,N_14117,N_14252);
xnor U14664 (N_14664,N_14014,N_14183);
or U14665 (N_14665,N_14083,N_14006);
nand U14666 (N_14666,N_14111,N_14047);
and U14667 (N_14667,N_14081,N_13942);
xor U14668 (N_14668,N_14386,N_14019);
nor U14669 (N_14669,N_13862,N_14243);
and U14670 (N_14670,N_13963,N_13938);
xor U14671 (N_14671,N_13937,N_13998);
nand U14672 (N_14672,N_14271,N_13865);
nand U14673 (N_14673,N_14382,N_14292);
and U14674 (N_14674,N_14142,N_14120);
or U14675 (N_14675,N_14015,N_14118);
nor U14676 (N_14676,N_14167,N_14298);
xor U14677 (N_14677,N_14369,N_14005);
and U14678 (N_14678,N_14121,N_14168);
nor U14679 (N_14679,N_14365,N_14359);
nand U14680 (N_14680,N_13933,N_13911);
or U14681 (N_14681,N_14384,N_13882);
nand U14682 (N_14682,N_13964,N_14360);
or U14683 (N_14683,N_14152,N_14309);
or U14684 (N_14684,N_13931,N_14155);
xor U14685 (N_14685,N_14242,N_14315);
xor U14686 (N_14686,N_13912,N_13990);
xnor U14687 (N_14687,N_14166,N_14380);
xnor U14688 (N_14688,N_13833,N_14248);
nand U14689 (N_14689,N_14092,N_14399);
and U14690 (N_14690,N_13999,N_14153);
nor U14691 (N_14691,N_14046,N_14287);
xnor U14692 (N_14692,N_13919,N_14288);
and U14693 (N_14693,N_14007,N_13952);
or U14694 (N_14694,N_13824,N_14125);
or U14695 (N_14695,N_14211,N_13876);
or U14696 (N_14696,N_14206,N_14124);
and U14697 (N_14697,N_14239,N_13967);
or U14698 (N_14698,N_14204,N_14277);
nand U14699 (N_14699,N_14104,N_14134);
or U14700 (N_14700,N_14364,N_13812);
nor U14701 (N_14701,N_13891,N_14303);
or U14702 (N_14702,N_14181,N_13838);
or U14703 (N_14703,N_14062,N_14082);
xor U14704 (N_14704,N_14125,N_13913);
nand U14705 (N_14705,N_14259,N_14043);
and U14706 (N_14706,N_14248,N_14246);
nand U14707 (N_14707,N_14252,N_14046);
xnor U14708 (N_14708,N_13817,N_13873);
and U14709 (N_14709,N_14199,N_13857);
and U14710 (N_14710,N_13882,N_13832);
nand U14711 (N_14711,N_14183,N_14310);
or U14712 (N_14712,N_14196,N_13965);
and U14713 (N_14713,N_14390,N_14103);
nor U14714 (N_14714,N_13875,N_14321);
nor U14715 (N_14715,N_14299,N_14386);
or U14716 (N_14716,N_14311,N_14004);
nor U14717 (N_14717,N_13990,N_14009);
xnor U14718 (N_14718,N_14398,N_14283);
or U14719 (N_14719,N_14079,N_14253);
xnor U14720 (N_14720,N_14092,N_14153);
and U14721 (N_14721,N_13825,N_14293);
nand U14722 (N_14722,N_14282,N_14230);
or U14723 (N_14723,N_14112,N_14350);
nand U14724 (N_14724,N_14244,N_13928);
xor U14725 (N_14725,N_14194,N_14266);
xnor U14726 (N_14726,N_13906,N_13914);
or U14727 (N_14727,N_14259,N_14373);
nor U14728 (N_14728,N_14380,N_14065);
nand U14729 (N_14729,N_13881,N_14018);
nand U14730 (N_14730,N_13817,N_13838);
nand U14731 (N_14731,N_14008,N_14043);
xnor U14732 (N_14732,N_14271,N_13844);
nand U14733 (N_14733,N_14349,N_14236);
xor U14734 (N_14734,N_14081,N_13886);
or U14735 (N_14735,N_13875,N_13969);
and U14736 (N_14736,N_13981,N_14323);
nand U14737 (N_14737,N_14122,N_14054);
xor U14738 (N_14738,N_14047,N_13806);
or U14739 (N_14739,N_14182,N_13952);
nand U14740 (N_14740,N_14126,N_13978);
and U14741 (N_14741,N_14244,N_13980);
xor U14742 (N_14742,N_14101,N_14277);
nand U14743 (N_14743,N_14398,N_14196);
xnor U14744 (N_14744,N_14384,N_13950);
nor U14745 (N_14745,N_14093,N_13815);
xnor U14746 (N_14746,N_14042,N_13834);
nor U14747 (N_14747,N_13946,N_14148);
or U14748 (N_14748,N_13846,N_14158);
xor U14749 (N_14749,N_13896,N_14241);
nor U14750 (N_14750,N_14095,N_14372);
and U14751 (N_14751,N_13853,N_13954);
nor U14752 (N_14752,N_14279,N_13951);
nand U14753 (N_14753,N_13831,N_14304);
nor U14754 (N_14754,N_13855,N_14056);
nand U14755 (N_14755,N_14011,N_14225);
or U14756 (N_14756,N_14077,N_14213);
xnor U14757 (N_14757,N_13866,N_13912);
and U14758 (N_14758,N_13850,N_14369);
xnor U14759 (N_14759,N_14215,N_14285);
xnor U14760 (N_14760,N_13916,N_13802);
or U14761 (N_14761,N_14229,N_14068);
and U14762 (N_14762,N_14113,N_14128);
and U14763 (N_14763,N_14312,N_14217);
nand U14764 (N_14764,N_14121,N_14084);
nor U14765 (N_14765,N_14181,N_13853);
nor U14766 (N_14766,N_14359,N_13961);
nand U14767 (N_14767,N_13865,N_14158);
or U14768 (N_14768,N_14059,N_14363);
and U14769 (N_14769,N_14041,N_13886);
and U14770 (N_14770,N_14171,N_13888);
nand U14771 (N_14771,N_13964,N_14138);
or U14772 (N_14772,N_14302,N_13946);
or U14773 (N_14773,N_14073,N_13899);
or U14774 (N_14774,N_14080,N_13979);
nor U14775 (N_14775,N_13991,N_14178);
nor U14776 (N_14776,N_14141,N_14101);
or U14777 (N_14777,N_13928,N_13939);
or U14778 (N_14778,N_14246,N_14259);
and U14779 (N_14779,N_13870,N_13919);
nor U14780 (N_14780,N_14065,N_14315);
or U14781 (N_14781,N_13953,N_14399);
and U14782 (N_14782,N_14292,N_14162);
xor U14783 (N_14783,N_14292,N_14155);
nand U14784 (N_14784,N_13994,N_14185);
nand U14785 (N_14785,N_14022,N_13871);
and U14786 (N_14786,N_13937,N_14201);
xnor U14787 (N_14787,N_13917,N_14182);
or U14788 (N_14788,N_14278,N_14066);
or U14789 (N_14789,N_14153,N_14016);
and U14790 (N_14790,N_14283,N_14341);
xor U14791 (N_14791,N_14028,N_14265);
xor U14792 (N_14792,N_14044,N_14314);
or U14793 (N_14793,N_14112,N_14046);
xnor U14794 (N_14794,N_14056,N_14279);
nor U14795 (N_14795,N_13931,N_14394);
or U14796 (N_14796,N_14183,N_14328);
nand U14797 (N_14797,N_14268,N_14096);
nand U14798 (N_14798,N_14237,N_14148);
and U14799 (N_14799,N_14035,N_14022);
nor U14800 (N_14800,N_13885,N_14183);
xnor U14801 (N_14801,N_14372,N_14245);
and U14802 (N_14802,N_14138,N_14318);
nand U14803 (N_14803,N_13951,N_14211);
nor U14804 (N_14804,N_13938,N_13946);
or U14805 (N_14805,N_13993,N_13914);
or U14806 (N_14806,N_14283,N_13941);
or U14807 (N_14807,N_14174,N_14327);
and U14808 (N_14808,N_13847,N_14097);
xor U14809 (N_14809,N_13964,N_14329);
nor U14810 (N_14810,N_13887,N_13933);
nand U14811 (N_14811,N_14348,N_13930);
or U14812 (N_14812,N_13800,N_13969);
nor U14813 (N_14813,N_14140,N_14357);
and U14814 (N_14814,N_13996,N_14271);
nand U14815 (N_14815,N_14367,N_14371);
xor U14816 (N_14816,N_14266,N_13853);
and U14817 (N_14817,N_14166,N_13932);
nor U14818 (N_14818,N_14373,N_13934);
and U14819 (N_14819,N_14063,N_14088);
nand U14820 (N_14820,N_14301,N_14343);
nand U14821 (N_14821,N_14203,N_14362);
nand U14822 (N_14822,N_14296,N_14071);
or U14823 (N_14823,N_14177,N_13910);
nor U14824 (N_14824,N_14305,N_14314);
nand U14825 (N_14825,N_14188,N_14023);
and U14826 (N_14826,N_14183,N_14131);
xor U14827 (N_14827,N_13872,N_14091);
and U14828 (N_14828,N_13932,N_14112);
nand U14829 (N_14829,N_13975,N_14255);
nor U14830 (N_14830,N_13801,N_14115);
nand U14831 (N_14831,N_14000,N_14227);
nand U14832 (N_14832,N_14081,N_14135);
nor U14833 (N_14833,N_14024,N_13807);
and U14834 (N_14834,N_14029,N_14019);
nand U14835 (N_14835,N_14076,N_14083);
or U14836 (N_14836,N_14110,N_14008);
nand U14837 (N_14837,N_14166,N_14137);
xor U14838 (N_14838,N_13908,N_14028);
nand U14839 (N_14839,N_14233,N_14360);
xor U14840 (N_14840,N_13878,N_14361);
xor U14841 (N_14841,N_14194,N_13824);
nor U14842 (N_14842,N_13876,N_14023);
nand U14843 (N_14843,N_14041,N_13890);
nor U14844 (N_14844,N_14269,N_14026);
or U14845 (N_14845,N_13996,N_14044);
nor U14846 (N_14846,N_14038,N_14092);
and U14847 (N_14847,N_14078,N_14317);
nor U14848 (N_14848,N_14115,N_14241);
and U14849 (N_14849,N_14098,N_14327);
and U14850 (N_14850,N_14295,N_14004);
and U14851 (N_14851,N_14288,N_14376);
nand U14852 (N_14852,N_14061,N_14350);
nor U14853 (N_14853,N_14256,N_13904);
nor U14854 (N_14854,N_13869,N_13870);
nor U14855 (N_14855,N_13820,N_14299);
nor U14856 (N_14856,N_14037,N_13865);
and U14857 (N_14857,N_14065,N_14063);
and U14858 (N_14858,N_14178,N_13838);
xor U14859 (N_14859,N_13815,N_14159);
and U14860 (N_14860,N_14328,N_13894);
and U14861 (N_14861,N_13839,N_14094);
and U14862 (N_14862,N_13995,N_13974);
or U14863 (N_14863,N_14088,N_14029);
xnor U14864 (N_14864,N_14389,N_14195);
xor U14865 (N_14865,N_13939,N_13803);
nand U14866 (N_14866,N_14222,N_14180);
and U14867 (N_14867,N_14307,N_14005);
and U14868 (N_14868,N_13987,N_13916);
or U14869 (N_14869,N_14068,N_13969);
or U14870 (N_14870,N_14302,N_13814);
and U14871 (N_14871,N_13850,N_14163);
nor U14872 (N_14872,N_14270,N_14394);
and U14873 (N_14873,N_14255,N_14335);
or U14874 (N_14874,N_13936,N_13905);
or U14875 (N_14875,N_13968,N_14243);
and U14876 (N_14876,N_14187,N_14082);
nand U14877 (N_14877,N_13903,N_13971);
and U14878 (N_14878,N_13840,N_13964);
and U14879 (N_14879,N_14276,N_14148);
xor U14880 (N_14880,N_14249,N_14338);
and U14881 (N_14881,N_14356,N_13850);
xor U14882 (N_14882,N_14212,N_13808);
nor U14883 (N_14883,N_14398,N_13917);
nand U14884 (N_14884,N_13872,N_14084);
nand U14885 (N_14885,N_14318,N_14028);
and U14886 (N_14886,N_14225,N_13879);
xor U14887 (N_14887,N_14052,N_13964);
xor U14888 (N_14888,N_14164,N_14214);
or U14889 (N_14889,N_13834,N_14031);
and U14890 (N_14890,N_14254,N_14190);
or U14891 (N_14891,N_14024,N_13914);
and U14892 (N_14892,N_14021,N_14006);
xnor U14893 (N_14893,N_14306,N_14276);
nand U14894 (N_14894,N_13912,N_14040);
nand U14895 (N_14895,N_14283,N_14194);
nand U14896 (N_14896,N_14158,N_14252);
xnor U14897 (N_14897,N_14275,N_14045);
or U14898 (N_14898,N_13896,N_14119);
nand U14899 (N_14899,N_14283,N_13893);
nor U14900 (N_14900,N_14191,N_14193);
xnor U14901 (N_14901,N_14171,N_14021);
and U14902 (N_14902,N_14320,N_14088);
nand U14903 (N_14903,N_14171,N_14117);
nand U14904 (N_14904,N_14047,N_14053);
and U14905 (N_14905,N_13856,N_14018);
xor U14906 (N_14906,N_14163,N_14337);
or U14907 (N_14907,N_13967,N_13948);
and U14908 (N_14908,N_13916,N_14065);
nor U14909 (N_14909,N_14257,N_14170);
xor U14910 (N_14910,N_13999,N_14035);
xnor U14911 (N_14911,N_14362,N_14120);
and U14912 (N_14912,N_14241,N_13801);
xor U14913 (N_14913,N_13998,N_14346);
nor U14914 (N_14914,N_14020,N_14369);
and U14915 (N_14915,N_13844,N_13994);
or U14916 (N_14916,N_14218,N_13803);
and U14917 (N_14917,N_13873,N_14057);
or U14918 (N_14918,N_13807,N_14048);
nand U14919 (N_14919,N_13918,N_14036);
xor U14920 (N_14920,N_14009,N_13924);
and U14921 (N_14921,N_14060,N_14086);
xor U14922 (N_14922,N_14254,N_14082);
and U14923 (N_14923,N_14199,N_14130);
nor U14924 (N_14924,N_14211,N_13804);
and U14925 (N_14925,N_14091,N_14066);
nor U14926 (N_14926,N_14237,N_13822);
and U14927 (N_14927,N_14366,N_14358);
and U14928 (N_14928,N_14138,N_14219);
and U14929 (N_14929,N_14114,N_14358);
nand U14930 (N_14930,N_14192,N_14089);
xor U14931 (N_14931,N_13921,N_14013);
nand U14932 (N_14932,N_14312,N_14151);
or U14933 (N_14933,N_13906,N_14376);
xnor U14934 (N_14934,N_13955,N_14082);
or U14935 (N_14935,N_14298,N_14270);
nor U14936 (N_14936,N_14136,N_13940);
nor U14937 (N_14937,N_13959,N_14132);
nand U14938 (N_14938,N_13967,N_14319);
nand U14939 (N_14939,N_14312,N_13922);
nor U14940 (N_14940,N_13828,N_14305);
nor U14941 (N_14941,N_13944,N_14125);
nor U14942 (N_14942,N_14340,N_14305);
nand U14943 (N_14943,N_13959,N_14260);
xnor U14944 (N_14944,N_14390,N_14277);
and U14945 (N_14945,N_14015,N_14395);
or U14946 (N_14946,N_14286,N_14365);
xnor U14947 (N_14947,N_13806,N_14130);
xor U14948 (N_14948,N_14325,N_14046);
nand U14949 (N_14949,N_14177,N_14080);
or U14950 (N_14950,N_13870,N_13993);
nor U14951 (N_14951,N_13884,N_14301);
and U14952 (N_14952,N_13945,N_13929);
and U14953 (N_14953,N_13955,N_14092);
and U14954 (N_14954,N_14288,N_14041);
xor U14955 (N_14955,N_13880,N_14149);
nor U14956 (N_14956,N_14007,N_14332);
nand U14957 (N_14957,N_14244,N_14009);
xnor U14958 (N_14958,N_13879,N_14123);
and U14959 (N_14959,N_14144,N_13904);
xor U14960 (N_14960,N_13994,N_13996);
nand U14961 (N_14961,N_14153,N_14355);
xnor U14962 (N_14962,N_14319,N_13826);
and U14963 (N_14963,N_14062,N_14146);
nand U14964 (N_14964,N_13959,N_13990);
or U14965 (N_14965,N_14152,N_13889);
and U14966 (N_14966,N_14364,N_13831);
nor U14967 (N_14967,N_13833,N_13979);
or U14968 (N_14968,N_14333,N_14383);
and U14969 (N_14969,N_13957,N_14168);
and U14970 (N_14970,N_14251,N_14045);
nor U14971 (N_14971,N_14282,N_13956);
nand U14972 (N_14972,N_13810,N_13807);
nor U14973 (N_14973,N_14143,N_14078);
xnor U14974 (N_14974,N_14248,N_14079);
xnor U14975 (N_14975,N_14006,N_13954);
nand U14976 (N_14976,N_14191,N_14352);
and U14977 (N_14977,N_14041,N_13991);
nand U14978 (N_14978,N_14201,N_13927);
or U14979 (N_14979,N_14373,N_14139);
nor U14980 (N_14980,N_14290,N_13811);
nand U14981 (N_14981,N_14136,N_14126);
and U14982 (N_14982,N_13836,N_14215);
or U14983 (N_14983,N_14262,N_14054);
or U14984 (N_14984,N_14344,N_13822);
or U14985 (N_14985,N_13934,N_14073);
and U14986 (N_14986,N_14394,N_13901);
and U14987 (N_14987,N_14344,N_14340);
xor U14988 (N_14988,N_14242,N_14257);
and U14989 (N_14989,N_14050,N_14040);
nor U14990 (N_14990,N_14016,N_14297);
xnor U14991 (N_14991,N_14002,N_14367);
and U14992 (N_14992,N_13828,N_13862);
and U14993 (N_14993,N_14372,N_14195);
or U14994 (N_14994,N_14030,N_14007);
or U14995 (N_14995,N_14114,N_14050);
nor U14996 (N_14996,N_14145,N_14255);
and U14997 (N_14997,N_14136,N_14394);
or U14998 (N_14998,N_14296,N_14098);
nand U14999 (N_14999,N_13888,N_14329);
or U15000 (N_15000,N_14819,N_14977);
xnor U15001 (N_15001,N_14452,N_14817);
nand U15002 (N_15002,N_14918,N_14432);
or U15003 (N_15003,N_14881,N_14462);
or U15004 (N_15004,N_14442,N_14764);
and U15005 (N_15005,N_14880,N_14969);
and U15006 (N_15006,N_14847,N_14607);
and U15007 (N_15007,N_14569,N_14448);
nor U15008 (N_15008,N_14699,N_14611);
nand U15009 (N_15009,N_14835,N_14676);
nand U15010 (N_15010,N_14713,N_14470);
nand U15011 (N_15011,N_14736,N_14600);
nor U15012 (N_15012,N_14976,N_14529);
xor U15013 (N_15013,N_14430,N_14993);
and U15014 (N_15014,N_14753,N_14842);
xnor U15015 (N_15015,N_14950,N_14721);
xnor U15016 (N_15016,N_14493,N_14453);
xnor U15017 (N_15017,N_14972,N_14863);
and U15018 (N_15018,N_14514,N_14694);
nor U15019 (N_15019,N_14771,N_14456);
xor U15020 (N_15020,N_14552,N_14719);
nor U15021 (N_15021,N_14733,N_14706);
nor U15022 (N_15022,N_14633,N_14823);
xnor U15023 (N_15023,N_14782,N_14518);
and U15024 (N_15024,N_14587,N_14696);
xnor U15025 (N_15025,N_14579,N_14801);
and U15026 (N_15026,N_14814,N_14886);
xnor U15027 (N_15027,N_14554,N_14659);
nand U15028 (N_15028,N_14454,N_14811);
xor U15029 (N_15029,N_14574,N_14476);
xor U15030 (N_15030,N_14698,N_14471);
and U15031 (N_15031,N_14522,N_14779);
and U15032 (N_15032,N_14562,N_14799);
xnor U15033 (N_15033,N_14517,N_14809);
nor U15034 (N_15034,N_14655,N_14887);
xor U15035 (N_15035,N_14744,N_14491);
and U15036 (N_15036,N_14830,N_14495);
and U15037 (N_15037,N_14509,N_14619);
xor U15038 (N_15038,N_14853,N_14612);
nand U15039 (N_15039,N_14878,N_14555);
nand U15040 (N_15040,N_14741,N_14783);
xor U15041 (N_15041,N_14610,N_14414);
nand U15042 (N_15042,N_14792,N_14730);
xor U15043 (N_15043,N_14685,N_14591);
or U15044 (N_15044,N_14731,N_14982);
xnor U15045 (N_15045,N_14434,N_14979);
or U15046 (N_15046,N_14499,N_14496);
xnor U15047 (N_15047,N_14987,N_14540);
or U15048 (N_15048,N_14994,N_14768);
or U15049 (N_15049,N_14578,N_14488);
and U15050 (N_15050,N_14841,N_14639);
and U15051 (N_15051,N_14505,N_14756);
nand U15052 (N_15052,N_14670,N_14871);
or U15053 (N_15053,N_14983,N_14966);
or U15054 (N_15054,N_14973,N_14464);
or U15055 (N_15055,N_14939,N_14838);
or U15056 (N_15056,N_14766,N_14691);
nand U15057 (N_15057,N_14791,N_14712);
nor U15058 (N_15058,N_14406,N_14455);
nand U15059 (N_15059,N_14752,N_14832);
and U15060 (N_15060,N_14565,N_14582);
or U15061 (N_15061,N_14739,N_14686);
and U15062 (N_15062,N_14946,N_14891);
or U15063 (N_15063,N_14647,N_14537);
xnor U15064 (N_15064,N_14978,N_14511);
xnor U15065 (N_15065,N_14897,N_14772);
nor U15066 (N_15066,N_14483,N_14563);
xor U15067 (N_15067,N_14411,N_14543);
or U15068 (N_15068,N_14703,N_14635);
xnor U15069 (N_15069,N_14457,N_14924);
xor U15070 (N_15070,N_14784,N_14571);
nor U15071 (N_15071,N_14873,N_14447);
xnor U15072 (N_15072,N_14513,N_14861);
nor U15073 (N_15073,N_14560,N_14620);
xnor U15074 (N_15074,N_14777,N_14535);
nor U15075 (N_15075,N_14584,N_14989);
nand U15076 (N_15076,N_14826,N_14849);
xor U15077 (N_15077,N_14931,N_14636);
nor U15078 (N_15078,N_14443,N_14466);
nor U15079 (N_15079,N_14804,N_14996);
nor U15080 (N_15080,N_14967,N_14705);
xor U15081 (N_15081,N_14460,N_14708);
xnor U15082 (N_15082,N_14908,N_14922);
and U15083 (N_15083,N_14604,N_14450);
or U15084 (N_15084,N_14688,N_14890);
nand U15085 (N_15085,N_14629,N_14478);
nand U15086 (N_15086,N_14729,N_14761);
xor U15087 (N_15087,N_14684,N_14742);
xor U15088 (N_15088,N_14843,N_14810);
nor U15089 (N_15089,N_14938,N_14524);
or U15090 (N_15090,N_14410,N_14428);
or U15091 (N_15091,N_14734,N_14762);
xor U15092 (N_15092,N_14913,N_14834);
xnor U15093 (N_15093,N_14767,N_14534);
xnor U15094 (N_15094,N_14479,N_14446);
xor U15095 (N_15095,N_14595,N_14815);
nand U15096 (N_15096,N_14451,N_14828);
nor U15097 (N_15097,N_14458,N_14836);
nor U15098 (N_15098,N_14566,N_14937);
xor U15099 (N_15099,N_14812,N_14882);
nor U15100 (N_15100,N_14904,N_14440);
nand U15101 (N_15101,N_14935,N_14785);
or U15102 (N_15102,N_14797,N_14586);
and U15103 (N_15103,N_14788,N_14401);
xnor U15104 (N_15104,N_14883,N_14846);
and U15105 (N_15105,N_14516,N_14519);
nand U15106 (N_15106,N_14542,N_14581);
xor U15107 (N_15107,N_14778,N_14644);
nor U15108 (N_15108,N_14870,N_14709);
xor U15109 (N_15109,N_14796,N_14921);
and U15110 (N_15110,N_14503,N_14985);
xnor U15111 (N_15111,N_14438,N_14527);
and U15112 (N_15112,N_14995,N_14902);
xnor U15113 (N_15113,N_14789,N_14421);
and U15114 (N_15114,N_14889,N_14775);
xor U15115 (N_15115,N_14833,N_14652);
or U15116 (N_15116,N_14588,N_14864);
nor U15117 (N_15117,N_14617,N_14926);
xor U15118 (N_15118,N_14749,N_14618);
and U15119 (N_15119,N_14678,N_14667);
or U15120 (N_15120,N_14824,N_14536);
or U15121 (N_15121,N_14634,N_14671);
nor U15122 (N_15122,N_14769,N_14765);
or U15123 (N_15123,N_14590,N_14933);
or U15124 (N_15124,N_14463,N_14793);
xor U15125 (N_15125,N_14609,N_14866);
or U15126 (N_15126,N_14592,N_14747);
xnor U15127 (N_15127,N_14855,N_14544);
or U15128 (N_15128,N_14914,N_14912);
or U15129 (N_15129,N_14541,N_14695);
and U15130 (N_15130,N_14640,N_14906);
nor U15131 (N_15131,N_14485,N_14533);
and U15132 (N_15132,N_14737,N_14895);
and U15133 (N_15133,N_14467,N_14875);
nand U15134 (N_15134,N_14480,N_14564);
xor U15135 (N_15135,N_14715,N_14910);
and U15136 (N_15136,N_14598,N_14472);
nor U15137 (N_15137,N_14474,N_14673);
xnor U15138 (N_15138,N_14837,N_14746);
or U15139 (N_15139,N_14649,N_14919);
nor U15140 (N_15140,N_14884,N_14940);
nand U15141 (N_15141,N_14669,N_14780);
nand U15142 (N_15142,N_14557,N_14420);
xnor U15143 (N_15143,N_14943,N_14745);
nor U15144 (N_15144,N_14538,N_14665);
nor U15145 (N_15145,N_14642,N_14431);
nand U15146 (N_15146,N_14991,N_14858);
or U15147 (N_15147,N_14876,N_14980);
and U15148 (N_15148,N_14510,N_14774);
and U15149 (N_15149,N_14660,N_14585);
nand U15150 (N_15150,N_14653,N_14613);
xnor U15151 (N_15151,N_14400,N_14512);
nand U15152 (N_15152,N_14905,N_14502);
or U15153 (N_15153,N_14682,N_14958);
and U15154 (N_15154,N_14484,N_14852);
or U15155 (N_15155,N_14738,N_14637);
nand U15156 (N_15156,N_14945,N_14627);
or U15157 (N_15157,N_14486,N_14622);
nor U15158 (N_15158,N_14413,N_14990);
and U15159 (N_15159,N_14929,N_14763);
or U15160 (N_15160,N_14657,N_14953);
and U15161 (N_15161,N_14487,N_14539);
nand U15162 (N_15162,N_14661,N_14520);
or U15163 (N_15163,N_14786,N_14839);
nand U15164 (N_15164,N_14621,N_14444);
or U15165 (N_15165,N_14602,N_14844);
or U15166 (N_15166,N_14422,N_14583);
nor U15167 (N_15167,N_14623,N_14805);
nand U15168 (N_15168,N_14680,N_14576);
and U15169 (N_15169,N_14603,N_14930);
or U15170 (N_15170,N_14903,N_14435);
or U15171 (N_15171,N_14795,N_14689);
or U15172 (N_15172,N_14758,N_14404);
xor U15173 (N_15173,N_14831,N_14662);
and U15174 (N_15174,N_14643,N_14992);
xor U15175 (N_15175,N_14975,N_14675);
nor U15176 (N_15176,N_14807,N_14429);
nand U15177 (N_15177,N_14498,N_14482);
xnor U15178 (N_15178,N_14885,N_14407);
nor U15179 (N_15179,N_14859,N_14526);
xor U15180 (N_15180,N_14947,N_14556);
or U15181 (N_15181,N_14868,N_14461);
xor U15182 (N_15182,N_14867,N_14567);
nor U15183 (N_15183,N_14412,N_14651);
nand U15184 (N_15184,N_14750,N_14957);
nand U15185 (N_15185,N_14711,N_14941);
xnor U15186 (N_15186,N_14515,N_14656);
or U15187 (N_15187,N_14949,N_14572);
nor U15188 (N_15188,N_14773,N_14625);
or U15189 (N_15189,N_14748,N_14909);
xor U15190 (N_15190,N_14965,N_14641);
and U15191 (N_15191,N_14477,N_14614);
nand U15192 (N_15192,N_14418,N_14672);
xor U15193 (N_15193,N_14650,N_14728);
and U15194 (N_15194,N_14959,N_14865);
nand U15195 (N_15195,N_14521,N_14437);
or U15196 (N_15196,N_14800,N_14722);
xor U15197 (N_15197,N_14690,N_14594);
or U15198 (N_15198,N_14893,N_14900);
nor U15199 (N_15199,N_14468,N_14894);
and U15200 (N_15200,N_14615,N_14829);
and U15201 (N_15201,N_14419,N_14551);
or U15202 (N_15202,N_14546,N_14605);
nor U15203 (N_15203,N_14559,N_14645);
and U15204 (N_15204,N_14449,N_14500);
xor U15205 (N_15205,N_14874,N_14692);
nand U15206 (N_15206,N_14821,N_14626);
or U15207 (N_15207,N_14794,N_14787);
xor U15208 (N_15208,N_14798,N_14528);
xnor U15209 (N_15209,N_14822,N_14506);
nand U15210 (N_15210,N_14716,N_14951);
or U15211 (N_15211,N_14917,N_14441);
xor U15212 (N_15212,N_14850,N_14986);
xor U15213 (N_15213,N_14948,N_14599);
and U15214 (N_15214,N_14936,N_14417);
and U15215 (N_15215,N_14664,N_14720);
nand U15216 (N_15216,N_14606,N_14962);
or U15217 (N_15217,N_14433,N_14654);
nand U15218 (N_15218,N_14648,N_14899);
nor U15219 (N_15219,N_14781,N_14963);
and U15220 (N_15220,N_14469,N_14674);
nor U15221 (N_15221,N_14702,N_14473);
nor U15222 (N_15222,N_14840,N_14803);
nand U15223 (N_15223,N_14439,N_14697);
nand U15224 (N_15224,N_14759,N_14727);
nor U15225 (N_15225,N_14423,N_14892);
nand U15226 (N_15226,N_14532,N_14492);
nor U15227 (N_15227,N_14628,N_14934);
or U15228 (N_15228,N_14666,N_14710);
nand U15229 (N_15229,N_14658,N_14501);
nand U15230 (N_15230,N_14997,N_14952);
and U15231 (N_15231,N_14631,N_14872);
nand U15232 (N_15232,N_14405,N_14459);
nand U15233 (N_15233,N_14955,N_14869);
xnor U15234 (N_15234,N_14888,N_14548);
or U15235 (N_15235,N_14907,N_14954);
and U15236 (N_15236,N_14577,N_14547);
and U15237 (N_15237,N_14550,N_14925);
xnor U15238 (N_15238,N_14570,N_14854);
nor U15239 (N_15239,N_14424,N_14687);
or U15240 (N_15240,N_14740,N_14724);
xnor U15241 (N_15241,N_14915,N_14663);
xnor U15242 (N_15242,N_14860,N_14408);
xnor U15243 (N_15243,N_14497,N_14984);
or U15244 (N_15244,N_14573,N_14568);
nand U15245 (N_15245,N_14726,N_14523);
and U15246 (N_15246,N_14402,N_14630);
nor U15247 (N_15247,N_14928,N_14960);
xor U15248 (N_15248,N_14549,N_14681);
xor U15249 (N_15249,N_14911,N_14942);
nor U15250 (N_15250,N_14508,N_14820);
or U15251 (N_15251,N_14856,N_14974);
nand U15252 (N_15252,N_14754,N_14475);
xnor U15253 (N_15253,N_14725,N_14923);
and U15254 (N_15254,N_14704,N_14755);
nand U15255 (N_15255,N_14545,N_14700);
xor U15256 (N_15256,N_14735,N_14760);
nor U15257 (N_15257,N_14677,N_14632);
nand U15258 (N_15258,N_14616,N_14751);
nor U15259 (N_15259,N_14558,N_14920);
nand U15260 (N_15260,N_14436,N_14507);
and U15261 (N_15261,N_14593,N_14668);
or U15262 (N_15262,N_14956,N_14723);
and U15263 (N_15263,N_14968,N_14597);
and U15264 (N_15264,N_14971,N_14403);
nand U15265 (N_15265,N_14999,N_14790);
xnor U15266 (N_15266,N_14596,N_14530);
nand U15267 (N_15267,N_14802,N_14679);
nand U15268 (N_15268,N_14415,N_14825);
xnor U15269 (N_15269,N_14757,N_14608);
xnor U15270 (N_15270,N_14525,N_14851);
xor U15271 (N_15271,N_14932,N_14575);
nand U15272 (N_15272,N_14732,N_14426);
and U15273 (N_15273,N_14580,N_14808);
or U15274 (N_15274,N_14504,N_14927);
and U15275 (N_15275,N_14770,N_14489);
and U15276 (N_15276,N_14445,N_14879);
xor U15277 (N_15277,N_14714,N_14465);
xor U15278 (N_15278,N_14998,N_14901);
xor U15279 (N_15279,N_14693,N_14813);
or U15280 (N_15280,N_14481,N_14988);
nor U15281 (N_15281,N_14427,N_14964);
and U15282 (N_15282,N_14494,N_14553);
and U15283 (N_15283,N_14877,N_14743);
or U15284 (N_15284,N_14646,N_14707);
xnor U15285 (N_15285,N_14981,N_14816);
xnor U15286 (N_15286,N_14896,N_14944);
nor U15287 (N_15287,N_14845,N_14601);
and U15288 (N_15288,N_14827,N_14898);
or U15289 (N_15289,N_14806,N_14961);
or U15290 (N_15290,N_14416,N_14862);
and U15291 (N_15291,N_14916,N_14531);
xnor U15292 (N_15292,N_14683,N_14589);
nor U15293 (N_15293,N_14776,N_14857);
or U15294 (N_15294,N_14970,N_14718);
nand U15295 (N_15295,N_14425,N_14409);
xor U15296 (N_15296,N_14717,N_14638);
and U15297 (N_15297,N_14701,N_14848);
and U15298 (N_15298,N_14490,N_14624);
xnor U15299 (N_15299,N_14818,N_14561);
nand U15300 (N_15300,N_14624,N_14948);
and U15301 (N_15301,N_14715,N_14757);
and U15302 (N_15302,N_14490,N_14698);
and U15303 (N_15303,N_14607,N_14832);
nor U15304 (N_15304,N_14709,N_14778);
or U15305 (N_15305,N_14803,N_14491);
xor U15306 (N_15306,N_14552,N_14678);
or U15307 (N_15307,N_14763,N_14962);
and U15308 (N_15308,N_14479,N_14719);
nand U15309 (N_15309,N_14641,N_14418);
xor U15310 (N_15310,N_14434,N_14472);
and U15311 (N_15311,N_14706,N_14866);
nand U15312 (N_15312,N_14421,N_14932);
xor U15313 (N_15313,N_14823,N_14734);
or U15314 (N_15314,N_14763,N_14524);
nor U15315 (N_15315,N_14538,N_14828);
xor U15316 (N_15316,N_14956,N_14840);
nor U15317 (N_15317,N_14430,N_14774);
xnor U15318 (N_15318,N_14961,N_14905);
and U15319 (N_15319,N_14470,N_14960);
nand U15320 (N_15320,N_14998,N_14557);
or U15321 (N_15321,N_14462,N_14566);
and U15322 (N_15322,N_14778,N_14607);
xnor U15323 (N_15323,N_14668,N_14876);
and U15324 (N_15324,N_14871,N_14798);
or U15325 (N_15325,N_14665,N_14724);
and U15326 (N_15326,N_14841,N_14678);
and U15327 (N_15327,N_14961,N_14833);
xnor U15328 (N_15328,N_14874,N_14477);
nor U15329 (N_15329,N_14689,N_14583);
xor U15330 (N_15330,N_14969,N_14538);
or U15331 (N_15331,N_14968,N_14499);
or U15332 (N_15332,N_14763,N_14472);
nand U15333 (N_15333,N_14467,N_14922);
and U15334 (N_15334,N_14599,N_14718);
or U15335 (N_15335,N_14759,N_14472);
nor U15336 (N_15336,N_14738,N_14785);
xor U15337 (N_15337,N_14533,N_14966);
nor U15338 (N_15338,N_14453,N_14893);
nand U15339 (N_15339,N_14699,N_14572);
xor U15340 (N_15340,N_14918,N_14881);
nand U15341 (N_15341,N_14684,N_14964);
nor U15342 (N_15342,N_14823,N_14660);
and U15343 (N_15343,N_14674,N_14412);
or U15344 (N_15344,N_14970,N_14431);
nand U15345 (N_15345,N_14606,N_14991);
nor U15346 (N_15346,N_14645,N_14983);
nand U15347 (N_15347,N_14512,N_14760);
nand U15348 (N_15348,N_14422,N_14747);
xor U15349 (N_15349,N_14872,N_14575);
nand U15350 (N_15350,N_14424,N_14497);
nand U15351 (N_15351,N_14525,N_14575);
nand U15352 (N_15352,N_14921,N_14479);
nand U15353 (N_15353,N_14711,N_14890);
nor U15354 (N_15354,N_14470,N_14846);
nand U15355 (N_15355,N_14458,N_14445);
and U15356 (N_15356,N_14828,N_14702);
nor U15357 (N_15357,N_14621,N_14698);
and U15358 (N_15358,N_14906,N_14403);
and U15359 (N_15359,N_14527,N_14956);
and U15360 (N_15360,N_14681,N_14741);
or U15361 (N_15361,N_14843,N_14721);
and U15362 (N_15362,N_14917,N_14944);
and U15363 (N_15363,N_14900,N_14890);
nor U15364 (N_15364,N_14930,N_14983);
nand U15365 (N_15365,N_14792,N_14668);
or U15366 (N_15366,N_14596,N_14721);
xor U15367 (N_15367,N_14934,N_14439);
or U15368 (N_15368,N_14734,N_14856);
xor U15369 (N_15369,N_14487,N_14881);
or U15370 (N_15370,N_14540,N_14502);
nor U15371 (N_15371,N_14882,N_14605);
or U15372 (N_15372,N_14762,N_14448);
nor U15373 (N_15373,N_14814,N_14701);
nor U15374 (N_15374,N_14796,N_14557);
or U15375 (N_15375,N_14626,N_14754);
and U15376 (N_15376,N_14856,N_14461);
or U15377 (N_15377,N_14795,N_14443);
nand U15378 (N_15378,N_14929,N_14768);
and U15379 (N_15379,N_14547,N_14694);
xnor U15380 (N_15380,N_14993,N_14466);
nand U15381 (N_15381,N_14891,N_14951);
or U15382 (N_15382,N_14645,N_14718);
xor U15383 (N_15383,N_14975,N_14874);
and U15384 (N_15384,N_14448,N_14621);
nor U15385 (N_15385,N_14848,N_14501);
and U15386 (N_15386,N_14615,N_14708);
or U15387 (N_15387,N_14426,N_14904);
or U15388 (N_15388,N_14628,N_14503);
and U15389 (N_15389,N_14904,N_14987);
or U15390 (N_15390,N_14577,N_14523);
or U15391 (N_15391,N_14612,N_14478);
nand U15392 (N_15392,N_14452,N_14746);
and U15393 (N_15393,N_14797,N_14510);
nand U15394 (N_15394,N_14457,N_14992);
and U15395 (N_15395,N_14805,N_14658);
nor U15396 (N_15396,N_14968,N_14625);
xnor U15397 (N_15397,N_14496,N_14403);
and U15398 (N_15398,N_14535,N_14520);
or U15399 (N_15399,N_14462,N_14969);
or U15400 (N_15400,N_14423,N_14889);
and U15401 (N_15401,N_14760,N_14753);
nand U15402 (N_15402,N_14444,N_14995);
or U15403 (N_15403,N_14542,N_14472);
nor U15404 (N_15404,N_14772,N_14642);
nor U15405 (N_15405,N_14464,N_14675);
and U15406 (N_15406,N_14883,N_14973);
nor U15407 (N_15407,N_14888,N_14802);
and U15408 (N_15408,N_14611,N_14914);
xnor U15409 (N_15409,N_14468,N_14434);
and U15410 (N_15410,N_14524,N_14482);
nand U15411 (N_15411,N_14778,N_14550);
and U15412 (N_15412,N_14456,N_14711);
nand U15413 (N_15413,N_14633,N_14497);
and U15414 (N_15414,N_14726,N_14779);
or U15415 (N_15415,N_14508,N_14430);
xor U15416 (N_15416,N_14643,N_14712);
and U15417 (N_15417,N_14754,N_14997);
nor U15418 (N_15418,N_14886,N_14894);
nand U15419 (N_15419,N_14728,N_14988);
nor U15420 (N_15420,N_14844,N_14707);
nor U15421 (N_15421,N_14427,N_14993);
or U15422 (N_15422,N_14818,N_14801);
and U15423 (N_15423,N_14652,N_14421);
and U15424 (N_15424,N_14964,N_14768);
xor U15425 (N_15425,N_14725,N_14689);
or U15426 (N_15426,N_14967,N_14946);
or U15427 (N_15427,N_14870,N_14672);
or U15428 (N_15428,N_14659,N_14475);
xnor U15429 (N_15429,N_14990,N_14479);
xor U15430 (N_15430,N_14625,N_14742);
or U15431 (N_15431,N_14922,N_14631);
nor U15432 (N_15432,N_14805,N_14870);
nor U15433 (N_15433,N_14672,N_14914);
nand U15434 (N_15434,N_14432,N_14836);
nand U15435 (N_15435,N_14825,N_14792);
and U15436 (N_15436,N_14476,N_14526);
and U15437 (N_15437,N_14523,N_14674);
nor U15438 (N_15438,N_14799,N_14435);
nand U15439 (N_15439,N_14488,N_14777);
nand U15440 (N_15440,N_14526,N_14563);
xnor U15441 (N_15441,N_14575,N_14798);
or U15442 (N_15442,N_14832,N_14768);
or U15443 (N_15443,N_14812,N_14500);
nand U15444 (N_15444,N_14687,N_14678);
nand U15445 (N_15445,N_14607,N_14732);
or U15446 (N_15446,N_14760,N_14994);
nor U15447 (N_15447,N_14537,N_14626);
nor U15448 (N_15448,N_14740,N_14776);
nand U15449 (N_15449,N_14543,N_14695);
and U15450 (N_15450,N_14679,N_14936);
nor U15451 (N_15451,N_14720,N_14544);
nor U15452 (N_15452,N_14748,N_14792);
or U15453 (N_15453,N_14460,N_14685);
xnor U15454 (N_15454,N_14656,N_14572);
nor U15455 (N_15455,N_14974,N_14988);
and U15456 (N_15456,N_14870,N_14731);
or U15457 (N_15457,N_14775,N_14621);
or U15458 (N_15458,N_14929,N_14471);
and U15459 (N_15459,N_14483,N_14844);
or U15460 (N_15460,N_14888,N_14755);
nor U15461 (N_15461,N_14883,N_14700);
or U15462 (N_15462,N_14693,N_14417);
xnor U15463 (N_15463,N_14407,N_14990);
nand U15464 (N_15464,N_14787,N_14473);
or U15465 (N_15465,N_14671,N_14568);
xor U15466 (N_15466,N_14679,N_14601);
nand U15467 (N_15467,N_14840,N_14489);
nor U15468 (N_15468,N_14638,N_14673);
nor U15469 (N_15469,N_14648,N_14974);
and U15470 (N_15470,N_14872,N_14929);
or U15471 (N_15471,N_14945,N_14733);
and U15472 (N_15472,N_14788,N_14825);
xor U15473 (N_15473,N_14632,N_14684);
xnor U15474 (N_15474,N_14778,N_14537);
nand U15475 (N_15475,N_14937,N_14542);
or U15476 (N_15476,N_14833,N_14700);
nor U15477 (N_15477,N_14814,N_14569);
and U15478 (N_15478,N_14634,N_14676);
nand U15479 (N_15479,N_14540,N_14523);
xor U15480 (N_15480,N_14898,N_14772);
xnor U15481 (N_15481,N_14783,N_14917);
xor U15482 (N_15482,N_14988,N_14530);
xor U15483 (N_15483,N_14649,N_14964);
and U15484 (N_15484,N_14433,N_14945);
or U15485 (N_15485,N_14819,N_14565);
xnor U15486 (N_15486,N_14532,N_14967);
nand U15487 (N_15487,N_14970,N_14590);
nand U15488 (N_15488,N_14848,N_14686);
nor U15489 (N_15489,N_14743,N_14709);
nand U15490 (N_15490,N_14895,N_14468);
xor U15491 (N_15491,N_14955,N_14490);
xnor U15492 (N_15492,N_14549,N_14690);
or U15493 (N_15493,N_14966,N_14985);
xor U15494 (N_15494,N_14750,N_14578);
nor U15495 (N_15495,N_14580,N_14889);
nand U15496 (N_15496,N_14457,N_14926);
nor U15497 (N_15497,N_14612,N_14828);
xnor U15498 (N_15498,N_14850,N_14421);
nand U15499 (N_15499,N_14981,N_14910);
or U15500 (N_15500,N_14545,N_14452);
xor U15501 (N_15501,N_14820,N_14533);
nor U15502 (N_15502,N_14913,N_14495);
nor U15503 (N_15503,N_14983,N_14512);
nor U15504 (N_15504,N_14915,N_14504);
xor U15505 (N_15505,N_14708,N_14882);
nor U15506 (N_15506,N_14938,N_14444);
nor U15507 (N_15507,N_14537,N_14672);
nor U15508 (N_15508,N_14545,N_14816);
or U15509 (N_15509,N_14949,N_14709);
or U15510 (N_15510,N_14739,N_14447);
and U15511 (N_15511,N_14438,N_14906);
and U15512 (N_15512,N_14467,N_14720);
or U15513 (N_15513,N_14942,N_14640);
or U15514 (N_15514,N_14907,N_14670);
nor U15515 (N_15515,N_14791,N_14777);
nor U15516 (N_15516,N_14481,N_14490);
or U15517 (N_15517,N_14702,N_14573);
xor U15518 (N_15518,N_14592,N_14892);
and U15519 (N_15519,N_14981,N_14437);
nand U15520 (N_15520,N_14738,N_14528);
nand U15521 (N_15521,N_14581,N_14932);
nand U15522 (N_15522,N_14599,N_14779);
and U15523 (N_15523,N_14705,N_14524);
and U15524 (N_15524,N_14659,N_14632);
xor U15525 (N_15525,N_14966,N_14521);
nor U15526 (N_15526,N_14745,N_14655);
xor U15527 (N_15527,N_14819,N_14763);
and U15528 (N_15528,N_14501,N_14811);
nor U15529 (N_15529,N_14973,N_14949);
and U15530 (N_15530,N_14413,N_14938);
and U15531 (N_15531,N_14819,N_14443);
nand U15532 (N_15532,N_14970,N_14568);
and U15533 (N_15533,N_14853,N_14601);
or U15534 (N_15534,N_14992,N_14506);
nor U15535 (N_15535,N_14605,N_14661);
and U15536 (N_15536,N_14523,N_14552);
or U15537 (N_15537,N_14620,N_14482);
xor U15538 (N_15538,N_14602,N_14705);
and U15539 (N_15539,N_14806,N_14488);
xor U15540 (N_15540,N_14846,N_14830);
nand U15541 (N_15541,N_14528,N_14672);
nand U15542 (N_15542,N_14845,N_14429);
nor U15543 (N_15543,N_14935,N_14700);
nand U15544 (N_15544,N_14611,N_14478);
nor U15545 (N_15545,N_14468,N_14764);
or U15546 (N_15546,N_14909,N_14760);
and U15547 (N_15547,N_14509,N_14686);
and U15548 (N_15548,N_14729,N_14512);
xnor U15549 (N_15549,N_14631,N_14514);
and U15550 (N_15550,N_14426,N_14572);
nor U15551 (N_15551,N_14745,N_14616);
or U15552 (N_15552,N_14588,N_14555);
xor U15553 (N_15553,N_14494,N_14617);
nor U15554 (N_15554,N_14882,N_14995);
or U15555 (N_15555,N_14588,N_14529);
or U15556 (N_15556,N_14600,N_14965);
xnor U15557 (N_15557,N_14612,N_14599);
nand U15558 (N_15558,N_14499,N_14638);
nand U15559 (N_15559,N_14974,N_14800);
or U15560 (N_15560,N_14498,N_14560);
nand U15561 (N_15561,N_14840,N_14859);
nand U15562 (N_15562,N_14881,N_14631);
nand U15563 (N_15563,N_14814,N_14919);
and U15564 (N_15564,N_14802,N_14819);
xnor U15565 (N_15565,N_14441,N_14515);
nor U15566 (N_15566,N_14625,N_14591);
and U15567 (N_15567,N_14468,N_14491);
and U15568 (N_15568,N_14944,N_14438);
or U15569 (N_15569,N_14731,N_14773);
xnor U15570 (N_15570,N_14959,N_14700);
nand U15571 (N_15571,N_14812,N_14658);
xor U15572 (N_15572,N_14705,N_14980);
and U15573 (N_15573,N_14651,N_14951);
nand U15574 (N_15574,N_14852,N_14415);
or U15575 (N_15575,N_14948,N_14480);
nor U15576 (N_15576,N_14616,N_14639);
xor U15577 (N_15577,N_14904,N_14744);
nand U15578 (N_15578,N_14403,N_14818);
or U15579 (N_15579,N_14494,N_14972);
xnor U15580 (N_15580,N_14600,N_14610);
and U15581 (N_15581,N_14934,N_14904);
nand U15582 (N_15582,N_14671,N_14674);
and U15583 (N_15583,N_14610,N_14704);
and U15584 (N_15584,N_14911,N_14941);
and U15585 (N_15585,N_14628,N_14554);
nand U15586 (N_15586,N_14428,N_14733);
nand U15587 (N_15587,N_14715,N_14481);
or U15588 (N_15588,N_14572,N_14586);
nand U15589 (N_15589,N_14625,N_14503);
nor U15590 (N_15590,N_14820,N_14878);
nand U15591 (N_15591,N_14822,N_14411);
nand U15592 (N_15592,N_14736,N_14925);
nand U15593 (N_15593,N_14698,N_14889);
xnor U15594 (N_15594,N_14965,N_14728);
nor U15595 (N_15595,N_14740,N_14581);
nand U15596 (N_15596,N_14915,N_14804);
and U15597 (N_15597,N_14439,N_14819);
xnor U15598 (N_15598,N_14762,N_14515);
or U15599 (N_15599,N_14619,N_14425);
xor U15600 (N_15600,N_15498,N_15387);
nand U15601 (N_15601,N_15118,N_15300);
xor U15602 (N_15602,N_15510,N_15474);
and U15603 (N_15603,N_15129,N_15362);
and U15604 (N_15604,N_15508,N_15313);
xor U15605 (N_15605,N_15316,N_15009);
or U15606 (N_15606,N_15022,N_15163);
nor U15607 (N_15607,N_15132,N_15098);
and U15608 (N_15608,N_15452,N_15228);
xnor U15609 (N_15609,N_15599,N_15516);
and U15610 (N_15610,N_15336,N_15564);
nand U15611 (N_15611,N_15295,N_15419);
nand U15612 (N_15612,N_15406,N_15094);
or U15613 (N_15613,N_15400,N_15032);
xnor U15614 (N_15614,N_15147,N_15287);
xnor U15615 (N_15615,N_15507,N_15397);
or U15616 (N_15616,N_15591,N_15082);
and U15617 (N_15617,N_15131,N_15284);
xnor U15618 (N_15618,N_15345,N_15558);
nor U15619 (N_15619,N_15398,N_15008);
and U15620 (N_15620,N_15236,N_15057);
nand U15621 (N_15621,N_15401,N_15451);
and U15622 (N_15622,N_15299,N_15254);
nor U15623 (N_15623,N_15159,N_15160);
nor U15624 (N_15624,N_15069,N_15093);
and U15625 (N_15625,N_15352,N_15246);
nor U15626 (N_15626,N_15531,N_15086);
xnor U15627 (N_15627,N_15480,N_15124);
nor U15628 (N_15628,N_15281,N_15413);
xnor U15629 (N_15629,N_15154,N_15115);
and U15630 (N_15630,N_15338,N_15371);
xor U15631 (N_15631,N_15309,N_15101);
or U15632 (N_15632,N_15056,N_15139);
xor U15633 (N_15633,N_15261,N_15590);
or U15634 (N_15634,N_15404,N_15497);
nand U15635 (N_15635,N_15321,N_15063);
and U15636 (N_15636,N_15412,N_15355);
and U15637 (N_15637,N_15211,N_15275);
or U15638 (N_15638,N_15052,N_15422);
xnor U15639 (N_15639,N_15088,N_15007);
nor U15640 (N_15640,N_15542,N_15396);
nand U15641 (N_15641,N_15249,N_15023);
and U15642 (N_15642,N_15453,N_15036);
nand U15643 (N_15643,N_15066,N_15125);
xnor U15644 (N_15644,N_15526,N_15193);
xor U15645 (N_15645,N_15500,N_15424);
nand U15646 (N_15646,N_15169,N_15204);
or U15647 (N_15647,N_15148,N_15006);
and U15648 (N_15648,N_15043,N_15378);
xor U15649 (N_15649,N_15178,N_15533);
nand U15650 (N_15650,N_15539,N_15015);
or U15651 (N_15651,N_15303,N_15501);
and U15652 (N_15652,N_15385,N_15201);
xnor U15653 (N_15653,N_15464,N_15174);
and U15654 (N_15654,N_15248,N_15183);
xor U15655 (N_15655,N_15024,N_15527);
or U15656 (N_15656,N_15065,N_15070);
or U15657 (N_15657,N_15179,N_15324);
and U15658 (N_15658,N_15367,N_15524);
and U15659 (N_15659,N_15012,N_15307);
nand U15660 (N_15660,N_15436,N_15105);
and U15661 (N_15661,N_15523,N_15005);
and U15662 (N_15662,N_15283,N_15374);
or U15663 (N_15663,N_15215,N_15540);
nor U15664 (N_15664,N_15266,N_15472);
or U15665 (N_15665,N_15432,N_15317);
or U15666 (N_15666,N_15091,N_15175);
nor U15667 (N_15667,N_15102,N_15077);
nand U15668 (N_15668,N_15586,N_15117);
xnor U15669 (N_15669,N_15176,N_15550);
nor U15670 (N_15670,N_15003,N_15414);
xor U15671 (N_15671,N_15133,N_15529);
xnor U15672 (N_15672,N_15241,N_15545);
nor U15673 (N_15673,N_15409,N_15209);
nand U15674 (N_15674,N_15037,N_15226);
nor U15675 (N_15675,N_15136,N_15020);
and U15676 (N_15676,N_15290,N_15503);
or U15677 (N_15677,N_15013,N_15106);
nor U15678 (N_15678,N_15061,N_15110);
and U15679 (N_15679,N_15348,N_15244);
nor U15680 (N_15680,N_15194,N_15479);
xor U15681 (N_15681,N_15572,N_15068);
and U15682 (N_15682,N_15173,N_15585);
nand U15683 (N_15683,N_15205,N_15121);
or U15684 (N_15684,N_15084,N_15016);
xor U15685 (N_15685,N_15319,N_15189);
nand U15686 (N_15686,N_15227,N_15269);
and U15687 (N_15687,N_15067,N_15502);
nor U15688 (N_15688,N_15337,N_15315);
and U15689 (N_15689,N_15033,N_15489);
nor U15690 (N_15690,N_15377,N_15430);
and U15691 (N_15691,N_15292,N_15334);
and U15692 (N_15692,N_15140,N_15191);
xor U15693 (N_15693,N_15206,N_15221);
and U15694 (N_15694,N_15238,N_15468);
nand U15695 (N_15695,N_15030,N_15286);
and U15696 (N_15696,N_15028,N_15113);
nor U15697 (N_15697,N_15518,N_15144);
nand U15698 (N_15698,N_15382,N_15096);
nand U15699 (N_15699,N_15198,N_15354);
and U15700 (N_15700,N_15492,N_15108);
nor U15701 (N_15701,N_15232,N_15368);
and U15702 (N_15702,N_15049,N_15351);
xnor U15703 (N_15703,N_15537,N_15549);
nor U15704 (N_15704,N_15567,N_15062);
nand U15705 (N_15705,N_15493,N_15104);
or U15706 (N_15706,N_15127,N_15343);
nand U15707 (N_15707,N_15310,N_15053);
or U15708 (N_15708,N_15212,N_15167);
and U15709 (N_15709,N_15214,N_15166);
nor U15710 (N_15710,N_15255,N_15584);
and U15711 (N_15711,N_15520,N_15554);
nor U15712 (N_15712,N_15234,N_15328);
nor U15713 (N_15713,N_15297,N_15044);
nor U15714 (N_15714,N_15568,N_15505);
xor U15715 (N_15715,N_15274,N_15389);
nand U15716 (N_15716,N_15509,N_15454);
and U15717 (N_15717,N_15188,N_15482);
or U15718 (N_15718,N_15279,N_15237);
nand U15719 (N_15719,N_15552,N_15207);
xor U15720 (N_15720,N_15320,N_15141);
or U15721 (N_15721,N_15029,N_15405);
and U15722 (N_15722,N_15597,N_15090);
or U15723 (N_15723,N_15285,N_15153);
or U15724 (N_15724,N_15532,N_15589);
and U15725 (N_15725,N_15277,N_15548);
or U15726 (N_15726,N_15031,N_15461);
nand U15727 (N_15727,N_15122,N_15119);
nand U15728 (N_15728,N_15087,N_15027);
nand U15729 (N_15729,N_15200,N_15380);
or U15730 (N_15730,N_15384,N_15410);
and U15731 (N_15731,N_15511,N_15571);
or U15732 (N_15732,N_15039,N_15562);
or U15733 (N_15733,N_15262,N_15535);
nand U15734 (N_15734,N_15434,N_15199);
nand U15735 (N_15735,N_15242,N_15187);
nand U15736 (N_15736,N_15534,N_15443);
xor U15737 (N_15737,N_15391,N_15379);
nor U15738 (N_15738,N_15038,N_15225);
nand U15739 (N_15739,N_15126,N_15460);
nor U15740 (N_15740,N_15557,N_15314);
or U15741 (N_15741,N_15517,N_15408);
and U15742 (N_15742,N_15473,N_15288);
xor U15743 (N_15743,N_15339,N_15559);
nor U15744 (N_15744,N_15109,N_15081);
nand U15745 (N_15745,N_15356,N_15340);
nor U15746 (N_15746,N_15580,N_15402);
or U15747 (N_15747,N_15040,N_15487);
nand U15748 (N_15748,N_15470,N_15363);
or U15749 (N_15749,N_15513,N_15318);
and U15750 (N_15750,N_15395,N_15325);
nor U15751 (N_15751,N_15270,N_15469);
and U15752 (N_15752,N_15440,N_15197);
xnor U15753 (N_15753,N_15230,N_15560);
and U15754 (N_15754,N_15569,N_15346);
nand U15755 (N_15755,N_15563,N_15311);
xor U15756 (N_15756,N_15393,N_15344);
nor U15757 (N_15757,N_15594,N_15465);
and U15758 (N_15758,N_15525,N_15095);
nand U15759 (N_15759,N_15018,N_15157);
and U15760 (N_15760,N_15298,N_15547);
xor U15761 (N_15761,N_15014,N_15078);
or U15762 (N_15762,N_15546,N_15411);
and U15763 (N_15763,N_15556,N_15239);
nand U15764 (N_15764,N_15579,N_15151);
or U15765 (N_15765,N_15566,N_15235);
and U15766 (N_15766,N_15483,N_15152);
nor U15767 (N_15767,N_15282,N_15172);
or U15768 (N_15768,N_15381,N_15467);
nand U15769 (N_15769,N_15047,N_15000);
nor U15770 (N_15770,N_15251,N_15418);
nand U15771 (N_15771,N_15494,N_15192);
and U15772 (N_15772,N_15437,N_15276);
xnor U15773 (N_15773,N_15046,N_15386);
nor U15774 (N_15774,N_15449,N_15264);
nand U15775 (N_15775,N_15265,N_15146);
or U15776 (N_15776,N_15514,N_15375);
and U15777 (N_15777,N_15025,N_15369);
xnor U15778 (N_15778,N_15100,N_15185);
xor U15779 (N_15779,N_15322,N_15574);
nand U15780 (N_15780,N_15538,N_15019);
and U15781 (N_15781,N_15582,N_15370);
nand U15782 (N_15782,N_15011,N_15528);
xnor U15783 (N_15783,N_15457,N_15233);
xor U15784 (N_15784,N_15010,N_15448);
xor U15785 (N_15785,N_15312,N_15123);
nor U15786 (N_15786,N_15263,N_15486);
nand U15787 (N_15787,N_15138,N_15331);
or U15788 (N_15788,N_15426,N_15485);
xnor U15789 (N_15789,N_15156,N_15196);
or U15790 (N_15790,N_15522,N_15074);
nand U15791 (N_15791,N_15596,N_15143);
nor U15792 (N_15792,N_15137,N_15353);
and U15793 (N_15793,N_15427,N_15471);
and U15794 (N_15794,N_15506,N_15423);
nor U15795 (N_15795,N_15092,N_15112);
and U15796 (N_15796,N_15210,N_15161);
or U15797 (N_15797,N_15330,N_15250);
nand U15798 (N_15798,N_15289,N_15271);
nand U15799 (N_15799,N_15541,N_15583);
nand U15800 (N_15800,N_15488,N_15403);
nand U15801 (N_15801,N_15213,N_15515);
or U15802 (N_15802,N_15359,N_15064);
xnor U15803 (N_15803,N_15577,N_15203);
xnor U15804 (N_15804,N_15543,N_15245);
xnor U15805 (N_15805,N_15588,N_15216);
or U15806 (N_15806,N_15327,N_15180);
and U15807 (N_15807,N_15111,N_15184);
or U15808 (N_15808,N_15442,N_15456);
and U15809 (N_15809,N_15155,N_15496);
xor U15810 (N_15810,N_15335,N_15222);
or U15811 (N_15811,N_15190,N_15182);
nor U15812 (N_15812,N_15120,N_15519);
and U15813 (N_15813,N_15438,N_15373);
nor U15814 (N_15814,N_15165,N_15475);
nand U15815 (N_15815,N_15202,N_15060);
nand U15816 (N_15816,N_15392,N_15581);
or U15817 (N_15817,N_15116,N_15079);
xor U15818 (N_15818,N_15323,N_15035);
nand U15819 (N_15819,N_15425,N_15598);
or U15820 (N_15820,N_15243,N_15421);
or U15821 (N_15821,N_15476,N_15595);
or U15822 (N_15822,N_15530,N_15058);
and U15823 (N_15823,N_15267,N_15051);
xnor U15824 (N_15824,N_15219,N_15376);
and U15825 (N_15825,N_15349,N_15195);
xor U15826 (N_15826,N_15168,N_15177);
xor U15827 (N_15827,N_15458,N_15341);
and U15828 (N_15828,N_15162,N_15252);
nand U15829 (N_15829,N_15158,N_15358);
and U15830 (N_15830,N_15347,N_15350);
xnor U15831 (N_15831,N_15099,N_15076);
or U15832 (N_15832,N_15455,N_15134);
xor U15833 (N_15833,N_15240,N_15578);
xor U15834 (N_15834,N_15441,N_15551);
nor U15835 (N_15835,N_15593,N_15364);
xor U15836 (N_15836,N_15268,N_15142);
or U15837 (N_15837,N_15229,N_15565);
or U15838 (N_15838,N_15459,N_15357);
or U15839 (N_15839,N_15208,N_15342);
or U15840 (N_15840,N_15048,N_15170);
nor U15841 (N_15841,N_15135,N_15326);
nor U15842 (N_15842,N_15536,N_15445);
xnor U15843 (N_15843,N_15223,N_15301);
xnor U15844 (N_15844,N_15466,N_15333);
nand U15845 (N_15845,N_15576,N_15561);
and U15846 (N_15846,N_15103,N_15499);
or U15847 (N_15847,N_15291,N_15075);
nand U15848 (N_15848,N_15329,N_15128);
xnor U15849 (N_15849,N_15383,N_15394);
nor U15850 (N_15850,N_15491,N_15302);
nor U15851 (N_15851,N_15420,N_15407);
xor U15852 (N_15852,N_15273,N_15450);
or U15853 (N_15853,N_15021,N_15388);
nor U15854 (N_15854,N_15257,N_15512);
xnor U15855 (N_15855,N_15484,N_15433);
xor U15856 (N_15856,N_15218,N_15073);
xor U15857 (N_15857,N_15042,N_15089);
and U15858 (N_15858,N_15463,N_15080);
or U15859 (N_15859,N_15372,N_15305);
and U15860 (N_15860,N_15365,N_15059);
xor U15861 (N_15861,N_15366,N_15575);
or U15862 (N_15862,N_15034,N_15293);
xnor U15863 (N_15863,N_15001,N_15041);
and U15864 (N_15864,N_15004,N_15495);
nand U15865 (N_15865,N_15258,N_15439);
nand U15866 (N_15866,N_15231,N_15478);
xnor U15867 (N_15867,N_15114,N_15573);
or U15868 (N_15868,N_15390,N_15431);
nand U15869 (N_15869,N_15083,N_15361);
nand U15870 (N_15870,N_15415,N_15435);
nand U15871 (N_15871,N_15017,N_15130);
or U15872 (N_15872,N_15587,N_15055);
and U15873 (N_15873,N_15304,N_15149);
or U15874 (N_15874,N_15278,N_15259);
or U15875 (N_15875,N_15555,N_15217);
nand U15876 (N_15876,N_15294,N_15477);
nand U15877 (N_15877,N_15553,N_15544);
xnor U15878 (N_15878,N_15360,N_15253);
or U15879 (N_15879,N_15429,N_15308);
nor U15880 (N_15880,N_15592,N_15097);
nor U15881 (N_15881,N_15260,N_15296);
nand U15882 (N_15882,N_15164,N_15002);
nor U15883 (N_15883,N_15462,N_15054);
nor U15884 (N_15884,N_15332,N_15280);
nor U15885 (N_15885,N_15181,N_15150);
xor U15886 (N_15886,N_15256,N_15521);
nor U15887 (N_15887,N_15428,N_15306);
nor U15888 (N_15888,N_15247,N_15272);
and U15889 (N_15889,N_15490,N_15071);
nand U15890 (N_15890,N_15045,N_15444);
nand U15891 (N_15891,N_15072,N_15446);
xor U15892 (N_15892,N_15504,N_15050);
xnor U15893 (N_15893,N_15085,N_15220);
and U15894 (N_15894,N_15417,N_15224);
and U15895 (N_15895,N_15570,N_15107);
nor U15896 (N_15896,N_15186,N_15416);
and U15897 (N_15897,N_15399,N_15481);
and U15898 (N_15898,N_15171,N_15145);
nand U15899 (N_15899,N_15026,N_15447);
xor U15900 (N_15900,N_15277,N_15456);
nand U15901 (N_15901,N_15146,N_15098);
nor U15902 (N_15902,N_15452,N_15390);
xnor U15903 (N_15903,N_15503,N_15540);
xnor U15904 (N_15904,N_15126,N_15368);
nor U15905 (N_15905,N_15004,N_15053);
and U15906 (N_15906,N_15042,N_15538);
or U15907 (N_15907,N_15366,N_15440);
nand U15908 (N_15908,N_15434,N_15292);
or U15909 (N_15909,N_15212,N_15171);
and U15910 (N_15910,N_15189,N_15463);
and U15911 (N_15911,N_15503,N_15396);
and U15912 (N_15912,N_15070,N_15202);
nor U15913 (N_15913,N_15373,N_15594);
nand U15914 (N_15914,N_15298,N_15078);
nor U15915 (N_15915,N_15531,N_15365);
or U15916 (N_15916,N_15231,N_15352);
and U15917 (N_15917,N_15476,N_15095);
nand U15918 (N_15918,N_15241,N_15151);
and U15919 (N_15919,N_15528,N_15181);
nor U15920 (N_15920,N_15451,N_15521);
xor U15921 (N_15921,N_15480,N_15536);
nand U15922 (N_15922,N_15240,N_15515);
or U15923 (N_15923,N_15435,N_15554);
and U15924 (N_15924,N_15202,N_15143);
nor U15925 (N_15925,N_15169,N_15486);
nand U15926 (N_15926,N_15152,N_15416);
nor U15927 (N_15927,N_15454,N_15222);
xnor U15928 (N_15928,N_15207,N_15592);
nand U15929 (N_15929,N_15404,N_15140);
and U15930 (N_15930,N_15166,N_15486);
or U15931 (N_15931,N_15569,N_15482);
nor U15932 (N_15932,N_15459,N_15018);
xnor U15933 (N_15933,N_15258,N_15503);
xor U15934 (N_15934,N_15435,N_15362);
and U15935 (N_15935,N_15098,N_15351);
nand U15936 (N_15936,N_15024,N_15541);
xor U15937 (N_15937,N_15440,N_15584);
xnor U15938 (N_15938,N_15288,N_15446);
nand U15939 (N_15939,N_15584,N_15281);
or U15940 (N_15940,N_15292,N_15000);
nand U15941 (N_15941,N_15485,N_15170);
xor U15942 (N_15942,N_15181,N_15393);
or U15943 (N_15943,N_15430,N_15525);
or U15944 (N_15944,N_15147,N_15455);
xor U15945 (N_15945,N_15355,N_15175);
and U15946 (N_15946,N_15525,N_15425);
or U15947 (N_15947,N_15405,N_15278);
xor U15948 (N_15948,N_15088,N_15148);
nor U15949 (N_15949,N_15180,N_15375);
and U15950 (N_15950,N_15595,N_15374);
or U15951 (N_15951,N_15028,N_15078);
xnor U15952 (N_15952,N_15542,N_15326);
and U15953 (N_15953,N_15227,N_15116);
nor U15954 (N_15954,N_15444,N_15079);
xnor U15955 (N_15955,N_15250,N_15574);
xor U15956 (N_15956,N_15563,N_15585);
nor U15957 (N_15957,N_15243,N_15057);
xnor U15958 (N_15958,N_15455,N_15259);
xor U15959 (N_15959,N_15043,N_15458);
nor U15960 (N_15960,N_15430,N_15213);
nor U15961 (N_15961,N_15056,N_15243);
or U15962 (N_15962,N_15159,N_15581);
and U15963 (N_15963,N_15048,N_15316);
xor U15964 (N_15964,N_15437,N_15568);
or U15965 (N_15965,N_15124,N_15519);
nor U15966 (N_15966,N_15116,N_15383);
xor U15967 (N_15967,N_15319,N_15350);
nor U15968 (N_15968,N_15038,N_15177);
nor U15969 (N_15969,N_15423,N_15439);
xor U15970 (N_15970,N_15194,N_15088);
and U15971 (N_15971,N_15240,N_15228);
and U15972 (N_15972,N_15062,N_15518);
nand U15973 (N_15973,N_15311,N_15347);
and U15974 (N_15974,N_15038,N_15035);
or U15975 (N_15975,N_15326,N_15440);
or U15976 (N_15976,N_15156,N_15009);
nor U15977 (N_15977,N_15389,N_15193);
and U15978 (N_15978,N_15292,N_15233);
nor U15979 (N_15979,N_15230,N_15422);
nand U15980 (N_15980,N_15282,N_15219);
and U15981 (N_15981,N_15223,N_15440);
and U15982 (N_15982,N_15259,N_15221);
xnor U15983 (N_15983,N_15355,N_15387);
nor U15984 (N_15984,N_15423,N_15547);
nor U15985 (N_15985,N_15040,N_15015);
xor U15986 (N_15986,N_15115,N_15587);
xnor U15987 (N_15987,N_15365,N_15573);
and U15988 (N_15988,N_15520,N_15097);
nor U15989 (N_15989,N_15093,N_15502);
and U15990 (N_15990,N_15578,N_15495);
or U15991 (N_15991,N_15211,N_15432);
and U15992 (N_15992,N_15438,N_15058);
xor U15993 (N_15993,N_15574,N_15314);
nand U15994 (N_15994,N_15118,N_15064);
or U15995 (N_15995,N_15572,N_15585);
or U15996 (N_15996,N_15095,N_15327);
nor U15997 (N_15997,N_15479,N_15553);
nand U15998 (N_15998,N_15348,N_15203);
and U15999 (N_15999,N_15565,N_15156);
or U16000 (N_16000,N_15374,N_15026);
nor U16001 (N_16001,N_15459,N_15195);
and U16002 (N_16002,N_15373,N_15051);
nand U16003 (N_16003,N_15448,N_15568);
xnor U16004 (N_16004,N_15378,N_15239);
xor U16005 (N_16005,N_15307,N_15089);
or U16006 (N_16006,N_15143,N_15193);
xnor U16007 (N_16007,N_15351,N_15039);
nand U16008 (N_16008,N_15031,N_15097);
nor U16009 (N_16009,N_15209,N_15014);
or U16010 (N_16010,N_15266,N_15171);
xor U16011 (N_16011,N_15526,N_15492);
nand U16012 (N_16012,N_15058,N_15488);
xnor U16013 (N_16013,N_15358,N_15408);
nor U16014 (N_16014,N_15031,N_15048);
xor U16015 (N_16015,N_15061,N_15311);
and U16016 (N_16016,N_15427,N_15253);
xor U16017 (N_16017,N_15537,N_15182);
or U16018 (N_16018,N_15049,N_15495);
and U16019 (N_16019,N_15156,N_15287);
and U16020 (N_16020,N_15066,N_15016);
or U16021 (N_16021,N_15516,N_15570);
nand U16022 (N_16022,N_15179,N_15298);
and U16023 (N_16023,N_15060,N_15342);
xnor U16024 (N_16024,N_15002,N_15498);
and U16025 (N_16025,N_15471,N_15587);
and U16026 (N_16026,N_15469,N_15554);
and U16027 (N_16027,N_15512,N_15244);
or U16028 (N_16028,N_15057,N_15029);
or U16029 (N_16029,N_15420,N_15073);
and U16030 (N_16030,N_15111,N_15451);
nand U16031 (N_16031,N_15598,N_15432);
and U16032 (N_16032,N_15143,N_15557);
xor U16033 (N_16033,N_15073,N_15549);
or U16034 (N_16034,N_15485,N_15329);
nand U16035 (N_16035,N_15029,N_15367);
xor U16036 (N_16036,N_15242,N_15177);
nand U16037 (N_16037,N_15194,N_15329);
xor U16038 (N_16038,N_15254,N_15185);
nand U16039 (N_16039,N_15236,N_15202);
xnor U16040 (N_16040,N_15488,N_15577);
and U16041 (N_16041,N_15559,N_15557);
nand U16042 (N_16042,N_15509,N_15103);
xnor U16043 (N_16043,N_15040,N_15386);
or U16044 (N_16044,N_15036,N_15309);
nand U16045 (N_16045,N_15059,N_15499);
nor U16046 (N_16046,N_15469,N_15095);
and U16047 (N_16047,N_15450,N_15425);
xnor U16048 (N_16048,N_15059,N_15109);
nand U16049 (N_16049,N_15294,N_15302);
or U16050 (N_16050,N_15363,N_15552);
xor U16051 (N_16051,N_15080,N_15466);
and U16052 (N_16052,N_15595,N_15199);
nand U16053 (N_16053,N_15539,N_15013);
nor U16054 (N_16054,N_15396,N_15401);
xor U16055 (N_16055,N_15581,N_15184);
or U16056 (N_16056,N_15259,N_15569);
nand U16057 (N_16057,N_15094,N_15563);
and U16058 (N_16058,N_15422,N_15196);
nor U16059 (N_16059,N_15261,N_15040);
nor U16060 (N_16060,N_15027,N_15471);
nor U16061 (N_16061,N_15262,N_15549);
nand U16062 (N_16062,N_15104,N_15294);
nand U16063 (N_16063,N_15323,N_15283);
nand U16064 (N_16064,N_15359,N_15129);
xor U16065 (N_16065,N_15176,N_15064);
and U16066 (N_16066,N_15129,N_15243);
nand U16067 (N_16067,N_15459,N_15392);
xor U16068 (N_16068,N_15135,N_15582);
xor U16069 (N_16069,N_15102,N_15176);
or U16070 (N_16070,N_15265,N_15307);
nand U16071 (N_16071,N_15396,N_15346);
nand U16072 (N_16072,N_15228,N_15291);
nand U16073 (N_16073,N_15234,N_15091);
nor U16074 (N_16074,N_15240,N_15133);
nor U16075 (N_16075,N_15546,N_15329);
and U16076 (N_16076,N_15527,N_15478);
nand U16077 (N_16077,N_15176,N_15248);
xnor U16078 (N_16078,N_15517,N_15545);
or U16079 (N_16079,N_15416,N_15362);
nand U16080 (N_16080,N_15366,N_15162);
and U16081 (N_16081,N_15278,N_15437);
or U16082 (N_16082,N_15110,N_15410);
xor U16083 (N_16083,N_15499,N_15418);
nand U16084 (N_16084,N_15324,N_15483);
nor U16085 (N_16085,N_15453,N_15574);
nor U16086 (N_16086,N_15140,N_15113);
xor U16087 (N_16087,N_15586,N_15191);
or U16088 (N_16088,N_15532,N_15426);
xnor U16089 (N_16089,N_15559,N_15084);
nor U16090 (N_16090,N_15422,N_15338);
xnor U16091 (N_16091,N_15407,N_15327);
and U16092 (N_16092,N_15439,N_15429);
xor U16093 (N_16093,N_15448,N_15351);
and U16094 (N_16094,N_15065,N_15190);
nand U16095 (N_16095,N_15166,N_15566);
nor U16096 (N_16096,N_15486,N_15274);
and U16097 (N_16097,N_15353,N_15226);
and U16098 (N_16098,N_15325,N_15427);
xnor U16099 (N_16099,N_15267,N_15531);
or U16100 (N_16100,N_15263,N_15391);
xnor U16101 (N_16101,N_15269,N_15332);
and U16102 (N_16102,N_15086,N_15231);
xor U16103 (N_16103,N_15225,N_15091);
xnor U16104 (N_16104,N_15061,N_15257);
nor U16105 (N_16105,N_15253,N_15550);
nand U16106 (N_16106,N_15251,N_15495);
xor U16107 (N_16107,N_15010,N_15443);
or U16108 (N_16108,N_15332,N_15450);
and U16109 (N_16109,N_15454,N_15332);
or U16110 (N_16110,N_15501,N_15561);
and U16111 (N_16111,N_15437,N_15233);
or U16112 (N_16112,N_15422,N_15449);
nor U16113 (N_16113,N_15345,N_15599);
or U16114 (N_16114,N_15549,N_15054);
nor U16115 (N_16115,N_15133,N_15408);
nor U16116 (N_16116,N_15474,N_15264);
or U16117 (N_16117,N_15266,N_15521);
or U16118 (N_16118,N_15468,N_15230);
nor U16119 (N_16119,N_15004,N_15231);
and U16120 (N_16120,N_15204,N_15107);
and U16121 (N_16121,N_15401,N_15237);
nor U16122 (N_16122,N_15012,N_15496);
nor U16123 (N_16123,N_15384,N_15190);
nand U16124 (N_16124,N_15261,N_15053);
nor U16125 (N_16125,N_15157,N_15462);
nor U16126 (N_16126,N_15084,N_15056);
and U16127 (N_16127,N_15596,N_15445);
or U16128 (N_16128,N_15365,N_15168);
and U16129 (N_16129,N_15292,N_15106);
nand U16130 (N_16130,N_15476,N_15453);
xnor U16131 (N_16131,N_15100,N_15546);
xor U16132 (N_16132,N_15250,N_15416);
xnor U16133 (N_16133,N_15060,N_15382);
and U16134 (N_16134,N_15068,N_15039);
nor U16135 (N_16135,N_15309,N_15181);
and U16136 (N_16136,N_15216,N_15239);
xor U16137 (N_16137,N_15044,N_15182);
and U16138 (N_16138,N_15192,N_15207);
nand U16139 (N_16139,N_15113,N_15329);
or U16140 (N_16140,N_15048,N_15377);
nor U16141 (N_16141,N_15505,N_15367);
xnor U16142 (N_16142,N_15151,N_15308);
nor U16143 (N_16143,N_15390,N_15388);
nor U16144 (N_16144,N_15460,N_15422);
nand U16145 (N_16145,N_15459,N_15368);
and U16146 (N_16146,N_15081,N_15312);
or U16147 (N_16147,N_15062,N_15504);
or U16148 (N_16148,N_15065,N_15462);
nor U16149 (N_16149,N_15015,N_15021);
or U16150 (N_16150,N_15000,N_15358);
and U16151 (N_16151,N_15584,N_15492);
xor U16152 (N_16152,N_15173,N_15017);
nand U16153 (N_16153,N_15230,N_15052);
nand U16154 (N_16154,N_15213,N_15104);
nand U16155 (N_16155,N_15172,N_15286);
or U16156 (N_16156,N_15122,N_15348);
nand U16157 (N_16157,N_15471,N_15046);
or U16158 (N_16158,N_15072,N_15232);
nand U16159 (N_16159,N_15588,N_15150);
nor U16160 (N_16160,N_15316,N_15574);
nand U16161 (N_16161,N_15110,N_15302);
xor U16162 (N_16162,N_15584,N_15061);
nor U16163 (N_16163,N_15390,N_15011);
xor U16164 (N_16164,N_15210,N_15236);
or U16165 (N_16165,N_15022,N_15577);
nor U16166 (N_16166,N_15163,N_15263);
nor U16167 (N_16167,N_15387,N_15460);
and U16168 (N_16168,N_15549,N_15582);
or U16169 (N_16169,N_15108,N_15415);
nor U16170 (N_16170,N_15180,N_15286);
nor U16171 (N_16171,N_15000,N_15462);
or U16172 (N_16172,N_15485,N_15308);
nor U16173 (N_16173,N_15260,N_15173);
nor U16174 (N_16174,N_15351,N_15264);
and U16175 (N_16175,N_15256,N_15486);
nor U16176 (N_16176,N_15025,N_15147);
nor U16177 (N_16177,N_15036,N_15491);
nor U16178 (N_16178,N_15160,N_15491);
xnor U16179 (N_16179,N_15476,N_15438);
xnor U16180 (N_16180,N_15111,N_15013);
nand U16181 (N_16181,N_15572,N_15546);
nand U16182 (N_16182,N_15134,N_15423);
or U16183 (N_16183,N_15404,N_15373);
xnor U16184 (N_16184,N_15267,N_15078);
xnor U16185 (N_16185,N_15493,N_15327);
or U16186 (N_16186,N_15108,N_15462);
xor U16187 (N_16187,N_15276,N_15014);
nand U16188 (N_16188,N_15212,N_15039);
nand U16189 (N_16189,N_15271,N_15460);
and U16190 (N_16190,N_15446,N_15285);
nand U16191 (N_16191,N_15100,N_15255);
nor U16192 (N_16192,N_15128,N_15411);
and U16193 (N_16193,N_15211,N_15166);
xor U16194 (N_16194,N_15073,N_15592);
and U16195 (N_16195,N_15447,N_15217);
or U16196 (N_16196,N_15421,N_15466);
nand U16197 (N_16197,N_15322,N_15246);
or U16198 (N_16198,N_15403,N_15119);
and U16199 (N_16199,N_15021,N_15296);
xnor U16200 (N_16200,N_15676,N_15876);
nand U16201 (N_16201,N_15942,N_15687);
xor U16202 (N_16202,N_16114,N_15672);
and U16203 (N_16203,N_16175,N_15803);
xnor U16204 (N_16204,N_15768,N_15807);
xnor U16205 (N_16205,N_15700,N_16132);
xnor U16206 (N_16206,N_15841,N_15826);
xnor U16207 (N_16207,N_16145,N_16079);
and U16208 (N_16208,N_16089,N_15724);
or U16209 (N_16209,N_15954,N_15656);
or U16210 (N_16210,N_15974,N_16118);
nor U16211 (N_16211,N_16099,N_16066);
nand U16212 (N_16212,N_15635,N_15604);
and U16213 (N_16213,N_15613,N_15994);
nor U16214 (N_16214,N_15797,N_15885);
nor U16215 (N_16215,N_15977,N_16037);
or U16216 (N_16216,N_15630,N_16000);
or U16217 (N_16217,N_16002,N_16019);
or U16218 (N_16218,N_15991,N_16195);
nand U16219 (N_16219,N_15927,N_15909);
xor U16220 (N_16220,N_15739,N_15867);
xnor U16221 (N_16221,N_16008,N_15605);
xor U16222 (N_16222,N_16108,N_16029);
and U16223 (N_16223,N_16072,N_15930);
and U16224 (N_16224,N_15881,N_15935);
or U16225 (N_16225,N_15607,N_15822);
or U16226 (N_16226,N_15821,N_16119);
nor U16227 (N_16227,N_15884,N_15854);
or U16228 (N_16228,N_15983,N_15618);
and U16229 (N_16229,N_15666,N_15784);
or U16230 (N_16230,N_15888,N_15653);
or U16231 (N_16231,N_15736,N_15939);
or U16232 (N_16232,N_15777,N_16182);
or U16233 (N_16233,N_15626,N_16070);
or U16234 (N_16234,N_15809,N_15861);
nand U16235 (N_16235,N_15926,N_15608);
nor U16236 (N_16236,N_15916,N_15793);
and U16237 (N_16237,N_16142,N_15897);
and U16238 (N_16238,N_15721,N_16125);
nand U16239 (N_16239,N_16170,N_15889);
nor U16240 (N_16240,N_15898,N_15691);
or U16241 (N_16241,N_16104,N_15675);
or U16242 (N_16242,N_15755,N_15840);
xnor U16243 (N_16243,N_15832,N_15874);
xor U16244 (N_16244,N_16107,N_15622);
nand U16245 (N_16245,N_15764,N_15895);
and U16246 (N_16246,N_16196,N_15998);
xnor U16247 (N_16247,N_15749,N_15640);
xor U16248 (N_16248,N_16111,N_15911);
xor U16249 (N_16249,N_15789,N_15646);
nor U16250 (N_16250,N_15649,N_15719);
nand U16251 (N_16251,N_16188,N_15752);
and U16252 (N_16252,N_15946,N_16160);
nand U16253 (N_16253,N_15726,N_15924);
nor U16254 (N_16254,N_15880,N_16046);
xnor U16255 (N_16255,N_16096,N_16052);
or U16256 (N_16256,N_15709,N_15728);
nor U16257 (N_16257,N_15651,N_15735);
or U16258 (N_16258,N_15667,N_15718);
nor U16259 (N_16259,N_15733,N_15619);
nand U16260 (N_16260,N_15714,N_16007);
nand U16261 (N_16261,N_16097,N_16130);
and U16262 (N_16262,N_15883,N_15668);
and U16263 (N_16263,N_15993,N_16167);
nor U16264 (N_16264,N_16058,N_15695);
xnor U16265 (N_16265,N_16056,N_15770);
xor U16266 (N_16266,N_16082,N_15810);
nand U16267 (N_16267,N_15844,N_15843);
or U16268 (N_16268,N_15694,N_15999);
nand U16269 (N_16269,N_16069,N_16087);
and U16270 (N_16270,N_16060,N_15616);
or U16271 (N_16271,N_15869,N_16077);
nor U16272 (N_16272,N_15917,N_16185);
and U16273 (N_16273,N_15959,N_15873);
nor U16274 (N_16274,N_15658,N_16115);
nand U16275 (N_16275,N_16031,N_15818);
xnor U16276 (N_16276,N_15820,N_16038);
or U16277 (N_16277,N_15940,N_16173);
nor U16278 (N_16278,N_15716,N_15913);
xnor U16279 (N_16279,N_16146,N_15890);
nor U16280 (N_16280,N_16152,N_15972);
nor U16281 (N_16281,N_15836,N_15894);
nand U16282 (N_16282,N_15919,N_15707);
and U16283 (N_16283,N_15842,N_15967);
nor U16284 (N_16284,N_16003,N_15837);
xnor U16285 (N_16285,N_15957,N_15754);
nor U16286 (N_16286,N_15688,N_16187);
and U16287 (N_16287,N_16006,N_15962);
xnor U16288 (N_16288,N_15979,N_15690);
and U16289 (N_16289,N_15639,N_16078);
nor U16290 (N_16290,N_15720,N_15738);
xnor U16291 (N_16291,N_16080,N_16180);
and U16292 (N_16292,N_15971,N_16061);
nand U16293 (N_16293,N_15730,N_15617);
nor U16294 (N_16294,N_15717,N_16179);
xnor U16295 (N_16295,N_16035,N_15796);
or U16296 (N_16296,N_15711,N_15624);
and U16297 (N_16297,N_16050,N_15771);
or U16298 (N_16298,N_15875,N_15931);
nor U16299 (N_16299,N_15813,N_15737);
nor U16300 (N_16300,N_16085,N_15902);
or U16301 (N_16301,N_15955,N_16098);
nor U16302 (N_16302,N_16094,N_15634);
nand U16303 (N_16303,N_15965,N_15825);
and U16304 (N_16304,N_15627,N_15664);
or U16305 (N_16305,N_15702,N_16015);
nor U16306 (N_16306,N_15838,N_15950);
xor U16307 (N_16307,N_16064,N_16122);
xnor U16308 (N_16308,N_15910,N_16168);
nor U16309 (N_16309,N_16140,N_15781);
nor U16310 (N_16310,N_15743,N_15985);
nor U16311 (N_16311,N_15703,N_15681);
nand U16312 (N_16312,N_15636,N_15866);
xnor U16313 (N_16313,N_16148,N_15907);
or U16314 (N_16314,N_15872,N_15833);
nor U16315 (N_16315,N_15632,N_15899);
and U16316 (N_16316,N_16149,N_15693);
nor U16317 (N_16317,N_15868,N_15980);
and U16318 (N_16318,N_15767,N_16101);
nand U16319 (N_16319,N_15683,N_16171);
nor U16320 (N_16320,N_16163,N_16156);
xnor U16321 (N_16321,N_16113,N_15637);
or U16322 (N_16322,N_15644,N_15712);
or U16323 (N_16323,N_15677,N_15660);
xnor U16324 (N_16324,N_16092,N_15629);
or U16325 (N_16325,N_15643,N_15633);
or U16326 (N_16326,N_15828,N_15747);
or U16327 (N_16327,N_15882,N_15699);
nor U16328 (N_16328,N_15773,N_16161);
or U16329 (N_16329,N_15900,N_16040);
nor U16330 (N_16330,N_16110,N_16041);
and U16331 (N_16331,N_15988,N_16053);
or U16332 (N_16332,N_15887,N_15751);
nor U16333 (N_16333,N_16004,N_16158);
or U16334 (N_16334,N_16018,N_15800);
nor U16335 (N_16335,N_15679,N_15745);
nor U16336 (N_16336,N_15976,N_16048);
or U16337 (N_16337,N_15775,N_15760);
and U16338 (N_16338,N_16021,N_15995);
and U16339 (N_16339,N_15665,N_16090);
xnor U16340 (N_16340,N_15852,N_16164);
xor U16341 (N_16341,N_15731,N_15798);
or U16342 (N_16342,N_15706,N_16009);
xor U16343 (N_16343,N_15951,N_15704);
xnor U16344 (N_16344,N_15830,N_15949);
and U16345 (N_16345,N_15641,N_15615);
and U16346 (N_16346,N_15863,N_15848);
xor U16347 (N_16347,N_15982,N_16150);
nor U16348 (N_16348,N_15602,N_16076);
nand U16349 (N_16349,N_16049,N_16102);
nand U16350 (N_16350,N_16131,N_16023);
xnor U16351 (N_16351,N_15878,N_16190);
xnor U16352 (N_16352,N_16042,N_16106);
nand U16353 (N_16353,N_16117,N_15879);
or U16354 (N_16354,N_16121,N_15970);
nand U16355 (N_16355,N_16025,N_16138);
nand U16356 (N_16356,N_16026,N_15765);
nor U16357 (N_16357,N_16093,N_16075);
xor U16358 (N_16358,N_15834,N_16024);
nor U16359 (N_16359,N_16045,N_15824);
and U16360 (N_16360,N_15722,N_15891);
nand U16361 (N_16361,N_16177,N_15662);
nor U16362 (N_16362,N_15984,N_16169);
nor U16363 (N_16363,N_15686,N_15859);
and U16364 (N_16364,N_16012,N_16027);
nand U16365 (N_16365,N_15996,N_15723);
nand U16366 (N_16366,N_16189,N_15932);
nor U16367 (N_16367,N_16095,N_16137);
nand U16368 (N_16368,N_15758,N_15941);
nor U16369 (N_16369,N_16028,N_15975);
nand U16370 (N_16370,N_15621,N_15601);
nand U16371 (N_16371,N_16051,N_15936);
and U16372 (N_16372,N_15966,N_15992);
or U16373 (N_16373,N_15925,N_15914);
nand U16374 (N_16374,N_16192,N_15968);
nand U16375 (N_16375,N_16186,N_15638);
or U16376 (N_16376,N_15877,N_15892);
xnor U16377 (N_16377,N_15990,N_16126);
nand U16378 (N_16378,N_15657,N_15774);
and U16379 (N_16379,N_15857,N_15670);
nand U16380 (N_16380,N_16071,N_16005);
and U16381 (N_16381,N_16047,N_15792);
nand U16382 (N_16382,N_15835,N_16063);
nor U16383 (N_16383,N_15997,N_16105);
nand U16384 (N_16384,N_16184,N_15948);
xor U16385 (N_16385,N_15987,N_16151);
and U16386 (N_16386,N_16181,N_16043);
nand U16387 (N_16387,N_16074,N_16030);
and U16388 (N_16388,N_15631,N_15870);
or U16389 (N_16389,N_15614,N_15969);
xnor U16390 (N_16390,N_15741,N_15928);
nor U16391 (N_16391,N_15696,N_16103);
xnor U16392 (N_16392,N_15804,N_15960);
and U16393 (N_16393,N_16127,N_15801);
nand U16394 (N_16394,N_15905,N_15645);
or U16395 (N_16395,N_15827,N_15839);
nand U16396 (N_16396,N_16044,N_16016);
nor U16397 (N_16397,N_16055,N_15851);
or U16398 (N_16398,N_15746,N_15692);
and U16399 (N_16399,N_16193,N_15655);
nor U16400 (N_16400,N_16141,N_15734);
nor U16401 (N_16401,N_16155,N_15915);
xor U16402 (N_16402,N_15938,N_15871);
xnor U16403 (N_16403,N_16083,N_15811);
xnor U16404 (N_16404,N_16086,N_16123);
nor U16405 (N_16405,N_15860,N_15756);
nor U16406 (N_16406,N_16174,N_15964);
nor U16407 (N_16407,N_16065,N_15762);
nor U16408 (N_16408,N_15937,N_15893);
xor U16409 (N_16409,N_15846,N_16194);
nor U16410 (N_16410,N_16199,N_15989);
or U16411 (N_16411,N_16153,N_16081);
nor U16412 (N_16412,N_16014,N_16036);
or U16413 (N_16413,N_15849,N_16162);
nand U16414 (N_16414,N_16134,N_15786);
or U16415 (N_16415,N_15750,N_15705);
nand U16416 (N_16416,N_16147,N_15823);
or U16417 (N_16417,N_15654,N_15904);
and U16418 (N_16418,N_15761,N_16197);
xor U16419 (N_16419,N_15780,N_15865);
nor U16420 (N_16420,N_15701,N_15682);
nor U16421 (N_16421,N_15732,N_15956);
or U16422 (N_16422,N_15603,N_15669);
and U16423 (N_16423,N_15791,N_15790);
xnor U16424 (N_16424,N_15923,N_15611);
or U16425 (N_16425,N_15986,N_15708);
xnor U16426 (N_16426,N_15788,N_16176);
xnor U16427 (N_16427,N_15772,N_16178);
xnor U16428 (N_16428,N_15906,N_15815);
nor U16429 (N_16429,N_15945,N_16135);
and U16430 (N_16430,N_15862,N_15819);
or U16431 (N_16431,N_15831,N_16054);
nand U16432 (N_16432,N_15778,N_15921);
and U16433 (N_16433,N_16057,N_15961);
and U16434 (N_16434,N_15678,N_15886);
and U16435 (N_16435,N_15753,N_16020);
nand U16436 (N_16436,N_15689,N_16011);
and U16437 (N_16437,N_15684,N_15783);
and U16438 (N_16438,N_16166,N_15609);
or U16439 (N_16439,N_15606,N_15958);
nor U16440 (N_16440,N_15806,N_15934);
and U16441 (N_16441,N_16157,N_16084);
nor U16442 (N_16442,N_15744,N_15953);
or U16443 (N_16443,N_15725,N_16088);
xnor U16444 (N_16444,N_15795,N_15787);
nand U16445 (N_16445,N_16133,N_16143);
and U16446 (N_16446,N_15901,N_16059);
nor U16447 (N_16447,N_15929,N_15612);
and U16448 (N_16448,N_16120,N_16010);
or U16449 (N_16449,N_16165,N_15808);
or U16450 (N_16450,N_16159,N_16100);
or U16451 (N_16451,N_16068,N_15673);
nand U16452 (N_16452,N_15600,N_15785);
xor U16453 (N_16453,N_15715,N_15650);
or U16454 (N_16454,N_15671,N_15981);
and U16455 (N_16455,N_15748,N_15661);
nor U16456 (N_16456,N_15620,N_15652);
nor U16457 (N_16457,N_15740,N_16073);
xor U16458 (N_16458,N_15978,N_15944);
nand U16459 (N_16459,N_16172,N_16033);
xor U16460 (N_16460,N_16198,N_15896);
nand U16461 (N_16461,N_16013,N_15685);
or U16462 (N_16462,N_16139,N_16034);
and U16463 (N_16463,N_15757,N_16109);
xnor U16464 (N_16464,N_15698,N_15952);
nor U16465 (N_16465,N_16116,N_16022);
nor U16466 (N_16466,N_16032,N_16191);
and U16467 (N_16467,N_15727,N_15648);
and U16468 (N_16468,N_16154,N_15853);
xor U16469 (N_16469,N_15623,N_15794);
or U16470 (N_16470,N_15829,N_15855);
or U16471 (N_16471,N_15812,N_15628);
or U16472 (N_16472,N_15817,N_15912);
nor U16473 (N_16473,N_15816,N_16112);
nor U16474 (N_16474,N_15729,N_15610);
nand U16475 (N_16475,N_15742,N_15766);
nor U16476 (N_16476,N_15759,N_15805);
and U16477 (N_16477,N_15659,N_16124);
and U16478 (N_16478,N_16039,N_15973);
or U16479 (N_16479,N_15763,N_15779);
nand U16480 (N_16480,N_16017,N_15908);
xor U16481 (N_16481,N_16136,N_15814);
xnor U16482 (N_16482,N_15680,N_15856);
and U16483 (N_16483,N_15864,N_15625);
xor U16484 (N_16484,N_15799,N_16183);
nand U16485 (N_16485,N_15918,N_15663);
and U16486 (N_16486,N_15674,N_15710);
nor U16487 (N_16487,N_15963,N_15713);
and U16488 (N_16488,N_15850,N_15903);
and U16489 (N_16489,N_16129,N_15647);
nor U16490 (N_16490,N_16062,N_15947);
or U16491 (N_16491,N_15802,N_16144);
nor U16492 (N_16492,N_15847,N_16001);
nand U16493 (N_16493,N_16128,N_16067);
and U16494 (N_16494,N_15922,N_15642);
nand U16495 (N_16495,N_15933,N_15858);
nor U16496 (N_16496,N_15769,N_15920);
nor U16497 (N_16497,N_15943,N_15776);
nand U16498 (N_16498,N_15845,N_15697);
and U16499 (N_16499,N_16091,N_15782);
xor U16500 (N_16500,N_16147,N_16000);
xnor U16501 (N_16501,N_16100,N_15753);
nand U16502 (N_16502,N_16094,N_15941);
nand U16503 (N_16503,N_16008,N_16131);
xor U16504 (N_16504,N_15670,N_15667);
xnor U16505 (N_16505,N_15810,N_15991);
xnor U16506 (N_16506,N_15921,N_16126);
nand U16507 (N_16507,N_16134,N_16141);
nand U16508 (N_16508,N_16025,N_15835);
or U16509 (N_16509,N_15864,N_15691);
and U16510 (N_16510,N_16069,N_15829);
and U16511 (N_16511,N_16068,N_15897);
xnor U16512 (N_16512,N_15866,N_16156);
xor U16513 (N_16513,N_15630,N_15647);
or U16514 (N_16514,N_16174,N_16123);
xnor U16515 (N_16515,N_15796,N_16077);
nor U16516 (N_16516,N_16137,N_15855);
xnor U16517 (N_16517,N_15655,N_16151);
xor U16518 (N_16518,N_16058,N_15749);
xor U16519 (N_16519,N_15990,N_16053);
nand U16520 (N_16520,N_15844,N_15800);
nor U16521 (N_16521,N_15914,N_16189);
xor U16522 (N_16522,N_15851,N_16042);
xnor U16523 (N_16523,N_15790,N_15836);
or U16524 (N_16524,N_15653,N_15791);
xnor U16525 (N_16525,N_16073,N_15941);
and U16526 (N_16526,N_15946,N_15866);
or U16527 (N_16527,N_15613,N_15736);
or U16528 (N_16528,N_15607,N_16030);
nand U16529 (N_16529,N_16168,N_15646);
nor U16530 (N_16530,N_16104,N_16144);
nand U16531 (N_16531,N_15768,N_16118);
xnor U16532 (N_16532,N_15882,N_15787);
and U16533 (N_16533,N_16070,N_15627);
or U16534 (N_16534,N_15722,N_15813);
xnor U16535 (N_16535,N_15886,N_15782);
nand U16536 (N_16536,N_16111,N_16031);
xor U16537 (N_16537,N_15791,N_16183);
or U16538 (N_16538,N_16048,N_16143);
nand U16539 (N_16539,N_15784,N_16053);
or U16540 (N_16540,N_15971,N_15871);
nand U16541 (N_16541,N_15664,N_15726);
nand U16542 (N_16542,N_16150,N_16175);
nor U16543 (N_16543,N_15863,N_15728);
nand U16544 (N_16544,N_15956,N_16073);
xor U16545 (N_16545,N_15928,N_15701);
nor U16546 (N_16546,N_16005,N_15837);
and U16547 (N_16547,N_15791,N_15893);
or U16548 (N_16548,N_16137,N_15610);
xnor U16549 (N_16549,N_15660,N_16021);
and U16550 (N_16550,N_15726,N_16185);
xnor U16551 (N_16551,N_15667,N_15829);
or U16552 (N_16552,N_15604,N_15866);
nor U16553 (N_16553,N_16065,N_15661);
nand U16554 (N_16554,N_15831,N_15925);
nor U16555 (N_16555,N_15995,N_15958);
nor U16556 (N_16556,N_15695,N_15910);
xor U16557 (N_16557,N_15728,N_15606);
and U16558 (N_16558,N_16127,N_16078);
or U16559 (N_16559,N_15781,N_15727);
and U16560 (N_16560,N_16117,N_15633);
or U16561 (N_16561,N_15855,N_15858);
and U16562 (N_16562,N_16018,N_15869);
or U16563 (N_16563,N_16188,N_15714);
nand U16564 (N_16564,N_15799,N_15931);
and U16565 (N_16565,N_15973,N_15996);
or U16566 (N_16566,N_15683,N_15734);
nor U16567 (N_16567,N_16165,N_16132);
nand U16568 (N_16568,N_16099,N_16058);
and U16569 (N_16569,N_15704,N_15745);
nor U16570 (N_16570,N_15631,N_15950);
or U16571 (N_16571,N_16139,N_15956);
nand U16572 (N_16572,N_15613,N_16170);
nand U16573 (N_16573,N_15620,N_15997);
or U16574 (N_16574,N_15990,N_15971);
nand U16575 (N_16575,N_15699,N_16179);
nand U16576 (N_16576,N_15869,N_15784);
xor U16577 (N_16577,N_15989,N_16016);
and U16578 (N_16578,N_15734,N_16150);
and U16579 (N_16579,N_15708,N_16081);
nor U16580 (N_16580,N_15887,N_16040);
xnor U16581 (N_16581,N_15914,N_15990);
and U16582 (N_16582,N_15915,N_15951);
nand U16583 (N_16583,N_15969,N_16154);
nand U16584 (N_16584,N_16087,N_15741);
or U16585 (N_16585,N_15947,N_16016);
nor U16586 (N_16586,N_15840,N_16124);
and U16587 (N_16587,N_15957,N_15617);
and U16588 (N_16588,N_15998,N_15731);
nand U16589 (N_16589,N_16148,N_15833);
or U16590 (N_16590,N_16024,N_15752);
nand U16591 (N_16591,N_15800,N_15915);
or U16592 (N_16592,N_15769,N_15997);
nor U16593 (N_16593,N_15737,N_15939);
xor U16594 (N_16594,N_15869,N_15873);
nand U16595 (N_16595,N_16149,N_15861);
nand U16596 (N_16596,N_16071,N_16197);
and U16597 (N_16597,N_15899,N_15916);
or U16598 (N_16598,N_15773,N_16023);
and U16599 (N_16599,N_15990,N_15839);
xor U16600 (N_16600,N_16108,N_15702);
nand U16601 (N_16601,N_16028,N_15940);
nand U16602 (N_16602,N_15785,N_16145);
and U16603 (N_16603,N_15956,N_16198);
or U16604 (N_16604,N_15927,N_15951);
or U16605 (N_16605,N_15731,N_15740);
and U16606 (N_16606,N_15900,N_16072);
xor U16607 (N_16607,N_15623,N_15660);
and U16608 (N_16608,N_15998,N_15855);
nor U16609 (N_16609,N_16154,N_16091);
nand U16610 (N_16610,N_15806,N_15924);
nor U16611 (N_16611,N_15930,N_15874);
or U16612 (N_16612,N_15608,N_15982);
and U16613 (N_16613,N_15871,N_16125);
xor U16614 (N_16614,N_15695,N_15620);
nand U16615 (N_16615,N_15779,N_16197);
nand U16616 (N_16616,N_16145,N_15751);
nand U16617 (N_16617,N_16068,N_15787);
or U16618 (N_16618,N_15703,N_15949);
or U16619 (N_16619,N_15813,N_15883);
nand U16620 (N_16620,N_16157,N_15721);
nor U16621 (N_16621,N_15761,N_15703);
and U16622 (N_16622,N_16002,N_15880);
xor U16623 (N_16623,N_15620,N_15771);
or U16624 (N_16624,N_15957,N_15821);
xnor U16625 (N_16625,N_15629,N_15870);
nor U16626 (N_16626,N_16070,N_15804);
nor U16627 (N_16627,N_16049,N_15847);
xnor U16628 (N_16628,N_16090,N_15836);
nand U16629 (N_16629,N_16001,N_16173);
nor U16630 (N_16630,N_15792,N_15633);
xor U16631 (N_16631,N_15967,N_15828);
xnor U16632 (N_16632,N_16006,N_15920);
and U16633 (N_16633,N_15718,N_15627);
and U16634 (N_16634,N_16041,N_15825);
xor U16635 (N_16635,N_15872,N_16022);
xor U16636 (N_16636,N_16019,N_16066);
and U16637 (N_16637,N_15723,N_16096);
nor U16638 (N_16638,N_15793,N_15904);
or U16639 (N_16639,N_15883,N_15893);
nand U16640 (N_16640,N_16109,N_15704);
xnor U16641 (N_16641,N_16105,N_16165);
or U16642 (N_16642,N_16151,N_16164);
and U16643 (N_16643,N_15641,N_15903);
and U16644 (N_16644,N_15615,N_15624);
xor U16645 (N_16645,N_16085,N_16119);
xnor U16646 (N_16646,N_15896,N_15651);
nor U16647 (N_16647,N_16058,N_15853);
and U16648 (N_16648,N_16163,N_15991);
and U16649 (N_16649,N_15695,N_15721);
nand U16650 (N_16650,N_16133,N_15823);
and U16651 (N_16651,N_16060,N_16067);
nand U16652 (N_16652,N_15950,N_15681);
nor U16653 (N_16653,N_16033,N_15755);
xor U16654 (N_16654,N_15727,N_16015);
or U16655 (N_16655,N_16143,N_16140);
nand U16656 (N_16656,N_16121,N_15947);
nor U16657 (N_16657,N_15601,N_16163);
nand U16658 (N_16658,N_16030,N_15615);
nand U16659 (N_16659,N_15656,N_15624);
xnor U16660 (N_16660,N_15657,N_15874);
nand U16661 (N_16661,N_15795,N_15807);
nor U16662 (N_16662,N_15618,N_16088);
or U16663 (N_16663,N_15822,N_15895);
or U16664 (N_16664,N_16093,N_15928);
nand U16665 (N_16665,N_15793,N_16102);
nor U16666 (N_16666,N_15885,N_16134);
xor U16667 (N_16667,N_16100,N_16097);
or U16668 (N_16668,N_16173,N_16069);
nand U16669 (N_16669,N_15674,N_15783);
or U16670 (N_16670,N_16118,N_15767);
or U16671 (N_16671,N_15818,N_16104);
or U16672 (N_16672,N_15639,N_15986);
xnor U16673 (N_16673,N_15849,N_15765);
and U16674 (N_16674,N_16081,N_16132);
and U16675 (N_16675,N_15760,N_16157);
or U16676 (N_16676,N_15934,N_16193);
nor U16677 (N_16677,N_16181,N_16021);
xor U16678 (N_16678,N_15920,N_15847);
nor U16679 (N_16679,N_15759,N_16144);
nand U16680 (N_16680,N_16157,N_15970);
or U16681 (N_16681,N_15972,N_15965);
or U16682 (N_16682,N_16157,N_15844);
and U16683 (N_16683,N_15876,N_15912);
or U16684 (N_16684,N_15925,N_16003);
nor U16685 (N_16685,N_15672,N_15967);
and U16686 (N_16686,N_15944,N_15919);
nand U16687 (N_16687,N_15721,N_15802);
nor U16688 (N_16688,N_15927,N_16132);
nor U16689 (N_16689,N_15671,N_16143);
and U16690 (N_16690,N_15656,N_15940);
or U16691 (N_16691,N_15901,N_16125);
and U16692 (N_16692,N_15843,N_15987);
xnor U16693 (N_16693,N_15947,N_15911);
and U16694 (N_16694,N_15786,N_16059);
nand U16695 (N_16695,N_15648,N_15968);
nand U16696 (N_16696,N_16198,N_16153);
and U16697 (N_16697,N_15822,N_15845);
and U16698 (N_16698,N_15941,N_16045);
nand U16699 (N_16699,N_15860,N_16087);
nor U16700 (N_16700,N_15826,N_15989);
or U16701 (N_16701,N_16061,N_15610);
nor U16702 (N_16702,N_15653,N_15668);
or U16703 (N_16703,N_15992,N_15646);
or U16704 (N_16704,N_15853,N_16040);
and U16705 (N_16705,N_15882,N_15712);
nor U16706 (N_16706,N_15647,N_15662);
and U16707 (N_16707,N_15704,N_16030);
nor U16708 (N_16708,N_15899,N_15610);
or U16709 (N_16709,N_16122,N_15869);
or U16710 (N_16710,N_15637,N_15658);
nand U16711 (N_16711,N_16032,N_15748);
nor U16712 (N_16712,N_15665,N_15766);
xor U16713 (N_16713,N_16028,N_15753);
nand U16714 (N_16714,N_15789,N_15942);
xnor U16715 (N_16715,N_15618,N_15984);
xor U16716 (N_16716,N_16176,N_15654);
nor U16717 (N_16717,N_16198,N_16122);
nor U16718 (N_16718,N_15907,N_15774);
and U16719 (N_16719,N_15692,N_15966);
or U16720 (N_16720,N_16173,N_15741);
nor U16721 (N_16721,N_15998,N_15784);
or U16722 (N_16722,N_15868,N_15846);
nand U16723 (N_16723,N_15967,N_15721);
and U16724 (N_16724,N_15832,N_15880);
nor U16725 (N_16725,N_16045,N_15821);
xor U16726 (N_16726,N_15868,N_15663);
or U16727 (N_16727,N_16027,N_15882);
nand U16728 (N_16728,N_15610,N_16010);
or U16729 (N_16729,N_16125,N_16193);
xor U16730 (N_16730,N_16056,N_16051);
or U16731 (N_16731,N_15662,N_16185);
or U16732 (N_16732,N_16155,N_15963);
and U16733 (N_16733,N_15888,N_16145);
or U16734 (N_16734,N_16015,N_16162);
nand U16735 (N_16735,N_15913,N_15735);
nor U16736 (N_16736,N_15722,N_15905);
xor U16737 (N_16737,N_16160,N_15676);
xnor U16738 (N_16738,N_15616,N_15791);
nand U16739 (N_16739,N_15746,N_15969);
xnor U16740 (N_16740,N_16130,N_15618);
and U16741 (N_16741,N_15917,N_16146);
nand U16742 (N_16742,N_15964,N_16053);
and U16743 (N_16743,N_15966,N_15789);
nor U16744 (N_16744,N_16197,N_15667);
xnor U16745 (N_16745,N_15825,N_15994);
nor U16746 (N_16746,N_16162,N_15981);
or U16747 (N_16747,N_15934,N_16102);
xor U16748 (N_16748,N_16057,N_15626);
xnor U16749 (N_16749,N_16002,N_15899);
nand U16750 (N_16750,N_15861,N_16107);
and U16751 (N_16751,N_15996,N_16012);
or U16752 (N_16752,N_15794,N_15772);
xor U16753 (N_16753,N_15719,N_15992);
nand U16754 (N_16754,N_16016,N_15697);
xor U16755 (N_16755,N_15824,N_15970);
or U16756 (N_16756,N_15787,N_15635);
nor U16757 (N_16757,N_16139,N_15845);
xor U16758 (N_16758,N_16080,N_15961);
nand U16759 (N_16759,N_15892,N_15653);
nor U16760 (N_16760,N_15835,N_16157);
nor U16761 (N_16761,N_15776,N_16053);
xnor U16762 (N_16762,N_15653,N_15794);
or U16763 (N_16763,N_16135,N_15877);
nand U16764 (N_16764,N_16103,N_15982);
nand U16765 (N_16765,N_15626,N_15947);
and U16766 (N_16766,N_15837,N_15726);
nor U16767 (N_16767,N_15698,N_15942);
nor U16768 (N_16768,N_16184,N_15923);
nor U16769 (N_16769,N_16031,N_15815);
and U16770 (N_16770,N_15979,N_15876);
and U16771 (N_16771,N_15772,N_15717);
nor U16772 (N_16772,N_16143,N_15724);
and U16773 (N_16773,N_16027,N_16132);
xor U16774 (N_16774,N_16085,N_15961);
nor U16775 (N_16775,N_15994,N_15614);
nor U16776 (N_16776,N_16193,N_15771);
nand U16777 (N_16777,N_15628,N_15903);
or U16778 (N_16778,N_15744,N_15917);
nand U16779 (N_16779,N_16089,N_15866);
or U16780 (N_16780,N_16178,N_15663);
and U16781 (N_16781,N_15801,N_15954);
or U16782 (N_16782,N_16197,N_16077);
xnor U16783 (N_16783,N_15931,N_16174);
and U16784 (N_16784,N_15710,N_15790);
nor U16785 (N_16785,N_16127,N_15967);
nor U16786 (N_16786,N_15608,N_15635);
or U16787 (N_16787,N_16040,N_15896);
and U16788 (N_16788,N_16024,N_16107);
or U16789 (N_16789,N_15815,N_15915);
or U16790 (N_16790,N_16053,N_15873);
xor U16791 (N_16791,N_15896,N_16036);
nand U16792 (N_16792,N_16007,N_16173);
xnor U16793 (N_16793,N_15946,N_16152);
nor U16794 (N_16794,N_16163,N_16181);
and U16795 (N_16795,N_15957,N_15614);
nor U16796 (N_16796,N_15816,N_15957);
xnor U16797 (N_16797,N_15811,N_16194);
and U16798 (N_16798,N_15873,N_15745);
nand U16799 (N_16799,N_15699,N_15931);
nand U16800 (N_16800,N_16638,N_16684);
xor U16801 (N_16801,N_16511,N_16489);
nor U16802 (N_16802,N_16367,N_16423);
xor U16803 (N_16803,N_16345,N_16709);
nand U16804 (N_16804,N_16412,N_16290);
nand U16805 (N_16805,N_16582,N_16749);
nand U16806 (N_16806,N_16569,N_16347);
nor U16807 (N_16807,N_16765,N_16581);
nand U16808 (N_16808,N_16401,N_16735);
and U16809 (N_16809,N_16524,N_16275);
nor U16810 (N_16810,N_16790,N_16535);
or U16811 (N_16811,N_16490,N_16289);
nand U16812 (N_16812,N_16518,N_16263);
nand U16813 (N_16813,N_16306,N_16388);
nand U16814 (N_16814,N_16291,N_16556);
and U16815 (N_16815,N_16646,N_16411);
nor U16816 (N_16816,N_16462,N_16369);
and U16817 (N_16817,N_16792,N_16598);
nor U16818 (N_16818,N_16757,N_16674);
and U16819 (N_16819,N_16705,N_16710);
xor U16820 (N_16820,N_16762,N_16526);
xor U16821 (N_16821,N_16766,N_16328);
and U16822 (N_16822,N_16285,N_16390);
and U16823 (N_16823,N_16726,N_16383);
nor U16824 (N_16824,N_16261,N_16316);
nor U16825 (N_16825,N_16441,N_16280);
xor U16826 (N_16826,N_16783,N_16795);
nand U16827 (N_16827,N_16601,N_16515);
or U16828 (N_16828,N_16586,N_16611);
or U16829 (N_16829,N_16459,N_16405);
xnor U16830 (N_16830,N_16561,N_16697);
xnor U16831 (N_16831,N_16558,N_16435);
nor U16832 (N_16832,N_16759,N_16568);
nand U16833 (N_16833,N_16440,N_16689);
xor U16834 (N_16834,N_16787,N_16623);
and U16835 (N_16835,N_16360,N_16476);
nand U16836 (N_16836,N_16782,N_16716);
nor U16837 (N_16837,N_16791,N_16225);
and U16838 (N_16838,N_16727,N_16610);
nand U16839 (N_16839,N_16607,N_16549);
and U16840 (N_16840,N_16382,N_16399);
nand U16841 (N_16841,N_16532,N_16536);
nor U16842 (N_16842,N_16723,N_16415);
xor U16843 (N_16843,N_16648,N_16510);
or U16844 (N_16844,N_16711,N_16438);
xnor U16845 (N_16845,N_16277,N_16577);
and U16846 (N_16846,N_16396,N_16756);
and U16847 (N_16847,N_16203,N_16721);
xor U16848 (N_16848,N_16690,N_16303);
or U16849 (N_16849,N_16769,N_16619);
or U16850 (N_16850,N_16310,N_16530);
nand U16851 (N_16851,N_16418,N_16338);
nor U16852 (N_16852,N_16429,N_16650);
nand U16853 (N_16853,N_16640,N_16724);
nor U16854 (N_16854,N_16617,N_16633);
and U16855 (N_16855,N_16269,N_16486);
nand U16856 (N_16856,N_16732,N_16230);
and U16857 (N_16857,N_16245,N_16737);
nor U16858 (N_16858,N_16753,N_16672);
nand U16859 (N_16859,N_16651,N_16589);
nor U16860 (N_16860,N_16470,N_16327);
and U16861 (N_16861,N_16293,N_16660);
nor U16862 (N_16862,N_16222,N_16478);
xnor U16863 (N_16863,N_16521,N_16579);
and U16864 (N_16864,N_16629,N_16381);
xor U16865 (N_16865,N_16520,N_16439);
nand U16866 (N_16866,N_16344,N_16428);
nand U16867 (N_16867,N_16608,N_16455);
nor U16868 (N_16868,N_16416,N_16797);
and U16869 (N_16869,N_16343,N_16449);
or U16870 (N_16870,N_16706,N_16599);
or U16871 (N_16871,N_16502,N_16529);
nor U16872 (N_16872,N_16323,N_16663);
and U16873 (N_16873,N_16352,N_16477);
xor U16874 (N_16874,N_16537,N_16249);
xor U16875 (N_16875,N_16346,N_16644);
or U16876 (N_16876,N_16278,N_16580);
nand U16877 (N_16877,N_16400,N_16202);
or U16878 (N_16878,N_16741,N_16223);
xnor U16879 (N_16879,N_16528,N_16761);
nand U16880 (N_16880,N_16484,N_16687);
or U16881 (N_16881,N_16567,N_16200);
nor U16882 (N_16882,N_16265,N_16417);
xnor U16883 (N_16883,N_16544,N_16313);
and U16884 (N_16884,N_16227,N_16754);
nor U16885 (N_16885,N_16666,N_16216);
nor U16886 (N_16886,N_16469,N_16768);
xor U16887 (N_16887,N_16512,N_16776);
or U16888 (N_16888,N_16519,N_16618);
and U16889 (N_16889,N_16395,N_16448);
and U16890 (N_16890,N_16686,N_16699);
nor U16891 (N_16891,N_16548,N_16321);
nor U16892 (N_16892,N_16314,N_16270);
nor U16893 (N_16893,N_16661,N_16593);
or U16894 (N_16894,N_16777,N_16466);
and U16895 (N_16895,N_16774,N_16793);
and U16896 (N_16896,N_16614,N_16335);
nor U16897 (N_16897,N_16786,N_16714);
and U16898 (N_16898,N_16295,N_16217);
or U16899 (N_16899,N_16479,N_16298);
or U16900 (N_16900,N_16665,N_16483);
nand U16901 (N_16901,N_16677,N_16755);
and U16902 (N_16902,N_16231,N_16342);
nand U16903 (N_16903,N_16679,N_16273);
xor U16904 (N_16904,N_16675,N_16377);
nand U16905 (N_16905,N_16523,N_16613);
nor U16906 (N_16906,N_16404,N_16540);
xnor U16907 (N_16907,N_16211,N_16514);
nor U16908 (N_16908,N_16264,N_16457);
nor U16909 (N_16909,N_16767,N_16334);
xnor U16910 (N_16910,N_16775,N_16372);
xor U16911 (N_16911,N_16788,N_16340);
nor U16912 (N_16912,N_16652,N_16364);
nor U16913 (N_16913,N_16332,N_16408);
nand U16914 (N_16914,N_16384,N_16320);
or U16915 (N_16915,N_16616,N_16373);
or U16916 (N_16916,N_16258,N_16595);
or U16917 (N_16917,N_16394,N_16212);
nand U16918 (N_16918,N_16432,N_16733);
nand U16919 (N_16919,N_16501,N_16325);
or U16920 (N_16920,N_16545,N_16664);
xor U16921 (N_16921,N_16257,N_16292);
xor U16922 (N_16922,N_16233,N_16503);
nor U16923 (N_16923,N_16253,N_16246);
nor U16924 (N_16924,N_16718,N_16739);
nand U16925 (N_16925,N_16734,N_16375);
or U16926 (N_16926,N_16682,N_16494);
or U16927 (N_16927,N_16240,N_16201);
or U16928 (N_16928,N_16659,N_16318);
and U16929 (N_16929,N_16557,N_16379);
nor U16930 (N_16930,N_16226,N_16385);
nand U16931 (N_16931,N_16221,N_16337);
xnor U16932 (N_16932,N_16588,N_16508);
or U16933 (N_16933,N_16256,N_16585);
or U16934 (N_16934,N_16683,N_16238);
xor U16935 (N_16935,N_16322,N_16612);
nor U16936 (N_16936,N_16630,N_16308);
nor U16937 (N_16937,N_16693,N_16299);
xor U16938 (N_16938,N_16229,N_16587);
xnor U16939 (N_16939,N_16274,N_16570);
xnor U16940 (N_16940,N_16239,N_16673);
or U16941 (N_16941,N_16622,N_16779);
or U16942 (N_16942,N_16413,N_16712);
and U16943 (N_16943,N_16228,N_16720);
nand U16944 (N_16944,N_16464,N_16444);
nand U16945 (N_16945,N_16252,N_16276);
or U16946 (N_16946,N_16563,N_16615);
nand U16947 (N_16947,N_16254,N_16424);
nand U16948 (N_16948,N_16604,N_16386);
or U16949 (N_16949,N_16669,N_16354);
nor U16950 (N_16950,N_16267,N_16309);
nand U16951 (N_16951,N_16546,N_16688);
xor U16952 (N_16952,N_16685,N_16205);
xnor U16953 (N_16953,N_16565,N_16368);
or U16954 (N_16954,N_16632,N_16625);
or U16955 (N_16955,N_16667,N_16780);
xor U16956 (N_16956,N_16363,N_16715);
nor U16957 (N_16957,N_16324,N_16410);
and U16958 (N_16958,N_16559,N_16255);
nor U16959 (N_16959,N_16358,N_16329);
and U16960 (N_16960,N_16407,N_16499);
nor U16961 (N_16961,N_16596,N_16642);
or U16962 (N_16962,N_16304,N_16422);
nor U16963 (N_16963,N_16771,N_16336);
nand U16964 (N_16964,N_16729,N_16763);
xor U16965 (N_16965,N_16764,N_16224);
nand U16966 (N_16966,N_16387,N_16402);
and U16967 (N_16967,N_16241,N_16606);
nand U16968 (N_16968,N_16218,N_16279);
or U16969 (N_16969,N_16398,N_16475);
and U16970 (N_16970,N_16305,N_16392);
xnor U16971 (N_16971,N_16431,N_16789);
nor U16972 (N_16972,N_16286,N_16208);
xor U16973 (N_16973,N_16592,N_16725);
nand U16974 (N_16974,N_16496,N_16708);
xor U16975 (N_16975,N_16206,N_16700);
nand U16976 (N_16976,N_16707,N_16695);
xnor U16977 (N_16977,N_16294,N_16473);
or U16978 (N_16978,N_16799,N_16434);
nor U16979 (N_16979,N_16717,N_16220);
nor U16980 (N_16980,N_16590,N_16566);
or U16981 (N_16981,N_16643,N_16597);
and U16982 (N_16982,N_16414,N_16636);
xnor U16983 (N_16983,N_16678,N_16751);
and U16984 (N_16984,N_16578,N_16728);
and U16985 (N_16985,N_16555,N_16425);
nand U16986 (N_16986,N_16624,N_16743);
xor U16987 (N_16987,N_16266,N_16430);
xor U16988 (N_16988,N_16272,N_16349);
nor U16989 (N_16989,N_16451,N_16676);
xnor U16990 (N_16990,N_16722,N_16333);
nand U16991 (N_16991,N_16785,N_16297);
and U16992 (N_16992,N_16366,N_16235);
or U16993 (N_16993,N_16282,N_16311);
and U16994 (N_16994,N_16738,N_16488);
nor U16995 (N_16995,N_16259,N_16692);
xor U16996 (N_16996,N_16406,N_16654);
and U16997 (N_16997,N_16271,N_16543);
or U16998 (N_16998,N_16210,N_16703);
xor U16999 (N_16999,N_16740,N_16621);
xor U17000 (N_17000,N_16359,N_16750);
nand U17001 (N_17001,N_16628,N_16620);
and U17002 (N_17002,N_16584,N_16420);
and U17003 (N_17003,N_16331,N_16542);
or U17004 (N_17004,N_16656,N_16748);
or U17005 (N_17005,N_16752,N_16248);
and U17006 (N_17006,N_16244,N_16436);
and U17007 (N_17007,N_16770,N_16350);
or U17008 (N_17008,N_16784,N_16452);
or U17009 (N_17009,N_16236,N_16232);
and U17010 (N_17010,N_16378,N_16798);
or U17011 (N_17011,N_16572,N_16641);
nand U17012 (N_17012,N_16370,N_16547);
or U17013 (N_17013,N_16433,N_16713);
or U17014 (N_17014,N_16554,N_16576);
and U17015 (N_17015,N_16517,N_16281);
xor U17016 (N_17016,N_16702,N_16627);
and U17017 (N_17017,N_16302,N_16247);
and U17018 (N_17018,N_16602,N_16376);
nand U17019 (N_17019,N_16355,N_16207);
nor U17020 (N_17020,N_16456,N_16639);
xnor U17021 (N_17021,N_16634,N_16560);
nand U17022 (N_17022,N_16453,N_16471);
or U17023 (N_17023,N_16296,N_16391);
or U17024 (N_17024,N_16730,N_16397);
nand U17025 (N_17025,N_16491,N_16482);
nand U17026 (N_17026,N_16746,N_16551);
and U17027 (N_17027,N_16487,N_16250);
nand U17028 (N_17028,N_16516,N_16330);
nor U17029 (N_17029,N_16507,N_16553);
xnor U17030 (N_17030,N_16284,N_16357);
or U17031 (N_17031,N_16758,N_16307);
nand U17032 (N_17032,N_16657,N_16583);
nand U17033 (N_17033,N_16301,N_16778);
or U17034 (N_17034,N_16742,N_16744);
or U17035 (N_17035,N_16450,N_16371);
nor U17036 (N_17036,N_16562,N_16326);
and U17037 (N_17037,N_16209,N_16319);
or U17038 (N_17038,N_16481,N_16704);
xnor U17039 (N_17039,N_16701,N_16609);
nand U17040 (N_17040,N_16681,N_16505);
or U17041 (N_17041,N_16214,N_16671);
nor U17042 (N_17042,N_16463,N_16437);
and U17043 (N_17043,N_16600,N_16362);
or U17044 (N_17044,N_16467,N_16513);
xor U17045 (N_17045,N_16389,N_16594);
nor U17046 (N_17046,N_16458,N_16541);
and U17047 (N_17047,N_16485,N_16351);
nor U17048 (N_17048,N_16747,N_16287);
or U17049 (N_17049,N_16772,N_16454);
xnor U17050 (N_17050,N_16461,N_16696);
nand U17051 (N_17051,N_16564,N_16234);
and U17052 (N_17052,N_16773,N_16760);
nor U17053 (N_17053,N_16575,N_16443);
nor U17054 (N_17054,N_16300,N_16315);
nand U17055 (N_17055,N_16492,N_16781);
and U17056 (N_17056,N_16504,N_16446);
or U17057 (N_17057,N_16403,N_16442);
nand U17058 (N_17058,N_16426,N_16506);
nand U17059 (N_17059,N_16731,N_16635);
nand U17060 (N_17060,N_16794,N_16670);
and U17061 (N_17061,N_16552,N_16288);
and U17062 (N_17062,N_16317,N_16447);
xnor U17063 (N_17063,N_16653,N_16525);
or U17064 (N_17064,N_16522,N_16348);
nand U17065 (N_17065,N_16237,N_16480);
nand U17066 (N_17066,N_16213,N_16380);
or U17067 (N_17067,N_16533,N_16419);
nand U17068 (N_17068,N_16465,N_16647);
and U17069 (N_17069,N_16495,N_16745);
and U17070 (N_17070,N_16312,N_16393);
nor U17071 (N_17071,N_16497,N_16460);
nand U17072 (N_17072,N_16468,N_16574);
or U17073 (N_17073,N_16571,N_16605);
nor U17074 (N_17074,N_16421,N_16531);
or U17075 (N_17075,N_16662,N_16409);
and U17076 (N_17076,N_16341,N_16365);
or U17077 (N_17077,N_16538,N_16215);
or U17078 (N_17078,N_16356,N_16474);
and U17079 (N_17079,N_16500,N_16353);
and U17080 (N_17080,N_16498,N_16268);
or U17081 (N_17081,N_16539,N_16680);
nand U17082 (N_17082,N_16534,N_16591);
nand U17083 (N_17083,N_16445,N_16796);
nand U17084 (N_17084,N_16719,N_16204);
nor U17085 (N_17085,N_16631,N_16527);
nor U17086 (N_17086,N_16736,N_16493);
or U17087 (N_17087,N_16573,N_16283);
nor U17088 (N_17088,N_16251,N_16645);
nor U17089 (N_17089,N_16658,N_16427);
nand U17090 (N_17090,N_16339,N_16374);
or U17091 (N_17091,N_16260,N_16698);
and U17092 (N_17092,N_16603,N_16262);
and U17093 (N_17093,N_16694,N_16655);
and U17094 (N_17094,N_16472,N_16691);
or U17095 (N_17095,N_16626,N_16509);
or U17096 (N_17096,N_16361,N_16550);
or U17097 (N_17097,N_16668,N_16637);
and U17098 (N_17098,N_16649,N_16242);
xnor U17099 (N_17099,N_16243,N_16219);
xor U17100 (N_17100,N_16788,N_16474);
xnor U17101 (N_17101,N_16758,N_16644);
and U17102 (N_17102,N_16626,N_16217);
xnor U17103 (N_17103,N_16768,N_16403);
or U17104 (N_17104,N_16710,N_16670);
and U17105 (N_17105,N_16581,N_16583);
and U17106 (N_17106,N_16604,N_16568);
or U17107 (N_17107,N_16207,N_16429);
nor U17108 (N_17108,N_16418,N_16391);
xor U17109 (N_17109,N_16479,N_16322);
or U17110 (N_17110,N_16419,N_16204);
nand U17111 (N_17111,N_16249,N_16513);
or U17112 (N_17112,N_16477,N_16731);
and U17113 (N_17113,N_16511,N_16534);
or U17114 (N_17114,N_16276,N_16655);
and U17115 (N_17115,N_16738,N_16330);
nor U17116 (N_17116,N_16735,N_16552);
xnor U17117 (N_17117,N_16291,N_16573);
nand U17118 (N_17118,N_16680,N_16319);
xnor U17119 (N_17119,N_16400,N_16574);
and U17120 (N_17120,N_16669,N_16504);
nor U17121 (N_17121,N_16467,N_16280);
nand U17122 (N_17122,N_16758,N_16650);
nor U17123 (N_17123,N_16359,N_16598);
or U17124 (N_17124,N_16342,N_16503);
xor U17125 (N_17125,N_16763,N_16400);
xnor U17126 (N_17126,N_16733,N_16583);
or U17127 (N_17127,N_16312,N_16293);
and U17128 (N_17128,N_16636,N_16580);
nor U17129 (N_17129,N_16544,N_16340);
nand U17130 (N_17130,N_16307,N_16224);
nor U17131 (N_17131,N_16624,N_16212);
or U17132 (N_17132,N_16657,N_16467);
nand U17133 (N_17133,N_16232,N_16608);
nor U17134 (N_17134,N_16676,N_16298);
nor U17135 (N_17135,N_16215,N_16592);
nand U17136 (N_17136,N_16648,N_16617);
nand U17137 (N_17137,N_16300,N_16280);
and U17138 (N_17138,N_16434,N_16649);
or U17139 (N_17139,N_16528,N_16329);
and U17140 (N_17140,N_16398,N_16759);
nand U17141 (N_17141,N_16713,N_16734);
nor U17142 (N_17142,N_16517,N_16665);
xnor U17143 (N_17143,N_16540,N_16231);
xor U17144 (N_17144,N_16694,N_16769);
nor U17145 (N_17145,N_16746,N_16652);
and U17146 (N_17146,N_16322,N_16628);
and U17147 (N_17147,N_16228,N_16750);
or U17148 (N_17148,N_16555,N_16742);
or U17149 (N_17149,N_16329,N_16620);
xor U17150 (N_17150,N_16299,N_16705);
or U17151 (N_17151,N_16755,N_16207);
nor U17152 (N_17152,N_16761,N_16269);
and U17153 (N_17153,N_16608,N_16523);
xor U17154 (N_17154,N_16520,N_16207);
xor U17155 (N_17155,N_16465,N_16702);
nand U17156 (N_17156,N_16414,N_16204);
nor U17157 (N_17157,N_16314,N_16498);
or U17158 (N_17158,N_16397,N_16748);
nor U17159 (N_17159,N_16205,N_16706);
or U17160 (N_17160,N_16572,N_16415);
xor U17161 (N_17161,N_16489,N_16522);
and U17162 (N_17162,N_16602,N_16231);
nor U17163 (N_17163,N_16219,N_16351);
and U17164 (N_17164,N_16286,N_16214);
nor U17165 (N_17165,N_16450,N_16705);
or U17166 (N_17166,N_16351,N_16560);
nor U17167 (N_17167,N_16540,N_16785);
xnor U17168 (N_17168,N_16477,N_16203);
xor U17169 (N_17169,N_16273,N_16473);
and U17170 (N_17170,N_16215,N_16569);
nand U17171 (N_17171,N_16391,N_16249);
or U17172 (N_17172,N_16368,N_16467);
nand U17173 (N_17173,N_16681,N_16736);
xor U17174 (N_17174,N_16257,N_16768);
xor U17175 (N_17175,N_16783,N_16754);
xor U17176 (N_17176,N_16590,N_16413);
nor U17177 (N_17177,N_16217,N_16581);
nand U17178 (N_17178,N_16298,N_16442);
xor U17179 (N_17179,N_16489,N_16779);
or U17180 (N_17180,N_16626,N_16748);
or U17181 (N_17181,N_16328,N_16312);
nand U17182 (N_17182,N_16530,N_16605);
nor U17183 (N_17183,N_16257,N_16497);
xnor U17184 (N_17184,N_16456,N_16541);
nor U17185 (N_17185,N_16442,N_16680);
nor U17186 (N_17186,N_16780,N_16732);
nor U17187 (N_17187,N_16378,N_16445);
nor U17188 (N_17188,N_16212,N_16728);
xor U17189 (N_17189,N_16612,N_16785);
xnor U17190 (N_17190,N_16793,N_16769);
or U17191 (N_17191,N_16385,N_16735);
nor U17192 (N_17192,N_16720,N_16543);
nor U17193 (N_17193,N_16407,N_16500);
or U17194 (N_17194,N_16751,N_16234);
nand U17195 (N_17195,N_16667,N_16377);
nor U17196 (N_17196,N_16662,N_16766);
and U17197 (N_17197,N_16352,N_16429);
and U17198 (N_17198,N_16485,N_16261);
nand U17199 (N_17199,N_16524,N_16449);
xor U17200 (N_17200,N_16379,N_16349);
xor U17201 (N_17201,N_16483,N_16628);
or U17202 (N_17202,N_16734,N_16702);
and U17203 (N_17203,N_16309,N_16306);
nor U17204 (N_17204,N_16256,N_16234);
nand U17205 (N_17205,N_16427,N_16581);
and U17206 (N_17206,N_16423,N_16647);
and U17207 (N_17207,N_16310,N_16728);
and U17208 (N_17208,N_16640,N_16565);
xor U17209 (N_17209,N_16534,N_16264);
and U17210 (N_17210,N_16418,N_16602);
nand U17211 (N_17211,N_16259,N_16659);
or U17212 (N_17212,N_16707,N_16756);
or U17213 (N_17213,N_16454,N_16750);
nor U17214 (N_17214,N_16541,N_16513);
or U17215 (N_17215,N_16538,N_16609);
nand U17216 (N_17216,N_16566,N_16341);
and U17217 (N_17217,N_16274,N_16366);
xnor U17218 (N_17218,N_16656,N_16302);
or U17219 (N_17219,N_16465,N_16267);
nor U17220 (N_17220,N_16674,N_16535);
or U17221 (N_17221,N_16654,N_16799);
and U17222 (N_17222,N_16560,N_16484);
and U17223 (N_17223,N_16404,N_16360);
nor U17224 (N_17224,N_16207,N_16319);
or U17225 (N_17225,N_16702,N_16420);
nand U17226 (N_17226,N_16625,N_16630);
xnor U17227 (N_17227,N_16383,N_16257);
nor U17228 (N_17228,N_16225,N_16416);
xor U17229 (N_17229,N_16546,N_16746);
or U17230 (N_17230,N_16444,N_16265);
xnor U17231 (N_17231,N_16700,N_16269);
or U17232 (N_17232,N_16348,N_16354);
xor U17233 (N_17233,N_16544,N_16716);
and U17234 (N_17234,N_16666,N_16775);
or U17235 (N_17235,N_16797,N_16353);
xor U17236 (N_17236,N_16708,N_16780);
nor U17237 (N_17237,N_16793,N_16751);
xor U17238 (N_17238,N_16522,N_16285);
nor U17239 (N_17239,N_16442,N_16643);
and U17240 (N_17240,N_16228,N_16717);
nand U17241 (N_17241,N_16392,N_16431);
and U17242 (N_17242,N_16421,N_16644);
nor U17243 (N_17243,N_16554,N_16590);
nor U17244 (N_17244,N_16302,N_16542);
or U17245 (N_17245,N_16692,N_16543);
or U17246 (N_17246,N_16339,N_16372);
nand U17247 (N_17247,N_16396,N_16786);
xnor U17248 (N_17248,N_16244,N_16542);
or U17249 (N_17249,N_16231,N_16317);
and U17250 (N_17250,N_16203,N_16639);
or U17251 (N_17251,N_16204,N_16571);
nor U17252 (N_17252,N_16687,N_16372);
nor U17253 (N_17253,N_16472,N_16345);
nor U17254 (N_17254,N_16653,N_16699);
nand U17255 (N_17255,N_16299,N_16420);
xor U17256 (N_17256,N_16393,N_16640);
or U17257 (N_17257,N_16593,N_16375);
nand U17258 (N_17258,N_16350,N_16693);
or U17259 (N_17259,N_16333,N_16380);
or U17260 (N_17260,N_16279,N_16697);
xor U17261 (N_17261,N_16261,N_16548);
nand U17262 (N_17262,N_16630,N_16709);
nor U17263 (N_17263,N_16622,N_16523);
nor U17264 (N_17264,N_16516,N_16607);
and U17265 (N_17265,N_16395,N_16238);
and U17266 (N_17266,N_16781,N_16210);
and U17267 (N_17267,N_16333,N_16309);
nor U17268 (N_17268,N_16286,N_16205);
xnor U17269 (N_17269,N_16297,N_16716);
nor U17270 (N_17270,N_16684,N_16581);
nand U17271 (N_17271,N_16361,N_16607);
and U17272 (N_17272,N_16338,N_16615);
and U17273 (N_17273,N_16548,N_16506);
nand U17274 (N_17274,N_16386,N_16312);
nor U17275 (N_17275,N_16614,N_16450);
xnor U17276 (N_17276,N_16463,N_16638);
nor U17277 (N_17277,N_16697,N_16499);
xnor U17278 (N_17278,N_16328,N_16347);
xnor U17279 (N_17279,N_16757,N_16368);
and U17280 (N_17280,N_16256,N_16491);
nor U17281 (N_17281,N_16223,N_16758);
nand U17282 (N_17282,N_16636,N_16696);
nand U17283 (N_17283,N_16750,N_16511);
nand U17284 (N_17284,N_16419,N_16714);
nand U17285 (N_17285,N_16582,N_16472);
xnor U17286 (N_17286,N_16755,N_16686);
and U17287 (N_17287,N_16707,N_16565);
nor U17288 (N_17288,N_16623,N_16403);
and U17289 (N_17289,N_16586,N_16257);
nand U17290 (N_17290,N_16482,N_16381);
xnor U17291 (N_17291,N_16646,N_16471);
nand U17292 (N_17292,N_16455,N_16406);
and U17293 (N_17293,N_16452,N_16730);
or U17294 (N_17294,N_16636,N_16638);
and U17295 (N_17295,N_16235,N_16477);
and U17296 (N_17296,N_16427,N_16380);
and U17297 (N_17297,N_16658,N_16501);
nand U17298 (N_17298,N_16339,N_16742);
and U17299 (N_17299,N_16558,N_16593);
nand U17300 (N_17300,N_16621,N_16732);
nor U17301 (N_17301,N_16700,N_16565);
nor U17302 (N_17302,N_16249,N_16750);
and U17303 (N_17303,N_16219,N_16687);
nor U17304 (N_17304,N_16583,N_16536);
or U17305 (N_17305,N_16779,N_16691);
nand U17306 (N_17306,N_16306,N_16568);
xnor U17307 (N_17307,N_16332,N_16458);
xnor U17308 (N_17308,N_16714,N_16473);
and U17309 (N_17309,N_16693,N_16342);
and U17310 (N_17310,N_16399,N_16675);
or U17311 (N_17311,N_16624,N_16723);
nor U17312 (N_17312,N_16672,N_16227);
nand U17313 (N_17313,N_16513,N_16255);
nand U17314 (N_17314,N_16568,N_16655);
or U17315 (N_17315,N_16279,N_16636);
and U17316 (N_17316,N_16607,N_16683);
or U17317 (N_17317,N_16579,N_16735);
and U17318 (N_17318,N_16632,N_16638);
and U17319 (N_17319,N_16685,N_16301);
or U17320 (N_17320,N_16267,N_16310);
nor U17321 (N_17321,N_16557,N_16645);
xnor U17322 (N_17322,N_16388,N_16447);
and U17323 (N_17323,N_16522,N_16527);
xnor U17324 (N_17324,N_16585,N_16744);
xor U17325 (N_17325,N_16582,N_16227);
nand U17326 (N_17326,N_16368,N_16647);
or U17327 (N_17327,N_16480,N_16678);
xor U17328 (N_17328,N_16283,N_16241);
or U17329 (N_17329,N_16267,N_16567);
nand U17330 (N_17330,N_16681,N_16511);
nor U17331 (N_17331,N_16526,N_16711);
or U17332 (N_17332,N_16799,N_16236);
or U17333 (N_17333,N_16274,N_16373);
nand U17334 (N_17334,N_16534,N_16442);
and U17335 (N_17335,N_16650,N_16546);
xor U17336 (N_17336,N_16639,N_16756);
xnor U17337 (N_17337,N_16516,N_16482);
or U17338 (N_17338,N_16559,N_16376);
nor U17339 (N_17339,N_16449,N_16420);
xor U17340 (N_17340,N_16744,N_16576);
nand U17341 (N_17341,N_16500,N_16421);
xor U17342 (N_17342,N_16727,N_16401);
nand U17343 (N_17343,N_16633,N_16703);
and U17344 (N_17344,N_16403,N_16585);
nor U17345 (N_17345,N_16406,N_16579);
and U17346 (N_17346,N_16392,N_16637);
xnor U17347 (N_17347,N_16644,N_16382);
nand U17348 (N_17348,N_16554,N_16765);
xnor U17349 (N_17349,N_16347,N_16436);
nor U17350 (N_17350,N_16464,N_16431);
or U17351 (N_17351,N_16224,N_16789);
xor U17352 (N_17352,N_16650,N_16527);
nor U17353 (N_17353,N_16556,N_16654);
xnor U17354 (N_17354,N_16797,N_16278);
nor U17355 (N_17355,N_16236,N_16538);
and U17356 (N_17356,N_16584,N_16553);
nand U17357 (N_17357,N_16562,N_16361);
nor U17358 (N_17358,N_16469,N_16748);
and U17359 (N_17359,N_16788,N_16451);
xor U17360 (N_17360,N_16248,N_16681);
and U17361 (N_17361,N_16226,N_16237);
or U17362 (N_17362,N_16377,N_16611);
nor U17363 (N_17363,N_16546,N_16413);
nor U17364 (N_17364,N_16640,N_16506);
and U17365 (N_17365,N_16741,N_16599);
nand U17366 (N_17366,N_16741,N_16352);
and U17367 (N_17367,N_16231,N_16213);
nand U17368 (N_17368,N_16369,N_16639);
nor U17369 (N_17369,N_16289,N_16493);
and U17370 (N_17370,N_16532,N_16366);
nand U17371 (N_17371,N_16517,N_16284);
nand U17372 (N_17372,N_16760,N_16527);
nand U17373 (N_17373,N_16235,N_16426);
or U17374 (N_17374,N_16364,N_16688);
nand U17375 (N_17375,N_16754,N_16647);
xnor U17376 (N_17376,N_16596,N_16517);
xor U17377 (N_17377,N_16769,N_16253);
nor U17378 (N_17378,N_16391,N_16265);
or U17379 (N_17379,N_16547,N_16407);
nand U17380 (N_17380,N_16788,N_16383);
xor U17381 (N_17381,N_16262,N_16553);
nor U17382 (N_17382,N_16723,N_16525);
nor U17383 (N_17383,N_16702,N_16240);
nor U17384 (N_17384,N_16212,N_16537);
nand U17385 (N_17385,N_16583,N_16462);
and U17386 (N_17386,N_16575,N_16623);
xnor U17387 (N_17387,N_16383,N_16282);
xor U17388 (N_17388,N_16326,N_16220);
nor U17389 (N_17389,N_16620,N_16422);
or U17390 (N_17390,N_16341,N_16493);
nand U17391 (N_17391,N_16300,N_16704);
nand U17392 (N_17392,N_16624,N_16333);
nand U17393 (N_17393,N_16281,N_16308);
and U17394 (N_17394,N_16398,N_16774);
or U17395 (N_17395,N_16241,N_16470);
or U17396 (N_17396,N_16550,N_16754);
or U17397 (N_17397,N_16749,N_16384);
or U17398 (N_17398,N_16470,N_16743);
or U17399 (N_17399,N_16360,N_16699);
nand U17400 (N_17400,N_17214,N_16898);
xnor U17401 (N_17401,N_17391,N_17284);
nand U17402 (N_17402,N_16987,N_17231);
xor U17403 (N_17403,N_17227,N_17126);
and U17404 (N_17404,N_17116,N_16849);
nand U17405 (N_17405,N_17183,N_16862);
or U17406 (N_17406,N_17179,N_16835);
and U17407 (N_17407,N_16954,N_17084);
and U17408 (N_17408,N_17259,N_17081);
nor U17409 (N_17409,N_16963,N_17119);
xnor U17410 (N_17410,N_17009,N_17289);
and U17411 (N_17411,N_17130,N_17364);
nand U17412 (N_17412,N_16989,N_16856);
nand U17413 (N_17413,N_17257,N_16929);
and U17414 (N_17414,N_17156,N_17033);
nand U17415 (N_17415,N_17275,N_17057);
and U17416 (N_17416,N_16827,N_17154);
xor U17417 (N_17417,N_16949,N_17170);
or U17418 (N_17418,N_17074,N_17345);
xnor U17419 (N_17419,N_16968,N_17120);
nand U17420 (N_17420,N_16994,N_16983);
or U17421 (N_17421,N_17038,N_17317);
and U17422 (N_17422,N_17213,N_17285);
nor U17423 (N_17423,N_16975,N_17082);
xnor U17424 (N_17424,N_16842,N_17316);
xor U17425 (N_17425,N_17110,N_17111);
nand U17426 (N_17426,N_16863,N_17080);
xnor U17427 (N_17427,N_16861,N_16804);
or U17428 (N_17428,N_17202,N_17191);
nor U17429 (N_17429,N_17143,N_17313);
and U17430 (N_17430,N_17205,N_17344);
xnor U17431 (N_17431,N_16906,N_17339);
nand U17432 (N_17432,N_17298,N_16834);
nand U17433 (N_17433,N_17189,N_16962);
nand U17434 (N_17434,N_17263,N_17046);
nand U17435 (N_17435,N_16915,N_17378);
nand U17436 (N_17436,N_16931,N_17019);
nand U17437 (N_17437,N_16953,N_16900);
nor U17438 (N_17438,N_17310,N_17078);
and U17439 (N_17439,N_17108,N_17000);
nor U17440 (N_17440,N_17247,N_17373);
or U17441 (N_17441,N_17328,N_17062);
and U17442 (N_17442,N_17255,N_16897);
xor U17443 (N_17443,N_17028,N_17077);
nand U17444 (N_17444,N_16896,N_16997);
and U17445 (N_17445,N_16951,N_17272);
and U17446 (N_17446,N_17321,N_16867);
xor U17447 (N_17447,N_16865,N_17195);
and U17448 (N_17448,N_16831,N_17161);
and U17449 (N_17449,N_16808,N_17278);
nand U17450 (N_17450,N_16993,N_16868);
or U17451 (N_17451,N_17357,N_16883);
nor U17452 (N_17452,N_17358,N_16969);
nor U17453 (N_17453,N_17058,N_16944);
nor U17454 (N_17454,N_17102,N_17204);
xnor U17455 (N_17455,N_16870,N_17260);
nor U17456 (N_17456,N_17301,N_17350);
or U17457 (N_17457,N_17376,N_17144);
and U17458 (N_17458,N_17300,N_17147);
nand U17459 (N_17459,N_17109,N_17017);
nor U17460 (N_17460,N_17209,N_16817);
nand U17461 (N_17461,N_17113,N_17211);
xnor U17462 (N_17462,N_17095,N_17125);
nor U17463 (N_17463,N_17290,N_16942);
nand U17464 (N_17464,N_16888,N_17016);
nor U17465 (N_17465,N_16967,N_16913);
and U17466 (N_17466,N_17224,N_16828);
nor U17467 (N_17467,N_17223,N_16947);
or U17468 (N_17468,N_17036,N_17248);
and U17469 (N_17469,N_17393,N_17256);
xor U17470 (N_17470,N_17387,N_16922);
nand U17471 (N_17471,N_17286,N_17150);
nand U17472 (N_17472,N_17309,N_17221);
and U17473 (N_17473,N_16902,N_17096);
nand U17474 (N_17474,N_17269,N_17382);
nand U17475 (N_17475,N_16977,N_17279);
and U17476 (N_17476,N_16806,N_17306);
or U17477 (N_17477,N_16818,N_17349);
or U17478 (N_17478,N_17106,N_16925);
or U17479 (N_17479,N_17145,N_17035);
xnor U17480 (N_17480,N_17199,N_16832);
nor U17481 (N_17481,N_17266,N_17359);
and U17482 (N_17482,N_17115,N_16823);
nor U17483 (N_17483,N_17105,N_17097);
or U17484 (N_17484,N_17064,N_17340);
and U17485 (N_17485,N_17308,N_16878);
or U17486 (N_17486,N_17388,N_17005);
and U17487 (N_17487,N_17249,N_17234);
or U17488 (N_17488,N_17068,N_17383);
nand U17489 (N_17489,N_16946,N_17222);
xnor U17490 (N_17490,N_17370,N_17245);
or U17491 (N_17491,N_16932,N_17201);
nand U17492 (N_17492,N_16958,N_17341);
xnor U17493 (N_17493,N_16839,N_17198);
xnor U17494 (N_17494,N_16923,N_17274);
or U17495 (N_17495,N_17335,N_16986);
and U17496 (N_17496,N_16860,N_17098);
or U17497 (N_17497,N_17165,N_17325);
xnor U17498 (N_17498,N_17287,N_16847);
or U17499 (N_17499,N_17217,N_17203);
and U17500 (N_17500,N_17187,N_17003);
and U17501 (N_17501,N_16805,N_17128);
or U17502 (N_17502,N_16801,N_17024);
and U17503 (N_17503,N_16838,N_16982);
xor U17504 (N_17504,N_16965,N_17190);
nor U17505 (N_17505,N_17398,N_17085);
nor U17506 (N_17506,N_17180,N_16879);
and U17507 (N_17507,N_17226,N_17394);
xor U17508 (N_17508,N_16841,N_17069);
or U17509 (N_17509,N_16943,N_17092);
xor U17510 (N_17510,N_17174,N_17244);
and U17511 (N_17511,N_17153,N_17208);
or U17512 (N_17512,N_17010,N_17379);
nand U17513 (N_17513,N_17242,N_16840);
or U17514 (N_17514,N_17021,N_17050);
xnor U17515 (N_17515,N_16984,N_16972);
nor U17516 (N_17516,N_16885,N_17206);
nor U17517 (N_17517,N_17250,N_17112);
nor U17518 (N_17518,N_17377,N_16966);
nor U17519 (N_17519,N_17066,N_17013);
xor U17520 (N_17520,N_17384,N_16903);
xor U17521 (N_17521,N_16973,N_16895);
nor U17522 (N_17522,N_16974,N_16936);
nand U17523 (N_17523,N_17194,N_16855);
nor U17524 (N_17524,N_16899,N_17372);
nand U17525 (N_17525,N_17163,N_17235);
or U17526 (N_17526,N_17338,N_16988);
nor U17527 (N_17527,N_16876,N_17129);
or U17528 (N_17528,N_17175,N_17396);
or U17529 (N_17529,N_17167,N_17014);
nor U17530 (N_17530,N_17314,N_17246);
nand U17531 (N_17531,N_17207,N_16803);
and U17532 (N_17532,N_16980,N_17271);
nor U17533 (N_17533,N_17363,N_17219);
nand U17534 (N_17534,N_17307,N_17299);
or U17535 (N_17535,N_17336,N_17261);
nor U17536 (N_17536,N_17353,N_17186);
nor U17537 (N_17537,N_16926,N_17166);
xnor U17538 (N_17538,N_17347,N_17216);
xnor U17539 (N_17539,N_17399,N_16952);
nand U17540 (N_17540,N_17090,N_16955);
nand U17541 (N_17541,N_16887,N_17210);
nor U17542 (N_17542,N_17149,N_17331);
nor U17543 (N_17543,N_17374,N_17103);
and U17544 (N_17544,N_17138,N_17040);
nor U17545 (N_17545,N_17196,N_16815);
and U17546 (N_17546,N_17160,N_17200);
nand U17547 (N_17547,N_16881,N_17100);
nor U17548 (N_17548,N_17146,N_16985);
and U17549 (N_17549,N_17232,N_16819);
nand U17550 (N_17550,N_16802,N_17293);
nor U17551 (N_17551,N_17094,N_17101);
or U17552 (N_17552,N_17368,N_17132);
and U17553 (N_17553,N_17323,N_16825);
nand U17554 (N_17554,N_17240,N_17041);
and U17555 (N_17555,N_17029,N_17291);
xor U17556 (N_17556,N_17079,N_16864);
or U17557 (N_17557,N_16837,N_16848);
or U17558 (N_17558,N_16882,N_17356);
and U17559 (N_17559,N_16941,N_17243);
xnor U17560 (N_17560,N_17073,N_17320);
nand U17561 (N_17561,N_16908,N_17133);
xor U17562 (N_17562,N_16919,N_17297);
nand U17563 (N_17563,N_17333,N_17020);
or U17564 (N_17564,N_17011,N_16914);
nor U17565 (N_17565,N_16886,N_16933);
nand U17566 (N_17566,N_16905,N_17239);
or U17567 (N_17567,N_17241,N_16981);
nor U17568 (N_17568,N_16996,N_17342);
or U17569 (N_17569,N_17076,N_17366);
and U17570 (N_17570,N_17311,N_17107);
or U17571 (N_17571,N_17367,N_17329);
xnor U17572 (N_17572,N_16976,N_16927);
nand U17573 (N_17573,N_16871,N_17008);
or U17574 (N_17574,N_17159,N_17052);
or U17575 (N_17575,N_16800,N_17151);
or U17576 (N_17576,N_16957,N_16911);
nor U17577 (N_17577,N_17193,N_17047);
and U17578 (N_17578,N_17185,N_16811);
and U17579 (N_17579,N_17343,N_17254);
nor U17580 (N_17580,N_16836,N_17181);
nand U17581 (N_17581,N_16894,N_16807);
or U17582 (N_17582,N_17086,N_17141);
nand U17583 (N_17583,N_17324,N_17381);
nand U17584 (N_17584,N_17385,N_17093);
nand U17585 (N_17585,N_17075,N_16934);
and U17586 (N_17586,N_17071,N_17006);
nand U17587 (N_17587,N_16833,N_16961);
xor U17588 (N_17588,N_17124,N_17139);
nor U17589 (N_17589,N_17360,N_16809);
xor U17590 (N_17590,N_17032,N_17001);
nor U17591 (N_17591,N_16964,N_17295);
and U17592 (N_17592,N_16938,N_16990);
xor U17593 (N_17593,N_16884,N_17045);
and U17594 (N_17594,N_17135,N_17276);
nor U17595 (N_17595,N_16916,N_16872);
or U17596 (N_17596,N_17089,N_17034);
or U17597 (N_17597,N_17192,N_16813);
nand U17598 (N_17598,N_17060,N_17212);
xor U17599 (N_17599,N_17330,N_16901);
and U17600 (N_17600,N_17365,N_17389);
xor U17601 (N_17601,N_17178,N_17055);
nor U17602 (N_17602,N_17039,N_17118);
nor U17603 (N_17603,N_17091,N_17164);
or U17604 (N_17604,N_16816,N_17351);
nor U17605 (N_17605,N_17137,N_16866);
and U17606 (N_17606,N_17072,N_17397);
xnor U17607 (N_17607,N_17121,N_17022);
xor U17608 (N_17608,N_17114,N_17294);
nand U17609 (N_17609,N_17265,N_17251);
nand U17610 (N_17610,N_17305,N_16810);
or U17611 (N_17611,N_16970,N_17122);
xor U17612 (N_17612,N_16851,N_17004);
xor U17613 (N_17613,N_16812,N_16814);
and U17614 (N_17614,N_17012,N_17348);
or U17615 (N_17615,N_17304,N_17168);
or U17616 (N_17616,N_17173,N_17334);
nor U17617 (N_17617,N_17322,N_17070);
and U17618 (N_17618,N_17127,N_16852);
xnor U17619 (N_17619,N_17140,N_17268);
or U17620 (N_17620,N_17326,N_16874);
or U17621 (N_17621,N_17197,N_17319);
and U17622 (N_17622,N_17162,N_16880);
nor U17623 (N_17623,N_17302,N_17327);
nand U17624 (N_17624,N_16889,N_17155);
xnor U17625 (N_17625,N_17283,N_17352);
or U17626 (N_17626,N_16910,N_16930);
or U17627 (N_17627,N_17264,N_17172);
nor U17628 (N_17628,N_17280,N_17061);
nand U17629 (N_17629,N_17152,N_17273);
or U17630 (N_17630,N_17053,N_17315);
nor U17631 (N_17631,N_16999,N_17288);
and U17632 (N_17632,N_16853,N_16950);
nand U17633 (N_17633,N_17371,N_17023);
nand U17634 (N_17634,N_16912,N_16830);
or U17635 (N_17635,N_16948,N_16909);
nand U17636 (N_17636,N_17395,N_17230);
xnor U17637 (N_17637,N_16939,N_17031);
nand U17638 (N_17638,N_17215,N_17088);
or U17639 (N_17639,N_16845,N_17346);
xor U17640 (N_17640,N_16821,N_16890);
nor U17641 (N_17641,N_17218,N_16844);
nor U17642 (N_17642,N_17281,N_17015);
xnor U17643 (N_17643,N_17332,N_16945);
and U17644 (N_17644,N_17148,N_17369);
nand U17645 (N_17645,N_17182,N_16904);
and U17646 (N_17646,N_17237,N_16921);
or U17647 (N_17647,N_17043,N_16956);
nand U17648 (N_17648,N_17312,N_16826);
nor U17649 (N_17649,N_17030,N_17253);
nor U17650 (N_17650,N_16992,N_17123);
or U17651 (N_17651,N_17177,N_16858);
nor U17652 (N_17652,N_17056,N_17362);
xnor U17653 (N_17653,N_17270,N_16893);
nor U17654 (N_17654,N_17262,N_17354);
nand U17655 (N_17655,N_16907,N_16940);
nor U17656 (N_17656,N_16846,N_17042);
and U17657 (N_17657,N_17049,N_17142);
or U17658 (N_17658,N_16820,N_17220);
and U17659 (N_17659,N_17018,N_17157);
nor U17660 (N_17660,N_16917,N_17277);
nor U17661 (N_17661,N_16991,N_16995);
nor U17662 (N_17662,N_17104,N_17303);
or U17663 (N_17663,N_17318,N_17296);
xnor U17664 (N_17664,N_17238,N_17065);
or U17665 (N_17665,N_16857,N_17252);
nand U17666 (N_17666,N_17236,N_17083);
or U17667 (N_17667,N_16998,N_17025);
and U17668 (N_17668,N_16854,N_17392);
xnor U17669 (N_17669,N_17267,N_16822);
and U17670 (N_17670,N_17099,N_17158);
xnor U17671 (N_17671,N_17228,N_17171);
xnor U17672 (N_17672,N_16935,N_17337);
and U17673 (N_17673,N_17051,N_17059);
nand U17674 (N_17674,N_16869,N_17225);
or U17675 (N_17675,N_17136,N_17169);
nor U17676 (N_17676,N_16924,N_17390);
nand U17677 (N_17677,N_16877,N_17375);
and U17678 (N_17678,N_17037,N_17048);
nand U17679 (N_17679,N_17063,N_16937);
and U17680 (N_17680,N_16920,N_17027);
nor U17681 (N_17681,N_16978,N_17380);
nand U17682 (N_17682,N_17176,N_16875);
xor U17683 (N_17683,N_17258,N_17131);
nor U17684 (N_17684,N_17282,N_17386);
and U17685 (N_17685,N_17134,N_17355);
xor U17686 (N_17686,N_17054,N_16979);
xnor U17687 (N_17687,N_17361,N_16824);
or U17688 (N_17688,N_17233,N_16959);
xor U17689 (N_17689,N_17184,N_16918);
nand U17690 (N_17690,N_16850,N_17007);
nor U17691 (N_17691,N_16971,N_16928);
or U17692 (N_17692,N_17087,N_16891);
nor U17693 (N_17693,N_16829,N_17229);
nand U17694 (N_17694,N_17292,N_16892);
xnor U17695 (N_17695,N_16843,N_17067);
and U17696 (N_17696,N_16960,N_16873);
nand U17697 (N_17697,N_17002,N_16859);
nor U17698 (N_17698,N_17044,N_17117);
nor U17699 (N_17699,N_17026,N_17188);
nand U17700 (N_17700,N_17172,N_16846);
nand U17701 (N_17701,N_17337,N_17161);
nand U17702 (N_17702,N_16976,N_17007);
nand U17703 (N_17703,N_17080,N_17304);
nor U17704 (N_17704,N_16921,N_17129);
and U17705 (N_17705,N_17250,N_17371);
nand U17706 (N_17706,N_17297,N_16977);
and U17707 (N_17707,N_16859,N_17257);
and U17708 (N_17708,N_16961,N_17187);
or U17709 (N_17709,N_16840,N_17195);
or U17710 (N_17710,N_17158,N_16862);
nor U17711 (N_17711,N_17348,N_16901);
and U17712 (N_17712,N_16906,N_16890);
or U17713 (N_17713,N_17149,N_16880);
or U17714 (N_17714,N_17234,N_16940);
xor U17715 (N_17715,N_16950,N_16825);
or U17716 (N_17716,N_16803,N_17099);
or U17717 (N_17717,N_17041,N_16838);
nor U17718 (N_17718,N_17194,N_17367);
xor U17719 (N_17719,N_16967,N_16850);
nor U17720 (N_17720,N_17196,N_16853);
nand U17721 (N_17721,N_17248,N_16804);
nor U17722 (N_17722,N_17026,N_17176);
xnor U17723 (N_17723,N_16988,N_17211);
and U17724 (N_17724,N_17238,N_17194);
and U17725 (N_17725,N_17047,N_17397);
xor U17726 (N_17726,N_16990,N_16907);
or U17727 (N_17727,N_16882,N_17257);
xnor U17728 (N_17728,N_17117,N_17243);
nand U17729 (N_17729,N_16836,N_17119);
xnor U17730 (N_17730,N_16911,N_17383);
or U17731 (N_17731,N_16890,N_17395);
nand U17732 (N_17732,N_16819,N_17213);
xor U17733 (N_17733,N_16818,N_16937);
and U17734 (N_17734,N_16959,N_17155);
nand U17735 (N_17735,N_17158,N_17226);
nand U17736 (N_17736,N_17370,N_17338);
and U17737 (N_17737,N_17153,N_16888);
and U17738 (N_17738,N_17030,N_17002);
xnor U17739 (N_17739,N_17362,N_16858);
nor U17740 (N_17740,N_17244,N_16923);
and U17741 (N_17741,N_17046,N_17049);
xnor U17742 (N_17742,N_17300,N_17237);
and U17743 (N_17743,N_17187,N_17015);
or U17744 (N_17744,N_17030,N_17026);
nor U17745 (N_17745,N_17257,N_16828);
or U17746 (N_17746,N_17251,N_16869);
and U17747 (N_17747,N_17237,N_16952);
and U17748 (N_17748,N_17147,N_17317);
or U17749 (N_17749,N_16854,N_17230);
and U17750 (N_17750,N_17244,N_17092);
xnor U17751 (N_17751,N_17089,N_16813);
and U17752 (N_17752,N_17161,N_16931);
xnor U17753 (N_17753,N_17382,N_16853);
nor U17754 (N_17754,N_17101,N_17184);
or U17755 (N_17755,N_16845,N_17281);
xnor U17756 (N_17756,N_17242,N_17132);
nor U17757 (N_17757,N_17302,N_16927);
or U17758 (N_17758,N_17344,N_16862);
nor U17759 (N_17759,N_17054,N_17196);
or U17760 (N_17760,N_16919,N_17104);
or U17761 (N_17761,N_17086,N_17185);
or U17762 (N_17762,N_17379,N_17117);
xor U17763 (N_17763,N_17080,N_16841);
or U17764 (N_17764,N_17297,N_17391);
xnor U17765 (N_17765,N_16887,N_17061);
or U17766 (N_17766,N_16978,N_16965);
and U17767 (N_17767,N_17232,N_17055);
nand U17768 (N_17768,N_16857,N_16979);
xnor U17769 (N_17769,N_16876,N_17067);
xnor U17770 (N_17770,N_17368,N_16940);
nand U17771 (N_17771,N_16996,N_17287);
xnor U17772 (N_17772,N_17221,N_17338);
nor U17773 (N_17773,N_17093,N_16935);
nor U17774 (N_17774,N_16975,N_16996);
nor U17775 (N_17775,N_16878,N_17203);
nor U17776 (N_17776,N_17014,N_17016);
or U17777 (N_17777,N_17081,N_17314);
and U17778 (N_17778,N_16991,N_16910);
and U17779 (N_17779,N_17257,N_17046);
xnor U17780 (N_17780,N_17020,N_17058);
nor U17781 (N_17781,N_17241,N_16906);
and U17782 (N_17782,N_17362,N_16885);
or U17783 (N_17783,N_17205,N_17372);
nor U17784 (N_17784,N_17390,N_17397);
xor U17785 (N_17785,N_17013,N_17156);
and U17786 (N_17786,N_17216,N_16823);
nor U17787 (N_17787,N_16845,N_17355);
nand U17788 (N_17788,N_16988,N_17062);
nand U17789 (N_17789,N_16938,N_16837);
and U17790 (N_17790,N_17252,N_16976);
xnor U17791 (N_17791,N_17249,N_16942);
nand U17792 (N_17792,N_17036,N_16818);
nand U17793 (N_17793,N_17394,N_17382);
nor U17794 (N_17794,N_16817,N_17045);
or U17795 (N_17795,N_17266,N_17219);
nor U17796 (N_17796,N_16803,N_17351);
and U17797 (N_17797,N_16999,N_17013);
nand U17798 (N_17798,N_16869,N_17302);
xnor U17799 (N_17799,N_17254,N_17076);
and U17800 (N_17800,N_17303,N_16993);
nor U17801 (N_17801,N_17391,N_17240);
nand U17802 (N_17802,N_17140,N_17252);
nor U17803 (N_17803,N_17204,N_16807);
and U17804 (N_17804,N_17169,N_16994);
xor U17805 (N_17805,N_17191,N_17091);
or U17806 (N_17806,N_17357,N_17035);
nand U17807 (N_17807,N_17093,N_16857);
nand U17808 (N_17808,N_17254,N_17198);
nor U17809 (N_17809,N_17089,N_17139);
xor U17810 (N_17810,N_17389,N_17223);
nor U17811 (N_17811,N_17196,N_17101);
nand U17812 (N_17812,N_17123,N_17014);
or U17813 (N_17813,N_17072,N_16863);
xor U17814 (N_17814,N_17206,N_17384);
xor U17815 (N_17815,N_17282,N_17325);
nand U17816 (N_17816,N_16952,N_16884);
and U17817 (N_17817,N_17308,N_17244);
or U17818 (N_17818,N_17284,N_17366);
and U17819 (N_17819,N_17158,N_17007);
nor U17820 (N_17820,N_16918,N_17349);
or U17821 (N_17821,N_16893,N_17282);
xor U17822 (N_17822,N_16838,N_16954);
xor U17823 (N_17823,N_17301,N_16959);
or U17824 (N_17824,N_16921,N_17226);
nand U17825 (N_17825,N_17301,N_17123);
nor U17826 (N_17826,N_16943,N_16863);
nor U17827 (N_17827,N_17248,N_16890);
nand U17828 (N_17828,N_17158,N_17271);
nand U17829 (N_17829,N_16925,N_16823);
and U17830 (N_17830,N_16963,N_17267);
and U17831 (N_17831,N_17279,N_17126);
or U17832 (N_17832,N_17088,N_17051);
xor U17833 (N_17833,N_16806,N_17112);
and U17834 (N_17834,N_17238,N_17394);
xnor U17835 (N_17835,N_17083,N_16818);
xnor U17836 (N_17836,N_17012,N_17327);
nor U17837 (N_17837,N_17238,N_17339);
xor U17838 (N_17838,N_17022,N_17303);
and U17839 (N_17839,N_17292,N_17157);
nor U17840 (N_17840,N_17358,N_16865);
or U17841 (N_17841,N_17009,N_17293);
nor U17842 (N_17842,N_17032,N_17249);
or U17843 (N_17843,N_16914,N_16886);
nor U17844 (N_17844,N_17276,N_17102);
and U17845 (N_17845,N_17385,N_16817);
nand U17846 (N_17846,N_17315,N_17012);
nand U17847 (N_17847,N_17239,N_16878);
or U17848 (N_17848,N_16817,N_16843);
nand U17849 (N_17849,N_17369,N_17008);
nor U17850 (N_17850,N_16850,N_16854);
and U17851 (N_17851,N_17200,N_17084);
and U17852 (N_17852,N_17006,N_17240);
and U17853 (N_17853,N_17330,N_17009);
xnor U17854 (N_17854,N_17160,N_17247);
nor U17855 (N_17855,N_17148,N_16899);
xnor U17856 (N_17856,N_16914,N_16907);
nor U17857 (N_17857,N_16916,N_16846);
xor U17858 (N_17858,N_17108,N_16852);
xnor U17859 (N_17859,N_17158,N_17035);
nand U17860 (N_17860,N_17041,N_16997);
or U17861 (N_17861,N_17361,N_16908);
nor U17862 (N_17862,N_16817,N_17364);
nor U17863 (N_17863,N_16955,N_16833);
and U17864 (N_17864,N_17097,N_17391);
and U17865 (N_17865,N_16919,N_17033);
xnor U17866 (N_17866,N_16805,N_17229);
nor U17867 (N_17867,N_17089,N_17379);
or U17868 (N_17868,N_17158,N_17133);
and U17869 (N_17869,N_17064,N_16926);
and U17870 (N_17870,N_16996,N_16941);
and U17871 (N_17871,N_17161,N_17151);
nand U17872 (N_17872,N_17234,N_17326);
and U17873 (N_17873,N_16828,N_17326);
and U17874 (N_17874,N_16822,N_17234);
xor U17875 (N_17875,N_16840,N_16950);
nand U17876 (N_17876,N_17278,N_16801);
and U17877 (N_17877,N_17394,N_17157);
or U17878 (N_17878,N_17188,N_17143);
or U17879 (N_17879,N_17044,N_16967);
and U17880 (N_17880,N_17055,N_17057);
nand U17881 (N_17881,N_17311,N_16872);
and U17882 (N_17882,N_17005,N_17214);
nand U17883 (N_17883,N_16900,N_17250);
and U17884 (N_17884,N_16810,N_17157);
or U17885 (N_17885,N_17120,N_16924);
xnor U17886 (N_17886,N_17274,N_17255);
and U17887 (N_17887,N_17070,N_16966);
xnor U17888 (N_17888,N_16998,N_17382);
nand U17889 (N_17889,N_16974,N_16935);
nor U17890 (N_17890,N_17370,N_16872);
or U17891 (N_17891,N_16947,N_17341);
nor U17892 (N_17892,N_17393,N_17126);
or U17893 (N_17893,N_17376,N_17389);
nand U17894 (N_17894,N_16941,N_17291);
and U17895 (N_17895,N_17019,N_17130);
and U17896 (N_17896,N_17016,N_16882);
and U17897 (N_17897,N_17288,N_17271);
nor U17898 (N_17898,N_17070,N_17352);
and U17899 (N_17899,N_17274,N_16821);
nand U17900 (N_17900,N_16947,N_17204);
and U17901 (N_17901,N_16916,N_16855);
nor U17902 (N_17902,N_16909,N_17080);
xnor U17903 (N_17903,N_17159,N_17146);
and U17904 (N_17904,N_17217,N_17040);
or U17905 (N_17905,N_16825,N_17046);
and U17906 (N_17906,N_17090,N_16888);
or U17907 (N_17907,N_16934,N_17225);
or U17908 (N_17908,N_17297,N_16999);
and U17909 (N_17909,N_17213,N_16907);
xor U17910 (N_17910,N_17225,N_17234);
nand U17911 (N_17911,N_16912,N_16832);
xnor U17912 (N_17912,N_17130,N_17162);
nand U17913 (N_17913,N_16840,N_17262);
or U17914 (N_17914,N_16869,N_17220);
nand U17915 (N_17915,N_16884,N_16983);
or U17916 (N_17916,N_17253,N_16895);
nand U17917 (N_17917,N_17020,N_16839);
or U17918 (N_17918,N_17357,N_17292);
and U17919 (N_17919,N_17058,N_16827);
nand U17920 (N_17920,N_16895,N_16825);
or U17921 (N_17921,N_16931,N_16982);
nand U17922 (N_17922,N_17075,N_16805);
nand U17923 (N_17923,N_17386,N_17184);
nand U17924 (N_17924,N_17290,N_17256);
nand U17925 (N_17925,N_16832,N_17010);
nand U17926 (N_17926,N_16974,N_17373);
or U17927 (N_17927,N_17356,N_16852);
nor U17928 (N_17928,N_17353,N_17140);
xnor U17929 (N_17929,N_17088,N_17059);
or U17930 (N_17930,N_17192,N_16978);
nor U17931 (N_17931,N_17179,N_17012);
xnor U17932 (N_17932,N_17348,N_16834);
or U17933 (N_17933,N_16934,N_17010);
and U17934 (N_17934,N_17129,N_17347);
or U17935 (N_17935,N_17353,N_17197);
or U17936 (N_17936,N_17025,N_17038);
xnor U17937 (N_17937,N_16816,N_16831);
and U17938 (N_17938,N_16894,N_17372);
xnor U17939 (N_17939,N_17292,N_16882);
xnor U17940 (N_17940,N_17180,N_17362);
nand U17941 (N_17941,N_16934,N_17355);
xor U17942 (N_17942,N_16857,N_17270);
nor U17943 (N_17943,N_17311,N_16893);
nor U17944 (N_17944,N_16867,N_17185);
xnor U17945 (N_17945,N_17337,N_17392);
and U17946 (N_17946,N_16980,N_17187);
or U17947 (N_17947,N_17257,N_17264);
xnor U17948 (N_17948,N_17139,N_17062);
nand U17949 (N_17949,N_17242,N_17201);
or U17950 (N_17950,N_16954,N_16875);
nor U17951 (N_17951,N_17013,N_17007);
nor U17952 (N_17952,N_16897,N_17223);
and U17953 (N_17953,N_16961,N_17234);
or U17954 (N_17954,N_16961,N_16835);
and U17955 (N_17955,N_17257,N_17190);
and U17956 (N_17956,N_17257,N_17090);
or U17957 (N_17957,N_16956,N_17206);
nor U17958 (N_17958,N_17316,N_16976);
nand U17959 (N_17959,N_17315,N_16849);
and U17960 (N_17960,N_17242,N_17214);
or U17961 (N_17961,N_16894,N_17287);
nor U17962 (N_17962,N_17067,N_16856);
xnor U17963 (N_17963,N_17197,N_17076);
nand U17964 (N_17964,N_16955,N_16805);
xnor U17965 (N_17965,N_17300,N_16862);
and U17966 (N_17966,N_16870,N_17174);
or U17967 (N_17967,N_17166,N_17244);
and U17968 (N_17968,N_16815,N_17140);
nand U17969 (N_17969,N_17129,N_17127);
or U17970 (N_17970,N_16884,N_17117);
or U17971 (N_17971,N_17079,N_17306);
nor U17972 (N_17972,N_16914,N_16882);
xor U17973 (N_17973,N_17091,N_17000);
nand U17974 (N_17974,N_17133,N_17377);
nor U17975 (N_17975,N_16898,N_17139);
nor U17976 (N_17976,N_17380,N_17353);
nand U17977 (N_17977,N_17090,N_17369);
nand U17978 (N_17978,N_16857,N_17112);
nand U17979 (N_17979,N_17123,N_16934);
xor U17980 (N_17980,N_17184,N_17354);
xor U17981 (N_17981,N_17394,N_17221);
or U17982 (N_17982,N_17157,N_16911);
and U17983 (N_17983,N_17286,N_17244);
nand U17984 (N_17984,N_16865,N_17259);
nand U17985 (N_17985,N_16813,N_17035);
nor U17986 (N_17986,N_16863,N_17331);
nor U17987 (N_17987,N_16937,N_17271);
and U17988 (N_17988,N_17035,N_16823);
xnor U17989 (N_17989,N_16941,N_16808);
or U17990 (N_17990,N_17147,N_17163);
xor U17991 (N_17991,N_17268,N_16843);
or U17992 (N_17992,N_17189,N_16872);
or U17993 (N_17993,N_17134,N_17318);
xor U17994 (N_17994,N_17279,N_17359);
nand U17995 (N_17995,N_17202,N_17330);
or U17996 (N_17996,N_17135,N_17166);
xor U17997 (N_17997,N_16878,N_16856);
nand U17998 (N_17998,N_17264,N_17185);
nor U17999 (N_17999,N_17274,N_16974);
nand U18000 (N_18000,N_17555,N_17737);
and U18001 (N_18001,N_17536,N_17569);
nor U18002 (N_18002,N_17979,N_17650);
xor U18003 (N_18003,N_17919,N_17873);
nand U18004 (N_18004,N_17710,N_17408);
nor U18005 (N_18005,N_17797,N_17869);
nand U18006 (N_18006,N_17912,N_17537);
xor U18007 (N_18007,N_17896,N_17744);
nand U18008 (N_18008,N_17692,N_17637);
and U18009 (N_18009,N_17841,N_17808);
and U18010 (N_18010,N_17551,N_17751);
and U18011 (N_18011,N_17681,N_17711);
nor U18012 (N_18012,N_17554,N_17724);
xor U18013 (N_18013,N_17830,N_17811);
or U18014 (N_18014,N_17431,N_17453);
or U18015 (N_18015,N_17831,N_17798);
xor U18016 (N_18016,N_17463,N_17634);
or U18017 (N_18017,N_17683,N_17604);
nor U18018 (N_18018,N_17496,N_17556);
xor U18019 (N_18019,N_17427,N_17660);
nor U18020 (N_18020,N_17937,N_17430);
and U18021 (N_18021,N_17647,N_17949);
and U18022 (N_18022,N_17789,N_17809);
xnor U18023 (N_18023,N_17868,N_17886);
nor U18024 (N_18024,N_17622,N_17516);
nor U18025 (N_18025,N_17471,N_17879);
nand U18026 (N_18026,N_17953,N_17617);
xor U18027 (N_18027,N_17701,N_17964);
nand U18028 (N_18028,N_17768,N_17638);
xor U18029 (N_18029,N_17497,N_17699);
nor U18030 (N_18030,N_17400,N_17917);
and U18031 (N_18031,N_17653,N_17455);
xor U18032 (N_18032,N_17958,N_17574);
and U18033 (N_18033,N_17575,N_17695);
and U18034 (N_18034,N_17872,N_17483);
and U18035 (N_18035,N_17926,N_17678);
xor U18036 (N_18036,N_17505,N_17515);
xnor U18037 (N_18037,N_17717,N_17754);
or U18038 (N_18038,N_17777,N_17719);
or U18039 (N_18039,N_17694,N_17942);
or U18040 (N_18040,N_17538,N_17527);
nand U18041 (N_18041,N_17928,N_17863);
and U18042 (N_18042,N_17693,N_17871);
nor U18043 (N_18043,N_17716,N_17757);
xor U18044 (N_18044,N_17742,N_17908);
and U18045 (N_18045,N_17761,N_17878);
xnor U18046 (N_18046,N_17741,N_17578);
xor U18047 (N_18047,N_17838,N_17685);
and U18048 (N_18048,N_17839,N_17881);
or U18049 (N_18049,N_17891,N_17880);
nor U18050 (N_18050,N_17974,N_17682);
and U18051 (N_18051,N_17429,N_17804);
nand U18052 (N_18052,N_17606,N_17907);
nor U18053 (N_18053,N_17733,N_17959);
xor U18054 (N_18054,N_17452,N_17985);
or U18055 (N_18055,N_17602,N_17619);
or U18056 (N_18056,N_17434,N_17465);
or U18057 (N_18057,N_17491,N_17406);
and U18058 (N_18058,N_17626,N_17528);
nand U18059 (N_18059,N_17844,N_17734);
and U18060 (N_18060,N_17627,N_17495);
nand U18061 (N_18061,N_17760,N_17616);
xnor U18062 (N_18062,N_17461,N_17725);
nor U18063 (N_18063,N_17915,N_17955);
xnor U18064 (N_18064,N_17920,N_17791);
and U18065 (N_18065,N_17781,N_17753);
nor U18066 (N_18066,N_17988,N_17864);
nor U18067 (N_18067,N_17680,N_17691);
xnor U18068 (N_18068,N_17600,N_17493);
and U18069 (N_18069,N_17425,N_17826);
nor U18070 (N_18070,N_17969,N_17727);
nand U18071 (N_18071,N_17519,N_17842);
and U18072 (N_18072,N_17906,N_17910);
and U18073 (N_18073,N_17747,N_17410);
and U18074 (N_18074,N_17549,N_17825);
and U18075 (N_18075,N_17518,N_17552);
nor U18076 (N_18076,N_17419,N_17480);
or U18077 (N_18077,N_17933,N_17892);
or U18078 (N_18078,N_17980,N_17870);
nand U18079 (N_18079,N_17944,N_17560);
xnor U18080 (N_18080,N_17963,N_17628);
or U18081 (N_18081,N_17846,N_17588);
nor U18082 (N_18082,N_17814,N_17758);
nor U18083 (N_18083,N_17584,N_17946);
or U18084 (N_18084,N_17581,N_17609);
or U18085 (N_18085,N_17776,N_17904);
or U18086 (N_18086,N_17561,N_17573);
or U18087 (N_18087,N_17509,N_17981);
xnor U18088 (N_18088,N_17404,N_17459);
and U18089 (N_18089,N_17477,N_17894);
or U18090 (N_18090,N_17925,N_17800);
and U18091 (N_18091,N_17921,N_17486);
nor U18092 (N_18092,N_17918,N_17531);
or U18093 (N_18093,N_17771,N_17572);
nor U18094 (N_18094,N_17625,N_17458);
nand U18095 (N_18095,N_17793,N_17952);
or U18096 (N_18096,N_17859,N_17828);
nand U18097 (N_18097,N_17893,N_17645);
or U18098 (N_18098,N_17792,N_17610);
or U18099 (N_18099,N_17690,N_17728);
nor U18100 (N_18100,N_17414,N_17684);
nor U18101 (N_18101,N_17655,N_17442);
xor U18102 (N_18102,N_17468,N_17855);
or U18103 (N_18103,N_17704,N_17905);
and U18104 (N_18104,N_17470,N_17848);
nand U18105 (N_18105,N_17794,N_17764);
and U18106 (N_18106,N_17767,N_17731);
and U18107 (N_18107,N_17931,N_17580);
xnor U18108 (N_18108,N_17759,N_17829);
nor U18109 (N_18109,N_17916,N_17909);
or U18110 (N_18110,N_17750,N_17577);
and U18111 (N_18111,N_17987,N_17526);
xor U18112 (N_18112,N_17624,N_17890);
and U18113 (N_18113,N_17436,N_17620);
xor U18114 (N_18114,N_17899,N_17428);
or U18115 (N_18115,N_17490,N_17709);
nor U18116 (N_18116,N_17854,N_17484);
or U18117 (N_18117,N_17752,N_17932);
xor U18118 (N_18118,N_17827,N_17562);
nor U18119 (N_18119,N_17721,N_17999);
nand U18120 (N_18120,N_17478,N_17521);
or U18121 (N_18121,N_17559,N_17822);
and U18122 (N_18122,N_17755,N_17674);
nand U18123 (N_18123,N_17523,N_17661);
nand U18124 (N_18124,N_17778,N_17707);
and U18125 (N_18125,N_17417,N_17457);
nand U18126 (N_18126,N_17849,N_17611);
or U18127 (N_18127,N_17499,N_17621);
xnor U18128 (N_18128,N_17927,N_17662);
or U18129 (N_18129,N_17762,N_17874);
nor U18130 (N_18130,N_17698,N_17433);
xor U18131 (N_18131,N_17903,N_17666);
nand U18132 (N_18132,N_17501,N_17677);
nand U18133 (N_18133,N_17550,N_17901);
nor U18134 (N_18134,N_17481,N_17877);
and U18135 (N_18135,N_17412,N_17913);
or U18136 (N_18136,N_17633,N_17663);
and U18137 (N_18137,N_17643,N_17595);
nor U18138 (N_18138,N_17875,N_17783);
or U18139 (N_18139,N_17858,N_17966);
nand U18140 (N_18140,N_17649,N_17943);
or U18141 (N_18141,N_17876,N_17902);
or U18142 (N_18142,N_17467,N_17494);
xor U18143 (N_18143,N_17785,N_17788);
and U18144 (N_18144,N_17997,N_17539);
and U18145 (N_18145,N_17743,N_17938);
and U18146 (N_18146,N_17437,N_17571);
nand U18147 (N_18147,N_17962,N_17658);
nand U18148 (N_18148,N_17968,N_17636);
nand U18149 (N_18149,N_17651,N_17608);
and U18150 (N_18150,N_17503,N_17508);
and U18151 (N_18151,N_17534,N_17813);
or U18152 (N_18152,N_17883,N_17590);
or U18153 (N_18153,N_17840,N_17469);
xor U18154 (N_18154,N_17605,N_17973);
xor U18155 (N_18155,N_17450,N_17506);
or U18156 (N_18156,N_17914,N_17948);
and U18157 (N_18157,N_17566,N_17451);
and U18158 (N_18158,N_17440,N_17697);
nor U18159 (N_18159,N_17441,N_17488);
nor U18160 (N_18160,N_17687,N_17887);
xnor U18161 (N_18161,N_17654,N_17945);
nand U18162 (N_18162,N_17796,N_17889);
and U18163 (N_18163,N_17866,N_17422);
and U18164 (N_18164,N_17565,N_17439);
nand U18165 (N_18165,N_17802,N_17558);
xor U18166 (N_18166,N_17736,N_17689);
nor U18167 (N_18167,N_17585,N_17473);
or U18168 (N_18168,N_17702,N_17991);
or U18169 (N_18169,N_17447,N_17517);
nand U18170 (N_18170,N_17639,N_17535);
nor U18171 (N_18171,N_17485,N_17756);
nor U18172 (N_18172,N_17888,N_17557);
or U18173 (N_18173,N_17489,N_17409);
and U18174 (N_18174,N_17775,N_17583);
xor U18175 (N_18175,N_17589,N_17564);
or U18176 (N_18176,N_17403,N_17712);
nor U18177 (N_18177,N_17487,N_17730);
or U18178 (N_18178,N_17543,N_17420);
nand U18179 (N_18179,N_17772,N_17718);
nand U18180 (N_18180,N_17786,N_17570);
nor U18181 (N_18181,N_17726,N_17510);
xnor U18182 (N_18182,N_17832,N_17615);
and U18183 (N_18183,N_17851,N_17445);
or U18184 (N_18184,N_17415,N_17923);
nor U18185 (N_18185,N_17976,N_17700);
and U18186 (N_18186,N_17579,N_17852);
nor U18187 (N_18187,N_17644,N_17567);
and U18188 (N_18188,N_17706,N_17446);
or U18189 (N_18189,N_17820,N_17462);
nor U18190 (N_18190,N_17970,N_17629);
or U18191 (N_18191,N_17703,N_17763);
nor U18192 (N_18192,N_17657,N_17476);
nor U18193 (N_18193,N_17464,N_17432);
nor U18194 (N_18194,N_17738,N_17965);
or U18195 (N_18195,N_17688,N_17454);
nor U18196 (N_18196,N_17546,N_17438);
xor U18197 (N_18197,N_17770,N_17834);
and U18198 (N_18198,N_17930,N_17421);
nor U18199 (N_18199,N_17669,N_17568);
or U18200 (N_18200,N_17790,N_17735);
nand U18201 (N_18201,N_17401,N_17635);
and U18202 (N_18202,N_17998,N_17835);
xor U18203 (N_18203,N_17500,N_17612);
xnor U18204 (N_18204,N_17641,N_17787);
or U18205 (N_18205,N_17652,N_17954);
nor U18206 (N_18206,N_17975,N_17823);
xor U18207 (N_18207,N_17847,N_17540);
xor U18208 (N_18208,N_17672,N_17774);
nor U18209 (N_18209,N_17676,N_17614);
and U18210 (N_18210,N_17411,N_17845);
xnor U18211 (N_18211,N_17642,N_17631);
xnor U18212 (N_18212,N_17522,N_17593);
or U18213 (N_18213,N_17824,N_17591);
xor U18214 (N_18214,N_17547,N_17897);
and U18215 (N_18215,N_17967,N_17670);
nor U18216 (N_18216,N_17746,N_17782);
nand U18217 (N_18217,N_17935,N_17984);
or U18218 (N_18218,N_17630,N_17860);
nor U18219 (N_18219,N_17837,N_17780);
nand U18220 (N_18220,N_17696,N_17582);
and U18221 (N_18221,N_17514,N_17597);
nand U18222 (N_18222,N_17934,N_17424);
nor U18223 (N_18223,N_17911,N_17990);
nor U18224 (N_18224,N_17773,N_17995);
nor U18225 (N_18225,N_17563,N_17989);
nor U18226 (N_18226,N_17607,N_17993);
and U18227 (N_18227,N_17407,N_17542);
xnor U18228 (N_18228,N_17882,N_17686);
nor U18229 (N_18229,N_17994,N_17951);
xnor U18230 (N_18230,N_17532,N_17548);
xor U18231 (N_18231,N_17795,N_17895);
and U18232 (N_18232,N_17807,N_17996);
xnor U18233 (N_18233,N_17596,N_17766);
and U18234 (N_18234,N_17603,N_17972);
nor U18235 (N_18235,N_17474,N_17599);
or U18236 (N_18236,N_17803,N_17833);
and U18237 (N_18237,N_17720,N_17623);
and U18238 (N_18238,N_17665,N_17957);
and U18239 (N_18239,N_17544,N_17405);
or U18240 (N_18240,N_17668,N_17507);
and U18241 (N_18241,N_17656,N_17664);
xor U18242 (N_18242,N_17836,N_17466);
xnor U18243 (N_18243,N_17511,N_17884);
nor U18244 (N_18244,N_17502,N_17817);
or U18245 (N_18245,N_17983,N_17520);
xor U18246 (N_18246,N_17533,N_17479);
and U18247 (N_18247,N_17857,N_17867);
or U18248 (N_18248,N_17805,N_17416);
nor U18249 (N_18249,N_17504,N_17861);
xnor U18250 (N_18250,N_17971,N_17856);
nor U18251 (N_18251,N_17667,N_17444);
xnor U18252 (N_18252,N_17413,N_17929);
and U18253 (N_18253,N_17482,N_17982);
and U18254 (N_18254,N_17806,N_17799);
nand U18255 (N_18255,N_17426,N_17940);
xnor U18256 (N_18256,N_17705,N_17443);
nand U18257 (N_18257,N_17545,N_17475);
or U18258 (N_18258,N_17449,N_17941);
nor U18259 (N_18259,N_17541,N_17819);
or U18260 (N_18260,N_17801,N_17865);
nand U18261 (N_18261,N_17749,N_17818);
xor U18262 (N_18262,N_17936,N_17922);
xnor U18263 (N_18263,N_17885,N_17722);
nand U18264 (N_18264,N_17423,N_17843);
nor U18265 (N_18265,N_17524,N_17853);
xnor U18266 (N_18266,N_17812,N_17513);
or U18267 (N_18267,N_17779,N_17769);
nor U18268 (N_18268,N_17810,N_17632);
nand U18269 (N_18269,N_17448,N_17598);
nor U18270 (N_18270,N_17950,N_17460);
or U18271 (N_18271,N_17529,N_17618);
and U18272 (N_18272,N_17530,N_17765);
and U18273 (N_18273,N_17498,N_17732);
xor U18274 (N_18274,N_17594,N_17472);
nand U18275 (N_18275,N_17418,N_17613);
and U18276 (N_18276,N_17402,N_17723);
and U18277 (N_18277,N_17850,N_17992);
nor U18278 (N_18278,N_17592,N_17715);
xor U18279 (N_18279,N_17714,N_17977);
and U18280 (N_18280,N_17956,N_17659);
and U18281 (N_18281,N_17947,N_17512);
and U18282 (N_18282,N_17961,N_17740);
xnor U18283 (N_18283,N_17745,N_17708);
nand U18284 (N_18284,N_17576,N_17587);
xnor U18285 (N_18285,N_17816,N_17815);
and U18286 (N_18286,N_17640,N_17675);
or U18287 (N_18287,N_17671,N_17586);
or U18288 (N_18288,N_17492,N_17784);
xnor U18289 (N_18289,N_17748,N_17646);
xor U18290 (N_18290,N_17939,N_17601);
nand U18291 (N_18291,N_17648,N_17456);
nand U18292 (N_18292,N_17986,N_17739);
nand U18293 (N_18293,N_17924,N_17673);
nor U18294 (N_18294,N_17713,N_17729);
nand U18295 (N_18295,N_17553,N_17978);
xnor U18296 (N_18296,N_17960,N_17525);
nor U18297 (N_18297,N_17679,N_17862);
and U18298 (N_18298,N_17821,N_17435);
and U18299 (N_18299,N_17900,N_17898);
and U18300 (N_18300,N_17598,N_17958);
xnor U18301 (N_18301,N_17822,N_17925);
and U18302 (N_18302,N_17427,N_17787);
or U18303 (N_18303,N_17444,N_17511);
xor U18304 (N_18304,N_17758,N_17871);
and U18305 (N_18305,N_17677,N_17785);
xnor U18306 (N_18306,N_17544,N_17713);
nand U18307 (N_18307,N_17494,N_17804);
xor U18308 (N_18308,N_17440,N_17530);
nand U18309 (N_18309,N_17912,N_17619);
and U18310 (N_18310,N_17943,N_17641);
xnor U18311 (N_18311,N_17687,N_17498);
and U18312 (N_18312,N_17898,N_17770);
nand U18313 (N_18313,N_17633,N_17634);
nor U18314 (N_18314,N_17689,N_17832);
nor U18315 (N_18315,N_17601,N_17986);
or U18316 (N_18316,N_17947,N_17953);
nand U18317 (N_18317,N_17655,N_17665);
and U18318 (N_18318,N_17812,N_17443);
nand U18319 (N_18319,N_17468,N_17470);
or U18320 (N_18320,N_17473,N_17508);
xnor U18321 (N_18321,N_17473,N_17990);
and U18322 (N_18322,N_17528,N_17620);
xor U18323 (N_18323,N_17435,N_17443);
and U18324 (N_18324,N_17426,N_17859);
and U18325 (N_18325,N_17647,N_17972);
and U18326 (N_18326,N_17410,N_17849);
or U18327 (N_18327,N_17932,N_17685);
xnor U18328 (N_18328,N_17610,N_17681);
nor U18329 (N_18329,N_17587,N_17673);
nand U18330 (N_18330,N_17825,N_17503);
nor U18331 (N_18331,N_17530,N_17713);
or U18332 (N_18332,N_17827,N_17756);
and U18333 (N_18333,N_17485,N_17526);
and U18334 (N_18334,N_17708,N_17815);
xor U18335 (N_18335,N_17857,N_17436);
nand U18336 (N_18336,N_17652,N_17513);
or U18337 (N_18337,N_17934,N_17444);
xnor U18338 (N_18338,N_17424,N_17907);
nand U18339 (N_18339,N_17698,N_17736);
or U18340 (N_18340,N_17814,N_17889);
nand U18341 (N_18341,N_17690,N_17469);
nand U18342 (N_18342,N_17416,N_17549);
nand U18343 (N_18343,N_17788,N_17547);
nand U18344 (N_18344,N_17679,N_17473);
nand U18345 (N_18345,N_17675,N_17908);
or U18346 (N_18346,N_17715,N_17678);
nand U18347 (N_18347,N_17620,N_17854);
nand U18348 (N_18348,N_17495,N_17976);
nor U18349 (N_18349,N_17898,N_17807);
or U18350 (N_18350,N_17475,N_17868);
or U18351 (N_18351,N_17421,N_17478);
nor U18352 (N_18352,N_17501,N_17782);
or U18353 (N_18353,N_17869,N_17926);
and U18354 (N_18354,N_17593,N_17874);
nand U18355 (N_18355,N_17466,N_17815);
nand U18356 (N_18356,N_17809,N_17896);
nand U18357 (N_18357,N_17489,N_17971);
and U18358 (N_18358,N_17449,N_17538);
and U18359 (N_18359,N_17632,N_17593);
nand U18360 (N_18360,N_17793,N_17858);
nand U18361 (N_18361,N_17737,N_17644);
or U18362 (N_18362,N_17968,N_17829);
nand U18363 (N_18363,N_17492,N_17448);
or U18364 (N_18364,N_17705,N_17922);
nand U18365 (N_18365,N_17864,N_17829);
nand U18366 (N_18366,N_17436,N_17628);
nand U18367 (N_18367,N_17764,N_17990);
or U18368 (N_18368,N_17535,N_17647);
or U18369 (N_18369,N_17576,N_17400);
or U18370 (N_18370,N_17917,N_17555);
nand U18371 (N_18371,N_17688,N_17976);
nor U18372 (N_18372,N_17806,N_17681);
nor U18373 (N_18373,N_17622,N_17962);
or U18374 (N_18374,N_17410,N_17798);
xor U18375 (N_18375,N_17598,N_17878);
nand U18376 (N_18376,N_17856,N_17952);
or U18377 (N_18377,N_17749,N_17786);
xnor U18378 (N_18378,N_17957,N_17697);
or U18379 (N_18379,N_17759,N_17808);
nor U18380 (N_18380,N_17683,N_17760);
and U18381 (N_18381,N_17663,N_17696);
and U18382 (N_18382,N_17898,N_17880);
or U18383 (N_18383,N_17843,N_17522);
and U18384 (N_18384,N_17412,N_17661);
xor U18385 (N_18385,N_17476,N_17920);
or U18386 (N_18386,N_17605,N_17923);
nor U18387 (N_18387,N_17911,N_17729);
and U18388 (N_18388,N_17628,N_17943);
xnor U18389 (N_18389,N_17708,N_17725);
xor U18390 (N_18390,N_17595,N_17641);
nand U18391 (N_18391,N_17539,N_17744);
or U18392 (N_18392,N_17685,N_17912);
xnor U18393 (N_18393,N_17901,N_17789);
nor U18394 (N_18394,N_17534,N_17527);
or U18395 (N_18395,N_17509,N_17445);
nand U18396 (N_18396,N_17456,N_17757);
and U18397 (N_18397,N_17850,N_17777);
or U18398 (N_18398,N_17437,N_17996);
and U18399 (N_18399,N_17469,N_17432);
and U18400 (N_18400,N_17482,N_17671);
and U18401 (N_18401,N_17852,N_17896);
nor U18402 (N_18402,N_17658,N_17947);
nor U18403 (N_18403,N_17720,N_17975);
nand U18404 (N_18404,N_17743,N_17616);
nand U18405 (N_18405,N_17444,N_17977);
nor U18406 (N_18406,N_17563,N_17678);
and U18407 (N_18407,N_17924,N_17500);
and U18408 (N_18408,N_17407,N_17732);
and U18409 (N_18409,N_17961,N_17631);
nand U18410 (N_18410,N_17680,N_17815);
and U18411 (N_18411,N_17509,N_17896);
or U18412 (N_18412,N_17858,N_17641);
nor U18413 (N_18413,N_17738,N_17929);
and U18414 (N_18414,N_17583,N_17826);
nand U18415 (N_18415,N_17789,N_17592);
or U18416 (N_18416,N_17870,N_17650);
nand U18417 (N_18417,N_17911,N_17901);
or U18418 (N_18418,N_17515,N_17831);
xor U18419 (N_18419,N_17539,N_17905);
nand U18420 (N_18420,N_17565,N_17400);
and U18421 (N_18421,N_17971,N_17478);
nor U18422 (N_18422,N_17937,N_17656);
and U18423 (N_18423,N_17697,N_17926);
and U18424 (N_18424,N_17422,N_17771);
or U18425 (N_18425,N_17455,N_17543);
xnor U18426 (N_18426,N_17920,N_17456);
xnor U18427 (N_18427,N_17655,N_17501);
xnor U18428 (N_18428,N_17731,N_17832);
nor U18429 (N_18429,N_17749,N_17510);
and U18430 (N_18430,N_17738,N_17628);
nand U18431 (N_18431,N_17569,N_17515);
nor U18432 (N_18432,N_17981,N_17776);
nor U18433 (N_18433,N_17477,N_17540);
and U18434 (N_18434,N_17706,N_17661);
or U18435 (N_18435,N_17699,N_17844);
or U18436 (N_18436,N_17722,N_17419);
or U18437 (N_18437,N_17669,N_17813);
xor U18438 (N_18438,N_17832,N_17500);
nor U18439 (N_18439,N_17956,N_17827);
nand U18440 (N_18440,N_17699,N_17995);
xor U18441 (N_18441,N_17977,N_17512);
nand U18442 (N_18442,N_17655,N_17836);
or U18443 (N_18443,N_17729,N_17842);
nand U18444 (N_18444,N_17529,N_17930);
nand U18445 (N_18445,N_17953,N_17680);
nand U18446 (N_18446,N_17599,N_17917);
or U18447 (N_18447,N_17924,N_17742);
or U18448 (N_18448,N_17438,N_17698);
nand U18449 (N_18449,N_17592,N_17455);
nor U18450 (N_18450,N_17514,N_17538);
nand U18451 (N_18451,N_17819,N_17652);
nand U18452 (N_18452,N_17407,N_17408);
nand U18453 (N_18453,N_17622,N_17514);
or U18454 (N_18454,N_17931,N_17601);
and U18455 (N_18455,N_17618,N_17999);
nor U18456 (N_18456,N_17559,N_17589);
nand U18457 (N_18457,N_17580,N_17681);
nand U18458 (N_18458,N_17573,N_17542);
nand U18459 (N_18459,N_17935,N_17458);
and U18460 (N_18460,N_17976,N_17729);
nor U18461 (N_18461,N_17568,N_17666);
nor U18462 (N_18462,N_17968,N_17551);
or U18463 (N_18463,N_17484,N_17848);
or U18464 (N_18464,N_17545,N_17496);
nand U18465 (N_18465,N_17936,N_17790);
and U18466 (N_18466,N_17632,N_17840);
or U18467 (N_18467,N_17703,N_17944);
or U18468 (N_18468,N_17978,N_17965);
xor U18469 (N_18469,N_17880,N_17853);
and U18470 (N_18470,N_17880,N_17496);
and U18471 (N_18471,N_17554,N_17692);
or U18472 (N_18472,N_17747,N_17975);
nand U18473 (N_18473,N_17497,N_17628);
and U18474 (N_18474,N_17994,N_17430);
nor U18475 (N_18475,N_17869,N_17542);
or U18476 (N_18476,N_17455,N_17559);
and U18477 (N_18477,N_17771,N_17436);
nor U18478 (N_18478,N_17687,N_17797);
nand U18479 (N_18479,N_17403,N_17703);
xnor U18480 (N_18480,N_17790,N_17795);
and U18481 (N_18481,N_17534,N_17726);
nand U18482 (N_18482,N_17726,N_17464);
nor U18483 (N_18483,N_17518,N_17634);
or U18484 (N_18484,N_17626,N_17448);
xnor U18485 (N_18485,N_17877,N_17680);
xnor U18486 (N_18486,N_17940,N_17680);
nor U18487 (N_18487,N_17788,N_17437);
or U18488 (N_18488,N_17834,N_17962);
or U18489 (N_18489,N_17700,N_17901);
and U18490 (N_18490,N_17753,N_17413);
nand U18491 (N_18491,N_17687,N_17828);
and U18492 (N_18492,N_17759,N_17897);
nand U18493 (N_18493,N_17571,N_17549);
nand U18494 (N_18494,N_17903,N_17777);
and U18495 (N_18495,N_17995,N_17402);
nor U18496 (N_18496,N_17923,N_17557);
xnor U18497 (N_18497,N_17658,N_17883);
nor U18498 (N_18498,N_17715,N_17958);
or U18499 (N_18499,N_17931,N_17517);
xnor U18500 (N_18500,N_17738,N_17749);
and U18501 (N_18501,N_17731,N_17476);
nor U18502 (N_18502,N_17604,N_17841);
and U18503 (N_18503,N_17492,N_17718);
nor U18504 (N_18504,N_17691,N_17659);
nand U18505 (N_18505,N_17702,N_17437);
nand U18506 (N_18506,N_17709,N_17851);
or U18507 (N_18507,N_17716,N_17958);
or U18508 (N_18508,N_17687,N_17561);
nand U18509 (N_18509,N_17973,N_17696);
nor U18510 (N_18510,N_17867,N_17441);
and U18511 (N_18511,N_17737,N_17846);
and U18512 (N_18512,N_17754,N_17618);
or U18513 (N_18513,N_17690,N_17454);
xor U18514 (N_18514,N_17724,N_17442);
nor U18515 (N_18515,N_17531,N_17746);
xnor U18516 (N_18516,N_17683,N_17485);
nor U18517 (N_18517,N_17402,N_17896);
or U18518 (N_18518,N_17952,N_17902);
xnor U18519 (N_18519,N_17516,N_17463);
nor U18520 (N_18520,N_17451,N_17542);
and U18521 (N_18521,N_17630,N_17877);
and U18522 (N_18522,N_17903,N_17754);
or U18523 (N_18523,N_17571,N_17676);
xor U18524 (N_18524,N_17628,N_17698);
nand U18525 (N_18525,N_17983,N_17931);
nor U18526 (N_18526,N_17420,N_17786);
nand U18527 (N_18527,N_17977,N_17824);
or U18528 (N_18528,N_17408,N_17516);
xnor U18529 (N_18529,N_17962,N_17585);
and U18530 (N_18530,N_17529,N_17636);
xor U18531 (N_18531,N_17945,N_17688);
xor U18532 (N_18532,N_17525,N_17689);
nor U18533 (N_18533,N_17497,N_17752);
nand U18534 (N_18534,N_17766,N_17845);
or U18535 (N_18535,N_17423,N_17993);
or U18536 (N_18536,N_17873,N_17406);
xor U18537 (N_18537,N_17852,N_17527);
or U18538 (N_18538,N_17975,N_17493);
or U18539 (N_18539,N_17994,N_17811);
xnor U18540 (N_18540,N_17610,N_17552);
xor U18541 (N_18541,N_17617,N_17949);
nor U18542 (N_18542,N_17520,N_17900);
and U18543 (N_18543,N_17885,N_17701);
or U18544 (N_18544,N_17445,N_17659);
or U18545 (N_18545,N_17963,N_17636);
and U18546 (N_18546,N_17806,N_17724);
xnor U18547 (N_18547,N_17456,N_17591);
nor U18548 (N_18548,N_17818,N_17647);
or U18549 (N_18549,N_17557,N_17592);
xnor U18550 (N_18550,N_17978,N_17805);
xor U18551 (N_18551,N_17429,N_17514);
or U18552 (N_18552,N_17481,N_17756);
or U18553 (N_18553,N_17572,N_17896);
nand U18554 (N_18554,N_17689,N_17670);
xor U18555 (N_18555,N_17840,N_17822);
or U18556 (N_18556,N_17500,N_17681);
or U18557 (N_18557,N_17700,N_17937);
or U18558 (N_18558,N_17465,N_17484);
nor U18559 (N_18559,N_17932,N_17978);
or U18560 (N_18560,N_17548,N_17526);
nand U18561 (N_18561,N_17836,N_17476);
nor U18562 (N_18562,N_17597,N_17625);
or U18563 (N_18563,N_17463,N_17459);
and U18564 (N_18564,N_17843,N_17466);
and U18565 (N_18565,N_17871,N_17477);
and U18566 (N_18566,N_17475,N_17846);
and U18567 (N_18567,N_17476,N_17923);
and U18568 (N_18568,N_17908,N_17890);
xnor U18569 (N_18569,N_17520,N_17730);
nand U18570 (N_18570,N_17417,N_17582);
nor U18571 (N_18571,N_17597,N_17576);
and U18572 (N_18572,N_17488,N_17871);
xor U18573 (N_18573,N_17883,N_17831);
nor U18574 (N_18574,N_17569,N_17974);
xnor U18575 (N_18575,N_17689,N_17785);
nand U18576 (N_18576,N_17783,N_17716);
xnor U18577 (N_18577,N_17770,N_17914);
and U18578 (N_18578,N_17459,N_17723);
nand U18579 (N_18579,N_17535,N_17822);
xnor U18580 (N_18580,N_17712,N_17759);
nor U18581 (N_18581,N_17755,N_17876);
nand U18582 (N_18582,N_17924,N_17611);
or U18583 (N_18583,N_17735,N_17593);
nor U18584 (N_18584,N_17677,N_17482);
xnor U18585 (N_18585,N_17502,N_17630);
xnor U18586 (N_18586,N_17440,N_17428);
xor U18587 (N_18587,N_17869,N_17848);
and U18588 (N_18588,N_17487,N_17510);
nand U18589 (N_18589,N_17598,N_17938);
xnor U18590 (N_18590,N_17431,N_17813);
and U18591 (N_18591,N_17730,N_17927);
and U18592 (N_18592,N_17689,N_17481);
and U18593 (N_18593,N_17979,N_17736);
nand U18594 (N_18594,N_17541,N_17833);
and U18595 (N_18595,N_17949,N_17983);
and U18596 (N_18596,N_17409,N_17807);
or U18597 (N_18597,N_17477,N_17743);
xnor U18598 (N_18598,N_17697,N_17566);
and U18599 (N_18599,N_17660,N_17743);
nor U18600 (N_18600,N_18106,N_18245);
nor U18601 (N_18601,N_18588,N_18034);
or U18602 (N_18602,N_18208,N_18472);
xnor U18603 (N_18603,N_18187,N_18394);
and U18604 (N_18604,N_18398,N_18199);
nand U18605 (N_18605,N_18100,N_18161);
and U18606 (N_18606,N_18184,N_18236);
nand U18607 (N_18607,N_18559,N_18082);
and U18608 (N_18608,N_18235,N_18003);
nor U18609 (N_18609,N_18299,N_18462);
xnor U18610 (N_18610,N_18572,N_18223);
and U18611 (N_18611,N_18586,N_18560);
nand U18612 (N_18612,N_18104,N_18538);
nand U18613 (N_18613,N_18160,N_18022);
xor U18614 (N_18614,N_18374,N_18469);
nor U18615 (N_18615,N_18585,N_18062);
xor U18616 (N_18616,N_18190,N_18259);
nor U18617 (N_18617,N_18308,N_18088);
and U18618 (N_18618,N_18587,N_18295);
nor U18619 (N_18619,N_18098,N_18416);
xor U18620 (N_18620,N_18101,N_18495);
nor U18621 (N_18621,N_18047,N_18116);
or U18622 (N_18622,N_18499,N_18211);
and U18623 (N_18623,N_18215,N_18217);
xnor U18624 (N_18624,N_18410,N_18340);
or U18625 (N_18625,N_18377,N_18146);
xnor U18626 (N_18626,N_18372,N_18253);
nand U18627 (N_18627,N_18352,N_18451);
nor U18628 (N_18628,N_18420,N_18418);
xnor U18629 (N_18629,N_18156,N_18511);
and U18630 (N_18630,N_18243,N_18168);
and U18631 (N_18631,N_18090,N_18431);
nor U18632 (N_18632,N_18520,N_18300);
xnor U18633 (N_18633,N_18458,N_18183);
and U18634 (N_18634,N_18118,N_18096);
and U18635 (N_18635,N_18388,N_18379);
and U18636 (N_18636,N_18207,N_18138);
nor U18637 (N_18637,N_18076,N_18396);
and U18638 (N_18638,N_18162,N_18565);
or U18639 (N_18639,N_18570,N_18525);
and U18640 (N_18640,N_18544,N_18290);
nand U18641 (N_18641,N_18338,N_18529);
or U18642 (N_18642,N_18046,N_18074);
nand U18643 (N_18643,N_18255,N_18467);
nand U18644 (N_18644,N_18204,N_18005);
and U18645 (N_18645,N_18256,N_18021);
nand U18646 (N_18646,N_18378,N_18288);
nor U18647 (N_18647,N_18030,N_18350);
and U18648 (N_18648,N_18287,N_18455);
nor U18649 (N_18649,N_18576,N_18368);
xnor U18650 (N_18650,N_18402,N_18342);
nor U18651 (N_18651,N_18522,N_18506);
nor U18652 (N_18652,N_18203,N_18250);
nor U18653 (N_18653,N_18234,N_18466);
or U18654 (N_18654,N_18513,N_18452);
nor U18655 (N_18655,N_18218,N_18397);
or U18656 (N_18656,N_18248,N_18284);
and U18657 (N_18657,N_18242,N_18508);
xor U18658 (N_18658,N_18122,N_18584);
xor U18659 (N_18659,N_18464,N_18423);
nor U18660 (N_18660,N_18233,N_18155);
nor U18661 (N_18661,N_18165,N_18043);
xor U18662 (N_18662,N_18442,N_18013);
and U18663 (N_18663,N_18282,N_18583);
nor U18664 (N_18664,N_18126,N_18360);
or U18665 (N_18665,N_18278,N_18450);
and U18666 (N_18666,N_18042,N_18011);
nand U18667 (N_18667,N_18346,N_18487);
and U18668 (N_18668,N_18305,N_18533);
or U18669 (N_18669,N_18335,N_18166);
nor U18670 (N_18670,N_18306,N_18093);
nor U18671 (N_18671,N_18505,N_18198);
or U18672 (N_18672,N_18044,N_18195);
or U18673 (N_18673,N_18324,N_18258);
and U18674 (N_18674,N_18542,N_18390);
and U18675 (N_18675,N_18473,N_18189);
nand U18676 (N_18676,N_18558,N_18114);
and U18677 (N_18677,N_18302,N_18337);
nand U18678 (N_18678,N_18261,N_18417);
nor U18679 (N_18679,N_18079,N_18169);
or U18680 (N_18680,N_18561,N_18105);
or U18681 (N_18681,N_18454,N_18547);
xnor U18682 (N_18682,N_18224,N_18485);
and U18683 (N_18683,N_18099,N_18072);
nand U18684 (N_18684,N_18521,N_18482);
nor U18685 (N_18685,N_18568,N_18170);
or U18686 (N_18686,N_18086,N_18019);
nor U18687 (N_18687,N_18322,N_18317);
and U18688 (N_18688,N_18070,N_18444);
or U18689 (N_18689,N_18094,N_18351);
or U18690 (N_18690,N_18141,N_18589);
nor U18691 (N_18691,N_18391,N_18202);
xor U18692 (N_18692,N_18361,N_18330);
or U18693 (N_18693,N_18219,N_18239);
xor U18694 (N_18694,N_18069,N_18554);
or U18695 (N_18695,N_18220,N_18073);
or U18696 (N_18696,N_18369,N_18212);
nand U18697 (N_18697,N_18075,N_18413);
or U18698 (N_18698,N_18550,N_18225);
nand U18699 (N_18699,N_18216,N_18263);
or U18700 (N_18700,N_18323,N_18051);
nand U18701 (N_18701,N_18310,N_18052);
and U18702 (N_18702,N_18497,N_18380);
and U18703 (N_18703,N_18384,N_18486);
and U18704 (N_18704,N_18392,N_18411);
nor U18705 (N_18705,N_18463,N_18084);
nand U18706 (N_18706,N_18582,N_18498);
nand U18707 (N_18707,N_18065,N_18244);
xnor U18708 (N_18708,N_18325,N_18033);
nand U18709 (N_18709,N_18465,N_18328);
or U18710 (N_18710,N_18415,N_18578);
and U18711 (N_18711,N_18480,N_18446);
and U18712 (N_18712,N_18474,N_18448);
nor U18713 (N_18713,N_18281,N_18347);
nor U18714 (N_18714,N_18481,N_18592);
and U18715 (N_18715,N_18140,N_18327);
or U18716 (N_18716,N_18557,N_18534);
nor U18717 (N_18717,N_18273,N_18006);
nor U18718 (N_18718,N_18389,N_18425);
nor U18719 (N_18719,N_18110,N_18336);
nand U18720 (N_18720,N_18036,N_18175);
nor U18721 (N_18721,N_18320,N_18232);
and U18722 (N_18722,N_18358,N_18018);
or U18723 (N_18723,N_18039,N_18016);
xor U18724 (N_18724,N_18158,N_18268);
and U18725 (N_18725,N_18029,N_18512);
nor U18726 (N_18726,N_18329,N_18428);
nor U18727 (N_18727,N_18265,N_18424);
xor U18728 (N_18728,N_18373,N_18238);
and U18729 (N_18729,N_18237,N_18080);
xnor U18730 (N_18730,N_18254,N_18440);
nor U18731 (N_18731,N_18293,N_18274);
nor U18732 (N_18732,N_18406,N_18004);
nand U18733 (N_18733,N_18438,N_18054);
xor U18734 (N_18734,N_18028,N_18260);
and U18735 (N_18735,N_18154,N_18436);
xor U18736 (N_18736,N_18171,N_18188);
xor U18737 (N_18737,N_18430,N_18083);
and U18738 (N_18738,N_18111,N_18127);
xnor U18739 (N_18739,N_18109,N_18151);
nand U18740 (N_18740,N_18501,N_18333);
xor U18741 (N_18741,N_18177,N_18103);
nand U18742 (N_18742,N_18279,N_18545);
and U18743 (N_18743,N_18055,N_18579);
or U18744 (N_18744,N_18112,N_18400);
nand U18745 (N_18745,N_18291,N_18353);
nor U18746 (N_18746,N_18283,N_18422);
and U18747 (N_18747,N_18546,N_18231);
nor U18748 (N_18748,N_18437,N_18067);
nand U18749 (N_18749,N_18020,N_18500);
and U18750 (N_18750,N_18014,N_18167);
nand U18751 (N_18751,N_18556,N_18599);
nor U18752 (N_18752,N_18569,N_18081);
and U18753 (N_18753,N_18027,N_18227);
and U18754 (N_18754,N_18147,N_18483);
xnor U18755 (N_18755,N_18562,N_18382);
or U18756 (N_18756,N_18364,N_18056);
and U18757 (N_18757,N_18296,N_18276);
or U18758 (N_18758,N_18552,N_18181);
and U18759 (N_18759,N_18386,N_18174);
xnor U18760 (N_18760,N_18385,N_18297);
and U18761 (N_18761,N_18490,N_18179);
nor U18762 (N_18762,N_18272,N_18514);
and U18763 (N_18763,N_18315,N_18157);
and U18764 (N_18764,N_18178,N_18510);
xor U18765 (N_18765,N_18426,N_18045);
and U18766 (N_18766,N_18381,N_18137);
xor U18767 (N_18767,N_18064,N_18148);
nand U18768 (N_18768,N_18433,N_18286);
nor U18769 (N_18769,N_18407,N_18403);
or U18770 (N_18770,N_18247,N_18564);
nand U18771 (N_18771,N_18535,N_18309);
or U18772 (N_18772,N_18077,N_18078);
and U18773 (N_18773,N_18349,N_18476);
nand U18774 (N_18774,N_18206,N_18432);
xnor U18775 (N_18775,N_18316,N_18228);
and U18776 (N_18776,N_18163,N_18097);
and U18777 (N_18777,N_18277,N_18210);
nor U18778 (N_18778,N_18549,N_18015);
xnor U18779 (N_18779,N_18571,N_18341);
xor U18780 (N_18780,N_18376,N_18144);
or U18781 (N_18781,N_18095,N_18230);
nand U18782 (N_18782,N_18201,N_18135);
or U18783 (N_18783,N_18492,N_18326);
or U18784 (N_18784,N_18214,N_18262);
nand U18785 (N_18785,N_18060,N_18577);
xnor U18786 (N_18786,N_18139,N_18573);
nand U18787 (N_18787,N_18401,N_18266);
xnor U18788 (N_18788,N_18257,N_18200);
xor U18789 (N_18789,N_18580,N_18128);
and U18790 (N_18790,N_18477,N_18457);
nand U18791 (N_18791,N_18108,N_18058);
and U18792 (N_18792,N_18197,N_18429);
nand U18793 (N_18793,N_18267,N_18125);
or U18794 (N_18794,N_18383,N_18150);
nor U18795 (N_18795,N_18527,N_18365);
nand U18796 (N_18796,N_18441,N_18493);
or U18797 (N_18797,N_18303,N_18304);
xor U18798 (N_18798,N_18345,N_18551);
xor U18799 (N_18799,N_18504,N_18226);
nor U18800 (N_18800,N_18526,N_18066);
nor U18801 (N_18801,N_18348,N_18123);
nand U18802 (N_18802,N_18598,N_18518);
and U18803 (N_18803,N_18134,N_18143);
nand U18804 (N_18804,N_18354,N_18539);
nand U18805 (N_18805,N_18484,N_18478);
xnor U18806 (N_18806,N_18024,N_18555);
and U18807 (N_18807,N_18591,N_18061);
and U18808 (N_18808,N_18312,N_18435);
nand U18809 (N_18809,N_18593,N_18318);
nand U18810 (N_18810,N_18405,N_18301);
nor U18811 (N_18811,N_18180,N_18581);
xnor U18812 (N_18812,N_18130,N_18121);
xor U18813 (N_18813,N_18037,N_18285);
and U18814 (N_18814,N_18294,N_18362);
nor U18815 (N_18815,N_18159,N_18092);
or U18816 (N_18816,N_18038,N_18087);
or U18817 (N_18817,N_18548,N_18532);
nand U18818 (N_18818,N_18017,N_18468);
nand U18819 (N_18819,N_18434,N_18566);
and U18820 (N_18820,N_18541,N_18205);
and U18821 (N_18821,N_18590,N_18149);
nand U18822 (N_18822,N_18319,N_18222);
nand U18823 (N_18823,N_18343,N_18479);
nand U18824 (N_18824,N_18164,N_18567);
nand U18825 (N_18825,N_18012,N_18192);
xor U18826 (N_18826,N_18241,N_18009);
nand U18827 (N_18827,N_18367,N_18503);
and U18828 (N_18828,N_18563,N_18313);
xor U18829 (N_18829,N_18597,N_18153);
xor U18830 (N_18830,N_18129,N_18445);
nor U18831 (N_18831,N_18289,N_18371);
nand U18832 (N_18832,N_18068,N_18528);
and U18833 (N_18833,N_18213,N_18270);
or U18834 (N_18834,N_18471,N_18307);
nand U18835 (N_18835,N_18404,N_18035);
nor U18836 (N_18836,N_18000,N_18496);
and U18837 (N_18837,N_18524,N_18408);
xnor U18838 (N_18838,N_18182,N_18449);
xnor U18839 (N_18839,N_18459,N_18516);
and U18840 (N_18840,N_18427,N_18530);
and U18841 (N_18841,N_18007,N_18523);
or U18842 (N_18842,N_18049,N_18421);
xnor U18843 (N_18843,N_18531,N_18439);
nor U18844 (N_18844,N_18475,N_18575);
xnor U18845 (N_18845,N_18298,N_18050);
and U18846 (N_18846,N_18387,N_18314);
nand U18847 (N_18847,N_18040,N_18331);
or U18848 (N_18848,N_18540,N_18246);
and U18849 (N_18849,N_18399,N_18023);
or U18850 (N_18850,N_18221,N_18393);
nor U18851 (N_18851,N_18193,N_18063);
nand U18852 (N_18852,N_18186,N_18536);
or U18853 (N_18853,N_18356,N_18113);
xnor U18854 (N_18854,N_18489,N_18395);
nand U18855 (N_18855,N_18332,N_18176);
nor U18856 (N_18856,N_18185,N_18240);
nor U18857 (N_18857,N_18057,N_18574);
or U18858 (N_18858,N_18229,N_18494);
or U18859 (N_18859,N_18488,N_18031);
nand U18860 (N_18860,N_18596,N_18249);
nor U18861 (N_18861,N_18001,N_18460);
or U18862 (N_18862,N_18002,N_18120);
xnor U18863 (N_18863,N_18515,N_18252);
and U18864 (N_18864,N_18537,N_18010);
nor U18865 (N_18865,N_18412,N_18269);
and U18866 (N_18866,N_18152,N_18025);
nor U18867 (N_18867,N_18366,N_18502);
nor U18868 (N_18868,N_18447,N_18131);
nor U18869 (N_18869,N_18119,N_18355);
and U18870 (N_18870,N_18102,N_18594);
or U18871 (N_18871,N_18048,N_18519);
or U18872 (N_18872,N_18370,N_18264);
xor U18873 (N_18873,N_18089,N_18507);
nor U18874 (N_18874,N_18173,N_18194);
or U18875 (N_18875,N_18543,N_18132);
nor U18876 (N_18876,N_18359,N_18311);
or U18877 (N_18877,N_18461,N_18145);
or U18878 (N_18878,N_18071,N_18491);
nand U18879 (N_18879,N_18209,N_18059);
nor U18880 (N_18880,N_18032,N_18595);
nand U18881 (N_18881,N_18453,N_18136);
or U18882 (N_18882,N_18419,N_18091);
xor U18883 (N_18883,N_18142,N_18172);
nor U18884 (N_18884,N_18344,N_18470);
nor U18885 (N_18885,N_18509,N_18280);
xor U18886 (N_18886,N_18133,N_18191);
nand U18887 (N_18887,N_18443,N_18053);
or U18888 (N_18888,N_18196,N_18375);
and U18889 (N_18889,N_18275,N_18357);
nand U18890 (N_18890,N_18334,N_18517);
xor U18891 (N_18891,N_18271,N_18292);
or U18892 (N_18892,N_18363,N_18251);
or U18893 (N_18893,N_18321,N_18107);
xnor U18894 (N_18894,N_18041,N_18115);
nor U18895 (N_18895,N_18339,N_18414);
or U18896 (N_18896,N_18124,N_18085);
xor U18897 (N_18897,N_18008,N_18117);
and U18898 (N_18898,N_18026,N_18409);
nand U18899 (N_18899,N_18456,N_18553);
and U18900 (N_18900,N_18344,N_18264);
and U18901 (N_18901,N_18191,N_18278);
and U18902 (N_18902,N_18347,N_18134);
and U18903 (N_18903,N_18071,N_18353);
and U18904 (N_18904,N_18461,N_18003);
and U18905 (N_18905,N_18320,N_18569);
nand U18906 (N_18906,N_18439,N_18047);
and U18907 (N_18907,N_18485,N_18075);
nor U18908 (N_18908,N_18439,N_18453);
nand U18909 (N_18909,N_18344,N_18110);
and U18910 (N_18910,N_18150,N_18055);
nand U18911 (N_18911,N_18451,N_18544);
nor U18912 (N_18912,N_18365,N_18574);
nor U18913 (N_18913,N_18051,N_18252);
nand U18914 (N_18914,N_18020,N_18478);
nor U18915 (N_18915,N_18441,N_18008);
nand U18916 (N_18916,N_18224,N_18018);
nand U18917 (N_18917,N_18589,N_18477);
nor U18918 (N_18918,N_18364,N_18264);
nand U18919 (N_18919,N_18582,N_18369);
and U18920 (N_18920,N_18003,N_18193);
xor U18921 (N_18921,N_18355,N_18359);
and U18922 (N_18922,N_18508,N_18524);
nor U18923 (N_18923,N_18388,N_18540);
or U18924 (N_18924,N_18502,N_18063);
nand U18925 (N_18925,N_18548,N_18238);
or U18926 (N_18926,N_18208,N_18410);
and U18927 (N_18927,N_18500,N_18212);
and U18928 (N_18928,N_18466,N_18389);
or U18929 (N_18929,N_18343,N_18404);
nor U18930 (N_18930,N_18221,N_18174);
or U18931 (N_18931,N_18557,N_18108);
nand U18932 (N_18932,N_18446,N_18187);
nor U18933 (N_18933,N_18359,N_18249);
xor U18934 (N_18934,N_18381,N_18569);
and U18935 (N_18935,N_18359,N_18357);
nor U18936 (N_18936,N_18193,N_18112);
and U18937 (N_18937,N_18559,N_18383);
xnor U18938 (N_18938,N_18338,N_18350);
xnor U18939 (N_18939,N_18570,N_18400);
nor U18940 (N_18940,N_18485,N_18105);
and U18941 (N_18941,N_18111,N_18391);
nand U18942 (N_18942,N_18343,N_18597);
nand U18943 (N_18943,N_18483,N_18460);
or U18944 (N_18944,N_18312,N_18334);
and U18945 (N_18945,N_18242,N_18049);
and U18946 (N_18946,N_18200,N_18277);
or U18947 (N_18947,N_18325,N_18541);
and U18948 (N_18948,N_18306,N_18118);
xnor U18949 (N_18949,N_18479,N_18280);
or U18950 (N_18950,N_18015,N_18481);
or U18951 (N_18951,N_18514,N_18399);
or U18952 (N_18952,N_18141,N_18096);
and U18953 (N_18953,N_18487,N_18370);
nor U18954 (N_18954,N_18524,N_18248);
nand U18955 (N_18955,N_18525,N_18517);
and U18956 (N_18956,N_18347,N_18145);
or U18957 (N_18957,N_18318,N_18225);
and U18958 (N_18958,N_18345,N_18504);
and U18959 (N_18959,N_18077,N_18520);
nor U18960 (N_18960,N_18312,N_18540);
and U18961 (N_18961,N_18092,N_18075);
and U18962 (N_18962,N_18230,N_18350);
or U18963 (N_18963,N_18105,N_18150);
and U18964 (N_18964,N_18284,N_18054);
or U18965 (N_18965,N_18540,N_18356);
nor U18966 (N_18966,N_18201,N_18463);
xnor U18967 (N_18967,N_18427,N_18599);
xnor U18968 (N_18968,N_18416,N_18213);
xnor U18969 (N_18969,N_18496,N_18272);
and U18970 (N_18970,N_18000,N_18105);
nand U18971 (N_18971,N_18105,N_18209);
nand U18972 (N_18972,N_18477,N_18326);
nor U18973 (N_18973,N_18153,N_18435);
nand U18974 (N_18974,N_18426,N_18162);
nand U18975 (N_18975,N_18565,N_18163);
nand U18976 (N_18976,N_18001,N_18035);
nand U18977 (N_18977,N_18103,N_18543);
nand U18978 (N_18978,N_18458,N_18030);
nor U18979 (N_18979,N_18584,N_18204);
and U18980 (N_18980,N_18333,N_18052);
xnor U18981 (N_18981,N_18352,N_18364);
or U18982 (N_18982,N_18570,N_18317);
and U18983 (N_18983,N_18394,N_18586);
nand U18984 (N_18984,N_18385,N_18033);
xor U18985 (N_18985,N_18127,N_18303);
and U18986 (N_18986,N_18442,N_18409);
and U18987 (N_18987,N_18347,N_18344);
nand U18988 (N_18988,N_18190,N_18103);
xor U18989 (N_18989,N_18240,N_18172);
xnor U18990 (N_18990,N_18010,N_18101);
xnor U18991 (N_18991,N_18195,N_18296);
xnor U18992 (N_18992,N_18551,N_18437);
or U18993 (N_18993,N_18555,N_18585);
xnor U18994 (N_18994,N_18082,N_18166);
or U18995 (N_18995,N_18461,N_18189);
or U18996 (N_18996,N_18319,N_18156);
and U18997 (N_18997,N_18309,N_18561);
and U18998 (N_18998,N_18293,N_18570);
xnor U18999 (N_18999,N_18175,N_18067);
or U19000 (N_19000,N_18103,N_18281);
or U19001 (N_19001,N_18216,N_18270);
and U19002 (N_19002,N_18528,N_18442);
nand U19003 (N_19003,N_18586,N_18100);
nor U19004 (N_19004,N_18226,N_18414);
or U19005 (N_19005,N_18170,N_18194);
xor U19006 (N_19006,N_18291,N_18585);
and U19007 (N_19007,N_18401,N_18173);
xnor U19008 (N_19008,N_18121,N_18162);
nand U19009 (N_19009,N_18169,N_18141);
nand U19010 (N_19010,N_18171,N_18521);
and U19011 (N_19011,N_18416,N_18382);
nand U19012 (N_19012,N_18523,N_18252);
or U19013 (N_19013,N_18029,N_18062);
nor U19014 (N_19014,N_18269,N_18507);
or U19015 (N_19015,N_18165,N_18429);
xor U19016 (N_19016,N_18325,N_18387);
nor U19017 (N_19017,N_18484,N_18066);
or U19018 (N_19018,N_18063,N_18436);
nor U19019 (N_19019,N_18285,N_18567);
nand U19020 (N_19020,N_18503,N_18338);
xnor U19021 (N_19021,N_18058,N_18114);
or U19022 (N_19022,N_18046,N_18584);
nand U19023 (N_19023,N_18454,N_18591);
nor U19024 (N_19024,N_18527,N_18219);
xnor U19025 (N_19025,N_18407,N_18022);
xnor U19026 (N_19026,N_18376,N_18476);
nor U19027 (N_19027,N_18539,N_18470);
xnor U19028 (N_19028,N_18588,N_18343);
or U19029 (N_19029,N_18499,N_18194);
xor U19030 (N_19030,N_18295,N_18134);
xor U19031 (N_19031,N_18045,N_18536);
nor U19032 (N_19032,N_18513,N_18255);
xor U19033 (N_19033,N_18438,N_18493);
nor U19034 (N_19034,N_18314,N_18165);
nand U19035 (N_19035,N_18444,N_18388);
xor U19036 (N_19036,N_18122,N_18532);
nor U19037 (N_19037,N_18517,N_18221);
xor U19038 (N_19038,N_18374,N_18303);
and U19039 (N_19039,N_18318,N_18284);
nor U19040 (N_19040,N_18590,N_18027);
xor U19041 (N_19041,N_18571,N_18503);
or U19042 (N_19042,N_18243,N_18144);
or U19043 (N_19043,N_18201,N_18255);
and U19044 (N_19044,N_18191,N_18480);
or U19045 (N_19045,N_18110,N_18460);
nor U19046 (N_19046,N_18035,N_18595);
and U19047 (N_19047,N_18256,N_18217);
xnor U19048 (N_19048,N_18120,N_18314);
or U19049 (N_19049,N_18259,N_18267);
xor U19050 (N_19050,N_18519,N_18075);
or U19051 (N_19051,N_18598,N_18278);
or U19052 (N_19052,N_18502,N_18189);
nor U19053 (N_19053,N_18568,N_18483);
nand U19054 (N_19054,N_18286,N_18191);
or U19055 (N_19055,N_18143,N_18296);
nand U19056 (N_19056,N_18456,N_18182);
nor U19057 (N_19057,N_18296,N_18339);
nor U19058 (N_19058,N_18180,N_18495);
or U19059 (N_19059,N_18261,N_18322);
and U19060 (N_19060,N_18316,N_18324);
or U19061 (N_19061,N_18394,N_18074);
nor U19062 (N_19062,N_18380,N_18567);
or U19063 (N_19063,N_18418,N_18285);
and U19064 (N_19064,N_18524,N_18416);
xor U19065 (N_19065,N_18123,N_18053);
nand U19066 (N_19066,N_18277,N_18183);
or U19067 (N_19067,N_18395,N_18246);
and U19068 (N_19068,N_18303,N_18491);
nor U19069 (N_19069,N_18546,N_18447);
nand U19070 (N_19070,N_18198,N_18544);
or U19071 (N_19071,N_18558,N_18354);
or U19072 (N_19072,N_18090,N_18563);
or U19073 (N_19073,N_18150,N_18044);
nor U19074 (N_19074,N_18501,N_18476);
and U19075 (N_19075,N_18544,N_18598);
or U19076 (N_19076,N_18401,N_18471);
nand U19077 (N_19077,N_18019,N_18145);
xnor U19078 (N_19078,N_18196,N_18248);
nor U19079 (N_19079,N_18187,N_18111);
or U19080 (N_19080,N_18336,N_18161);
xor U19081 (N_19081,N_18556,N_18562);
and U19082 (N_19082,N_18304,N_18475);
xnor U19083 (N_19083,N_18098,N_18408);
and U19084 (N_19084,N_18261,N_18364);
nand U19085 (N_19085,N_18177,N_18473);
nand U19086 (N_19086,N_18278,N_18244);
xor U19087 (N_19087,N_18086,N_18122);
xnor U19088 (N_19088,N_18555,N_18533);
xor U19089 (N_19089,N_18120,N_18377);
xnor U19090 (N_19090,N_18519,N_18165);
nor U19091 (N_19091,N_18222,N_18571);
xor U19092 (N_19092,N_18292,N_18463);
nand U19093 (N_19093,N_18322,N_18027);
nor U19094 (N_19094,N_18373,N_18340);
nand U19095 (N_19095,N_18122,N_18339);
or U19096 (N_19096,N_18155,N_18572);
nand U19097 (N_19097,N_18249,N_18244);
and U19098 (N_19098,N_18567,N_18572);
nor U19099 (N_19099,N_18362,N_18003);
nor U19100 (N_19100,N_18290,N_18493);
or U19101 (N_19101,N_18545,N_18572);
nand U19102 (N_19102,N_18334,N_18577);
or U19103 (N_19103,N_18168,N_18039);
xor U19104 (N_19104,N_18517,N_18381);
nor U19105 (N_19105,N_18588,N_18288);
xor U19106 (N_19106,N_18157,N_18074);
nand U19107 (N_19107,N_18391,N_18055);
nand U19108 (N_19108,N_18290,N_18266);
nand U19109 (N_19109,N_18532,N_18062);
xnor U19110 (N_19110,N_18521,N_18467);
and U19111 (N_19111,N_18595,N_18274);
nor U19112 (N_19112,N_18276,N_18254);
or U19113 (N_19113,N_18111,N_18491);
nor U19114 (N_19114,N_18093,N_18071);
nor U19115 (N_19115,N_18198,N_18156);
nor U19116 (N_19116,N_18442,N_18349);
and U19117 (N_19117,N_18050,N_18041);
and U19118 (N_19118,N_18557,N_18526);
nor U19119 (N_19119,N_18121,N_18198);
nor U19120 (N_19120,N_18222,N_18581);
or U19121 (N_19121,N_18438,N_18027);
and U19122 (N_19122,N_18100,N_18398);
xnor U19123 (N_19123,N_18262,N_18391);
and U19124 (N_19124,N_18235,N_18341);
or U19125 (N_19125,N_18026,N_18565);
nor U19126 (N_19126,N_18048,N_18497);
nor U19127 (N_19127,N_18468,N_18061);
xnor U19128 (N_19128,N_18271,N_18016);
xnor U19129 (N_19129,N_18053,N_18581);
and U19130 (N_19130,N_18094,N_18118);
nand U19131 (N_19131,N_18161,N_18588);
nor U19132 (N_19132,N_18408,N_18293);
nor U19133 (N_19133,N_18215,N_18597);
nor U19134 (N_19134,N_18590,N_18243);
nor U19135 (N_19135,N_18180,N_18471);
nor U19136 (N_19136,N_18516,N_18019);
xnor U19137 (N_19137,N_18378,N_18092);
or U19138 (N_19138,N_18249,N_18111);
nor U19139 (N_19139,N_18019,N_18039);
nand U19140 (N_19140,N_18314,N_18249);
nand U19141 (N_19141,N_18087,N_18398);
nor U19142 (N_19142,N_18017,N_18200);
or U19143 (N_19143,N_18133,N_18593);
or U19144 (N_19144,N_18033,N_18218);
xor U19145 (N_19145,N_18273,N_18475);
or U19146 (N_19146,N_18438,N_18486);
xor U19147 (N_19147,N_18157,N_18318);
and U19148 (N_19148,N_18574,N_18147);
and U19149 (N_19149,N_18051,N_18538);
or U19150 (N_19150,N_18555,N_18160);
nor U19151 (N_19151,N_18594,N_18191);
nand U19152 (N_19152,N_18501,N_18368);
or U19153 (N_19153,N_18117,N_18422);
and U19154 (N_19154,N_18150,N_18378);
nand U19155 (N_19155,N_18447,N_18536);
or U19156 (N_19156,N_18480,N_18179);
and U19157 (N_19157,N_18102,N_18533);
or U19158 (N_19158,N_18277,N_18336);
and U19159 (N_19159,N_18557,N_18003);
or U19160 (N_19160,N_18270,N_18200);
and U19161 (N_19161,N_18548,N_18497);
xnor U19162 (N_19162,N_18469,N_18161);
xor U19163 (N_19163,N_18475,N_18266);
or U19164 (N_19164,N_18080,N_18575);
nand U19165 (N_19165,N_18074,N_18355);
nor U19166 (N_19166,N_18155,N_18394);
nor U19167 (N_19167,N_18005,N_18359);
xnor U19168 (N_19168,N_18123,N_18362);
xnor U19169 (N_19169,N_18447,N_18252);
or U19170 (N_19170,N_18138,N_18307);
or U19171 (N_19171,N_18499,N_18314);
nor U19172 (N_19172,N_18207,N_18586);
xor U19173 (N_19173,N_18481,N_18466);
and U19174 (N_19174,N_18185,N_18389);
xor U19175 (N_19175,N_18311,N_18264);
xor U19176 (N_19176,N_18348,N_18039);
nor U19177 (N_19177,N_18426,N_18535);
nor U19178 (N_19178,N_18022,N_18220);
and U19179 (N_19179,N_18598,N_18526);
xnor U19180 (N_19180,N_18250,N_18151);
nand U19181 (N_19181,N_18186,N_18086);
xor U19182 (N_19182,N_18511,N_18018);
xnor U19183 (N_19183,N_18168,N_18110);
nor U19184 (N_19184,N_18011,N_18099);
nor U19185 (N_19185,N_18262,N_18008);
xnor U19186 (N_19186,N_18016,N_18061);
or U19187 (N_19187,N_18445,N_18237);
nand U19188 (N_19188,N_18349,N_18286);
nor U19189 (N_19189,N_18135,N_18496);
xnor U19190 (N_19190,N_18577,N_18119);
nor U19191 (N_19191,N_18238,N_18253);
nor U19192 (N_19192,N_18101,N_18395);
or U19193 (N_19193,N_18252,N_18028);
or U19194 (N_19194,N_18084,N_18419);
and U19195 (N_19195,N_18572,N_18059);
nand U19196 (N_19196,N_18404,N_18455);
or U19197 (N_19197,N_18010,N_18550);
xor U19198 (N_19198,N_18192,N_18551);
or U19199 (N_19199,N_18266,N_18131);
and U19200 (N_19200,N_19050,N_18998);
xor U19201 (N_19201,N_18959,N_18688);
nor U19202 (N_19202,N_18610,N_19041);
and U19203 (N_19203,N_18710,N_18720);
nand U19204 (N_19204,N_19018,N_19065);
nor U19205 (N_19205,N_18616,N_19022);
nand U19206 (N_19206,N_18747,N_18807);
or U19207 (N_19207,N_18672,N_19043);
or U19208 (N_19208,N_19006,N_19099);
nor U19209 (N_19209,N_19167,N_18728);
nor U19210 (N_19210,N_19100,N_18966);
nor U19211 (N_19211,N_18676,N_19111);
nor U19212 (N_19212,N_19097,N_18945);
and U19213 (N_19213,N_18934,N_18729);
nand U19214 (N_19214,N_19117,N_18857);
and U19215 (N_19215,N_18699,N_19148);
and U19216 (N_19216,N_18772,N_18844);
and U19217 (N_19217,N_18642,N_18768);
xnor U19218 (N_19218,N_18798,N_18647);
nand U19219 (N_19219,N_19095,N_18939);
xor U19220 (N_19220,N_18816,N_19162);
nor U19221 (N_19221,N_18948,N_18872);
and U19222 (N_19222,N_18722,N_19102);
nand U19223 (N_19223,N_18740,N_19092);
nor U19224 (N_19224,N_19136,N_18810);
xor U19225 (N_19225,N_18894,N_18875);
and U19226 (N_19226,N_18916,N_18615);
and U19227 (N_19227,N_18895,N_19188);
xor U19228 (N_19228,N_18759,N_18848);
xnor U19229 (N_19229,N_18698,N_19123);
xor U19230 (N_19230,N_18755,N_19048);
nand U19231 (N_19231,N_18629,N_19121);
nand U19232 (N_19232,N_18746,N_18622);
nand U19233 (N_19233,N_18835,N_18985);
and U19234 (N_19234,N_19032,N_18803);
nor U19235 (N_19235,N_19197,N_19016);
nor U19236 (N_19236,N_18712,N_19187);
and U19237 (N_19237,N_18708,N_19130);
and U19238 (N_19238,N_18602,N_18984);
nand U19239 (N_19239,N_18704,N_19154);
nor U19240 (N_19240,N_18987,N_18797);
nor U19241 (N_19241,N_18983,N_19038);
nand U19242 (N_19242,N_18656,N_18785);
or U19243 (N_19243,N_19008,N_18689);
or U19244 (N_19244,N_18600,N_18748);
xnor U19245 (N_19245,N_18653,N_18972);
nor U19246 (N_19246,N_19066,N_18936);
nor U19247 (N_19247,N_19172,N_19047);
xor U19248 (N_19248,N_18633,N_18905);
or U19249 (N_19249,N_18717,N_18873);
or U19250 (N_19250,N_19035,N_18626);
nand U19251 (N_19251,N_18751,N_18639);
nand U19252 (N_19252,N_18684,N_18775);
xor U19253 (N_19253,N_19107,N_18767);
nor U19254 (N_19254,N_18809,N_18766);
and U19255 (N_19255,N_18737,N_19078);
xnor U19256 (N_19256,N_18881,N_18799);
or U19257 (N_19257,N_19103,N_18837);
or U19258 (N_19258,N_18938,N_18765);
nand U19259 (N_19259,N_19105,N_19104);
or U19260 (N_19260,N_19181,N_18643);
xnor U19261 (N_19261,N_18757,N_18743);
and U19262 (N_19262,N_19039,N_18679);
nor U19263 (N_19263,N_18625,N_18957);
nand U19264 (N_19264,N_18804,N_18820);
xor U19265 (N_19265,N_19151,N_18640);
or U19266 (N_19266,N_19005,N_18665);
nor U19267 (N_19267,N_18999,N_19182);
or U19268 (N_19268,N_18904,N_18861);
or U19269 (N_19269,N_18669,N_18635);
or U19270 (N_19270,N_18659,N_19176);
nor U19271 (N_19271,N_19033,N_18780);
nor U19272 (N_19272,N_18836,N_18661);
xor U19273 (N_19273,N_19169,N_18801);
or U19274 (N_19274,N_19115,N_18877);
xor U19275 (N_19275,N_18947,N_18833);
or U19276 (N_19276,N_18986,N_18893);
xor U19277 (N_19277,N_18822,N_18874);
xor U19278 (N_19278,N_19088,N_18982);
or U19279 (N_19279,N_19090,N_19113);
nand U19280 (N_19280,N_18745,N_19158);
xnor U19281 (N_19281,N_18879,N_19046);
xor U19282 (N_19282,N_19164,N_19067);
or U19283 (N_19283,N_18834,N_19037);
nand U19284 (N_19284,N_18750,N_19080);
nor U19285 (N_19285,N_18968,N_18981);
or U19286 (N_19286,N_18702,N_18738);
nor U19287 (N_19287,N_19119,N_18670);
or U19288 (N_19288,N_19076,N_18891);
xor U19289 (N_19289,N_18830,N_18707);
xor U19290 (N_19290,N_19152,N_18946);
nand U19291 (N_19291,N_18620,N_19146);
xor U19292 (N_19292,N_18989,N_18652);
xor U19293 (N_19293,N_19021,N_18869);
nor U19294 (N_19294,N_18693,N_18863);
and U19295 (N_19295,N_19185,N_18988);
xor U19296 (N_19296,N_18865,N_18858);
or U19297 (N_19297,N_18763,N_18645);
nor U19298 (N_19298,N_18923,N_18695);
or U19299 (N_19299,N_18995,N_18903);
xor U19300 (N_19300,N_18931,N_19009);
nor U19301 (N_19301,N_18828,N_19083);
nand U19302 (N_19302,N_19174,N_19141);
nand U19303 (N_19303,N_18992,N_18974);
and U19304 (N_19304,N_18976,N_18808);
and U19305 (N_19305,N_18641,N_18686);
or U19306 (N_19306,N_18912,N_18673);
xnor U19307 (N_19307,N_19196,N_18680);
nor U19308 (N_19308,N_18624,N_19007);
and U19309 (N_19309,N_19085,N_19135);
nand U19310 (N_19310,N_18927,N_18827);
nor U19311 (N_19311,N_18812,N_18787);
nand U19312 (N_19312,N_18734,N_19000);
and U19313 (N_19313,N_18818,N_18733);
xor U19314 (N_19314,N_18762,N_18648);
xor U19315 (N_19315,N_18991,N_18721);
nand U19316 (N_19316,N_18847,N_19057);
or U19317 (N_19317,N_19068,N_18941);
xnor U19318 (N_19318,N_18978,N_19064);
xnor U19319 (N_19319,N_18663,N_18849);
and U19320 (N_19320,N_19098,N_18630);
and U19321 (N_19321,N_18897,N_18632);
nor U19322 (N_19322,N_19109,N_18609);
nand U19323 (N_19323,N_18921,N_18860);
nand U19324 (N_19324,N_18918,N_18681);
nand U19325 (N_19325,N_19144,N_18853);
xnor U19326 (N_19326,N_19186,N_18691);
and U19327 (N_19327,N_18782,N_18924);
nand U19328 (N_19328,N_18650,N_19096);
xor U19329 (N_19329,N_18842,N_19044);
nand U19330 (N_19330,N_19153,N_19110);
and U19331 (N_19331,N_18614,N_19142);
xnor U19332 (N_19332,N_19051,N_18962);
or U19333 (N_19333,N_19063,N_18658);
nand U19334 (N_19334,N_18783,N_18973);
and U19335 (N_19335,N_19112,N_18971);
or U19336 (N_19336,N_19194,N_19086);
nand U19337 (N_19337,N_18711,N_18727);
and U19338 (N_19338,N_19101,N_18876);
and U19339 (N_19339,N_19093,N_19177);
and U19340 (N_19340,N_19161,N_18651);
nand U19341 (N_19341,N_18928,N_19053);
nor U19342 (N_19342,N_18845,N_18664);
or U19343 (N_19343,N_19091,N_18649);
or U19344 (N_19344,N_18674,N_18926);
and U19345 (N_19345,N_18714,N_19191);
nor U19346 (N_19346,N_18718,N_18890);
and U19347 (N_19347,N_18880,N_18898);
and U19348 (N_19348,N_19155,N_18975);
or U19349 (N_19349,N_18675,N_18900);
nand U19350 (N_19350,N_18888,N_18823);
nand U19351 (N_19351,N_19012,N_18932);
or U19352 (N_19352,N_19138,N_18843);
nor U19353 (N_19353,N_18942,N_19055);
and U19354 (N_19354,N_18911,N_18949);
and U19355 (N_19355,N_18758,N_18773);
xnor U19356 (N_19356,N_19134,N_19163);
nor U19357 (N_19357,N_18852,N_19143);
nor U19358 (N_19358,N_18952,N_18965);
nor U19359 (N_19359,N_18846,N_19131);
or U19360 (N_19360,N_19133,N_18760);
or U19361 (N_19361,N_18859,N_18646);
nor U19362 (N_19362,N_18940,N_19189);
or U19363 (N_19363,N_18725,N_18781);
nor U19364 (N_19364,N_19079,N_19168);
or U19365 (N_19365,N_19028,N_18901);
and U19366 (N_19366,N_19084,N_18732);
xor U19367 (N_19367,N_19001,N_19140);
xnor U19368 (N_19368,N_18754,N_18944);
xnor U19369 (N_19369,N_18805,N_18613);
nor U19370 (N_19370,N_18950,N_18703);
nor U19371 (N_19371,N_18892,N_19026);
and U19372 (N_19372,N_19193,N_19081);
and U19373 (N_19373,N_19015,N_18933);
or U19374 (N_19374,N_19075,N_18606);
xor U19375 (N_19375,N_18969,N_18997);
xnor U19376 (N_19376,N_18779,N_19198);
or U19377 (N_19377,N_18790,N_18685);
nor U19378 (N_19378,N_18896,N_18739);
or U19379 (N_19379,N_18716,N_18637);
nand U19380 (N_19380,N_18619,N_18771);
and U19381 (N_19381,N_18603,N_18607);
nor U19382 (N_19382,N_19060,N_18825);
and U19383 (N_19383,N_18899,N_18631);
and U19384 (N_19384,N_19069,N_18761);
nand U19385 (N_19385,N_18902,N_18953);
nor U19386 (N_19386,N_18730,N_18817);
and U19387 (N_19387,N_18819,N_18692);
or U19388 (N_19388,N_19195,N_18870);
xnor U19389 (N_19389,N_19072,N_18851);
and U19390 (N_19390,N_19157,N_18826);
nand U19391 (N_19391,N_19183,N_19118);
or U19392 (N_19392,N_18967,N_18618);
nor U19393 (N_19393,N_18886,N_18735);
and U19394 (N_19394,N_18914,N_18784);
nand U19395 (N_19395,N_19010,N_18829);
and U19396 (N_19396,N_18667,N_18838);
nand U19397 (N_19397,N_18617,N_18638);
nand U19398 (N_19398,N_18937,N_19002);
or U19399 (N_19399,N_18868,N_18655);
nand U19400 (N_19400,N_19027,N_18970);
nand U19401 (N_19401,N_18700,N_18994);
xor U19402 (N_19402,N_19127,N_18697);
nand U19403 (N_19403,N_18910,N_18854);
nand U19404 (N_19404,N_18715,N_18915);
nand U19405 (N_19405,N_19071,N_19052);
or U19406 (N_19406,N_18705,N_19126);
nor U19407 (N_19407,N_19094,N_19025);
or U19408 (N_19408,N_18815,N_18791);
or U19409 (N_19409,N_18884,N_18996);
xnor U19410 (N_19410,N_19054,N_19108);
or U19411 (N_19411,N_18839,N_18832);
nand U19412 (N_19412,N_19190,N_18623);
or U19413 (N_19413,N_18611,N_18954);
xnor U19414 (N_19414,N_19014,N_18668);
or U19415 (N_19415,N_18929,N_18956);
xor U19416 (N_19416,N_19040,N_19173);
nor U19417 (N_19417,N_18883,N_18795);
or U19418 (N_19418,N_19145,N_19034);
or U19419 (N_19419,N_18867,N_18917);
xnor U19420 (N_19420,N_19178,N_19030);
xor U19421 (N_19421,N_19082,N_18964);
or U19422 (N_19422,N_19170,N_18960);
or U19423 (N_19423,N_18789,N_18605);
xnor U19424 (N_19424,N_19129,N_18701);
or U19425 (N_19425,N_18919,N_18908);
xnor U19426 (N_19426,N_18723,N_18612);
nand U19427 (N_19427,N_19124,N_18777);
and U19428 (N_19428,N_19180,N_18811);
nor U19429 (N_19429,N_18906,N_18993);
nand U19430 (N_19430,N_18687,N_18749);
nand U19431 (N_19431,N_18840,N_18706);
xnor U19432 (N_19432,N_18636,N_19159);
nand U19433 (N_19433,N_18621,N_19011);
or U19434 (N_19434,N_19139,N_18864);
nand U19435 (N_19435,N_18608,N_18913);
and U19436 (N_19436,N_18736,N_18980);
xor U19437 (N_19437,N_19087,N_18683);
and U19438 (N_19438,N_19004,N_19049);
nand U19439 (N_19439,N_18634,N_18909);
and U19440 (N_19440,N_19019,N_18713);
or U19441 (N_19441,N_18831,N_18709);
nor U19442 (N_19442,N_19137,N_18802);
and U19443 (N_19443,N_18694,N_19045);
nand U19444 (N_19444,N_18682,N_18770);
xnor U19445 (N_19445,N_18862,N_19042);
nand U19446 (N_19446,N_19165,N_18604);
and U19447 (N_19447,N_19059,N_19120);
nand U19448 (N_19448,N_18690,N_18943);
xnor U19449 (N_19449,N_18814,N_18677);
or U19450 (N_19450,N_18821,N_18601);
nand U19451 (N_19451,N_18741,N_18792);
and U19452 (N_19452,N_18935,N_18990);
nand U19453 (N_19453,N_19147,N_19184);
xor U19454 (N_19454,N_18979,N_18889);
nor U19455 (N_19455,N_18958,N_18788);
nor U19456 (N_19456,N_19132,N_18678);
nand U19457 (N_19457,N_18977,N_18719);
and U19458 (N_19458,N_19128,N_18850);
and U19459 (N_19459,N_18878,N_18866);
nand U19460 (N_19460,N_19171,N_18907);
and U19461 (N_19461,N_19089,N_18724);
and U19462 (N_19462,N_18776,N_19077);
or U19463 (N_19463,N_18753,N_18871);
nor U19464 (N_19464,N_18731,N_19199);
xor U19465 (N_19465,N_18813,N_19031);
xnor U19466 (N_19466,N_18963,N_18726);
and U19467 (N_19467,N_18806,N_18885);
nor U19468 (N_19468,N_18671,N_19150);
nand U19469 (N_19469,N_18627,N_18951);
nand U19470 (N_19470,N_19061,N_19122);
xnor U19471 (N_19471,N_18752,N_18744);
xor U19472 (N_19472,N_18756,N_19125);
nand U19473 (N_19473,N_19003,N_19175);
nor U19474 (N_19474,N_19058,N_18666);
nand U19475 (N_19475,N_19116,N_18824);
xnor U19476 (N_19476,N_19114,N_19179);
nand U19477 (N_19477,N_19020,N_19156);
nand U19478 (N_19478,N_18793,N_18796);
nor U19479 (N_19479,N_18856,N_19106);
nor U19480 (N_19480,N_18794,N_18696);
nand U19481 (N_19481,N_18769,N_18800);
nor U19482 (N_19482,N_18654,N_19160);
or U19483 (N_19483,N_19149,N_18742);
xor U19484 (N_19484,N_18882,N_18855);
and U19485 (N_19485,N_18887,N_18660);
and U19486 (N_19486,N_18961,N_19166);
or U19487 (N_19487,N_19056,N_18662);
nor U19488 (N_19488,N_19029,N_19036);
xor U19489 (N_19489,N_18955,N_18786);
or U19490 (N_19490,N_18657,N_19017);
or U19491 (N_19491,N_19013,N_18644);
and U19492 (N_19492,N_19062,N_18774);
xnor U19493 (N_19493,N_18925,N_18778);
nand U19494 (N_19494,N_19074,N_19024);
and U19495 (N_19495,N_19023,N_19192);
or U19496 (N_19496,N_18764,N_19070);
xnor U19497 (N_19497,N_18922,N_18930);
nand U19498 (N_19498,N_19073,N_18628);
and U19499 (N_19499,N_18841,N_18920);
nor U19500 (N_19500,N_18747,N_18711);
xor U19501 (N_19501,N_18811,N_18951);
nand U19502 (N_19502,N_18807,N_18766);
or U19503 (N_19503,N_19033,N_18749);
or U19504 (N_19504,N_19057,N_18833);
nand U19505 (N_19505,N_18969,N_18755);
or U19506 (N_19506,N_18808,N_19064);
nor U19507 (N_19507,N_18823,N_18790);
and U19508 (N_19508,N_18813,N_18741);
xnor U19509 (N_19509,N_18770,N_18760);
xnor U19510 (N_19510,N_18612,N_18966);
xor U19511 (N_19511,N_18925,N_19103);
or U19512 (N_19512,N_18851,N_18871);
xor U19513 (N_19513,N_18706,N_18618);
and U19514 (N_19514,N_18851,N_18687);
and U19515 (N_19515,N_18751,N_18769);
nand U19516 (N_19516,N_18737,N_19115);
and U19517 (N_19517,N_19042,N_18763);
nand U19518 (N_19518,N_18643,N_19197);
and U19519 (N_19519,N_18993,N_18628);
or U19520 (N_19520,N_18790,N_19199);
nand U19521 (N_19521,N_18754,N_19004);
nor U19522 (N_19522,N_19171,N_18914);
xor U19523 (N_19523,N_19028,N_18712);
xor U19524 (N_19524,N_19142,N_18929);
or U19525 (N_19525,N_18666,N_18613);
nor U19526 (N_19526,N_19068,N_18629);
nand U19527 (N_19527,N_18788,N_18861);
nor U19528 (N_19528,N_18893,N_19068);
nor U19529 (N_19529,N_19111,N_18914);
xnor U19530 (N_19530,N_18876,N_18872);
nor U19531 (N_19531,N_18855,N_18778);
nor U19532 (N_19532,N_18865,N_18843);
nor U19533 (N_19533,N_18822,N_18602);
nor U19534 (N_19534,N_18696,N_18658);
xnor U19535 (N_19535,N_18970,N_18677);
and U19536 (N_19536,N_19179,N_18668);
or U19537 (N_19537,N_18814,N_18994);
nor U19538 (N_19538,N_19045,N_19066);
and U19539 (N_19539,N_19078,N_19133);
or U19540 (N_19540,N_18710,N_18604);
and U19541 (N_19541,N_18667,N_19179);
xnor U19542 (N_19542,N_18896,N_19175);
xnor U19543 (N_19543,N_19087,N_18634);
xor U19544 (N_19544,N_18860,N_18893);
or U19545 (N_19545,N_18932,N_19028);
xor U19546 (N_19546,N_18668,N_18674);
and U19547 (N_19547,N_19173,N_18922);
nand U19548 (N_19548,N_19010,N_18990);
nand U19549 (N_19549,N_18912,N_18795);
nor U19550 (N_19550,N_18937,N_18900);
xor U19551 (N_19551,N_19031,N_19141);
or U19552 (N_19552,N_18914,N_19099);
and U19553 (N_19553,N_19178,N_18744);
or U19554 (N_19554,N_18689,N_18611);
or U19555 (N_19555,N_18712,N_19142);
or U19556 (N_19556,N_18738,N_19088);
nor U19557 (N_19557,N_18773,N_18820);
nor U19558 (N_19558,N_18655,N_18790);
or U19559 (N_19559,N_18836,N_18706);
nor U19560 (N_19560,N_19101,N_19015);
nor U19561 (N_19561,N_18778,N_18672);
xnor U19562 (N_19562,N_18977,N_18729);
or U19563 (N_19563,N_18888,N_18939);
and U19564 (N_19564,N_18664,N_18979);
or U19565 (N_19565,N_19021,N_18836);
nand U19566 (N_19566,N_18769,N_18779);
and U19567 (N_19567,N_18609,N_18726);
xor U19568 (N_19568,N_18934,N_18917);
xor U19569 (N_19569,N_18727,N_18985);
xor U19570 (N_19570,N_18652,N_19177);
xor U19571 (N_19571,N_18644,N_18830);
or U19572 (N_19572,N_19003,N_18712);
xnor U19573 (N_19573,N_18934,N_18624);
nand U19574 (N_19574,N_18919,N_18743);
or U19575 (N_19575,N_18877,N_18842);
nand U19576 (N_19576,N_18889,N_18635);
xor U19577 (N_19577,N_19079,N_18721);
xor U19578 (N_19578,N_19198,N_18869);
nand U19579 (N_19579,N_19076,N_18642);
nor U19580 (N_19580,N_19125,N_18656);
nand U19581 (N_19581,N_18757,N_18885);
nand U19582 (N_19582,N_18922,N_18986);
nand U19583 (N_19583,N_19128,N_18935);
xnor U19584 (N_19584,N_18610,N_18995);
nor U19585 (N_19585,N_19015,N_18817);
nand U19586 (N_19586,N_18624,N_19167);
nand U19587 (N_19587,N_18857,N_18938);
or U19588 (N_19588,N_18780,N_18874);
nor U19589 (N_19589,N_18836,N_19043);
and U19590 (N_19590,N_19112,N_19113);
and U19591 (N_19591,N_18812,N_19133);
xor U19592 (N_19592,N_18982,N_18753);
nand U19593 (N_19593,N_18855,N_18602);
and U19594 (N_19594,N_18748,N_18773);
nand U19595 (N_19595,N_18849,N_19131);
nand U19596 (N_19596,N_18955,N_18669);
xor U19597 (N_19597,N_19025,N_18992);
xnor U19598 (N_19598,N_18999,N_19019);
or U19599 (N_19599,N_18988,N_18853);
and U19600 (N_19600,N_19113,N_19064);
xnor U19601 (N_19601,N_18926,N_18795);
or U19602 (N_19602,N_18767,N_18730);
or U19603 (N_19603,N_18740,N_18756);
xnor U19604 (N_19604,N_18940,N_19130);
xor U19605 (N_19605,N_19073,N_18828);
and U19606 (N_19606,N_18937,N_19064);
xnor U19607 (N_19607,N_19093,N_18901);
nand U19608 (N_19608,N_18647,N_19179);
or U19609 (N_19609,N_18706,N_18799);
or U19610 (N_19610,N_18902,N_18841);
and U19611 (N_19611,N_19037,N_18982);
nor U19612 (N_19612,N_18837,N_19140);
nand U19613 (N_19613,N_19094,N_18763);
nand U19614 (N_19614,N_18940,N_18891);
and U19615 (N_19615,N_18723,N_18824);
nand U19616 (N_19616,N_18801,N_19127);
nand U19617 (N_19617,N_18978,N_18973);
or U19618 (N_19618,N_19140,N_19065);
nor U19619 (N_19619,N_19020,N_18922);
or U19620 (N_19620,N_19105,N_18675);
and U19621 (N_19621,N_18725,N_18647);
xnor U19622 (N_19622,N_18719,N_19125);
xnor U19623 (N_19623,N_18964,N_19007);
or U19624 (N_19624,N_19047,N_18610);
or U19625 (N_19625,N_19179,N_19076);
xnor U19626 (N_19626,N_18701,N_18901);
nand U19627 (N_19627,N_19199,N_18727);
and U19628 (N_19628,N_18673,N_18855);
xor U19629 (N_19629,N_19009,N_19040);
or U19630 (N_19630,N_18617,N_19035);
nor U19631 (N_19631,N_19171,N_18949);
and U19632 (N_19632,N_19169,N_18743);
xor U19633 (N_19633,N_18906,N_18650);
and U19634 (N_19634,N_18624,N_18998);
or U19635 (N_19635,N_18892,N_19082);
nor U19636 (N_19636,N_19100,N_18887);
or U19637 (N_19637,N_19115,N_19037);
and U19638 (N_19638,N_19132,N_19117);
xnor U19639 (N_19639,N_18883,N_18904);
or U19640 (N_19640,N_19192,N_18696);
xor U19641 (N_19641,N_18999,N_18760);
xor U19642 (N_19642,N_18878,N_18879);
nand U19643 (N_19643,N_19155,N_18981);
xor U19644 (N_19644,N_18883,N_18778);
or U19645 (N_19645,N_18805,N_18811);
and U19646 (N_19646,N_18797,N_18768);
or U19647 (N_19647,N_19121,N_18793);
or U19648 (N_19648,N_19150,N_18635);
nor U19649 (N_19649,N_18956,N_19107);
and U19650 (N_19650,N_19043,N_18710);
nor U19651 (N_19651,N_19002,N_19155);
nor U19652 (N_19652,N_18844,N_18780);
xnor U19653 (N_19653,N_19035,N_18817);
nand U19654 (N_19654,N_18729,N_18804);
nand U19655 (N_19655,N_18768,N_18953);
nor U19656 (N_19656,N_19010,N_18959);
or U19657 (N_19657,N_18614,N_18796);
and U19658 (N_19658,N_18996,N_18769);
nor U19659 (N_19659,N_19139,N_18678);
nand U19660 (N_19660,N_18943,N_19056);
and U19661 (N_19661,N_19101,N_18635);
nand U19662 (N_19662,N_19007,N_18650);
xor U19663 (N_19663,N_18642,N_18829);
or U19664 (N_19664,N_18683,N_19037);
or U19665 (N_19665,N_19121,N_19170);
and U19666 (N_19666,N_18882,N_18985);
or U19667 (N_19667,N_18823,N_19058);
or U19668 (N_19668,N_18688,N_19167);
nand U19669 (N_19669,N_18889,N_18672);
nand U19670 (N_19670,N_19010,N_18803);
nand U19671 (N_19671,N_18646,N_18785);
or U19672 (N_19672,N_18635,N_19019);
nand U19673 (N_19673,N_19070,N_18650);
or U19674 (N_19674,N_18854,N_18952);
and U19675 (N_19675,N_18864,N_18701);
nor U19676 (N_19676,N_18882,N_19008);
nand U19677 (N_19677,N_18997,N_18944);
nor U19678 (N_19678,N_18765,N_18679);
nor U19679 (N_19679,N_19103,N_18603);
or U19680 (N_19680,N_19080,N_19114);
or U19681 (N_19681,N_18843,N_18618);
nor U19682 (N_19682,N_18600,N_18977);
xnor U19683 (N_19683,N_18872,N_18673);
or U19684 (N_19684,N_18781,N_18903);
nand U19685 (N_19685,N_18921,N_18930);
nand U19686 (N_19686,N_18916,N_19159);
or U19687 (N_19687,N_19073,N_18724);
nand U19688 (N_19688,N_19008,N_18718);
nand U19689 (N_19689,N_19159,N_18997);
or U19690 (N_19690,N_18824,N_19199);
nor U19691 (N_19691,N_19018,N_19003);
xnor U19692 (N_19692,N_18665,N_18626);
nand U19693 (N_19693,N_19088,N_19057);
or U19694 (N_19694,N_18637,N_19177);
nand U19695 (N_19695,N_18943,N_19160);
nor U19696 (N_19696,N_18899,N_18966);
xnor U19697 (N_19697,N_18913,N_19153);
and U19698 (N_19698,N_19112,N_19189);
and U19699 (N_19699,N_18755,N_18771);
xnor U19700 (N_19700,N_18770,N_19194);
nor U19701 (N_19701,N_19160,N_18800);
or U19702 (N_19702,N_18768,N_18705);
or U19703 (N_19703,N_19020,N_18939);
nor U19704 (N_19704,N_18627,N_18821);
nand U19705 (N_19705,N_18882,N_18960);
nand U19706 (N_19706,N_18882,N_18776);
and U19707 (N_19707,N_18603,N_19047);
nand U19708 (N_19708,N_18910,N_19111);
nor U19709 (N_19709,N_18605,N_18613);
nand U19710 (N_19710,N_19115,N_19157);
nand U19711 (N_19711,N_19166,N_18730);
xnor U19712 (N_19712,N_19110,N_18789);
xnor U19713 (N_19713,N_18872,N_18672);
nand U19714 (N_19714,N_19105,N_18966);
nand U19715 (N_19715,N_18805,N_18827);
and U19716 (N_19716,N_18694,N_18897);
nor U19717 (N_19717,N_18955,N_18993);
nor U19718 (N_19718,N_18733,N_18784);
nor U19719 (N_19719,N_18883,N_18678);
nor U19720 (N_19720,N_18657,N_19157);
xnor U19721 (N_19721,N_18930,N_18854);
xnor U19722 (N_19722,N_18627,N_18769);
xnor U19723 (N_19723,N_18912,N_19159);
xnor U19724 (N_19724,N_19106,N_18661);
xnor U19725 (N_19725,N_18763,N_18766);
xor U19726 (N_19726,N_18744,N_18644);
or U19727 (N_19727,N_18855,N_19151);
xnor U19728 (N_19728,N_18910,N_18770);
xnor U19729 (N_19729,N_18938,N_18769);
and U19730 (N_19730,N_19120,N_19134);
nand U19731 (N_19731,N_18638,N_18671);
and U19732 (N_19732,N_18774,N_18645);
and U19733 (N_19733,N_18789,N_18617);
or U19734 (N_19734,N_19161,N_18798);
nor U19735 (N_19735,N_18722,N_19155);
or U19736 (N_19736,N_19080,N_18980);
nor U19737 (N_19737,N_19050,N_19180);
nor U19738 (N_19738,N_19034,N_18922);
nor U19739 (N_19739,N_18839,N_19066);
nand U19740 (N_19740,N_18916,N_18831);
nand U19741 (N_19741,N_18967,N_19151);
or U19742 (N_19742,N_19007,N_18812);
or U19743 (N_19743,N_19179,N_19083);
nand U19744 (N_19744,N_18618,N_18960);
xor U19745 (N_19745,N_19122,N_18696);
or U19746 (N_19746,N_18719,N_18822);
nand U19747 (N_19747,N_18649,N_18896);
xnor U19748 (N_19748,N_18709,N_18992);
xor U19749 (N_19749,N_18772,N_18889);
nand U19750 (N_19750,N_18759,N_18752);
xnor U19751 (N_19751,N_19120,N_18924);
and U19752 (N_19752,N_19197,N_19185);
xor U19753 (N_19753,N_19085,N_18600);
nand U19754 (N_19754,N_19175,N_19109);
nand U19755 (N_19755,N_19158,N_19110);
xnor U19756 (N_19756,N_19109,N_18619);
nor U19757 (N_19757,N_18899,N_19145);
and U19758 (N_19758,N_18741,N_18830);
and U19759 (N_19759,N_18627,N_19187);
or U19760 (N_19760,N_18610,N_18713);
and U19761 (N_19761,N_19186,N_19035);
nand U19762 (N_19762,N_18712,N_18631);
or U19763 (N_19763,N_18971,N_18703);
and U19764 (N_19764,N_18891,N_19188);
xor U19765 (N_19765,N_18753,N_18751);
xor U19766 (N_19766,N_19104,N_19029);
or U19767 (N_19767,N_18847,N_19072);
or U19768 (N_19768,N_18642,N_19001);
or U19769 (N_19769,N_18967,N_18770);
nor U19770 (N_19770,N_18656,N_18725);
nor U19771 (N_19771,N_18961,N_19141);
or U19772 (N_19772,N_18604,N_18745);
nand U19773 (N_19773,N_19032,N_19031);
xor U19774 (N_19774,N_19057,N_18808);
xor U19775 (N_19775,N_18723,N_18736);
xor U19776 (N_19776,N_18826,N_19001);
or U19777 (N_19777,N_19180,N_18818);
nor U19778 (N_19778,N_18796,N_18907);
or U19779 (N_19779,N_18931,N_18933);
and U19780 (N_19780,N_18629,N_18823);
or U19781 (N_19781,N_18696,N_18934);
or U19782 (N_19782,N_18909,N_18677);
xor U19783 (N_19783,N_19076,N_19021);
and U19784 (N_19784,N_18808,N_18861);
and U19785 (N_19785,N_18796,N_18809);
or U19786 (N_19786,N_19173,N_18971);
xor U19787 (N_19787,N_18806,N_19152);
nand U19788 (N_19788,N_19120,N_18913);
nand U19789 (N_19789,N_18652,N_19120);
xor U19790 (N_19790,N_18697,N_18982);
or U19791 (N_19791,N_19078,N_19052);
and U19792 (N_19792,N_19011,N_18741);
or U19793 (N_19793,N_19043,N_18972);
and U19794 (N_19794,N_18897,N_18642);
nand U19795 (N_19795,N_18758,N_18606);
or U19796 (N_19796,N_18644,N_18783);
nor U19797 (N_19797,N_18904,N_18689);
nor U19798 (N_19798,N_19128,N_19122);
nand U19799 (N_19799,N_19029,N_19001);
or U19800 (N_19800,N_19713,N_19403);
nand U19801 (N_19801,N_19383,N_19491);
or U19802 (N_19802,N_19729,N_19231);
nor U19803 (N_19803,N_19679,N_19634);
or U19804 (N_19804,N_19688,N_19718);
nand U19805 (N_19805,N_19682,N_19340);
xnor U19806 (N_19806,N_19237,N_19702);
xor U19807 (N_19807,N_19677,N_19609);
and U19808 (N_19808,N_19648,N_19370);
nand U19809 (N_19809,N_19304,N_19243);
and U19810 (N_19810,N_19664,N_19581);
nor U19811 (N_19811,N_19326,N_19208);
and U19812 (N_19812,N_19375,N_19396);
nand U19813 (N_19813,N_19350,N_19201);
nor U19814 (N_19814,N_19267,N_19500);
xor U19815 (N_19815,N_19797,N_19235);
xnor U19816 (N_19816,N_19446,N_19359);
nand U19817 (N_19817,N_19552,N_19458);
and U19818 (N_19818,N_19335,N_19788);
nor U19819 (N_19819,N_19625,N_19590);
xnor U19820 (N_19820,N_19752,N_19269);
nand U19821 (N_19821,N_19381,N_19576);
and U19822 (N_19822,N_19541,N_19731);
and U19823 (N_19823,N_19654,N_19285);
and U19824 (N_19824,N_19268,N_19447);
nand U19825 (N_19825,N_19344,N_19621);
nand U19826 (N_19826,N_19532,N_19308);
and U19827 (N_19827,N_19264,N_19619);
or U19828 (N_19828,N_19583,N_19436);
or U19829 (N_19829,N_19617,N_19368);
or U19830 (N_19830,N_19706,N_19596);
xor U19831 (N_19831,N_19493,N_19555);
or U19832 (N_19832,N_19780,N_19223);
nor U19833 (N_19833,N_19227,N_19736);
and U19834 (N_19834,N_19572,N_19672);
and U19835 (N_19835,N_19431,N_19520);
nand U19836 (N_19836,N_19354,N_19464);
and U19837 (N_19837,N_19506,N_19412);
xnor U19838 (N_19838,N_19781,N_19758);
nor U19839 (N_19839,N_19507,N_19275);
nor U19840 (N_19840,N_19761,N_19579);
or U19841 (N_19841,N_19616,N_19360);
nor U19842 (N_19842,N_19330,N_19432);
or U19843 (N_19843,N_19252,N_19485);
nand U19844 (N_19844,N_19347,N_19787);
or U19845 (N_19845,N_19380,N_19647);
nor U19846 (N_19846,N_19349,N_19577);
xor U19847 (N_19847,N_19321,N_19454);
and U19848 (N_19848,N_19624,N_19795);
xnor U19849 (N_19849,N_19226,N_19741);
or U19850 (N_19850,N_19734,N_19336);
or U19851 (N_19851,N_19589,N_19261);
nand U19852 (N_19852,N_19723,N_19700);
xor U19853 (N_19853,N_19440,N_19641);
nor U19854 (N_19854,N_19292,N_19525);
nor U19855 (N_19855,N_19317,N_19694);
xor U19856 (N_19856,N_19470,N_19385);
nor U19857 (N_19857,N_19435,N_19288);
or U19858 (N_19858,N_19279,N_19662);
nand U19859 (N_19859,N_19659,N_19676);
nand U19860 (N_19860,N_19778,N_19430);
or U19861 (N_19861,N_19759,N_19508);
xor U19862 (N_19862,N_19523,N_19484);
nor U19863 (N_19863,N_19522,N_19299);
nand U19864 (N_19864,N_19595,N_19324);
or U19865 (N_19865,N_19796,N_19389);
xor U19866 (N_19866,N_19366,N_19627);
nor U19867 (N_19867,N_19241,N_19398);
or U19868 (N_19868,N_19351,N_19737);
or U19869 (N_19869,N_19692,N_19757);
nor U19870 (N_19870,N_19224,N_19730);
and U19871 (N_19871,N_19253,N_19674);
or U19872 (N_19872,N_19450,N_19701);
and U19873 (N_19873,N_19533,N_19559);
nand U19874 (N_19874,N_19206,N_19384);
nand U19875 (N_19875,N_19756,N_19695);
nor U19876 (N_19876,N_19482,N_19281);
nand U19877 (N_19877,N_19260,N_19382);
xnor U19878 (N_19878,N_19521,N_19420);
nor U19879 (N_19879,N_19371,N_19671);
and U19880 (N_19880,N_19418,N_19537);
nor U19881 (N_19881,N_19284,N_19526);
nand U19882 (N_19882,N_19274,N_19417);
or U19883 (N_19883,N_19293,N_19785);
xor U19884 (N_19884,N_19545,N_19301);
nor U19885 (N_19885,N_19428,N_19652);
nand U19886 (N_19886,N_19327,N_19512);
or U19887 (N_19887,N_19710,N_19228);
and U19888 (N_19888,N_19764,N_19789);
nor U19889 (N_19889,N_19610,N_19316);
and U19890 (N_19890,N_19345,N_19578);
or U19891 (N_19891,N_19635,N_19314);
nor U19892 (N_19892,N_19587,N_19691);
xnor U19893 (N_19893,N_19546,N_19471);
xor U19894 (N_19894,N_19580,N_19307);
or U19895 (N_19895,N_19711,N_19423);
nand U19896 (N_19896,N_19518,N_19593);
nand U19897 (N_19897,N_19215,N_19549);
nand U19898 (N_19898,N_19251,N_19755);
xnor U19899 (N_19899,N_19653,N_19209);
and U19900 (N_19900,N_19575,N_19313);
nor U19901 (N_19901,N_19438,N_19277);
nor U19902 (N_19902,N_19643,N_19312);
and U19903 (N_19903,N_19405,N_19468);
or U19904 (N_19904,N_19250,N_19407);
nor U19905 (N_19905,N_19722,N_19282);
nand U19906 (N_19906,N_19232,N_19218);
and U19907 (N_19907,N_19400,N_19727);
nand U19908 (N_19908,N_19735,N_19716);
xor U19909 (N_19909,N_19379,N_19399);
and U19910 (N_19910,N_19239,N_19531);
xnor U19911 (N_19911,N_19510,N_19479);
nor U19912 (N_19912,N_19753,N_19775);
and U19913 (N_19913,N_19358,N_19728);
and U19914 (N_19914,N_19703,N_19406);
and U19915 (N_19915,N_19453,N_19684);
or U19916 (N_19916,N_19513,N_19763);
and U19917 (N_19917,N_19637,N_19465);
and U19918 (N_19918,N_19352,N_19733);
nor U19919 (N_19919,N_19489,N_19568);
xor U19920 (N_19920,N_19517,N_19230);
nor U19921 (N_19921,N_19337,N_19481);
nor U19922 (N_19922,N_19516,N_19649);
nand U19923 (N_19923,N_19540,N_19690);
xor U19924 (N_19924,N_19445,N_19614);
xor U19925 (N_19925,N_19622,N_19615);
nor U19926 (N_19926,N_19698,N_19678);
nor U19927 (N_19927,N_19413,N_19469);
nor U19928 (N_19928,N_19739,N_19318);
or U19929 (N_19929,N_19768,N_19630);
xnor U19930 (N_19930,N_19636,N_19644);
xor U19931 (N_19931,N_19750,N_19426);
nand U19932 (N_19932,N_19202,N_19663);
or U19933 (N_19933,N_19502,N_19628);
nor U19934 (N_19934,N_19501,N_19437);
or U19935 (N_19935,N_19666,N_19488);
or U19936 (N_19936,N_19278,N_19565);
and U19937 (N_19937,N_19592,N_19311);
nand U19938 (N_19938,N_19222,N_19717);
xnor U19939 (N_19939,N_19212,N_19640);
xor U19940 (N_19940,N_19563,N_19234);
or U19941 (N_19941,N_19362,N_19289);
or U19942 (N_19942,N_19490,N_19601);
nand U19943 (N_19943,N_19276,N_19598);
nor U19944 (N_19944,N_19262,N_19325);
nand U19945 (N_19945,N_19242,N_19548);
and U19946 (N_19946,N_19402,N_19509);
nor U19947 (N_19947,N_19642,N_19338);
xnor U19948 (N_19948,N_19594,N_19608);
nor U19949 (N_19949,N_19773,N_19499);
nor U19950 (N_19950,N_19455,N_19320);
nand U19951 (N_19951,N_19602,N_19497);
nor U19952 (N_19952,N_19305,N_19461);
nand U19953 (N_19953,N_19618,N_19708);
xnor U19954 (N_19954,N_19646,N_19794);
and U19955 (N_19955,N_19607,N_19667);
nand U19956 (N_19956,N_19534,N_19689);
nor U19957 (N_19957,N_19254,N_19528);
or U19958 (N_19958,N_19751,N_19462);
nand U19959 (N_19959,N_19342,N_19393);
and U19960 (N_19960,N_19255,N_19777);
xor U19961 (N_19961,N_19505,N_19765);
nand U19962 (N_19962,N_19749,N_19738);
xnor U19963 (N_19963,N_19527,N_19709);
nand U19964 (N_19964,N_19207,N_19632);
nand U19965 (N_19965,N_19422,N_19448);
nor U19966 (N_19966,N_19626,N_19374);
and U19967 (N_19967,N_19770,N_19503);
xor U19968 (N_19968,N_19744,N_19270);
nand U19969 (N_19969,N_19651,N_19638);
or U19970 (N_19970,N_19424,N_19564);
nand U19971 (N_19971,N_19495,N_19460);
nand U19972 (N_19972,N_19558,N_19287);
or U19973 (N_19973,N_19323,N_19556);
and U19974 (N_19974,N_19742,N_19378);
or U19975 (N_19975,N_19771,N_19754);
xnor U19976 (N_19976,N_19233,N_19599);
nand U19977 (N_19977,N_19225,N_19258);
nor U19978 (N_19978,N_19200,N_19762);
nand U19979 (N_19979,N_19514,N_19245);
xnor U19980 (N_19980,N_19585,N_19449);
or U19981 (N_19981,N_19363,N_19259);
nor U19982 (N_19982,N_19786,N_19560);
xnor U19983 (N_19983,N_19566,N_19792);
or U19984 (N_19984,N_19386,N_19570);
or U19985 (N_19985,N_19213,N_19669);
or U19986 (N_19986,N_19515,N_19740);
and U19987 (N_19987,N_19410,N_19743);
and U19988 (N_19988,N_19769,N_19219);
or U19989 (N_19989,N_19249,N_19551);
and U19990 (N_19990,N_19343,N_19790);
nor U19991 (N_19991,N_19720,N_19680);
and U19992 (N_19992,N_19466,N_19726);
nand U19993 (N_19993,N_19256,N_19356);
xnor U19994 (N_19994,N_19273,N_19496);
and U19995 (N_19995,N_19421,N_19395);
or U19996 (N_19996,N_19612,N_19291);
nor U19997 (N_19997,N_19306,N_19456);
and U19998 (N_19998,N_19613,N_19714);
nand U19999 (N_19999,N_19369,N_19332);
and U20000 (N_20000,N_19238,N_19766);
nor U20001 (N_20001,N_19504,N_19645);
nand U20002 (N_20002,N_19220,N_19685);
nor U20003 (N_20003,N_19732,N_19452);
nand U20004 (N_20004,N_19543,N_19429);
or U20005 (N_20005,N_19597,N_19473);
xnor U20006 (N_20006,N_19390,N_19300);
nand U20007 (N_20007,N_19286,N_19524);
nor U20008 (N_20008,N_19433,N_19247);
nand U20009 (N_20009,N_19550,N_19302);
nor U20010 (N_20010,N_19475,N_19683);
xnor U20011 (N_20011,N_19416,N_19799);
nand U20012 (N_20012,N_19606,N_19444);
xor U20013 (N_20013,N_19639,N_19760);
and U20014 (N_20014,N_19748,N_19603);
xor U20015 (N_20015,N_19704,N_19476);
xnor U20016 (N_20016,N_19784,N_19459);
and U20017 (N_20017,N_19588,N_19442);
nand U20018 (N_20018,N_19280,N_19296);
or U20019 (N_20019,N_19236,N_19623);
or U20020 (N_20020,N_19408,N_19721);
xor U20021 (N_20021,N_19361,N_19419);
xor U20022 (N_20022,N_19229,N_19376);
nand U20023 (N_20023,N_19687,N_19611);
xnor U20024 (N_20024,N_19257,N_19745);
nand U20025 (N_20025,N_19357,N_19620);
or U20026 (N_20026,N_19341,N_19411);
xnor U20027 (N_20027,N_19547,N_19474);
or U20028 (N_20028,N_19725,N_19567);
xnor U20029 (N_20029,N_19793,N_19244);
nand U20030 (N_20030,N_19303,N_19519);
nor U20031 (N_20031,N_19346,N_19216);
xor U20032 (N_20032,N_19333,N_19569);
or U20033 (N_20033,N_19605,N_19409);
and U20034 (N_20034,N_19310,N_19486);
and U20035 (N_20035,N_19322,N_19204);
nor U20036 (N_20036,N_19427,N_19539);
nor U20037 (N_20037,N_19571,N_19657);
nand U20038 (N_20038,N_19660,N_19415);
nand U20039 (N_20039,N_19661,N_19655);
or U20040 (N_20040,N_19772,N_19295);
or U20041 (N_20041,N_19791,N_19290);
nand U20042 (N_20042,N_19367,N_19483);
xor U20043 (N_20043,N_19463,N_19712);
xnor U20044 (N_20044,N_19562,N_19414);
and U20045 (N_20045,N_19707,N_19348);
or U20046 (N_20046,N_19451,N_19719);
xor U20047 (N_20047,N_19246,N_19600);
and U20048 (N_20048,N_19650,N_19441);
nand U20049 (N_20049,N_19434,N_19355);
or U20050 (N_20050,N_19498,N_19699);
xor U20051 (N_20051,N_19266,N_19265);
xor U20052 (N_20052,N_19554,N_19214);
xnor U20053 (N_20053,N_19783,N_19782);
nand U20054 (N_20054,N_19401,N_19397);
and U20055 (N_20055,N_19315,N_19553);
nand U20056 (N_20056,N_19776,N_19582);
or U20057 (N_20057,N_19217,N_19573);
nor U20058 (N_20058,N_19364,N_19715);
xnor U20059 (N_20059,N_19494,N_19387);
or U20060 (N_20060,N_19779,N_19629);
nand U20061 (N_20061,N_19675,N_19205);
xor U20062 (N_20062,N_19658,N_19457);
nand U20063 (N_20063,N_19604,N_19724);
xnor U20064 (N_20064,N_19561,N_19388);
or U20065 (N_20065,N_19696,N_19681);
nor U20066 (N_20066,N_19365,N_19331);
nor U20067 (N_20067,N_19746,N_19248);
or U20068 (N_20068,N_19240,N_19697);
or U20069 (N_20069,N_19530,N_19297);
nand U20070 (N_20070,N_19705,N_19487);
and U20071 (N_20071,N_19263,N_19665);
nand U20072 (N_20072,N_19377,N_19478);
or U20073 (N_20073,N_19353,N_19538);
nand U20074 (N_20074,N_19467,N_19536);
or U20075 (N_20075,N_19544,N_19319);
xnor U20076 (N_20076,N_19391,N_19439);
nand U20077 (N_20077,N_19211,N_19767);
nor U20078 (N_20078,N_19294,N_19774);
and U20079 (N_20079,N_19480,N_19492);
or U20080 (N_20080,N_19584,N_19557);
and U20081 (N_20081,N_19221,N_19668);
or U20082 (N_20082,N_19443,N_19298);
nand U20083 (N_20083,N_19656,N_19511);
nor U20084 (N_20084,N_19673,N_19404);
and U20085 (N_20085,N_19586,N_19477);
nor U20086 (N_20086,N_19210,N_19394);
nor U20087 (N_20087,N_19591,N_19529);
and U20088 (N_20088,N_19309,N_19798);
nor U20089 (N_20089,N_19272,N_19329);
xor U20090 (N_20090,N_19283,N_19271);
xor U20091 (N_20091,N_19631,N_19693);
and U20092 (N_20092,N_19747,N_19392);
nand U20093 (N_20093,N_19203,N_19574);
and U20094 (N_20094,N_19372,N_19542);
and U20095 (N_20095,N_19373,N_19328);
nor U20096 (N_20096,N_19633,N_19339);
nand U20097 (N_20097,N_19670,N_19334);
nand U20098 (N_20098,N_19535,N_19425);
nor U20099 (N_20099,N_19686,N_19472);
and U20100 (N_20100,N_19331,N_19362);
and U20101 (N_20101,N_19448,N_19759);
and U20102 (N_20102,N_19259,N_19269);
nor U20103 (N_20103,N_19320,N_19663);
nor U20104 (N_20104,N_19202,N_19528);
or U20105 (N_20105,N_19270,N_19301);
xnor U20106 (N_20106,N_19680,N_19351);
xnor U20107 (N_20107,N_19406,N_19245);
xor U20108 (N_20108,N_19348,N_19536);
or U20109 (N_20109,N_19302,N_19476);
xor U20110 (N_20110,N_19416,N_19436);
and U20111 (N_20111,N_19309,N_19436);
and U20112 (N_20112,N_19251,N_19237);
nor U20113 (N_20113,N_19528,N_19328);
nor U20114 (N_20114,N_19485,N_19795);
or U20115 (N_20115,N_19533,N_19200);
and U20116 (N_20116,N_19455,N_19218);
nand U20117 (N_20117,N_19536,N_19743);
xor U20118 (N_20118,N_19710,N_19644);
and U20119 (N_20119,N_19415,N_19406);
nor U20120 (N_20120,N_19712,N_19667);
and U20121 (N_20121,N_19463,N_19330);
nand U20122 (N_20122,N_19502,N_19620);
xnor U20123 (N_20123,N_19356,N_19640);
and U20124 (N_20124,N_19207,N_19293);
or U20125 (N_20125,N_19262,N_19296);
or U20126 (N_20126,N_19327,N_19398);
xor U20127 (N_20127,N_19725,N_19227);
nand U20128 (N_20128,N_19695,N_19393);
and U20129 (N_20129,N_19336,N_19434);
and U20130 (N_20130,N_19780,N_19739);
xnor U20131 (N_20131,N_19627,N_19575);
xnor U20132 (N_20132,N_19571,N_19741);
nor U20133 (N_20133,N_19390,N_19653);
xor U20134 (N_20134,N_19503,N_19638);
or U20135 (N_20135,N_19569,N_19487);
or U20136 (N_20136,N_19500,N_19690);
or U20137 (N_20137,N_19208,N_19333);
or U20138 (N_20138,N_19331,N_19248);
nand U20139 (N_20139,N_19350,N_19362);
xor U20140 (N_20140,N_19599,N_19275);
nor U20141 (N_20141,N_19217,N_19413);
nor U20142 (N_20142,N_19474,N_19214);
nand U20143 (N_20143,N_19203,N_19439);
nor U20144 (N_20144,N_19576,N_19377);
nor U20145 (N_20145,N_19401,N_19466);
and U20146 (N_20146,N_19553,N_19312);
xnor U20147 (N_20147,N_19214,N_19696);
nand U20148 (N_20148,N_19497,N_19502);
nand U20149 (N_20149,N_19700,N_19390);
nor U20150 (N_20150,N_19720,N_19778);
xnor U20151 (N_20151,N_19283,N_19477);
nor U20152 (N_20152,N_19395,N_19788);
or U20153 (N_20153,N_19377,N_19613);
xor U20154 (N_20154,N_19202,N_19373);
and U20155 (N_20155,N_19605,N_19398);
xnor U20156 (N_20156,N_19535,N_19514);
nor U20157 (N_20157,N_19521,N_19792);
xor U20158 (N_20158,N_19582,N_19307);
nand U20159 (N_20159,N_19448,N_19496);
xnor U20160 (N_20160,N_19466,N_19372);
and U20161 (N_20161,N_19270,N_19306);
and U20162 (N_20162,N_19461,N_19798);
nand U20163 (N_20163,N_19591,N_19377);
nand U20164 (N_20164,N_19692,N_19227);
nand U20165 (N_20165,N_19421,N_19252);
xor U20166 (N_20166,N_19298,N_19779);
or U20167 (N_20167,N_19372,N_19723);
nor U20168 (N_20168,N_19668,N_19518);
or U20169 (N_20169,N_19620,N_19652);
xnor U20170 (N_20170,N_19656,N_19368);
xnor U20171 (N_20171,N_19289,N_19738);
and U20172 (N_20172,N_19756,N_19356);
nand U20173 (N_20173,N_19699,N_19684);
nor U20174 (N_20174,N_19201,N_19320);
and U20175 (N_20175,N_19550,N_19273);
xor U20176 (N_20176,N_19584,N_19324);
or U20177 (N_20177,N_19459,N_19708);
or U20178 (N_20178,N_19657,N_19495);
nand U20179 (N_20179,N_19358,N_19260);
nor U20180 (N_20180,N_19654,N_19602);
or U20181 (N_20181,N_19455,N_19673);
xor U20182 (N_20182,N_19558,N_19566);
or U20183 (N_20183,N_19361,N_19662);
and U20184 (N_20184,N_19641,N_19599);
nand U20185 (N_20185,N_19464,N_19201);
xor U20186 (N_20186,N_19216,N_19546);
nand U20187 (N_20187,N_19558,N_19470);
and U20188 (N_20188,N_19778,N_19234);
nor U20189 (N_20189,N_19617,N_19572);
xnor U20190 (N_20190,N_19654,N_19248);
nand U20191 (N_20191,N_19399,N_19768);
nor U20192 (N_20192,N_19218,N_19702);
xor U20193 (N_20193,N_19440,N_19269);
nand U20194 (N_20194,N_19241,N_19618);
and U20195 (N_20195,N_19712,N_19304);
nand U20196 (N_20196,N_19534,N_19238);
nor U20197 (N_20197,N_19568,N_19359);
nor U20198 (N_20198,N_19795,N_19428);
nor U20199 (N_20199,N_19354,N_19261);
xor U20200 (N_20200,N_19603,N_19461);
or U20201 (N_20201,N_19286,N_19482);
and U20202 (N_20202,N_19725,N_19208);
and U20203 (N_20203,N_19543,N_19551);
or U20204 (N_20204,N_19661,N_19700);
nor U20205 (N_20205,N_19690,N_19391);
nor U20206 (N_20206,N_19246,N_19567);
xnor U20207 (N_20207,N_19348,N_19546);
nor U20208 (N_20208,N_19211,N_19603);
or U20209 (N_20209,N_19753,N_19702);
and U20210 (N_20210,N_19768,N_19472);
nor U20211 (N_20211,N_19263,N_19408);
or U20212 (N_20212,N_19490,N_19211);
xnor U20213 (N_20213,N_19540,N_19686);
nor U20214 (N_20214,N_19671,N_19482);
or U20215 (N_20215,N_19493,N_19264);
xnor U20216 (N_20216,N_19242,N_19662);
or U20217 (N_20217,N_19541,N_19442);
xnor U20218 (N_20218,N_19578,N_19640);
nand U20219 (N_20219,N_19280,N_19629);
nand U20220 (N_20220,N_19652,N_19598);
xnor U20221 (N_20221,N_19233,N_19203);
xnor U20222 (N_20222,N_19298,N_19610);
and U20223 (N_20223,N_19579,N_19433);
and U20224 (N_20224,N_19428,N_19444);
or U20225 (N_20225,N_19454,N_19392);
nand U20226 (N_20226,N_19745,N_19324);
and U20227 (N_20227,N_19752,N_19680);
or U20228 (N_20228,N_19553,N_19687);
nor U20229 (N_20229,N_19603,N_19255);
nor U20230 (N_20230,N_19212,N_19369);
nand U20231 (N_20231,N_19528,N_19644);
nor U20232 (N_20232,N_19234,N_19442);
or U20233 (N_20233,N_19731,N_19264);
xnor U20234 (N_20234,N_19757,N_19669);
nor U20235 (N_20235,N_19765,N_19257);
nand U20236 (N_20236,N_19515,N_19228);
nor U20237 (N_20237,N_19236,N_19515);
nand U20238 (N_20238,N_19204,N_19332);
nor U20239 (N_20239,N_19284,N_19466);
or U20240 (N_20240,N_19754,N_19390);
xor U20241 (N_20241,N_19271,N_19560);
nand U20242 (N_20242,N_19599,N_19729);
xnor U20243 (N_20243,N_19757,N_19479);
and U20244 (N_20244,N_19727,N_19281);
nand U20245 (N_20245,N_19237,N_19374);
nor U20246 (N_20246,N_19760,N_19710);
or U20247 (N_20247,N_19228,N_19611);
or U20248 (N_20248,N_19755,N_19633);
nand U20249 (N_20249,N_19434,N_19221);
nor U20250 (N_20250,N_19479,N_19587);
and U20251 (N_20251,N_19670,N_19357);
xor U20252 (N_20252,N_19743,N_19555);
or U20253 (N_20253,N_19427,N_19516);
xor U20254 (N_20254,N_19389,N_19463);
xor U20255 (N_20255,N_19430,N_19571);
nand U20256 (N_20256,N_19687,N_19720);
or U20257 (N_20257,N_19453,N_19741);
xor U20258 (N_20258,N_19760,N_19400);
or U20259 (N_20259,N_19218,N_19766);
nor U20260 (N_20260,N_19325,N_19555);
and U20261 (N_20261,N_19331,N_19319);
xnor U20262 (N_20262,N_19799,N_19432);
and U20263 (N_20263,N_19568,N_19206);
nor U20264 (N_20264,N_19330,N_19783);
nand U20265 (N_20265,N_19316,N_19459);
nand U20266 (N_20266,N_19322,N_19481);
and U20267 (N_20267,N_19413,N_19448);
xor U20268 (N_20268,N_19359,N_19554);
nor U20269 (N_20269,N_19642,N_19428);
and U20270 (N_20270,N_19574,N_19789);
nand U20271 (N_20271,N_19367,N_19749);
nand U20272 (N_20272,N_19401,N_19325);
or U20273 (N_20273,N_19304,N_19448);
nand U20274 (N_20274,N_19443,N_19567);
nor U20275 (N_20275,N_19390,N_19736);
nor U20276 (N_20276,N_19497,N_19429);
xnor U20277 (N_20277,N_19584,N_19655);
and U20278 (N_20278,N_19539,N_19398);
or U20279 (N_20279,N_19429,N_19395);
nand U20280 (N_20280,N_19460,N_19472);
nand U20281 (N_20281,N_19330,N_19763);
nor U20282 (N_20282,N_19509,N_19236);
nand U20283 (N_20283,N_19439,N_19319);
nor U20284 (N_20284,N_19767,N_19755);
and U20285 (N_20285,N_19683,N_19315);
nand U20286 (N_20286,N_19771,N_19625);
xnor U20287 (N_20287,N_19611,N_19640);
or U20288 (N_20288,N_19563,N_19501);
or U20289 (N_20289,N_19550,N_19453);
nand U20290 (N_20290,N_19487,N_19227);
xnor U20291 (N_20291,N_19227,N_19313);
or U20292 (N_20292,N_19540,N_19367);
nor U20293 (N_20293,N_19298,N_19434);
or U20294 (N_20294,N_19671,N_19266);
nor U20295 (N_20295,N_19401,N_19573);
and U20296 (N_20296,N_19255,N_19575);
and U20297 (N_20297,N_19461,N_19317);
nand U20298 (N_20298,N_19243,N_19310);
and U20299 (N_20299,N_19401,N_19399);
nor U20300 (N_20300,N_19322,N_19211);
or U20301 (N_20301,N_19532,N_19779);
nand U20302 (N_20302,N_19491,N_19753);
nor U20303 (N_20303,N_19411,N_19471);
or U20304 (N_20304,N_19560,N_19338);
or U20305 (N_20305,N_19445,N_19495);
nor U20306 (N_20306,N_19272,N_19590);
or U20307 (N_20307,N_19658,N_19246);
nand U20308 (N_20308,N_19556,N_19698);
xnor U20309 (N_20309,N_19320,N_19750);
nor U20310 (N_20310,N_19588,N_19225);
and U20311 (N_20311,N_19341,N_19203);
xor U20312 (N_20312,N_19502,N_19742);
nor U20313 (N_20313,N_19517,N_19340);
xor U20314 (N_20314,N_19517,N_19774);
nand U20315 (N_20315,N_19258,N_19416);
or U20316 (N_20316,N_19338,N_19650);
or U20317 (N_20317,N_19666,N_19750);
or U20318 (N_20318,N_19618,N_19739);
and U20319 (N_20319,N_19707,N_19534);
or U20320 (N_20320,N_19619,N_19623);
nand U20321 (N_20321,N_19412,N_19772);
xor U20322 (N_20322,N_19344,N_19433);
or U20323 (N_20323,N_19764,N_19747);
nand U20324 (N_20324,N_19622,N_19752);
nor U20325 (N_20325,N_19201,N_19388);
nor U20326 (N_20326,N_19526,N_19546);
xor U20327 (N_20327,N_19588,N_19628);
and U20328 (N_20328,N_19628,N_19513);
nor U20329 (N_20329,N_19557,N_19581);
or U20330 (N_20330,N_19792,N_19321);
and U20331 (N_20331,N_19561,N_19640);
and U20332 (N_20332,N_19595,N_19741);
or U20333 (N_20333,N_19483,N_19776);
and U20334 (N_20334,N_19350,N_19709);
and U20335 (N_20335,N_19421,N_19631);
nor U20336 (N_20336,N_19595,N_19776);
nand U20337 (N_20337,N_19718,N_19436);
nor U20338 (N_20338,N_19294,N_19694);
nor U20339 (N_20339,N_19229,N_19725);
nand U20340 (N_20340,N_19306,N_19729);
nand U20341 (N_20341,N_19241,N_19673);
nor U20342 (N_20342,N_19739,N_19726);
and U20343 (N_20343,N_19217,N_19668);
nand U20344 (N_20344,N_19420,N_19346);
and U20345 (N_20345,N_19645,N_19755);
nor U20346 (N_20346,N_19228,N_19580);
nand U20347 (N_20347,N_19548,N_19333);
nand U20348 (N_20348,N_19646,N_19781);
xor U20349 (N_20349,N_19314,N_19706);
nand U20350 (N_20350,N_19524,N_19232);
nor U20351 (N_20351,N_19728,N_19205);
or U20352 (N_20352,N_19226,N_19478);
and U20353 (N_20353,N_19292,N_19655);
or U20354 (N_20354,N_19281,N_19765);
nand U20355 (N_20355,N_19325,N_19773);
nand U20356 (N_20356,N_19342,N_19385);
nand U20357 (N_20357,N_19583,N_19287);
xnor U20358 (N_20358,N_19445,N_19640);
xor U20359 (N_20359,N_19595,N_19609);
nand U20360 (N_20360,N_19553,N_19799);
and U20361 (N_20361,N_19658,N_19368);
xnor U20362 (N_20362,N_19470,N_19474);
and U20363 (N_20363,N_19673,N_19716);
nor U20364 (N_20364,N_19609,N_19429);
nand U20365 (N_20365,N_19693,N_19221);
nand U20366 (N_20366,N_19798,N_19474);
or U20367 (N_20367,N_19520,N_19616);
nand U20368 (N_20368,N_19636,N_19318);
nand U20369 (N_20369,N_19507,N_19571);
xnor U20370 (N_20370,N_19344,N_19480);
nor U20371 (N_20371,N_19519,N_19328);
nor U20372 (N_20372,N_19647,N_19656);
and U20373 (N_20373,N_19396,N_19644);
nor U20374 (N_20374,N_19486,N_19425);
or U20375 (N_20375,N_19779,N_19581);
xnor U20376 (N_20376,N_19564,N_19364);
nand U20377 (N_20377,N_19625,N_19703);
or U20378 (N_20378,N_19423,N_19376);
nor U20379 (N_20379,N_19323,N_19601);
nor U20380 (N_20380,N_19213,N_19644);
and U20381 (N_20381,N_19273,N_19261);
nand U20382 (N_20382,N_19718,N_19754);
nor U20383 (N_20383,N_19653,N_19749);
or U20384 (N_20384,N_19696,N_19512);
and U20385 (N_20385,N_19313,N_19649);
or U20386 (N_20386,N_19504,N_19621);
nand U20387 (N_20387,N_19408,N_19325);
or U20388 (N_20388,N_19495,N_19601);
xnor U20389 (N_20389,N_19316,N_19485);
xnor U20390 (N_20390,N_19751,N_19492);
nor U20391 (N_20391,N_19383,N_19682);
or U20392 (N_20392,N_19674,N_19669);
and U20393 (N_20393,N_19638,N_19431);
nand U20394 (N_20394,N_19561,N_19301);
or U20395 (N_20395,N_19418,N_19404);
xnor U20396 (N_20396,N_19514,N_19567);
nor U20397 (N_20397,N_19575,N_19284);
and U20398 (N_20398,N_19274,N_19743);
nand U20399 (N_20399,N_19658,N_19314);
and U20400 (N_20400,N_19983,N_20021);
nor U20401 (N_20401,N_20133,N_20104);
nor U20402 (N_20402,N_20385,N_20320);
nand U20403 (N_20403,N_19894,N_20022);
and U20404 (N_20404,N_19886,N_19833);
nand U20405 (N_20405,N_20028,N_19847);
nand U20406 (N_20406,N_19980,N_19997);
or U20407 (N_20407,N_20398,N_19982);
nor U20408 (N_20408,N_20006,N_19908);
nand U20409 (N_20409,N_20185,N_20077);
nand U20410 (N_20410,N_20357,N_20205);
nand U20411 (N_20411,N_20075,N_20298);
or U20412 (N_20412,N_20321,N_19859);
nand U20413 (N_20413,N_20295,N_20181);
xor U20414 (N_20414,N_20146,N_20217);
xor U20415 (N_20415,N_19905,N_19897);
xnor U20416 (N_20416,N_19920,N_20305);
or U20417 (N_20417,N_20102,N_20358);
xor U20418 (N_20418,N_20086,N_20340);
and U20419 (N_20419,N_20203,N_20176);
nand U20420 (N_20420,N_19856,N_20277);
or U20421 (N_20421,N_19973,N_19870);
xor U20422 (N_20422,N_19869,N_20148);
nand U20423 (N_20423,N_20281,N_20116);
xnor U20424 (N_20424,N_20239,N_19801);
nor U20425 (N_20425,N_20323,N_20338);
or U20426 (N_20426,N_19955,N_19954);
and U20427 (N_20427,N_20184,N_19812);
and U20428 (N_20428,N_20063,N_20393);
or U20429 (N_20429,N_20200,N_20352);
nor U20430 (N_20430,N_19951,N_20317);
or U20431 (N_20431,N_20384,N_20128);
and U20432 (N_20432,N_20225,N_20078);
nand U20433 (N_20433,N_19975,N_20353);
nand U20434 (N_20434,N_20160,N_19946);
and U20435 (N_20435,N_19860,N_20315);
nand U20436 (N_20436,N_19826,N_20057);
nand U20437 (N_20437,N_19825,N_19985);
nand U20438 (N_20438,N_20129,N_19978);
nor U20439 (N_20439,N_20227,N_20339);
xnor U20440 (N_20440,N_19800,N_19844);
and U20441 (N_20441,N_20049,N_20241);
nor U20442 (N_20442,N_20346,N_19810);
xor U20443 (N_20443,N_19994,N_20334);
nor U20444 (N_20444,N_20264,N_19879);
nor U20445 (N_20445,N_19814,N_20061);
or U20446 (N_20446,N_19881,N_20190);
nor U20447 (N_20447,N_20262,N_20388);
or U20448 (N_20448,N_20103,N_20294);
nand U20449 (N_20449,N_20003,N_20117);
and U20450 (N_20450,N_20301,N_20223);
nand U20451 (N_20451,N_20072,N_19872);
xor U20452 (N_20452,N_20267,N_20114);
xor U20453 (N_20453,N_20329,N_19930);
or U20454 (N_20454,N_19827,N_19952);
and U20455 (N_20455,N_20178,N_20081);
and U20456 (N_20456,N_19862,N_19883);
or U20457 (N_20457,N_20067,N_20194);
xnor U20458 (N_20458,N_20261,N_20259);
and U20459 (N_20459,N_19807,N_19922);
nand U20460 (N_20460,N_20130,N_20382);
nor U20461 (N_20461,N_19803,N_19857);
xor U20462 (N_20462,N_19838,N_20328);
xor U20463 (N_20463,N_20379,N_20175);
nand U20464 (N_20464,N_20371,N_19903);
or U20465 (N_20465,N_20150,N_20218);
nor U20466 (N_20466,N_19926,N_20232);
nor U20467 (N_20467,N_20091,N_20009);
nor U20468 (N_20468,N_20345,N_20138);
nor U20469 (N_20469,N_20054,N_20202);
xor U20470 (N_20470,N_20216,N_20020);
xnor U20471 (N_20471,N_20083,N_20173);
nand U20472 (N_20472,N_19972,N_19828);
and U20473 (N_20473,N_20044,N_20052);
and U20474 (N_20474,N_19840,N_20390);
nor U20475 (N_20475,N_19836,N_20155);
nand U20476 (N_20476,N_20271,N_20397);
nand U20477 (N_20477,N_20013,N_19910);
nor U20478 (N_20478,N_20221,N_20197);
or U20479 (N_20479,N_19839,N_20211);
and U20480 (N_20480,N_20363,N_20389);
nand U20481 (N_20481,N_20122,N_19895);
or U20482 (N_20482,N_20163,N_20399);
nor U20483 (N_20483,N_20387,N_19864);
nand U20484 (N_20484,N_19964,N_20159);
or U20485 (N_20485,N_20204,N_19988);
and U20486 (N_20486,N_20378,N_20153);
xor U20487 (N_20487,N_20235,N_20237);
nand U20488 (N_20488,N_20268,N_20325);
xnor U20489 (N_20489,N_20099,N_20210);
and U20490 (N_20490,N_20326,N_20011);
and U20491 (N_20491,N_19877,N_20302);
xor U20492 (N_20492,N_19932,N_20288);
nand U20493 (N_20493,N_19884,N_20018);
and U20494 (N_20494,N_20125,N_19929);
nand U20495 (N_20495,N_20079,N_20025);
xnor U20496 (N_20496,N_20347,N_20036);
xnor U20497 (N_20497,N_20359,N_19842);
xor U20498 (N_20498,N_19928,N_20220);
nor U20499 (N_20499,N_19934,N_20166);
xor U20500 (N_20500,N_20004,N_19942);
and U20501 (N_20501,N_20058,N_20222);
xnor U20502 (N_20502,N_20010,N_19949);
xor U20503 (N_20503,N_19958,N_20139);
or U20504 (N_20504,N_20002,N_19945);
xor U20505 (N_20505,N_19849,N_20141);
xor U20506 (N_20506,N_19907,N_20219);
and U20507 (N_20507,N_20350,N_20215);
or U20508 (N_20508,N_20073,N_20364);
xor U20509 (N_20509,N_20319,N_20233);
and U20510 (N_20510,N_20123,N_19937);
xor U20511 (N_20511,N_19850,N_20135);
or U20512 (N_20512,N_20093,N_20087);
and U20513 (N_20513,N_19858,N_19813);
and U20514 (N_20514,N_20132,N_20307);
and U20515 (N_20515,N_20381,N_20206);
nor U20516 (N_20516,N_20266,N_20105);
nor U20517 (N_20517,N_20292,N_20279);
or U20518 (N_20518,N_20048,N_20253);
xnor U20519 (N_20519,N_20275,N_19999);
xnor U20520 (N_20520,N_20098,N_20213);
or U20521 (N_20521,N_20245,N_20270);
nor U20522 (N_20522,N_19968,N_20107);
and U20523 (N_20523,N_20088,N_20349);
and U20524 (N_20524,N_20084,N_20053);
or U20525 (N_20525,N_20019,N_20059);
and U20526 (N_20526,N_19868,N_19984);
xnor U20527 (N_20527,N_20318,N_20256);
nand U20528 (N_20528,N_19967,N_20108);
and U20529 (N_20529,N_20195,N_20312);
or U20530 (N_20530,N_19866,N_19936);
or U20531 (N_20531,N_19939,N_19888);
xor U20532 (N_20532,N_20171,N_19875);
nand U20533 (N_20533,N_20137,N_20240);
nand U20534 (N_20534,N_20276,N_20333);
nand U20535 (N_20535,N_20322,N_20042);
xnor U20536 (N_20536,N_19899,N_19986);
or U20537 (N_20537,N_20030,N_20074);
nor U20538 (N_20538,N_19818,N_20395);
and U20539 (N_20539,N_20386,N_20014);
nor U20540 (N_20540,N_19918,N_20001);
nor U20541 (N_20541,N_20291,N_20335);
nor U20542 (N_20542,N_20287,N_19824);
and U20543 (N_20543,N_19965,N_20273);
xor U20544 (N_20544,N_19811,N_20110);
and U20545 (N_20545,N_20174,N_20115);
or U20546 (N_20546,N_20283,N_20118);
and U20547 (N_20547,N_19969,N_19874);
and U20548 (N_20548,N_19890,N_20066);
nor U20549 (N_20549,N_20265,N_20039);
nand U20550 (N_20550,N_19846,N_20300);
nand U20551 (N_20551,N_19933,N_20119);
nor U20552 (N_20552,N_20188,N_20306);
or U20553 (N_20553,N_19919,N_19817);
and U20554 (N_20554,N_20070,N_19804);
or U20555 (N_20555,N_20289,N_19898);
and U20556 (N_20556,N_20196,N_19896);
or U20557 (N_20557,N_20201,N_20165);
or U20558 (N_20558,N_20244,N_19809);
and U20559 (N_20559,N_20127,N_20280);
xor U20560 (N_20560,N_19876,N_20154);
or U20561 (N_20561,N_19855,N_20076);
nor U20562 (N_20562,N_19921,N_19863);
or U20563 (N_20563,N_19923,N_19829);
nor U20564 (N_20564,N_20258,N_19887);
xor U20565 (N_20565,N_19831,N_20140);
and U20566 (N_20566,N_19943,N_20156);
nor U20567 (N_20567,N_19971,N_19996);
nor U20568 (N_20568,N_20332,N_20182);
and U20569 (N_20569,N_20016,N_20094);
nor U20570 (N_20570,N_20231,N_20372);
and U20571 (N_20571,N_19916,N_20136);
and U20572 (N_20572,N_19808,N_20193);
nor U20573 (N_20573,N_19832,N_20354);
or U20574 (N_20574,N_20278,N_19802);
xor U20575 (N_20575,N_20282,N_19950);
nand U20576 (N_20576,N_19901,N_20254);
and U20577 (N_20577,N_20164,N_19885);
xnor U20578 (N_20578,N_20012,N_19822);
nor U20579 (N_20579,N_19956,N_20041);
nand U20580 (N_20580,N_19957,N_20391);
and U20581 (N_20581,N_20090,N_20029);
xor U20582 (N_20582,N_20369,N_19873);
xnor U20583 (N_20583,N_20224,N_20069);
or U20584 (N_20584,N_20064,N_20170);
nand U20585 (N_20585,N_20285,N_20242);
xnor U20586 (N_20586,N_20131,N_20027);
xor U20587 (N_20587,N_19959,N_20269);
xnor U20588 (N_20588,N_20272,N_20361);
xor U20589 (N_20589,N_19977,N_20297);
or U20590 (N_20590,N_20327,N_20167);
and U20591 (N_20591,N_19806,N_20043);
nor U20592 (N_20592,N_19947,N_19998);
nor U20593 (N_20593,N_19906,N_19991);
or U20594 (N_20594,N_20299,N_20296);
or U20595 (N_20595,N_20038,N_19990);
nor U20596 (N_20596,N_19880,N_19837);
nor U20597 (N_20597,N_20375,N_20007);
xnor U20598 (N_20598,N_20208,N_19892);
nor U20599 (N_20599,N_20092,N_19834);
xor U20600 (N_20600,N_20168,N_20362);
xnor U20601 (N_20601,N_20366,N_20144);
and U20602 (N_20602,N_20311,N_20226);
or U20603 (N_20603,N_20274,N_19995);
or U20604 (N_20604,N_20095,N_20290);
and U20605 (N_20605,N_20121,N_19893);
and U20606 (N_20606,N_20032,N_20343);
nand U20607 (N_20607,N_19976,N_20047);
nand U20608 (N_20608,N_20045,N_20157);
xnor U20609 (N_20609,N_20065,N_20341);
nor U20610 (N_20610,N_20192,N_19963);
nor U20611 (N_20611,N_20100,N_20096);
xnor U20612 (N_20612,N_19845,N_20180);
nand U20613 (N_20613,N_20199,N_20189);
and U20614 (N_20614,N_20152,N_19835);
or U20615 (N_20615,N_20330,N_20026);
nand U20616 (N_20616,N_19953,N_20005);
nor U20617 (N_20617,N_19843,N_20324);
or U20618 (N_20618,N_20255,N_20071);
nand U20619 (N_20619,N_19815,N_20106);
and U20620 (N_20620,N_19924,N_20313);
xor U20621 (N_20621,N_19913,N_19851);
or U20622 (N_20622,N_20172,N_20304);
xnor U20623 (N_20623,N_19981,N_19940);
or U20624 (N_20624,N_20342,N_19992);
xnor U20625 (N_20625,N_19917,N_20250);
nand U20626 (N_20626,N_19871,N_20394);
and U20627 (N_20627,N_20257,N_20344);
nand U20628 (N_20628,N_20260,N_20023);
and U20629 (N_20629,N_20068,N_19889);
nand U20630 (N_20630,N_19948,N_20310);
nand U20631 (N_20631,N_20238,N_20198);
nor U20632 (N_20632,N_20249,N_20368);
and U20633 (N_20633,N_20120,N_20143);
xor U20634 (N_20634,N_20112,N_19974);
nor U20635 (N_20635,N_19935,N_20314);
xor U20636 (N_20636,N_20050,N_20251);
and U20637 (N_20637,N_19993,N_20089);
and U20638 (N_20638,N_20024,N_20035);
nand U20639 (N_20639,N_20337,N_20179);
and U20640 (N_20640,N_20230,N_19961);
xor U20641 (N_20641,N_20355,N_19878);
or U20642 (N_20642,N_20284,N_19987);
xnor U20643 (N_20643,N_20263,N_19861);
nor U20644 (N_20644,N_20101,N_20046);
or U20645 (N_20645,N_20008,N_20097);
xor U20646 (N_20646,N_20331,N_20017);
nor U20647 (N_20647,N_20209,N_20082);
or U20648 (N_20648,N_19962,N_20034);
and U20649 (N_20649,N_20374,N_20365);
nor U20650 (N_20650,N_20085,N_20062);
nor U20651 (N_20651,N_20126,N_19882);
nor U20652 (N_20652,N_20396,N_20336);
and U20653 (N_20653,N_20243,N_20348);
nor U20654 (N_20654,N_20111,N_20351);
xor U20655 (N_20655,N_20316,N_19820);
and U20656 (N_20656,N_20370,N_20383);
and U20657 (N_20657,N_19853,N_20303);
xor U20658 (N_20658,N_19841,N_19902);
nor U20659 (N_20659,N_20113,N_20234);
nand U20660 (N_20660,N_20367,N_19823);
nor U20661 (N_20661,N_19912,N_20247);
nand U20662 (N_20662,N_20214,N_20124);
nand U20663 (N_20663,N_19891,N_19970);
nand U20664 (N_20664,N_20145,N_19915);
nand U20665 (N_20665,N_19925,N_19960);
nand U20666 (N_20666,N_20246,N_19966);
xnor U20667 (N_20667,N_20228,N_20293);
or U20668 (N_20668,N_19805,N_19867);
nor U20669 (N_20669,N_20248,N_20309);
and U20670 (N_20670,N_20177,N_20080);
nor U20671 (N_20671,N_20147,N_20033);
and U20672 (N_20672,N_19904,N_20376);
nand U20673 (N_20673,N_20037,N_20392);
xnor U20674 (N_20674,N_20109,N_19865);
nand U20675 (N_20675,N_19938,N_19927);
xnor U20676 (N_20676,N_20187,N_20183);
xnor U20677 (N_20677,N_19819,N_19821);
and U20678 (N_20678,N_19911,N_20055);
nand U20679 (N_20679,N_20191,N_20134);
xor U20680 (N_20680,N_20373,N_19944);
nand U20681 (N_20681,N_19830,N_19979);
xnor U20682 (N_20682,N_20149,N_20252);
nor U20683 (N_20683,N_19900,N_20031);
or U20684 (N_20684,N_19909,N_20380);
or U20685 (N_20685,N_20212,N_20308);
nor U20686 (N_20686,N_20151,N_19848);
nor U20687 (N_20687,N_19941,N_20162);
nor U20688 (N_20688,N_20229,N_20056);
or U20689 (N_20689,N_20051,N_20060);
and U20690 (N_20690,N_20000,N_20356);
nand U20691 (N_20691,N_19852,N_20161);
nor U20692 (N_20692,N_20186,N_20286);
xor U20693 (N_20693,N_19914,N_20040);
and U20694 (N_20694,N_19816,N_19931);
or U20695 (N_20695,N_20207,N_20015);
or U20696 (N_20696,N_20377,N_20158);
and U20697 (N_20697,N_20360,N_20236);
nand U20698 (N_20698,N_19989,N_20169);
nand U20699 (N_20699,N_19854,N_20142);
nand U20700 (N_20700,N_20172,N_20077);
xor U20701 (N_20701,N_20066,N_20109);
xnor U20702 (N_20702,N_20151,N_19865);
nor U20703 (N_20703,N_19856,N_20249);
nor U20704 (N_20704,N_20316,N_20131);
xnor U20705 (N_20705,N_20035,N_19863);
nand U20706 (N_20706,N_20181,N_20252);
nor U20707 (N_20707,N_20387,N_20329);
nor U20708 (N_20708,N_19821,N_20056);
nand U20709 (N_20709,N_20003,N_20178);
xor U20710 (N_20710,N_20187,N_20102);
xor U20711 (N_20711,N_19975,N_19861);
nor U20712 (N_20712,N_20121,N_19904);
nand U20713 (N_20713,N_20208,N_19873);
nand U20714 (N_20714,N_19896,N_20161);
nor U20715 (N_20715,N_20263,N_19832);
xnor U20716 (N_20716,N_19924,N_20113);
nand U20717 (N_20717,N_20383,N_20232);
or U20718 (N_20718,N_20153,N_19990);
nor U20719 (N_20719,N_20132,N_20090);
or U20720 (N_20720,N_19951,N_20047);
nand U20721 (N_20721,N_19845,N_20149);
xnor U20722 (N_20722,N_19918,N_19992);
xor U20723 (N_20723,N_19900,N_20379);
nand U20724 (N_20724,N_20208,N_20325);
and U20725 (N_20725,N_20340,N_19938);
or U20726 (N_20726,N_20128,N_20071);
and U20727 (N_20727,N_20036,N_19944);
nand U20728 (N_20728,N_20192,N_20025);
and U20729 (N_20729,N_20052,N_20383);
xor U20730 (N_20730,N_19899,N_20346);
and U20731 (N_20731,N_20270,N_20389);
nand U20732 (N_20732,N_20305,N_20348);
nand U20733 (N_20733,N_19854,N_19942);
nand U20734 (N_20734,N_19898,N_20104);
xor U20735 (N_20735,N_20290,N_20283);
nand U20736 (N_20736,N_19865,N_20272);
or U20737 (N_20737,N_19895,N_20242);
xnor U20738 (N_20738,N_20345,N_20350);
nor U20739 (N_20739,N_19837,N_20246);
and U20740 (N_20740,N_20044,N_19884);
nand U20741 (N_20741,N_20399,N_19839);
and U20742 (N_20742,N_20155,N_20134);
nand U20743 (N_20743,N_20203,N_20163);
xnor U20744 (N_20744,N_20056,N_19957);
or U20745 (N_20745,N_19822,N_20302);
and U20746 (N_20746,N_19867,N_19880);
and U20747 (N_20747,N_20335,N_20127);
nor U20748 (N_20748,N_20220,N_19961);
or U20749 (N_20749,N_20245,N_20127);
xor U20750 (N_20750,N_20134,N_19984);
nand U20751 (N_20751,N_20114,N_19863);
xnor U20752 (N_20752,N_20399,N_19812);
nor U20753 (N_20753,N_19946,N_20029);
or U20754 (N_20754,N_20202,N_20295);
xor U20755 (N_20755,N_20105,N_20294);
and U20756 (N_20756,N_20076,N_20279);
nand U20757 (N_20757,N_20204,N_20054);
nand U20758 (N_20758,N_20065,N_20382);
nand U20759 (N_20759,N_20209,N_20057);
nand U20760 (N_20760,N_19930,N_20274);
nor U20761 (N_20761,N_20088,N_20314);
and U20762 (N_20762,N_20045,N_20341);
nand U20763 (N_20763,N_20103,N_19887);
nand U20764 (N_20764,N_19839,N_20240);
xnor U20765 (N_20765,N_20399,N_20386);
and U20766 (N_20766,N_20067,N_20138);
or U20767 (N_20767,N_20342,N_19938);
or U20768 (N_20768,N_19923,N_19955);
nand U20769 (N_20769,N_19937,N_20092);
nand U20770 (N_20770,N_20070,N_19904);
and U20771 (N_20771,N_20222,N_19934);
or U20772 (N_20772,N_20263,N_19807);
and U20773 (N_20773,N_20362,N_19915);
or U20774 (N_20774,N_19838,N_19992);
nand U20775 (N_20775,N_20376,N_20044);
xnor U20776 (N_20776,N_19852,N_20041);
nor U20777 (N_20777,N_20380,N_19823);
or U20778 (N_20778,N_20080,N_20354);
xor U20779 (N_20779,N_20070,N_20232);
nand U20780 (N_20780,N_20025,N_19858);
and U20781 (N_20781,N_20036,N_20213);
and U20782 (N_20782,N_20393,N_19980);
xnor U20783 (N_20783,N_20302,N_20298);
nor U20784 (N_20784,N_20350,N_20094);
and U20785 (N_20785,N_20397,N_20216);
nand U20786 (N_20786,N_19967,N_20258);
and U20787 (N_20787,N_20183,N_20201);
or U20788 (N_20788,N_20139,N_20152);
nand U20789 (N_20789,N_20097,N_20277);
xnor U20790 (N_20790,N_20244,N_20152);
xnor U20791 (N_20791,N_19918,N_20037);
nor U20792 (N_20792,N_20126,N_20394);
nor U20793 (N_20793,N_20372,N_19977);
nand U20794 (N_20794,N_19865,N_20306);
or U20795 (N_20795,N_20309,N_19929);
xnor U20796 (N_20796,N_20073,N_20113);
and U20797 (N_20797,N_20201,N_19813);
nor U20798 (N_20798,N_19997,N_19888);
xnor U20799 (N_20799,N_19886,N_19928);
xnor U20800 (N_20800,N_20332,N_20305);
nor U20801 (N_20801,N_20306,N_19827);
nor U20802 (N_20802,N_19836,N_20163);
nor U20803 (N_20803,N_20041,N_19868);
or U20804 (N_20804,N_20244,N_19857);
or U20805 (N_20805,N_20288,N_20380);
xor U20806 (N_20806,N_19809,N_20014);
and U20807 (N_20807,N_20389,N_19928);
and U20808 (N_20808,N_20038,N_20371);
xnor U20809 (N_20809,N_19907,N_20233);
xnor U20810 (N_20810,N_20227,N_19909);
xor U20811 (N_20811,N_19841,N_20309);
or U20812 (N_20812,N_20059,N_20379);
nor U20813 (N_20813,N_19859,N_19844);
nor U20814 (N_20814,N_19918,N_20207);
nand U20815 (N_20815,N_19846,N_20225);
nand U20816 (N_20816,N_19913,N_19908);
xor U20817 (N_20817,N_20119,N_20093);
nor U20818 (N_20818,N_20063,N_19869);
nand U20819 (N_20819,N_19987,N_20309);
nor U20820 (N_20820,N_19840,N_20040);
xor U20821 (N_20821,N_20029,N_19811);
or U20822 (N_20822,N_19952,N_20135);
or U20823 (N_20823,N_20278,N_20177);
xor U20824 (N_20824,N_20160,N_19887);
and U20825 (N_20825,N_20191,N_20027);
xnor U20826 (N_20826,N_20107,N_20158);
or U20827 (N_20827,N_20017,N_20071);
xnor U20828 (N_20828,N_20296,N_20230);
nand U20829 (N_20829,N_19976,N_20348);
and U20830 (N_20830,N_20343,N_20223);
xnor U20831 (N_20831,N_19937,N_20109);
nand U20832 (N_20832,N_20235,N_20053);
nor U20833 (N_20833,N_20333,N_20045);
xnor U20834 (N_20834,N_19908,N_20041);
and U20835 (N_20835,N_20169,N_19924);
xor U20836 (N_20836,N_20098,N_19931);
nor U20837 (N_20837,N_20091,N_20063);
and U20838 (N_20838,N_19843,N_20359);
nand U20839 (N_20839,N_19881,N_20055);
xor U20840 (N_20840,N_20289,N_20185);
xnor U20841 (N_20841,N_19991,N_19976);
and U20842 (N_20842,N_19864,N_20038);
nand U20843 (N_20843,N_20263,N_19804);
nand U20844 (N_20844,N_20074,N_20108);
nor U20845 (N_20845,N_20033,N_20298);
nand U20846 (N_20846,N_20087,N_20329);
nor U20847 (N_20847,N_20138,N_19806);
or U20848 (N_20848,N_19995,N_19944);
xnor U20849 (N_20849,N_19968,N_19908);
nand U20850 (N_20850,N_20264,N_19972);
nand U20851 (N_20851,N_19949,N_20066);
nand U20852 (N_20852,N_19815,N_20293);
and U20853 (N_20853,N_20016,N_20001);
nand U20854 (N_20854,N_20192,N_20135);
nor U20855 (N_20855,N_20152,N_20064);
and U20856 (N_20856,N_20006,N_20266);
or U20857 (N_20857,N_20186,N_19803);
nand U20858 (N_20858,N_19948,N_19975);
nor U20859 (N_20859,N_19870,N_19949);
nor U20860 (N_20860,N_20281,N_20126);
and U20861 (N_20861,N_20081,N_20358);
nor U20862 (N_20862,N_19914,N_20227);
xnor U20863 (N_20863,N_20266,N_20054);
xnor U20864 (N_20864,N_20080,N_20025);
nand U20865 (N_20865,N_20389,N_20294);
or U20866 (N_20866,N_20338,N_20227);
xor U20867 (N_20867,N_20318,N_20352);
or U20868 (N_20868,N_20371,N_20313);
xnor U20869 (N_20869,N_20063,N_20060);
and U20870 (N_20870,N_19894,N_20356);
or U20871 (N_20871,N_20319,N_20081);
or U20872 (N_20872,N_20176,N_20268);
nor U20873 (N_20873,N_20330,N_20256);
and U20874 (N_20874,N_19906,N_20300);
nor U20875 (N_20875,N_20135,N_19812);
xor U20876 (N_20876,N_20091,N_20020);
nand U20877 (N_20877,N_20331,N_20372);
nand U20878 (N_20878,N_20225,N_20291);
xnor U20879 (N_20879,N_20281,N_19976);
nor U20880 (N_20880,N_19863,N_19954);
or U20881 (N_20881,N_20321,N_19881);
xnor U20882 (N_20882,N_20107,N_19826);
xnor U20883 (N_20883,N_20297,N_19846);
nor U20884 (N_20884,N_20265,N_20228);
or U20885 (N_20885,N_20185,N_20247);
nor U20886 (N_20886,N_20250,N_19859);
nand U20887 (N_20887,N_19905,N_20060);
nand U20888 (N_20888,N_19819,N_19897);
nand U20889 (N_20889,N_20061,N_20195);
xor U20890 (N_20890,N_20182,N_20057);
or U20891 (N_20891,N_19862,N_20285);
xnor U20892 (N_20892,N_19966,N_19909);
and U20893 (N_20893,N_20304,N_20227);
nand U20894 (N_20894,N_20240,N_19843);
nand U20895 (N_20895,N_20027,N_20235);
nand U20896 (N_20896,N_20393,N_19863);
and U20897 (N_20897,N_19806,N_19891);
nand U20898 (N_20898,N_20132,N_20243);
and U20899 (N_20899,N_20098,N_20123);
nand U20900 (N_20900,N_20026,N_20146);
nand U20901 (N_20901,N_19994,N_20097);
nand U20902 (N_20902,N_20115,N_20395);
nand U20903 (N_20903,N_20000,N_19873);
nor U20904 (N_20904,N_20305,N_19872);
xor U20905 (N_20905,N_20177,N_20210);
xor U20906 (N_20906,N_20057,N_20173);
xnor U20907 (N_20907,N_20122,N_19892);
nor U20908 (N_20908,N_20094,N_19840);
xnor U20909 (N_20909,N_20088,N_20221);
xor U20910 (N_20910,N_20014,N_20140);
nor U20911 (N_20911,N_19941,N_19944);
xor U20912 (N_20912,N_20089,N_20375);
xor U20913 (N_20913,N_19815,N_20100);
or U20914 (N_20914,N_19961,N_20047);
xnor U20915 (N_20915,N_19868,N_20223);
or U20916 (N_20916,N_19890,N_20055);
nor U20917 (N_20917,N_20198,N_20258);
or U20918 (N_20918,N_19924,N_20106);
or U20919 (N_20919,N_20209,N_19954);
and U20920 (N_20920,N_20184,N_19921);
nor U20921 (N_20921,N_20125,N_20352);
and U20922 (N_20922,N_20029,N_19813);
xnor U20923 (N_20923,N_19840,N_20082);
nand U20924 (N_20924,N_20031,N_20052);
and U20925 (N_20925,N_20222,N_19905);
nand U20926 (N_20926,N_19953,N_19875);
or U20927 (N_20927,N_20022,N_20032);
or U20928 (N_20928,N_19899,N_19939);
nor U20929 (N_20929,N_20076,N_20251);
xor U20930 (N_20930,N_19959,N_20173);
or U20931 (N_20931,N_20198,N_19891);
nand U20932 (N_20932,N_20250,N_19885);
nand U20933 (N_20933,N_20261,N_19978);
or U20934 (N_20934,N_20125,N_20192);
nor U20935 (N_20935,N_19996,N_19808);
and U20936 (N_20936,N_20229,N_19947);
xor U20937 (N_20937,N_20383,N_19856);
nand U20938 (N_20938,N_19944,N_19950);
or U20939 (N_20939,N_20013,N_20383);
nor U20940 (N_20940,N_19823,N_20090);
or U20941 (N_20941,N_20348,N_19871);
or U20942 (N_20942,N_19854,N_20368);
nor U20943 (N_20943,N_19838,N_20067);
or U20944 (N_20944,N_19852,N_20056);
nor U20945 (N_20945,N_20390,N_20394);
nand U20946 (N_20946,N_19923,N_20381);
and U20947 (N_20947,N_19867,N_19891);
nand U20948 (N_20948,N_19890,N_19856);
nand U20949 (N_20949,N_20116,N_19914);
and U20950 (N_20950,N_20095,N_20211);
nor U20951 (N_20951,N_19915,N_20310);
nor U20952 (N_20952,N_19980,N_19820);
nor U20953 (N_20953,N_19893,N_20211);
nand U20954 (N_20954,N_20085,N_19848);
nand U20955 (N_20955,N_20221,N_20279);
or U20956 (N_20956,N_19836,N_19845);
and U20957 (N_20957,N_20054,N_20397);
or U20958 (N_20958,N_20353,N_20356);
xor U20959 (N_20959,N_20002,N_20364);
and U20960 (N_20960,N_20252,N_19809);
or U20961 (N_20961,N_19924,N_20386);
or U20962 (N_20962,N_20300,N_19894);
and U20963 (N_20963,N_19822,N_19867);
nand U20964 (N_20964,N_19944,N_19815);
nor U20965 (N_20965,N_19814,N_20267);
and U20966 (N_20966,N_20361,N_19905);
xnor U20967 (N_20967,N_20382,N_19858);
and U20968 (N_20968,N_20015,N_20051);
nor U20969 (N_20969,N_20240,N_20022);
or U20970 (N_20970,N_19826,N_20200);
nor U20971 (N_20971,N_19984,N_20064);
and U20972 (N_20972,N_20040,N_19972);
xnor U20973 (N_20973,N_20035,N_20101);
nand U20974 (N_20974,N_20251,N_20198);
xor U20975 (N_20975,N_19843,N_20329);
nor U20976 (N_20976,N_20062,N_20315);
nor U20977 (N_20977,N_20011,N_20213);
nand U20978 (N_20978,N_20297,N_19884);
or U20979 (N_20979,N_20204,N_20005);
xor U20980 (N_20980,N_19816,N_20378);
nand U20981 (N_20981,N_20361,N_19877);
nand U20982 (N_20982,N_20160,N_19866);
nand U20983 (N_20983,N_20147,N_20048);
xor U20984 (N_20984,N_20298,N_20062);
and U20985 (N_20985,N_19976,N_20157);
or U20986 (N_20986,N_20307,N_19904);
nor U20987 (N_20987,N_20081,N_20247);
and U20988 (N_20988,N_20289,N_20252);
xnor U20989 (N_20989,N_20199,N_20299);
nor U20990 (N_20990,N_19991,N_19864);
nor U20991 (N_20991,N_20366,N_20044);
nor U20992 (N_20992,N_20224,N_20172);
xnor U20993 (N_20993,N_19920,N_19866);
or U20994 (N_20994,N_20223,N_20013);
or U20995 (N_20995,N_19895,N_20068);
or U20996 (N_20996,N_19800,N_19950);
xnor U20997 (N_20997,N_20138,N_20177);
nand U20998 (N_20998,N_20297,N_20261);
and U20999 (N_20999,N_19968,N_20390);
nand U21000 (N_21000,N_20902,N_20643);
or U21001 (N_21001,N_20919,N_20800);
xor U21002 (N_21002,N_20869,N_20593);
nor U21003 (N_21003,N_20415,N_20577);
and U21004 (N_21004,N_20708,N_20583);
nor U21005 (N_21005,N_20949,N_20457);
and U21006 (N_21006,N_20839,N_20900);
xor U21007 (N_21007,N_20984,N_20827);
and U21008 (N_21008,N_20719,N_20526);
or U21009 (N_21009,N_20615,N_20463);
xnor U21010 (N_21010,N_20845,N_20512);
xnor U21011 (N_21011,N_20901,N_20429);
nor U21012 (N_21012,N_20649,N_20933);
or U21013 (N_21013,N_20724,N_20702);
xor U21014 (N_21014,N_20689,N_20776);
or U21015 (N_21015,N_20444,N_20936);
and U21016 (N_21016,N_20796,N_20622);
xor U21017 (N_21017,N_20482,N_20992);
or U21018 (N_21018,N_20611,N_20728);
nand U21019 (N_21019,N_20767,N_20939);
and U21020 (N_21020,N_20645,N_20422);
or U21021 (N_21021,N_20935,N_20772);
nor U21022 (N_21022,N_20671,N_20748);
nand U21023 (N_21023,N_20676,N_20911);
xor U21024 (N_21024,N_20913,N_20674);
or U21025 (N_21025,N_20856,N_20417);
nand U21026 (N_21026,N_20882,N_20514);
xnor U21027 (N_21027,N_20407,N_20754);
or U21028 (N_21028,N_20757,N_20995);
or U21029 (N_21029,N_20559,N_20918);
xnor U21030 (N_21030,N_20730,N_20453);
or U21031 (N_21031,N_20535,N_20779);
nor U21032 (N_21032,N_20642,N_20921);
nor U21033 (N_21033,N_20541,N_20553);
nand U21034 (N_21034,N_20979,N_20928);
nand U21035 (N_21035,N_20519,N_20894);
nand U21036 (N_21036,N_20993,N_20937);
nand U21037 (N_21037,N_20833,N_20585);
xor U21038 (N_21038,N_20687,N_20923);
and U21039 (N_21039,N_20785,N_20692);
or U21040 (N_21040,N_20626,N_20634);
xor U21041 (N_21041,N_20837,N_20743);
nand U21042 (N_21042,N_20737,N_20638);
nor U21043 (N_21043,N_20847,N_20771);
xnor U21044 (N_21044,N_20840,N_20443);
nand U21045 (N_21045,N_20711,N_20467);
and U21046 (N_21046,N_20665,N_20545);
and U21047 (N_21047,N_20852,N_20732);
and U21048 (N_21048,N_20828,N_20486);
or U21049 (N_21049,N_20694,N_20400);
and U21050 (N_21050,N_20706,N_20814);
nand U21051 (N_21051,N_20838,N_20784);
nor U21052 (N_21052,N_20974,N_20798);
or U21053 (N_21053,N_20720,N_20770);
or U21054 (N_21054,N_20925,N_20616);
nor U21055 (N_21055,N_20549,N_20922);
nand U21056 (N_21056,N_20860,N_20903);
nand U21057 (N_21057,N_20971,N_20441);
and U21058 (N_21058,N_20880,N_20461);
or U21059 (N_21059,N_20803,N_20774);
nand U21060 (N_21060,N_20862,N_20945);
nand U21061 (N_21061,N_20801,N_20603);
or U21062 (N_21062,N_20538,N_20758);
or U21063 (N_21063,N_20663,N_20744);
xnor U21064 (N_21064,N_20909,N_20656);
and U21065 (N_21065,N_20605,N_20517);
xor U21066 (N_21066,N_20607,N_20496);
nor U21067 (N_21067,N_20419,N_20973);
nor U21068 (N_21068,N_20818,N_20652);
or U21069 (N_21069,N_20968,N_20899);
nor U21070 (N_21070,N_20588,N_20410);
nand U21071 (N_21071,N_20586,N_20418);
nand U21072 (N_21072,N_20520,N_20910);
xnor U21073 (N_21073,N_20953,N_20980);
or U21074 (N_21074,N_20853,N_20946);
and U21075 (N_21075,N_20815,N_20963);
nand U21076 (N_21076,N_20734,N_20797);
or U21077 (N_21077,N_20842,N_20879);
or U21078 (N_21078,N_20411,N_20749);
and U21079 (N_21079,N_20836,N_20620);
and U21080 (N_21080,N_20917,N_20602);
nand U21081 (N_21081,N_20807,N_20460);
nand U21082 (N_21082,N_20491,N_20502);
xnor U21083 (N_21083,N_20983,N_20637);
or U21084 (N_21084,N_20769,N_20621);
or U21085 (N_21085,N_20695,N_20760);
xor U21086 (N_21086,N_20431,N_20644);
xnor U21087 (N_21087,N_20717,N_20698);
or U21088 (N_21088,N_20488,N_20716);
nand U21089 (N_21089,N_20686,N_20670);
or U21090 (N_21090,N_20926,N_20497);
xor U21091 (N_21091,N_20557,N_20599);
nor U21092 (N_21092,N_20843,N_20568);
or U21093 (N_21093,N_20906,N_20857);
xnor U21094 (N_21094,N_20793,N_20693);
nor U21095 (N_21095,N_20948,N_20891);
nor U21096 (N_21096,N_20966,N_20524);
and U21097 (N_21097,N_20532,N_20594);
nor U21098 (N_21098,N_20863,N_20556);
nor U21099 (N_21099,N_20989,N_20576);
or U21100 (N_21100,N_20485,N_20952);
and U21101 (N_21101,N_20528,N_20941);
nand U21102 (N_21102,N_20614,N_20484);
nand U21103 (N_21103,N_20783,N_20490);
nor U21104 (N_21104,N_20503,N_20624);
or U21105 (N_21105,N_20550,N_20592);
and U21106 (N_21106,N_20756,N_20629);
and U21107 (N_21107,N_20481,N_20878);
or U21108 (N_21108,N_20835,N_20780);
or U21109 (N_21109,N_20747,N_20721);
and U21110 (N_21110,N_20961,N_20679);
nor U21111 (N_21111,N_20546,N_20709);
or U21112 (N_21112,N_20628,N_20864);
nor U21113 (N_21113,N_20813,N_20883);
nand U21114 (N_21114,N_20867,N_20534);
or U21115 (N_21115,N_20570,N_20572);
or U21116 (N_21116,N_20792,N_20582);
and U21117 (N_21117,N_20672,N_20782);
nor U21118 (N_21118,N_20499,N_20691);
and U21119 (N_21119,N_20817,N_20950);
nor U21120 (N_21120,N_20487,N_20977);
nor U21121 (N_21121,N_20723,N_20483);
and U21122 (N_21122,N_20822,N_20808);
nor U21123 (N_21123,N_20661,N_20507);
nand U21124 (N_21124,N_20439,N_20960);
xor U21125 (N_21125,N_20425,N_20537);
xnor U21126 (N_21126,N_20947,N_20738);
xnor U21127 (N_21127,N_20868,N_20580);
or U21128 (N_21128,N_20998,N_20877);
nand U21129 (N_21129,N_20462,N_20861);
nor U21130 (N_21130,N_20428,N_20456);
nor U21131 (N_21131,N_20531,N_20521);
or U21132 (N_21132,N_20561,N_20908);
and U21133 (N_21133,N_20573,N_20420);
xor U21134 (N_21134,N_20632,N_20625);
nand U21135 (N_21135,N_20449,N_20543);
nand U21136 (N_21136,N_20454,N_20606);
and U21137 (N_21137,N_20493,N_20646);
nor U21138 (N_21138,N_20802,N_20981);
nand U21139 (N_21139,N_20970,N_20612);
xor U21140 (N_21140,N_20508,N_20562);
xor U21141 (N_21141,N_20701,N_20834);
and U21142 (N_21142,N_20819,N_20763);
nand U21143 (N_21143,N_20700,N_20608);
xnor U21144 (N_21144,N_20731,N_20405);
xor U21145 (N_21145,N_20871,N_20904);
or U21146 (N_21146,N_20951,N_20495);
or U21147 (N_21147,N_20450,N_20434);
xor U21148 (N_21148,N_20563,N_20773);
and U21149 (N_21149,N_20500,N_20492);
xor U21150 (N_21150,N_20799,N_20551);
nor U21151 (N_21151,N_20722,N_20542);
nor U21152 (N_21152,N_20832,N_20437);
nand U21153 (N_21153,N_20962,N_20826);
or U21154 (N_21154,N_20712,N_20859);
nand U21155 (N_21155,N_20511,N_20848);
or U21156 (N_21156,N_20858,N_20846);
nand U21157 (N_21157,N_20750,N_20574);
and U21158 (N_21158,N_20618,N_20787);
or U21159 (N_21159,N_20725,N_20735);
xor U21160 (N_21160,N_20768,N_20727);
and U21161 (N_21161,N_20416,N_20682);
and U21162 (N_21162,N_20759,N_20681);
nor U21163 (N_21163,N_20726,N_20515);
xor U21164 (N_21164,N_20794,N_20912);
nor U21165 (N_21165,N_20558,N_20751);
or U21166 (N_21166,N_20965,N_20470);
nand U21167 (N_21167,N_20778,N_20413);
or U21168 (N_21168,N_20955,N_20504);
nand U21169 (N_21169,N_20930,N_20897);
nand U21170 (N_21170,N_20775,N_20591);
nor U21171 (N_21171,N_20786,N_20890);
and U21172 (N_21172,N_20421,N_20884);
nand U21173 (N_21173,N_20680,N_20990);
nor U21174 (N_21174,N_20885,N_20736);
xnor U21175 (N_21175,N_20844,N_20564);
and U21176 (N_21176,N_20408,N_20442);
or U21177 (N_21177,N_20433,N_20660);
or U21178 (N_21178,N_20565,N_20888);
xnor U21179 (N_21179,N_20659,N_20469);
nor U21180 (N_21180,N_20954,N_20889);
nor U21181 (N_21181,N_20886,N_20544);
xnor U21182 (N_21182,N_20975,N_20790);
nor U21183 (N_21183,N_20409,N_20423);
or U21184 (N_21184,N_20403,N_20655);
nor U21185 (N_21185,N_20445,N_20639);
xor U21186 (N_21186,N_20875,N_20667);
nor U21187 (N_21187,N_20942,N_20851);
and U21188 (N_21188,N_20657,N_20539);
nand U21189 (N_21189,N_20745,N_20873);
or U21190 (N_21190,N_20959,N_20617);
or U21191 (N_21191,N_20478,N_20536);
or U21192 (N_21192,N_20458,N_20587);
nor U21193 (N_21193,N_20956,N_20406);
and U21194 (N_21194,N_20677,N_20887);
or U21195 (N_21195,N_20424,N_20619);
nor U21196 (N_21196,N_20505,N_20976);
and U21197 (N_21197,N_20964,N_20569);
or U21198 (N_21198,N_20865,N_20440);
nand U21199 (N_21199,N_20739,N_20929);
nand U21200 (N_21200,N_20554,N_20464);
nand U21201 (N_21201,N_20755,N_20829);
xnor U21202 (N_21202,N_20713,N_20579);
and U21203 (N_21203,N_20881,N_20566);
and U21204 (N_21204,N_20489,N_20506);
xnor U21205 (N_21205,N_20402,N_20943);
nor U21206 (N_21206,N_20631,N_20468);
or U21207 (N_21207,N_20525,N_20841);
nor U21208 (N_21208,N_20972,N_20651);
and U21209 (N_21209,N_20893,N_20824);
and U21210 (N_21210,N_20601,N_20791);
nor U21211 (N_21211,N_20916,N_20675);
and U21212 (N_21212,N_20648,N_20789);
nand U21213 (N_21213,N_20640,N_20704);
or U21214 (N_21214,N_20872,N_20811);
and U21215 (N_21215,N_20560,N_20613);
nand U21216 (N_21216,N_20684,N_20914);
xor U21217 (N_21217,N_20806,N_20430);
or U21218 (N_21218,N_20690,N_20664);
nor U21219 (N_21219,N_20915,N_20596);
nor U21220 (N_21220,N_20633,N_20927);
xor U21221 (N_21221,N_20494,N_20934);
and U21222 (N_21222,N_20666,N_20940);
or U21223 (N_21223,N_20969,N_20623);
or U21224 (N_21224,N_20471,N_20764);
or U21225 (N_21225,N_20635,N_20752);
nor U21226 (N_21226,N_20938,N_20527);
nand U21227 (N_21227,N_20533,N_20510);
nand U21228 (N_21228,N_20435,N_20830);
nor U21229 (N_21229,N_20477,N_20412);
nor U21230 (N_21230,N_20513,N_20597);
or U21231 (N_21231,N_20475,N_20427);
and U21232 (N_21232,N_20994,N_20473);
and U21233 (N_21233,N_20476,N_20697);
and U21234 (N_21234,N_20555,N_20781);
nand U21235 (N_21235,N_20523,N_20991);
or U21236 (N_21236,N_20459,N_20590);
nand U21237 (N_21237,N_20761,N_20448);
nor U21238 (N_21238,N_20850,N_20571);
xnor U21239 (N_21239,N_20825,N_20501);
nor U21240 (N_21240,N_20831,N_20600);
or U21241 (N_21241,N_20997,N_20465);
nand U21242 (N_21242,N_20436,N_20641);
or U21243 (N_21243,N_20540,N_20474);
nand U21244 (N_21244,N_20729,N_20820);
or U21245 (N_21245,N_20907,N_20683);
nor U21246 (N_21246,N_20924,N_20809);
nand U21247 (N_21247,N_20876,N_20703);
nor U21248 (N_21248,N_20788,N_20714);
and U21249 (N_21249,N_20892,N_20999);
nand U21250 (N_21250,N_20447,N_20931);
xor U21251 (N_21251,N_20895,N_20740);
and U21252 (N_21252,N_20548,N_20581);
and U21253 (N_21253,N_20777,N_20518);
xor U21254 (N_21254,N_20530,N_20766);
and U21255 (N_21255,N_20905,N_20987);
nor U21256 (N_21256,N_20707,N_20401);
or U21257 (N_21257,N_20715,N_20647);
xor U21258 (N_21258,N_20746,N_20627);
and U21259 (N_21259,N_20438,N_20958);
or U21260 (N_21260,N_20636,N_20414);
xor U21261 (N_21261,N_20733,N_20604);
and U21262 (N_21262,N_20896,N_20765);
and U21263 (N_21263,N_20699,N_20529);
and U21264 (N_21264,N_20710,N_20451);
nand U21265 (N_21265,N_20944,N_20654);
xnor U21266 (N_21266,N_20567,N_20718);
nand U21267 (N_21267,N_20452,N_20996);
and U21268 (N_21268,N_20653,N_20985);
nor U21269 (N_21269,N_20432,N_20522);
nor U21270 (N_21270,N_20821,N_20595);
or U21271 (N_21271,N_20967,N_20920);
nor U21272 (N_21272,N_20480,N_20753);
nor U21273 (N_21273,N_20696,N_20804);
and U21274 (N_21274,N_20705,N_20742);
xnor U21275 (N_21275,N_20849,N_20609);
nand U21276 (N_21276,N_20552,N_20472);
nor U21277 (N_21277,N_20662,N_20610);
xnor U21278 (N_21278,N_20650,N_20578);
xnor U21279 (N_21279,N_20455,N_20669);
nand U21280 (N_21280,N_20812,N_20982);
nand U21281 (N_21281,N_20673,N_20823);
xor U21282 (N_21282,N_20630,N_20584);
nor U21283 (N_21283,N_20816,N_20466);
nand U21284 (N_21284,N_20426,N_20957);
xor U21285 (N_21285,N_20898,N_20795);
nand U21286 (N_21286,N_20870,N_20589);
or U21287 (N_21287,N_20762,N_20986);
nor U21288 (N_21288,N_20988,N_20547);
and U21289 (N_21289,N_20866,N_20404);
nor U21290 (N_21290,N_20685,N_20479);
or U21291 (N_21291,N_20446,N_20678);
and U21292 (N_21292,N_20658,N_20855);
and U21293 (N_21293,N_20668,N_20978);
and U21294 (N_21294,N_20805,N_20854);
or U21295 (N_21295,N_20498,N_20598);
nor U21296 (N_21296,N_20688,N_20932);
or U21297 (N_21297,N_20810,N_20509);
or U21298 (N_21298,N_20741,N_20516);
nand U21299 (N_21299,N_20874,N_20575);
or U21300 (N_21300,N_20892,N_20610);
or U21301 (N_21301,N_20640,N_20494);
nor U21302 (N_21302,N_20480,N_20886);
or U21303 (N_21303,N_20784,N_20673);
nand U21304 (N_21304,N_20579,N_20408);
xor U21305 (N_21305,N_20816,N_20489);
xnor U21306 (N_21306,N_20715,N_20841);
or U21307 (N_21307,N_20508,N_20521);
or U21308 (N_21308,N_20655,N_20556);
xnor U21309 (N_21309,N_20554,N_20631);
and U21310 (N_21310,N_20709,N_20668);
nor U21311 (N_21311,N_20570,N_20886);
xnor U21312 (N_21312,N_20595,N_20786);
xnor U21313 (N_21313,N_20987,N_20516);
or U21314 (N_21314,N_20571,N_20794);
or U21315 (N_21315,N_20417,N_20655);
nor U21316 (N_21316,N_20779,N_20437);
nor U21317 (N_21317,N_20891,N_20505);
or U21318 (N_21318,N_20566,N_20762);
nand U21319 (N_21319,N_20776,N_20753);
nand U21320 (N_21320,N_20684,N_20971);
or U21321 (N_21321,N_20678,N_20434);
nand U21322 (N_21322,N_20829,N_20625);
nand U21323 (N_21323,N_20938,N_20655);
and U21324 (N_21324,N_20892,N_20469);
nor U21325 (N_21325,N_20753,N_20999);
xor U21326 (N_21326,N_20474,N_20669);
nand U21327 (N_21327,N_20922,N_20904);
or U21328 (N_21328,N_20570,N_20901);
xor U21329 (N_21329,N_20605,N_20899);
and U21330 (N_21330,N_20805,N_20915);
nand U21331 (N_21331,N_20703,N_20791);
and U21332 (N_21332,N_20507,N_20428);
nand U21333 (N_21333,N_20579,N_20795);
or U21334 (N_21334,N_20727,N_20878);
nor U21335 (N_21335,N_20449,N_20903);
nor U21336 (N_21336,N_20421,N_20622);
xnor U21337 (N_21337,N_20568,N_20675);
nand U21338 (N_21338,N_20880,N_20596);
nor U21339 (N_21339,N_20868,N_20715);
nor U21340 (N_21340,N_20955,N_20480);
or U21341 (N_21341,N_20623,N_20544);
xnor U21342 (N_21342,N_20900,N_20668);
and U21343 (N_21343,N_20806,N_20816);
nor U21344 (N_21344,N_20890,N_20974);
xor U21345 (N_21345,N_20512,N_20414);
or U21346 (N_21346,N_20866,N_20418);
nor U21347 (N_21347,N_20927,N_20967);
nand U21348 (N_21348,N_20701,N_20680);
and U21349 (N_21349,N_20732,N_20588);
and U21350 (N_21350,N_20986,N_20953);
or U21351 (N_21351,N_20912,N_20666);
xor U21352 (N_21352,N_20543,N_20682);
or U21353 (N_21353,N_20930,N_20505);
nor U21354 (N_21354,N_20541,N_20924);
or U21355 (N_21355,N_20817,N_20583);
xnor U21356 (N_21356,N_20651,N_20647);
or U21357 (N_21357,N_20560,N_20740);
nand U21358 (N_21358,N_20423,N_20505);
nand U21359 (N_21359,N_20587,N_20734);
xnor U21360 (N_21360,N_20791,N_20401);
or U21361 (N_21361,N_20875,N_20523);
nand U21362 (N_21362,N_20713,N_20959);
nor U21363 (N_21363,N_20492,N_20955);
and U21364 (N_21364,N_20524,N_20660);
nand U21365 (N_21365,N_20550,N_20643);
nand U21366 (N_21366,N_20530,N_20940);
nor U21367 (N_21367,N_20720,N_20754);
and U21368 (N_21368,N_20939,N_20408);
and U21369 (N_21369,N_20550,N_20744);
or U21370 (N_21370,N_20707,N_20581);
xor U21371 (N_21371,N_20472,N_20689);
nand U21372 (N_21372,N_20846,N_20532);
nor U21373 (N_21373,N_20702,N_20459);
nand U21374 (N_21374,N_20732,N_20707);
nand U21375 (N_21375,N_20564,N_20738);
and U21376 (N_21376,N_20750,N_20549);
xor U21377 (N_21377,N_20697,N_20600);
nor U21378 (N_21378,N_20823,N_20605);
or U21379 (N_21379,N_20910,N_20594);
or U21380 (N_21380,N_20757,N_20791);
and U21381 (N_21381,N_20972,N_20642);
nor U21382 (N_21382,N_20961,N_20882);
nand U21383 (N_21383,N_20956,N_20623);
xor U21384 (N_21384,N_20528,N_20576);
and U21385 (N_21385,N_20828,N_20767);
nor U21386 (N_21386,N_20971,N_20462);
or U21387 (N_21387,N_20425,N_20684);
and U21388 (N_21388,N_20821,N_20959);
and U21389 (N_21389,N_20493,N_20867);
xnor U21390 (N_21390,N_20883,N_20405);
nor U21391 (N_21391,N_20619,N_20539);
nand U21392 (N_21392,N_20701,N_20539);
nand U21393 (N_21393,N_20753,N_20649);
xor U21394 (N_21394,N_20788,N_20635);
nor U21395 (N_21395,N_20770,N_20595);
or U21396 (N_21396,N_20748,N_20914);
and U21397 (N_21397,N_20827,N_20773);
xnor U21398 (N_21398,N_20917,N_20977);
nand U21399 (N_21399,N_20832,N_20746);
or U21400 (N_21400,N_20485,N_20910);
xor U21401 (N_21401,N_20610,N_20956);
nand U21402 (N_21402,N_20858,N_20768);
nor U21403 (N_21403,N_20946,N_20689);
nor U21404 (N_21404,N_20701,N_20854);
and U21405 (N_21405,N_20674,N_20666);
nand U21406 (N_21406,N_20657,N_20431);
xor U21407 (N_21407,N_20539,N_20454);
nand U21408 (N_21408,N_20452,N_20942);
xnor U21409 (N_21409,N_20620,N_20977);
or U21410 (N_21410,N_20554,N_20717);
xor U21411 (N_21411,N_20866,N_20909);
nor U21412 (N_21412,N_20761,N_20727);
nor U21413 (N_21413,N_20784,N_20579);
or U21414 (N_21414,N_20845,N_20500);
nor U21415 (N_21415,N_20939,N_20929);
nor U21416 (N_21416,N_20583,N_20662);
or U21417 (N_21417,N_20712,N_20847);
xor U21418 (N_21418,N_20511,N_20828);
nand U21419 (N_21419,N_20711,N_20659);
xnor U21420 (N_21420,N_20640,N_20403);
nand U21421 (N_21421,N_20846,N_20753);
or U21422 (N_21422,N_20493,N_20556);
nor U21423 (N_21423,N_20752,N_20446);
xor U21424 (N_21424,N_20918,N_20940);
xor U21425 (N_21425,N_20908,N_20909);
xor U21426 (N_21426,N_20623,N_20441);
or U21427 (N_21427,N_20902,N_20603);
nor U21428 (N_21428,N_20894,N_20596);
nand U21429 (N_21429,N_20590,N_20661);
nand U21430 (N_21430,N_20700,N_20887);
nor U21431 (N_21431,N_20826,N_20983);
xor U21432 (N_21432,N_20755,N_20498);
xnor U21433 (N_21433,N_20540,N_20475);
xnor U21434 (N_21434,N_20883,N_20470);
nor U21435 (N_21435,N_20457,N_20443);
xnor U21436 (N_21436,N_20415,N_20556);
nor U21437 (N_21437,N_20886,N_20433);
nor U21438 (N_21438,N_20451,N_20934);
or U21439 (N_21439,N_20693,N_20862);
nand U21440 (N_21440,N_20795,N_20969);
xor U21441 (N_21441,N_20908,N_20528);
xor U21442 (N_21442,N_20888,N_20750);
or U21443 (N_21443,N_20533,N_20927);
nand U21444 (N_21444,N_20914,N_20486);
nor U21445 (N_21445,N_20980,N_20867);
xnor U21446 (N_21446,N_20736,N_20453);
nor U21447 (N_21447,N_20733,N_20559);
nand U21448 (N_21448,N_20763,N_20938);
and U21449 (N_21449,N_20573,N_20722);
or U21450 (N_21450,N_20704,N_20939);
xor U21451 (N_21451,N_20650,N_20475);
and U21452 (N_21452,N_20892,N_20932);
or U21453 (N_21453,N_20565,N_20403);
and U21454 (N_21454,N_20706,N_20405);
or U21455 (N_21455,N_20435,N_20729);
nor U21456 (N_21456,N_20578,N_20455);
xnor U21457 (N_21457,N_20955,N_20712);
or U21458 (N_21458,N_20496,N_20535);
xnor U21459 (N_21459,N_20574,N_20438);
nor U21460 (N_21460,N_20836,N_20923);
nand U21461 (N_21461,N_20873,N_20458);
nor U21462 (N_21462,N_20410,N_20634);
nand U21463 (N_21463,N_20592,N_20826);
or U21464 (N_21464,N_20456,N_20823);
or U21465 (N_21465,N_20433,N_20867);
nor U21466 (N_21466,N_20660,N_20620);
nor U21467 (N_21467,N_20884,N_20982);
nor U21468 (N_21468,N_20589,N_20885);
xnor U21469 (N_21469,N_20892,N_20813);
xor U21470 (N_21470,N_20420,N_20423);
or U21471 (N_21471,N_20451,N_20731);
nor U21472 (N_21472,N_20694,N_20900);
and U21473 (N_21473,N_20836,N_20809);
or U21474 (N_21474,N_20816,N_20758);
and U21475 (N_21475,N_20984,N_20663);
nand U21476 (N_21476,N_20753,N_20980);
nor U21477 (N_21477,N_20459,N_20735);
or U21478 (N_21478,N_20709,N_20455);
nand U21479 (N_21479,N_20559,N_20424);
and U21480 (N_21480,N_20961,N_20809);
nor U21481 (N_21481,N_20672,N_20450);
xnor U21482 (N_21482,N_20965,N_20444);
or U21483 (N_21483,N_20412,N_20475);
nor U21484 (N_21484,N_20647,N_20484);
nand U21485 (N_21485,N_20634,N_20533);
nand U21486 (N_21486,N_20803,N_20438);
and U21487 (N_21487,N_20949,N_20498);
or U21488 (N_21488,N_20838,N_20820);
or U21489 (N_21489,N_20623,N_20633);
and U21490 (N_21490,N_20666,N_20968);
and U21491 (N_21491,N_20683,N_20816);
nor U21492 (N_21492,N_20913,N_20406);
nand U21493 (N_21493,N_20933,N_20740);
or U21494 (N_21494,N_20868,N_20818);
nand U21495 (N_21495,N_20560,N_20680);
nor U21496 (N_21496,N_20728,N_20400);
and U21497 (N_21497,N_20509,N_20551);
xnor U21498 (N_21498,N_20937,N_20680);
nand U21499 (N_21499,N_20797,N_20921);
xnor U21500 (N_21500,N_20772,N_20811);
nand U21501 (N_21501,N_20618,N_20736);
and U21502 (N_21502,N_20787,N_20443);
nand U21503 (N_21503,N_20413,N_20544);
nand U21504 (N_21504,N_20969,N_20641);
and U21505 (N_21505,N_20550,N_20680);
xnor U21506 (N_21506,N_20538,N_20565);
or U21507 (N_21507,N_20751,N_20658);
xor U21508 (N_21508,N_20708,N_20991);
or U21509 (N_21509,N_20968,N_20508);
xor U21510 (N_21510,N_20540,N_20995);
and U21511 (N_21511,N_20891,N_20974);
nor U21512 (N_21512,N_20900,N_20569);
and U21513 (N_21513,N_20688,N_20867);
xor U21514 (N_21514,N_20464,N_20409);
or U21515 (N_21515,N_20908,N_20935);
nor U21516 (N_21516,N_20682,N_20934);
and U21517 (N_21517,N_20532,N_20446);
or U21518 (N_21518,N_20519,N_20951);
and U21519 (N_21519,N_20416,N_20665);
xnor U21520 (N_21520,N_20548,N_20771);
xnor U21521 (N_21521,N_20863,N_20516);
nand U21522 (N_21522,N_20666,N_20453);
nor U21523 (N_21523,N_20736,N_20875);
xor U21524 (N_21524,N_20463,N_20687);
xor U21525 (N_21525,N_20977,N_20669);
nor U21526 (N_21526,N_20584,N_20909);
nor U21527 (N_21527,N_20792,N_20617);
and U21528 (N_21528,N_20478,N_20756);
and U21529 (N_21529,N_20956,N_20944);
nor U21530 (N_21530,N_20552,N_20648);
and U21531 (N_21531,N_20751,N_20866);
nand U21532 (N_21532,N_20570,N_20560);
nor U21533 (N_21533,N_20427,N_20905);
xor U21534 (N_21534,N_20721,N_20484);
and U21535 (N_21535,N_20769,N_20732);
nand U21536 (N_21536,N_20661,N_20435);
nor U21537 (N_21537,N_20588,N_20977);
xnor U21538 (N_21538,N_20910,N_20633);
nor U21539 (N_21539,N_20525,N_20717);
nand U21540 (N_21540,N_20573,N_20941);
nand U21541 (N_21541,N_20631,N_20649);
and U21542 (N_21542,N_20796,N_20433);
nand U21543 (N_21543,N_20629,N_20498);
nor U21544 (N_21544,N_20455,N_20494);
nor U21545 (N_21545,N_20400,N_20726);
nand U21546 (N_21546,N_20942,N_20516);
xnor U21547 (N_21547,N_20816,N_20866);
xnor U21548 (N_21548,N_20703,N_20509);
and U21549 (N_21549,N_20618,N_20872);
nor U21550 (N_21550,N_20605,N_20902);
or U21551 (N_21551,N_20543,N_20761);
nor U21552 (N_21552,N_20910,N_20727);
nand U21553 (N_21553,N_20946,N_20488);
and U21554 (N_21554,N_20478,N_20739);
xor U21555 (N_21555,N_20464,N_20556);
xor U21556 (N_21556,N_20894,N_20612);
and U21557 (N_21557,N_20521,N_20945);
and U21558 (N_21558,N_20506,N_20662);
or U21559 (N_21559,N_20573,N_20667);
and U21560 (N_21560,N_20699,N_20961);
xor U21561 (N_21561,N_20865,N_20767);
xor U21562 (N_21562,N_20540,N_20441);
and U21563 (N_21563,N_20592,N_20724);
nand U21564 (N_21564,N_20857,N_20659);
nor U21565 (N_21565,N_20733,N_20513);
nor U21566 (N_21566,N_20676,N_20541);
xnor U21567 (N_21567,N_20947,N_20892);
and U21568 (N_21568,N_20797,N_20408);
nand U21569 (N_21569,N_20491,N_20510);
nand U21570 (N_21570,N_20709,N_20417);
xnor U21571 (N_21571,N_20620,N_20828);
nand U21572 (N_21572,N_20733,N_20914);
xor U21573 (N_21573,N_20672,N_20853);
nand U21574 (N_21574,N_20713,N_20636);
and U21575 (N_21575,N_20688,N_20695);
xnor U21576 (N_21576,N_20977,N_20582);
and U21577 (N_21577,N_20812,N_20553);
nand U21578 (N_21578,N_20787,N_20478);
or U21579 (N_21579,N_20961,N_20848);
or U21580 (N_21580,N_20725,N_20878);
or U21581 (N_21581,N_20445,N_20763);
or U21582 (N_21582,N_20766,N_20838);
nor U21583 (N_21583,N_20554,N_20433);
nand U21584 (N_21584,N_20520,N_20610);
xor U21585 (N_21585,N_20535,N_20814);
or U21586 (N_21586,N_20810,N_20552);
nor U21587 (N_21587,N_20447,N_20517);
and U21588 (N_21588,N_20638,N_20927);
or U21589 (N_21589,N_20708,N_20959);
or U21590 (N_21590,N_20415,N_20529);
and U21591 (N_21591,N_20414,N_20790);
xor U21592 (N_21592,N_20921,N_20528);
xnor U21593 (N_21593,N_20872,N_20714);
nand U21594 (N_21594,N_20432,N_20934);
nor U21595 (N_21595,N_20412,N_20870);
nor U21596 (N_21596,N_20839,N_20457);
nor U21597 (N_21597,N_20779,N_20835);
xnor U21598 (N_21598,N_20440,N_20439);
nand U21599 (N_21599,N_20884,N_20515);
or U21600 (N_21600,N_21195,N_21251);
xnor U21601 (N_21601,N_21391,N_21530);
or U21602 (N_21602,N_21449,N_21159);
nand U21603 (N_21603,N_21241,N_21470);
nand U21604 (N_21604,N_21343,N_21539);
and U21605 (N_21605,N_21411,N_21002);
and U21606 (N_21606,N_21192,N_21074);
nand U21607 (N_21607,N_21542,N_21441);
nor U21608 (N_21608,N_21164,N_21418);
or U21609 (N_21609,N_21124,N_21131);
or U21610 (N_21610,N_21256,N_21357);
nand U21611 (N_21611,N_21080,N_21452);
or U21612 (N_21612,N_21171,N_21030);
and U21613 (N_21613,N_21584,N_21060);
xor U21614 (N_21614,N_21176,N_21172);
and U21615 (N_21615,N_21269,N_21005);
xnor U21616 (N_21616,N_21268,N_21011);
nand U21617 (N_21617,N_21087,N_21336);
or U21618 (N_21618,N_21404,N_21578);
nand U21619 (N_21619,N_21358,N_21324);
and U21620 (N_21620,N_21346,N_21473);
and U21621 (N_21621,N_21254,N_21147);
and U21622 (N_21622,N_21550,N_21496);
or U21623 (N_21623,N_21423,N_21055);
xnor U21624 (N_21624,N_21231,N_21194);
xnor U21625 (N_21625,N_21386,N_21430);
and U21626 (N_21626,N_21039,N_21564);
or U21627 (N_21627,N_21599,N_21144);
xor U21628 (N_21628,N_21295,N_21491);
nand U21629 (N_21629,N_21366,N_21260);
xor U21630 (N_21630,N_21058,N_21132);
nand U21631 (N_21631,N_21092,N_21137);
and U21632 (N_21632,N_21454,N_21403);
and U21633 (N_21633,N_21553,N_21013);
or U21634 (N_21634,N_21433,N_21414);
or U21635 (N_21635,N_21024,N_21401);
nand U21636 (N_21636,N_21279,N_21071);
xor U21637 (N_21637,N_21179,N_21489);
nor U21638 (N_21638,N_21512,N_21543);
and U21639 (N_21639,N_21243,N_21010);
and U21640 (N_21640,N_21204,N_21227);
xnor U21641 (N_21641,N_21276,N_21363);
and U21642 (N_21642,N_21486,N_21218);
xor U21643 (N_21643,N_21421,N_21582);
xnor U21644 (N_21644,N_21485,N_21196);
and U21645 (N_21645,N_21151,N_21261);
xor U21646 (N_21646,N_21133,N_21238);
and U21647 (N_21647,N_21375,N_21077);
and U21648 (N_21648,N_21432,N_21163);
nor U21649 (N_21649,N_21275,N_21367);
or U21650 (N_21650,N_21004,N_21001);
xnor U21651 (N_21651,N_21398,N_21368);
nand U21652 (N_21652,N_21580,N_21347);
nand U21653 (N_21653,N_21424,N_21208);
and U21654 (N_21654,N_21081,N_21395);
xor U21655 (N_21655,N_21157,N_21465);
and U21656 (N_21656,N_21456,N_21116);
nand U21657 (N_21657,N_21146,N_21558);
or U21658 (N_21658,N_21323,N_21112);
nand U21659 (N_21659,N_21337,N_21283);
or U21660 (N_21660,N_21334,N_21222);
and U21661 (N_21661,N_21274,N_21221);
nand U21662 (N_21662,N_21228,N_21447);
nand U21663 (N_21663,N_21211,N_21242);
or U21664 (N_21664,N_21101,N_21119);
or U21665 (N_21665,N_21481,N_21528);
or U21666 (N_21666,N_21202,N_21108);
nand U21667 (N_21667,N_21448,N_21301);
and U21668 (N_21668,N_21174,N_21434);
nor U21669 (N_21669,N_21115,N_21380);
or U21670 (N_21670,N_21427,N_21145);
nand U21671 (N_21671,N_21583,N_21259);
and U21672 (N_21672,N_21237,N_21096);
nor U21673 (N_21673,N_21110,N_21422);
nand U21674 (N_21674,N_21289,N_21351);
xor U21675 (N_21675,N_21111,N_21245);
nand U21676 (N_21676,N_21502,N_21170);
xnor U21677 (N_21677,N_21050,N_21574);
nand U21678 (N_21678,N_21405,N_21105);
or U21679 (N_21679,N_21420,N_21069);
and U21680 (N_21680,N_21464,N_21579);
and U21681 (N_21681,N_21244,N_21271);
nand U21682 (N_21682,N_21526,N_21522);
nand U21683 (N_21683,N_21498,N_21278);
nor U21684 (N_21684,N_21135,N_21122);
nor U21685 (N_21685,N_21349,N_21199);
xnor U21686 (N_21686,N_21121,N_21296);
or U21687 (N_21687,N_21381,N_21136);
or U21688 (N_21688,N_21044,N_21090);
and U21689 (N_21689,N_21478,N_21355);
or U21690 (N_21690,N_21288,N_21093);
and U21691 (N_21691,N_21045,N_21314);
and U21692 (N_21692,N_21472,N_21240);
and U21693 (N_21693,N_21047,N_21359);
nor U21694 (N_21694,N_21460,N_21061);
and U21695 (N_21695,N_21210,N_21340);
xnor U21696 (N_21696,N_21161,N_21178);
xor U21697 (N_21697,N_21258,N_21138);
nor U21698 (N_21698,N_21562,N_21372);
and U21699 (N_21699,N_21419,N_21500);
and U21700 (N_21700,N_21028,N_21309);
and U21701 (N_21701,N_21376,N_21064);
nor U21702 (N_21702,N_21225,N_21130);
and U21703 (N_21703,N_21142,N_21057);
nand U21704 (N_21704,N_21223,N_21262);
nor U21705 (N_21705,N_21306,N_21284);
nor U21706 (N_21706,N_21467,N_21286);
nand U21707 (N_21707,N_21361,N_21330);
nand U21708 (N_21708,N_21084,N_21000);
and U21709 (N_21709,N_21070,N_21480);
xor U21710 (N_21710,N_21073,N_21117);
nor U21711 (N_21711,N_21017,N_21120);
xor U21712 (N_21712,N_21495,N_21206);
nor U21713 (N_21713,N_21033,N_21444);
xnor U21714 (N_21714,N_21139,N_21463);
nand U21715 (N_21715,N_21127,N_21352);
or U21716 (N_21716,N_21134,N_21402);
xnor U21717 (N_21717,N_21152,N_21513);
nor U21718 (N_21718,N_21338,N_21332);
nor U21719 (N_21719,N_21325,N_21400);
nor U21720 (N_21720,N_21319,N_21577);
nor U21721 (N_21721,N_21248,N_21003);
nor U21722 (N_21722,N_21183,N_21345);
nand U21723 (N_21723,N_21415,N_21075);
nor U21724 (N_21724,N_21287,N_21506);
or U21725 (N_21725,N_21531,N_21062);
xnor U21726 (N_21726,N_21089,N_21440);
nand U21727 (N_21727,N_21412,N_21588);
and U21728 (N_21728,N_21012,N_21519);
or U21729 (N_21729,N_21590,N_21469);
nand U21730 (N_21730,N_21200,N_21406);
or U21731 (N_21731,N_21229,N_21257);
nand U21732 (N_21732,N_21078,N_21014);
or U21733 (N_21733,N_21255,N_21126);
xor U21734 (N_21734,N_21369,N_21079);
or U21735 (N_21735,N_21514,N_21342);
nand U21736 (N_21736,N_21552,N_21515);
nand U21737 (N_21737,N_21560,N_21317);
xor U21738 (N_21738,N_21523,N_21143);
xor U21739 (N_21739,N_21468,N_21354);
nor U21740 (N_21740,N_21507,N_21474);
xor U21741 (N_21741,N_21410,N_21233);
and U21742 (N_21742,N_21499,N_21082);
and U21743 (N_21743,N_21216,N_21246);
nor U21744 (N_21744,N_21350,N_21021);
and U21745 (N_21745,N_21428,N_21471);
nor U21746 (N_21746,N_21032,N_21594);
nor U21747 (N_21747,N_21326,N_21593);
xnor U21748 (N_21748,N_21224,N_21168);
and U21749 (N_21749,N_21335,N_21492);
and U21750 (N_21750,N_21546,N_21532);
nor U21751 (N_21751,N_21303,N_21438);
or U21752 (N_21752,N_21102,N_21446);
nor U21753 (N_21753,N_21592,N_21313);
or U21754 (N_21754,N_21100,N_21023);
and U21755 (N_21755,N_21015,N_21165);
nor U21756 (N_21756,N_21088,N_21148);
nor U21757 (N_21757,N_21370,N_21393);
and U21758 (N_21758,N_21150,N_21517);
xor U21759 (N_21759,N_21031,N_21181);
and U21760 (N_21760,N_21298,N_21520);
and U21761 (N_21761,N_21308,N_21597);
and U21762 (N_21762,N_21409,N_21426);
and U21763 (N_21763,N_21569,N_21049);
and U21764 (N_21764,N_21232,N_21025);
and U21765 (N_21765,N_21360,N_21408);
nor U21766 (N_21766,N_21189,N_21095);
and U21767 (N_21767,N_21307,N_21453);
and U21768 (N_21768,N_21394,N_21559);
and U21769 (N_21769,N_21020,N_21160);
or U21770 (N_21770,N_21253,N_21016);
and U21771 (N_21771,N_21570,N_21356);
nor U21772 (N_21772,N_21109,N_21598);
nand U21773 (N_21773,N_21576,N_21377);
nor U21774 (N_21774,N_21521,N_21292);
xnor U21775 (N_21775,N_21477,N_21445);
nor U21776 (N_21776,N_21333,N_21234);
or U21777 (N_21777,N_21185,N_21555);
xor U21778 (N_21778,N_21267,N_21572);
xor U21779 (N_21779,N_21321,N_21266);
and U21780 (N_21780,N_21504,N_21329);
nand U21781 (N_21781,N_21508,N_21399);
nor U21782 (N_21782,N_21320,N_21373);
or U21783 (N_21783,N_21544,N_21548);
or U21784 (N_21784,N_21379,N_21040);
nand U21785 (N_21785,N_21128,N_21476);
xnor U21786 (N_21786,N_21575,N_21297);
xor U21787 (N_21787,N_21006,N_21518);
xor U21788 (N_21788,N_21201,N_21215);
nand U21789 (N_21789,N_21029,N_21220);
xor U21790 (N_21790,N_21557,N_21382);
and U21791 (N_21791,N_21053,N_21561);
or U21792 (N_21792,N_21534,N_21129);
nor U21793 (N_21793,N_21524,N_21173);
or U21794 (N_21794,N_21273,N_21591);
nor U21795 (N_21795,N_21525,N_21007);
nand U21796 (N_21796,N_21059,N_21396);
xor U21797 (N_21797,N_21203,N_21595);
nor U21798 (N_21798,N_21086,N_21416);
xnor U21799 (N_21799,N_21545,N_21429);
xor U21800 (N_21800,N_21535,N_21461);
nor U21801 (N_21801,N_21365,N_21387);
nor U21802 (N_21802,N_21459,N_21091);
nand U21803 (N_21803,N_21188,N_21511);
xnor U21804 (N_21804,N_21209,N_21328);
and U21805 (N_21805,N_21046,N_21487);
nand U21806 (N_21806,N_21312,N_21378);
and U21807 (N_21807,N_21106,N_21198);
nor U21808 (N_21808,N_21219,N_21140);
and U21809 (N_21809,N_21439,N_21156);
xor U21810 (N_21810,N_21250,N_21388);
and U21811 (N_21811,N_21034,N_21596);
and U21812 (N_21812,N_21290,N_21155);
xor U21813 (N_21813,N_21063,N_21493);
nand U21814 (N_21814,N_21235,N_21212);
or U21815 (N_21815,N_21565,N_21207);
and U21816 (N_21816,N_21516,N_21180);
nand U21817 (N_21817,N_21277,N_21425);
nand U21818 (N_21818,N_21019,N_21540);
xnor U21819 (N_21819,N_21270,N_21280);
and U21820 (N_21820,N_21099,N_21217);
xnor U21821 (N_21821,N_21264,N_21450);
nor U21822 (N_21822,N_21247,N_21187);
nor U21823 (N_21823,N_21587,N_21417);
nand U21824 (N_21824,N_21153,N_21536);
or U21825 (N_21825,N_21265,N_21167);
xor U21826 (N_21826,N_21175,N_21041);
nor U21827 (N_21827,N_21567,N_21586);
nor U21828 (N_21828,N_21385,N_21384);
nor U21829 (N_21829,N_21158,N_21304);
and U21830 (N_21830,N_21497,N_21466);
nand U21831 (N_21831,N_21085,N_21281);
nand U21832 (N_21832,N_21483,N_21056);
nor U21833 (N_21833,N_21374,N_21437);
xnor U21834 (N_21834,N_21505,N_21475);
and U21835 (N_21835,N_21451,N_21533);
nand U21836 (N_21836,N_21503,N_21008);
or U21837 (N_21837,N_21177,N_21318);
nand U21838 (N_21838,N_21383,N_21252);
nand U21839 (N_21839,N_21066,N_21263);
nand U21840 (N_21840,N_21103,N_21205);
nand U21841 (N_21841,N_21556,N_21573);
and U21842 (N_21842,N_21037,N_21322);
xnor U21843 (N_21843,N_21482,N_21067);
xor U21844 (N_21844,N_21097,N_21299);
and U21845 (N_21845,N_21113,N_21214);
xor U21846 (N_21846,N_21118,N_21344);
nand U21847 (N_21847,N_21581,N_21018);
or U21848 (N_21848,N_21538,N_21510);
and U21849 (N_21849,N_21098,N_21027);
nor U21850 (N_21850,N_21009,N_21154);
xor U21851 (N_21851,N_21191,N_21094);
and U21852 (N_21852,N_21457,N_21193);
xnor U21853 (N_21853,N_21362,N_21291);
xnor U21854 (N_21854,N_21537,N_21166);
xor U21855 (N_21855,N_21315,N_21038);
nand U21856 (N_21856,N_21311,N_21436);
and U21857 (N_21857,N_21076,N_21230);
nor U21858 (N_21858,N_21068,N_21490);
nor U21859 (N_21859,N_21282,N_21442);
or U21860 (N_21860,N_21272,N_21563);
or U21861 (N_21861,N_21397,N_21353);
nand U21862 (N_21862,N_21554,N_21339);
nand U21863 (N_21863,N_21529,N_21036);
and U21864 (N_21864,N_21568,N_21083);
xor U21865 (N_21865,N_21509,N_21035);
and U21866 (N_21866,N_21190,N_21149);
or U21867 (N_21867,N_21541,N_21052);
nor U21868 (N_21868,N_21407,N_21431);
nand U21869 (N_21869,N_21392,N_21316);
and U21870 (N_21870,N_21455,N_21389);
nand U21871 (N_21871,N_21104,N_21302);
nand U21872 (N_21872,N_21042,N_21549);
nor U21873 (N_21873,N_21054,N_21197);
and U21874 (N_21874,N_21494,N_21186);
nor U21875 (N_21875,N_21458,N_21213);
nand U21876 (N_21876,N_21327,N_21048);
xnor U21877 (N_21877,N_21141,N_21547);
nor U21878 (N_21878,N_21293,N_21571);
nand U21879 (N_21879,N_21479,N_21294);
and U21880 (N_21880,N_21169,N_21501);
xor U21881 (N_21881,N_21348,N_21488);
nand U21882 (N_21882,N_21300,N_21364);
xor U21883 (N_21883,N_21341,N_21239);
or U21884 (N_21884,N_21589,N_21413);
or U21885 (N_21885,N_21566,N_21182);
nand U21886 (N_21886,N_21051,N_21123);
nor U21887 (N_21887,N_21065,N_21107);
and U21888 (N_21888,N_21026,N_21551);
or U21889 (N_21889,N_21435,N_21484);
nand U21890 (N_21890,N_21236,N_21162);
xor U21891 (N_21891,N_21527,N_21331);
or U21892 (N_21892,N_21390,N_21125);
nand U21893 (N_21893,N_21226,N_21371);
or U21894 (N_21894,N_21305,N_21443);
and U21895 (N_21895,N_21184,N_21114);
xnor U21896 (N_21896,N_21249,N_21462);
xnor U21897 (N_21897,N_21585,N_21043);
and U21898 (N_21898,N_21022,N_21310);
and U21899 (N_21899,N_21072,N_21285);
or U21900 (N_21900,N_21449,N_21270);
xor U21901 (N_21901,N_21500,N_21507);
xor U21902 (N_21902,N_21324,N_21485);
xor U21903 (N_21903,N_21550,N_21028);
and U21904 (N_21904,N_21381,N_21101);
or U21905 (N_21905,N_21582,N_21113);
and U21906 (N_21906,N_21311,N_21526);
and U21907 (N_21907,N_21290,N_21481);
or U21908 (N_21908,N_21355,N_21497);
and U21909 (N_21909,N_21467,N_21522);
nor U21910 (N_21910,N_21012,N_21441);
nand U21911 (N_21911,N_21548,N_21344);
nand U21912 (N_21912,N_21167,N_21591);
nand U21913 (N_21913,N_21272,N_21506);
and U21914 (N_21914,N_21363,N_21596);
and U21915 (N_21915,N_21264,N_21413);
xor U21916 (N_21916,N_21452,N_21408);
xor U21917 (N_21917,N_21123,N_21112);
nand U21918 (N_21918,N_21437,N_21031);
xnor U21919 (N_21919,N_21195,N_21523);
or U21920 (N_21920,N_21386,N_21122);
xnor U21921 (N_21921,N_21051,N_21287);
and U21922 (N_21922,N_21500,N_21240);
nand U21923 (N_21923,N_21501,N_21579);
xor U21924 (N_21924,N_21366,N_21240);
nor U21925 (N_21925,N_21467,N_21208);
and U21926 (N_21926,N_21576,N_21391);
and U21927 (N_21927,N_21482,N_21226);
or U21928 (N_21928,N_21533,N_21225);
xnor U21929 (N_21929,N_21301,N_21274);
nor U21930 (N_21930,N_21413,N_21497);
and U21931 (N_21931,N_21572,N_21336);
nor U21932 (N_21932,N_21318,N_21126);
and U21933 (N_21933,N_21555,N_21523);
and U21934 (N_21934,N_21189,N_21526);
or U21935 (N_21935,N_21391,N_21312);
nand U21936 (N_21936,N_21389,N_21126);
nor U21937 (N_21937,N_21389,N_21394);
and U21938 (N_21938,N_21545,N_21506);
nor U21939 (N_21939,N_21427,N_21233);
nor U21940 (N_21940,N_21007,N_21485);
nor U21941 (N_21941,N_21461,N_21082);
or U21942 (N_21942,N_21227,N_21203);
xnor U21943 (N_21943,N_21355,N_21230);
and U21944 (N_21944,N_21338,N_21450);
or U21945 (N_21945,N_21206,N_21518);
nor U21946 (N_21946,N_21208,N_21046);
or U21947 (N_21947,N_21559,N_21201);
nand U21948 (N_21948,N_21119,N_21436);
and U21949 (N_21949,N_21016,N_21279);
nand U21950 (N_21950,N_21534,N_21262);
nand U21951 (N_21951,N_21174,N_21316);
and U21952 (N_21952,N_21424,N_21225);
and U21953 (N_21953,N_21527,N_21519);
nand U21954 (N_21954,N_21512,N_21505);
nand U21955 (N_21955,N_21386,N_21280);
xnor U21956 (N_21956,N_21144,N_21201);
xor U21957 (N_21957,N_21241,N_21183);
or U21958 (N_21958,N_21169,N_21476);
or U21959 (N_21959,N_21539,N_21487);
and U21960 (N_21960,N_21075,N_21077);
xnor U21961 (N_21961,N_21265,N_21204);
nand U21962 (N_21962,N_21106,N_21350);
nand U21963 (N_21963,N_21293,N_21551);
or U21964 (N_21964,N_21091,N_21592);
nand U21965 (N_21965,N_21418,N_21474);
xnor U21966 (N_21966,N_21020,N_21350);
nor U21967 (N_21967,N_21195,N_21191);
or U21968 (N_21968,N_21446,N_21250);
nor U21969 (N_21969,N_21382,N_21357);
xnor U21970 (N_21970,N_21373,N_21236);
nand U21971 (N_21971,N_21130,N_21196);
or U21972 (N_21972,N_21027,N_21147);
xor U21973 (N_21973,N_21457,N_21476);
or U21974 (N_21974,N_21235,N_21239);
and U21975 (N_21975,N_21576,N_21075);
nand U21976 (N_21976,N_21022,N_21109);
nor U21977 (N_21977,N_21418,N_21280);
nor U21978 (N_21978,N_21463,N_21582);
nand U21979 (N_21979,N_21043,N_21093);
nand U21980 (N_21980,N_21476,N_21244);
xnor U21981 (N_21981,N_21338,N_21342);
or U21982 (N_21982,N_21005,N_21270);
nor U21983 (N_21983,N_21568,N_21054);
nand U21984 (N_21984,N_21117,N_21365);
or U21985 (N_21985,N_21221,N_21098);
nand U21986 (N_21986,N_21058,N_21032);
nor U21987 (N_21987,N_21485,N_21398);
xnor U21988 (N_21988,N_21329,N_21417);
xor U21989 (N_21989,N_21522,N_21362);
or U21990 (N_21990,N_21577,N_21006);
nor U21991 (N_21991,N_21462,N_21573);
and U21992 (N_21992,N_21087,N_21070);
nand U21993 (N_21993,N_21243,N_21438);
xor U21994 (N_21994,N_21303,N_21183);
nand U21995 (N_21995,N_21075,N_21151);
xor U21996 (N_21996,N_21377,N_21244);
and U21997 (N_21997,N_21471,N_21375);
nand U21998 (N_21998,N_21352,N_21335);
or U21999 (N_21999,N_21086,N_21453);
and U22000 (N_22000,N_21414,N_21169);
xnor U22001 (N_22001,N_21286,N_21221);
and U22002 (N_22002,N_21479,N_21400);
and U22003 (N_22003,N_21210,N_21530);
or U22004 (N_22004,N_21587,N_21533);
nor U22005 (N_22005,N_21378,N_21023);
nand U22006 (N_22006,N_21208,N_21318);
and U22007 (N_22007,N_21334,N_21373);
or U22008 (N_22008,N_21203,N_21324);
xnor U22009 (N_22009,N_21402,N_21482);
nand U22010 (N_22010,N_21240,N_21270);
nand U22011 (N_22011,N_21425,N_21552);
and U22012 (N_22012,N_21411,N_21518);
nand U22013 (N_22013,N_21172,N_21363);
and U22014 (N_22014,N_21353,N_21437);
or U22015 (N_22015,N_21536,N_21463);
nand U22016 (N_22016,N_21036,N_21413);
nand U22017 (N_22017,N_21441,N_21234);
nand U22018 (N_22018,N_21297,N_21201);
nor U22019 (N_22019,N_21514,N_21433);
nand U22020 (N_22020,N_21440,N_21236);
and U22021 (N_22021,N_21116,N_21573);
or U22022 (N_22022,N_21103,N_21381);
nand U22023 (N_22023,N_21083,N_21048);
nor U22024 (N_22024,N_21444,N_21548);
nor U22025 (N_22025,N_21575,N_21558);
nand U22026 (N_22026,N_21024,N_21357);
nand U22027 (N_22027,N_21486,N_21404);
xor U22028 (N_22028,N_21112,N_21495);
and U22029 (N_22029,N_21110,N_21564);
nand U22030 (N_22030,N_21177,N_21065);
xnor U22031 (N_22031,N_21097,N_21044);
nand U22032 (N_22032,N_21209,N_21308);
nor U22033 (N_22033,N_21189,N_21064);
and U22034 (N_22034,N_21426,N_21140);
or U22035 (N_22035,N_21104,N_21292);
nor U22036 (N_22036,N_21494,N_21447);
xor U22037 (N_22037,N_21205,N_21399);
nor U22038 (N_22038,N_21310,N_21323);
xnor U22039 (N_22039,N_21438,N_21100);
nor U22040 (N_22040,N_21585,N_21219);
nor U22041 (N_22041,N_21596,N_21315);
or U22042 (N_22042,N_21293,N_21369);
and U22043 (N_22043,N_21317,N_21407);
xnor U22044 (N_22044,N_21239,N_21522);
and U22045 (N_22045,N_21387,N_21059);
nor U22046 (N_22046,N_21382,N_21521);
xnor U22047 (N_22047,N_21084,N_21072);
or U22048 (N_22048,N_21452,N_21068);
nor U22049 (N_22049,N_21552,N_21068);
or U22050 (N_22050,N_21186,N_21060);
and U22051 (N_22051,N_21131,N_21474);
or U22052 (N_22052,N_21156,N_21527);
nor U22053 (N_22053,N_21479,N_21061);
nand U22054 (N_22054,N_21400,N_21513);
nor U22055 (N_22055,N_21142,N_21000);
xor U22056 (N_22056,N_21378,N_21221);
xnor U22057 (N_22057,N_21373,N_21155);
or U22058 (N_22058,N_21516,N_21595);
and U22059 (N_22059,N_21279,N_21225);
nand U22060 (N_22060,N_21401,N_21229);
or U22061 (N_22061,N_21131,N_21458);
nor U22062 (N_22062,N_21357,N_21291);
and U22063 (N_22063,N_21401,N_21147);
xnor U22064 (N_22064,N_21345,N_21024);
and U22065 (N_22065,N_21166,N_21497);
nand U22066 (N_22066,N_21136,N_21405);
nand U22067 (N_22067,N_21064,N_21330);
or U22068 (N_22068,N_21349,N_21260);
xnor U22069 (N_22069,N_21026,N_21108);
and U22070 (N_22070,N_21573,N_21596);
xnor U22071 (N_22071,N_21030,N_21107);
and U22072 (N_22072,N_21459,N_21151);
or U22073 (N_22073,N_21280,N_21260);
nor U22074 (N_22074,N_21320,N_21439);
xor U22075 (N_22075,N_21058,N_21201);
or U22076 (N_22076,N_21372,N_21310);
nand U22077 (N_22077,N_21517,N_21146);
nor U22078 (N_22078,N_21030,N_21234);
xnor U22079 (N_22079,N_21018,N_21119);
or U22080 (N_22080,N_21098,N_21485);
xnor U22081 (N_22081,N_21493,N_21234);
nand U22082 (N_22082,N_21564,N_21533);
nor U22083 (N_22083,N_21273,N_21425);
and U22084 (N_22084,N_21534,N_21139);
nand U22085 (N_22085,N_21441,N_21418);
xnor U22086 (N_22086,N_21102,N_21136);
nor U22087 (N_22087,N_21350,N_21130);
and U22088 (N_22088,N_21506,N_21466);
xnor U22089 (N_22089,N_21210,N_21394);
nand U22090 (N_22090,N_21005,N_21034);
nand U22091 (N_22091,N_21544,N_21291);
nor U22092 (N_22092,N_21004,N_21123);
and U22093 (N_22093,N_21581,N_21311);
or U22094 (N_22094,N_21392,N_21035);
and U22095 (N_22095,N_21593,N_21529);
nor U22096 (N_22096,N_21196,N_21166);
nor U22097 (N_22097,N_21037,N_21519);
and U22098 (N_22098,N_21351,N_21509);
or U22099 (N_22099,N_21380,N_21029);
nor U22100 (N_22100,N_21352,N_21242);
and U22101 (N_22101,N_21393,N_21055);
nor U22102 (N_22102,N_21500,N_21510);
and U22103 (N_22103,N_21331,N_21552);
and U22104 (N_22104,N_21572,N_21399);
nor U22105 (N_22105,N_21543,N_21169);
nand U22106 (N_22106,N_21390,N_21459);
nand U22107 (N_22107,N_21362,N_21172);
and U22108 (N_22108,N_21113,N_21466);
or U22109 (N_22109,N_21079,N_21487);
xnor U22110 (N_22110,N_21468,N_21347);
nand U22111 (N_22111,N_21227,N_21164);
nor U22112 (N_22112,N_21301,N_21226);
and U22113 (N_22113,N_21491,N_21022);
and U22114 (N_22114,N_21171,N_21482);
nand U22115 (N_22115,N_21333,N_21133);
or U22116 (N_22116,N_21287,N_21097);
nor U22117 (N_22117,N_21200,N_21414);
or U22118 (N_22118,N_21239,N_21216);
nand U22119 (N_22119,N_21097,N_21093);
and U22120 (N_22120,N_21348,N_21059);
or U22121 (N_22121,N_21492,N_21100);
nor U22122 (N_22122,N_21028,N_21105);
or U22123 (N_22123,N_21271,N_21260);
nor U22124 (N_22124,N_21201,N_21158);
nor U22125 (N_22125,N_21400,N_21183);
nand U22126 (N_22126,N_21254,N_21226);
and U22127 (N_22127,N_21059,N_21125);
or U22128 (N_22128,N_21440,N_21002);
xor U22129 (N_22129,N_21328,N_21262);
xnor U22130 (N_22130,N_21131,N_21496);
xor U22131 (N_22131,N_21115,N_21247);
or U22132 (N_22132,N_21227,N_21142);
or U22133 (N_22133,N_21503,N_21326);
xor U22134 (N_22134,N_21573,N_21212);
or U22135 (N_22135,N_21535,N_21115);
nand U22136 (N_22136,N_21084,N_21157);
and U22137 (N_22137,N_21301,N_21568);
xor U22138 (N_22138,N_21574,N_21020);
or U22139 (N_22139,N_21565,N_21582);
xnor U22140 (N_22140,N_21388,N_21288);
nand U22141 (N_22141,N_21284,N_21329);
nor U22142 (N_22142,N_21469,N_21059);
nand U22143 (N_22143,N_21146,N_21487);
and U22144 (N_22144,N_21123,N_21195);
xnor U22145 (N_22145,N_21203,N_21207);
xnor U22146 (N_22146,N_21570,N_21233);
or U22147 (N_22147,N_21305,N_21139);
nor U22148 (N_22148,N_21469,N_21047);
and U22149 (N_22149,N_21446,N_21499);
nor U22150 (N_22150,N_21279,N_21307);
or U22151 (N_22151,N_21312,N_21110);
or U22152 (N_22152,N_21315,N_21357);
xor U22153 (N_22153,N_21269,N_21565);
or U22154 (N_22154,N_21364,N_21387);
and U22155 (N_22155,N_21565,N_21208);
nor U22156 (N_22156,N_21228,N_21160);
or U22157 (N_22157,N_21490,N_21517);
nand U22158 (N_22158,N_21520,N_21412);
or U22159 (N_22159,N_21138,N_21527);
nand U22160 (N_22160,N_21426,N_21597);
nand U22161 (N_22161,N_21080,N_21040);
xor U22162 (N_22162,N_21529,N_21300);
nand U22163 (N_22163,N_21089,N_21108);
nand U22164 (N_22164,N_21358,N_21552);
or U22165 (N_22165,N_21291,N_21200);
nor U22166 (N_22166,N_21451,N_21226);
or U22167 (N_22167,N_21117,N_21124);
nor U22168 (N_22168,N_21246,N_21482);
nor U22169 (N_22169,N_21223,N_21120);
and U22170 (N_22170,N_21410,N_21148);
nand U22171 (N_22171,N_21291,N_21332);
nand U22172 (N_22172,N_21012,N_21475);
and U22173 (N_22173,N_21360,N_21464);
or U22174 (N_22174,N_21021,N_21416);
and U22175 (N_22175,N_21277,N_21048);
nand U22176 (N_22176,N_21595,N_21381);
nor U22177 (N_22177,N_21131,N_21276);
and U22178 (N_22178,N_21109,N_21112);
nand U22179 (N_22179,N_21380,N_21534);
nor U22180 (N_22180,N_21314,N_21377);
xor U22181 (N_22181,N_21230,N_21296);
and U22182 (N_22182,N_21311,N_21367);
nor U22183 (N_22183,N_21103,N_21467);
nand U22184 (N_22184,N_21540,N_21330);
or U22185 (N_22185,N_21228,N_21420);
xnor U22186 (N_22186,N_21423,N_21209);
or U22187 (N_22187,N_21446,N_21467);
and U22188 (N_22188,N_21124,N_21438);
xor U22189 (N_22189,N_21163,N_21373);
nor U22190 (N_22190,N_21146,N_21032);
or U22191 (N_22191,N_21169,N_21321);
xor U22192 (N_22192,N_21234,N_21201);
xnor U22193 (N_22193,N_21195,N_21043);
and U22194 (N_22194,N_21411,N_21364);
xnor U22195 (N_22195,N_21410,N_21416);
xnor U22196 (N_22196,N_21116,N_21079);
and U22197 (N_22197,N_21592,N_21147);
xor U22198 (N_22198,N_21445,N_21362);
or U22199 (N_22199,N_21174,N_21436);
nor U22200 (N_22200,N_21727,N_22140);
xnor U22201 (N_22201,N_22026,N_22019);
xor U22202 (N_22202,N_21692,N_22094);
and U22203 (N_22203,N_21702,N_22043);
and U22204 (N_22204,N_22083,N_21623);
xor U22205 (N_22205,N_21807,N_21696);
xnor U22206 (N_22206,N_21875,N_22169);
xor U22207 (N_22207,N_21643,N_21866);
and U22208 (N_22208,N_21862,N_21611);
or U22209 (N_22209,N_21870,N_22000);
nand U22210 (N_22210,N_22049,N_22034);
and U22211 (N_22211,N_21867,N_22001);
and U22212 (N_22212,N_21794,N_21934);
nand U22213 (N_22213,N_21806,N_21826);
xor U22214 (N_22214,N_21832,N_21812);
or U22215 (N_22215,N_21805,N_22171);
nand U22216 (N_22216,N_21881,N_22078);
nor U22217 (N_22217,N_22192,N_21697);
or U22218 (N_22218,N_21726,N_22128);
xnor U22219 (N_22219,N_22161,N_21746);
or U22220 (N_22220,N_22136,N_21993);
and U22221 (N_22221,N_22058,N_21690);
nor U22222 (N_22222,N_21943,N_22070);
nand U22223 (N_22223,N_21885,N_22084);
xnor U22224 (N_22224,N_21648,N_21985);
nor U22225 (N_22225,N_21714,N_21616);
nor U22226 (N_22226,N_21653,N_22120);
or U22227 (N_22227,N_21990,N_22007);
xnor U22228 (N_22228,N_21937,N_21755);
xnor U22229 (N_22229,N_21986,N_21811);
or U22230 (N_22230,N_21845,N_22130);
nor U22231 (N_22231,N_22087,N_21822);
or U22232 (N_22232,N_21821,N_21860);
and U22233 (N_22233,N_21841,N_21961);
or U22234 (N_22234,N_21838,N_21799);
nand U22235 (N_22235,N_21905,N_21914);
nand U22236 (N_22236,N_21863,N_22177);
xor U22237 (N_22237,N_21602,N_22009);
or U22238 (N_22238,N_21886,N_21922);
xor U22239 (N_22239,N_21667,N_21903);
nor U22240 (N_22240,N_21979,N_21780);
xor U22241 (N_22241,N_22173,N_22011);
or U22242 (N_22242,N_21820,N_21716);
nand U22243 (N_22243,N_21703,N_21786);
nand U22244 (N_22244,N_22164,N_21778);
nor U22245 (N_22245,N_21808,N_21837);
and U22246 (N_22246,N_22198,N_21906);
nor U22247 (N_22247,N_22146,N_22153);
or U22248 (N_22248,N_21916,N_21765);
or U22249 (N_22249,N_22071,N_22048);
or U22250 (N_22250,N_21917,N_21936);
and U22251 (N_22251,N_21710,N_21946);
and U22252 (N_22252,N_21883,N_21952);
nand U22253 (N_22253,N_21694,N_21728);
and U22254 (N_22254,N_22193,N_21941);
or U22255 (N_22255,N_21843,N_22158);
nor U22256 (N_22256,N_22039,N_21959);
nand U22257 (N_22257,N_21745,N_21717);
and U22258 (N_22258,N_21898,N_22135);
xnor U22259 (N_22259,N_21685,N_21974);
or U22260 (N_22260,N_21782,N_22187);
nor U22261 (N_22261,N_21802,N_22138);
or U22262 (N_22262,N_21718,N_21868);
nor U22263 (N_22263,N_21774,N_21908);
nor U22264 (N_22264,N_21713,N_22156);
nand U22265 (N_22265,N_21854,N_21955);
nand U22266 (N_22266,N_21664,N_22099);
or U22267 (N_22267,N_21999,N_21938);
nand U22268 (N_22268,N_21646,N_22097);
or U22269 (N_22269,N_22038,N_22176);
nand U22270 (N_22270,N_21689,N_21677);
or U22271 (N_22271,N_21632,N_22086);
nor U22272 (N_22272,N_22137,N_22121);
xnor U22273 (N_22273,N_22040,N_21925);
or U22274 (N_22274,N_21833,N_21607);
nand U22275 (N_22275,N_21736,N_21700);
xor U22276 (N_22276,N_21801,N_21666);
nor U22277 (N_22277,N_22190,N_21850);
or U22278 (N_22278,N_21784,N_22015);
xnor U22279 (N_22279,N_21661,N_21682);
nand U22280 (N_22280,N_21939,N_21958);
and U22281 (N_22281,N_21608,N_22144);
xnor U22282 (N_22282,N_21753,N_21707);
nand U22283 (N_22283,N_22091,N_21779);
and U22284 (N_22284,N_21940,N_21688);
and U22285 (N_22285,N_21858,N_22059);
xor U22286 (N_22286,N_22032,N_21600);
or U22287 (N_22287,N_22013,N_21751);
xor U22288 (N_22288,N_22103,N_21754);
nand U22289 (N_22289,N_22055,N_21988);
nand U22290 (N_22290,N_21948,N_21629);
or U22291 (N_22291,N_22141,N_21855);
or U22292 (N_22292,N_21884,N_21676);
or U22293 (N_22293,N_22003,N_21894);
nor U22294 (N_22294,N_22054,N_21798);
xnor U22295 (N_22295,N_21642,N_22018);
nand U22296 (N_22296,N_21732,N_21861);
or U22297 (N_22297,N_22062,N_22079);
xnor U22298 (N_22298,N_21951,N_21633);
nand U22299 (N_22299,N_21725,N_21947);
xnor U22300 (N_22300,N_21790,N_21731);
xor U22301 (N_22301,N_21724,N_21735);
xnor U22302 (N_22302,N_21647,N_21781);
nor U22303 (N_22303,N_21721,N_21966);
xnor U22304 (N_22304,N_21889,N_21859);
and U22305 (N_22305,N_21998,N_22104);
nor U22306 (N_22306,N_21771,N_21686);
xor U22307 (N_22307,N_21815,N_21758);
or U22308 (N_22308,N_21891,N_21788);
xnor U22309 (N_22309,N_21827,N_21665);
nand U22310 (N_22310,N_22021,N_22122);
nand U22311 (N_22311,N_21994,N_21787);
xnor U22312 (N_22312,N_21762,N_21683);
or U22313 (N_22313,N_21670,N_22178);
nand U22314 (N_22314,N_21738,N_22030);
and U22315 (N_22315,N_22124,N_21928);
xnor U22316 (N_22316,N_21704,N_21913);
or U22317 (N_22317,N_22063,N_21847);
nand U22318 (N_22318,N_21626,N_21612);
xor U22319 (N_22319,N_21622,N_21747);
xor U22320 (N_22320,N_21831,N_21896);
nor U22321 (N_22321,N_21679,N_22166);
and U22322 (N_22322,N_21942,N_22085);
and U22323 (N_22323,N_22133,N_21969);
or U22324 (N_22324,N_21671,N_21856);
nand U22325 (N_22325,N_22194,N_21605);
or U22326 (N_22326,N_21888,N_21953);
xor U22327 (N_22327,N_22139,N_22186);
xnor U22328 (N_22328,N_22060,N_21950);
nor U22329 (N_22329,N_22196,N_22113);
or U22330 (N_22330,N_22061,N_22115);
or U22331 (N_22331,N_21711,N_21921);
xnor U22332 (N_22332,N_21759,N_21730);
and U22333 (N_22333,N_21907,N_21800);
or U22334 (N_22334,N_22175,N_21723);
and U22335 (N_22335,N_21920,N_22167);
and U22336 (N_22336,N_21699,N_21835);
xor U22337 (N_22337,N_22075,N_21639);
nand U22338 (N_22338,N_22143,N_21624);
nand U22339 (N_22339,N_21931,N_22065);
xor U22340 (N_22340,N_22081,N_21764);
and U22341 (N_22341,N_21628,N_21972);
nand U22342 (N_22342,N_21744,N_21637);
and U22343 (N_22343,N_21901,N_22107);
nor U22344 (N_22344,N_22082,N_21963);
xor U22345 (N_22345,N_21695,N_21772);
and U22346 (N_22346,N_21962,N_22183);
nand U22347 (N_22347,N_21880,N_21627);
nand U22348 (N_22348,N_21823,N_21836);
xnor U22349 (N_22349,N_21978,N_21680);
and U22350 (N_22350,N_21967,N_21892);
and U22351 (N_22351,N_21949,N_21797);
nor U22352 (N_22352,N_21621,N_21849);
nand U22353 (N_22353,N_21640,N_21672);
and U22354 (N_22354,N_21842,N_21681);
and U22355 (N_22355,N_22014,N_21877);
nor U22356 (N_22356,N_22093,N_22008);
xor U22357 (N_22357,N_21663,N_22147);
nand U22358 (N_22358,N_21975,N_21748);
nor U22359 (N_22359,N_21630,N_21659);
and U22360 (N_22360,N_21846,N_21853);
and U22361 (N_22361,N_21882,N_22096);
nand U22362 (N_22362,N_21770,N_22126);
xnor U22363 (N_22363,N_21674,N_21840);
xnor U22364 (N_22364,N_21918,N_22041);
xnor U22365 (N_22365,N_21625,N_22046);
nand U22366 (N_22366,N_22073,N_22116);
nand U22367 (N_22367,N_22064,N_21954);
and U22368 (N_22368,N_21698,N_21618);
xnor U22369 (N_22369,N_22145,N_22101);
xor U22370 (N_22370,N_22072,N_21701);
nand U22371 (N_22371,N_22052,N_21777);
xnor U22372 (N_22372,N_21852,N_22182);
nand U22373 (N_22373,N_21749,N_22056);
xor U22374 (N_22374,N_21829,N_21851);
xnor U22375 (N_22375,N_21752,N_22191);
xor U22376 (N_22376,N_22108,N_21857);
nor U22377 (N_22377,N_21926,N_21601);
or U22378 (N_22378,N_21933,N_22037);
xnor U22379 (N_22379,N_21684,N_22023);
or U22380 (N_22380,N_22155,N_21957);
xnor U22381 (N_22381,N_22105,N_22163);
or U22382 (N_22382,N_22119,N_21654);
nor U22383 (N_22383,N_22112,N_22195);
nor U22384 (N_22384,N_21935,N_21923);
xnor U22385 (N_22385,N_21878,N_22131);
and U22386 (N_22386,N_21817,N_21776);
or U22387 (N_22387,N_21742,N_21615);
nand U22388 (N_22388,N_21660,N_21810);
nand U22389 (N_22389,N_21613,N_22031);
and U22390 (N_22390,N_21791,N_22162);
nor U22391 (N_22391,N_22022,N_22016);
xor U22392 (N_22392,N_21641,N_22024);
and U22393 (N_22393,N_22102,N_22074);
nand U22394 (N_22394,N_22125,N_22159);
and U22395 (N_22395,N_21973,N_21828);
and U22396 (N_22396,N_22127,N_22017);
nor U22397 (N_22397,N_21793,N_22095);
and U22398 (N_22398,N_21971,N_21981);
xor U22399 (N_22399,N_21919,N_22006);
xnor U22400 (N_22400,N_21818,N_21864);
or U22401 (N_22401,N_22152,N_21768);
or U22402 (N_22402,N_21869,N_21789);
nor U22403 (N_22403,N_22118,N_21708);
and U22404 (N_22404,N_21729,N_21669);
and U22405 (N_22405,N_21650,N_21893);
or U22406 (N_22406,N_21634,N_21709);
xnor U22407 (N_22407,N_21652,N_21995);
and U22408 (N_22408,N_22106,N_22134);
and U22409 (N_22409,N_21814,N_22168);
nand U22410 (N_22410,N_22027,N_21945);
or U22411 (N_22411,N_21756,N_22165);
nor U22412 (N_22412,N_22033,N_21636);
nor U22413 (N_22413,N_21638,N_22184);
nor U22414 (N_22414,N_21606,N_21783);
or U22415 (N_22415,N_21987,N_21750);
or U22416 (N_22416,N_22154,N_21733);
and U22417 (N_22417,N_22090,N_21819);
xnor U22418 (N_22418,N_21792,N_21911);
and U22419 (N_22419,N_22174,N_22111);
xnor U22420 (N_22420,N_21960,N_22098);
xnor U22421 (N_22421,N_22029,N_21769);
xor U22422 (N_22422,N_21839,N_21909);
or U22423 (N_22423,N_22179,N_21757);
nor U22424 (N_22424,N_22028,N_22088);
or U22425 (N_22425,N_22148,N_21649);
nor U22426 (N_22426,N_21968,N_22010);
nand U22427 (N_22427,N_21675,N_21720);
and U22428 (N_22428,N_21743,N_22157);
nor U22429 (N_22429,N_21897,N_22012);
xor U22430 (N_22430,N_21982,N_21900);
and U22431 (N_22431,N_21610,N_21773);
xnor U22432 (N_22432,N_21740,N_22002);
or U22433 (N_22433,N_21706,N_21910);
and U22434 (N_22434,N_21767,N_21984);
nor U22435 (N_22435,N_21609,N_21887);
and U22436 (N_22436,N_22092,N_21992);
nor U22437 (N_22437,N_22180,N_22110);
nand U22438 (N_22438,N_21956,N_21809);
or U22439 (N_22439,N_21977,N_21983);
xnor U22440 (N_22440,N_21631,N_21619);
nand U22441 (N_22441,N_21796,N_22077);
xnor U22442 (N_22442,N_21865,N_21929);
xor U22443 (N_22443,N_21876,N_21614);
or U22444 (N_22444,N_21693,N_21927);
nor U22445 (N_22445,N_22150,N_22160);
and U22446 (N_22446,N_21924,N_21873);
and U22447 (N_22447,N_21687,N_21691);
nor U22448 (N_22448,N_22035,N_22004);
nor U22449 (N_22449,N_21719,N_21871);
and U22450 (N_22450,N_22080,N_21915);
and U22451 (N_22451,N_21813,N_22044);
or U22452 (N_22452,N_22123,N_21932);
nor U22453 (N_22453,N_22047,N_21673);
xor U22454 (N_22454,N_21997,N_21804);
xor U22455 (N_22455,N_21964,N_22188);
xor U22456 (N_22456,N_22067,N_21761);
nand U22457 (N_22457,N_22053,N_22005);
xor U22458 (N_22458,N_21658,N_21879);
nor U22459 (N_22459,N_21816,N_21890);
nand U22460 (N_22460,N_22066,N_21976);
nand U22461 (N_22461,N_21734,N_21912);
nand U22462 (N_22462,N_22151,N_21848);
nand U22463 (N_22463,N_22189,N_21644);
nand U22464 (N_22464,N_22170,N_21899);
xnor U22465 (N_22465,N_21980,N_21844);
or U22466 (N_22466,N_22068,N_22114);
nor U22467 (N_22467,N_21996,N_22149);
nor U22468 (N_22468,N_22197,N_22109);
nor U22469 (N_22469,N_22036,N_21705);
or U22470 (N_22470,N_21712,N_21678);
or U22471 (N_22471,N_21657,N_21904);
and U22472 (N_22472,N_22051,N_21737);
xor U22473 (N_22473,N_22199,N_22076);
xor U22474 (N_22474,N_21651,N_21874);
xnor U22475 (N_22475,N_22045,N_22057);
xnor U22476 (N_22476,N_22025,N_21825);
nand U22477 (N_22477,N_21775,N_21872);
or U22478 (N_22478,N_22172,N_21785);
nand U22479 (N_22479,N_22050,N_21635);
and U22480 (N_22480,N_22117,N_21766);
or U22481 (N_22481,N_22185,N_21655);
and U22482 (N_22482,N_21763,N_21989);
nand U22483 (N_22483,N_21944,N_21965);
or U22484 (N_22484,N_21715,N_21760);
xor U22485 (N_22485,N_22142,N_22129);
nand U22486 (N_22486,N_22181,N_21830);
nor U22487 (N_22487,N_21741,N_21722);
or U22488 (N_22488,N_22132,N_21895);
xnor U22489 (N_22489,N_22089,N_21620);
or U22490 (N_22490,N_21603,N_21604);
nand U22491 (N_22491,N_21902,N_22042);
xor U22492 (N_22492,N_21739,N_21834);
nor U22493 (N_22493,N_21991,N_22020);
or U22494 (N_22494,N_21668,N_22100);
or U22495 (N_22495,N_21795,N_22069);
or U22496 (N_22496,N_21662,N_21930);
nand U22497 (N_22497,N_21617,N_21970);
and U22498 (N_22498,N_21803,N_21824);
and U22499 (N_22499,N_21656,N_21645);
nand U22500 (N_22500,N_21775,N_21918);
nor U22501 (N_22501,N_21955,N_22129);
xor U22502 (N_22502,N_22050,N_22090);
xnor U22503 (N_22503,N_21825,N_21652);
nand U22504 (N_22504,N_21898,N_21700);
nand U22505 (N_22505,N_22188,N_21921);
or U22506 (N_22506,N_21685,N_22184);
nor U22507 (N_22507,N_21950,N_22199);
xnor U22508 (N_22508,N_22136,N_21888);
and U22509 (N_22509,N_21772,N_22046);
nand U22510 (N_22510,N_22082,N_22059);
nor U22511 (N_22511,N_21794,N_22083);
nand U22512 (N_22512,N_22166,N_21698);
and U22513 (N_22513,N_22010,N_21622);
or U22514 (N_22514,N_21968,N_22187);
and U22515 (N_22515,N_21905,N_22139);
nand U22516 (N_22516,N_21855,N_21947);
or U22517 (N_22517,N_21851,N_21665);
or U22518 (N_22518,N_21824,N_21652);
nor U22519 (N_22519,N_21925,N_21860);
and U22520 (N_22520,N_22043,N_22012);
nor U22521 (N_22521,N_22056,N_22027);
xnor U22522 (N_22522,N_21743,N_21896);
and U22523 (N_22523,N_21943,N_22097);
and U22524 (N_22524,N_21611,N_22137);
or U22525 (N_22525,N_21932,N_22152);
nor U22526 (N_22526,N_21737,N_21728);
xnor U22527 (N_22527,N_21796,N_21623);
xor U22528 (N_22528,N_21753,N_21627);
xor U22529 (N_22529,N_22090,N_22045);
nor U22530 (N_22530,N_21663,N_22065);
and U22531 (N_22531,N_21923,N_22195);
or U22532 (N_22532,N_21628,N_21694);
nor U22533 (N_22533,N_21648,N_22145);
or U22534 (N_22534,N_22108,N_22085);
and U22535 (N_22535,N_21983,N_21804);
nor U22536 (N_22536,N_21677,N_21814);
or U22537 (N_22537,N_22137,N_21921);
xor U22538 (N_22538,N_21848,N_21611);
nor U22539 (N_22539,N_21841,N_22060);
nor U22540 (N_22540,N_21739,N_22006);
and U22541 (N_22541,N_21886,N_21825);
and U22542 (N_22542,N_21695,N_21641);
and U22543 (N_22543,N_21765,N_21755);
or U22544 (N_22544,N_21717,N_21867);
nand U22545 (N_22545,N_21895,N_21998);
xor U22546 (N_22546,N_21934,N_21780);
and U22547 (N_22547,N_21772,N_21933);
or U22548 (N_22548,N_22112,N_21947);
and U22549 (N_22549,N_21952,N_21827);
and U22550 (N_22550,N_21700,N_21969);
nand U22551 (N_22551,N_21829,N_21736);
and U22552 (N_22552,N_21717,N_21776);
or U22553 (N_22553,N_22119,N_22110);
xnor U22554 (N_22554,N_21824,N_21783);
xor U22555 (N_22555,N_21759,N_21710);
or U22556 (N_22556,N_22005,N_22130);
nor U22557 (N_22557,N_22049,N_21913);
nand U22558 (N_22558,N_21823,N_22104);
and U22559 (N_22559,N_21831,N_21936);
or U22560 (N_22560,N_21636,N_21754);
or U22561 (N_22561,N_21681,N_22018);
xor U22562 (N_22562,N_21768,N_21795);
nand U22563 (N_22563,N_22086,N_21707);
xor U22564 (N_22564,N_22164,N_21655);
nor U22565 (N_22565,N_21823,N_22018);
and U22566 (N_22566,N_21821,N_22120);
nor U22567 (N_22567,N_22164,N_21606);
or U22568 (N_22568,N_22084,N_21699);
and U22569 (N_22569,N_21900,N_22023);
and U22570 (N_22570,N_21866,N_21885);
xor U22571 (N_22571,N_21927,N_21943);
and U22572 (N_22572,N_22015,N_21891);
and U22573 (N_22573,N_22010,N_21954);
and U22574 (N_22574,N_21722,N_21664);
xnor U22575 (N_22575,N_21736,N_21972);
nor U22576 (N_22576,N_21962,N_22158);
nand U22577 (N_22577,N_21891,N_21835);
and U22578 (N_22578,N_21889,N_21609);
xnor U22579 (N_22579,N_21959,N_21792);
and U22580 (N_22580,N_21760,N_21786);
nand U22581 (N_22581,N_21821,N_22112);
nand U22582 (N_22582,N_21893,N_22122);
nor U22583 (N_22583,N_21699,N_21760);
nand U22584 (N_22584,N_22045,N_21796);
and U22585 (N_22585,N_21889,N_21659);
and U22586 (N_22586,N_22186,N_21605);
nor U22587 (N_22587,N_22088,N_21988);
and U22588 (N_22588,N_21901,N_22027);
nor U22589 (N_22589,N_21985,N_21888);
xor U22590 (N_22590,N_22055,N_21689);
xnor U22591 (N_22591,N_21858,N_21652);
nand U22592 (N_22592,N_21755,N_21996);
nor U22593 (N_22593,N_21785,N_21908);
or U22594 (N_22594,N_22199,N_21864);
xor U22595 (N_22595,N_22005,N_22075);
nor U22596 (N_22596,N_21818,N_21607);
nor U22597 (N_22597,N_22029,N_21725);
xnor U22598 (N_22598,N_21781,N_21905);
or U22599 (N_22599,N_21903,N_22098);
nand U22600 (N_22600,N_21876,N_22196);
and U22601 (N_22601,N_22040,N_22156);
nor U22602 (N_22602,N_21779,N_22108);
nand U22603 (N_22603,N_21999,N_21830);
nand U22604 (N_22604,N_22004,N_22142);
and U22605 (N_22605,N_21987,N_21716);
xnor U22606 (N_22606,N_21768,N_21862);
xnor U22607 (N_22607,N_21910,N_21618);
and U22608 (N_22608,N_21987,N_21688);
and U22609 (N_22609,N_21683,N_22149);
nor U22610 (N_22610,N_22034,N_21699);
and U22611 (N_22611,N_22157,N_21970);
and U22612 (N_22612,N_22127,N_21870);
nand U22613 (N_22613,N_22040,N_22012);
or U22614 (N_22614,N_21663,N_21786);
or U22615 (N_22615,N_21900,N_21799);
xnor U22616 (N_22616,N_21853,N_21903);
xnor U22617 (N_22617,N_21866,N_21610);
xor U22618 (N_22618,N_22158,N_21981);
nor U22619 (N_22619,N_22129,N_21978);
or U22620 (N_22620,N_21606,N_21691);
or U22621 (N_22621,N_21767,N_21988);
nand U22622 (N_22622,N_21934,N_21779);
and U22623 (N_22623,N_21634,N_21773);
xor U22624 (N_22624,N_21870,N_22082);
nor U22625 (N_22625,N_21685,N_21914);
xor U22626 (N_22626,N_22193,N_21911);
xor U22627 (N_22627,N_21657,N_22138);
nor U22628 (N_22628,N_22109,N_22060);
xnor U22629 (N_22629,N_21748,N_22095);
nor U22630 (N_22630,N_22138,N_21999);
xor U22631 (N_22631,N_21852,N_22159);
nor U22632 (N_22632,N_22172,N_21988);
nor U22633 (N_22633,N_21743,N_21899);
or U22634 (N_22634,N_21953,N_21790);
or U22635 (N_22635,N_21920,N_22114);
xnor U22636 (N_22636,N_21853,N_21883);
and U22637 (N_22637,N_21865,N_22124);
or U22638 (N_22638,N_21811,N_22170);
and U22639 (N_22639,N_21903,N_21804);
and U22640 (N_22640,N_22141,N_21705);
or U22641 (N_22641,N_22110,N_21986);
xor U22642 (N_22642,N_21822,N_22101);
xor U22643 (N_22643,N_21927,N_22004);
and U22644 (N_22644,N_21639,N_22145);
nor U22645 (N_22645,N_21938,N_22092);
and U22646 (N_22646,N_21738,N_22091);
nand U22647 (N_22647,N_21818,N_22141);
nor U22648 (N_22648,N_21602,N_21805);
xnor U22649 (N_22649,N_21746,N_21890);
nor U22650 (N_22650,N_21994,N_22070);
nor U22651 (N_22651,N_21861,N_21641);
and U22652 (N_22652,N_22100,N_21660);
and U22653 (N_22653,N_21809,N_21858);
xnor U22654 (N_22654,N_21762,N_21677);
or U22655 (N_22655,N_21937,N_22185);
or U22656 (N_22656,N_21799,N_21756);
nand U22657 (N_22657,N_22172,N_22002);
or U22658 (N_22658,N_22095,N_21609);
nor U22659 (N_22659,N_22048,N_21614);
or U22660 (N_22660,N_21958,N_21839);
nand U22661 (N_22661,N_22118,N_21621);
or U22662 (N_22662,N_21608,N_21739);
xnor U22663 (N_22663,N_21845,N_22033);
nand U22664 (N_22664,N_21834,N_22077);
and U22665 (N_22665,N_22133,N_21797);
or U22666 (N_22666,N_22152,N_21861);
xnor U22667 (N_22667,N_22106,N_21902);
and U22668 (N_22668,N_21673,N_21862);
xor U22669 (N_22669,N_21825,N_21829);
and U22670 (N_22670,N_21772,N_21750);
nand U22671 (N_22671,N_22123,N_21886);
nor U22672 (N_22672,N_21669,N_21981);
nand U22673 (N_22673,N_21820,N_21754);
nor U22674 (N_22674,N_21721,N_21919);
nand U22675 (N_22675,N_22025,N_21613);
or U22676 (N_22676,N_21725,N_22122);
nand U22677 (N_22677,N_21977,N_21759);
nor U22678 (N_22678,N_21909,N_22073);
nand U22679 (N_22679,N_22183,N_22175);
or U22680 (N_22680,N_21799,N_22091);
or U22681 (N_22681,N_21900,N_21718);
and U22682 (N_22682,N_21627,N_22158);
and U22683 (N_22683,N_21734,N_21702);
and U22684 (N_22684,N_21774,N_21743);
nor U22685 (N_22685,N_21752,N_22041);
nor U22686 (N_22686,N_22041,N_22167);
nand U22687 (N_22687,N_21818,N_21815);
nor U22688 (N_22688,N_21821,N_21629);
nand U22689 (N_22689,N_22083,N_22132);
and U22690 (N_22690,N_21627,N_21977);
xor U22691 (N_22691,N_21800,N_21910);
nand U22692 (N_22692,N_21648,N_22036);
xnor U22693 (N_22693,N_21983,N_22144);
or U22694 (N_22694,N_21779,N_21750);
xor U22695 (N_22695,N_21885,N_21986);
and U22696 (N_22696,N_21965,N_21797);
and U22697 (N_22697,N_22021,N_22105);
nand U22698 (N_22698,N_21954,N_21686);
nor U22699 (N_22699,N_21850,N_21742);
and U22700 (N_22700,N_21944,N_21711);
and U22701 (N_22701,N_22006,N_21664);
xnor U22702 (N_22702,N_21745,N_22135);
nor U22703 (N_22703,N_21928,N_21706);
or U22704 (N_22704,N_22126,N_21842);
xor U22705 (N_22705,N_21651,N_22123);
nor U22706 (N_22706,N_21623,N_21722);
or U22707 (N_22707,N_22033,N_22134);
and U22708 (N_22708,N_22134,N_21641);
xnor U22709 (N_22709,N_22001,N_21927);
nand U22710 (N_22710,N_22031,N_21971);
nand U22711 (N_22711,N_22096,N_21949);
xor U22712 (N_22712,N_21754,N_21756);
nor U22713 (N_22713,N_22110,N_21770);
xor U22714 (N_22714,N_21714,N_22046);
and U22715 (N_22715,N_22044,N_21672);
and U22716 (N_22716,N_21891,N_21949);
and U22717 (N_22717,N_21849,N_21725);
nor U22718 (N_22718,N_22010,N_21949);
and U22719 (N_22719,N_21865,N_22127);
nor U22720 (N_22720,N_21685,N_21709);
and U22721 (N_22721,N_21670,N_21819);
and U22722 (N_22722,N_21874,N_21972);
xor U22723 (N_22723,N_21634,N_22163);
nand U22724 (N_22724,N_21639,N_21736);
or U22725 (N_22725,N_21655,N_21992);
nand U22726 (N_22726,N_21678,N_21766);
nor U22727 (N_22727,N_21808,N_21749);
xor U22728 (N_22728,N_21767,N_21738);
nand U22729 (N_22729,N_21928,N_22108);
and U22730 (N_22730,N_21674,N_21901);
and U22731 (N_22731,N_21959,N_21769);
and U22732 (N_22732,N_21947,N_21687);
xor U22733 (N_22733,N_21642,N_21921);
nand U22734 (N_22734,N_21808,N_21948);
and U22735 (N_22735,N_21942,N_21878);
nand U22736 (N_22736,N_21994,N_21902);
nand U22737 (N_22737,N_21693,N_21999);
nor U22738 (N_22738,N_21626,N_21680);
xor U22739 (N_22739,N_21983,N_22000);
or U22740 (N_22740,N_21800,N_21994);
xor U22741 (N_22741,N_21859,N_21773);
nor U22742 (N_22742,N_22067,N_21949);
nor U22743 (N_22743,N_22155,N_21779);
nand U22744 (N_22744,N_21801,N_21789);
xor U22745 (N_22745,N_21830,N_22040);
xor U22746 (N_22746,N_22016,N_21615);
nor U22747 (N_22747,N_22047,N_22161);
nand U22748 (N_22748,N_21960,N_21907);
and U22749 (N_22749,N_21725,N_21937);
nand U22750 (N_22750,N_22164,N_21821);
nand U22751 (N_22751,N_22013,N_21872);
nand U22752 (N_22752,N_21894,N_21984);
xor U22753 (N_22753,N_21683,N_21890);
nand U22754 (N_22754,N_21911,N_22005);
xnor U22755 (N_22755,N_21774,N_21909);
nand U22756 (N_22756,N_21898,N_21790);
nand U22757 (N_22757,N_21699,N_21662);
or U22758 (N_22758,N_21706,N_21830);
nand U22759 (N_22759,N_22069,N_22097);
nand U22760 (N_22760,N_22174,N_21861);
and U22761 (N_22761,N_21646,N_22102);
xor U22762 (N_22762,N_22177,N_21913);
xnor U22763 (N_22763,N_21650,N_21640);
nor U22764 (N_22764,N_21945,N_22071);
and U22765 (N_22765,N_22012,N_21760);
nor U22766 (N_22766,N_21942,N_21692);
and U22767 (N_22767,N_22112,N_21710);
or U22768 (N_22768,N_22035,N_21801);
nand U22769 (N_22769,N_21948,N_22062);
and U22770 (N_22770,N_22085,N_22180);
or U22771 (N_22771,N_21856,N_21617);
or U22772 (N_22772,N_21954,N_21628);
or U22773 (N_22773,N_21796,N_22078);
nand U22774 (N_22774,N_21987,N_21720);
and U22775 (N_22775,N_22174,N_21969);
xor U22776 (N_22776,N_21760,N_22130);
or U22777 (N_22777,N_22053,N_21779);
nor U22778 (N_22778,N_21979,N_21694);
and U22779 (N_22779,N_21665,N_21998);
or U22780 (N_22780,N_21955,N_21666);
xor U22781 (N_22781,N_21883,N_22022);
nor U22782 (N_22782,N_21778,N_22045);
or U22783 (N_22783,N_22083,N_21747);
xnor U22784 (N_22784,N_22174,N_21965);
or U22785 (N_22785,N_21832,N_21729);
or U22786 (N_22786,N_22137,N_22146);
nor U22787 (N_22787,N_22076,N_21781);
and U22788 (N_22788,N_21960,N_21824);
nor U22789 (N_22789,N_21756,N_21969);
xnor U22790 (N_22790,N_21777,N_21844);
and U22791 (N_22791,N_21617,N_21849);
or U22792 (N_22792,N_22175,N_22132);
and U22793 (N_22793,N_22182,N_21889);
nand U22794 (N_22794,N_21840,N_21960);
nand U22795 (N_22795,N_21936,N_22091);
xor U22796 (N_22796,N_21844,N_21933);
and U22797 (N_22797,N_21748,N_21798);
xnor U22798 (N_22798,N_21860,N_21729);
nand U22799 (N_22799,N_22130,N_22132);
xnor U22800 (N_22800,N_22702,N_22323);
and U22801 (N_22801,N_22455,N_22428);
or U22802 (N_22802,N_22623,N_22287);
xor U22803 (N_22803,N_22424,N_22570);
xnor U22804 (N_22804,N_22648,N_22572);
nand U22805 (N_22805,N_22232,N_22320);
xnor U22806 (N_22806,N_22466,N_22574);
or U22807 (N_22807,N_22666,N_22449);
xnor U22808 (N_22808,N_22334,N_22563);
nor U22809 (N_22809,N_22504,N_22625);
xnor U22810 (N_22810,N_22763,N_22213);
nand U22811 (N_22811,N_22452,N_22490);
or U22812 (N_22812,N_22719,N_22674);
xor U22813 (N_22813,N_22523,N_22367);
xor U22814 (N_22814,N_22537,N_22283);
nand U22815 (N_22815,N_22661,N_22254);
xor U22816 (N_22816,N_22778,N_22344);
and U22817 (N_22817,N_22549,N_22796);
and U22818 (N_22818,N_22772,N_22352);
nor U22819 (N_22819,N_22407,N_22732);
nor U22820 (N_22820,N_22280,N_22225);
or U22821 (N_22821,N_22598,N_22451);
nor U22822 (N_22822,N_22429,N_22382);
nand U22823 (N_22823,N_22212,N_22560);
or U22824 (N_22824,N_22445,N_22418);
xor U22825 (N_22825,N_22370,N_22681);
and U22826 (N_22826,N_22359,N_22410);
nand U22827 (N_22827,N_22608,N_22353);
xnor U22828 (N_22828,N_22652,N_22491);
and U22829 (N_22829,N_22383,N_22745);
and U22830 (N_22830,N_22618,N_22337);
and U22831 (N_22831,N_22708,N_22580);
nand U22832 (N_22832,N_22274,N_22416);
nand U22833 (N_22833,N_22567,N_22789);
nand U22834 (N_22834,N_22326,N_22715);
or U22835 (N_22835,N_22516,N_22612);
and U22836 (N_22836,N_22725,N_22253);
or U22837 (N_22837,N_22436,N_22741);
nor U22838 (N_22838,N_22750,N_22602);
or U22839 (N_22839,N_22768,N_22622);
nor U22840 (N_22840,N_22378,N_22300);
or U22841 (N_22841,N_22659,N_22203);
xor U22842 (N_22842,N_22356,N_22527);
xnor U22843 (N_22843,N_22722,N_22564);
nor U22844 (N_22844,N_22311,N_22538);
or U22845 (N_22845,N_22517,N_22706);
or U22846 (N_22846,N_22403,N_22400);
nor U22847 (N_22847,N_22626,N_22257);
nand U22848 (N_22848,N_22374,N_22228);
and U22849 (N_22849,N_22209,N_22554);
xor U22850 (N_22850,N_22506,N_22686);
or U22851 (N_22851,N_22372,N_22373);
or U22852 (N_22852,N_22649,N_22781);
nand U22853 (N_22853,N_22525,N_22774);
and U22854 (N_22854,N_22733,N_22237);
and U22855 (N_22855,N_22476,N_22399);
or U22856 (N_22856,N_22728,N_22753);
or U22857 (N_22857,N_22278,N_22387);
xnor U22858 (N_22858,N_22575,N_22521);
nand U22859 (N_22859,N_22683,N_22543);
or U22860 (N_22860,N_22559,N_22611);
xnor U22861 (N_22861,N_22555,N_22472);
or U22862 (N_22862,N_22247,N_22454);
and U22863 (N_22863,N_22251,N_22229);
xnor U22864 (N_22864,N_22531,N_22680);
or U22865 (N_22865,N_22737,N_22204);
xnor U22866 (N_22866,N_22477,N_22634);
nor U22867 (N_22867,N_22261,N_22388);
or U22868 (N_22868,N_22246,N_22565);
nand U22869 (N_22869,N_22718,N_22364);
nor U22870 (N_22870,N_22566,N_22233);
nand U22871 (N_22871,N_22430,N_22499);
or U22872 (N_22872,N_22709,N_22316);
and U22873 (N_22873,N_22534,N_22606);
and U22874 (N_22874,N_22262,N_22200);
nor U22875 (N_22875,N_22519,N_22294);
xor U22876 (N_22876,N_22551,N_22628);
or U22877 (N_22877,N_22640,N_22758);
and U22878 (N_22878,N_22583,N_22295);
or U22879 (N_22879,N_22780,N_22770);
nand U22880 (N_22880,N_22779,N_22284);
xnor U22881 (N_22881,N_22665,N_22302);
nor U22882 (N_22882,N_22275,N_22214);
and U22883 (N_22883,N_22577,N_22614);
nor U22884 (N_22884,N_22217,N_22569);
nand U22885 (N_22885,N_22390,N_22518);
xor U22886 (N_22886,N_22647,N_22546);
and U22887 (N_22887,N_22272,N_22775);
nand U22888 (N_22888,N_22720,N_22699);
nand U22889 (N_22889,N_22593,N_22432);
nor U22890 (N_22890,N_22268,N_22201);
nor U22891 (N_22891,N_22426,N_22646);
nand U22892 (N_22892,N_22524,N_22279);
and U22893 (N_22893,N_22401,N_22587);
or U22894 (N_22894,N_22662,N_22724);
and U22895 (N_22895,N_22713,N_22277);
or U22896 (N_22896,N_22288,N_22485);
and U22897 (N_22897,N_22696,N_22548);
and U22898 (N_22898,N_22714,N_22791);
or U22899 (N_22899,N_22306,N_22742);
xnor U22900 (N_22900,N_22630,N_22743);
and U22901 (N_22901,N_22363,N_22433);
xnor U22902 (N_22902,N_22371,N_22589);
or U22903 (N_22903,N_22496,N_22557);
or U22904 (N_22904,N_22729,N_22245);
xor U22905 (N_22905,N_22438,N_22369);
xor U22906 (N_22906,N_22776,N_22619);
xor U22907 (N_22907,N_22480,N_22329);
nor U22908 (N_22908,N_22206,N_22345);
and U22909 (N_22909,N_22324,N_22486);
nand U22910 (N_22910,N_22797,N_22785);
nor U22911 (N_22911,N_22461,N_22421);
nor U22912 (N_22912,N_22473,N_22297);
or U22913 (N_22913,N_22641,N_22793);
xor U22914 (N_22914,N_22705,N_22435);
xor U22915 (N_22915,N_22457,N_22375);
and U22916 (N_22916,N_22230,N_22511);
nand U22917 (N_22917,N_22467,N_22483);
or U22918 (N_22918,N_22735,N_22386);
nand U22919 (N_22919,N_22777,N_22604);
nor U22920 (N_22920,N_22597,N_22520);
or U22921 (N_22921,N_22547,N_22500);
and U22922 (N_22922,N_22234,N_22571);
xnor U22923 (N_22923,N_22515,N_22226);
nand U22924 (N_22924,N_22631,N_22498);
nand U22925 (N_22925,N_22299,N_22795);
nor U22926 (N_22926,N_22761,N_22282);
and U22927 (N_22927,N_22409,N_22687);
nor U22928 (N_22928,N_22423,N_22317);
nor U22929 (N_22929,N_22405,N_22769);
nand U22930 (N_22930,N_22248,N_22624);
or U22931 (N_22931,N_22545,N_22727);
nand U22932 (N_22932,N_22322,N_22503);
and U22933 (N_22933,N_22752,N_22269);
or U22934 (N_22934,N_22760,N_22258);
nor U22935 (N_22935,N_22292,N_22573);
xor U22936 (N_22936,N_22354,N_22310);
and U22937 (N_22937,N_22585,N_22717);
nor U22938 (N_22938,N_22787,N_22747);
or U22939 (N_22939,N_22601,N_22495);
nand U22940 (N_22940,N_22227,N_22544);
nor U22941 (N_22941,N_22402,N_22734);
and U22942 (N_22942,N_22319,N_22756);
and U22943 (N_22943,N_22347,N_22252);
nand U22944 (N_22944,N_22450,N_22790);
and U22945 (N_22945,N_22568,N_22783);
xor U22946 (N_22946,N_22341,N_22362);
nand U22947 (N_22947,N_22798,N_22693);
and U22948 (N_22948,N_22427,N_22417);
xor U22949 (N_22949,N_22443,N_22526);
or U22950 (N_22950,N_22398,N_22672);
xnor U22951 (N_22951,N_22629,N_22657);
and U22952 (N_22952,N_22749,N_22255);
nor U22953 (N_22953,N_22420,N_22238);
nor U22954 (N_22954,N_22671,N_22459);
nor U22955 (N_22955,N_22360,N_22757);
and U22956 (N_22956,N_22408,N_22469);
nor U22957 (N_22957,N_22730,N_22670);
xor U22958 (N_22958,N_22723,N_22361);
nor U22959 (N_22959,N_22348,N_22357);
nand U22960 (N_22960,N_22609,N_22210);
nand U22961 (N_22961,N_22350,N_22256);
xor U22962 (N_22962,N_22250,N_22677);
nand U22963 (N_22963,N_22249,N_22532);
and U22964 (N_22964,N_22607,N_22340);
nor U22965 (N_22965,N_22484,N_22638);
and U22966 (N_22966,N_22492,N_22312);
or U22967 (N_22967,N_22271,N_22765);
xnor U22968 (N_22968,N_22773,N_22578);
or U22969 (N_22969,N_22509,N_22539);
nand U22970 (N_22970,N_22782,N_22298);
nor U22971 (N_22971,N_22296,N_22381);
or U22972 (N_22972,N_22599,N_22366);
and U22973 (N_22973,N_22605,N_22510);
and U22974 (N_22974,N_22642,N_22639);
nor U22975 (N_22975,N_22712,N_22707);
xor U22976 (N_22976,N_22422,N_22305);
and U22977 (N_22977,N_22654,N_22658);
and U22978 (N_22978,N_22241,N_22487);
xor U22979 (N_22979,N_22281,N_22441);
and U22980 (N_22980,N_22235,N_22505);
xor U22981 (N_22981,N_22412,N_22703);
nand U22982 (N_22982,N_22692,N_22309);
nand U22983 (N_22983,N_22285,N_22293);
nor U22984 (N_22984,N_22220,N_22389);
nand U22985 (N_22985,N_22541,N_22444);
or U22986 (N_22986,N_22384,N_22231);
and U22987 (N_22987,N_22447,N_22411);
nand U22988 (N_22988,N_22488,N_22478);
or U22989 (N_22989,N_22704,N_22327);
nand U22990 (N_22990,N_22380,N_22202);
nor U22991 (N_22991,N_22244,N_22437);
xnor U22992 (N_22992,N_22385,N_22465);
and U22993 (N_22993,N_22695,N_22222);
xnor U22994 (N_22994,N_22346,N_22304);
nor U22995 (N_22995,N_22243,N_22394);
and U22996 (N_22996,N_22600,N_22470);
or U22997 (N_22997,N_22205,N_22731);
nor U22998 (N_22998,N_22318,N_22536);
nand U22999 (N_22999,N_22425,N_22603);
nand U23000 (N_23000,N_22512,N_22377);
xnor U23001 (N_23001,N_22396,N_22682);
or U23002 (N_23002,N_22542,N_22358);
and U23003 (N_23003,N_22522,N_22588);
and U23004 (N_23004,N_22751,N_22215);
and U23005 (N_23005,N_22754,N_22794);
xor U23006 (N_23006,N_22489,N_22664);
and U23007 (N_23007,N_22415,N_22270);
xnor U23008 (N_23008,N_22471,N_22307);
or U23009 (N_23009,N_22540,N_22239);
nand U23010 (N_23010,N_22482,N_22463);
nand U23011 (N_23011,N_22721,N_22335);
and U23012 (N_23012,N_22656,N_22637);
or U23013 (N_23013,N_22627,N_22332);
nand U23014 (N_23014,N_22303,N_22576);
nand U23015 (N_23015,N_22259,N_22330);
xor U23016 (N_23016,N_22739,N_22550);
and U23017 (N_23017,N_22221,N_22660);
or U23018 (N_23018,N_22558,N_22468);
xor U23019 (N_23019,N_22351,N_22328);
nor U23020 (N_23020,N_22655,N_22442);
nor U23021 (N_23021,N_22528,N_22265);
or U23022 (N_23022,N_22592,N_22616);
xnor U23023 (N_23023,N_22208,N_22759);
xor U23024 (N_23024,N_22736,N_22501);
and U23025 (N_23025,N_22448,N_22644);
or U23026 (N_23026,N_22404,N_22650);
or U23027 (N_23027,N_22218,N_22494);
xnor U23028 (N_23028,N_22207,N_22349);
or U23029 (N_23029,N_22553,N_22475);
xnor U23030 (N_23030,N_22762,N_22533);
xnor U23031 (N_23031,N_22236,N_22746);
xor U23032 (N_23032,N_22325,N_22508);
and U23033 (N_23033,N_22273,N_22513);
or U23034 (N_23034,N_22635,N_22529);
or U23035 (N_23035,N_22764,N_22771);
nand U23036 (N_23036,N_22679,N_22391);
or U23037 (N_23037,N_22700,N_22434);
or U23038 (N_23038,N_22651,N_22342);
nand U23039 (N_23039,N_22698,N_22633);
nand U23040 (N_23040,N_22767,N_22610);
and U23041 (N_23041,N_22308,N_22621);
and U23042 (N_23042,N_22474,N_22458);
or U23043 (N_23043,N_22581,N_22395);
or U23044 (N_23044,N_22464,N_22643);
nand U23045 (N_23045,N_22701,N_22440);
xor U23046 (N_23046,N_22788,N_22343);
xor U23047 (N_23047,N_22688,N_22419);
nor U23048 (N_23048,N_22211,N_22414);
and U23049 (N_23049,N_22406,N_22333);
nand U23050 (N_23050,N_22615,N_22336);
and U23051 (N_23051,N_22667,N_22591);
xnor U23052 (N_23052,N_22338,N_22596);
and U23053 (N_23053,N_22514,N_22266);
nor U23054 (N_23054,N_22240,N_22590);
nand U23055 (N_23055,N_22497,N_22276);
nand U23056 (N_23056,N_22691,N_22579);
nor U23057 (N_23057,N_22339,N_22697);
nor U23058 (N_23058,N_22711,N_22613);
nand U23059 (N_23059,N_22223,N_22552);
and U23060 (N_23060,N_22690,N_22291);
nor U23061 (N_23061,N_22446,N_22726);
nand U23062 (N_23062,N_22586,N_22582);
xor U23063 (N_23063,N_22289,N_22784);
xor U23064 (N_23064,N_22556,N_22355);
nor U23065 (N_23065,N_22594,N_22632);
nand U23066 (N_23066,N_22313,N_22331);
and U23067 (N_23067,N_22493,N_22479);
nand U23068 (N_23068,N_22748,N_22595);
nand U23069 (N_23069,N_22620,N_22755);
and U23070 (N_23070,N_22264,N_22507);
nand U23071 (N_23071,N_22684,N_22397);
nor U23072 (N_23072,N_22219,N_22716);
and U23073 (N_23073,N_22799,N_22456);
nor U23074 (N_23074,N_22766,N_22413);
and U23075 (N_23075,N_22694,N_22584);
nor U23076 (N_23076,N_22676,N_22321);
and U23077 (N_23077,N_22675,N_22617);
nor U23078 (N_23078,N_22535,N_22653);
and U23079 (N_23079,N_22744,N_22453);
nand U23080 (N_23080,N_22286,N_22260);
nor U23081 (N_23081,N_22267,N_22669);
nand U23082 (N_23082,N_22431,N_22786);
xnor U23083 (N_23083,N_22530,N_22224);
nor U23084 (N_23084,N_22636,N_22376);
nand U23085 (N_23085,N_22710,N_22392);
nor U23086 (N_23086,N_22738,N_22393);
and U23087 (N_23087,N_22365,N_22685);
or U23088 (N_23088,N_22645,N_22242);
xor U23089 (N_23089,N_22481,N_22792);
xor U23090 (N_23090,N_22502,N_22689);
xnor U23091 (N_23091,N_22379,N_22663);
nor U23092 (N_23092,N_22561,N_22668);
or U23093 (N_23093,N_22439,N_22301);
nand U23094 (N_23094,N_22562,N_22678);
nor U23095 (N_23095,N_22460,N_22740);
xnor U23096 (N_23096,N_22462,N_22263);
nand U23097 (N_23097,N_22673,N_22290);
and U23098 (N_23098,N_22368,N_22314);
and U23099 (N_23099,N_22216,N_22315);
or U23100 (N_23100,N_22595,N_22472);
nand U23101 (N_23101,N_22404,N_22474);
xnor U23102 (N_23102,N_22666,N_22702);
or U23103 (N_23103,N_22794,N_22498);
or U23104 (N_23104,N_22344,N_22637);
nor U23105 (N_23105,N_22527,N_22310);
nand U23106 (N_23106,N_22227,N_22714);
or U23107 (N_23107,N_22337,N_22344);
or U23108 (N_23108,N_22278,N_22705);
and U23109 (N_23109,N_22616,N_22720);
and U23110 (N_23110,N_22743,N_22476);
and U23111 (N_23111,N_22694,N_22703);
xor U23112 (N_23112,N_22242,N_22369);
xnor U23113 (N_23113,N_22419,N_22451);
nand U23114 (N_23114,N_22726,N_22669);
nor U23115 (N_23115,N_22237,N_22621);
or U23116 (N_23116,N_22658,N_22586);
nor U23117 (N_23117,N_22677,N_22732);
nand U23118 (N_23118,N_22579,N_22789);
and U23119 (N_23119,N_22462,N_22674);
nor U23120 (N_23120,N_22298,N_22598);
nand U23121 (N_23121,N_22649,N_22728);
xor U23122 (N_23122,N_22430,N_22324);
xor U23123 (N_23123,N_22253,N_22358);
nor U23124 (N_23124,N_22563,N_22504);
and U23125 (N_23125,N_22429,N_22591);
nand U23126 (N_23126,N_22561,N_22275);
and U23127 (N_23127,N_22774,N_22713);
or U23128 (N_23128,N_22520,N_22684);
xor U23129 (N_23129,N_22421,N_22714);
nand U23130 (N_23130,N_22513,N_22719);
nor U23131 (N_23131,N_22316,N_22543);
nand U23132 (N_23132,N_22598,N_22521);
nor U23133 (N_23133,N_22506,N_22500);
nor U23134 (N_23134,N_22308,N_22297);
or U23135 (N_23135,N_22701,N_22569);
or U23136 (N_23136,N_22563,N_22705);
nor U23137 (N_23137,N_22333,N_22543);
xnor U23138 (N_23138,N_22595,N_22651);
nor U23139 (N_23139,N_22778,N_22772);
and U23140 (N_23140,N_22460,N_22584);
xnor U23141 (N_23141,N_22663,N_22475);
or U23142 (N_23142,N_22534,N_22224);
nand U23143 (N_23143,N_22239,N_22260);
or U23144 (N_23144,N_22741,N_22760);
nand U23145 (N_23145,N_22598,N_22353);
nand U23146 (N_23146,N_22418,N_22285);
xnor U23147 (N_23147,N_22657,N_22679);
nand U23148 (N_23148,N_22300,N_22600);
nand U23149 (N_23149,N_22652,N_22534);
xnor U23150 (N_23150,N_22468,N_22262);
nor U23151 (N_23151,N_22298,N_22449);
nand U23152 (N_23152,N_22645,N_22490);
and U23153 (N_23153,N_22684,N_22512);
and U23154 (N_23154,N_22408,N_22200);
and U23155 (N_23155,N_22417,N_22278);
nor U23156 (N_23156,N_22693,N_22635);
and U23157 (N_23157,N_22543,N_22340);
or U23158 (N_23158,N_22765,N_22620);
or U23159 (N_23159,N_22273,N_22284);
and U23160 (N_23160,N_22502,N_22538);
xor U23161 (N_23161,N_22411,N_22688);
xnor U23162 (N_23162,N_22649,N_22501);
nor U23163 (N_23163,N_22639,N_22660);
nor U23164 (N_23164,N_22317,N_22379);
xnor U23165 (N_23165,N_22407,N_22214);
nor U23166 (N_23166,N_22522,N_22317);
and U23167 (N_23167,N_22431,N_22272);
nand U23168 (N_23168,N_22625,N_22546);
xor U23169 (N_23169,N_22741,N_22329);
nor U23170 (N_23170,N_22314,N_22603);
nor U23171 (N_23171,N_22401,N_22379);
nor U23172 (N_23172,N_22770,N_22250);
nand U23173 (N_23173,N_22253,N_22592);
nor U23174 (N_23174,N_22707,N_22723);
nand U23175 (N_23175,N_22479,N_22697);
and U23176 (N_23176,N_22756,N_22667);
nand U23177 (N_23177,N_22707,N_22762);
or U23178 (N_23178,N_22607,N_22355);
nor U23179 (N_23179,N_22546,N_22719);
nor U23180 (N_23180,N_22202,N_22623);
nand U23181 (N_23181,N_22459,N_22732);
nor U23182 (N_23182,N_22227,N_22422);
nand U23183 (N_23183,N_22278,N_22659);
and U23184 (N_23184,N_22295,N_22727);
xnor U23185 (N_23185,N_22763,N_22387);
xnor U23186 (N_23186,N_22728,N_22351);
and U23187 (N_23187,N_22711,N_22313);
nor U23188 (N_23188,N_22452,N_22407);
or U23189 (N_23189,N_22408,N_22571);
nand U23190 (N_23190,N_22545,N_22319);
nor U23191 (N_23191,N_22592,N_22335);
and U23192 (N_23192,N_22570,N_22416);
or U23193 (N_23193,N_22513,N_22369);
nor U23194 (N_23194,N_22395,N_22551);
nand U23195 (N_23195,N_22267,N_22790);
nor U23196 (N_23196,N_22276,N_22645);
and U23197 (N_23197,N_22665,N_22624);
nor U23198 (N_23198,N_22486,N_22367);
and U23199 (N_23199,N_22735,N_22207);
nand U23200 (N_23200,N_22703,N_22231);
nand U23201 (N_23201,N_22408,N_22750);
or U23202 (N_23202,N_22675,N_22529);
or U23203 (N_23203,N_22688,N_22467);
nor U23204 (N_23204,N_22240,N_22379);
xor U23205 (N_23205,N_22269,N_22700);
or U23206 (N_23206,N_22498,N_22336);
xnor U23207 (N_23207,N_22203,N_22291);
or U23208 (N_23208,N_22454,N_22532);
nor U23209 (N_23209,N_22627,N_22330);
nand U23210 (N_23210,N_22401,N_22293);
or U23211 (N_23211,N_22358,N_22399);
xor U23212 (N_23212,N_22303,N_22596);
nand U23213 (N_23213,N_22411,N_22637);
xnor U23214 (N_23214,N_22702,N_22782);
nand U23215 (N_23215,N_22212,N_22231);
nor U23216 (N_23216,N_22764,N_22443);
nand U23217 (N_23217,N_22683,N_22513);
or U23218 (N_23218,N_22477,N_22330);
and U23219 (N_23219,N_22757,N_22525);
and U23220 (N_23220,N_22668,N_22443);
and U23221 (N_23221,N_22238,N_22326);
nor U23222 (N_23222,N_22430,N_22662);
and U23223 (N_23223,N_22589,N_22561);
nand U23224 (N_23224,N_22780,N_22448);
nand U23225 (N_23225,N_22264,N_22523);
xor U23226 (N_23226,N_22787,N_22320);
and U23227 (N_23227,N_22622,N_22378);
or U23228 (N_23228,N_22507,N_22471);
xor U23229 (N_23229,N_22583,N_22206);
and U23230 (N_23230,N_22612,N_22694);
nor U23231 (N_23231,N_22285,N_22277);
xor U23232 (N_23232,N_22600,N_22253);
and U23233 (N_23233,N_22339,N_22773);
xor U23234 (N_23234,N_22585,N_22218);
or U23235 (N_23235,N_22238,N_22630);
and U23236 (N_23236,N_22346,N_22275);
nor U23237 (N_23237,N_22734,N_22612);
nand U23238 (N_23238,N_22569,N_22653);
xnor U23239 (N_23239,N_22337,N_22530);
nand U23240 (N_23240,N_22569,N_22568);
nor U23241 (N_23241,N_22648,N_22408);
nand U23242 (N_23242,N_22591,N_22341);
or U23243 (N_23243,N_22713,N_22566);
nand U23244 (N_23244,N_22225,N_22201);
and U23245 (N_23245,N_22297,N_22503);
or U23246 (N_23246,N_22249,N_22713);
nor U23247 (N_23247,N_22793,N_22420);
and U23248 (N_23248,N_22722,N_22254);
xor U23249 (N_23249,N_22389,N_22782);
or U23250 (N_23250,N_22588,N_22544);
nand U23251 (N_23251,N_22683,N_22416);
xor U23252 (N_23252,N_22516,N_22413);
nor U23253 (N_23253,N_22443,N_22543);
nand U23254 (N_23254,N_22763,N_22557);
xor U23255 (N_23255,N_22647,N_22430);
nand U23256 (N_23256,N_22358,N_22498);
or U23257 (N_23257,N_22687,N_22390);
nand U23258 (N_23258,N_22503,N_22686);
xnor U23259 (N_23259,N_22695,N_22405);
nor U23260 (N_23260,N_22703,N_22418);
xnor U23261 (N_23261,N_22497,N_22740);
nor U23262 (N_23262,N_22730,N_22416);
nand U23263 (N_23263,N_22751,N_22622);
and U23264 (N_23264,N_22280,N_22330);
nand U23265 (N_23265,N_22618,N_22377);
xor U23266 (N_23266,N_22574,N_22551);
xnor U23267 (N_23267,N_22263,N_22463);
or U23268 (N_23268,N_22259,N_22606);
xor U23269 (N_23269,N_22217,N_22563);
xor U23270 (N_23270,N_22453,N_22570);
or U23271 (N_23271,N_22533,N_22353);
xor U23272 (N_23272,N_22360,N_22487);
and U23273 (N_23273,N_22421,N_22666);
nand U23274 (N_23274,N_22300,N_22271);
or U23275 (N_23275,N_22738,N_22762);
xor U23276 (N_23276,N_22705,N_22283);
nand U23277 (N_23277,N_22515,N_22664);
xnor U23278 (N_23278,N_22324,N_22709);
nand U23279 (N_23279,N_22711,N_22465);
xnor U23280 (N_23280,N_22364,N_22608);
and U23281 (N_23281,N_22598,N_22582);
nand U23282 (N_23282,N_22674,N_22539);
nor U23283 (N_23283,N_22509,N_22608);
nor U23284 (N_23284,N_22777,N_22367);
or U23285 (N_23285,N_22670,N_22640);
nand U23286 (N_23286,N_22501,N_22532);
nand U23287 (N_23287,N_22558,N_22282);
or U23288 (N_23288,N_22650,N_22709);
xnor U23289 (N_23289,N_22309,N_22344);
and U23290 (N_23290,N_22725,N_22500);
or U23291 (N_23291,N_22652,N_22346);
nand U23292 (N_23292,N_22503,N_22424);
xor U23293 (N_23293,N_22776,N_22762);
xnor U23294 (N_23294,N_22738,N_22291);
nand U23295 (N_23295,N_22593,N_22316);
and U23296 (N_23296,N_22456,N_22361);
and U23297 (N_23297,N_22364,N_22604);
or U23298 (N_23298,N_22427,N_22366);
and U23299 (N_23299,N_22515,N_22731);
xor U23300 (N_23300,N_22714,N_22284);
nand U23301 (N_23301,N_22417,N_22548);
nand U23302 (N_23302,N_22487,N_22758);
or U23303 (N_23303,N_22413,N_22231);
nand U23304 (N_23304,N_22633,N_22531);
or U23305 (N_23305,N_22294,N_22760);
xnor U23306 (N_23306,N_22299,N_22394);
and U23307 (N_23307,N_22746,N_22528);
nor U23308 (N_23308,N_22350,N_22371);
nand U23309 (N_23309,N_22612,N_22209);
or U23310 (N_23310,N_22695,N_22365);
xor U23311 (N_23311,N_22758,N_22282);
and U23312 (N_23312,N_22769,N_22381);
nor U23313 (N_23313,N_22789,N_22554);
xor U23314 (N_23314,N_22466,N_22495);
xnor U23315 (N_23315,N_22666,N_22412);
xor U23316 (N_23316,N_22690,N_22714);
nor U23317 (N_23317,N_22262,N_22589);
xor U23318 (N_23318,N_22796,N_22255);
xnor U23319 (N_23319,N_22488,N_22685);
nand U23320 (N_23320,N_22229,N_22486);
or U23321 (N_23321,N_22749,N_22320);
nand U23322 (N_23322,N_22782,N_22277);
or U23323 (N_23323,N_22765,N_22663);
nor U23324 (N_23324,N_22672,N_22302);
and U23325 (N_23325,N_22578,N_22737);
or U23326 (N_23326,N_22788,N_22358);
xnor U23327 (N_23327,N_22793,N_22785);
or U23328 (N_23328,N_22651,N_22485);
nand U23329 (N_23329,N_22347,N_22294);
nand U23330 (N_23330,N_22422,N_22315);
nor U23331 (N_23331,N_22483,N_22397);
or U23332 (N_23332,N_22306,N_22585);
xnor U23333 (N_23333,N_22495,N_22627);
xnor U23334 (N_23334,N_22470,N_22273);
nand U23335 (N_23335,N_22564,N_22200);
xor U23336 (N_23336,N_22699,N_22331);
or U23337 (N_23337,N_22464,N_22720);
xnor U23338 (N_23338,N_22416,N_22279);
or U23339 (N_23339,N_22294,N_22446);
or U23340 (N_23340,N_22611,N_22680);
nor U23341 (N_23341,N_22441,N_22710);
and U23342 (N_23342,N_22314,N_22780);
nand U23343 (N_23343,N_22562,N_22355);
nand U23344 (N_23344,N_22284,N_22481);
or U23345 (N_23345,N_22598,N_22453);
nand U23346 (N_23346,N_22624,N_22336);
and U23347 (N_23347,N_22407,N_22429);
or U23348 (N_23348,N_22267,N_22465);
or U23349 (N_23349,N_22377,N_22430);
or U23350 (N_23350,N_22621,N_22354);
xnor U23351 (N_23351,N_22426,N_22782);
nor U23352 (N_23352,N_22600,N_22424);
nand U23353 (N_23353,N_22790,N_22429);
nand U23354 (N_23354,N_22282,N_22559);
nor U23355 (N_23355,N_22782,N_22303);
or U23356 (N_23356,N_22599,N_22568);
and U23357 (N_23357,N_22399,N_22393);
and U23358 (N_23358,N_22742,N_22745);
or U23359 (N_23359,N_22292,N_22238);
nor U23360 (N_23360,N_22322,N_22372);
nor U23361 (N_23361,N_22432,N_22528);
nor U23362 (N_23362,N_22224,N_22711);
and U23363 (N_23363,N_22529,N_22452);
nand U23364 (N_23364,N_22773,N_22412);
nand U23365 (N_23365,N_22224,N_22730);
nand U23366 (N_23366,N_22553,N_22237);
nand U23367 (N_23367,N_22248,N_22417);
nor U23368 (N_23368,N_22548,N_22310);
or U23369 (N_23369,N_22617,N_22357);
and U23370 (N_23370,N_22200,N_22763);
nor U23371 (N_23371,N_22374,N_22591);
nand U23372 (N_23372,N_22355,N_22353);
or U23373 (N_23373,N_22455,N_22601);
nand U23374 (N_23374,N_22538,N_22524);
or U23375 (N_23375,N_22423,N_22774);
nor U23376 (N_23376,N_22460,N_22783);
nand U23377 (N_23377,N_22748,N_22772);
nor U23378 (N_23378,N_22750,N_22766);
and U23379 (N_23379,N_22666,N_22743);
and U23380 (N_23380,N_22705,N_22204);
or U23381 (N_23381,N_22701,N_22729);
nand U23382 (N_23382,N_22609,N_22375);
or U23383 (N_23383,N_22678,N_22590);
or U23384 (N_23384,N_22776,N_22328);
or U23385 (N_23385,N_22428,N_22460);
nor U23386 (N_23386,N_22398,N_22673);
or U23387 (N_23387,N_22675,N_22739);
xnor U23388 (N_23388,N_22257,N_22394);
and U23389 (N_23389,N_22529,N_22380);
or U23390 (N_23390,N_22571,N_22484);
xor U23391 (N_23391,N_22461,N_22531);
xor U23392 (N_23392,N_22229,N_22559);
or U23393 (N_23393,N_22536,N_22613);
or U23394 (N_23394,N_22662,N_22449);
nand U23395 (N_23395,N_22235,N_22518);
nand U23396 (N_23396,N_22697,N_22735);
nand U23397 (N_23397,N_22517,N_22495);
nand U23398 (N_23398,N_22460,N_22637);
xnor U23399 (N_23399,N_22615,N_22241);
xnor U23400 (N_23400,N_23368,N_23080);
nor U23401 (N_23401,N_23384,N_23030);
nor U23402 (N_23402,N_23092,N_22849);
nand U23403 (N_23403,N_22838,N_23215);
or U23404 (N_23404,N_23222,N_23023);
nor U23405 (N_23405,N_23225,N_23003);
nor U23406 (N_23406,N_23367,N_22935);
or U23407 (N_23407,N_23325,N_23362);
nand U23408 (N_23408,N_23358,N_22803);
and U23409 (N_23409,N_22978,N_22806);
nor U23410 (N_23410,N_23178,N_23143);
xnor U23411 (N_23411,N_22828,N_22931);
and U23412 (N_23412,N_22897,N_23000);
or U23413 (N_23413,N_22951,N_22873);
nor U23414 (N_23414,N_23087,N_22966);
nor U23415 (N_23415,N_23017,N_23145);
nor U23416 (N_23416,N_23345,N_22834);
nand U23417 (N_23417,N_23252,N_23088);
nor U23418 (N_23418,N_22864,N_23068);
nand U23419 (N_23419,N_23112,N_22800);
and U23420 (N_23420,N_22807,N_23175);
xnor U23421 (N_23421,N_23194,N_23011);
xnor U23422 (N_23422,N_23221,N_22816);
nor U23423 (N_23423,N_23301,N_22840);
nor U23424 (N_23424,N_23163,N_22945);
and U23425 (N_23425,N_23277,N_22982);
or U23426 (N_23426,N_22832,N_23341);
xnor U23427 (N_23427,N_23209,N_23138);
xnor U23428 (N_23428,N_23234,N_23122);
or U23429 (N_23429,N_22959,N_23352);
xnor U23430 (N_23430,N_23107,N_23149);
xnor U23431 (N_23431,N_23237,N_23328);
and U23432 (N_23432,N_22862,N_23361);
nor U23433 (N_23433,N_23395,N_23022);
nor U23434 (N_23434,N_23201,N_23116);
xor U23435 (N_23435,N_23075,N_22998);
or U23436 (N_23436,N_23266,N_23263);
nor U23437 (N_23437,N_23039,N_23074);
or U23438 (N_23438,N_23284,N_23398);
and U23439 (N_23439,N_23244,N_23396);
or U23440 (N_23440,N_23243,N_23162);
nor U23441 (N_23441,N_23025,N_23388);
nand U23442 (N_23442,N_23048,N_22955);
nor U23443 (N_23443,N_23264,N_23129);
nor U23444 (N_23444,N_23223,N_22843);
nand U23445 (N_23445,N_23317,N_23172);
nor U23446 (N_23446,N_23235,N_22989);
and U23447 (N_23447,N_23051,N_23012);
or U23448 (N_23448,N_23191,N_23248);
or U23449 (N_23449,N_23097,N_23110);
and U23450 (N_23450,N_23079,N_22993);
or U23451 (N_23451,N_23132,N_23106);
or U23452 (N_23452,N_23290,N_23306);
or U23453 (N_23453,N_23102,N_22990);
nor U23454 (N_23454,N_22995,N_22808);
nand U23455 (N_23455,N_22872,N_23044);
and U23456 (N_23456,N_23180,N_22884);
or U23457 (N_23457,N_23285,N_23016);
or U23458 (N_23458,N_23381,N_22914);
nand U23459 (N_23459,N_23089,N_23208);
nor U23460 (N_23460,N_23128,N_23391);
nand U23461 (N_23461,N_23257,N_23117);
and U23462 (N_23462,N_23064,N_22973);
xor U23463 (N_23463,N_22852,N_23049);
or U23464 (N_23464,N_23188,N_23307);
xnor U23465 (N_23465,N_22942,N_23108);
nor U23466 (N_23466,N_23158,N_23329);
nor U23467 (N_23467,N_22880,N_22819);
and U23468 (N_23468,N_23249,N_22985);
xor U23469 (N_23469,N_23333,N_23347);
xnor U23470 (N_23470,N_22888,N_22854);
or U23471 (N_23471,N_23004,N_23084);
and U23472 (N_23472,N_23386,N_23014);
xnor U23473 (N_23473,N_22837,N_23036);
nand U23474 (N_23474,N_23046,N_22920);
and U23475 (N_23475,N_23365,N_23183);
nor U23476 (N_23476,N_22824,N_23309);
xor U23477 (N_23477,N_23268,N_23137);
xor U23478 (N_23478,N_23115,N_22892);
and U23479 (N_23479,N_22981,N_22980);
nor U23480 (N_23480,N_23019,N_23148);
xnor U23481 (N_23481,N_23216,N_23171);
or U23482 (N_23482,N_22814,N_22830);
or U23483 (N_23483,N_22938,N_23065);
and U23484 (N_23484,N_23281,N_22836);
nand U23485 (N_23485,N_23118,N_23207);
nand U23486 (N_23486,N_23043,N_23189);
xor U23487 (N_23487,N_22963,N_23399);
nand U23488 (N_23488,N_23173,N_23002);
xnor U23489 (N_23489,N_23184,N_23392);
xnor U23490 (N_23490,N_22918,N_23071);
and U23491 (N_23491,N_23350,N_23348);
or U23492 (N_23492,N_22850,N_23247);
nand U23493 (N_23493,N_22833,N_23192);
nand U23494 (N_23494,N_23226,N_23010);
or U23495 (N_23495,N_22825,N_23327);
xnor U23496 (N_23496,N_22970,N_22802);
and U23497 (N_23497,N_22908,N_23008);
nor U23498 (N_23498,N_23385,N_22911);
xor U23499 (N_23499,N_23300,N_22969);
and U23500 (N_23500,N_22889,N_22986);
nor U23501 (N_23501,N_23276,N_22905);
nand U23502 (N_23502,N_23369,N_22956);
nand U23503 (N_23503,N_23136,N_23186);
nor U23504 (N_23504,N_22907,N_23182);
nor U23505 (N_23505,N_23139,N_23273);
and U23506 (N_23506,N_23187,N_23330);
and U23507 (N_23507,N_23370,N_23177);
and U23508 (N_23508,N_23259,N_22804);
xor U23509 (N_23509,N_23037,N_23041);
xor U23510 (N_23510,N_22826,N_23357);
and U23511 (N_23511,N_22853,N_23072);
or U23512 (N_23512,N_23166,N_23360);
or U23513 (N_23513,N_23363,N_22976);
xor U23514 (N_23514,N_22876,N_23331);
nand U23515 (N_23515,N_22952,N_23093);
or U23516 (N_23516,N_23305,N_22874);
and U23517 (N_23517,N_23035,N_22894);
xor U23518 (N_23518,N_23340,N_23343);
nor U23519 (N_23519,N_22867,N_23220);
and U23520 (N_23520,N_23297,N_23389);
nand U23521 (N_23521,N_23121,N_23200);
nand U23522 (N_23522,N_22813,N_23324);
nor U23523 (N_23523,N_23038,N_23314);
xnor U23524 (N_23524,N_22967,N_22823);
nand U23525 (N_23525,N_22860,N_23058);
or U23526 (N_23526,N_22987,N_22858);
or U23527 (N_23527,N_23001,N_23313);
xnor U23528 (N_23528,N_22988,N_22968);
xnor U23529 (N_23529,N_22939,N_23167);
or U23530 (N_23530,N_22922,N_23150);
and U23531 (N_23531,N_22857,N_22801);
nand U23532 (N_23532,N_23203,N_22847);
and U23533 (N_23533,N_23344,N_22941);
nand U23534 (N_23534,N_23308,N_23125);
xnor U23535 (N_23535,N_22805,N_22870);
nor U23536 (N_23536,N_23169,N_23380);
or U23537 (N_23537,N_23170,N_23359);
nand U23538 (N_23538,N_23081,N_23262);
or U23539 (N_23539,N_22861,N_23293);
and U23540 (N_23540,N_22891,N_23119);
nor U23541 (N_23541,N_23230,N_22902);
nor U23542 (N_23542,N_23042,N_23337);
nor U23543 (N_23543,N_23390,N_22954);
and U23544 (N_23544,N_23312,N_23278);
nand U23545 (N_23545,N_23111,N_23311);
nand U23546 (N_23546,N_23303,N_23077);
nor U23547 (N_23547,N_22940,N_23056);
or U23548 (N_23548,N_23383,N_23214);
or U23549 (N_23549,N_23349,N_22821);
and U23550 (N_23550,N_22979,N_23224);
and U23551 (N_23551,N_22877,N_23168);
or U23552 (N_23552,N_23336,N_23031);
nor U23553 (N_23553,N_22900,N_23013);
or U23554 (N_23554,N_22996,N_23355);
and U23555 (N_23555,N_22879,N_23227);
nor U23556 (N_23556,N_23164,N_23316);
or U23557 (N_23557,N_22999,N_23176);
nand U23558 (N_23558,N_22923,N_23083);
xnor U23559 (N_23559,N_23069,N_23378);
and U23560 (N_23560,N_22831,N_23135);
or U23561 (N_23561,N_22871,N_23040);
xnor U23562 (N_23562,N_23134,N_22896);
nor U23563 (N_23563,N_23339,N_22881);
nor U23564 (N_23564,N_23090,N_23335);
nor U23565 (N_23565,N_23261,N_22972);
xor U23566 (N_23566,N_23377,N_22977);
xor U23567 (N_23567,N_22904,N_23179);
nor U23568 (N_23568,N_22953,N_23205);
xnor U23569 (N_23569,N_22878,N_23321);
xnor U23570 (N_23570,N_23258,N_22997);
and U23571 (N_23571,N_23238,N_23326);
nand U23572 (N_23572,N_23219,N_23236);
and U23573 (N_23573,N_23159,N_22851);
and U23574 (N_23574,N_23241,N_22839);
nor U23575 (N_23575,N_23332,N_23060);
or U23576 (N_23576,N_23130,N_23157);
xor U23577 (N_23577,N_22958,N_22820);
and U23578 (N_23578,N_23098,N_23232);
or U23579 (N_23579,N_23212,N_22925);
nor U23580 (N_23580,N_22994,N_23152);
nand U23581 (N_23581,N_23260,N_23161);
xor U23582 (N_23582,N_23015,N_23033);
nand U23583 (N_23583,N_22949,N_23275);
nor U23584 (N_23584,N_22912,N_23382);
nand U23585 (N_23585,N_22974,N_23020);
nor U23586 (N_23586,N_22926,N_23354);
nand U23587 (N_23587,N_22946,N_23005);
and U23588 (N_23588,N_22811,N_22898);
nor U23589 (N_23589,N_23196,N_22865);
nand U23590 (N_23590,N_22818,N_23288);
and U23591 (N_23591,N_23376,N_23298);
nor U23592 (N_23592,N_23142,N_22829);
xnor U23593 (N_23593,N_23120,N_23299);
xor U23594 (N_23594,N_23185,N_23063);
nor U23595 (N_23595,N_23140,N_22937);
or U23596 (N_23596,N_22885,N_23151);
nand U23597 (N_23597,N_22913,N_22863);
and U23598 (N_23598,N_23195,N_23006);
nand U23599 (N_23599,N_23109,N_23029);
xor U23600 (N_23600,N_23197,N_23296);
xor U23601 (N_23601,N_23127,N_23211);
xnor U23602 (N_23602,N_22866,N_22915);
xnor U23603 (N_23603,N_23342,N_23034);
xor U23604 (N_23604,N_23302,N_23206);
or U23605 (N_23605,N_23146,N_22842);
or U23606 (N_23606,N_23156,N_23123);
nor U23607 (N_23607,N_22948,N_22932);
and U23608 (N_23608,N_23141,N_23315);
or U23609 (N_23609,N_23070,N_23032);
or U23610 (N_23610,N_23114,N_23052);
nand U23611 (N_23611,N_23155,N_23217);
nor U23612 (N_23612,N_22975,N_23371);
nor U23613 (N_23613,N_22883,N_22859);
nor U23614 (N_23614,N_23274,N_23181);
xnor U23615 (N_23615,N_23021,N_23291);
nand U23616 (N_23616,N_23364,N_23295);
xor U23617 (N_23617,N_23334,N_23242);
and U23618 (N_23618,N_22835,N_23283);
or U23619 (N_23619,N_22895,N_23346);
or U23620 (N_23620,N_22927,N_23353);
nor U23621 (N_23621,N_22848,N_23253);
nor U23622 (N_23622,N_23066,N_22930);
or U23623 (N_23623,N_23320,N_22890);
or U23624 (N_23624,N_23190,N_23292);
xnor U23625 (N_23625,N_23096,N_23373);
nand U23626 (N_23626,N_23280,N_22809);
nand U23627 (N_23627,N_22950,N_22844);
nor U23628 (N_23628,N_23104,N_23387);
and U23629 (N_23629,N_23054,N_23279);
nand U23630 (N_23630,N_23265,N_23199);
or U23631 (N_23631,N_22841,N_22812);
or U23632 (N_23632,N_22964,N_23269);
xor U23633 (N_23633,N_23085,N_23310);
and U23634 (N_23634,N_23153,N_22919);
nand U23635 (N_23635,N_23160,N_23374);
and U23636 (N_23636,N_23076,N_22921);
and U23637 (N_23637,N_23318,N_23202);
nand U23638 (N_23638,N_23282,N_22992);
nand U23639 (N_23639,N_23009,N_23147);
nor U23640 (N_23640,N_22899,N_22845);
and U23641 (N_23641,N_22936,N_23086);
nand U23642 (N_23642,N_23289,N_23270);
nor U23643 (N_23643,N_23271,N_22947);
xor U23644 (N_23644,N_23272,N_23256);
or U23645 (N_23645,N_23061,N_22901);
xor U23646 (N_23646,N_23053,N_23250);
nand U23647 (N_23647,N_23067,N_22924);
xor U23648 (N_23648,N_23251,N_23091);
nor U23649 (N_23649,N_22943,N_23287);
nor U23650 (N_23650,N_22909,N_22971);
xnor U23651 (N_23651,N_22984,N_23028);
nand U23652 (N_23652,N_23113,N_23245);
nor U23653 (N_23653,N_23133,N_23027);
and U23654 (N_23654,N_23233,N_22810);
nor U23655 (N_23655,N_23026,N_23229);
and U23656 (N_23656,N_23240,N_23131);
nand U23657 (N_23657,N_23319,N_22934);
and U23658 (N_23658,N_23228,N_22957);
nand U23659 (N_23659,N_23231,N_22893);
nand U23660 (N_23660,N_23045,N_23322);
nand U23661 (N_23661,N_23239,N_23126);
nor U23662 (N_23662,N_23394,N_23255);
xnor U23663 (N_23663,N_23294,N_22933);
or U23664 (N_23664,N_22815,N_23267);
and U23665 (N_23665,N_22827,N_23254);
or U23666 (N_23666,N_23210,N_23204);
and U23667 (N_23667,N_22855,N_22875);
and U23668 (N_23668,N_22917,N_23198);
or U23669 (N_23669,N_23379,N_22991);
and U23670 (N_23670,N_22869,N_23073);
nor U23671 (N_23671,N_23101,N_22868);
nand U23672 (N_23672,N_23007,N_23304);
xor U23673 (N_23673,N_22887,N_22929);
nand U23674 (N_23674,N_23078,N_23372);
nand U23675 (N_23675,N_23338,N_23105);
nor U23676 (N_23676,N_23059,N_23154);
nand U23677 (N_23677,N_23094,N_23351);
nor U23678 (N_23678,N_23024,N_22916);
nand U23679 (N_23679,N_23144,N_22817);
nand U23680 (N_23680,N_23082,N_23050);
and U23681 (N_23681,N_23100,N_23397);
nand U23682 (N_23682,N_22906,N_22846);
nor U23683 (N_23683,N_23356,N_22856);
nand U23684 (N_23684,N_23286,N_22910);
nor U23685 (N_23685,N_23062,N_22882);
nand U23686 (N_23686,N_23366,N_22965);
nor U23687 (N_23687,N_23099,N_23103);
and U23688 (N_23688,N_23124,N_22983);
and U23689 (N_23689,N_23174,N_22928);
nor U23690 (N_23690,N_23055,N_23393);
xor U23691 (N_23691,N_22822,N_22944);
nand U23692 (N_23692,N_22962,N_23375);
and U23693 (N_23693,N_23218,N_23057);
and U23694 (N_23694,N_22903,N_23095);
nand U23695 (N_23695,N_23323,N_23213);
and U23696 (N_23696,N_23165,N_23018);
nand U23697 (N_23697,N_22960,N_23047);
xnor U23698 (N_23698,N_23193,N_23246);
and U23699 (N_23699,N_22886,N_22961);
nor U23700 (N_23700,N_22897,N_23240);
nand U23701 (N_23701,N_23372,N_22940);
and U23702 (N_23702,N_23330,N_23116);
and U23703 (N_23703,N_23359,N_23391);
nand U23704 (N_23704,N_23163,N_22819);
nand U23705 (N_23705,N_22884,N_23365);
nand U23706 (N_23706,N_22934,N_23086);
xnor U23707 (N_23707,N_22826,N_22932);
and U23708 (N_23708,N_23184,N_23356);
nor U23709 (N_23709,N_22816,N_23287);
xnor U23710 (N_23710,N_23051,N_22946);
or U23711 (N_23711,N_22837,N_22992);
or U23712 (N_23712,N_22811,N_22871);
or U23713 (N_23713,N_22996,N_23304);
or U23714 (N_23714,N_23020,N_22816);
xnor U23715 (N_23715,N_23107,N_23221);
nor U23716 (N_23716,N_22909,N_23264);
or U23717 (N_23717,N_23106,N_23350);
nor U23718 (N_23718,N_23240,N_23301);
nand U23719 (N_23719,N_22957,N_23385);
xnor U23720 (N_23720,N_22944,N_23270);
nand U23721 (N_23721,N_23362,N_23123);
nand U23722 (N_23722,N_23000,N_22879);
nor U23723 (N_23723,N_23221,N_23391);
xnor U23724 (N_23724,N_23047,N_22949);
nor U23725 (N_23725,N_23299,N_23098);
xnor U23726 (N_23726,N_23184,N_22885);
nor U23727 (N_23727,N_22940,N_22971);
nand U23728 (N_23728,N_23328,N_23107);
xnor U23729 (N_23729,N_23021,N_23267);
nor U23730 (N_23730,N_23171,N_23047);
nor U23731 (N_23731,N_22950,N_22831);
nand U23732 (N_23732,N_23204,N_23326);
or U23733 (N_23733,N_23295,N_23158);
xnor U23734 (N_23734,N_22939,N_23262);
xnor U23735 (N_23735,N_23129,N_22869);
nand U23736 (N_23736,N_22887,N_22930);
nand U23737 (N_23737,N_23062,N_23308);
nor U23738 (N_23738,N_23194,N_23224);
and U23739 (N_23739,N_23123,N_22927);
nor U23740 (N_23740,N_22951,N_22882);
nand U23741 (N_23741,N_23354,N_23211);
nand U23742 (N_23742,N_23007,N_22866);
and U23743 (N_23743,N_23320,N_22861);
xnor U23744 (N_23744,N_23071,N_23159);
or U23745 (N_23745,N_23035,N_23270);
nand U23746 (N_23746,N_23064,N_23030);
xnor U23747 (N_23747,N_22819,N_22805);
and U23748 (N_23748,N_22821,N_23282);
and U23749 (N_23749,N_23095,N_23039);
nand U23750 (N_23750,N_22831,N_23072);
or U23751 (N_23751,N_23397,N_22948);
nand U23752 (N_23752,N_23340,N_22865);
nand U23753 (N_23753,N_23014,N_23284);
and U23754 (N_23754,N_22964,N_23060);
or U23755 (N_23755,N_22884,N_23106);
xnor U23756 (N_23756,N_22908,N_22816);
or U23757 (N_23757,N_23075,N_22953);
nor U23758 (N_23758,N_23145,N_23371);
xnor U23759 (N_23759,N_23371,N_23235);
or U23760 (N_23760,N_23147,N_23356);
or U23761 (N_23761,N_22912,N_23354);
and U23762 (N_23762,N_23234,N_23317);
and U23763 (N_23763,N_23031,N_23352);
nor U23764 (N_23764,N_23228,N_23385);
nor U23765 (N_23765,N_23321,N_23133);
xnor U23766 (N_23766,N_23172,N_22829);
and U23767 (N_23767,N_23273,N_23003);
and U23768 (N_23768,N_23082,N_23255);
or U23769 (N_23769,N_23190,N_23303);
nor U23770 (N_23770,N_23347,N_23042);
or U23771 (N_23771,N_22904,N_22924);
xor U23772 (N_23772,N_23379,N_22849);
or U23773 (N_23773,N_22878,N_22881);
and U23774 (N_23774,N_23105,N_23317);
nor U23775 (N_23775,N_23367,N_23254);
nand U23776 (N_23776,N_23137,N_23193);
or U23777 (N_23777,N_23393,N_22973);
xnor U23778 (N_23778,N_23359,N_23384);
nand U23779 (N_23779,N_22893,N_23016);
xnor U23780 (N_23780,N_22897,N_23107);
xor U23781 (N_23781,N_23008,N_23313);
and U23782 (N_23782,N_23264,N_23340);
xnor U23783 (N_23783,N_23057,N_22875);
or U23784 (N_23784,N_23250,N_23340);
xor U23785 (N_23785,N_23102,N_23235);
xnor U23786 (N_23786,N_23080,N_23254);
or U23787 (N_23787,N_23071,N_23358);
or U23788 (N_23788,N_22932,N_22911);
nand U23789 (N_23789,N_23056,N_23284);
nor U23790 (N_23790,N_23121,N_23217);
nor U23791 (N_23791,N_23066,N_23189);
nand U23792 (N_23792,N_22986,N_22974);
xnor U23793 (N_23793,N_23373,N_22896);
nand U23794 (N_23794,N_23028,N_22911);
nand U23795 (N_23795,N_23070,N_23239);
nor U23796 (N_23796,N_22855,N_23363);
nand U23797 (N_23797,N_23263,N_23143);
and U23798 (N_23798,N_23207,N_22893);
or U23799 (N_23799,N_23325,N_23029);
nor U23800 (N_23800,N_23389,N_23260);
or U23801 (N_23801,N_22985,N_22847);
xor U23802 (N_23802,N_23375,N_23067);
or U23803 (N_23803,N_23361,N_23159);
nor U23804 (N_23804,N_22970,N_23328);
nand U23805 (N_23805,N_23396,N_23389);
or U23806 (N_23806,N_22965,N_22813);
and U23807 (N_23807,N_23335,N_23110);
xor U23808 (N_23808,N_23177,N_23315);
nor U23809 (N_23809,N_22851,N_22900);
or U23810 (N_23810,N_23027,N_22853);
nor U23811 (N_23811,N_23085,N_23386);
nand U23812 (N_23812,N_23310,N_23097);
or U23813 (N_23813,N_23290,N_22917);
nor U23814 (N_23814,N_22985,N_23160);
and U23815 (N_23815,N_22832,N_23363);
xor U23816 (N_23816,N_23040,N_23209);
nor U23817 (N_23817,N_23102,N_23162);
xnor U23818 (N_23818,N_22931,N_22925);
nand U23819 (N_23819,N_23168,N_23089);
or U23820 (N_23820,N_23348,N_23329);
nor U23821 (N_23821,N_22845,N_23206);
and U23822 (N_23822,N_22921,N_22907);
nand U23823 (N_23823,N_22900,N_22973);
xnor U23824 (N_23824,N_23309,N_23363);
and U23825 (N_23825,N_23055,N_23228);
nand U23826 (N_23826,N_23301,N_23105);
or U23827 (N_23827,N_22993,N_22989);
nor U23828 (N_23828,N_23247,N_23136);
and U23829 (N_23829,N_23259,N_23385);
xor U23830 (N_23830,N_23324,N_22926);
xor U23831 (N_23831,N_23091,N_23263);
or U23832 (N_23832,N_22916,N_23088);
nor U23833 (N_23833,N_23228,N_23356);
nor U23834 (N_23834,N_23171,N_23065);
xnor U23835 (N_23835,N_23173,N_23025);
or U23836 (N_23836,N_23346,N_22958);
nor U23837 (N_23837,N_23048,N_23327);
xnor U23838 (N_23838,N_23388,N_22868);
or U23839 (N_23839,N_23287,N_22904);
nand U23840 (N_23840,N_23107,N_23374);
xnor U23841 (N_23841,N_23238,N_22886);
xor U23842 (N_23842,N_23385,N_22935);
xnor U23843 (N_23843,N_23140,N_23097);
and U23844 (N_23844,N_23081,N_23203);
nor U23845 (N_23845,N_22818,N_23389);
xnor U23846 (N_23846,N_23398,N_23168);
and U23847 (N_23847,N_23324,N_22885);
and U23848 (N_23848,N_23018,N_22857);
nand U23849 (N_23849,N_23141,N_22948);
nand U23850 (N_23850,N_22865,N_23031);
xor U23851 (N_23851,N_23092,N_23358);
nand U23852 (N_23852,N_23390,N_23243);
xor U23853 (N_23853,N_22909,N_23262);
nor U23854 (N_23854,N_23211,N_22940);
nand U23855 (N_23855,N_23053,N_23226);
xnor U23856 (N_23856,N_23039,N_22985);
and U23857 (N_23857,N_23319,N_22902);
or U23858 (N_23858,N_23028,N_22858);
nor U23859 (N_23859,N_22845,N_23334);
or U23860 (N_23860,N_22836,N_23197);
nand U23861 (N_23861,N_23024,N_23265);
xnor U23862 (N_23862,N_23042,N_22962);
xor U23863 (N_23863,N_23129,N_23254);
nor U23864 (N_23864,N_23271,N_22935);
or U23865 (N_23865,N_23202,N_23003);
nor U23866 (N_23866,N_22817,N_23021);
and U23867 (N_23867,N_23232,N_23190);
nor U23868 (N_23868,N_23121,N_22901);
or U23869 (N_23869,N_23239,N_22890);
nor U23870 (N_23870,N_22984,N_23177);
xnor U23871 (N_23871,N_23136,N_23331);
xnor U23872 (N_23872,N_23364,N_23244);
xnor U23873 (N_23873,N_22852,N_23107);
and U23874 (N_23874,N_23255,N_23104);
and U23875 (N_23875,N_22813,N_23292);
nand U23876 (N_23876,N_23206,N_23040);
and U23877 (N_23877,N_23237,N_23042);
nand U23878 (N_23878,N_22826,N_23371);
xnor U23879 (N_23879,N_22808,N_22812);
xor U23880 (N_23880,N_23044,N_23315);
or U23881 (N_23881,N_23250,N_23338);
xnor U23882 (N_23882,N_23079,N_23255);
nor U23883 (N_23883,N_23234,N_23178);
or U23884 (N_23884,N_23364,N_23236);
xnor U23885 (N_23885,N_23182,N_23161);
and U23886 (N_23886,N_23004,N_23313);
or U23887 (N_23887,N_23330,N_22910);
or U23888 (N_23888,N_23387,N_23235);
or U23889 (N_23889,N_23217,N_23115);
nor U23890 (N_23890,N_23138,N_22983);
xnor U23891 (N_23891,N_22958,N_22950);
or U23892 (N_23892,N_22930,N_23304);
nand U23893 (N_23893,N_22809,N_23208);
nor U23894 (N_23894,N_23078,N_23346);
nand U23895 (N_23895,N_22925,N_23023);
nor U23896 (N_23896,N_22936,N_23204);
nand U23897 (N_23897,N_23194,N_23239);
or U23898 (N_23898,N_23219,N_22843);
xnor U23899 (N_23899,N_23316,N_22977);
nor U23900 (N_23900,N_23064,N_22838);
or U23901 (N_23901,N_22924,N_22930);
xnor U23902 (N_23902,N_23371,N_23378);
and U23903 (N_23903,N_23352,N_23088);
nand U23904 (N_23904,N_22831,N_23079);
and U23905 (N_23905,N_23050,N_22926);
nor U23906 (N_23906,N_23110,N_23158);
or U23907 (N_23907,N_22846,N_23130);
xnor U23908 (N_23908,N_22992,N_23141);
nand U23909 (N_23909,N_23360,N_22822);
nor U23910 (N_23910,N_22843,N_23040);
nand U23911 (N_23911,N_22928,N_22901);
nor U23912 (N_23912,N_22873,N_23065);
and U23913 (N_23913,N_23212,N_22920);
nor U23914 (N_23914,N_23372,N_23028);
or U23915 (N_23915,N_23114,N_23337);
and U23916 (N_23916,N_23256,N_22861);
nand U23917 (N_23917,N_22806,N_23175);
and U23918 (N_23918,N_23103,N_22919);
and U23919 (N_23919,N_23208,N_22882);
or U23920 (N_23920,N_23337,N_23382);
nand U23921 (N_23921,N_22987,N_23192);
xnor U23922 (N_23922,N_22830,N_23215);
and U23923 (N_23923,N_23105,N_22933);
nor U23924 (N_23924,N_22931,N_23307);
and U23925 (N_23925,N_22887,N_23080);
or U23926 (N_23926,N_23092,N_23343);
xnor U23927 (N_23927,N_22896,N_22876);
xnor U23928 (N_23928,N_23005,N_22895);
nor U23929 (N_23929,N_23105,N_22818);
nor U23930 (N_23930,N_23079,N_23184);
xor U23931 (N_23931,N_22904,N_23021);
and U23932 (N_23932,N_23170,N_23182);
and U23933 (N_23933,N_22948,N_23061);
and U23934 (N_23934,N_23025,N_22890);
xnor U23935 (N_23935,N_23250,N_23163);
nor U23936 (N_23936,N_22964,N_23164);
or U23937 (N_23937,N_23335,N_23316);
nand U23938 (N_23938,N_23035,N_23026);
xnor U23939 (N_23939,N_23150,N_22972);
nor U23940 (N_23940,N_23316,N_22838);
or U23941 (N_23941,N_23353,N_22907);
nand U23942 (N_23942,N_22851,N_22818);
nor U23943 (N_23943,N_23240,N_23030);
and U23944 (N_23944,N_23377,N_22837);
nand U23945 (N_23945,N_22931,N_23296);
xnor U23946 (N_23946,N_23314,N_22984);
xor U23947 (N_23947,N_23132,N_22979);
or U23948 (N_23948,N_22957,N_23312);
or U23949 (N_23949,N_22822,N_23191);
or U23950 (N_23950,N_23285,N_23346);
or U23951 (N_23951,N_23202,N_23263);
nand U23952 (N_23952,N_23075,N_22900);
nand U23953 (N_23953,N_23101,N_23123);
nand U23954 (N_23954,N_23251,N_22867);
nor U23955 (N_23955,N_23344,N_23343);
and U23956 (N_23956,N_22980,N_22927);
nor U23957 (N_23957,N_23238,N_23209);
or U23958 (N_23958,N_23325,N_22842);
nand U23959 (N_23959,N_23101,N_22802);
xor U23960 (N_23960,N_22931,N_23084);
nand U23961 (N_23961,N_22808,N_23088);
nor U23962 (N_23962,N_22844,N_22816);
or U23963 (N_23963,N_23182,N_23048);
or U23964 (N_23964,N_23095,N_23041);
and U23965 (N_23965,N_23013,N_23270);
or U23966 (N_23966,N_22857,N_23285);
nor U23967 (N_23967,N_22987,N_23076);
xor U23968 (N_23968,N_23055,N_23158);
xor U23969 (N_23969,N_23118,N_22944);
or U23970 (N_23970,N_22999,N_22982);
nor U23971 (N_23971,N_23370,N_23097);
nor U23972 (N_23972,N_22881,N_22880);
nor U23973 (N_23973,N_22802,N_23289);
xor U23974 (N_23974,N_23370,N_23379);
nand U23975 (N_23975,N_23094,N_23241);
or U23976 (N_23976,N_23123,N_23303);
nor U23977 (N_23977,N_23216,N_23102);
and U23978 (N_23978,N_23079,N_23273);
or U23979 (N_23979,N_23301,N_22837);
nand U23980 (N_23980,N_22959,N_23275);
nor U23981 (N_23981,N_22995,N_23190);
nor U23982 (N_23982,N_23290,N_22863);
nor U23983 (N_23983,N_23090,N_22955);
xor U23984 (N_23984,N_22918,N_22841);
nor U23985 (N_23985,N_23360,N_23020);
and U23986 (N_23986,N_22999,N_22821);
and U23987 (N_23987,N_23066,N_23240);
and U23988 (N_23988,N_22821,N_23037);
nor U23989 (N_23989,N_23037,N_23078);
nor U23990 (N_23990,N_23119,N_23112);
nand U23991 (N_23991,N_22945,N_23008);
nor U23992 (N_23992,N_23398,N_22945);
xor U23993 (N_23993,N_23352,N_23034);
nand U23994 (N_23994,N_23194,N_22807);
nor U23995 (N_23995,N_23335,N_23338);
nand U23996 (N_23996,N_23179,N_23322);
xnor U23997 (N_23997,N_23026,N_23361);
nand U23998 (N_23998,N_23192,N_23264);
xnor U23999 (N_23999,N_23141,N_22994);
nor U24000 (N_24000,N_23645,N_23677);
nor U24001 (N_24001,N_23570,N_23464);
xor U24002 (N_24002,N_23528,N_23632);
and U24003 (N_24003,N_23861,N_23634);
nand U24004 (N_24004,N_23899,N_23990);
xnor U24005 (N_24005,N_23991,N_23710);
xor U24006 (N_24006,N_23611,N_23964);
xnor U24007 (N_24007,N_23689,N_23944);
nand U24008 (N_24008,N_23694,N_23993);
nand U24009 (N_24009,N_23994,N_23806);
and U24010 (N_24010,N_23875,N_23532);
nand U24011 (N_24011,N_23736,N_23636);
and U24012 (N_24012,N_23697,N_23984);
or U24013 (N_24013,N_23921,N_23562);
xor U24014 (N_24014,N_23959,N_23950);
nor U24015 (N_24015,N_23801,N_23661);
and U24016 (N_24016,N_23704,N_23855);
xor U24017 (N_24017,N_23913,N_23617);
or U24018 (N_24018,N_23483,N_23792);
or U24019 (N_24019,N_23401,N_23529);
or U24020 (N_24020,N_23598,N_23545);
or U24021 (N_24021,N_23893,N_23638);
or U24022 (N_24022,N_23523,N_23682);
xor U24023 (N_24023,N_23556,N_23916);
nor U24024 (N_24024,N_23750,N_23582);
xor U24025 (N_24025,N_23847,N_23476);
nor U24026 (N_24026,N_23663,N_23621);
and U24027 (N_24027,N_23650,N_23633);
nor U24028 (N_24028,N_23918,N_23961);
or U24029 (N_24029,N_23488,N_23563);
nand U24030 (N_24030,N_23826,N_23596);
or U24031 (N_24031,N_23492,N_23434);
nor U24032 (N_24032,N_23500,N_23683);
nand U24033 (N_24033,N_23724,N_23738);
xor U24034 (N_24034,N_23837,N_23760);
nand U24035 (N_24035,N_23431,N_23456);
xnor U24036 (N_24036,N_23997,N_23443);
or U24037 (N_24037,N_23930,N_23781);
nor U24038 (N_24038,N_23654,N_23752);
and U24039 (N_24039,N_23606,N_23735);
nor U24040 (N_24040,N_23739,N_23519);
or U24041 (N_24041,N_23776,N_23771);
xnor U24042 (N_24042,N_23762,N_23437);
and U24043 (N_24043,N_23469,N_23446);
or U24044 (N_24044,N_23815,N_23924);
xor U24045 (N_24045,N_23473,N_23883);
or U24046 (N_24046,N_23936,N_23414);
nor U24047 (N_24047,N_23722,N_23402);
xnor U24048 (N_24048,N_23573,N_23881);
or U24049 (N_24049,N_23513,N_23729);
xor U24050 (N_24050,N_23419,N_23898);
nor U24051 (N_24051,N_23868,N_23769);
nand U24052 (N_24052,N_23974,N_23856);
xor U24053 (N_24053,N_23681,N_23400);
and U24054 (N_24054,N_23442,N_23809);
nand U24055 (N_24055,N_23779,N_23509);
xor U24056 (N_24056,N_23471,N_23770);
and U24057 (N_24057,N_23583,N_23745);
and U24058 (N_24058,N_23879,N_23934);
and U24059 (N_24059,N_23648,N_23825);
nor U24060 (N_24060,N_23901,N_23538);
xor U24061 (N_24061,N_23678,N_23450);
nand U24062 (N_24062,N_23499,N_23592);
and U24063 (N_24063,N_23628,N_23639);
nor U24064 (N_24064,N_23876,N_23914);
nor U24065 (N_24065,N_23740,N_23518);
or U24066 (N_24066,N_23448,N_23629);
and U24067 (N_24067,N_23413,N_23841);
or U24068 (N_24068,N_23664,N_23882);
nand U24069 (N_24069,N_23641,N_23527);
nand U24070 (N_24070,N_23466,N_23965);
or U24071 (N_24071,N_23960,N_23676);
and U24072 (N_24072,N_23671,N_23428);
xor U24073 (N_24073,N_23708,N_23884);
nand U24074 (N_24074,N_23426,N_23851);
nor U24075 (N_24075,N_23758,N_23498);
nand U24076 (N_24076,N_23418,N_23834);
and U24077 (N_24077,N_23853,N_23701);
nor U24078 (N_24078,N_23968,N_23477);
and U24079 (N_24079,N_23858,N_23764);
xor U24080 (N_24080,N_23668,N_23586);
or U24081 (N_24081,N_23813,N_23590);
xor U24082 (N_24082,N_23917,N_23656);
or U24083 (N_24083,N_23608,N_23555);
and U24084 (N_24084,N_23880,N_23695);
nand U24085 (N_24085,N_23441,N_23995);
nor U24086 (N_24086,N_23604,N_23470);
xnor U24087 (N_24087,N_23415,N_23662);
and U24088 (N_24088,N_23620,N_23566);
and U24089 (N_24089,N_23747,N_23686);
nor U24090 (N_24090,N_23975,N_23808);
xor U24091 (N_24091,N_23790,N_23980);
xor U24092 (N_24092,N_23978,N_23507);
nor U24093 (N_24093,N_23521,N_23933);
nand U24094 (N_24094,N_23553,N_23833);
and U24095 (N_24095,N_23940,N_23484);
and U24096 (N_24096,N_23605,N_23755);
nand U24097 (N_24097,N_23811,N_23560);
and U24098 (N_24098,N_23603,N_23494);
and U24099 (N_24099,N_23593,N_23669);
nand U24100 (N_24100,N_23478,N_23777);
or U24101 (N_24101,N_23999,N_23992);
nor U24102 (N_24102,N_23907,N_23873);
nor U24103 (N_24103,N_23547,N_23440);
xor U24104 (N_24104,N_23807,N_23599);
xor U24105 (N_24105,N_23627,N_23712);
nand U24106 (N_24106,N_23859,N_23463);
xnor U24107 (N_24107,N_23939,N_23888);
nand U24108 (N_24108,N_23646,N_23761);
xnor U24109 (N_24109,N_23577,N_23778);
and U24110 (N_24110,N_23820,N_23430);
nor U24111 (N_24111,N_23886,N_23536);
and U24112 (N_24112,N_23989,N_23839);
xnor U24113 (N_24113,N_23460,N_23969);
nor U24114 (N_24114,N_23404,N_23998);
nor U24115 (N_24115,N_23465,N_23832);
nor U24116 (N_24116,N_23958,N_23455);
or U24117 (N_24117,N_23673,N_23626);
or U24118 (N_24118,N_23895,N_23850);
and U24119 (N_24119,N_23848,N_23584);
and U24120 (N_24120,N_23571,N_23516);
and U24121 (N_24121,N_23459,N_23725);
and U24122 (N_24122,N_23951,N_23515);
xor U24123 (N_24123,N_23892,N_23702);
nor U24124 (N_24124,N_23618,N_23726);
and U24125 (N_24125,N_23927,N_23533);
nand U24126 (N_24126,N_23672,N_23572);
nand U24127 (N_24127,N_23458,N_23727);
nand U24128 (N_24128,N_23407,N_23754);
nand U24129 (N_24129,N_23445,N_23630);
nand U24130 (N_24130,N_23835,N_23530);
or U24131 (N_24131,N_23496,N_23731);
nor U24132 (N_24132,N_23773,N_23782);
nand U24133 (N_24133,N_23922,N_23955);
nor U24134 (N_24134,N_23580,N_23869);
nand U24135 (N_24135,N_23561,N_23453);
nand U24136 (N_24136,N_23526,N_23952);
nor U24137 (N_24137,N_23728,N_23768);
and U24138 (N_24138,N_23763,N_23957);
or U24139 (N_24139,N_23438,N_23432);
nand U24140 (N_24140,N_23552,N_23569);
and U24141 (N_24141,N_23447,N_23878);
nor U24142 (N_24142,N_23711,N_23775);
or U24143 (N_24143,N_23439,N_23693);
xnor U24144 (N_24144,N_23667,N_23684);
nor U24145 (N_24145,N_23581,N_23915);
xor U24146 (N_24146,N_23549,N_23436);
xnor U24147 (N_24147,N_23709,N_23979);
or U24148 (N_24148,N_23690,N_23597);
nand U24149 (N_24149,N_23900,N_23749);
or U24150 (N_24150,N_23746,N_23482);
and U24151 (N_24151,N_23405,N_23877);
and U24152 (N_24152,N_23817,N_23904);
xnor U24153 (N_24153,N_23688,N_23600);
or U24154 (N_24154,N_23798,N_23416);
and U24155 (N_24155,N_23522,N_23602);
nor U24156 (N_24156,N_23786,N_23919);
xnor U24157 (N_24157,N_23417,N_23559);
nand U24158 (N_24158,N_23823,N_23720);
xor U24159 (N_24159,N_23637,N_23505);
nand U24160 (N_24160,N_23653,N_23824);
xor U24161 (N_24161,N_23793,N_23557);
or U24162 (N_24162,N_23860,N_23640);
and U24163 (N_24163,N_23647,N_23759);
and U24164 (N_24164,N_23624,N_23977);
nand U24165 (N_24165,N_23472,N_23838);
and U24166 (N_24166,N_23737,N_23887);
nand U24167 (N_24167,N_23967,N_23796);
nand U24168 (N_24168,N_23550,N_23982);
xnor U24169 (N_24169,N_23732,N_23475);
nor U24170 (N_24170,N_23774,N_23435);
xor U24171 (N_24171,N_23829,N_23937);
or U24172 (N_24172,N_23468,N_23985);
or U24173 (N_24173,N_23408,N_23819);
or U24174 (N_24174,N_23751,N_23451);
and U24175 (N_24175,N_23912,N_23902);
and U24176 (N_24176,N_23942,N_23954);
nor U24177 (N_24177,N_23714,N_23539);
and U24178 (N_24178,N_23842,N_23956);
or U24179 (N_24179,N_23585,N_23474);
xnor U24180 (N_24180,N_23578,N_23929);
or U24181 (N_24181,N_23409,N_23631);
and U24182 (N_24182,N_23461,N_23718);
nand U24183 (N_24183,N_23616,N_23791);
nor U24184 (N_24184,N_23574,N_23652);
nand U24185 (N_24185,N_23411,N_23715);
nand U24186 (N_24186,N_23795,N_23429);
xnor U24187 (N_24187,N_23659,N_23923);
or U24188 (N_24188,N_23733,N_23591);
or U24189 (N_24189,N_23423,N_23772);
and U24190 (N_24190,N_23564,N_23613);
and U24191 (N_24191,N_23846,N_23512);
or U24192 (N_24192,N_23454,N_23666);
xnor U24193 (N_24193,N_23988,N_23742);
xnor U24194 (N_24194,N_23502,N_23609);
and U24195 (N_24195,N_23818,N_23589);
nand U24196 (N_24196,N_23534,N_23462);
xor U24197 (N_24197,N_23481,N_23544);
and U24198 (N_24198,N_23679,N_23698);
nand U24199 (N_24199,N_23849,N_23962);
and U24200 (N_24200,N_23981,N_23949);
and U24201 (N_24201,N_23787,N_23852);
nor U24202 (N_24202,N_23457,N_23511);
nor U24203 (N_24203,N_23976,N_23830);
xnor U24204 (N_24204,N_23812,N_23643);
or U24205 (N_24205,N_23433,N_23894);
or U24206 (N_24206,N_23495,N_23854);
nand U24207 (N_24207,N_23487,N_23932);
nor U24208 (N_24208,N_23660,N_23963);
nand U24209 (N_24209,N_23615,N_23575);
nor U24210 (N_24210,N_23928,N_23703);
nand U24211 (N_24211,N_23612,N_23685);
or U24212 (N_24212,N_23506,N_23588);
nand U24213 (N_24213,N_23767,N_23635);
nor U24214 (N_24214,N_23905,N_23541);
and U24215 (N_24215,N_23804,N_23579);
and U24216 (N_24216,N_23622,N_23822);
xnor U24217 (N_24217,N_23467,N_23799);
or U24218 (N_24218,N_23524,N_23614);
nor U24219 (N_24219,N_23421,N_23783);
and U24220 (N_24220,N_23814,N_23707);
or U24221 (N_24221,N_23425,N_23816);
or U24222 (N_24222,N_23424,N_23497);
nand U24223 (N_24223,N_23508,N_23744);
xnor U24224 (N_24224,N_23642,N_23412);
or U24225 (N_24225,N_23696,N_23665);
xor U24226 (N_24226,N_23651,N_23721);
xnor U24227 (N_24227,N_23890,N_23734);
xor U24228 (N_24228,N_23871,N_23863);
xor U24229 (N_24229,N_23568,N_23805);
xor U24230 (N_24230,N_23657,N_23510);
nand U24231 (N_24231,N_23802,N_23836);
xor U24232 (N_24232,N_23784,N_23889);
nand U24233 (N_24233,N_23931,N_23903);
or U24234 (N_24234,N_23452,N_23948);
nor U24235 (N_24235,N_23909,N_23674);
nor U24236 (N_24236,N_23576,N_23493);
or U24237 (N_24237,N_23780,N_23925);
xnor U24238 (N_24238,N_23910,N_23716);
xor U24239 (N_24239,N_23986,N_23619);
xnor U24240 (N_24240,N_23870,N_23691);
nand U24241 (N_24241,N_23403,N_23427);
xnor U24242 (N_24242,N_23803,N_23514);
and U24243 (N_24243,N_23687,N_23595);
xor U24244 (N_24244,N_23789,N_23983);
or U24245 (N_24245,N_23862,N_23810);
or U24246 (N_24246,N_23594,N_23486);
and U24247 (N_24247,N_23766,N_23670);
or U24248 (N_24248,N_23865,N_23610);
xor U24249 (N_24249,N_23490,N_23741);
nor U24250 (N_24250,N_23908,N_23730);
or U24251 (N_24251,N_23794,N_23601);
or U24252 (N_24252,N_23947,N_23542);
nor U24253 (N_24253,N_23479,N_23866);
and U24254 (N_24254,N_23845,N_23719);
or U24255 (N_24255,N_23874,N_23788);
xor U24256 (N_24256,N_23885,N_23531);
xor U24257 (N_24257,N_23644,N_23587);
xor U24258 (N_24258,N_23680,N_23422);
xor U24259 (N_24259,N_23535,N_23540);
nor U24260 (N_24260,N_23480,N_23554);
nor U24261 (N_24261,N_23987,N_23996);
nor U24262 (N_24262,N_23489,N_23558);
or U24263 (N_24263,N_23946,N_23966);
and U24264 (N_24264,N_23953,N_23491);
or U24265 (N_24265,N_23843,N_23551);
and U24266 (N_24266,N_23941,N_23748);
xnor U24267 (N_24267,N_23517,N_23857);
nor U24268 (N_24268,N_23543,N_23757);
or U24269 (N_24269,N_23717,N_23623);
xor U24270 (N_24270,N_23525,N_23872);
nand U24271 (N_24271,N_23406,N_23844);
nand U24272 (N_24272,N_23449,N_23785);
or U24273 (N_24273,N_23800,N_23504);
or U24274 (N_24274,N_23658,N_23546);
xnor U24275 (N_24275,N_23971,N_23896);
nor U24276 (N_24276,N_23444,N_23537);
xnor U24277 (N_24277,N_23625,N_23565);
xor U24278 (N_24278,N_23864,N_23973);
nor U24279 (N_24279,N_23743,N_23938);
nor U24280 (N_24280,N_23607,N_23503);
or U24281 (N_24281,N_23821,N_23705);
xor U24282 (N_24282,N_23706,N_23692);
and U24283 (N_24283,N_23655,N_23926);
and U24284 (N_24284,N_23649,N_23827);
xor U24285 (N_24285,N_23797,N_23831);
nor U24286 (N_24286,N_23723,N_23675);
nor U24287 (N_24287,N_23753,N_23713);
nand U24288 (N_24288,N_23699,N_23867);
xnor U24289 (N_24289,N_23972,N_23485);
xor U24290 (N_24290,N_23756,N_23943);
xnor U24291 (N_24291,N_23840,N_23548);
and U24292 (N_24292,N_23700,N_23920);
or U24293 (N_24293,N_23765,N_23501);
nor U24294 (N_24294,N_23891,N_23906);
and U24295 (N_24295,N_23410,N_23828);
nand U24296 (N_24296,N_23911,N_23897);
or U24297 (N_24297,N_23520,N_23935);
nor U24298 (N_24298,N_23970,N_23567);
xor U24299 (N_24299,N_23945,N_23420);
nor U24300 (N_24300,N_23754,N_23923);
or U24301 (N_24301,N_23705,N_23872);
or U24302 (N_24302,N_23785,N_23544);
nand U24303 (N_24303,N_23638,N_23607);
and U24304 (N_24304,N_23602,N_23815);
and U24305 (N_24305,N_23920,N_23946);
or U24306 (N_24306,N_23778,N_23744);
xnor U24307 (N_24307,N_23649,N_23502);
nor U24308 (N_24308,N_23723,N_23851);
and U24309 (N_24309,N_23885,N_23715);
nand U24310 (N_24310,N_23830,N_23772);
nor U24311 (N_24311,N_23642,N_23763);
or U24312 (N_24312,N_23741,N_23996);
xor U24313 (N_24313,N_23909,N_23496);
xnor U24314 (N_24314,N_23460,N_23993);
nor U24315 (N_24315,N_23813,N_23796);
nor U24316 (N_24316,N_23442,N_23810);
xor U24317 (N_24317,N_23640,N_23475);
xor U24318 (N_24318,N_23749,N_23695);
nand U24319 (N_24319,N_23821,N_23714);
and U24320 (N_24320,N_23608,N_23794);
or U24321 (N_24321,N_23764,N_23824);
nand U24322 (N_24322,N_23651,N_23647);
nor U24323 (N_24323,N_23754,N_23909);
nand U24324 (N_24324,N_23402,N_23413);
or U24325 (N_24325,N_23488,N_23415);
nand U24326 (N_24326,N_23565,N_23662);
nand U24327 (N_24327,N_23843,N_23620);
nand U24328 (N_24328,N_23665,N_23910);
or U24329 (N_24329,N_23765,N_23990);
nand U24330 (N_24330,N_23836,N_23880);
or U24331 (N_24331,N_23954,N_23845);
nand U24332 (N_24332,N_23665,N_23470);
xor U24333 (N_24333,N_23746,N_23415);
xnor U24334 (N_24334,N_23890,N_23599);
and U24335 (N_24335,N_23973,N_23818);
or U24336 (N_24336,N_23515,N_23720);
and U24337 (N_24337,N_23477,N_23480);
nor U24338 (N_24338,N_23528,N_23736);
nand U24339 (N_24339,N_23668,N_23582);
and U24340 (N_24340,N_23939,N_23990);
nand U24341 (N_24341,N_23720,N_23475);
nand U24342 (N_24342,N_23558,N_23642);
nand U24343 (N_24343,N_23716,N_23621);
nor U24344 (N_24344,N_23827,N_23631);
and U24345 (N_24345,N_23582,N_23456);
nand U24346 (N_24346,N_23749,N_23436);
xor U24347 (N_24347,N_23502,N_23443);
or U24348 (N_24348,N_23812,N_23551);
nor U24349 (N_24349,N_23736,N_23517);
nand U24350 (N_24350,N_23946,N_23485);
xnor U24351 (N_24351,N_23692,N_23940);
or U24352 (N_24352,N_23947,N_23744);
xor U24353 (N_24353,N_23809,N_23404);
xor U24354 (N_24354,N_23560,N_23969);
nor U24355 (N_24355,N_23793,N_23801);
nand U24356 (N_24356,N_23698,N_23418);
or U24357 (N_24357,N_23552,N_23882);
nand U24358 (N_24358,N_23885,N_23713);
nor U24359 (N_24359,N_23572,N_23741);
nor U24360 (N_24360,N_23935,N_23757);
xor U24361 (N_24361,N_23548,N_23735);
or U24362 (N_24362,N_23722,N_23612);
xor U24363 (N_24363,N_23712,N_23769);
and U24364 (N_24364,N_23714,N_23560);
or U24365 (N_24365,N_23887,N_23747);
and U24366 (N_24366,N_23680,N_23540);
or U24367 (N_24367,N_23638,N_23927);
nand U24368 (N_24368,N_23501,N_23979);
or U24369 (N_24369,N_23924,N_23874);
nor U24370 (N_24370,N_23871,N_23711);
xnor U24371 (N_24371,N_23810,N_23677);
xnor U24372 (N_24372,N_23998,N_23956);
nor U24373 (N_24373,N_23956,N_23510);
xor U24374 (N_24374,N_23985,N_23644);
xor U24375 (N_24375,N_23837,N_23895);
nand U24376 (N_24376,N_23473,N_23493);
nand U24377 (N_24377,N_23921,N_23441);
and U24378 (N_24378,N_23819,N_23852);
xor U24379 (N_24379,N_23456,N_23921);
nor U24380 (N_24380,N_23638,N_23717);
or U24381 (N_24381,N_23998,N_23583);
or U24382 (N_24382,N_23783,N_23757);
and U24383 (N_24383,N_23777,N_23891);
nand U24384 (N_24384,N_23471,N_23438);
xor U24385 (N_24385,N_23897,N_23652);
nand U24386 (N_24386,N_23440,N_23782);
nor U24387 (N_24387,N_23756,N_23896);
or U24388 (N_24388,N_23923,N_23619);
and U24389 (N_24389,N_23721,N_23948);
and U24390 (N_24390,N_23952,N_23517);
xor U24391 (N_24391,N_23941,N_23963);
nand U24392 (N_24392,N_23667,N_23478);
xor U24393 (N_24393,N_23521,N_23560);
or U24394 (N_24394,N_23408,N_23808);
and U24395 (N_24395,N_23635,N_23771);
or U24396 (N_24396,N_23914,N_23890);
and U24397 (N_24397,N_23887,N_23926);
or U24398 (N_24398,N_23737,N_23871);
and U24399 (N_24399,N_23904,N_23730);
nor U24400 (N_24400,N_23418,N_23604);
and U24401 (N_24401,N_23942,N_23815);
or U24402 (N_24402,N_23840,N_23989);
and U24403 (N_24403,N_23532,N_23797);
xor U24404 (N_24404,N_23488,N_23604);
nor U24405 (N_24405,N_23928,N_23637);
xor U24406 (N_24406,N_23704,N_23957);
nand U24407 (N_24407,N_23615,N_23671);
or U24408 (N_24408,N_23992,N_23784);
and U24409 (N_24409,N_23921,N_23868);
or U24410 (N_24410,N_23661,N_23912);
nor U24411 (N_24411,N_23651,N_23432);
xnor U24412 (N_24412,N_23986,N_23787);
and U24413 (N_24413,N_23501,N_23859);
or U24414 (N_24414,N_23693,N_23924);
and U24415 (N_24415,N_23814,N_23938);
or U24416 (N_24416,N_23947,N_23896);
and U24417 (N_24417,N_23845,N_23767);
or U24418 (N_24418,N_23779,N_23732);
and U24419 (N_24419,N_23696,N_23740);
nand U24420 (N_24420,N_23829,N_23708);
xnor U24421 (N_24421,N_23743,N_23983);
or U24422 (N_24422,N_23850,N_23945);
nand U24423 (N_24423,N_23835,N_23685);
and U24424 (N_24424,N_23721,N_23446);
and U24425 (N_24425,N_23401,N_23889);
nand U24426 (N_24426,N_23713,N_23584);
or U24427 (N_24427,N_23866,N_23797);
or U24428 (N_24428,N_23435,N_23952);
nor U24429 (N_24429,N_23617,N_23689);
nand U24430 (N_24430,N_23580,N_23678);
nor U24431 (N_24431,N_23625,N_23436);
or U24432 (N_24432,N_23878,N_23523);
nor U24433 (N_24433,N_23707,N_23942);
nand U24434 (N_24434,N_23818,N_23446);
or U24435 (N_24435,N_23839,N_23718);
nor U24436 (N_24436,N_23813,N_23919);
nor U24437 (N_24437,N_23452,N_23538);
xor U24438 (N_24438,N_23544,N_23728);
xor U24439 (N_24439,N_23819,N_23718);
nand U24440 (N_24440,N_23484,N_23755);
xor U24441 (N_24441,N_23439,N_23449);
xor U24442 (N_24442,N_23448,N_23484);
and U24443 (N_24443,N_23999,N_23550);
or U24444 (N_24444,N_23948,N_23578);
or U24445 (N_24445,N_23505,N_23508);
and U24446 (N_24446,N_23539,N_23931);
xnor U24447 (N_24447,N_23659,N_23541);
nand U24448 (N_24448,N_23416,N_23441);
xnor U24449 (N_24449,N_23765,N_23830);
nor U24450 (N_24450,N_23867,N_23604);
and U24451 (N_24451,N_23741,N_23783);
and U24452 (N_24452,N_23892,N_23812);
or U24453 (N_24453,N_23824,N_23668);
nor U24454 (N_24454,N_23892,N_23507);
nor U24455 (N_24455,N_23661,N_23827);
xnor U24456 (N_24456,N_23885,N_23810);
nand U24457 (N_24457,N_23987,N_23687);
nand U24458 (N_24458,N_23828,N_23956);
nand U24459 (N_24459,N_23517,N_23794);
and U24460 (N_24460,N_23785,N_23873);
or U24461 (N_24461,N_23839,N_23545);
nor U24462 (N_24462,N_23531,N_23788);
or U24463 (N_24463,N_23593,N_23730);
or U24464 (N_24464,N_23803,N_23460);
nor U24465 (N_24465,N_23827,N_23772);
or U24466 (N_24466,N_23906,N_23863);
nor U24467 (N_24467,N_23533,N_23634);
nor U24468 (N_24468,N_23942,N_23421);
nand U24469 (N_24469,N_23554,N_23743);
nor U24470 (N_24470,N_23904,N_23794);
xnor U24471 (N_24471,N_23474,N_23997);
nor U24472 (N_24472,N_23582,N_23919);
xor U24473 (N_24473,N_23814,N_23575);
nor U24474 (N_24474,N_23550,N_23985);
xnor U24475 (N_24475,N_23521,N_23463);
or U24476 (N_24476,N_23589,N_23449);
nand U24477 (N_24477,N_23600,N_23661);
xnor U24478 (N_24478,N_23812,N_23994);
nor U24479 (N_24479,N_23684,N_23844);
or U24480 (N_24480,N_23844,N_23619);
nor U24481 (N_24481,N_23661,N_23896);
nor U24482 (N_24482,N_23766,N_23897);
nand U24483 (N_24483,N_23735,N_23567);
nand U24484 (N_24484,N_23887,N_23433);
xor U24485 (N_24485,N_23593,N_23733);
nor U24486 (N_24486,N_23436,N_23445);
nor U24487 (N_24487,N_23658,N_23667);
and U24488 (N_24488,N_23633,N_23940);
nor U24489 (N_24489,N_23959,N_23540);
and U24490 (N_24490,N_23452,N_23544);
and U24491 (N_24491,N_23949,N_23716);
nand U24492 (N_24492,N_23974,N_23992);
and U24493 (N_24493,N_23436,N_23613);
nor U24494 (N_24494,N_23695,N_23933);
xnor U24495 (N_24495,N_23544,N_23942);
nor U24496 (N_24496,N_23527,N_23643);
nand U24497 (N_24497,N_23906,N_23526);
xor U24498 (N_24498,N_23765,N_23522);
nor U24499 (N_24499,N_23808,N_23699);
xor U24500 (N_24500,N_23494,N_23796);
nor U24501 (N_24501,N_23550,N_23770);
xor U24502 (N_24502,N_23903,N_23938);
nor U24503 (N_24503,N_23626,N_23780);
and U24504 (N_24504,N_23777,N_23623);
or U24505 (N_24505,N_23993,N_23521);
xor U24506 (N_24506,N_23510,N_23494);
nor U24507 (N_24507,N_23427,N_23938);
or U24508 (N_24508,N_23595,N_23912);
nand U24509 (N_24509,N_23589,N_23924);
nand U24510 (N_24510,N_23712,N_23700);
xor U24511 (N_24511,N_23827,N_23412);
nor U24512 (N_24512,N_23842,N_23875);
xnor U24513 (N_24513,N_23526,N_23439);
xor U24514 (N_24514,N_23792,N_23804);
or U24515 (N_24515,N_23790,N_23842);
and U24516 (N_24516,N_23599,N_23404);
nor U24517 (N_24517,N_23480,N_23838);
nand U24518 (N_24518,N_23928,N_23748);
nand U24519 (N_24519,N_23442,N_23577);
xnor U24520 (N_24520,N_23819,N_23585);
and U24521 (N_24521,N_23793,N_23415);
xor U24522 (N_24522,N_23681,N_23951);
and U24523 (N_24523,N_23711,N_23809);
nor U24524 (N_24524,N_23973,N_23887);
and U24525 (N_24525,N_23626,N_23850);
nor U24526 (N_24526,N_23885,N_23923);
and U24527 (N_24527,N_23590,N_23773);
nor U24528 (N_24528,N_23843,N_23443);
nor U24529 (N_24529,N_23470,N_23666);
and U24530 (N_24530,N_23573,N_23862);
and U24531 (N_24531,N_23474,N_23724);
and U24532 (N_24532,N_23934,N_23756);
xor U24533 (N_24533,N_23806,N_23940);
nand U24534 (N_24534,N_23829,N_23710);
and U24535 (N_24535,N_23594,N_23501);
nand U24536 (N_24536,N_23814,N_23621);
nor U24537 (N_24537,N_23768,N_23729);
and U24538 (N_24538,N_23749,N_23704);
nand U24539 (N_24539,N_23872,N_23839);
or U24540 (N_24540,N_23658,N_23712);
nor U24541 (N_24541,N_23799,N_23803);
xor U24542 (N_24542,N_23892,N_23620);
xnor U24543 (N_24543,N_23718,N_23945);
or U24544 (N_24544,N_23909,N_23753);
and U24545 (N_24545,N_23549,N_23432);
nand U24546 (N_24546,N_23446,N_23966);
or U24547 (N_24547,N_23749,N_23575);
nand U24548 (N_24548,N_23636,N_23640);
xor U24549 (N_24549,N_23516,N_23774);
or U24550 (N_24550,N_23616,N_23486);
nand U24551 (N_24551,N_23773,N_23976);
or U24552 (N_24552,N_23703,N_23537);
nor U24553 (N_24553,N_23459,N_23843);
nand U24554 (N_24554,N_23858,N_23893);
and U24555 (N_24555,N_23512,N_23529);
or U24556 (N_24556,N_23871,N_23616);
and U24557 (N_24557,N_23850,N_23914);
xor U24558 (N_24558,N_23587,N_23755);
and U24559 (N_24559,N_23996,N_23652);
xor U24560 (N_24560,N_23722,N_23485);
nor U24561 (N_24561,N_23709,N_23962);
or U24562 (N_24562,N_23725,N_23527);
or U24563 (N_24563,N_23771,N_23621);
nor U24564 (N_24564,N_23975,N_23575);
and U24565 (N_24565,N_23597,N_23796);
nor U24566 (N_24566,N_23446,N_23606);
xnor U24567 (N_24567,N_23530,N_23851);
nand U24568 (N_24568,N_23412,N_23534);
xor U24569 (N_24569,N_23616,N_23951);
and U24570 (N_24570,N_23430,N_23542);
or U24571 (N_24571,N_23543,N_23476);
nor U24572 (N_24572,N_23805,N_23551);
nand U24573 (N_24573,N_23561,N_23923);
nand U24574 (N_24574,N_23769,N_23846);
and U24575 (N_24575,N_23898,N_23417);
nor U24576 (N_24576,N_23844,N_23631);
xnor U24577 (N_24577,N_23578,N_23527);
nor U24578 (N_24578,N_23556,N_23874);
or U24579 (N_24579,N_23534,N_23855);
or U24580 (N_24580,N_23565,N_23484);
xnor U24581 (N_24581,N_23646,N_23560);
nand U24582 (N_24582,N_23513,N_23567);
or U24583 (N_24583,N_23443,N_23512);
nand U24584 (N_24584,N_23963,N_23410);
and U24585 (N_24585,N_23956,N_23808);
and U24586 (N_24586,N_23667,N_23955);
and U24587 (N_24587,N_23854,N_23819);
and U24588 (N_24588,N_23932,N_23871);
and U24589 (N_24589,N_23728,N_23855);
xnor U24590 (N_24590,N_23966,N_23891);
or U24591 (N_24591,N_23795,N_23857);
nand U24592 (N_24592,N_23434,N_23732);
nand U24593 (N_24593,N_23449,N_23606);
nand U24594 (N_24594,N_23756,N_23420);
and U24595 (N_24595,N_23879,N_23636);
xor U24596 (N_24596,N_23741,N_23593);
and U24597 (N_24597,N_23500,N_23631);
nor U24598 (N_24598,N_23573,N_23565);
nor U24599 (N_24599,N_23696,N_23457);
nand U24600 (N_24600,N_24137,N_24131);
nand U24601 (N_24601,N_24157,N_24335);
nand U24602 (N_24602,N_24149,N_24322);
or U24603 (N_24603,N_24105,N_24435);
or U24604 (N_24604,N_24141,N_24204);
xor U24605 (N_24605,N_24573,N_24410);
and U24606 (N_24606,N_24519,N_24097);
or U24607 (N_24607,N_24400,N_24262);
nor U24608 (N_24608,N_24499,N_24295);
xnor U24609 (N_24609,N_24445,N_24046);
nand U24610 (N_24610,N_24473,N_24255);
xor U24611 (N_24611,N_24050,N_24200);
nor U24612 (N_24612,N_24249,N_24480);
or U24613 (N_24613,N_24414,N_24083);
nor U24614 (N_24614,N_24011,N_24551);
nor U24615 (N_24615,N_24516,N_24508);
nor U24616 (N_24616,N_24206,N_24133);
and U24617 (N_24617,N_24224,N_24502);
and U24618 (N_24618,N_24201,N_24416);
nand U24619 (N_24619,N_24265,N_24254);
xnor U24620 (N_24620,N_24507,N_24504);
nand U24621 (N_24621,N_24205,N_24483);
xnor U24622 (N_24622,N_24260,N_24013);
nand U24623 (N_24623,N_24116,N_24577);
or U24624 (N_24624,N_24117,N_24037);
and U24625 (N_24625,N_24509,N_24014);
or U24626 (N_24626,N_24188,N_24309);
or U24627 (N_24627,N_24549,N_24110);
xnor U24628 (N_24628,N_24251,N_24066);
or U24629 (N_24629,N_24367,N_24020);
nor U24630 (N_24630,N_24015,N_24227);
nor U24631 (N_24631,N_24540,N_24217);
xor U24632 (N_24632,N_24554,N_24491);
nand U24633 (N_24633,N_24167,N_24271);
nand U24634 (N_24634,N_24183,N_24337);
nand U24635 (N_24635,N_24300,N_24542);
xnor U24636 (N_24636,N_24085,N_24379);
and U24637 (N_24637,N_24489,N_24594);
xor U24638 (N_24638,N_24590,N_24058);
or U24639 (N_24639,N_24510,N_24475);
xnor U24640 (N_24640,N_24144,N_24537);
nor U24641 (N_24641,N_24333,N_24469);
nor U24642 (N_24642,N_24592,N_24560);
nand U24643 (N_24643,N_24166,N_24041);
nand U24644 (N_24644,N_24082,N_24478);
nand U24645 (N_24645,N_24346,N_24017);
nor U24646 (N_24646,N_24488,N_24569);
nor U24647 (N_24647,N_24316,N_24004);
and U24648 (N_24648,N_24056,N_24016);
and U24649 (N_24649,N_24456,N_24222);
and U24650 (N_24650,N_24296,N_24436);
xor U24651 (N_24651,N_24425,N_24539);
nor U24652 (N_24652,N_24127,N_24282);
or U24653 (N_24653,N_24287,N_24395);
and U24654 (N_24654,N_24591,N_24186);
nand U24655 (N_24655,N_24274,N_24040);
xor U24656 (N_24656,N_24417,N_24595);
or U24657 (N_24657,N_24384,N_24026);
and U24658 (N_24658,N_24253,N_24360);
and U24659 (N_24659,N_24311,N_24428);
nand U24660 (N_24660,N_24567,N_24369);
nor U24661 (N_24661,N_24408,N_24441);
xnor U24662 (N_24662,N_24568,N_24241);
and U24663 (N_24663,N_24345,N_24124);
and U24664 (N_24664,N_24151,N_24107);
nor U24665 (N_24665,N_24388,N_24599);
and U24666 (N_24666,N_24429,N_24392);
xnor U24667 (N_24667,N_24242,N_24168);
or U24668 (N_24668,N_24520,N_24329);
and U24669 (N_24669,N_24457,N_24596);
nand U24670 (N_24670,N_24069,N_24459);
or U24671 (N_24671,N_24398,N_24315);
nor U24672 (N_24672,N_24263,N_24455);
and U24673 (N_24673,N_24012,N_24318);
and U24674 (N_24674,N_24173,N_24076);
nand U24675 (N_24675,N_24331,N_24356);
nand U24676 (N_24676,N_24177,N_24492);
nand U24677 (N_24677,N_24450,N_24299);
xnor U24678 (N_24678,N_24522,N_24405);
and U24679 (N_24679,N_24272,N_24449);
or U24680 (N_24680,N_24411,N_24008);
nand U24681 (N_24681,N_24171,N_24019);
nand U24682 (N_24682,N_24055,N_24108);
nor U24683 (N_24683,N_24024,N_24277);
and U24684 (N_24684,N_24039,N_24174);
xnor U24685 (N_24685,N_24317,N_24547);
and U24686 (N_24686,N_24556,N_24075);
nand U24687 (N_24687,N_24080,N_24303);
nor U24688 (N_24688,N_24098,N_24493);
nor U24689 (N_24689,N_24461,N_24434);
or U24690 (N_24690,N_24385,N_24028);
xor U24691 (N_24691,N_24235,N_24582);
nand U24692 (N_24692,N_24072,N_24348);
xor U24693 (N_24693,N_24120,N_24464);
xor U24694 (N_24694,N_24589,N_24094);
nor U24695 (N_24695,N_24021,N_24430);
xor U24696 (N_24696,N_24401,N_24158);
xnor U24697 (N_24697,N_24187,N_24529);
and U24698 (N_24698,N_24358,N_24324);
xor U24699 (N_24699,N_24178,N_24269);
xnor U24700 (N_24700,N_24454,N_24297);
or U24701 (N_24701,N_24139,N_24218);
nand U24702 (N_24702,N_24000,N_24472);
and U24703 (N_24703,N_24498,N_24555);
and U24704 (N_24704,N_24307,N_24354);
and U24705 (N_24705,N_24115,N_24340);
and U24706 (N_24706,N_24320,N_24285);
xnor U24707 (N_24707,N_24419,N_24163);
or U24708 (N_24708,N_24099,N_24409);
or U24709 (N_24709,N_24583,N_24598);
nor U24710 (N_24710,N_24413,N_24534);
xor U24711 (N_24711,N_24518,N_24128);
and U24712 (N_24712,N_24140,N_24258);
and U24713 (N_24713,N_24289,N_24193);
and U24714 (N_24714,N_24433,N_24361);
nor U24715 (N_24715,N_24372,N_24202);
nand U24716 (N_24716,N_24135,N_24197);
nand U24717 (N_24717,N_24334,N_24302);
nand U24718 (N_24718,N_24546,N_24572);
xnor U24719 (N_24719,N_24093,N_24484);
xnor U24720 (N_24720,N_24245,N_24383);
nand U24721 (N_24721,N_24264,N_24452);
xnor U24722 (N_24722,N_24138,N_24482);
or U24723 (N_24723,N_24387,N_24561);
xor U24724 (N_24724,N_24153,N_24389);
xor U24725 (N_24725,N_24581,N_24023);
nand U24726 (N_24726,N_24159,N_24181);
and U24727 (N_24727,N_24121,N_24172);
nor U24728 (N_24728,N_24544,N_24029);
nand U24729 (N_24729,N_24152,N_24091);
or U24730 (N_24730,N_24404,N_24347);
nand U24731 (N_24731,N_24460,N_24090);
or U24732 (N_24732,N_24330,N_24426);
nor U24733 (N_24733,N_24113,N_24027);
nor U24734 (N_24734,N_24286,N_24497);
nand U24735 (N_24735,N_24378,N_24585);
and U24736 (N_24736,N_24564,N_24043);
xor U24737 (N_24737,N_24374,N_24049);
or U24738 (N_24738,N_24463,N_24194);
nor U24739 (N_24739,N_24035,N_24240);
nand U24740 (N_24740,N_24382,N_24566);
and U24741 (N_24741,N_24146,N_24231);
nand U24742 (N_24742,N_24275,N_24185);
or U24743 (N_24743,N_24230,N_24095);
nor U24744 (N_24744,N_24225,N_24100);
and U24745 (N_24745,N_24437,N_24365);
nor U24746 (N_24746,N_24150,N_24246);
or U24747 (N_24747,N_24423,N_24009);
and U24748 (N_24748,N_24313,N_24057);
nand U24749 (N_24749,N_24070,N_24476);
or U24750 (N_24750,N_24189,N_24371);
nand U24751 (N_24751,N_24575,N_24030);
or U24752 (N_24752,N_24527,N_24326);
and U24753 (N_24753,N_24487,N_24524);
nand U24754 (N_24754,N_24276,N_24477);
nor U24755 (N_24755,N_24530,N_24068);
xnor U24756 (N_24756,N_24521,N_24310);
nor U24757 (N_24757,N_24257,N_24501);
xnor U24758 (N_24758,N_24448,N_24515);
nand U24759 (N_24759,N_24424,N_24281);
nand U24760 (N_24760,N_24001,N_24366);
nor U24761 (N_24761,N_24588,N_24526);
xnor U24762 (N_24762,N_24233,N_24535);
xor U24763 (N_24763,N_24044,N_24078);
and U24764 (N_24764,N_24129,N_24160);
and U24765 (N_24765,N_24209,N_24396);
nor U24766 (N_24766,N_24288,N_24081);
or U24767 (N_24767,N_24394,N_24215);
or U24768 (N_24768,N_24574,N_24418);
and U24769 (N_24769,N_24444,N_24119);
nor U24770 (N_24770,N_24471,N_24261);
xnor U24771 (N_24771,N_24351,N_24292);
or U24772 (N_24772,N_24352,N_24114);
and U24773 (N_24773,N_24208,N_24243);
nand U24774 (N_24774,N_24580,N_24031);
xnor U24775 (N_24775,N_24165,N_24213);
nand U24776 (N_24776,N_24373,N_24415);
or U24777 (N_24777,N_24237,N_24106);
nor U24778 (N_24778,N_24375,N_24370);
and U24779 (N_24779,N_24393,N_24479);
nand U24780 (N_24780,N_24247,N_24325);
nor U24781 (N_24781,N_24336,N_24118);
xor U24782 (N_24782,N_24362,N_24376);
nor U24783 (N_24783,N_24304,N_24431);
nand U24784 (N_24784,N_24164,N_24586);
nor U24785 (N_24785,N_24192,N_24350);
nor U24786 (N_24786,N_24503,N_24191);
xnor U24787 (N_24787,N_24543,N_24219);
nor U24788 (N_24788,N_24306,N_24481);
xor U24789 (N_24789,N_24541,N_24377);
and U24790 (N_24790,N_24273,N_24467);
nor U24791 (N_24791,N_24349,N_24528);
and U24792 (N_24792,N_24221,N_24060);
xor U24793 (N_24793,N_24147,N_24390);
nor U24794 (N_24794,N_24067,N_24584);
nor U24795 (N_24795,N_24223,N_24062);
xnor U24796 (N_24796,N_24368,N_24134);
nand U24797 (N_24797,N_24079,N_24283);
or U24798 (N_24798,N_24155,N_24406);
nand U24799 (N_24799,N_24339,N_24294);
and U24800 (N_24800,N_24517,N_24511);
xor U24801 (N_24801,N_24045,N_24111);
nand U24802 (N_24802,N_24018,N_24565);
nand U24803 (N_24803,N_24112,N_24327);
xnor U24804 (N_24804,N_24559,N_24064);
or U24805 (N_24805,N_24343,N_24136);
nand U24806 (N_24806,N_24447,N_24074);
or U24807 (N_24807,N_24293,N_24439);
nand U24808 (N_24808,N_24088,N_24195);
or U24809 (N_24809,N_24440,N_24196);
nand U24810 (N_24810,N_24451,N_24407);
xor U24811 (N_24811,N_24270,N_24256);
nand U24812 (N_24812,N_24006,N_24126);
and U24813 (N_24813,N_24506,N_24259);
and U24814 (N_24814,N_24156,N_24207);
xor U24815 (N_24815,N_24252,N_24402);
and U24816 (N_24816,N_24268,N_24130);
xor U24817 (N_24817,N_24513,N_24494);
or U24818 (N_24818,N_24446,N_24123);
nand U24819 (N_24819,N_24391,N_24470);
or U24820 (N_24820,N_24432,N_24438);
nor U24821 (N_24821,N_24364,N_24047);
nor U24822 (N_24822,N_24148,N_24280);
nor U24823 (N_24823,N_24397,N_24005);
nand U24824 (N_24824,N_24033,N_24442);
xnor U24825 (N_24825,N_24279,N_24234);
nand U24826 (N_24826,N_24571,N_24420);
or U24827 (N_24827,N_24216,N_24179);
and U24828 (N_24828,N_24576,N_24244);
and U24829 (N_24829,N_24278,N_24025);
nand U24830 (N_24830,N_24532,N_24175);
nand U24831 (N_24831,N_24063,N_24102);
or U24832 (N_24832,N_24579,N_24169);
or U24833 (N_24833,N_24089,N_24036);
nand U24834 (N_24834,N_24353,N_24465);
nand U24835 (N_24835,N_24061,N_24308);
and U24836 (N_24836,N_24338,N_24342);
nand U24837 (N_24837,N_24003,N_24236);
xor U24838 (N_24838,N_24239,N_24587);
nor U24839 (N_24839,N_24380,N_24314);
and U24840 (N_24840,N_24548,N_24474);
or U24841 (N_24841,N_24051,N_24466);
nor U24842 (N_24842,N_24512,N_24550);
nor U24843 (N_24843,N_24034,N_24284);
nor U24844 (N_24844,N_24570,N_24578);
nand U24845 (N_24845,N_24180,N_24562);
nor U24846 (N_24846,N_24162,N_24053);
nand U24847 (N_24847,N_24170,N_24220);
nand U24848 (N_24848,N_24022,N_24399);
and U24849 (N_24849,N_24104,N_24557);
nand U24850 (N_24850,N_24495,N_24238);
or U24851 (N_24851,N_24210,N_24531);
xor U24852 (N_24852,N_24533,N_24199);
and U24853 (N_24853,N_24002,N_24305);
nor U24854 (N_24854,N_24109,N_24071);
nor U24855 (N_24855,N_24563,N_24267);
nand U24856 (N_24856,N_24103,N_24010);
or U24857 (N_24857,N_24007,N_24505);
and U24858 (N_24858,N_24154,N_24077);
nand U24859 (N_24859,N_24341,N_24125);
nand U24860 (N_24860,N_24427,N_24212);
and U24861 (N_24861,N_24381,N_24176);
nor U24862 (N_24862,N_24211,N_24323);
nor U24863 (N_24863,N_24332,N_24096);
xnor U24864 (N_24864,N_24514,N_24558);
nand U24865 (N_24865,N_24232,N_24298);
xnor U24866 (N_24866,N_24048,N_24355);
nand U24867 (N_24867,N_24190,N_24363);
and U24868 (N_24868,N_24073,N_24228);
and U24869 (N_24869,N_24468,N_24143);
xnor U24870 (N_24870,N_24321,N_24038);
or U24871 (N_24871,N_24145,N_24301);
or U24872 (N_24872,N_24122,N_24182);
or U24873 (N_24873,N_24290,N_24065);
or U24874 (N_24874,N_24593,N_24042);
or U24875 (N_24875,N_24536,N_24403);
nand U24876 (N_24876,N_24291,N_24486);
or U24877 (N_24877,N_24059,N_24319);
nor U24878 (N_24878,N_24443,N_24086);
xnor U24879 (N_24879,N_24250,N_24490);
or U24880 (N_24880,N_24229,N_24184);
and U24881 (N_24881,N_24054,N_24084);
nand U24882 (N_24882,N_24421,N_24132);
nor U24883 (N_24883,N_24101,N_24525);
nand U24884 (N_24884,N_24226,N_24142);
nor U24885 (N_24885,N_24453,N_24500);
nand U24886 (N_24886,N_24422,N_24266);
or U24887 (N_24887,N_24553,N_24052);
nand U24888 (N_24888,N_24538,N_24032);
nand U24889 (N_24889,N_24496,N_24203);
and U24890 (N_24890,N_24328,N_24161);
xor U24891 (N_24891,N_24087,N_24523);
nand U24892 (N_24892,N_24458,N_24312);
xnor U24893 (N_24893,N_24597,N_24545);
or U24894 (N_24894,N_24248,N_24359);
or U24895 (N_24895,N_24198,N_24092);
nor U24896 (N_24896,N_24412,N_24462);
nand U24897 (N_24897,N_24552,N_24485);
nand U24898 (N_24898,N_24357,N_24344);
nand U24899 (N_24899,N_24214,N_24386);
nand U24900 (N_24900,N_24513,N_24448);
and U24901 (N_24901,N_24411,N_24439);
and U24902 (N_24902,N_24545,N_24397);
xnor U24903 (N_24903,N_24317,N_24262);
or U24904 (N_24904,N_24148,N_24551);
nand U24905 (N_24905,N_24336,N_24370);
or U24906 (N_24906,N_24084,N_24571);
xor U24907 (N_24907,N_24398,N_24341);
nand U24908 (N_24908,N_24073,N_24491);
or U24909 (N_24909,N_24330,N_24325);
and U24910 (N_24910,N_24175,N_24318);
and U24911 (N_24911,N_24198,N_24173);
xor U24912 (N_24912,N_24432,N_24426);
nor U24913 (N_24913,N_24251,N_24331);
nor U24914 (N_24914,N_24052,N_24327);
nand U24915 (N_24915,N_24501,N_24368);
nand U24916 (N_24916,N_24260,N_24155);
nor U24917 (N_24917,N_24417,N_24445);
xor U24918 (N_24918,N_24374,N_24227);
xnor U24919 (N_24919,N_24282,N_24027);
xnor U24920 (N_24920,N_24427,N_24114);
and U24921 (N_24921,N_24012,N_24265);
and U24922 (N_24922,N_24559,N_24209);
nor U24923 (N_24923,N_24194,N_24466);
or U24924 (N_24924,N_24320,N_24044);
xor U24925 (N_24925,N_24508,N_24315);
xnor U24926 (N_24926,N_24045,N_24583);
nand U24927 (N_24927,N_24162,N_24280);
and U24928 (N_24928,N_24517,N_24014);
or U24929 (N_24929,N_24362,N_24373);
and U24930 (N_24930,N_24501,N_24311);
or U24931 (N_24931,N_24013,N_24229);
xnor U24932 (N_24932,N_24160,N_24373);
nor U24933 (N_24933,N_24014,N_24433);
or U24934 (N_24934,N_24141,N_24309);
or U24935 (N_24935,N_24561,N_24312);
or U24936 (N_24936,N_24314,N_24050);
and U24937 (N_24937,N_24117,N_24074);
nand U24938 (N_24938,N_24178,N_24361);
or U24939 (N_24939,N_24581,N_24070);
and U24940 (N_24940,N_24453,N_24032);
xnor U24941 (N_24941,N_24477,N_24273);
or U24942 (N_24942,N_24528,N_24477);
or U24943 (N_24943,N_24415,N_24074);
xor U24944 (N_24944,N_24433,N_24136);
and U24945 (N_24945,N_24505,N_24281);
or U24946 (N_24946,N_24386,N_24502);
xor U24947 (N_24947,N_24548,N_24517);
or U24948 (N_24948,N_24371,N_24283);
nand U24949 (N_24949,N_24229,N_24505);
nor U24950 (N_24950,N_24583,N_24219);
nand U24951 (N_24951,N_24203,N_24098);
or U24952 (N_24952,N_24113,N_24404);
and U24953 (N_24953,N_24458,N_24459);
or U24954 (N_24954,N_24469,N_24405);
xor U24955 (N_24955,N_24391,N_24573);
or U24956 (N_24956,N_24198,N_24204);
or U24957 (N_24957,N_24357,N_24011);
nor U24958 (N_24958,N_24356,N_24132);
nor U24959 (N_24959,N_24439,N_24355);
or U24960 (N_24960,N_24312,N_24581);
or U24961 (N_24961,N_24115,N_24250);
and U24962 (N_24962,N_24144,N_24412);
nand U24963 (N_24963,N_24103,N_24226);
xnor U24964 (N_24964,N_24490,N_24346);
and U24965 (N_24965,N_24588,N_24210);
and U24966 (N_24966,N_24540,N_24054);
and U24967 (N_24967,N_24474,N_24371);
or U24968 (N_24968,N_24095,N_24399);
or U24969 (N_24969,N_24543,N_24235);
and U24970 (N_24970,N_24414,N_24221);
xnor U24971 (N_24971,N_24313,N_24170);
nand U24972 (N_24972,N_24254,N_24245);
nand U24973 (N_24973,N_24165,N_24591);
nor U24974 (N_24974,N_24307,N_24168);
xor U24975 (N_24975,N_24356,N_24351);
nand U24976 (N_24976,N_24293,N_24224);
and U24977 (N_24977,N_24209,N_24571);
nand U24978 (N_24978,N_24153,N_24272);
nor U24979 (N_24979,N_24362,N_24456);
xnor U24980 (N_24980,N_24329,N_24254);
xnor U24981 (N_24981,N_24114,N_24129);
or U24982 (N_24982,N_24467,N_24161);
or U24983 (N_24983,N_24306,N_24572);
nand U24984 (N_24984,N_24354,N_24246);
or U24985 (N_24985,N_24448,N_24158);
nor U24986 (N_24986,N_24324,N_24044);
or U24987 (N_24987,N_24232,N_24360);
nor U24988 (N_24988,N_24024,N_24390);
and U24989 (N_24989,N_24329,N_24188);
or U24990 (N_24990,N_24566,N_24240);
or U24991 (N_24991,N_24564,N_24490);
nand U24992 (N_24992,N_24454,N_24395);
or U24993 (N_24993,N_24212,N_24317);
xor U24994 (N_24994,N_24268,N_24008);
or U24995 (N_24995,N_24409,N_24165);
or U24996 (N_24996,N_24053,N_24033);
xor U24997 (N_24997,N_24434,N_24051);
xor U24998 (N_24998,N_24010,N_24527);
xnor U24999 (N_24999,N_24573,N_24464);
nor U25000 (N_25000,N_24132,N_24417);
or U25001 (N_25001,N_24539,N_24176);
and U25002 (N_25002,N_24531,N_24480);
and U25003 (N_25003,N_24042,N_24450);
or U25004 (N_25004,N_24350,N_24215);
nand U25005 (N_25005,N_24233,N_24343);
nand U25006 (N_25006,N_24015,N_24567);
xor U25007 (N_25007,N_24011,N_24314);
or U25008 (N_25008,N_24513,N_24088);
nor U25009 (N_25009,N_24072,N_24365);
nand U25010 (N_25010,N_24471,N_24175);
xnor U25011 (N_25011,N_24032,N_24465);
or U25012 (N_25012,N_24160,N_24387);
and U25013 (N_25013,N_24055,N_24143);
nor U25014 (N_25014,N_24599,N_24387);
and U25015 (N_25015,N_24375,N_24068);
nor U25016 (N_25016,N_24357,N_24184);
nand U25017 (N_25017,N_24197,N_24360);
or U25018 (N_25018,N_24358,N_24315);
nor U25019 (N_25019,N_24390,N_24076);
nor U25020 (N_25020,N_24038,N_24008);
nor U25021 (N_25021,N_24192,N_24032);
or U25022 (N_25022,N_24194,N_24175);
nand U25023 (N_25023,N_24197,N_24597);
and U25024 (N_25024,N_24272,N_24445);
nor U25025 (N_25025,N_24103,N_24204);
nand U25026 (N_25026,N_24129,N_24597);
and U25027 (N_25027,N_24063,N_24428);
nor U25028 (N_25028,N_24338,N_24276);
nand U25029 (N_25029,N_24368,N_24040);
or U25030 (N_25030,N_24214,N_24507);
or U25031 (N_25031,N_24214,N_24562);
or U25032 (N_25032,N_24576,N_24227);
nand U25033 (N_25033,N_24170,N_24528);
xnor U25034 (N_25034,N_24430,N_24234);
or U25035 (N_25035,N_24055,N_24278);
xnor U25036 (N_25036,N_24347,N_24352);
nor U25037 (N_25037,N_24186,N_24351);
and U25038 (N_25038,N_24393,N_24248);
and U25039 (N_25039,N_24356,N_24403);
nor U25040 (N_25040,N_24225,N_24569);
and U25041 (N_25041,N_24221,N_24257);
and U25042 (N_25042,N_24296,N_24020);
nand U25043 (N_25043,N_24365,N_24381);
and U25044 (N_25044,N_24149,N_24536);
nor U25045 (N_25045,N_24585,N_24327);
and U25046 (N_25046,N_24176,N_24528);
nand U25047 (N_25047,N_24141,N_24491);
nand U25048 (N_25048,N_24452,N_24350);
xnor U25049 (N_25049,N_24467,N_24217);
and U25050 (N_25050,N_24053,N_24152);
and U25051 (N_25051,N_24370,N_24159);
and U25052 (N_25052,N_24061,N_24113);
xnor U25053 (N_25053,N_24281,N_24096);
xor U25054 (N_25054,N_24035,N_24310);
and U25055 (N_25055,N_24552,N_24031);
or U25056 (N_25056,N_24379,N_24054);
or U25057 (N_25057,N_24090,N_24137);
nand U25058 (N_25058,N_24515,N_24194);
xnor U25059 (N_25059,N_24215,N_24137);
and U25060 (N_25060,N_24420,N_24132);
xnor U25061 (N_25061,N_24031,N_24041);
nand U25062 (N_25062,N_24290,N_24087);
or U25063 (N_25063,N_24352,N_24326);
or U25064 (N_25064,N_24441,N_24314);
or U25065 (N_25065,N_24021,N_24524);
or U25066 (N_25066,N_24167,N_24228);
and U25067 (N_25067,N_24131,N_24293);
and U25068 (N_25068,N_24510,N_24590);
and U25069 (N_25069,N_24320,N_24550);
xor U25070 (N_25070,N_24364,N_24198);
or U25071 (N_25071,N_24563,N_24352);
nor U25072 (N_25072,N_24441,N_24530);
nand U25073 (N_25073,N_24332,N_24458);
nand U25074 (N_25074,N_24340,N_24276);
and U25075 (N_25075,N_24204,N_24497);
nand U25076 (N_25076,N_24393,N_24208);
xor U25077 (N_25077,N_24530,N_24317);
xor U25078 (N_25078,N_24175,N_24109);
nor U25079 (N_25079,N_24582,N_24176);
or U25080 (N_25080,N_24560,N_24391);
nor U25081 (N_25081,N_24477,N_24383);
xor U25082 (N_25082,N_24514,N_24248);
nand U25083 (N_25083,N_24226,N_24562);
and U25084 (N_25084,N_24549,N_24139);
nand U25085 (N_25085,N_24569,N_24537);
nor U25086 (N_25086,N_24138,N_24313);
xor U25087 (N_25087,N_24213,N_24520);
xor U25088 (N_25088,N_24020,N_24532);
or U25089 (N_25089,N_24553,N_24411);
xor U25090 (N_25090,N_24454,N_24393);
xnor U25091 (N_25091,N_24367,N_24414);
nor U25092 (N_25092,N_24073,N_24406);
and U25093 (N_25093,N_24081,N_24061);
and U25094 (N_25094,N_24239,N_24584);
nand U25095 (N_25095,N_24201,N_24370);
or U25096 (N_25096,N_24147,N_24379);
xnor U25097 (N_25097,N_24434,N_24370);
xor U25098 (N_25098,N_24081,N_24012);
nor U25099 (N_25099,N_24410,N_24058);
nand U25100 (N_25100,N_24073,N_24355);
nor U25101 (N_25101,N_24211,N_24534);
xnor U25102 (N_25102,N_24199,N_24166);
nor U25103 (N_25103,N_24384,N_24048);
or U25104 (N_25104,N_24455,N_24213);
nand U25105 (N_25105,N_24307,N_24541);
xnor U25106 (N_25106,N_24223,N_24520);
or U25107 (N_25107,N_24174,N_24210);
and U25108 (N_25108,N_24262,N_24072);
xor U25109 (N_25109,N_24574,N_24437);
nand U25110 (N_25110,N_24009,N_24203);
nor U25111 (N_25111,N_24351,N_24217);
nor U25112 (N_25112,N_24385,N_24159);
nor U25113 (N_25113,N_24251,N_24403);
or U25114 (N_25114,N_24429,N_24407);
nor U25115 (N_25115,N_24575,N_24193);
nand U25116 (N_25116,N_24428,N_24127);
nor U25117 (N_25117,N_24170,N_24188);
nor U25118 (N_25118,N_24542,N_24367);
nand U25119 (N_25119,N_24344,N_24496);
nor U25120 (N_25120,N_24204,N_24243);
xor U25121 (N_25121,N_24117,N_24150);
or U25122 (N_25122,N_24547,N_24424);
or U25123 (N_25123,N_24428,N_24189);
xor U25124 (N_25124,N_24462,N_24591);
or U25125 (N_25125,N_24253,N_24120);
xnor U25126 (N_25126,N_24420,N_24027);
nor U25127 (N_25127,N_24293,N_24240);
nand U25128 (N_25128,N_24135,N_24334);
nor U25129 (N_25129,N_24457,N_24350);
or U25130 (N_25130,N_24476,N_24593);
xnor U25131 (N_25131,N_24480,N_24171);
xor U25132 (N_25132,N_24339,N_24302);
or U25133 (N_25133,N_24584,N_24295);
xor U25134 (N_25134,N_24231,N_24077);
or U25135 (N_25135,N_24501,N_24417);
nor U25136 (N_25136,N_24033,N_24591);
or U25137 (N_25137,N_24404,N_24365);
nor U25138 (N_25138,N_24269,N_24128);
nor U25139 (N_25139,N_24438,N_24433);
nand U25140 (N_25140,N_24226,N_24409);
xnor U25141 (N_25141,N_24157,N_24238);
and U25142 (N_25142,N_24497,N_24285);
xnor U25143 (N_25143,N_24120,N_24582);
and U25144 (N_25144,N_24081,N_24080);
and U25145 (N_25145,N_24293,N_24053);
xor U25146 (N_25146,N_24450,N_24018);
xnor U25147 (N_25147,N_24478,N_24326);
or U25148 (N_25148,N_24410,N_24057);
and U25149 (N_25149,N_24268,N_24155);
nor U25150 (N_25150,N_24370,N_24012);
and U25151 (N_25151,N_24329,N_24420);
xnor U25152 (N_25152,N_24211,N_24117);
nor U25153 (N_25153,N_24332,N_24021);
nand U25154 (N_25154,N_24002,N_24438);
nor U25155 (N_25155,N_24320,N_24065);
nor U25156 (N_25156,N_24539,N_24025);
nor U25157 (N_25157,N_24471,N_24176);
xor U25158 (N_25158,N_24309,N_24348);
nand U25159 (N_25159,N_24180,N_24078);
and U25160 (N_25160,N_24014,N_24396);
and U25161 (N_25161,N_24479,N_24236);
or U25162 (N_25162,N_24238,N_24359);
nand U25163 (N_25163,N_24007,N_24252);
and U25164 (N_25164,N_24348,N_24269);
and U25165 (N_25165,N_24499,N_24158);
and U25166 (N_25166,N_24316,N_24503);
nand U25167 (N_25167,N_24178,N_24364);
or U25168 (N_25168,N_24414,N_24403);
and U25169 (N_25169,N_24262,N_24585);
or U25170 (N_25170,N_24357,N_24335);
xor U25171 (N_25171,N_24403,N_24415);
or U25172 (N_25172,N_24486,N_24397);
xor U25173 (N_25173,N_24112,N_24429);
nand U25174 (N_25174,N_24047,N_24159);
or U25175 (N_25175,N_24201,N_24406);
nor U25176 (N_25176,N_24091,N_24367);
xor U25177 (N_25177,N_24363,N_24205);
nor U25178 (N_25178,N_24515,N_24388);
nor U25179 (N_25179,N_24255,N_24097);
or U25180 (N_25180,N_24431,N_24395);
nand U25181 (N_25181,N_24455,N_24479);
nand U25182 (N_25182,N_24494,N_24220);
nand U25183 (N_25183,N_24291,N_24347);
nand U25184 (N_25184,N_24473,N_24531);
or U25185 (N_25185,N_24287,N_24118);
nor U25186 (N_25186,N_24515,N_24127);
nand U25187 (N_25187,N_24230,N_24418);
or U25188 (N_25188,N_24018,N_24163);
xnor U25189 (N_25189,N_24181,N_24574);
nor U25190 (N_25190,N_24254,N_24225);
or U25191 (N_25191,N_24242,N_24301);
or U25192 (N_25192,N_24592,N_24389);
and U25193 (N_25193,N_24441,N_24578);
nor U25194 (N_25194,N_24385,N_24213);
nor U25195 (N_25195,N_24588,N_24069);
nor U25196 (N_25196,N_24163,N_24438);
and U25197 (N_25197,N_24252,N_24055);
nor U25198 (N_25198,N_24592,N_24024);
and U25199 (N_25199,N_24114,N_24381);
xnor U25200 (N_25200,N_24639,N_24940);
nor U25201 (N_25201,N_25095,N_25100);
nand U25202 (N_25202,N_25121,N_25105);
and U25203 (N_25203,N_24776,N_24739);
nor U25204 (N_25204,N_25139,N_24964);
or U25205 (N_25205,N_24990,N_24633);
nor U25206 (N_25206,N_24852,N_25012);
nand U25207 (N_25207,N_24996,N_24773);
or U25208 (N_25208,N_25190,N_25074);
and U25209 (N_25209,N_24758,N_25193);
nand U25210 (N_25210,N_25102,N_24982);
nor U25211 (N_25211,N_25017,N_24975);
nand U25212 (N_25212,N_24709,N_25091);
nand U25213 (N_25213,N_24632,N_24705);
and U25214 (N_25214,N_25056,N_24960);
nor U25215 (N_25215,N_24795,N_25134);
nor U25216 (N_25216,N_24707,N_24708);
xnor U25217 (N_25217,N_24903,N_24959);
nand U25218 (N_25218,N_24907,N_25042);
or U25219 (N_25219,N_25079,N_24906);
nand U25220 (N_25220,N_25089,N_25065);
and U25221 (N_25221,N_24703,N_24833);
and U25222 (N_25222,N_24650,N_24798);
xor U25223 (N_25223,N_24831,N_24863);
or U25224 (N_25224,N_25161,N_24944);
xor U25225 (N_25225,N_24896,N_24669);
xor U25226 (N_25226,N_25130,N_24656);
and U25227 (N_25227,N_25162,N_25137);
nor U25228 (N_25228,N_24814,N_24729);
nor U25229 (N_25229,N_25035,N_24718);
nand U25230 (N_25230,N_24929,N_25026);
and U25231 (N_25231,N_24822,N_25004);
nor U25232 (N_25232,N_24752,N_24989);
xnor U25233 (N_25233,N_24911,N_25033);
nor U25234 (N_25234,N_24726,N_24608);
nor U25235 (N_25235,N_24868,N_24934);
nand U25236 (N_25236,N_24757,N_24673);
nor U25237 (N_25237,N_25087,N_24775);
and U25238 (N_25238,N_25187,N_24979);
and U25239 (N_25239,N_24704,N_25093);
xnor U25240 (N_25240,N_25063,N_25126);
or U25241 (N_25241,N_25044,N_24935);
or U25242 (N_25242,N_25142,N_24654);
nor U25243 (N_25243,N_24671,N_24972);
nand U25244 (N_25244,N_24610,N_25133);
nor U25245 (N_25245,N_24751,N_24793);
and U25246 (N_25246,N_24600,N_25104);
xor U25247 (N_25247,N_24685,N_24987);
xnor U25248 (N_25248,N_25184,N_24785);
or U25249 (N_25249,N_24637,N_24862);
xor U25250 (N_25250,N_24895,N_24651);
xnor U25251 (N_25251,N_24627,N_25029);
xor U25252 (N_25252,N_24675,N_25173);
xnor U25253 (N_25253,N_24662,N_24614);
or U25254 (N_25254,N_24642,N_24908);
nand U25255 (N_25255,N_24869,N_24784);
or U25256 (N_25256,N_25051,N_24921);
xor U25257 (N_25257,N_25185,N_24783);
nor U25258 (N_25258,N_24786,N_24937);
and U25259 (N_25259,N_24838,N_24800);
nand U25260 (N_25260,N_24841,N_24927);
and U25261 (N_25261,N_25024,N_25101);
xnor U25262 (N_25262,N_24645,N_25103);
xor U25263 (N_25263,N_25144,N_24936);
and U25264 (N_25264,N_24950,N_24803);
nor U25265 (N_25265,N_24872,N_24667);
and U25266 (N_25266,N_25014,N_25171);
nor U25267 (N_25267,N_24696,N_25108);
nand U25268 (N_25268,N_24954,N_24680);
nor U25269 (N_25269,N_25107,N_24998);
nor U25270 (N_25270,N_25020,N_25088);
or U25271 (N_25271,N_24792,N_24628);
nor U25272 (N_25272,N_24962,N_25117);
xor U25273 (N_25273,N_24899,N_24794);
nand U25274 (N_25274,N_25048,N_25150);
and U25275 (N_25275,N_25147,N_24874);
xor U25276 (N_25276,N_24724,N_24860);
and U25277 (N_25277,N_25008,N_24687);
nand U25278 (N_25278,N_24678,N_25094);
nand U25279 (N_25279,N_25181,N_25077);
xor U25280 (N_25280,N_24988,N_25128);
and U25281 (N_25281,N_24859,N_24805);
and U25282 (N_25282,N_24603,N_24842);
nor U25283 (N_25283,N_25145,N_25198);
or U25284 (N_25284,N_25160,N_24880);
and U25285 (N_25285,N_24881,N_24867);
nor U25286 (N_25286,N_24605,N_25057);
or U25287 (N_25287,N_24712,N_24780);
nand U25288 (N_25288,N_24976,N_24985);
nor U25289 (N_25289,N_24886,N_25053);
nand U25290 (N_25290,N_24961,N_25152);
xnor U25291 (N_25291,N_25165,N_25006);
nor U25292 (N_25292,N_24636,N_24742);
nor U25293 (N_25293,N_24973,N_24733);
xor U25294 (N_25294,N_25169,N_24722);
or U25295 (N_25295,N_24723,N_24809);
nor U25296 (N_25296,N_24698,N_24821);
nor U25297 (N_25297,N_24778,N_24755);
nand U25298 (N_25298,N_24955,N_25052);
xor U25299 (N_25299,N_24661,N_24890);
and U25300 (N_25300,N_25143,N_24837);
and U25301 (N_25301,N_25031,N_25163);
or U25302 (N_25302,N_24725,N_24894);
xnor U25303 (N_25303,N_24966,N_24827);
and U25304 (N_25304,N_25156,N_24980);
nor U25305 (N_25305,N_24657,N_24682);
nand U25306 (N_25306,N_25076,N_25188);
nor U25307 (N_25307,N_24858,N_24690);
nor U25308 (N_25308,N_24735,N_24918);
or U25309 (N_25309,N_25129,N_24760);
nand U25310 (N_25310,N_25084,N_24638);
and U25311 (N_25311,N_25036,N_24931);
nor U25312 (N_25312,N_24787,N_25111);
and U25313 (N_25313,N_24801,N_25096);
or U25314 (N_25314,N_25039,N_24816);
or U25315 (N_25315,N_24702,N_24848);
and U25316 (N_25316,N_25009,N_24676);
nor U25317 (N_25317,N_24613,N_25168);
and U25318 (N_25318,N_25194,N_25186);
nor U25319 (N_25319,N_24963,N_25177);
xor U25320 (N_25320,N_25116,N_24953);
nor U25321 (N_25321,N_24655,N_25025);
nor U25322 (N_25322,N_25154,N_24991);
nand U25323 (N_25323,N_24641,N_24952);
xor U25324 (N_25324,N_24799,N_24635);
nand U25325 (N_25325,N_24909,N_24700);
nor U25326 (N_25326,N_25085,N_25131);
nand U25327 (N_25327,N_24839,N_25118);
or U25328 (N_25328,N_25183,N_24693);
or U25329 (N_25329,N_24728,N_24769);
or U25330 (N_25330,N_25174,N_24779);
xor U25331 (N_25331,N_24818,N_25010);
nor U25332 (N_25332,N_24802,N_24905);
nor U25333 (N_25333,N_24897,N_25066);
nor U25334 (N_25334,N_24796,N_25097);
xnor U25335 (N_25335,N_24840,N_24847);
or U25336 (N_25336,N_24994,N_24901);
nor U25337 (N_25337,N_24925,N_24995);
or U25338 (N_25338,N_25099,N_24932);
xor U25339 (N_25339,N_24766,N_24791);
or U25340 (N_25340,N_24813,N_24992);
and U25341 (N_25341,N_24767,N_24631);
nand U25342 (N_25342,N_25064,N_25112);
or U25343 (N_25343,N_24710,N_24970);
nor U25344 (N_25344,N_24744,N_24782);
or U25345 (N_25345,N_25070,N_25125);
and U25346 (N_25346,N_25019,N_24892);
nor U25347 (N_25347,N_24873,N_24745);
nand U25348 (N_25348,N_25069,N_25081);
nand U25349 (N_25349,N_24697,N_25197);
xnor U25350 (N_25350,N_24888,N_25092);
xnor U25351 (N_25351,N_24984,N_24734);
xnor U25352 (N_25352,N_24923,N_25192);
nand U25353 (N_25353,N_24889,N_24826);
or U25354 (N_25354,N_24945,N_24983);
nand U25355 (N_25355,N_25127,N_24715);
nor U25356 (N_25356,N_24753,N_25005);
xnor U25357 (N_25357,N_25027,N_24617);
or U25358 (N_25358,N_24939,N_25003);
nor U25359 (N_25359,N_24772,N_25106);
or U25360 (N_25360,N_24756,N_24870);
xnor U25361 (N_25361,N_24914,N_25001);
and U25362 (N_25362,N_24913,N_25062);
or U25363 (N_25363,N_24683,N_24618);
nor U25364 (N_25364,N_24777,N_25175);
xor U25365 (N_25365,N_24615,N_25055);
nor U25366 (N_25366,N_24688,N_24644);
or U25367 (N_25367,N_25196,N_24686);
nand U25368 (N_25368,N_24922,N_24653);
nand U25369 (N_25369,N_24928,N_24943);
nor U25370 (N_25370,N_25110,N_25155);
nor U25371 (N_25371,N_24851,N_24737);
nor U25372 (N_25372,N_24740,N_25030);
and U25373 (N_25373,N_24699,N_24967);
and U25374 (N_25374,N_24763,N_24820);
xnor U25375 (N_25375,N_25158,N_25141);
xor U25376 (N_25376,N_25086,N_24815);
nand U25377 (N_25377,N_24974,N_24789);
and U25378 (N_25378,N_24612,N_25140);
nor U25379 (N_25379,N_24665,N_25002);
nand U25380 (N_25380,N_24971,N_24659);
nor U25381 (N_25381,N_24692,N_25199);
xnor U25382 (N_25382,N_24843,N_24956);
or U25383 (N_25383,N_25123,N_24946);
nand U25384 (N_25384,N_24986,N_24817);
and U25385 (N_25385,N_24646,N_24717);
and U25386 (N_25386,N_25013,N_24706);
nor U25387 (N_25387,N_25159,N_24668);
or U25388 (N_25388,N_24748,N_25178);
nand U25389 (N_25389,N_24917,N_25045);
xnor U25390 (N_25390,N_24684,N_25059);
nand U25391 (N_25391,N_24749,N_24957);
nor U25392 (N_25392,N_24844,N_25195);
xor U25393 (N_25393,N_24711,N_24900);
or U25394 (N_25394,N_24808,N_25068);
nand U25395 (N_25395,N_24738,N_24611);
and U25396 (N_25396,N_25018,N_24604);
xor U25397 (N_25397,N_25061,N_24602);
nor U25398 (N_25398,N_24865,N_24915);
or U25399 (N_25399,N_24746,N_24884);
nand U25400 (N_25400,N_24965,N_24861);
nor U25401 (N_25401,N_24670,N_24771);
nor U25402 (N_25402,N_25016,N_24629);
and U25403 (N_25403,N_24770,N_24806);
or U25404 (N_25404,N_24616,N_24811);
nand U25405 (N_25405,N_25124,N_25000);
nor U25406 (N_25406,N_24910,N_24630);
nand U25407 (N_25407,N_25083,N_25149);
nor U25408 (N_25408,N_24864,N_25073);
nand U25409 (N_25409,N_24853,N_24649);
nor U25410 (N_25410,N_25176,N_24882);
nand U25411 (N_25411,N_25151,N_25109);
xor U25412 (N_25412,N_24621,N_24866);
xnor U25413 (N_25413,N_25034,N_25028);
nand U25414 (N_25414,N_24743,N_24926);
xnor U25415 (N_25415,N_24977,N_24804);
nand U25416 (N_25416,N_24930,N_24924);
or U25417 (N_25417,N_24878,N_25180);
xor U25418 (N_25418,N_24920,N_24741);
nor U25419 (N_25419,N_25040,N_24810);
nand U25420 (N_25420,N_24601,N_24713);
or U25421 (N_25421,N_25072,N_24736);
and U25422 (N_25422,N_24885,N_24640);
nor U25423 (N_25423,N_25078,N_24854);
nor U25424 (N_25424,N_25041,N_25120);
nand U25425 (N_25425,N_24781,N_25049);
and U25426 (N_25426,N_24647,N_24981);
nor U25427 (N_25427,N_25032,N_24902);
or U25428 (N_25428,N_24942,N_24807);
and U25429 (N_25429,N_24893,N_24721);
nor U25430 (N_25430,N_24879,N_24624);
xnor U25431 (N_25431,N_24819,N_24606);
and U25432 (N_25432,N_24919,N_25119);
nand U25433 (N_25433,N_24948,N_25037);
xnor U25434 (N_25434,N_25071,N_25090);
nand U25435 (N_25435,N_25167,N_24877);
nand U25436 (N_25436,N_24999,N_25075);
xor U25437 (N_25437,N_24949,N_24968);
and U25438 (N_25438,N_24719,N_24947);
or U25439 (N_25439,N_24625,N_25043);
nand U25440 (N_25440,N_24689,N_24658);
nand U25441 (N_25441,N_25113,N_24727);
xor U25442 (N_25442,N_24788,N_24828);
and U25443 (N_25443,N_24978,N_24695);
or U25444 (N_25444,N_24845,N_24761);
xor U25445 (N_25445,N_24876,N_25047);
xnor U25446 (N_25446,N_24857,N_25058);
or U25447 (N_25447,N_24823,N_25153);
or U25448 (N_25448,N_24829,N_24634);
nor U25449 (N_25449,N_25115,N_24648);
and U25450 (N_25450,N_24716,N_24730);
and U25451 (N_25451,N_25054,N_25038);
or U25452 (N_25452,N_25132,N_25011);
or U25453 (N_25453,N_24912,N_24679);
and U25454 (N_25454,N_25015,N_25060);
nand U25455 (N_25455,N_25138,N_24871);
nand U25456 (N_25456,N_24849,N_24732);
nand U25457 (N_25457,N_24855,N_24933);
and U25458 (N_25458,N_24835,N_24938);
nand U25459 (N_25459,N_24620,N_24759);
nand U25460 (N_25460,N_25082,N_25164);
and U25461 (N_25461,N_24754,N_25148);
or U25462 (N_25462,N_24666,N_24790);
xor U25463 (N_25463,N_25098,N_25007);
nand U25464 (N_25464,N_24875,N_25146);
and U25465 (N_25465,N_25080,N_24850);
nand U25466 (N_25466,N_24643,N_24660);
nor U25467 (N_25467,N_24887,N_24652);
or U25468 (N_25468,N_24694,N_24764);
and U25469 (N_25469,N_25172,N_24768);
xor U25470 (N_25470,N_24904,N_24836);
or U25471 (N_25471,N_24720,N_24731);
nand U25472 (N_25472,N_24762,N_24663);
nand U25473 (N_25473,N_24832,N_24672);
or U25474 (N_25474,N_25050,N_24714);
nor U25475 (N_25475,N_25179,N_24750);
nand U25476 (N_25476,N_25166,N_24993);
nor U25477 (N_25477,N_24997,N_24691);
and U25478 (N_25478,N_24969,N_24898);
xnor U25479 (N_25479,N_24747,N_24797);
xnor U25480 (N_25480,N_24765,N_25157);
nor U25481 (N_25481,N_25191,N_24677);
xnor U25482 (N_25482,N_24626,N_25135);
xnor U25483 (N_25483,N_25122,N_24916);
xnor U25484 (N_25484,N_25189,N_25170);
xnor U25485 (N_25485,N_24951,N_25136);
nand U25486 (N_25486,N_25021,N_24623);
nor U25487 (N_25487,N_24830,N_24622);
nand U25488 (N_25488,N_24846,N_24812);
nand U25489 (N_25489,N_24674,N_24681);
xnor U25490 (N_25490,N_25022,N_24883);
nor U25491 (N_25491,N_25067,N_24701);
xnor U25492 (N_25492,N_24834,N_25023);
or U25493 (N_25493,N_25046,N_24824);
nor U25494 (N_25494,N_24619,N_24958);
nor U25495 (N_25495,N_25114,N_24774);
and U25496 (N_25496,N_24609,N_25182);
or U25497 (N_25497,N_24941,N_24664);
xnor U25498 (N_25498,N_24891,N_24856);
nand U25499 (N_25499,N_24825,N_24607);
xor U25500 (N_25500,N_25111,N_25028);
nor U25501 (N_25501,N_25196,N_25085);
nor U25502 (N_25502,N_25169,N_24620);
or U25503 (N_25503,N_24759,N_24667);
nor U25504 (N_25504,N_25148,N_24669);
xnor U25505 (N_25505,N_24980,N_24721);
and U25506 (N_25506,N_24861,N_24701);
nor U25507 (N_25507,N_24699,N_24951);
or U25508 (N_25508,N_25039,N_24981);
or U25509 (N_25509,N_24862,N_24853);
and U25510 (N_25510,N_24719,N_24801);
nand U25511 (N_25511,N_25153,N_24738);
or U25512 (N_25512,N_24930,N_25002);
nor U25513 (N_25513,N_24799,N_25152);
xnor U25514 (N_25514,N_24621,N_25132);
nor U25515 (N_25515,N_25087,N_24744);
xor U25516 (N_25516,N_25142,N_24978);
and U25517 (N_25517,N_24743,N_24628);
xnor U25518 (N_25518,N_25159,N_24824);
and U25519 (N_25519,N_24802,N_24769);
xor U25520 (N_25520,N_24626,N_24606);
xor U25521 (N_25521,N_24896,N_24620);
nor U25522 (N_25522,N_24641,N_25121);
nor U25523 (N_25523,N_24856,N_24827);
nor U25524 (N_25524,N_24984,N_24649);
nand U25525 (N_25525,N_24858,N_25028);
nand U25526 (N_25526,N_25096,N_24645);
nand U25527 (N_25527,N_24973,N_24724);
xor U25528 (N_25528,N_24769,N_25037);
or U25529 (N_25529,N_24705,N_24810);
xor U25530 (N_25530,N_24952,N_24925);
xnor U25531 (N_25531,N_24772,N_24728);
nor U25532 (N_25532,N_25060,N_24624);
nand U25533 (N_25533,N_24819,N_25182);
nor U25534 (N_25534,N_25004,N_24703);
and U25535 (N_25535,N_24748,N_24632);
nand U25536 (N_25536,N_25151,N_24775);
nand U25537 (N_25537,N_25019,N_24796);
nand U25538 (N_25538,N_25180,N_24755);
or U25539 (N_25539,N_24980,N_24836);
xor U25540 (N_25540,N_24786,N_24902);
nand U25541 (N_25541,N_25039,N_24791);
or U25542 (N_25542,N_24627,N_25148);
and U25543 (N_25543,N_25016,N_24614);
nand U25544 (N_25544,N_24834,N_25119);
or U25545 (N_25545,N_24765,N_25026);
nand U25546 (N_25546,N_24636,N_24827);
nand U25547 (N_25547,N_24957,N_24603);
and U25548 (N_25548,N_25094,N_25021);
or U25549 (N_25549,N_24784,N_25070);
nor U25550 (N_25550,N_25085,N_24649);
or U25551 (N_25551,N_25010,N_24725);
and U25552 (N_25552,N_24806,N_25065);
nand U25553 (N_25553,N_25022,N_24909);
nor U25554 (N_25554,N_24752,N_24987);
nand U25555 (N_25555,N_24671,N_24717);
nand U25556 (N_25556,N_24603,N_25006);
or U25557 (N_25557,N_25170,N_24953);
xor U25558 (N_25558,N_25168,N_25015);
and U25559 (N_25559,N_25160,N_25034);
and U25560 (N_25560,N_24675,N_24708);
xnor U25561 (N_25561,N_24720,N_25028);
and U25562 (N_25562,N_24827,N_25102);
or U25563 (N_25563,N_24729,N_25043);
nor U25564 (N_25564,N_24996,N_24809);
or U25565 (N_25565,N_24678,N_24792);
or U25566 (N_25566,N_25001,N_25121);
nor U25567 (N_25567,N_25030,N_25098);
nor U25568 (N_25568,N_24742,N_24889);
nor U25569 (N_25569,N_24693,N_24608);
nor U25570 (N_25570,N_25101,N_24900);
nor U25571 (N_25571,N_24859,N_24695);
nor U25572 (N_25572,N_24618,N_24865);
xnor U25573 (N_25573,N_25129,N_24846);
nor U25574 (N_25574,N_24793,N_24891);
or U25575 (N_25575,N_25008,N_24793);
and U25576 (N_25576,N_24733,N_25046);
xor U25577 (N_25577,N_24881,N_24701);
or U25578 (N_25578,N_24908,N_24762);
or U25579 (N_25579,N_25103,N_25157);
or U25580 (N_25580,N_24863,N_24743);
nor U25581 (N_25581,N_24845,N_24984);
and U25582 (N_25582,N_25081,N_25194);
nor U25583 (N_25583,N_24634,N_24873);
nand U25584 (N_25584,N_25105,N_24996);
or U25585 (N_25585,N_25027,N_25048);
and U25586 (N_25586,N_24811,N_24878);
or U25587 (N_25587,N_25017,N_24710);
xnor U25588 (N_25588,N_25116,N_24728);
and U25589 (N_25589,N_24822,N_24962);
or U25590 (N_25590,N_24714,N_24976);
nor U25591 (N_25591,N_25149,N_24748);
xnor U25592 (N_25592,N_24733,N_24667);
nand U25593 (N_25593,N_24955,N_25103);
nand U25594 (N_25594,N_24887,N_25144);
nor U25595 (N_25595,N_25044,N_24868);
or U25596 (N_25596,N_25121,N_24998);
nand U25597 (N_25597,N_24738,N_24980);
nor U25598 (N_25598,N_25059,N_24833);
xor U25599 (N_25599,N_25023,N_25054);
nor U25600 (N_25600,N_25004,N_24684);
and U25601 (N_25601,N_25081,N_25115);
or U25602 (N_25602,N_25046,N_24709);
nand U25603 (N_25603,N_24740,N_24937);
nand U25604 (N_25604,N_24791,N_24690);
and U25605 (N_25605,N_25122,N_24696);
xnor U25606 (N_25606,N_24723,N_24669);
and U25607 (N_25607,N_25132,N_24738);
nand U25608 (N_25608,N_24851,N_24696);
nand U25609 (N_25609,N_24772,N_24828);
and U25610 (N_25610,N_24989,N_25060);
or U25611 (N_25611,N_25105,N_24859);
nor U25612 (N_25612,N_25110,N_25056);
nand U25613 (N_25613,N_25076,N_24678);
nand U25614 (N_25614,N_24709,N_24998);
xnor U25615 (N_25615,N_24817,N_24715);
nand U25616 (N_25616,N_24880,N_24841);
or U25617 (N_25617,N_24867,N_24703);
nand U25618 (N_25618,N_24798,N_25148);
nand U25619 (N_25619,N_25123,N_25199);
and U25620 (N_25620,N_24917,N_25142);
nor U25621 (N_25621,N_25057,N_24720);
or U25622 (N_25622,N_25140,N_25146);
xor U25623 (N_25623,N_24982,N_25157);
nand U25624 (N_25624,N_25193,N_24737);
nor U25625 (N_25625,N_24709,N_24724);
or U25626 (N_25626,N_24794,N_24647);
or U25627 (N_25627,N_24781,N_24870);
nand U25628 (N_25628,N_24755,N_24835);
xnor U25629 (N_25629,N_25026,N_24960);
xor U25630 (N_25630,N_24828,N_24633);
and U25631 (N_25631,N_25036,N_25014);
nand U25632 (N_25632,N_24743,N_24928);
nand U25633 (N_25633,N_24923,N_24638);
xnor U25634 (N_25634,N_24971,N_24741);
and U25635 (N_25635,N_24852,N_25185);
or U25636 (N_25636,N_24833,N_24999);
and U25637 (N_25637,N_25016,N_24806);
nor U25638 (N_25638,N_24742,N_25003);
nand U25639 (N_25639,N_25196,N_24876);
or U25640 (N_25640,N_25135,N_24723);
xnor U25641 (N_25641,N_24681,N_24652);
and U25642 (N_25642,N_25012,N_25195);
or U25643 (N_25643,N_24884,N_24677);
nor U25644 (N_25644,N_24868,N_25158);
xor U25645 (N_25645,N_25115,N_24806);
nand U25646 (N_25646,N_24801,N_24611);
and U25647 (N_25647,N_25066,N_25167);
and U25648 (N_25648,N_25096,N_25074);
xnor U25649 (N_25649,N_25010,N_25131);
and U25650 (N_25650,N_25059,N_25128);
xor U25651 (N_25651,N_24685,N_24821);
nand U25652 (N_25652,N_24854,N_24849);
nand U25653 (N_25653,N_24741,N_24661);
or U25654 (N_25654,N_24775,N_25138);
or U25655 (N_25655,N_24902,N_24710);
or U25656 (N_25656,N_24865,N_25058);
or U25657 (N_25657,N_24677,N_24934);
or U25658 (N_25658,N_25154,N_24820);
nor U25659 (N_25659,N_25036,N_24988);
and U25660 (N_25660,N_25080,N_24891);
or U25661 (N_25661,N_24820,N_25016);
and U25662 (N_25662,N_25087,N_25014);
nand U25663 (N_25663,N_24966,N_25198);
xnor U25664 (N_25664,N_25178,N_24712);
nand U25665 (N_25665,N_24727,N_25119);
or U25666 (N_25666,N_24869,N_25141);
or U25667 (N_25667,N_24853,N_25127);
or U25668 (N_25668,N_24818,N_24629);
nand U25669 (N_25669,N_25169,N_24909);
xor U25670 (N_25670,N_25194,N_25066);
or U25671 (N_25671,N_24703,N_25196);
and U25672 (N_25672,N_25085,N_25117);
or U25673 (N_25673,N_25114,N_25129);
xor U25674 (N_25674,N_24956,N_24661);
nand U25675 (N_25675,N_25036,N_24742);
nand U25676 (N_25676,N_24808,N_24713);
and U25677 (N_25677,N_24946,N_24934);
nor U25678 (N_25678,N_24785,N_25116);
nor U25679 (N_25679,N_25177,N_24873);
nor U25680 (N_25680,N_25058,N_24958);
xor U25681 (N_25681,N_25064,N_24608);
nor U25682 (N_25682,N_24969,N_24748);
or U25683 (N_25683,N_24668,N_25151);
xor U25684 (N_25684,N_24764,N_24681);
or U25685 (N_25685,N_24757,N_24813);
nand U25686 (N_25686,N_25189,N_25071);
and U25687 (N_25687,N_24774,N_24936);
and U25688 (N_25688,N_24705,N_25097);
nand U25689 (N_25689,N_24625,N_24982);
or U25690 (N_25690,N_24646,N_24682);
or U25691 (N_25691,N_25047,N_25027);
xor U25692 (N_25692,N_24655,N_24864);
nor U25693 (N_25693,N_25058,N_25169);
and U25694 (N_25694,N_24641,N_24779);
and U25695 (N_25695,N_24760,N_24627);
xnor U25696 (N_25696,N_24818,N_24724);
nand U25697 (N_25697,N_24892,N_24916);
or U25698 (N_25698,N_25144,N_24934);
and U25699 (N_25699,N_24774,N_25132);
nand U25700 (N_25700,N_24989,N_24691);
and U25701 (N_25701,N_25075,N_25151);
and U25702 (N_25702,N_24621,N_24826);
or U25703 (N_25703,N_25095,N_24904);
and U25704 (N_25704,N_24677,N_25179);
nand U25705 (N_25705,N_24863,N_25050);
nor U25706 (N_25706,N_24657,N_24666);
and U25707 (N_25707,N_24750,N_25173);
and U25708 (N_25708,N_25155,N_24891);
nor U25709 (N_25709,N_25017,N_24916);
nand U25710 (N_25710,N_25104,N_24800);
or U25711 (N_25711,N_25044,N_25001);
and U25712 (N_25712,N_24851,N_24991);
xor U25713 (N_25713,N_24946,N_24853);
nand U25714 (N_25714,N_25040,N_24910);
and U25715 (N_25715,N_24935,N_24684);
and U25716 (N_25716,N_24733,N_25033);
nor U25717 (N_25717,N_25131,N_24831);
xnor U25718 (N_25718,N_25146,N_24861);
xor U25719 (N_25719,N_25121,N_24936);
and U25720 (N_25720,N_25041,N_25103);
nor U25721 (N_25721,N_24835,N_25124);
nand U25722 (N_25722,N_24619,N_25135);
xor U25723 (N_25723,N_24997,N_24925);
nand U25724 (N_25724,N_24877,N_24938);
or U25725 (N_25725,N_24627,N_25006);
nand U25726 (N_25726,N_24814,N_25182);
xor U25727 (N_25727,N_25110,N_25003);
nor U25728 (N_25728,N_24701,N_24992);
nand U25729 (N_25729,N_24944,N_24987);
nand U25730 (N_25730,N_24773,N_24983);
nor U25731 (N_25731,N_25066,N_25128);
xor U25732 (N_25732,N_24711,N_25049);
xor U25733 (N_25733,N_24629,N_24604);
xor U25734 (N_25734,N_24881,N_24618);
nand U25735 (N_25735,N_24717,N_25011);
and U25736 (N_25736,N_25087,N_25139);
xnor U25737 (N_25737,N_24866,N_24878);
xor U25738 (N_25738,N_24904,N_25100);
or U25739 (N_25739,N_24620,N_24993);
nor U25740 (N_25740,N_24897,N_25044);
or U25741 (N_25741,N_25155,N_24986);
or U25742 (N_25742,N_24934,N_24861);
or U25743 (N_25743,N_24760,N_24675);
or U25744 (N_25744,N_24863,N_25138);
xor U25745 (N_25745,N_25193,N_24917);
nand U25746 (N_25746,N_24932,N_24794);
nand U25747 (N_25747,N_25089,N_24823);
nand U25748 (N_25748,N_24991,N_24968);
nand U25749 (N_25749,N_25166,N_24728);
and U25750 (N_25750,N_24917,N_24849);
xnor U25751 (N_25751,N_25066,N_24715);
nor U25752 (N_25752,N_24794,N_24702);
or U25753 (N_25753,N_24884,N_24982);
or U25754 (N_25754,N_24961,N_24653);
or U25755 (N_25755,N_25190,N_24706);
xor U25756 (N_25756,N_24865,N_24690);
or U25757 (N_25757,N_25132,N_24812);
nand U25758 (N_25758,N_25088,N_24817);
xor U25759 (N_25759,N_24744,N_24639);
nand U25760 (N_25760,N_24962,N_24788);
and U25761 (N_25761,N_24684,N_24747);
nor U25762 (N_25762,N_24986,N_25146);
and U25763 (N_25763,N_24760,N_24605);
or U25764 (N_25764,N_24760,N_24632);
or U25765 (N_25765,N_24875,N_24821);
nor U25766 (N_25766,N_24897,N_24853);
xor U25767 (N_25767,N_25097,N_24710);
xnor U25768 (N_25768,N_25096,N_24894);
and U25769 (N_25769,N_24893,N_25074);
or U25770 (N_25770,N_24795,N_24652);
xnor U25771 (N_25771,N_24975,N_24629);
xnor U25772 (N_25772,N_24783,N_25142);
and U25773 (N_25773,N_25054,N_25172);
or U25774 (N_25774,N_25112,N_24811);
or U25775 (N_25775,N_25161,N_25010);
xor U25776 (N_25776,N_25015,N_24994);
nand U25777 (N_25777,N_24663,N_24764);
and U25778 (N_25778,N_25062,N_24711);
and U25779 (N_25779,N_24758,N_24963);
and U25780 (N_25780,N_24951,N_24903);
and U25781 (N_25781,N_25000,N_24731);
nor U25782 (N_25782,N_24930,N_24732);
nand U25783 (N_25783,N_24984,N_24819);
nand U25784 (N_25784,N_24718,N_24866);
nand U25785 (N_25785,N_25180,N_25020);
and U25786 (N_25786,N_24924,N_25056);
xnor U25787 (N_25787,N_25169,N_24622);
and U25788 (N_25788,N_24952,N_25081);
nand U25789 (N_25789,N_24806,N_24826);
nor U25790 (N_25790,N_24930,N_24831);
nor U25791 (N_25791,N_24960,N_25042);
or U25792 (N_25792,N_24753,N_24691);
and U25793 (N_25793,N_24982,N_25138);
xor U25794 (N_25794,N_24604,N_25104);
and U25795 (N_25795,N_24868,N_24816);
nor U25796 (N_25796,N_24789,N_24899);
nor U25797 (N_25797,N_25010,N_24816);
and U25798 (N_25798,N_24969,N_25084);
or U25799 (N_25799,N_25151,N_24828);
and U25800 (N_25800,N_25485,N_25555);
or U25801 (N_25801,N_25597,N_25638);
or U25802 (N_25802,N_25502,N_25657);
nand U25803 (N_25803,N_25232,N_25786);
xor U25804 (N_25804,N_25358,N_25513);
xor U25805 (N_25805,N_25600,N_25571);
and U25806 (N_25806,N_25373,N_25443);
xor U25807 (N_25807,N_25576,N_25713);
nor U25808 (N_25808,N_25499,N_25315);
nand U25809 (N_25809,N_25663,N_25464);
or U25810 (N_25810,N_25265,N_25678);
xor U25811 (N_25811,N_25715,N_25740);
xor U25812 (N_25812,N_25533,N_25267);
xor U25813 (N_25813,N_25343,N_25551);
nand U25814 (N_25814,N_25703,N_25460);
or U25815 (N_25815,N_25418,N_25325);
or U25816 (N_25816,N_25553,N_25396);
xnor U25817 (N_25817,N_25369,N_25483);
nand U25818 (N_25818,N_25585,N_25293);
nor U25819 (N_25819,N_25581,N_25436);
nor U25820 (N_25820,N_25324,N_25428);
or U25821 (N_25821,N_25558,N_25213);
nand U25822 (N_25822,N_25363,N_25599);
and U25823 (N_25823,N_25276,N_25449);
and U25824 (N_25824,N_25775,N_25593);
nor U25825 (N_25825,N_25275,N_25298);
xor U25826 (N_25826,N_25210,N_25763);
nor U25827 (N_25827,N_25212,N_25783);
and U25828 (N_25828,N_25417,N_25227);
or U25829 (N_25829,N_25208,N_25580);
and U25830 (N_25830,N_25321,N_25257);
nor U25831 (N_25831,N_25730,N_25494);
or U25832 (N_25832,N_25221,N_25538);
nor U25833 (N_25833,N_25463,N_25525);
or U25834 (N_25834,N_25754,N_25259);
nor U25835 (N_25835,N_25587,N_25320);
or U25836 (N_25836,N_25468,N_25535);
nor U25837 (N_25837,N_25514,N_25640);
xnor U25838 (N_25838,N_25224,N_25313);
and U25839 (N_25839,N_25361,N_25731);
nor U25840 (N_25840,N_25537,N_25621);
nand U25841 (N_25841,N_25458,N_25771);
or U25842 (N_25842,N_25311,N_25602);
nand U25843 (N_25843,N_25431,N_25415);
xnor U25844 (N_25844,N_25302,N_25403);
or U25845 (N_25845,N_25500,N_25595);
nand U25846 (N_25846,N_25778,N_25798);
nor U25847 (N_25847,N_25296,N_25416);
nor U25848 (N_25848,N_25634,N_25242);
nor U25849 (N_25849,N_25498,N_25596);
or U25850 (N_25850,N_25491,N_25346);
nor U25851 (N_25851,N_25550,N_25256);
nor U25852 (N_25852,N_25216,N_25748);
and U25853 (N_25853,N_25618,N_25654);
and U25854 (N_25854,N_25753,N_25342);
and U25855 (N_25855,N_25479,N_25478);
or U25856 (N_25856,N_25223,N_25422);
nor U25857 (N_25857,N_25252,N_25359);
xnor U25858 (N_25858,N_25757,N_25307);
nand U25859 (N_25859,N_25531,N_25762);
or U25860 (N_25860,N_25316,N_25441);
nor U25861 (N_25861,N_25387,N_25787);
xnor U25862 (N_25862,N_25702,N_25374);
or U25863 (N_25863,N_25780,N_25506);
xor U25864 (N_25864,N_25345,N_25310);
xnor U25865 (N_25865,N_25523,N_25610);
or U25866 (N_25866,N_25413,N_25694);
nand U25867 (N_25867,N_25285,N_25706);
nor U25868 (N_25868,N_25250,N_25306);
and U25869 (N_25869,N_25240,N_25592);
or U25870 (N_25870,N_25288,N_25327);
nor U25871 (N_25871,N_25495,N_25652);
nor U25872 (N_25872,N_25639,N_25238);
and U25873 (N_25873,N_25789,N_25779);
xor U25874 (N_25874,N_25598,N_25386);
xnor U25875 (N_25875,N_25711,N_25727);
nand U25876 (N_25876,N_25329,N_25260);
and U25877 (N_25877,N_25318,N_25248);
nand U25878 (N_25878,N_25554,N_25527);
and U25879 (N_25879,N_25548,N_25644);
xnor U25880 (N_25880,N_25445,N_25247);
xor U25881 (N_25881,N_25225,N_25541);
nand U25882 (N_25882,N_25556,N_25718);
or U25883 (N_25883,N_25565,N_25628);
nand U25884 (N_25884,N_25701,N_25466);
nand U25885 (N_25885,N_25251,N_25394);
nand U25886 (N_25886,N_25672,N_25414);
nor U25887 (N_25887,N_25630,N_25734);
xor U25888 (N_25888,N_25666,N_25280);
or U25889 (N_25889,N_25217,N_25669);
xor U25890 (N_25890,N_25430,N_25360);
or U25891 (N_25891,N_25427,N_25381);
xor U25892 (N_25892,N_25222,N_25705);
nand U25893 (N_25893,N_25230,N_25620);
nand U25894 (N_25894,N_25425,N_25650);
nand U25895 (N_25895,N_25473,N_25333);
nor U25896 (N_25896,N_25658,N_25546);
nor U25897 (N_25897,N_25508,N_25207);
nor U25898 (N_25898,N_25467,N_25738);
nand U25899 (N_25899,N_25526,N_25680);
or U25900 (N_25900,N_25765,N_25564);
nand U25901 (N_25901,N_25661,N_25435);
or U25902 (N_25902,N_25612,N_25397);
and U25903 (N_25903,N_25563,N_25725);
xor U25904 (N_25904,N_25743,N_25235);
nor U25905 (N_25905,N_25690,N_25515);
nor U25906 (N_25906,N_25246,N_25699);
xor U25907 (N_25907,N_25660,N_25737);
nand U25908 (N_25908,N_25444,N_25291);
xnor U25909 (N_25909,N_25382,N_25354);
nor U25910 (N_25910,N_25736,N_25759);
nand U25911 (N_25911,N_25493,N_25542);
nand U25912 (N_25912,N_25557,N_25337);
or U25913 (N_25913,N_25351,N_25410);
and U25914 (N_25914,N_25352,N_25411);
or U25915 (N_25915,N_25398,N_25301);
and U25916 (N_25916,N_25206,N_25465);
and U25917 (N_25917,N_25353,N_25772);
nor U25918 (N_25918,N_25279,N_25512);
xor U25919 (N_25919,N_25401,N_25322);
nand U25920 (N_25920,N_25659,N_25627);
or U25921 (N_25921,N_25331,N_25745);
nand U25922 (N_25922,N_25579,N_25350);
xor U25923 (N_25923,N_25588,N_25231);
and U25924 (N_25924,N_25461,N_25481);
nor U25925 (N_25925,N_25237,N_25497);
nor U25926 (N_25926,N_25489,N_25408);
nor U25927 (N_25927,N_25670,N_25419);
and U25928 (N_25928,N_25604,N_25708);
nand U25929 (N_25929,N_25673,N_25214);
or U25930 (N_25930,N_25439,N_25603);
xnor U25931 (N_25931,N_25682,N_25613);
xor U25932 (N_25932,N_25539,N_25476);
xor U25933 (N_25933,N_25273,N_25501);
or U25934 (N_25934,N_25522,N_25685);
or U25935 (N_25935,N_25274,N_25510);
nor U25936 (N_25936,N_25590,N_25785);
and U25937 (N_25937,N_25283,N_25648);
nor U25938 (N_25938,N_25616,N_25761);
nor U25939 (N_25939,N_25432,N_25211);
or U25940 (N_25940,N_25450,N_25393);
xnor U25941 (N_25941,N_25392,N_25790);
nand U25942 (N_25942,N_25689,N_25543);
nor U25943 (N_25943,N_25426,N_25475);
xnor U25944 (N_25944,N_25601,N_25545);
and U25945 (N_25945,N_25304,N_25516);
or U25946 (N_25946,N_25675,N_25649);
xnor U25947 (N_25947,N_25243,N_25691);
and U25948 (N_25948,N_25496,N_25200);
nor U25949 (N_25949,N_25364,N_25295);
xnor U25950 (N_25950,N_25378,N_25536);
xnor U25951 (N_25951,N_25719,N_25629);
or U25952 (N_25952,N_25517,N_25794);
and U25953 (N_25953,N_25735,N_25299);
nor U25954 (N_25954,N_25375,N_25262);
nand U25955 (N_25955,N_25582,N_25334);
nand U25956 (N_25956,N_25755,N_25692);
or U25957 (N_25957,N_25693,N_25341);
or U25958 (N_25958,N_25561,N_25488);
and U25959 (N_25959,N_25747,N_25245);
nor U25960 (N_25960,N_25752,N_25606);
and U25961 (N_25961,N_25338,N_25609);
and U25962 (N_25962,N_25226,N_25560);
xor U25963 (N_25963,N_25671,N_25524);
and U25964 (N_25964,N_25717,N_25376);
nor U25965 (N_25965,N_25462,N_25332);
nand U25966 (N_25966,N_25688,N_25442);
or U25967 (N_25967,N_25277,N_25266);
or U25968 (N_25968,N_25455,N_25459);
nor U25969 (N_25969,N_25261,N_25319);
or U25970 (N_25970,N_25229,N_25328);
xor U25971 (N_25971,N_25236,N_25544);
xor U25972 (N_25972,N_25799,N_25647);
and U25973 (N_25973,N_25404,N_25440);
nand U25974 (N_25974,N_25220,N_25366);
nand U25975 (N_25975,N_25797,N_25684);
nor U25976 (N_25976,N_25710,N_25472);
xnor U25977 (N_25977,N_25339,N_25305);
or U25978 (N_25978,N_25656,N_25709);
nand U25979 (N_25979,N_25424,N_25782);
nand U25980 (N_25980,N_25619,N_25681);
xnor U25981 (N_25981,N_25309,N_25796);
and U25982 (N_25982,N_25480,N_25284);
nand U25983 (N_25983,N_25589,N_25287);
nand U25984 (N_25984,N_25389,N_25573);
xor U25985 (N_25985,N_25792,N_25697);
and U25986 (N_25986,N_25776,N_25509);
and U25987 (N_25987,N_25349,N_25570);
nand U25988 (N_25988,N_25209,N_25429);
nand U25989 (N_25989,N_25477,N_25269);
or U25990 (N_25990,N_25788,N_25712);
and U25991 (N_25991,N_25751,N_25739);
nand U25992 (N_25992,N_25335,N_25448);
xnor U25993 (N_25993,N_25219,N_25383);
xnor U25994 (N_25994,N_25294,N_25317);
xnor U25995 (N_25995,N_25552,N_25281);
xor U25996 (N_25996,N_25662,N_25664);
or U25997 (N_25997,N_25519,N_25744);
and U25998 (N_25998,N_25244,N_25676);
and U25999 (N_25999,N_25732,N_25340);
nor U26000 (N_26000,N_25434,N_25379);
or U26001 (N_26001,N_25559,N_25268);
xnor U26002 (N_26002,N_25721,N_25482);
xnor U26003 (N_26003,N_25453,N_25679);
xor U26004 (N_26004,N_25733,N_25380);
or U26005 (N_26005,N_25674,N_25258);
and U26006 (N_26006,N_25370,N_25578);
and U26007 (N_26007,N_25204,N_25687);
and U26008 (N_26008,N_25365,N_25764);
or U26009 (N_26009,N_25594,N_25653);
or U26010 (N_26010,N_25700,N_25270);
xor U26011 (N_26011,N_25769,N_25623);
and U26012 (N_26012,N_25577,N_25614);
nand U26013 (N_26013,N_25504,N_25202);
xnor U26014 (N_26014,N_25407,N_25749);
nor U26015 (N_26015,N_25271,N_25683);
nand U26016 (N_26016,N_25770,N_25726);
and U26017 (N_26017,N_25234,N_25724);
xnor U26018 (N_26018,N_25228,N_25547);
or U26019 (N_26019,N_25395,N_25469);
and U26020 (N_26020,N_25584,N_25507);
or U26021 (N_26021,N_25239,N_25312);
xnor U26022 (N_26022,N_25774,N_25323);
xnor U26023 (N_26023,N_25344,N_25487);
nor U26024 (N_26024,N_25528,N_25297);
nor U26025 (N_26025,N_25486,N_25446);
and U26026 (N_26026,N_25253,N_25503);
nand U26027 (N_26027,N_25384,N_25784);
nand U26028 (N_26028,N_25390,N_25409);
xor U26029 (N_26029,N_25300,N_25720);
or U26030 (N_26030,N_25677,N_25518);
xor U26031 (N_26031,N_25696,N_25750);
or U26032 (N_26032,N_25423,N_25215);
xor U26033 (N_26033,N_25474,N_25773);
nor U26034 (N_26034,N_25626,N_25583);
nor U26035 (N_26035,N_25308,N_25562);
nor U26036 (N_26036,N_25534,N_25686);
nor U26037 (N_26037,N_25406,N_25716);
nand U26038 (N_26038,N_25367,N_25420);
and U26039 (N_26039,N_25625,N_25667);
and U26040 (N_26040,N_25532,N_25767);
nand U26041 (N_26041,N_25633,N_25348);
nand U26042 (N_26042,N_25391,N_25605);
nor U26043 (N_26043,N_25303,N_25203);
nor U26044 (N_26044,N_25357,N_25549);
or U26045 (N_26045,N_25651,N_25611);
nand U26046 (N_26046,N_25540,N_25695);
and U26047 (N_26047,N_25723,N_25668);
and U26048 (N_26048,N_25632,N_25704);
nand U26049 (N_26049,N_25385,N_25286);
nand U26050 (N_26050,N_25766,N_25254);
and U26051 (N_26051,N_25511,N_25336);
nor U26052 (N_26052,N_25330,N_25452);
or U26053 (N_26053,N_25457,N_25471);
nor U26054 (N_26054,N_25362,N_25530);
nor U26055 (N_26055,N_25529,N_25567);
xnor U26056 (N_26056,N_25400,N_25249);
xnor U26057 (N_26057,N_25607,N_25746);
nand U26058 (N_26058,N_25722,N_25631);
or U26059 (N_26059,N_25665,N_25756);
or U26060 (N_26060,N_25314,N_25264);
or U26061 (N_26061,N_25290,N_25635);
xor U26062 (N_26062,N_25637,N_25728);
or U26063 (N_26063,N_25521,N_25470);
xnor U26064 (N_26064,N_25278,N_25624);
or U26065 (N_26065,N_25289,N_25622);
and U26066 (N_26066,N_25569,N_25201);
nor U26067 (N_26067,N_25641,N_25586);
or U26068 (N_26068,N_25795,N_25282);
and U26069 (N_26069,N_25575,N_25255);
and U26070 (N_26070,N_25456,N_25758);
nor U26071 (N_26071,N_25505,N_25781);
or U26072 (N_26072,N_25447,N_25572);
or U26073 (N_26073,N_25326,N_25741);
or U26074 (N_26074,N_25405,N_25272);
xnor U26075 (N_26075,N_25591,N_25402);
or U26076 (N_26076,N_25484,N_25388);
and U26077 (N_26077,N_25233,N_25791);
or U26078 (N_26078,N_25377,N_25642);
xor U26079 (N_26079,N_25421,N_25368);
nor U26080 (N_26080,N_25645,N_25454);
nor U26081 (N_26081,N_25437,N_25646);
nor U26082 (N_26082,N_25355,N_25714);
xor U26083 (N_26083,N_25636,N_25608);
nor U26084 (N_26084,N_25263,N_25615);
xnor U26085 (N_26085,N_25742,N_25574);
and U26086 (N_26086,N_25729,N_25371);
or U26087 (N_26087,N_25205,N_25707);
nand U26088 (N_26088,N_25218,N_25490);
nor U26089 (N_26089,N_25698,N_25372);
nand U26090 (N_26090,N_25655,N_25399);
and U26091 (N_26091,N_25768,N_25438);
or U26092 (N_26092,N_25777,N_25760);
nand U26093 (N_26093,N_25292,N_25566);
and U26094 (N_26094,N_25643,N_25568);
xor U26095 (N_26095,N_25520,N_25793);
xnor U26096 (N_26096,N_25433,N_25617);
nand U26097 (N_26097,N_25356,N_25241);
and U26098 (N_26098,N_25347,N_25412);
xor U26099 (N_26099,N_25451,N_25492);
xnor U26100 (N_26100,N_25644,N_25708);
nor U26101 (N_26101,N_25503,N_25771);
nor U26102 (N_26102,N_25757,N_25686);
nand U26103 (N_26103,N_25586,N_25471);
nand U26104 (N_26104,N_25617,N_25344);
or U26105 (N_26105,N_25295,N_25425);
xor U26106 (N_26106,N_25534,N_25675);
xnor U26107 (N_26107,N_25750,N_25370);
xnor U26108 (N_26108,N_25761,N_25361);
xnor U26109 (N_26109,N_25606,N_25699);
and U26110 (N_26110,N_25521,N_25239);
xnor U26111 (N_26111,N_25546,N_25206);
xor U26112 (N_26112,N_25541,N_25553);
nand U26113 (N_26113,N_25751,N_25772);
nand U26114 (N_26114,N_25431,N_25752);
or U26115 (N_26115,N_25646,N_25483);
xor U26116 (N_26116,N_25658,N_25540);
and U26117 (N_26117,N_25386,N_25585);
nor U26118 (N_26118,N_25484,N_25551);
or U26119 (N_26119,N_25783,N_25381);
nand U26120 (N_26120,N_25395,N_25258);
or U26121 (N_26121,N_25727,N_25737);
nand U26122 (N_26122,N_25589,N_25259);
xor U26123 (N_26123,N_25715,N_25675);
or U26124 (N_26124,N_25664,N_25631);
and U26125 (N_26125,N_25742,N_25480);
xor U26126 (N_26126,N_25581,N_25673);
nand U26127 (N_26127,N_25522,N_25382);
nand U26128 (N_26128,N_25570,N_25578);
nand U26129 (N_26129,N_25410,N_25419);
nand U26130 (N_26130,N_25421,N_25386);
and U26131 (N_26131,N_25530,N_25773);
or U26132 (N_26132,N_25618,N_25494);
nor U26133 (N_26133,N_25593,N_25306);
and U26134 (N_26134,N_25590,N_25255);
xnor U26135 (N_26135,N_25624,N_25558);
nand U26136 (N_26136,N_25673,N_25613);
xnor U26137 (N_26137,N_25230,N_25223);
and U26138 (N_26138,N_25735,N_25522);
nand U26139 (N_26139,N_25336,N_25364);
and U26140 (N_26140,N_25612,N_25419);
xnor U26141 (N_26141,N_25326,N_25581);
xnor U26142 (N_26142,N_25263,N_25572);
nand U26143 (N_26143,N_25749,N_25300);
nand U26144 (N_26144,N_25780,N_25744);
nor U26145 (N_26145,N_25461,N_25202);
and U26146 (N_26146,N_25614,N_25285);
and U26147 (N_26147,N_25300,N_25526);
xor U26148 (N_26148,N_25498,N_25617);
nor U26149 (N_26149,N_25671,N_25644);
xor U26150 (N_26150,N_25325,N_25450);
xnor U26151 (N_26151,N_25212,N_25581);
xor U26152 (N_26152,N_25367,N_25218);
nor U26153 (N_26153,N_25473,N_25290);
nand U26154 (N_26154,N_25251,N_25618);
nor U26155 (N_26155,N_25229,N_25430);
xnor U26156 (N_26156,N_25740,N_25335);
nor U26157 (N_26157,N_25712,N_25314);
nand U26158 (N_26158,N_25381,N_25236);
xnor U26159 (N_26159,N_25600,N_25583);
nand U26160 (N_26160,N_25610,N_25721);
xor U26161 (N_26161,N_25373,N_25642);
or U26162 (N_26162,N_25656,N_25466);
nor U26163 (N_26163,N_25311,N_25210);
or U26164 (N_26164,N_25765,N_25471);
and U26165 (N_26165,N_25539,N_25626);
xnor U26166 (N_26166,N_25483,N_25457);
and U26167 (N_26167,N_25784,N_25507);
or U26168 (N_26168,N_25462,N_25322);
and U26169 (N_26169,N_25353,N_25514);
xor U26170 (N_26170,N_25554,N_25773);
nand U26171 (N_26171,N_25539,N_25326);
or U26172 (N_26172,N_25535,N_25295);
or U26173 (N_26173,N_25588,N_25408);
nand U26174 (N_26174,N_25220,N_25590);
xor U26175 (N_26175,N_25708,N_25584);
or U26176 (N_26176,N_25594,N_25658);
nand U26177 (N_26177,N_25210,N_25559);
xor U26178 (N_26178,N_25285,N_25391);
or U26179 (N_26179,N_25509,N_25616);
nor U26180 (N_26180,N_25773,N_25223);
nand U26181 (N_26181,N_25204,N_25313);
nor U26182 (N_26182,N_25506,N_25390);
nor U26183 (N_26183,N_25386,N_25216);
xnor U26184 (N_26184,N_25503,N_25434);
or U26185 (N_26185,N_25757,N_25701);
nor U26186 (N_26186,N_25266,N_25642);
and U26187 (N_26187,N_25493,N_25480);
nor U26188 (N_26188,N_25688,N_25755);
and U26189 (N_26189,N_25691,N_25672);
xnor U26190 (N_26190,N_25708,N_25527);
and U26191 (N_26191,N_25613,N_25739);
nand U26192 (N_26192,N_25542,N_25223);
nor U26193 (N_26193,N_25456,N_25418);
and U26194 (N_26194,N_25444,N_25674);
or U26195 (N_26195,N_25633,N_25290);
nand U26196 (N_26196,N_25252,N_25612);
and U26197 (N_26197,N_25275,N_25664);
nand U26198 (N_26198,N_25517,N_25529);
nand U26199 (N_26199,N_25577,N_25285);
xor U26200 (N_26200,N_25285,N_25425);
or U26201 (N_26201,N_25614,N_25483);
nand U26202 (N_26202,N_25296,N_25669);
xnor U26203 (N_26203,N_25272,N_25701);
and U26204 (N_26204,N_25606,N_25246);
and U26205 (N_26205,N_25201,N_25206);
or U26206 (N_26206,N_25685,N_25289);
nor U26207 (N_26207,N_25674,N_25710);
nand U26208 (N_26208,N_25751,N_25448);
nand U26209 (N_26209,N_25740,N_25732);
and U26210 (N_26210,N_25442,N_25323);
and U26211 (N_26211,N_25251,N_25614);
xor U26212 (N_26212,N_25498,N_25299);
nor U26213 (N_26213,N_25221,N_25391);
nand U26214 (N_26214,N_25523,N_25749);
and U26215 (N_26215,N_25290,N_25202);
or U26216 (N_26216,N_25707,N_25570);
or U26217 (N_26217,N_25660,N_25495);
or U26218 (N_26218,N_25788,N_25477);
nand U26219 (N_26219,N_25357,N_25691);
or U26220 (N_26220,N_25556,N_25750);
and U26221 (N_26221,N_25573,N_25612);
and U26222 (N_26222,N_25705,N_25321);
and U26223 (N_26223,N_25536,N_25229);
and U26224 (N_26224,N_25548,N_25443);
and U26225 (N_26225,N_25555,N_25560);
nand U26226 (N_26226,N_25716,N_25732);
nand U26227 (N_26227,N_25470,N_25223);
nor U26228 (N_26228,N_25521,N_25455);
nand U26229 (N_26229,N_25459,N_25638);
nand U26230 (N_26230,N_25460,N_25713);
nand U26231 (N_26231,N_25596,N_25506);
and U26232 (N_26232,N_25322,N_25289);
nand U26233 (N_26233,N_25526,N_25213);
or U26234 (N_26234,N_25283,N_25708);
nand U26235 (N_26235,N_25223,N_25551);
xor U26236 (N_26236,N_25272,N_25461);
nand U26237 (N_26237,N_25253,N_25283);
and U26238 (N_26238,N_25306,N_25797);
or U26239 (N_26239,N_25361,N_25376);
or U26240 (N_26240,N_25791,N_25459);
xor U26241 (N_26241,N_25691,N_25579);
nor U26242 (N_26242,N_25709,N_25293);
nor U26243 (N_26243,N_25460,N_25421);
or U26244 (N_26244,N_25372,N_25533);
nor U26245 (N_26245,N_25575,N_25472);
and U26246 (N_26246,N_25392,N_25232);
or U26247 (N_26247,N_25426,N_25653);
nand U26248 (N_26248,N_25218,N_25586);
xnor U26249 (N_26249,N_25622,N_25368);
and U26250 (N_26250,N_25246,N_25357);
nand U26251 (N_26251,N_25587,N_25770);
nor U26252 (N_26252,N_25284,N_25265);
xor U26253 (N_26253,N_25564,N_25334);
or U26254 (N_26254,N_25464,N_25360);
xor U26255 (N_26255,N_25313,N_25493);
nor U26256 (N_26256,N_25287,N_25352);
and U26257 (N_26257,N_25682,N_25509);
nand U26258 (N_26258,N_25784,N_25270);
or U26259 (N_26259,N_25496,N_25771);
nand U26260 (N_26260,N_25265,N_25767);
nand U26261 (N_26261,N_25676,N_25442);
xnor U26262 (N_26262,N_25373,N_25410);
nand U26263 (N_26263,N_25721,N_25411);
or U26264 (N_26264,N_25354,N_25270);
and U26265 (N_26265,N_25722,N_25450);
xor U26266 (N_26266,N_25278,N_25320);
or U26267 (N_26267,N_25686,N_25500);
nand U26268 (N_26268,N_25763,N_25757);
or U26269 (N_26269,N_25200,N_25459);
and U26270 (N_26270,N_25685,N_25367);
nand U26271 (N_26271,N_25475,N_25248);
nand U26272 (N_26272,N_25395,N_25413);
nand U26273 (N_26273,N_25659,N_25334);
or U26274 (N_26274,N_25717,N_25444);
nand U26275 (N_26275,N_25230,N_25494);
nand U26276 (N_26276,N_25315,N_25568);
and U26277 (N_26277,N_25233,N_25439);
nor U26278 (N_26278,N_25440,N_25792);
nand U26279 (N_26279,N_25667,N_25243);
or U26280 (N_26280,N_25445,N_25208);
xnor U26281 (N_26281,N_25380,N_25283);
nor U26282 (N_26282,N_25421,N_25352);
and U26283 (N_26283,N_25562,N_25318);
nand U26284 (N_26284,N_25267,N_25552);
nand U26285 (N_26285,N_25651,N_25255);
and U26286 (N_26286,N_25318,N_25331);
or U26287 (N_26287,N_25781,N_25219);
nor U26288 (N_26288,N_25663,N_25558);
nor U26289 (N_26289,N_25656,N_25777);
nand U26290 (N_26290,N_25380,N_25445);
and U26291 (N_26291,N_25329,N_25297);
or U26292 (N_26292,N_25466,N_25532);
xor U26293 (N_26293,N_25329,N_25356);
or U26294 (N_26294,N_25523,N_25545);
and U26295 (N_26295,N_25731,N_25501);
nor U26296 (N_26296,N_25630,N_25249);
and U26297 (N_26297,N_25584,N_25344);
nand U26298 (N_26298,N_25749,N_25629);
or U26299 (N_26299,N_25670,N_25745);
or U26300 (N_26300,N_25408,N_25532);
and U26301 (N_26301,N_25470,N_25203);
nand U26302 (N_26302,N_25303,N_25419);
nor U26303 (N_26303,N_25555,N_25594);
nand U26304 (N_26304,N_25530,N_25560);
or U26305 (N_26305,N_25248,N_25660);
and U26306 (N_26306,N_25479,N_25436);
xor U26307 (N_26307,N_25502,N_25540);
and U26308 (N_26308,N_25467,N_25306);
and U26309 (N_26309,N_25388,N_25650);
xnor U26310 (N_26310,N_25638,N_25250);
nand U26311 (N_26311,N_25717,N_25499);
xnor U26312 (N_26312,N_25460,N_25363);
nand U26313 (N_26313,N_25620,N_25292);
and U26314 (N_26314,N_25666,N_25785);
xnor U26315 (N_26315,N_25253,N_25454);
or U26316 (N_26316,N_25709,N_25335);
or U26317 (N_26317,N_25535,N_25247);
or U26318 (N_26318,N_25762,N_25606);
nor U26319 (N_26319,N_25479,N_25713);
xor U26320 (N_26320,N_25767,N_25255);
or U26321 (N_26321,N_25720,N_25257);
nor U26322 (N_26322,N_25784,N_25799);
xnor U26323 (N_26323,N_25465,N_25425);
nor U26324 (N_26324,N_25384,N_25296);
xnor U26325 (N_26325,N_25331,N_25489);
xnor U26326 (N_26326,N_25508,N_25721);
or U26327 (N_26327,N_25486,N_25349);
xnor U26328 (N_26328,N_25665,N_25383);
nand U26329 (N_26329,N_25256,N_25618);
or U26330 (N_26330,N_25464,N_25739);
nor U26331 (N_26331,N_25600,N_25260);
and U26332 (N_26332,N_25525,N_25445);
or U26333 (N_26333,N_25422,N_25640);
xnor U26334 (N_26334,N_25432,N_25469);
nor U26335 (N_26335,N_25576,N_25761);
nand U26336 (N_26336,N_25652,N_25347);
or U26337 (N_26337,N_25279,N_25340);
nand U26338 (N_26338,N_25680,N_25525);
and U26339 (N_26339,N_25401,N_25603);
nand U26340 (N_26340,N_25281,N_25465);
nor U26341 (N_26341,N_25793,N_25546);
xnor U26342 (N_26342,N_25218,N_25294);
and U26343 (N_26343,N_25216,N_25549);
nand U26344 (N_26344,N_25389,N_25346);
nor U26345 (N_26345,N_25270,N_25319);
xor U26346 (N_26346,N_25343,N_25363);
and U26347 (N_26347,N_25206,N_25704);
nor U26348 (N_26348,N_25248,N_25641);
or U26349 (N_26349,N_25473,N_25363);
and U26350 (N_26350,N_25320,N_25752);
and U26351 (N_26351,N_25607,N_25631);
or U26352 (N_26352,N_25311,N_25459);
nand U26353 (N_26353,N_25414,N_25523);
or U26354 (N_26354,N_25346,N_25259);
nand U26355 (N_26355,N_25263,N_25697);
and U26356 (N_26356,N_25578,N_25580);
and U26357 (N_26357,N_25281,N_25667);
and U26358 (N_26358,N_25526,N_25401);
and U26359 (N_26359,N_25606,N_25375);
and U26360 (N_26360,N_25546,N_25290);
nand U26361 (N_26361,N_25623,N_25557);
and U26362 (N_26362,N_25716,N_25619);
nor U26363 (N_26363,N_25586,N_25648);
nor U26364 (N_26364,N_25393,N_25485);
nand U26365 (N_26365,N_25675,N_25523);
and U26366 (N_26366,N_25215,N_25717);
nor U26367 (N_26367,N_25431,N_25744);
xor U26368 (N_26368,N_25428,N_25561);
or U26369 (N_26369,N_25499,N_25746);
nand U26370 (N_26370,N_25731,N_25690);
nand U26371 (N_26371,N_25355,N_25748);
xnor U26372 (N_26372,N_25231,N_25787);
xnor U26373 (N_26373,N_25465,N_25357);
or U26374 (N_26374,N_25442,N_25371);
or U26375 (N_26375,N_25567,N_25214);
nor U26376 (N_26376,N_25544,N_25520);
nor U26377 (N_26377,N_25579,N_25322);
nor U26378 (N_26378,N_25768,N_25478);
xnor U26379 (N_26379,N_25713,N_25760);
or U26380 (N_26380,N_25498,N_25283);
and U26381 (N_26381,N_25458,N_25592);
nand U26382 (N_26382,N_25720,N_25629);
or U26383 (N_26383,N_25368,N_25718);
xnor U26384 (N_26384,N_25525,N_25497);
or U26385 (N_26385,N_25511,N_25750);
and U26386 (N_26386,N_25757,N_25488);
nand U26387 (N_26387,N_25573,N_25295);
and U26388 (N_26388,N_25309,N_25421);
or U26389 (N_26389,N_25532,N_25477);
nor U26390 (N_26390,N_25619,N_25356);
nand U26391 (N_26391,N_25747,N_25735);
xnor U26392 (N_26392,N_25792,N_25267);
nor U26393 (N_26393,N_25625,N_25583);
and U26394 (N_26394,N_25744,N_25279);
nor U26395 (N_26395,N_25767,N_25706);
nor U26396 (N_26396,N_25247,N_25497);
or U26397 (N_26397,N_25524,N_25286);
xor U26398 (N_26398,N_25290,N_25710);
nor U26399 (N_26399,N_25553,N_25712);
or U26400 (N_26400,N_25938,N_26217);
or U26401 (N_26401,N_26260,N_26091);
nor U26402 (N_26402,N_25931,N_26181);
or U26403 (N_26403,N_26030,N_25853);
xor U26404 (N_26404,N_25915,N_25945);
and U26405 (N_26405,N_26279,N_26148);
nor U26406 (N_26406,N_26241,N_26079);
nand U26407 (N_26407,N_26287,N_26055);
xnor U26408 (N_26408,N_25862,N_26142);
xnor U26409 (N_26409,N_25998,N_25811);
and U26410 (N_26410,N_26113,N_26196);
nor U26411 (N_26411,N_26311,N_26045);
nor U26412 (N_26412,N_26345,N_26304);
or U26413 (N_26413,N_26035,N_26203);
nor U26414 (N_26414,N_25967,N_25819);
xnor U26415 (N_26415,N_25993,N_25806);
nand U26416 (N_26416,N_25863,N_26152);
nor U26417 (N_26417,N_25954,N_25810);
xnor U26418 (N_26418,N_25939,N_26183);
nand U26419 (N_26419,N_25884,N_25930);
nor U26420 (N_26420,N_26115,N_26036);
nor U26421 (N_26421,N_26277,N_26065);
nor U26422 (N_26422,N_26157,N_26374);
or U26423 (N_26423,N_25836,N_26349);
nand U26424 (N_26424,N_26054,N_26352);
nor U26425 (N_26425,N_25844,N_25825);
nor U26426 (N_26426,N_25902,N_26368);
nor U26427 (N_26427,N_25981,N_25868);
nor U26428 (N_26428,N_26249,N_25969);
and U26429 (N_26429,N_25999,N_25929);
nand U26430 (N_26430,N_26110,N_26158);
nand U26431 (N_26431,N_26151,N_26307);
xor U26432 (N_26432,N_26117,N_26319);
xor U26433 (N_26433,N_26395,N_25928);
or U26434 (N_26434,N_25846,N_26165);
or U26435 (N_26435,N_26326,N_26250);
xnor U26436 (N_26436,N_26088,N_25943);
or U26437 (N_26437,N_25837,N_25818);
nor U26438 (N_26438,N_25947,N_25976);
nor U26439 (N_26439,N_25864,N_25869);
or U26440 (N_26440,N_25896,N_26338);
nor U26441 (N_26441,N_26232,N_26007);
and U26442 (N_26442,N_25879,N_26121);
or U26443 (N_26443,N_25962,N_26182);
and U26444 (N_26444,N_25982,N_26060);
xor U26445 (N_26445,N_25855,N_26147);
nor U26446 (N_26446,N_26206,N_26162);
nand U26447 (N_26447,N_25813,N_25859);
nor U26448 (N_26448,N_26372,N_26202);
and U26449 (N_26449,N_25833,N_26258);
nor U26450 (N_26450,N_26061,N_25804);
or U26451 (N_26451,N_26012,N_26118);
xor U26452 (N_26452,N_26062,N_25870);
or U26453 (N_26453,N_25839,N_26313);
nand U26454 (N_26454,N_25857,N_26233);
and U26455 (N_26455,N_26144,N_26131);
nor U26456 (N_26456,N_25906,N_25985);
nand U26457 (N_26457,N_26078,N_26041);
or U26458 (N_26458,N_26334,N_25914);
or U26459 (N_26459,N_26123,N_26024);
nor U26460 (N_26460,N_26090,N_25824);
or U26461 (N_26461,N_25838,N_25965);
xnor U26462 (N_26462,N_26263,N_26093);
nor U26463 (N_26463,N_26040,N_25856);
nor U26464 (N_26464,N_26239,N_26386);
nand U26465 (N_26465,N_26322,N_26316);
and U26466 (N_26466,N_26213,N_26317);
xnor U26467 (N_26467,N_25889,N_26120);
or U26468 (N_26468,N_26259,N_26101);
nor U26469 (N_26469,N_25968,N_25899);
and U26470 (N_26470,N_26300,N_26220);
nand U26471 (N_26471,N_26194,N_26132);
or U26472 (N_26472,N_26379,N_26298);
nor U26473 (N_26473,N_25877,N_26327);
nor U26474 (N_26474,N_26283,N_26017);
nand U26475 (N_26475,N_26247,N_25827);
and U26476 (N_26476,N_26265,N_26272);
and U26477 (N_26477,N_26029,N_25822);
xnor U26478 (N_26478,N_25988,N_26373);
or U26479 (N_26479,N_26053,N_26236);
xnor U26480 (N_26480,N_26080,N_26254);
nor U26481 (N_26481,N_26067,N_26375);
nor U26482 (N_26482,N_26240,N_26331);
nand U26483 (N_26483,N_26064,N_26310);
xor U26484 (N_26484,N_26149,N_25923);
xnor U26485 (N_26485,N_26398,N_26363);
and U26486 (N_26486,N_26177,N_26022);
and U26487 (N_26487,N_26021,N_26384);
nor U26488 (N_26488,N_26137,N_26222);
xor U26489 (N_26489,N_26167,N_26034);
nor U26490 (N_26490,N_26252,N_26256);
and U26491 (N_26491,N_25958,N_26002);
nand U26492 (N_26492,N_25867,N_25960);
nor U26493 (N_26493,N_26388,N_26225);
and U26494 (N_26494,N_26380,N_26290);
nor U26495 (N_26495,N_26377,N_26185);
nand U26496 (N_26496,N_26295,N_26020);
or U26497 (N_26497,N_25917,N_26369);
and U26498 (N_26498,N_26199,N_25955);
or U26499 (N_26499,N_25919,N_26156);
xnor U26500 (N_26500,N_26106,N_26362);
and U26501 (N_26501,N_25949,N_26336);
and U26502 (N_26502,N_25873,N_26238);
or U26503 (N_26503,N_25893,N_26235);
or U26504 (N_26504,N_25878,N_25886);
or U26505 (N_26505,N_26333,N_26321);
nor U26506 (N_26506,N_25888,N_26288);
nor U26507 (N_26507,N_26270,N_26178);
nand U26508 (N_26508,N_26297,N_25882);
nand U26509 (N_26509,N_25974,N_25934);
nand U26510 (N_26510,N_26069,N_26228);
xnor U26511 (N_26511,N_26130,N_26318);
and U26512 (N_26512,N_26289,N_25817);
nor U26513 (N_26513,N_25812,N_26072);
nand U26514 (N_26514,N_26046,N_26073);
nor U26515 (N_26515,N_26397,N_25894);
xor U26516 (N_26516,N_25950,N_26224);
or U26517 (N_26517,N_26248,N_26218);
nor U26518 (N_26518,N_26396,N_25875);
nand U26519 (N_26519,N_25858,N_26392);
and U26520 (N_26520,N_26221,N_26286);
and U26521 (N_26521,N_25935,N_25883);
and U26522 (N_26522,N_26089,N_26099);
xor U26523 (N_26523,N_26399,N_26096);
nand U26524 (N_26524,N_26074,N_26173);
xnor U26525 (N_26525,N_25995,N_25829);
or U26526 (N_26526,N_25924,N_25820);
nand U26527 (N_26527,N_25957,N_25849);
or U26528 (N_26528,N_26160,N_26006);
or U26529 (N_26529,N_26343,N_26138);
xor U26530 (N_26530,N_26100,N_26341);
or U26531 (N_26531,N_26266,N_26219);
xor U26532 (N_26532,N_25826,N_26269);
and U26533 (N_26533,N_25861,N_26299);
nor U26534 (N_26534,N_25892,N_26039);
and U26535 (N_26535,N_26105,N_25854);
xnor U26536 (N_26536,N_25904,N_26033);
and U26537 (N_26537,N_25800,N_25978);
xnor U26538 (N_26538,N_26284,N_26129);
xnor U26539 (N_26539,N_26070,N_26346);
and U26540 (N_26540,N_26009,N_26193);
nor U26541 (N_26541,N_26087,N_26174);
or U26542 (N_26542,N_25852,N_26107);
nor U26543 (N_26543,N_26223,N_25832);
nand U26544 (N_26544,N_25895,N_26214);
nand U26545 (N_26545,N_25953,N_26257);
nand U26546 (N_26546,N_25994,N_26188);
nor U26547 (N_26547,N_26303,N_26207);
nor U26548 (N_26548,N_25916,N_26348);
and U26549 (N_26549,N_26201,N_26355);
xor U26550 (N_26550,N_26198,N_26143);
or U26551 (N_26551,N_26075,N_25881);
xnor U26552 (N_26552,N_26382,N_26357);
and U26553 (N_26553,N_25921,N_25992);
xnor U26554 (N_26554,N_25940,N_26042);
nor U26555 (N_26555,N_26128,N_26013);
xnor U26556 (N_26556,N_26262,N_26049);
xor U26557 (N_26557,N_26347,N_25956);
and U26558 (N_26558,N_26216,N_26003);
xnor U26559 (N_26559,N_25808,N_25847);
nand U26560 (N_26560,N_25927,N_26351);
nor U26561 (N_26561,N_25959,N_26209);
xnor U26562 (N_26562,N_26164,N_26376);
nand U26563 (N_26563,N_25874,N_26169);
or U26564 (N_26564,N_26119,N_26367);
nor U26565 (N_26565,N_26385,N_26339);
xnor U26566 (N_26566,N_26251,N_25971);
nor U26567 (N_26567,N_26077,N_25807);
or U26568 (N_26568,N_26330,N_26175);
or U26569 (N_26569,N_26329,N_26011);
and U26570 (N_26570,N_26166,N_26189);
or U26571 (N_26571,N_25909,N_26186);
and U26572 (N_26572,N_26356,N_26378);
xor U26573 (N_26573,N_26212,N_26294);
or U26574 (N_26574,N_26058,N_26146);
nor U26575 (N_26575,N_25865,N_26155);
xnor U26576 (N_26576,N_25866,N_25823);
nand U26577 (N_26577,N_26387,N_26323);
xnor U26578 (N_26578,N_26227,N_26135);
nand U26579 (N_26579,N_26271,N_26141);
nor U26580 (N_26580,N_25880,N_25913);
and U26581 (N_26581,N_26028,N_26306);
nor U26582 (N_26582,N_26281,N_26163);
xnor U26583 (N_26583,N_25834,N_25845);
or U26584 (N_26584,N_26000,N_26176);
nand U26585 (N_26585,N_26004,N_26309);
or U26586 (N_26586,N_26047,N_25821);
xnor U26587 (N_26587,N_26057,N_26305);
or U26588 (N_26588,N_26255,N_25872);
nand U26589 (N_26589,N_26102,N_26342);
or U26590 (N_26590,N_26122,N_25871);
nor U26591 (N_26591,N_25805,N_25951);
xnor U26592 (N_26592,N_26001,N_26192);
nor U26593 (N_26593,N_25977,N_26094);
and U26594 (N_26594,N_26125,N_26184);
or U26595 (N_26595,N_25803,N_25876);
xnor U26596 (N_26596,N_25802,N_26180);
or U26597 (N_26597,N_25890,N_25941);
nand U26598 (N_26598,N_26126,N_26264);
nand U26599 (N_26599,N_26044,N_26237);
nand U26600 (N_26600,N_26320,N_25975);
or U26601 (N_26601,N_26086,N_25973);
nor U26602 (N_26602,N_26391,N_26145);
and U26603 (N_26603,N_25910,N_25987);
nand U26604 (N_26604,N_26084,N_25830);
nor U26605 (N_26605,N_26019,N_26066);
or U26606 (N_26606,N_26246,N_26280);
and U26607 (N_26607,N_26337,N_26171);
nor U26608 (N_26608,N_25936,N_26112);
and U26609 (N_26609,N_25848,N_25841);
nand U26610 (N_26610,N_25932,N_25897);
or U26611 (N_26611,N_25851,N_26393);
or U26612 (N_26612,N_26153,N_25952);
nor U26613 (N_26613,N_26332,N_26204);
or U26614 (N_26614,N_26063,N_26274);
xor U26615 (N_26615,N_26293,N_25963);
nor U26616 (N_26616,N_26353,N_25903);
and U26617 (N_26617,N_26302,N_26292);
nand U26618 (N_26618,N_26370,N_26104);
or U26619 (N_26619,N_26015,N_25925);
nor U26620 (N_26620,N_26031,N_25905);
xor U26621 (N_26621,N_26190,N_26010);
nor U26622 (N_26622,N_26200,N_26179);
and U26623 (N_26623,N_26359,N_26076);
nand U26624 (N_26624,N_26390,N_26159);
xnor U26625 (N_26625,N_25908,N_26161);
and U26626 (N_26626,N_26234,N_26325);
xor U26627 (N_26627,N_25937,N_26085);
nand U26628 (N_26628,N_26092,N_26328);
xnor U26629 (N_26629,N_26083,N_26139);
and U26630 (N_26630,N_25961,N_25997);
xor U26631 (N_26631,N_25991,N_26268);
nor U26632 (N_26632,N_26243,N_25814);
xnor U26633 (N_26633,N_26134,N_25986);
xnor U26634 (N_26634,N_26276,N_26038);
and U26635 (N_26635,N_26187,N_25801);
nand U26636 (N_26636,N_26071,N_26208);
xor U26637 (N_26637,N_26095,N_25933);
or U26638 (N_26638,N_25912,N_26026);
and U26639 (N_26639,N_26267,N_26050);
or U26640 (N_26640,N_25996,N_25920);
or U26641 (N_26641,N_26043,N_26124);
or U26642 (N_26642,N_25948,N_25887);
or U26643 (N_26643,N_26205,N_25850);
nand U26644 (N_26644,N_25840,N_25944);
xnor U26645 (N_26645,N_25835,N_26018);
xor U26646 (N_26646,N_26136,N_25891);
or U26647 (N_26647,N_26383,N_26114);
or U26648 (N_26648,N_26097,N_26324);
and U26649 (N_26649,N_25966,N_25972);
and U26650 (N_26650,N_25942,N_26282);
or U26651 (N_26651,N_26358,N_26344);
nand U26652 (N_26652,N_25970,N_26098);
or U26653 (N_26653,N_25860,N_26335);
xor U26654 (N_26654,N_25885,N_26168);
xor U26655 (N_26655,N_26261,N_25843);
or U26656 (N_26656,N_26048,N_26111);
nand U26657 (N_26657,N_26127,N_26230);
or U26658 (N_26658,N_26361,N_26366);
or U26659 (N_26659,N_25989,N_26301);
or U26660 (N_26660,N_25901,N_25815);
nor U26661 (N_26661,N_25980,N_25809);
nand U26662 (N_26662,N_26226,N_26025);
and U26663 (N_26663,N_26103,N_25964);
xor U26664 (N_26664,N_25911,N_26032);
and U26665 (N_26665,N_26244,N_25984);
and U26666 (N_26666,N_26014,N_25990);
nand U26667 (N_26667,N_25926,N_25907);
and U26668 (N_26668,N_25983,N_26016);
or U26669 (N_26669,N_26312,N_26210);
xnor U26670 (N_26670,N_26364,N_26037);
nor U26671 (N_26671,N_26197,N_26005);
and U26672 (N_26672,N_26215,N_26354);
and U26673 (N_26673,N_26109,N_25900);
xor U26674 (N_26674,N_25946,N_26023);
and U26675 (N_26675,N_26350,N_25979);
nor U26676 (N_26676,N_26315,N_25816);
or U26677 (N_26677,N_26273,N_26195);
or U26678 (N_26678,N_26108,N_26150);
nor U26679 (N_26679,N_26154,N_26371);
and U26680 (N_26680,N_26231,N_26081);
and U26681 (N_26681,N_26229,N_26056);
nor U26682 (N_26682,N_26116,N_26360);
xor U26683 (N_26683,N_25922,N_26245);
and U26684 (N_26684,N_25842,N_26172);
and U26685 (N_26685,N_26291,N_26278);
or U26686 (N_26686,N_26394,N_26051);
xnor U26687 (N_26687,N_26191,N_26340);
xor U26688 (N_26688,N_26253,N_26170);
xnor U26689 (N_26689,N_26068,N_26296);
and U26690 (N_26690,N_26381,N_26052);
xor U26691 (N_26691,N_26140,N_26211);
or U26692 (N_26692,N_25898,N_26059);
or U26693 (N_26693,N_25831,N_26008);
xor U26694 (N_26694,N_26027,N_26389);
or U26695 (N_26695,N_26133,N_26242);
xnor U26696 (N_26696,N_26082,N_25828);
xnor U26697 (N_26697,N_26365,N_26275);
nand U26698 (N_26698,N_26314,N_26285);
and U26699 (N_26699,N_25918,N_26308);
or U26700 (N_26700,N_26204,N_26253);
and U26701 (N_26701,N_25907,N_26311);
nand U26702 (N_26702,N_26140,N_25883);
and U26703 (N_26703,N_26043,N_26120);
nand U26704 (N_26704,N_25867,N_26180);
or U26705 (N_26705,N_26223,N_26059);
xnor U26706 (N_26706,N_26304,N_26134);
xor U26707 (N_26707,N_26247,N_26045);
nor U26708 (N_26708,N_26154,N_25804);
nand U26709 (N_26709,N_26050,N_26397);
xor U26710 (N_26710,N_26227,N_26365);
xnor U26711 (N_26711,N_26297,N_25874);
nand U26712 (N_26712,N_26356,N_25940);
xnor U26713 (N_26713,N_26019,N_25844);
and U26714 (N_26714,N_25899,N_26016);
nand U26715 (N_26715,N_26280,N_26040);
nor U26716 (N_26716,N_26025,N_26229);
xnor U26717 (N_26717,N_26280,N_25913);
xor U26718 (N_26718,N_25981,N_25948);
xor U26719 (N_26719,N_26311,N_26073);
or U26720 (N_26720,N_25857,N_25819);
or U26721 (N_26721,N_25991,N_26095);
or U26722 (N_26722,N_25865,N_26317);
or U26723 (N_26723,N_26003,N_26335);
xor U26724 (N_26724,N_26305,N_25834);
nor U26725 (N_26725,N_25916,N_25903);
nor U26726 (N_26726,N_25911,N_25914);
and U26727 (N_26727,N_26208,N_26001);
nor U26728 (N_26728,N_26215,N_25819);
xnor U26729 (N_26729,N_26167,N_25963);
xor U26730 (N_26730,N_26034,N_25939);
and U26731 (N_26731,N_26173,N_25961);
nor U26732 (N_26732,N_26392,N_26338);
or U26733 (N_26733,N_26223,N_26030);
nand U26734 (N_26734,N_26374,N_26186);
xnor U26735 (N_26735,N_25830,N_26008);
nor U26736 (N_26736,N_25998,N_26035);
nor U26737 (N_26737,N_26398,N_26243);
or U26738 (N_26738,N_26114,N_26297);
and U26739 (N_26739,N_25860,N_26327);
nor U26740 (N_26740,N_26328,N_25843);
xor U26741 (N_26741,N_26355,N_26082);
nand U26742 (N_26742,N_25859,N_26027);
and U26743 (N_26743,N_26230,N_25830);
nor U26744 (N_26744,N_26163,N_25982);
or U26745 (N_26745,N_26388,N_25848);
or U26746 (N_26746,N_25803,N_25836);
nand U26747 (N_26747,N_26272,N_25811);
xnor U26748 (N_26748,N_26188,N_26066);
or U26749 (N_26749,N_26112,N_26275);
xnor U26750 (N_26750,N_26249,N_26026);
and U26751 (N_26751,N_25813,N_26145);
nand U26752 (N_26752,N_25933,N_26326);
or U26753 (N_26753,N_25998,N_26167);
nand U26754 (N_26754,N_26368,N_26043);
xnor U26755 (N_26755,N_26294,N_25838);
xor U26756 (N_26756,N_25803,N_26342);
nand U26757 (N_26757,N_26226,N_26269);
and U26758 (N_26758,N_26304,N_26159);
nor U26759 (N_26759,N_26333,N_26265);
nand U26760 (N_26760,N_26379,N_25990);
and U26761 (N_26761,N_26277,N_26191);
or U26762 (N_26762,N_26098,N_26120);
and U26763 (N_26763,N_26354,N_26122);
or U26764 (N_26764,N_26030,N_26204);
xnor U26765 (N_26765,N_25870,N_25895);
nand U26766 (N_26766,N_25901,N_26352);
nor U26767 (N_26767,N_26046,N_26118);
xnor U26768 (N_26768,N_25835,N_26162);
xor U26769 (N_26769,N_25818,N_26207);
and U26770 (N_26770,N_25819,N_26279);
nand U26771 (N_26771,N_26345,N_26165);
nand U26772 (N_26772,N_25977,N_26194);
xnor U26773 (N_26773,N_25878,N_26293);
nand U26774 (N_26774,N_26261,N_26221);
nor U26775 (N_26775,N_26322,N_25909);
nand U26776 (N_26776,N_26246,N_25805);
and U26777 (N_26777,N_26310,N_26195);
or U26778 (N_26778,N_26006,N_26142);
and U26779 (N_26779,N_26180,N_25944);
nor U26780 (N_26780,N_26061,N_26019);
nor U26781 (N_26781,N_26365,N_25871);
xnor U26782 (N_26782,N_26014,N_26224);
nand U26783 (N_26783,N_25825,N_26389);
or U26784 (N_26784,N_26107,N_26123);
and U26785 (N_26785,N_25924,N_26214);
and U26786 (N_26786,N_26324,N_26211);
and U26787 (N_26787,N_26042,N_25960);
nor U26788 (N_26788,N_26371,N_26235);
or U26789 (N_26789,N_26027,N_26235);
or U26790 (N_26790,N_26248,N_25974);
nor U26791 (N_26791,N_26061,N_26345);
and U26792 (N_26792,N_26248,N_26247);
nand U26793 (N_26793,N_26187,N_26302);
nor U26794 (N_26794,N_26077,N_25860);
and U26795 (N_26795,N_25800,N_26346);
nand U26796 (N_26796,N_25831,N_26379);
or U26797 (N_26797,N_26390,N_25822);
or U26798 (N_26798,N_26336,N_25832);
and U26799 (N_26799,N_26360,N_26007);
and U26800 (N_26800,N_26300,N_25812);
or U26801 (N_26801,N_25828,N_26028);
or U26802 (N_26802,N_26197,N_25867);
and U26803 (N_26803,N_25886,N_26285);
nand U26804 (N_26804,N_25992,N_26010);
and U26805 (N_26805,N_26054,N_26332);
xnor U26806 (N_26806,N_25889,N_25966);
or U26807 (N_26807,N_26090,N_25879);
nand U26808 (N_26808,N_25920,N_26110);
and U26809 (N_26809,N_25952,N_26232);
xnor U26810 (N_26810,N_25972,N_25807);
nor U26811 (N_26811,N_26078,N_26161);
nor U26812 (N_26812,N_25830,N_26083);
or U26813 (N_26813,N_26259,N_25912);
or U26814 (N_26814,N_26112,N_26029);
xnor U26815 (N_26815,N_26241,N_25880);
nor U26816 (N_26816,N_26041,N_26030);
nor U26817 (N_26817,N_26098,N_25835);
and U26818 (N_26818,N_26171,N_25917);
nor U26819 (N_26819,N_25838,N_26338);
nor U26820 (N_26820,N_26214,N_26381);
or U26821 (N_26821,N_25894,N_26163);
nor U26822 (N_26822,N_26211,N_25909);
nor U26823 (N_26823,N_26056,N_25954);
nand U26824 (N_26824,N_25910,N_26061);
and U26825 (N_26825,N_26156,N_26242);
and U26826 (N_26826,N_26243,N_25948);
and U26827 (N_26827,N_26051,N_26119);
xor U26828 (N_26828,N_25804,N_25945);
nor U26829 (N_26829,N_26274,N_26318);
nor U26830 (N_26830,N_25817,N_26293);
xnor U26831 (N_26831,N_25885,N_26071);
nand U26832 (N_26832,N_26351,N_26339);
or U26833 (N_26833,N_26060,N_26071);
and U26834 (N_26834,N_25824,N_26064);
xor U26835 (N_26835,N_26170,N_26305);
and U26836 (N_26836,N_26268,N_26299);
xor U26837 (N_26837,N_26235,N_26236);
xnor U26838 (N_26838,N_26114,N_25838);
or U26839 (N_26839,N_26185,N_25807);
and U26840 (N_26840,N_26030,N_26392);
or U26841 (N_26841,N_26155,N_25862);
xor U26842 (N_26842,N_25822,N_25823);
or U26843 (N_26843,N_26202,N_25847);
or U26844 (N_26844,N_25878,N_25991);
or U26845 (N_26845,N_26027,N_26065);
nand U26846 (N_26846,N_26368,N_26196);
xor U26847 (N_26847,N_26198,N_26350);
or U26848 (N_26848,N_26116,N_26219);
or U26849 (N_26849,N_26243,N_26371);
or U26850 (N_26850,N_25977,N_25973);
nand U26851 (N_26851,N_26301,N_25928);
or U26852 (N_26852,N_25936,N_25909);
or U26853 (N_26853,N_25923,N_25816);
or U26854 (N_26854,N_26048,N_25980);
nor U26855 (N_26855,N_26008,N_26110);
or U26856 (N_26856,N_26336,N_26398);
nand U26857 (N_26857,N_25819,N_26267);
or U26858 (N_26858,N_26282,N_25918);
nor U26859 (N_26859,N_25819,N_25843);
or U26860 (N_26860,N_25801,N_26213);
xnor U26861 (N_26861,N_26198,N_26294);
nand U26862 (N_26862,N_26361,N_26151);
nor U26863 (N_26863,N_25944,N_25964);
and U26864 (N_26864,N_25897,N_26303);
xnor U26865 (N_26865,N_26238,N_26263);
or U26866 (N_26866,N_26162,N_25873);
nor U26867 (N_26867,N_26033,N_25841);
nor U26868 (N_26868,N_26257,N_26129);
xor U26869 (N_26869,N_26194,N_26136);
nor U26870 (N_26870,N_26331,N_25876);
nor U26871 (N_26871,N_26161,N_26238);
xnor U26872 (N_26872,N_26236,N_25927);
nand U26873 (N_26873,N_26107,N_26006);
or U26874 (N_26874,N_26373,N_25985);
or U26875 (N_26875,N_25809,N_26175);
xor U26876 (N_26876,N_26066,N_26228);
xnor U26877 (N_26877,N_26233,N_26058);
or U26878 (N_26878,N_26252,N_26217);
and U26879 (N_26879,N_26178,N_26321);
and U26880 (N_26880,N_26158,N_25865);
nand U26881 (N_26881,N_26295,N_26209);
nor U26882 (N_26882,N_26033,N_26160);
nor U26883 (N_26883,N_25900,N_26337);
or U26884 (N_26884,N_26187,N_26176);
and U26885 (N_26885,N_26310,N_26171);
nand U26886 (N_26886,N_26145,N_26253);
or U26887 (N_26887,N_26264,N_26226);
xor U26888 (N_26888,N_26103,N_26151);
nor U26889 (N_26889,N_26062,N_26050);
nand U26890 (N_26890,N_26049,N_26156);
nand U26891 (N_26891,N_26390,N_25992);
and U26892 (N_26892,N_25895,N_26035);
nor U26893 (N_26893,N_26005,N_26204);
and U26894 (N_26894,N_26170,N_26306);
or U26895 (N_26895,N_25885,N_25818);
or U26896 (N_26896,N_26376,N_26072);
nand U26897 (N_26897,N_26116,N_25910);
nor U26898 (N_26898,N_25982,N_26212);
nor U26899 (N_26899,N_26320,N_26140);
xor U26900 (N_26900,N_25814,N_26299);
xor U26901 (N_26901,N_26156,N_25813);
nor U26902 (N_26902,N_26319,N_26134);
xnor U26903 (N_26903,N_25880,N_26340);
nand U26904 (N_26904,N_26044,N_26293);
nand U26905 (N_26905,N_26292,N_26200);
or U26906 (N_26906,N_26053,N_26077);
or U26907 (N_26907,N_25890,N_26292);
and U26908 (N_26908,N_26063,N_26020);
nand U26909 (N_26909,N_26168,N_26045);
and U26910 (N_26910,N_26360,N_25942);
nand U26911 (N_26911,N_26142,N_26306);
nor U26912 (N_26912,N_25803,N_26027);
and U26913 (N_26913,N_26342,N_25944);
and U26914 (N_26914,N_25887,N_26218);
nor U26915 (N_26915,N_26075,N_25892);
nor U26916 (N_26916,N_26005,N_26306);
nor U26917 (N_26917,N_26050,N_26226);
xor U26918 (N_26918,N_26155,N_26267);
nand U26919 (N_26919,N_26298,N_26136);
and U26920 (N_26920,N_26335,N_26290);
or U26921 (N_26921,N_26214,N_26138);
or U26922 (N_26922,N_26286,N_26004);
or U26923 (N_26923,N_26043,N_25851);
xor U26924 (N_26924,N_25983,N_26213);
and U26925 (N_26925,N_26198,N_25916);
nand U26926 (N_26926,N_26131,N_25929);
or U26927 (N_26927,N_26137,N_26348);
and U26928 (N_26928,N_26335,N_26190);
or U26929 (N_26929,N_26180,N_26375);
or U26930 (N_26930,N_26375,N_25981);
or U26931 (N_26931,N_25991,N_25837);
xor U26932 (N_26932,N_25871,N_26035);
and U26933 (N_26933,N_26050,N_26204);
and U26934 (N_26934,N_25842,N_26292);
nor U26935 (N_26935,N_26246,N_26022);
or U26936 (N_26936,N_25867,N_25841);
or U26937 (N_26937,N_26178,N_26359);
or U26938 (N_26938,N_26015,N_25805);
or U26939 (N_26939,N_26064,N_26088);
nand U26940 (N_26940,N_25895,N_25857);
or U26941 (N_26941,N_26365,N_25820);
or U26942 (N_26942,N_26147,N_26310);
xor U26943 (N_26943,N_25884,N_25969);
nor U26944 (N_26944,N_25990,N_25833);
nor U26945 (N_26945,N_26381,N_26229);
or U26946 (N_26946,N_26340,N_26321);
and U26947 (N_26947,N_26081,N_26015);
xnor U26948 (N_26948,N_26117,N_25993);
nor U26949 (N_26949,N_25926,N_26219);
and U26950 (N_26950,N_26395,N_25919);
or U26951 (N_26951,N_25969,N_26221);
nor U26952 (N_26952,N_26399,N_25951);
nor U26953 (N_26953,N_26170,N_26120);
or U26954 (N_26954,N_26192,N_26126);
nor U26955 (N_26955,N_26110,N_26397);
or U26956 (N_26956,N_26353,N_25976);
and U26957 (N_26957,N_26249,N_26137);
nor U26958 (N_26958,N_26117,N_26278);
xnor U26959 (N_26959,N_26380,N_26187);
nand U26960 (N_26960,N_26123,N_26271);
xnor U26961 (N_26961,N_26355,N_25863);
or U26962 (N_26962,N_26092,N_26168);
nor U26963 (N_26963,N_26328,N_26121);
nor U26964 (N_26964,N_26093,N_26295);
xnor U26965 (N_26965,N_26391,N_26248);
nor U26966 (N_26966,N_25994,N_26311);
and U26967 (N_26967,N_25940,N_26119);
nor U26968 (N_26968,N_25969,N_26195);
nor U26969 (N_26969,N_26161,N_26223);
nand U26970 (N_26970,N_26178,N_26028);
xor U26971 (N_26971,N_25925,N_26144);
and U26972 (N_26972,N_26199,N_26061);
nand U26973 (N_26973,N_25963,N_26005);
nor U26974 (N_26974,N_26149,N_26130);
or U26975 (N_26975,N_26384,N_26072);
nor U26976 (N_26976,N_26076,N_26114);
and U26977 (N_26977,N_25991,N_26194);
nand U26978 (N_26978,N_25867,N_26385);
or U26979 (N_26979,N_26278,N_26235);
xnor U26980 (N_26980,N_26399,N_26087);
and U26981 (N_26981,N_25926,N_26321);
nor U26982 (N_26982,N_25955,N_26018);
and U26983 (N_26983,N_26206,N_25884);
or U26984 (N_26984,N_25989,N_25968);
or U26985 (N_26985,N_26306,N_25941);
xor U26986 (N_26986,N_25978,N_26231);
nor U26987 (N_26987,N_26319,N_26077);
xor U26988 (N_26988,N_25940,N_26096);
and U26989 (N_26989,N_26224,N_26313);
xor U26990 (N_26990,N_25989,N_25942);
or U26991 (N_26991,N_26159,N_25815);
nor U26992 (N_26992,N_26091,N_25862);
nand U26993 (N_26993,N_26199,N_25987);
xnor U26994 (N_26994,N_25827,N_26242);
nor U26995 (N_26995,N_26011,N_25906);
nand U26996 (N_26996,N_25944,N_25930);
or U26997 (N_26997,N_26032,N_26352);
nor U26998 (N_26998,N_26352,N_25924);
nand U26999 (N_26999,N_25989,N_25963);
and U27000 (N_27000,N_26924,N_26414);
or U27001 (N_27001,N_26996,N_26491);
xnor U27002 (N_27002,N_26881,N_26547);
nor U27003 (N_27003,N_26577,N_26821);
xor U27004 (N_27004,N_26570,N_26668);
or U27005 (N_27005,N_26463,N_26890);
nor U27006 (N_27006,N_26887,N_26681);
nor U27007 (N_27007,N_26567,N_26932);
nor U27008 (N_27008,N_26593,N_26427);
nor U27009 (N_27009,N_26471,N_26473);
nor U27010 (N_27010,N_26696,N_26861);
nand U27011 (N_27011,N_26852,N_26559);
or U27012 (N_27012,N_26906,N_26889);
nand U27013 (N_27013,N_26413,N_26512);
or U27014 (N_27014,N_26978,N_26905);
nand U27015 (N_27015,N_26498,N_26937);
nand U27016 (N_27016,N_26594,N_26921);
xnor U27017 (N_27017,N_26869,N_26481);
xnor U27018 (N_27018,N_26453,N_26475);
xor U27019 (N_27019,N_26597,N_26408);
and U27020 (N_27020,N_26918,N_26812);
xnor U27021 (N_27021,N_26666,N_26785);
xnor U27022 (N_27022,N_26566,N_26802);
and U27023 (N_27023,N_26831,N_26535);
nand U27024 (N_27024,N_26472,N_26857);
and U27025 (N_27025,N_26579,N_26718);
xor U27026 (N_27026,N_26879,N_26914);
nor U27027 (N_27027,N_26662,N_26588);
or U27028 (N_27028,N_26529,N_26706);
nand U27029 (N_27029,N_26965,N_26883);
nand U27030 (N_27030,N_26532,N_26817);
nor U27031 (N_27031,N_26929,N_26515);
nand U27032 (N_27032,N_26652,N_26572);
nor U27033 (N_27033,N_26739,N_26563);
and U27034 (N_27034,N_26781,N_26493);
or U27035 (N_27035,N_26651,N_26749);
xnor U27036 (N_27036,N_26665,N_26780);
and U27037 (N_27037,N_26990,N_26659);
xor U27038 (N_27038,N_26561,N_26900);
nor U27039 (N_27039,N_26891,N_26528);
and U27040 (N_27040,N_26671,N_26683);
xor U27041 (N_27041,N_26590,N_26946);
xor U27042 (N_27042,N_26587,N_26745);
xor U27043 (N_27043,N_26620,N_26851);
and U27044 (N_27044,N_26727,N_26959);
or U27045 (N_27045,N_26439,N_26970);
xor U27046 (N_27046,N_26949,N_26508);
and U27047 (N_27047,N_26462,N_26539);
or U27048 (N_27048,N_26574,N_26947);
xnor U27049 (N_27049,N_26777,N_26797);
xnor U27050 (N_27050,N_26656,N_26488);
nand U27051 (N_27051,N_26614,N_26627);
and U27052 (N_27052,N_26884,N_26950);
or U27053 (N_27053,N_26499,N_26839);
or U27054 (N_27054,N_26615,N_26700);
or U27055 (N_27055,N_26728,N_26420);
and U27056 (N_27056,N_26913,N_26447);
nor U27057 (N_27057,N_26873,N_26582);
nor U27058 (N_27058,N_26800,N_26938);
nor U27059 (N_27059,N_26448,N_26854);
nand U27060 (N_27060,N_26935,N_26557);
nor U27061 (N_27061,N_26772,N_26476);
nand U27062 (N_27062,N_26536,N_26417);
or U27063 (N_27063,N_26554,N_26892);
xor U27064 (N_27064,N_26541,N_26510);
or U27065 (N_27065,N_26433,N_26810);
or U27066 (N_27066,N_26858,N_26443);
nor U27067 (N_27067,N_26863,N_26859);
nor U27068 (N_27068,N_26964,N_26560);
or U27069 (N_27069,N_26993,N_26490);
nand U27070 (N_27070,N_26682,N_26699);
and U27071 (N_27071,N_26865,N_26633);
xnor U27072 (N_27072,N_26667,N_26416);
or U27073 (N_27073,N_26621,N_26595);
or U27074 (N_27074,N_26792,N_26422);
nand U27075 (N_27075,N_26804,N_26544);
and U27076 (N_27076,N_26632,N_26530);
and U27077 (N_27077,N_26465,N_26717);
and U27078 (N_27078,N_26680,N_26432);
xnor U27079 (N_27079,N_26603,N_26919);
xnor U27080 (N_27080,N_26992,N_26838);
or U27081 (N_27081,N_26872,N_26917);
nand U27082 (N_27082,N_26705,N_26407);
nand U27083 (N_27083,N_26446,N_26436);
xor U27084 (N_27084,N_26725,N_26737);
or U27085 (N_27085,N_26972,N_26822);
nand U27086 (N_27086,N_26923,N_26989);
and U27087 (N_27087,N_26786,N_26457);
and U27088 (N_27088,N_26591,N_26653);
xnor U27089 (N_27089,N_26486,N_26634);
nand U27090 (N_27090,N_26966,N_26648);
nor U27091 (N_27091,N_26719,N_26550);
or U27092 (N_27092,N_26760,N_26789);
or U27093 (N_27093,N_26675,N_26808);
nand U27094 (N_27094,N_26679,N_26776);
xnor U27095 (N_27095,N_26755,N_26870);
xor U27096 (N_27096,N_26685,N_26741);
xor U27097 (N_27097,N_26751,N_26956);
and U27098 (N_27098,N_26431,N_26916);
nand U27099 (N_27099,N_26610,N_26429);
or U27100 (N_27100,N_26456,N_26411);
xor U27101 (N_27101,N_26543,N_26548);
nor U27102 (N_27102,N_26692,N_26955);
nor U27103 (N_27103,N_26895,N_26624);
and U27104 (N_27104,N_26423,N_26807);
nand U27105 (N_27105,N_26787,N_26801);
xor U27106 (N_27106,N_26455,N_26762);
xor U27107 (N_27107,N_26445,N_26437);
xnor U27108 (N_27108,N_26690,N_26885);
and U27109 (N_27109,N_26805,N_26520);
and U27110 (N_27110,N_26622,N_26503);
nor U27111 (N_27111,N_26980,N_26672);
nand U27112 (N_27112,N_26747,N_26971);
xnor U27113 (N_27113,N_26649,N_26819);
xor U27114 (N_27114,N_26864,N_26589);
or U27115 (N_27115,N_26984,N_26825);
nand U27116 (N_27116,N_26688,N_26855);
or U27117 (N_27117,N_26898,N_26596);
nor U27118 (N_27118,N_26833,N_26744);
xor U27119 (N_27119,N_26722,N_26948);
xor U27120 (N_27120,N_26968,N_26623);
xor U27121 (N_27121,N_26421,N_26791);
nand U27122 (N_27122,N_26911,N_26927);
nand U27123 (N_27123,N_26874,N_26977);
nand U27124 (N_27124,N_26998,N_26640);
and U27125 (N_27125,N_26779,N_26832);
or U27126 (N_27126,N_26714,N_26523);
nand U27127 (N_27127,N_26729,N_26979);
and U27128 (N_27128,N_26910,N_26827);
xor U27129 (N_27129,N_26886,N_26504);
or U27130 (N_27130,N_26495,N_26551);
nand U27131 (N_27131,N_26403,N_26641);
nand U27132 (N_27132,N_26840,N_26545);
and U27133 (N_27133,N_26412,N_26466);
nor U27134 (N_27134,N_26794,N_26790);
nor U27135 (N_27135,N_26643,N_26754);
xnor U27136 (N_27136,N_26555,N_26829);
and U27137 (N_27137,N_26487,N_26987);
nor U27138 (N_27138,N_26928,N_26568);
nor U27139 (N_27139,N_26584,N_26846);
nor U27140 (N_27140,N_26516,N_26771);
nor U27141 (N_27141,N_26761,N_26880);
nand U27142 (N_27142,N_26406,N_26664);
nor U27143 (N_27143,N_26454,N_26740);
nand U27144 (N_27144,N_26766,N_26876);
nand U27145 (N_27145,N_26995,N_26769);
and U27146 (N_27146,N_26517,N_26438);
or U27147 (N_27147,N_26999,N_26957);
xor U27148 (N_27148,N_26811,N_26856);
and U27149 (N_27149,N_26799,N_26502);
nand U27150 (N_27150,N_26960,N_26449);
and U27151 (N_27151,N_26850,N_26575);
nand U27152 (N_27152,N_26875,N_26991);
or U27153 (N_27153,N_26894,N_26708);
or U27154 (N_27154,N_26518,N_26470);
or U27155 (N_27155,N_26496,N_26592);
xor U27156 (N_27156,N_26904,N_26757);
and U27157 (N_27157,N_26556,N_26997);
xnor U27158 (N_27158,N_26730,N_26616);
nor U27159 (N_27159,N_26451,N_26841);
nand U27160 (N_27160,N_26480,N_26670);
nand U27161 (N_27161,N_26585,N_26501);
and U27162 (N_27162,N_26424,N_26908);
and U27163 (N_27163,N_26763,N_26669);
and U27164 (N_27164,N_26742,N_26639);
nand U27165 (N_27165,N_26720,N_26707);
or U27166 (N_27166,N_26691,N_26571);
and U27167 (N_27167,N_26882,N_26695);
and U27168 (N_27168,N_26638,N_26715);
nor U27169 (N_27169,N_26697,N_26409);
xnor U27170 (N_27170,N_26626,N_26724);
or U27171 (N_27171,N_26494,N_26617);
nor U27172 (N_27172,N_26569,N_26922);
xnor U27173 (N_27173,N_26866,N_26435);
and U27174 (N_27174,N_26542,N_26525);
nor U27175 (N_27175,N_26468,N_26844);
xor U27176 (N_27176,N_26767,N_26847);
xnor U27177 (N_27177,N_26778,N_26458);
and U27178 (N_27178,N_26853,N_26482);
xor U27179 (N_27179,N_26830,N_26743);
xor U27180 (N_27180,N_26425,N_26673);
or U27181 (N_27181,N_26644,N_26818);
and U27182 (N_27182,N_26986,N_26686);
or U27183 (N_27183,N_26565,N_26553);
nor U27184 (N_27184,N_26636,N_26952);
and U27185 (N_27185,N_26934,N_26521);
xor U27186 (N_27186,N_26912,N_26444);
and U27187 (N_27187,N_26676,N_26862);
nor U27188 (N_27188,N_26401,N_26721);
nand U27189 (N_27189,N_26513,N_26835);
nand U27190 (N_27190,N_26578,N_26461);
and U27191 (N_27191,N_26460,N_26759);
xor U27192 (N_27192,N_26732,N_26868);
or U27193 (N_27193,N_26902,N_26689);
xnor U27194 (N_27194,N_26606,N_26712);
nor U27195 (N_27195,N_26897,N_26783);
or U27196 (N_27196,N_26635,N_26843);
or U27197 (N_27197,N_26576,N_26793);
or U27198 (N_27198,N_26752,N_26940);
and U27199 (N_27199,N_26511,N_26803);
nor U27200 (N_27200,N_26974,N_26925);
or U27201 (N_27201,N_26824,N_26798);
and U27202 (N_27202,N_26611,N_26598);
nand U27203 (N_27203,N_26507,N_26430);
xor U27204 (N_27204,N_26726,N_26684);
xor U27205 (N_27205,N_26573,N_26519);
and U27206 (N_27206,N_26537,N_26526);
nand U27207 (N_27207,N_26764,N_26711);
nor U27208 (N_27208,N_26506,N_26848);
and U27209 (N_27209,N_26618,N_26703);
or U27210 (N_27210,N_26936,N_26775);
or U27211 (N_27211,N_26975,N_26450);
and U27212 (N_27212,N_26784,N_26531);
nand U27213 (N_27213,N_26985,N_26586);
nand U27214 (N_27214,N_26926,N_26753);
nor U27215 (N_27215,N_26694,N_26467);
xnor U27216 (N_27216,N_26888,N_26645);
nand U27217 (N_27217,N_26723,N_26602);
xnor U27218 (N_27218,N_26702,N_26909);
xnor U27219 (N_27219,N_26806,N_26893);
or U27220 (N_27220,N_26629,N_26509);
nand U27221 (N_27221,N_26750,N_26698);
nor U27222 (N_27222,N_26674,N_26538);
xnor U27223 (N_27223,N_26628,N_26534);
xor U27224 (N_27224,N_26533,N_26736);
xor U27225 (N_27225,N_26410,N_26601);
or U27226 (N_27226,N_26583,N_26903);
nand U27227 (N_27227,N_26600,N_26637);
and U27228 (N_27228,N_26828,N_26654);
or U27229 (N_27229,N_26484,N_26522);
nand U27230 (N_27230,N_26663,N_26404);
nor U27231 (N_27231,N_26489,N_26580);
and U27232 (N_27232,N_26815,N_26963);
or U27233 (N_27233,N_26546,N_26469);
nand U27234 (N_27234,N_26713,N_26479);
xor U27235 (N_27235,N_26564,N_26660);
nand U27236 (N_27236,N_26746,N_26655);
nand U27237 (N_27237,N_26930,N_26607);
nand U27238 (N_27238,N_26939,N_26434);
nand U27239 (N_27239,N_26619,N_26581);
nand U27240 (N_27240,N_26505,N_26796);
nor U27241 (N_27241,N_26400,N_26836);
and U27242 (N_27242,N_26871,N_26524);
or U27243 (N_27243,N_26734,N_26452);
nand U27244 (N_27244,N_26402,N_26849);
or U27245 (N_27245,N_26405,N_26677);
nand U27246 (N_27246,N_26733,N_26773);
xnor U27247 (N_27247,N_26562,N_26931);
and U27248 (N_27248,N_26500,N_26958);
xor U27249 (N_27249,N_26768,N_26613);
nor U27250 (N_27250,N_26704,N_26945);
xor U27251 (N_27251,N_26599,N_26497);
nand U27252 (N_27252,N_26549,N_26442);
and U27253 (N_27253,N_26933,N_26969);
and U27254 (N_27254,N_26944,N_26428);
nand U27255 (N_27255,N_26492,N_26826);
nor U27256 (N_27256,N_26441,N_26459);
and U27257 (N_27257,N_26514,N_26657);
and U27258 (N_27258,N_26967,N_26820);
and U27259 (N_27259,N_26687,N_26474);
nor U27260 (N_27260,N_26774,N_26605);
nor U27261 (N_27261,N_26953,N_26878);
nor U27262 (N_27262,N_26941,N_26612);
and U27263 (N_27263,N_26642,N_26899);
and U27264 (N_27264,N_26609,N_26860);
and U27265 (N_27265,N_26415,N_26478);
nor U27266 (N_27266,N_26795,N_26758);
or U27267 (N_27267,N_26558,N_26814);
nor U27268 (N_27268,N_26658,N_26962);
or U27269 (N_27269,N_26994,N_26661);
or U27270 (N_27270,N_26527,N_26625);
and U27271 (N_27271,N_26765,N_26982);
and U27272 (N_27272,N_26419,N_26901);
or U27273 (N_27273,N_26896,N_26716);
nand U27274 (N_27274,N_26630,N_26748);
or U27275 (N_27275,N_26477,N_26920);
nand U27276 (N_27276,N_26915,N_26943);
nor U27277 (N_27277,N_26464,N_26954);
and U27278 (N_27278,N_26735,N_26842);
nand U27279 (N_27279,N_26710,N_26709);
and U27280 (N_27280,N_26770,N_26782);
and U27281 (N_27281,N_26845,N_26961);
nand U27282 (N_27282,N_26823,N_26942);
nand U27283 (N_27283,N_26426,N_26983);
xnor U27284 (N_27284,N_26973,N_26907);
nor U27285 (N_27285,N_26976,N_26604);
nor U27286 (N_27286,N_26867,N_26646);
nor U27287 (N_27287,N_26988,N_26738);
nand U27288 (N_27288,N_26552,N_26816);
and U27289 (N_27289,N_26834,N_26540);
or U27290 (N_27290,N_26418,N_26631);
xor U27291 (N_27291,N_26809,N_26837);
and U27292 (N_27292,N_26788,N_26756);
xnor U27293 (N_27293,N_26483,N_26877);
nor U27294 (N_27294,N_26650,N_26647);
and U27295 (N_27295,N_26678,N_26951);
or U27296 (N_27296,N_26981,N_26701);
and U27297 (N_27297,N_26731,N_26693);
nor U27298 (N_27298,N_26608,N_26813);
nor U27299 (N_27299,N_26485,N_26440);
xnor U27300 (N_27300,N_26650,N_26976);
nor U27301 (N_27301,N_26813,N_26503);
nor U27302 (N_27302,N_26965,N_26782);
and U27303 (N_27303,N_26950,N_26664);
nor U27304 (N_27304,N_26569,N_26671);
nor U27305 (N_27305,N_26778,N_26466);
nand U27306 (N_27306,N_26511,N_26827);
nand U27307 (N_27307,N_26649,N_26811);
xor U27308 (N_27308,N_26949,N_26515);
xor U27309 (N_27309,N_26601,N_26451);
xnor U27310 (N_27310,N_26565,N_26809);
nor U27311 (N_27311,N_26583,N_26500);
nor U27312 (N_27312,N_26989,N_26785);
or U27313 (N_27313,N_26577,N_26493);
or U27314 (N_27314,N_26646,N_26471);
and U27315 (N_27315,N_26446,N_26455);
and U27316 (N_27316,N_26565,N_26513);
or U27317 (N_27317,N_26783,N_26680);
or U27318 (N_27318,N_26518,N_26627);
xor U27319 (N_27319,N_26777,N_26539);
nor U27320 (N_27320,N_26631,N_26588);
or U27321 (N_27321,N_26750,N_26843);
or U27322 (N_27322,N_26677,N_26971);
xor U27323 (N_27323,N_26513,N_26844);
nand U27324 (N_27324,N_26913,N_26551);
nand U27325 (N_27325,N_26935,N_26907);
or U27326 (N_27326,N_26658,N_26726);
and U27327 (N_27327,N_26443,N_26881);
nor U27328 (N_27328,N_26879,N_26555);
nand U27329 (N_27329,N_26430,N_26735);
or U27330 (N_27330,N_26680,N_26450);
nand U27331 (N_27331,N_26567,N_26727);
and U27332 (N_27332,N_26784,N_26543);
nand U27333 (N_27333,N_26619,N_26764);
nor U27334 (N_27334,N_26459,N_26727);
and U27335 (N_27335,N_26929,N_26879);
or U27336 (N_27336,N_26763,N_26526);
xnor U27337 (N_27337,N_26745,N_26617);
and U27338 (N_27338,N_26500,N_26938);
nor U27339 (N_27339,N_26439,N_26598);
nand U27340 (N_27340,N_26766,N_26811);
nand U27341 (N_27341,N_26624,N_26556);
xor U27342 (N_27342,N_26469,N_26639);
or U27343 (N_27343,N_26484,N_26609);
and U27344 (N_27344,N_26875,N_26665);
or U27345 (N_27345,N_26418,N_26835);
nor U27346 (N_27346,N_26517,N_26956);
xnor U27347 (N_27347,N_26634,N_26874);
nor U27348 (N_27348,N_26428,N_26673);
and U27349 (N_27349,N_26890,N_26830);
or U27350 (N_27350,N_26537,N_26543);
nand U27351 (N_27351,N_26567,N_26454);
nor U27352 (N_27352,N_26438,N_26511);
nor U27353 (N_27353,N_26747,N_26699);
and U27354 (N_27354,N_26446,N_26422);
nand U27355 (N_27355,N_26639,N_26999);
and U27356 (N_27356,N_26808,N_26604);
xor U27357 (N_27357,N_26453,N_26829);
xor U27358 (N_27358,N_26750,N_26581);
xnor U27359 (N_27359,N_26421,N_26653);
xnor U27360 (N_27360,N_26853,N_26526);
or U27361 (N_27361,N_26951,N_26746);
nand U27362 (N_27362,N_26799,N_26881);
and U27363 (N_27363,N_26666,N_26833);
or U27364 (N_27364,N_26542,N_26789);
and U27365 (N_27365,N_26916,N_26855);
nand U27366 (N_27366,N_26494,N_26414);
xor U27367 (N_27367,N_26485,N_26703);
and U27368 (N_27368,N_26799,N_26820);
and U27369 (N_27369,N_26770,N_26456);
or U27370 (N_27370,N_26707,N_26846);
nand U27371 (N_27371,N_26871,N_26737);
xnor U27372 (N_27372,N_26990,N_26466);
or U27373 (N_27373,N_26425,N_26712);
and U27374 (N_27374,N_26722,N_26713);
xor U27375 (N_27375,N_26626,N_26515);
xor U27376 (N_27376,N_26799,N_26526);
nor U27377 (N_27377,N_26745,N_26601);
nor U27378 (N_27378,N_26814,N_26720);
nand U27379 (N_27379,N_26967,N_26523);
or U27380 (N_27380,N_26573,N_26892);
or U27381 (N_27381,N_26856,N_26701);
xor U27382 (N_27382,N_26923,N_26771);
nor U27383 (N_27383,N_26929,N_26721);
nor U27384 (N_27384,N_26967,N_26516);
nand U27385 (N_27385,N_26615,N_26786);
and U27386 (N_27386,N_26707,N_26664);
xor U27387 (N_27387,N_26855,N_26489);
nand U27388 (N_27388,N_26861,N_26921);
nor U27389 (N_27389,N_26505,N_26434);
or U27390 (N_27390,N_26406,N_26464);
nand U27391 (N_27391,N_26714,N_26823);
xor U27392 (N_27392,N_26602,N_26920);
xor U27393 (N_27393,N_26677,N_26562);
and U27394 (N_27394,N_26841,N_26737);
xnor U27395 (N_27395,N_26442,N_26565);
and U27396 (N_27396,N_26439,N_26878);
nor U27397 (N_27397,N_26696,N_26422);
nand U27398 (N_27398,N_26549,N_26674);
and U27399 (N_27399,N_26518,N_26752);
xnor U27400 (N_27400,N_26940,N_26965);
nor U27401 (N_27401,N_26573,N_26485);
and U27402 (N_27402,N_26415,N_26564);
nor U27403 (N_27403,N_26926,N_26400);
nor U27404 (N_27404,N_26478,N_26708);
xnor U27405 (N_27405,N_26550,N_26406);
nor U27406 (N_27406,N_26424,N_26632);
and U27407 (N_27407,N_26481,N_26688);
and U27408 (N_27408,N_26411,N_26434);
nor U27409 (N_27409,N_26419,N_26622);
and U27410 (N_27410,N_26575,N_26979);
and U27411 (N_27411,N_26410,N_26416);
nand U27412 (N_27412,N_26782,N_26452);
nor U27413 (N_27413,N_26832,N_26600);
and U27414 (N_27414,N_26620,N_26568);
nor U27415 (N_27415,N_26842,N_26881);
and U27416 (N_27416,N_26545,N_26570);
xnor U27417 (N_27417,N_26772,N_26468);
or U27418 (N_27418,N_26458,N_26841);
nand U27419 (N_27419,N_26906,N_26753);
xor U27420 (N_27420,N_26929,N_26766);
nand U27421 (N_27421,N_26939,N_26497);
and U27422 (N_27422,N_26525,N_26663);
and U27423 (N_27423,N_26958,N_26722);
nand U27424 (N_27424,N_26885,N_26752);
xor U27425 (N_27425,N_26813,N_26477);
nand U27426 (N_27426,N_26998,N_26409);
or U27427 (N_27427,N_26741,N_26505);
nor U27428 (N_27428,N_26761,N_26771);
xnor U27429 (N_27429,N_26555,N_26989);
or U27430 (N_27430,N_26994,N_26738);
xor U27431 (N_27431,N_26648,N_26996);
xor U27432 (N_27432,N_26433,N_26807);
nand U27433 (N_27433,N_26466,N_26482);
and U27434 (N_27434,N_26811,N_26608);
nand U27435 (N_27435,N_26551,N_26505);
nand U27436 (N_27436,N_26981,N_26469);
nand U27437 (N_27437,N_26969,N_26762);
nor U27438 (N_27438,N_26604,N_26446);
and U27439 (N_27439,N_26771,N_26401);
xor U27440 (N_27440,N_26772,N_26424);
nor U27441 (N_27441,N_26754,N_26589);
xnor U27442 (N_27442,N_26846,N_26662);
nor U27443 (N_27443,N_26611,N_26961);
nor U27444 (N_27444,N_26614,N_26548);
and U27445 (N_27445,N_26483,N_26461);
and U27446 (N_27446,N_26916,N_26648);
or U27447 (N_27447,N_26974,N_26668);
nor U27448 (N_27448,N_26847,N_26811);
nand U27449 (N_27449,N_26825,N_26712);
xnor U27450 (N_27450,N_26574,N_26447);
or U27451 (N_27451,N_26606,N_26895);
nor U27452 (N_27452,N_26544,N_26673);
nor U27453 (N_27453,N_26698,N_26974);
nor U27454 (N_27454,N_26750,N_26527);
nor U27455 (N_27455,N_26649,N_26603);
and U27456 (N_27456,N_26517,N_26699);
nor U27457 (N_27457,N_26669,N_26655);
xnor U27458 (N_27458,N_26945,N_26953);
nand U27459 (N_27459,N_26702,N_26405);
nor U27460 (N_27460,N_26505,N_26746);
and U27461 (N_27461,N_26897,N_26923);
nand U27462 (N_27462,N_26909,N_26731);
nand U27463 (N_27463,N_26766,N_26545);
nand U27464 (N_27464,N_26823,N_26635);
or U27465 (N_27465,N_26580,N_26409);
or U27466 (N_27466,N_26980,N_26650);
nand U27467 (N_27467,N_26860,N_26537);
or U27468 (N_27468,N_26774,N_26807);
xor U27469 (N_27469,N_26986,N_26592);
and U27470 (N_27470,N_26652,N_26772);
nand U27471 (N_27471,N_26517,N_26511);
or U27472 (N_27472,N_26581,N_26762);
and U27473 (N_27473,N_26617,N_26766);
nor U27474 (N_27474,N_26967,N_26615);
nand U27475 (N_27475,N_26425,N_26686);
or U27476 (N_27476,N_26927,N_26925);
and U27477 (N_27477,N_26637,N_26481);
nand U27478 (N_27478,N_26476,N_26844);
nor U27479 (N_27479,N_26900,N_26954);
nor U27480 (N_27480,N_26798,N_26862);
or U27481 (N_27481,N_26859,N_26624);
xnor U27482 (N_27482,N_26602,N_26959);
nand U27483 (N_27483,N_26997,N_26982);
xor U27484 (N_27484,N_26915,N_26871);
nand U27485 (N_27485,N_26712,N_26940);
nand U27486 (N_27486,N_26985,N_26465);
nor U27487 (N_27487,N_26806,N_26530);
xnor U27488 (N_27488,N_26834,N_26622);
nand U27489 (N_27489,N_26841,N_26860);
nand U27490 (N_27490,N_26949,N_26903);
xor U27491 (N_27491,N_26850,N_26820);
and U27492 (N_27492,N_26718,N_26414);
or U27493 (N_27493,N_26944,N_26668);
nor U27494 (N_27494,N_26610,N_26495);
and U27495 (N_27495,N_26956,N_26737);
or U27496 (N_27496,N_26512,N_26809);
nand U27497 (N_27497,N_26479,N_26922);
nor U27498 (N_27498,N_26488,N_26846);
or U27499 (N_27499,N_26972,N_26431);
nand U27500 (N_27500,N_26946,N_26899);
xnor U27501 (N_27501,N_26840,N_26929);
xnor U27502 (N_27502,N_26980,N_26589);
or U27503 (N_27503,N_26450,N_26907);
or U27504 (N_27504,N_26865,N_26742);
nor U27505 (N_27505,N_26907,N_26900);
and U27506 (N_27506,N_26993,N_26531);
nand U27507 (N_27507,N_26563,N_26423);
xor U27508 (N_27508,N_26969,N_26991);
nor U27509 (N_27509,N_26596,N_26670);
nor U27510 (N_27510,N_26733,N_26623);
nor U27511 (N_27511,N_26530,N_26412);
nor U27512 (N_27512,N_26463,N_26501);
xor U27513 (N_27513,N_26490,N_26611);
nand U27514 (N_27514,N_26748,N_26491);
and U27515 (N_27515,N_26992,N_26866);
nor U27516 (N_27516,N_26666,N_26904);
xor U27517 (N_27517,N_26474,N_26423);
nor U27518 (N_27518,N_26788,N_26950);
or U27519 (N_27519,N_26996,N_26577);
nand U27520 (N_27520,N_26783,N_26559);
nor U27521 (N_27521,N_26451,N_26892);
nor U27522 (N_27522,N_26868,N_26910);
nor U27523 (N_27523,N_26439,N_26505);
or U27524 (N_27524,N_26782,N_26516);
xnor U27525 (N_27525,N_26811,N_26596);
nor U27526 (N_27526,N_26966,N_26827);
nand U27527 (N_27527,N_26906,N_26631);
and U27528 (N_27528,N_26545,N_26554);
or U27529 (N_27529,N_26435,N_26618);
and U27530 (N_27530,N_26476,N_26880);
nand U27531 (N_27531,N_26736,N_26552);
and U27532 (N_27532,N_26939,N_26961);
and U27533 (N_27533,N_26790,N_26893);
and U27534 (N_27534,N_26477,N_26544);
and U27535 (N_27535,N_26453,N_26607);
nor U27536 (N_27536,N_26645,N_26959);
xnor U27537 (N_27537,N_26671,N_26721);
nand U27538 (N_27538,N_26593,N_26990);
nand U27539 (N_27539,N_26576,N_26486);
nand U27540 (N_27540,N_26796,N_26608);
or U27541 (N_27541,N_26421,N_26565);
and U27542 (N_27542,N_26452,N_26722);
nor U27543 (N_27543,N_26527,N_26773);
nor U27544 (N_27544,N_26773,N_26413);
nand U27545 (N_27545,N_26401,N_26973);
and U27546 (N_27546,N_26575,N_26660);
or U27547 (N_27547,N_26425,N_26792);
xor U27548 (N_27548,N_26407,N_26444);
or U27549 (N_27549,N_26923,N_26676);
and U27550 (N_27550,N_26922,N_26862);
and U27551 (N_27551,N_26943,N_26490);
nor U27552 (N_27552,N_26687,N_26802);
or U27553 (N_27553,N_26711,N_26600);
or U27554 (N_27554,N_26811,N_26537);
xnor U27555 (N_27555,N_26954,N_26460);
xnor U27556 (N_27556,N_26623,N_26774);
nand U27557 (N_27557,N_26890,N_26785);
or U27558 (N_27558,N_26887,N_26954);
and U27559 (N_27559,N_26588,N_26645);
nor U27560 (N_27560,N_26981,N_26413);
nand U27561 (N_27561,N_26848,N_26413);
nor U27562 (N_27562,N_26758,N_26623);
nor U27563 (N_27563,N_26917,N_26593);
or U27564 (N_27564,N_26406,N_26803);
and U27565 (N_27565,N_26978,N_26960);
and U27566 (N_27566,N_26857,N_26705);
nor U27567 (N_27567,N_26431,N_26708);
xnor U27568 (N_27568,N_26757,N_26625);
and U27569 (N_27569,N_26478,N_26432);
nand U27570 (N_27570,N_26962,N_26421);
or U27571 (N_27571,N_26472,N_26869);
and U27572 (N_27572,N_26669,N_26890);
or U27573 (N_27573,N_26495,N_26402);
xor U27574 (N_27574,N_26834,N_26418);
nor U27575 (N_27575,N_26708,N_26535);
xor U27576 (N_27576,N_26458,N_26657);
nand U27577 (N_27577,N_26588,N_26660);
nor U27578 (N_27578,N_26810,N_26747);
and U27579 (N_27579,N_26655,N_26458);
or U27580 (N_27580,N_26870,N_26541);
and U27581 (N_27581,N_26809,N_26448);
nand U27582 (N_27582,N_26533,N_26932);
and U27583 (N_27583,N_26515,N_26975);
or U27584 (N_27584,N_26672,N_26785);
nor U27585 (N_27585,N_26815,N_26753);
or U27586 (N_27586,N_26840,N_26921);
or U27587 (N_27587,N_26578,N_26621);
and U27588 (N_27588,N_26821,N_26456);
nor U27589 (N_27589,N_26839,N_26643);
or U27590 (N_27590,N_26675,N_26868);
and U27591 (N_27591,N_26682,N_26470);
nand U27592 (N_27592,N_26659,N_26805);
xnor U27593 (N_27593,N_26687,N_26433);
or U27594 (N_27594,N_26947,N_26880);
nand U27595 (N_27595,N_26561,N_26465);
or U27596 (N_27596,N_26967,N_26527);
xor U27597 (N_27597,N_26541,N_26663);
nand U27598 (N_27598,N_26722,N_26550);
or U27599 (N_27599,N_26564,N_26910);
nand U27600 (N_27600,N_27085,N_27215);
nor U27601 (N_27601,N_27507,N_27343);
and U27602 (N_27602,N_27288,N_27247);
or U27603 (N_27603,N_27303,N_27279);
and U27604 (N_27604,N_27446,N_27023);
and U27605 (N_27605,N_27052,N_27425);
xnor U27606 (N_27606,N_27504,N_27136);
nor U27607 (N_27607,N_27494,N_27436);
nand U27608 (N_27608,N_27244,N_27135);
nor U27609 (N_27609,N_27584,N_27535);
nand U27610 (N_27610,N_27409,N_27368);
and U27611 (N_27611,N_27417,N_27435);
nor U27612 (N_27612,N_27219,N_27223);
xnor U27613 (N_27613,N_27198,N_27291);
xor U27614 (N_27614,N_27466,N_27034);
nand U27615 (N_27615,N_27537,N_27220);
or U27616 (N_27616,N_27360,N_27150);
and U27617 (N_27617,N_27207,N_27108);
xor U27618 (N_27618,N_27339,N_27255);
xor U27619 (N_27619,N_27415,N_27462);
nor U27620 (N_27620,N_27470,N_27277);
nand U27621 (N_27621,N_27497,N_27204);
or U27622 (N_27622,N_27526,N_27329);
nor U27623 (N_27623,N_27389,N_27556);
xor U27624 (N_27624,N_27451,N_27473);
or U27625 (N_27625,N_27027,N_27580);
and U27626 (N_27626,N_27426,N_27089);
nand U27627 (N_27627,N_27463,N_27132);
xor U27628 (N_27628,N_27499,N_27233);
nand U27629 (N_27629,N_27503,N_27016);
xnor U27630 (N_27630,N_27010,N_27289);
nor U27631 (N_27631,N_27159,N_27116);
nand U27632 (N_27632,N_27483,N_27391);
and U27633 (N_27633,N_27599,N_27283);
nor U27634 (N_27634,N_27160,N_27254);
or U27635 (N_27635,N_27053,N_27572);
or U27636 (N_27636,N_27182,N_27505);
or U27637 (N_27637,N_27450,N_27379);
and U27638 (N_27638,N_27138,N_27325);
or U27639 (N_27639,N_27024,N_27530);
nand U27640 (N_27640,N_27000,N_27259);
nand U27641 (N_27641,N_27115,N_27284);
and U27642 (N_27642,N_27544,N_27054);
xnor U27643 (N_27643,N_27165,N_27495);
nor U27644 (N_27644,N_27093,N_27468);
xor U27645 (N_27645,N_27552,N_27441);
xor U27646 (N_27646,N_27057,N_27130);
and U27647 (N_27647,N_27351,N_27532);
nand U27648 (N_27648,N_27529,N_27512);
nor U27649 (N_27649,N_27140,N_27175);
nand U27650 (N_27650,N_27020,N_27107);
nor U27651 (N_27651,N_27217,N_27437);
xor U27652 (N_27652,N_27313,N_27307);
or U27653 (N_27653,N_27066,N_27492);
nor U27654 (N_27654,N_27231,N_27190);
nand U27655 (N_27655,N_27500,N_27056);
and U27656 (N_27656,N_27420,N_27253);
xor U27657 (N_27657,N_27464,N_27591);
xnor U27658 (N_27658,N_27346,N_27364);
and U27659 (N_27659,N_27075,N_27548);
nor U27660 (N_27660,N_27469,N_27498);
nand U27661 (N_27661,N_27311,N_27001);
nand U27662 (N_27662,N_27021,N_27101);
nand U27663 (N_27663,N_27587,N_27092);
xor U27664 (N_27664,N_27597,N_27044);
or U27665 (N_27665,N_27439,N_27332);
nand U27666 (N_27666,N_27251,N_27012);
or U27667 (N_27667,N_27088,N_27145);
and U27668 (N_27668,N_27413,N_27367);
nor U27669 (N_27669,N_27102,N_27402);
or U27670 (N_27670,N_27035,N_27039);
and U27671 (N_27671,N_27594,N_27128);
xor U27672 (N_27672,N_27336,N_27476);
or U27673 (N_27673,N_27058,N_27246);
and U27674 (N_27674,N_27200,N_27296);
nor U27675 (N_27675,N_27265,N_27199);
nand U27676 (N_27676,N_27534,N_27392);
or U27677 (N_27677,N_27163,N_27146);
nor U27678 (N_27678,N_27459,N_27576);
nor U27679 (N_27679,N_27376,N_27008);
and U27680 (N_27680,N_27270,N_27273);
or U27681 (N_27681,N_27352,N_27558);
and U27682 (N_27682,N_27334,N_27046);
or U27683 (N_27683,N_27185,N_27267);
xnor U27684 (N_27684,N_27186,N_27281);
nand U27685 (N_27685,N_27224,N_27388);
nor U27686 (N_27686,N_27210,N_27151);
nand U27687 (N_27687,N_27406,N_27328);
xor U27688 (N_27688,N_27557,N_27348);
nand U27689 (N_27689,N_27427,N_27453);
xor U27690 (N_27690,N_27086,N_27314);
and U27691 (N_27691,N_27033,N_27258);
nand U27692 (N_27692,N_27068,N_27372);
nor U27693 (N_27693,N_27589,N_27161);
nor U27694 (N_27694,N_27117,N_27490);
nand U27695 (N_27695,N_27422,N_27511);
nor U27696 (N_27696,N_27211,N_27479);
and U27697 (N_27697,N_27015,N_27235);
xnor U27698 (N_27698,N_27380,N_27318);
xnor U27699 (N_27699,N_27443,N_27100);
xor U27700 (N_27700,N_27440,N_27410);
nor U27701 (N_27701,N_27004,N_27338);
xnor U27702 (N_27702,N_27104,N_27395);
xor U27703 (N_27703,N_27261,N_27516);
nand U27704 (N_27704,N_27359,N_27598);
and U27705 (N_27705,N_27485,N_27096);
nor U27706 (N_27706,N_27322,N_27149);
xnor U27707 (N_27707,N_27384,N_27448);
nor U27708 (N_27708,N_27375,N_27230);
or U27709 (N_27709,N_27240,N_27205);
and U27710 (N_27710,N_27245,N_27588);
or U27711 (N_27711,N_27278,N_27162);
xor U27712 (N_27712,N_27356,N_27091);
xor U27713 (N_27713,N_27465,N_27310);
and U27714 (N_27714,N_27127,N_27141);
or U27715 (N_27715,N_27358,N_27517);
nor U27716 (N_27716,N_27043,N_27518);
nand U27717 (N_27717,N_27263,N_27103);
xor U27718 (N_27718,N_27378,N_27038);
and U27719 (N_27719,N_27565,N_27069);
nand U27720 (N_27720,N_27579,N_27112);
nand U27721 (N_27721,N_27546,N_27137);
nor U27722 (N_27722,N_27513,N_27166);
nand U27723 (N_27723,N_27386,N_27302);
nand U27724 (N_27724,N_27578,N_27026);
nor U27725 (N_27725,N_27363,N_27369);
xor U27726 (N_27726,N_27194,N_27256);
nor U27727 (N_27727,N_27340,N_27361);
nand U27728 (N_27728,N_27341,N_27113);
or U27729 (N_27729,N_27502,N_27070);
xor U27730 (N_27730,N_27394,N_27218);
xor U27731 (N_27731,N_27337,N_27025);
xor U27732 (N_27732,N_27519,N_27506);
nand U27733 (N_27733,N_27032,N_27125);
xor U27734 (N_27734,N_27124,N_27133);
nor U27735 (N_27735,N_27488,N_27226);
xnor U27736 (N_27736,N_27158,N_27292);
xnor U27737 (N_27737,N_27590,N_27531);
nand U27738 (N_27738,N_27357,N_27569);
xor U27739 (N_27739,N_27030,N_27390);
nor U27740 (N_27740,N_27401,N_27065);
nand U27741 (N_27741,N_27111,N_27174);
nand U27742 (N_27742,N_27275,N_27472);
and U27743 (N_27743,N_27430,N_27084);
or U27744 (N_27744,N_27509,N_27005);
or U27745 (N_27745,N_27126,N_27491);
or U27746 (N_27746,N_27119,N_27407);
nor U27747 (N_27747,N_27383,N_27022);
or U27748 (N_27748,N_27216,N_27154);
and U27749 (N_27749,N_27209,N_27252);
nor U27750 (N_27750,N_27480,N_27041);
nand U27751 (N_27751,N_27201,N_27382);
and U27752 (N_27752,N_27192,N_27449);
nor U27753 (N_27753,N_27482,N_27344);
nand U27754 (N_27754,N_27374,N_27538);
and U27755 (N_27755,N_27342,N_27304);
nand U27756 (N_27756,N_27481,N_27458);
nor U27757 (N_27757,N_27447,N_27345);
xor U27758 (N_27758,N_27076,N_27560);
or U27759 (N_27759,N_27109,N_27434);
xnor U27760 (N_27760,N_27571,N_27110);
and U27761 (N_27761,N_27286,N_27055);
and U27762 (N_27762,N_27444,N_27403);
nor U27763 (N_27763,N_27196,N_27168);
nand U27764 (N_27764,N_27051,N_27202);
nor U27765 (N_27765,N_27316,N_27250);
nor U27766 (N_27766,N_27234,N_27206);
nor U27767 (N_27767,N_27431,N_27272);
nand U27768 (N_27768,N_27399,N_27009);
and U27769 (N_27769,N_27524,N_27408);
nand U27770 (N_27770,N_27129,N_27063);
nor U27771 (N_27771,N_27595,N_27114);
and U27772 (N_27772,N_27049,N_27582);
nor U27773 (N_27773,N_27098,N_27180);
and U27774 (N_27774,N_27048,N_27521);
xnor U27775 (N_27775,N_27370,N_27428);
and U27776 (N_27776,N_27236,N_27148);
nand U27777 (N_27777,N_27164,N_27079);
or U27778 (N_27778,N_27072,N_27551);
nand U27779 (N_27779,N_27295,N_27147);
nor U27780 (N_27780,N_27221,N_27564);
and U27781 (N_27781,N_27282,N_27373);
xnor U27782 (N_27782,N_27404,N_27319);
nor U27783 (N_27783,N_27484,N_27002);
or U27784 (N_27784,N_27522,N_27539);
nor U27785 (N_27785,N_27040,N_27559);
or U27786 (N_27786,N_27242,N_27228);
and U27787 (N_27787,N_27019,N_27268);
and U27788 (N_27788,N_27312,N_27181);
or U27789 (N_27789,N_27131,N_27299);
xor U27790 (N_27790,N_27398,N_27324);
xnor U27791 (N_27791,N_27028,N_27416);
nor U27792 (N_27792,N_27396,N_27433);
or U27793 (N_27793,N_27097,N_27120);
or U27794 (N_27794,N_27156,N_27520);
and U27795 (N_27795,N_27169,N_27018);
and U27796 (N_27796,N_27142,N_27424);
xor U27797 (N_27797,N_27596,N_27570);
nand U27798 (N_27798,N_27387,N_27554);
and U27799 (N_27799,N_27118,N_27347);
or U27800 (N_27800,N_27331,N_27081);
nand U27801 (N_27801,N_27553,N_27561);
nor U27802 (N_27802,N_27155,N_27095);
and U27803 (N_27803,N_27320,N_27438);
and U27804 (N_27804,N_27285,N_27074);
or U27805 (N_27805,N_27349,N_27550);
or U27806 (N_27806,N_27575,N_27173);
or U27807 (N_27807,N_27067,N_27523);
nand U27808 (N_27808,N_27017,N_27188);
nor U27809 (N_27809,N_27400,N_27232);
xnor U27810 (N_27810,N_27460,N_27144);
xnor U27811 (N_27811,N_27029,N_27036);
xor U27812 (N_27812,N_27179,N_27060);
xnor U27813 (N_27813,N_27266,N_27062);
xnor U27814 (N_27814,N_27143,N_27555);
nor U27815 (N_27815,N_27264,N_27461);
nor U27816 (N_27816,N_27045,N_27123);
xor U27817 (N_27817,N_27077,N_27003);
and U27818 (N_27818,N_27195,N_27229);
and U27819 (N_27819,N_27385,N_27064);
nand U27820 (N_27820,N_27157,N_27583);
or U27821 (N_27821,N_27547,N_27031);
nand U27822 (N_27822,N_27477,N_27566);
and U27823 (N_27823,N_27442,N_27193);
or U27824 (N_27824,N_27527,N_27405);
nor U27825 (N_27825,N_27260,N_27269);
xnor U27826 (N_27826,N_27419,N_27414);
xor U27827 (N_27827,N_27421,N_27536);
xor U27828 (N_27828,N_27290,N_27167);
xnor U27829 (N_27829,N_27541,N_27330);
nand U27830 (N_27830,N_27540,N_27457);
nand U27831 (N_27831,N_27397,N_27099);
nor U27832 (N_27832,N_27381,N_27350);
or U27833 (N_27833,N_27214,N_27280);
xor U27834 (N_27834,N_27287,N_27423);
and U27835 (N_27835,N_27317,N_27013);
xor U27836 (N_27836,N_27105,N_27323);
xor U27837 (N_27837,N_27592,N_27208);
and U27838 (N_27838,N_27327,N_27486);
or U27839 (N_27839,N_27455,N_27257);
nand U27840 (N_27840,N_27050,N_27262);
xor U27841 (N_27841,N_27362,N_27071);
nor U27842 (N_27842,N_27326,N_27073);
or U27843 (N_27843,N_27471,N_27212);
xor U27844 (N_27844,N_27335,N_27191);
nand U27845 (N_27845,N_27300,N_27542);
nor U27846 (N_27846,N_27134,N_27082);
and U27847 (N_27847,N_27237,N_27011);
and U27848 (N_27848,N_27309,N_27515);
and U27849 (N_27849,N_27078,N_27189);
nor U27850 (N_27850,N_27543,N_27365);
nor U27851 (N_27851,N_27298,N_27581);
nor U27852 (N_27852,N_27297,N_27249);
xor U27853 (N_27853,N_27042,N_27080);
xor U27854 (N_27854,N_27510,N_27475);
and U27855 (N_27855,N_27377,N_27549);
nand U27856 (N_27856,N_27321,N_27152);
nand U27857 (N_27857,N_27577,N_27176);
nor U27858 (N_27858,N_27306,N_27121);
nand U27859 (N_27859,N_27474,N_27371);
xor U27860 (N_27860,N_27271,N_27178);
xor U27861 (N_27861,N_27445,N_27333);
and U27862 (N_27862,N_27456,N_27187);
xnor U27863 (N_27863,N_27094,N_27037);
xor U27864 (N_27864,N_27454,N_27274);
nor U27865 (N_27865,N_27183,N_27308);
nand U27866 (N_27866,N_27171,N_27355);
nor U27867 (N_27867,N_27574,N_27429);
xor U27868 (N_27868,N_27418,N_27083);
nand U27869 (N_27869,N_27528,N_27493);
nor U27870 (N_27870,N_27061,N_27585);
or U27871 (N_27871,N_27563,N_27545);
and U27872 (N_27872,N_27294,N_27139);
nand U27873 (N_27873,N_27172,N_27059);
and U27874 (N_27874,N_27203,N_27366);
nand U27875 (N_27875,N_27467,N_27184);
nor U27876 (N_27876,N_27238,N_27573);
nor U27877 (N_27877,N_27153,N_27293);
or U27878 (N_27878,N_27170,N_27007);
and U27879 (N_27879,N_27225,N_27276);
nand U27880 (N_27880,N_27197,N_27087);
or U27881 (N_27881,N_27090,N_27586);
and U27882 (N_27882,N_27222,N_27411);
or U27883 (N_27883,N_27496,N_27508);
or U27884 (N_27884,N_27213,N_27487);
or U27885 (N_27885,N_27006,N_27501);
nor U27886 (N_27886,N_27243,N_27593);
nor U27887 (N_27887,N_27533,N_27122);
xnor U27888 (N_27888,N_27568,N_27489);
or U27889 (N_27889,N_27514,N_27353);
xnor U27890 (N_27890,N_27315,N_27014);
xnor U27891 (N_27891,N_27562,N_27227);
or U27892 (N_27892,N_27047,N_27239);
and U27893 (N_27893,N_27301,N_27177);
and U27894 (N_27894,N_27106,N_27525);
and U27895 (N_27895,N_27393,N_27452);
nand U27896 (N_27896,N_27567,N_27241);
or U27897 (N_27897,N_27305,N_27478);
and U27898 (N_27898,N_27248,N_27412);
nor U27899 (N_27899,N_27432,N_27354);
xnor U27900 (N_27900,N_27345,N_27556);
nor U27901 (N_27901,N_27030,N_27418);
nor U27902 (N_27902,N_27482,N_27533);
or U27903 (N_27903,N_27141,N_27211);
nor U27904 (N_27904,N_27516,N_27196);
nand U27905 (N_27905,N_27542,N_27255);
or U27906 (N_27906,N_27188,N_27250);
xnor U27907 (N_27907,N_27329,N_27165);
nand U27908 (N_27908,N_27050,N_27229);
xnor U27909 (N_27909,N_27429,N_27081);
nor U27910 (N_27910,N_27187,N_27511);
and U27911 (N_27911,N_27086,N_27523);
xor U27912 (N_27912,N_27175,N_27017);
nor U27913 (N_27913,N_27170,N_27195);
or U27914 (N_27914,N_27192,N_27281);
and U27915 (N_27915,N_27106,N_27129);
xnor U27916 (N_27916,N_27226,N_27534);
nand U27917 (N_27917,N_27049,N_27574);
nor U27918 (N_27918,N_27360,N_27137);
and U27919 (N_27919,N_27008,N_27026);
xnor U27920 (N_27920,N_27026,N_27489);
nand U27921 (N_27921,N_27513,N_27052);
xor U27922 (N_27922,N_27538,N_27246);
nand U27923 (N_27923,N_27306,N_27463);
nor U27924 (N_27924,N_27221,N_27171);
xor U27925 (N_27925,N_27470,N_27382);
or U27926 (N_27926,N_27448,N_27043);
nand U27927 (N_27927,N_27531,N_27130);
xor U27928 (N_27928,N_27006,N_27362);
and U27929 (N_27929,N_27084,N_27407);
or U27930 (N_27930,N_27487,N_27590);
nand U27931 (N_27931,N_27260,N_27066);
nor U27932 (N_27932,N_27117,N_27168);
nand U27933 (N_27933,N_27263,N_27179);
xor U27934 (N_27934,N_27062,N_27421);
and U27935 (N_27935,N_27237,N_27551);
nand U27936 (N_27936,N_27075,N_27514);
nand U27937 (N_27937,N_27520,N_27357);
and U27938 (N_27938,N_27249,N_27158);
and U27939 (N_27939,N_27151,N_27447);
nor U27940 (N_27940,N_27526,N_27475);
nand U27941 (N_27941,N_27384,N_27315);
or U27942 (N_27942,N_27548,N_27222);
nand U27943 (N_27943,N_27383,N_27019);
nand U27944 (N_27944,N_27177,N_27495);
nand U27945 (N_27945,N_27318,N_27403);
nand U27946 (N_27946,N_27174,N_27535);
or U27947 (N_27947,N_27493,N_27458);
or U27948 (N_27948,N_27024,N_27384);
and U27949 (N_27949,N_27317,N_27145);
or U27950 (N_27950,N_27466,N_27126);
and U27951 (N_27951,N_27132,N_27323);
nand U27952 (N_27952,N_27211,N_27066);
and U27953 (N_27953,N_27312,N_27021);
nor U27954 (N_27954,N_27089,N_27178);
nor U27955 (N_27955,N_27050,N_27129);
nor U27956 (N_27956,N_27174,N_27477);
or U27957 (N_27957,N_27271,N_27102);
nand U27958 (N_27958,N_27495,N_27143);
xnor U27959 (N_27959,N_27527,N_27141);
or U27960 (N_27960,N_27014,N_27162);
nand U27961 (N_27961,N_27472,N_27508);
nor U27962 (N_27962,N_27092,N_27593);
nand U27963 (N_27963,N_27301,N_27362);
and U27964 (N_27964,N_27586,N_27572);
and U27965 (N_27965,N_27324,N_27176);
or U27966 (N_27966,N_27063,N_27319);
nor U27967 (N_27967,N_27302,N_27080);
or U27968 (N_27968,N_27538,N_27197);
nand U27969 (N_27969,N_27354,N_27453);
nor U27970 (N_27970,N_27338,N_27003);
nand U27971 (N_27971,N_27422,N_27250);
and U27972 (N_27972,N_27196,N_27500);
nor U27973 (N_27973,N_27492,N_27146);
or U27974 (N_27974,N_27334,N_27341);
xnor U27975 (N_27975,N_27467,N_27480);
nor U27976 (N_27976,N_27515,N_27275);
and U27977 (N_27977,N_27537,N_27058);
nor U27978 (N_27978,N_27163,N_27316);
nor U27979 (N_27979,N_27560,N_27592);
nand U27980 (N_27980,N_27177,N_27043);
nor U27981 (N_27981,N_27217,N_27377);
nand U27982 (N_27982,N_27006,N_27316);
and U27983 (N_27983,N_27027,N_27300);
nor U27984 (N_27984,N_27054,N_27467);
nor U27985 (N_27985,N_27314,N_27139);
nor U27986 (N_27986,N_27382,N_27243);
nor U27987 (N_27987,N_27015,N_27098);
or U27988 (N_27988,N_27422,N_27234);
or U27989 (N_27989,N_27540,N_27001);
and U27990 (N_27990,N_27086,N_27043);
or U27991 (N_27991,N_27293,N_27583);
xnor U27992 (N_27992,N_27193,N_27093);
and U27993 (N_27993,N_27326,N_27005);
nor U27994 (N_27994,N_27195,N_27225);
and U27995 (N_27995,N_27324,N_27578);
nand U27996 (N_27996,N_27154,N_27537);
or U27997 (N_27997,N_27376,N_27042);
or U27998 (N_27998,N_27503,N_27007);
and U27999 (N_27999,N_27414,N_27558);
and U28000 (N_28000,N_27141,N_27136);
or U28001 (N_28001,N_27324,N_27434);
xnor U28002 (N_28002,N_27549,N_27421);
nor U28003 (N_28003,N_27474,N_27410);
nor U28004 (N_28004,N_27087,N_27149);
nor U28005 (N_28005,N_27597,N_27396);
nor U28006 (N_28006,N_27419,N_27296);
and U28007 (N_28007,N_27321,N_27105);
or U28008 (N_28008,N_27286,N_27283);
nand U28009 (N_28009,N_27257,N_27213);
nor U28010 (N_28010,N_27356,N_27041);
xor U28011 (N_28011,N_27574,N_27148);
nor U28012 (N_28012,N_27574,N_27367);
nand U28013 (N_28013,N_27315,N_27067);
nand U28014 (N_28014,N_27112,N_27570);
or U28015 (N_28015,N_27285,N_27107);
xor U28016 (N_28016,N_27488,N_27041);
or U28017 (N_28017,N_27359,N_27508);
nand U28018 (N_28018,N_27412,N_27511);
and U28019 (N_28019,N_27038,N_27413);
nor U28020 (N_28020,N_27198,N_27354);
nor U28021 (N_28021,N_27378,N_27517);
and U28022 (N_28022,N_27480,N_27275);
nand U28023 (N_28023,N_27217,N_27192);
xnor U28024 (N_28024,N_27378,N_27424);
xnor U28025 (N_28025,N_27494,N_27386);
nand U28026 (N_28026,N_27084,N_27426);
xnor U28027 (N_28027,N_27590,N_27217);
and U28028 (N_28028,N_27159,N_27563);
xnor U28029 (N_28029,N_27473,N_27434);
or U28030 (N_28030,N_27217,N_27552);
xor U28031 (N_28031,N_27553,N_27102);
and U28032 (N_28032,N_27001,N_27459);
nand U28033 (N_28033,N_27068,N_27129);
and U28034 (N_28034,N_27001,N_27027);
nor U28035 (N_28035,N_27455,N_27396);
or U28036 (N_28036,N_27444,N_27331);
or U28037 (N_28037,N_27342,N_27572);
or U28038 (N_28038,N_27318,N_27127);
nor U28039 (N_28039,N_27347,N_27583);
and U28040 (N_28040,N_27251,N_27011);
and U28041 (N_28041,N_27032,N_27049);
and U28042 (N_28042,N_27301,N_27265);
nor U28043 (N_28043,N_27259,N_27554);
xor U28044 (N_28044,N_27561,N_27583);
and U28045 (N_28045,N_27181,N_27056);
and U28046 (N_28046,N_27112,N_27027);
and U28047 (N_28047,N_27216,N_27203);
nor U28048 (N_28048,N_27581,N_27141);
nor U28049 (N_28049,N_27217,N_27309);
xor U28050 (N_28050,N_27058,N_27070);
nor U28051 (N_28051,N_27378,N_27191);
and U28052 (N_28052,N_27183,N_27454);
nand U28053 (N_28053,N_27390,N_27023);
or U28054 (N_28054,N_27106,N_27231);
xor U28055 (N_28055,N_27225,N_27269);
and U28056 (N_28056,N_27381,N_27316);
or U28057 (N_28057,N_27415,N_27273);
or U28058 (N_28058,N_27473,N_27013);
or U28059 (N_28059,N_27429,N_27074);
or U28060 (N_28060,N_27238,N_27121);
and U28061 (N_28061,N_27450,N_27573);
or U28062 (N_28062,N_27581,N_27222);
or U28063 (N_28063,N_27073,N_27368);
xnor U28064 (N_28064,N_27559,N_27402);
or U28065 (N_28065,N_27556,N_27179);
nor U28066 (N_28066,N_27098,N_27361);
xnor U28067 (N_28067,N_27555,N_27171);
xnor U28068 (N_28068,N_27181,N_27296);
nor U28069 (N_28069,N_27562,N_27316);
nor U28070 (N_28070,N_27480,N_27487);
xor U28071 (N_28071,N_27256,N_27317);
and U28072 (N_28072,N_27487,N_27206);
nand U28073 (N_28073,N_27327,N_27123);
nor U28074 (N_28074,N_27199,N_27248);
nand U28075 (N_28075,N_27261,N_27519);
xnor U28076 (N_28076,N_27246,N_27402);
or U28077 (N_28077,N_27406,N_27476);
or U28078 (N_28078,N_27459,N_27451);
and U28079 (N_28079,N_27249,N_27241);
nand U28080 (N_28080,N_27474,N_27212);
and U28081 (N_28081,N_27190,N_27586);
or U28082 (N_28082,N_27379,N_27324);
nor U28083 (N_28083,N_27550,N_27317);
and U28084 (N_28084,N_27559,N_27082);
nor U28085 (N_28085,N_27358,N_27553);
nor U28086 (N_28086,N_27135,N_27064);
or U28087 (N_28087,N_27239,N_27144);
nand U28088 (N_28088,N_27247,N_27566);
nand U28089 (N_28089,N_27209,N_27257);
xor U28090 (N_28090,N_27530,N_27173);
xor U28091 (N_28091,N_27415,N_27320);
nand U28092 (N_28092,N_27081,N_27179);
nand U28093 (N_28093,N_27159,N_27067);
nand U28094 (N_28094,N_27214,N_27087);
nand U28095 (N_28095,N_27071,N_27400);
and U28096 (N_28096,N_27439,N_27212);
nand U28097 (N_28097,N_27287,N_27467);
nand U28098 (N_28098,N_27523,N_27185);
xnor U28099 (N_28099,N_27494,N_27052);
nand U28100 (N_28100,N_27341,N_27259);
xnor U28101 (N_28101,N_27556,N_27534);
nand U28102 (N_28102,N_27010,N_27371);
nand U28103 (N_28103,N_27521,N_27569);
nand U28104 (N_28104,N_27112,N_27559);
nor U28105 (N_28105,N_27407,N_27123);
or U28106 (N_28106,N_27079,N_27255);
or U28107 (N_28107,N_27344,N_27257);
nand U28108 (N_28108,N_27019,N_27473);
nor U28109 (N_28109,N_27561,N_27086);
nor U28110 (N_28110,N_27415,N_27092);
nor U28111 (N_28111,N_27006,N_27236);
nand U28112 (N_28112,N_27044,N_27105);
and U28113 (N_28113,N_27379,N_27174);
nand U28114 (N_28114,N_27293,N_27445);
and U28115 (N_28115,N_27026,N_27239);
nor U28116 (N_28116,N_27120,N_27194);
and U28117 (N_28117,N_27590,N_27324);
or U28118 (N_28118,N_27584,N_27155);
xnor U28119 (N_28119,N_27015,N_27171);
xor U28120 (N_28120,N_27241,N_27481);
nand U28121 (N_28121,N_27014,N_27394);
nor U28122 (N_28122,N_27271,N_27011);
and U28123 (N_28123,N_27458,N_27577);
xor U28124 (N_28124,N_27479,N_27103);
and U28125 (N_28125,N_27043,N_27171);
nor U28126 (N_28126,N_27425,N_27250);
xnor U28127 (N_28127,N_27223,N_27440);
nand U28128 (N_28128,N_27260,N_27587);
xor U28129 (N_28129,N_27099,N_27169);
nand U28130 (N_28130,N_27112,N_27101);
and U28131 (N_28131,N_27018,N_27462);
or U28132 (N_28132,N_27201,N_27170);
xor U28133 (N_28133,N_27146,N_27324);
nand U28134 (N_28134,N_27456,N_27359);
and U28135 (N_28135,N_27393,N_27282);
nand U28136 (N_28136,N_27312,N_27517);
nor U28137 (N_28137,N_27289,N_27316);
nor U28138 (N_28138,N_27576,N_27545);
or U28139 (N_28139,N_27108,N_27060);
xor U28140 (N_28140,N_27429,N_27082);
or U28141 (N_28141,N_27342,N_27386);
or U28142 (N_28142,N_27364,N_27545);
or U28143 (N_28143,N_27261,N_27127);
nand U28144 (N_28144,N_27587,N_27140);
nor U28145 (N_28145,N_27512,N_27261);
nor U28146 (N_28146,N_27553,N_27182);
or U28147 (N_28147,N_27047,N_27320);
or U28148 (N_28148,N_27428,N_27238);
or U28149 (N_28149,N_27182,N_27300);
nand U28150 (N_28150,N_27210,N_27303);
xor U28151 (N_28151,N_27437,N_27034);
nand U28152 (N_28152,N_27018,N_27221);
nand U28153 (N_28153,N_27104,N_27219);
nand U28154 (N_28154,N_27185,N_27124);
and U28155 (N_28155,N_27004,N_27509);
nand U28156 (N_28156,N_27569,N_27359);
xnor U28157 (N_28157,N_27373,N_27386);
nand U28158 (N_28158,N_27029,N_27535);
and U28159 (N_28159,N_27133,N_27253);
nand U28160 (N_28160,N_27399,N_27263);
xnor U28161 (N_28161,N_27114,N_27306);
xor U28162 (N_28162,N_27243,N_27042);
and U28163 (N_28163,N_27501,N_27168);
or U28164 (N_28164,N_27472,N_27262);
and U28165 (N_28165,N_27359,N_27382);
and U28166 (N_28166,N_27118,N_27463);
xor U28167 (N_28167,N_27323,N_27501);
or U28168 (N_28168,N_27560,N_27596);
and U28169 (N_28169,N_27232,N_27007);
or U28170 (N_28170,N_27548,N_27436);
and U28171 (N_28171,N_27079,N_27540);
nand U28172 (N_28172,N_27112,N_27524);
xor U28173 (N_28173,N_27447,N_27558);
and U28174 (N_28174,N_27269,N_27588);
or U28175 (N_28175,N_27004,N_27160);
nand U28176 (N_28176,N_27024,N_27147);
nor U28177 (N_28177,N_27576,N_27219);
and U28178 (N_28178,N_27206,N_27491);
xor U28179 (N_28179,N_27206,N_27095);
nand U28180 (N_28180,N_27327,N_27257);
nor U28181 (N_28181,N_27011,N_27301);
xor U28182 (N_28182,N_27245,N_27002);
nor U28183 (N_28183,N_27408,N_27582);
xnor U28184 (N_28184,N_27167,N_27599);
nor U28185 (N_28185,N_27584,N_27285);
nand U28186 (N_28186,N_27532,N_27549);
and U28187 (N_28187,N_27166,N_27583);
or U28188 (N_28188,N_27292,N_27476);
xor U28189 (N_28189,N_27232,N_27051);
xnor U28190 (N_28190,N_27286,N_27371);
and U28191 (N_28191,N_27485,N_27512);
xor U28192 (N_28192,N_27192,N_27594);
nand U28193 (N_28193,N_27243,N_27537);
or U28194 (N_28194,N_27264,N_27190);
or U28195 (N_28195,N_27149,N_27281);
nand U28196 (N_28196,N_27366,N_27303);
or U28197 (N_28197,N_27443,N_27315);
xor U28198 (N_28198,N_27037,N_27523);
or U28199 (N_28199,N_27116,N_27275);
and U28200 (N_28200,N_28186,N_28008);
nor U28201 (N_28201,N_28047,N_28141);
and U28202 (N_28202,N_27840,N_27749);
or U28203 (N_28203,N_28016,N_27848);
nor U28204 (N_28204,N_27913,N_28143);
and U28205 (N_28205,N_27744,N_27951);
or U28206 (N_28206,N_27740,N_27900);
nand U28207 (N_28207,N_27783,N_27958);
nand U28208 (N_28208,N_28136,N_28063);
and U28209 (N_28209,N_28086,N_28028);
and U28210 (N_28210,N_27683,N_28198);
nand U28211 (N_28211,N_27982,N_28105);
or U28212 (N_28212,N_28101,N_27624);
nor U28213 (N_28213,N_27894,N_27704);
nand U28214 (N_28214,N_27604,N_27633);
nor U28215 (N_28215,N_28004,N_27901);
nor U28216 (N_28216,N_27876,N_28079);
nand U28217 (N_28217,N_27794,N_28187);
xnor U28218 (N_28218,N_27696,N_27795);
and U28219 (N_28219,N_28133,N_28171);
or U28220 (N_28220,N_27738,N_27760);
nor U28221 (N_28221,N_27917,N_27694);
or U28222 (N_28222,N_27879,N_27774);
xor U28223 (N_28223,N_28024,N_27882);
xor U28224 (N_28224,N_27851,N_27976);
or U28225 (N_28225,N_28191,N_28075);
xor U28226 (N_28226,N_27811,N_27810);
or U28227 (N_28227,N_27733,N_27784);
or U28228 (N_28228,N_27943,N_27763);
xnor U28229 (N_28229,N_28166,N_27718);
and U28230 (N_28230,N_27945,N_27643);
and U28231 (N_28231,N_27875,N_27865);
xor U28232 (N_28232,N_27804,N_27939);
and U28233 (N_28233,N_27620,N_27909);
and U28234 (N_28234,N_27841,N_28159);
and U28235 (N_28235,N_27727,N_28072);
xnor U28236 (N_28236,N_27995,N_27666);
nand U28237 (N_28237,N_28054,N_27896);
and U28238 (N_28238,N_28115,N_28123);
and U28239 (N_28239,N_28029,N_27628);
or U28240 (N_28240,N_27916,N_27717);
nand U28241 (N_28241,N_27924,N_27856);
xnor U28242 (N_28242,N_27753,N_27651);
and U28243 (N_28243,N_27824,N_27602);
or U28244 (N_28244,N_27797,N_27729);
nand U28245 (N_28245,N_27808,N_27722);
xnor U28246 (N_28246,N_27748,N_27790);
nand U28247 (N_28247,N_27761,N_27708);
or U28248 (N_28248,N_28089,N_27664);
xnor U28249 (N_28249,N_27908,N_27912);
nor U28250 (N_28250,N_27706,N_27796);
or U28251 (N_28251,N_28144,N_27789);
or U28252 (N_28252,N_27667,N_28190);
or U28253 (N_28253,N_27889,N_27906);
nor U28254 (N_28254,N_27755,N_28062);
and U28255 (N_28255,N_27747,N_27737);
and U28256 (N_28256,N_28006,N_28070);
xnor U28257 (N_28257,N_27685,N_27846);
nand U28258 (N_28258,N_28129,N_27885);
or U28259 (N_28259,N_27746,N_28050);
and U28260 (N_28260,N_27860,N_28180);
xnor U28261 (N_28261,N_27647,N_28130);
nor U28262 (N_28262,N_27881,N_27800);
xnor U28263 (N_28263,N_27682,N_27925);
nor U28264 (N_28264,N_27607,N_28014);
or U28265 (N_28265,N_28027,N_28169);
nand U28266 (N_28266,N_28137,N_27758);
xnor U28267 (N_28267,N_28139,N_27690);
and U28268 (N_28268,N_27726,N_28057);
or U28269 (N_28269,N_27861,N_27780);
and U28270 (N_28270,N_27845,N_28069);
nand U28271 (N_28271,N_27781,N_27741);
or U28272 (N_28272,N_28118,N_28002);
xnor U28273 (N_28273,N_27874,N_28122);
nand U28274 (N_28274,N_28104,N_27688);
or U28275 (N_28275,N_28088,N_27926);
nand U28276 (N_28276,N_28117,N_27970);
xor U28277 (N_28277,N_27921,N_27701);
and U28278 (N_28278,N_28066,N_28087);
nand U28279 (N_28279,N_27999,N_28150);
nor U28280 (N_28280,N_27842,N_27793);
and U28281 (N_28281,N_27659,N_28194);
nor U28282 (N_28282,N_27614,N_28099);
nand U28283 (N_28283,N_27713,N_28055);
and U28284 (N_28284,N_28116,N_28152);
and U28285 (N_28285,N_28102,N_28173);
and U28286 (N_28286,N_28003,N_27960);
or U28287 (N_28287,N_27745,N_28000);
nor U28288 (N_28288,N_27855,N_27836);
nor U28289 (N_28289,N_28084,N_27905);
and U28290 (N_28290,N_28037,N_27806);
nor U28291 (N_28291,N_27634,N_27967);
xnor U28292 (N_28292,N_28012,N_27962);
nor U28293 (N_28293,N_27979,N_27698);
nand U28294 (N_28294,N_27693,N_28030);
or U28295 (N_28295,N_27971,N_28128);
or U28296 (N_28296,N_28042,N_27993);
nand U28297 (N_28297,N_27974,N_27676);
and U28298 (N_28298,N_28167,N_28043);
xor U28299 (N_28299,N_27853,N_27835);
or U28300 (N_28300,N_27692,N_28182);
or U28301 (N_28301,N_28126,N_27644);
xnor U28302 (N_28302,N_27648,N_28013);
and U28303 (N_28303,N_27772,N_27799);
nor U28304 (N_28304,N_27991,N_27878);
nand U28305 (N_28305,N_27764,N_28076);
or U28306 (N_28306,N_27869,N_27877);
or U28307 (N_28307,N_27703,N_28157);
xnor U28308 (N_28308,N_27765,N_28023);
nor U28309 (N_28309,N_27631,N_27898);
nor U28310 (N_28310,N_27966,N_28052);
and U28311 (N_28311,N_27655,N_27972);
or U28312 (N_28312,N_28082,N_27639);
nand U28313 (N_28313,N_28156,N_27981);
nand U28314 (N_28314,N_27814,N_27606);
and U28315 (N_28315,N_28077,N_28192);
and U28316 (N_28316,N_28018,N_28085);
and U28317 (N_28317,N_27801,N_27839);
and U28318 (N_28318,N_28053,N_27903);
and U28319 (N_28319,N_27674,N_27942);
xnor U28320 (N_28320,N_28015,N_28199);
xnor U28321 (N_28321,N_28010,N_27997);
nand U28322 (N_28322,N_27762,N_28036);
nand U28323 (N_28323,N_27719,N_27759);
nor U28324 (N_28324,N_28146,N_27689);
nor U28325 (N_28325,N_27870,N_27857);
xor U28326 (N_28326,N_28090,N_27989);
nor U28327 (N_28327,N_27618,N_27817);
xnor U28328 (N_28328,N_27679,N_28155);
or U28329 (N_28329,N_28138,N_27769);
nand U28330 (N_28330,N_28177,N_27990);
nor U28331 (N_28331,N_27767,N_28021);
and U28332 (N_28332,N_27615,N_27658);
and U28333 (N_28333,N_27669,N_28162);
and U28334 (N_28334,N_27931,N_27968);
nand U28335 (N_28335,N_27776,N_27770);
and U28336 (N_28336,N_28149,N_28196);
or U28337 (N_28337,N_27973,N_27854);
nand U28338 (N_28338,N_27673,N_27986);
nand U28339 (N_28339,N_27725,N_27994);
xnor U28340 (N_28340,N_27757,N_28168);
nand U28341 (N_28341,N_28114,N_27734);
nand U28342 (N_28342,N_27754,N_27812);
or U28343 (N_28343,N_27635,N_27630);
or U28344 (N_28344,N_27697,N_27601);
nand U28345 (N_28345,N_27961,N_27805);
or U28346 (N_28346,N_28151,N_27695);
nand U28347 (N_28347,N_27775,N_27732);
or U28348 (N_28348,N_27975,N_27867);
nor U28349 (N_28349,N_28046,N_28125);
or U28350 (N_28350,N_27935,N_28161);
nand U28351 (N_28351,N_27652,N_27743);
and U28352 (N_28352,N_28051,N_27678);
and U28353 (N_28353,N_27807,N_27700);
nand U28354 (N_28354,N_27815,N_28153);
nand U28355 (N_28355,N_27965,N_27709);
nand U28356 (N_28356,N_27936,N_27619);
nor U28357 (N_28357,N_27629,N_27645);
or U28358 (N_28358,N_27720,N_27863);
nor U28359 (N_28359,N_28098,N_27895);
xnor U28360 (N_28360,N_28103,N_27904);
nor U28361 (N_28361,N_28031,N_27803);
or U28362 (N_28362,N_27985,N_27608);
and U28363 (N_28363,N_27650,N_27665);
and U28364 (N_28364,N_27886,N_28060);
xnor U28365 (N_28365,N_27662,N_27777);
and U28366 (N_28366,N_28121,N_28148);
nor U28367 (N_28367,N_27640,N_27829);
xor U28368 (N_28368,N_28080,N_27788);
and U28369 (N_28369,N_27778,N_27914);
nor U28370 (N_28370,N_27712,N_28174);
or U28371 (N_28371,N_28093,N_27929);
and U28372 (N_28372,N_27837,N_27707);
nor U28373 (N_28373,N_27826,N_27899);
or U28374 (N_28374,N_27978,N_27933);
or U28375 (N_28375,N_27668,N_27786);
or U28376 (N_28376,N_27963,N_27956);
nand U28377 (N_28377,N_28134,N_28179);
xnor U28378 (N_28378,N_28067,N_27792);
nor U28379 (N_28379,N_27819,N_28061);
and U28380 (N_28380,N_27802,N_27821);
nor U28381 (N_28381,N_27852,N_27736);
nand U28382 (N_28382,N_27616,N_27779);
or U28383 (N_28383,N_28007,N_28183);
xor U28384 (N_28384,N_27957,N_28193);
nor U28385 (N_28385,N_28108,N_27605);
or U28386 (N_28386,N_27730,N_28044);
xnor U28387 (N_28387,N_28033,N_28112);
xnor U28388 (N_28388,N_28113,N_27827);
nand U28389 (N_28389,N_28058,N_27897);
xnor U28390 (N_28390,N_27996,N_28059);
or U28391 (N_28391,N_28096,N_27813);
nor U28392 (N_28392,N_28120,N_28100);
xor U28393 (N_28393,N_27686,N_27934);
or U28394 (N_28394,N_27773,N_27623);
xnor U28395 (N_28395,N_27663,N_27626);
and U28396 (N_28396,N_27980,N_28020);
xor U28397 (N_28397,N_27656,N_28025);
nor U28398 (N_28398,N_27910,N_28092);
nor U28399 (N_28399,N_28035,N_27822);
nor U28400 (N_28400,N_28009,N_28165);
nand U28401 (N_28401,N_28064,N_27723);
and U28402 (N_28402,N_28040,N_27834);
nor U28403 (N_28403,N_27959,N_27646);
xor U28404 (N_28404,N_27661,N_27735);
and U28405 (N_28405,N_27883,N_27617);
and U28406 (N_28406,N_27715,N_28189);
nor U28407 (N_28407,N_28073,N_28163);
xor U28408 (N_28408,N_27654,N_27642);
nor U28409 (N_28409,N_27681,N_27907);
and U28410 (N_28410,N_27785,N_27705);
or U28411 (N_28411,N_28124,N_28097);
nand U28412 (N_28412,N_27750,N_28041);
nor U28413 (N_28413,N_28074,N_28140);
or U28414 (N_28414,N_28127,N_28175);
nand U28415 (N_28415,N_27838,N_28065);
nor U28416 (N_28416,N_27809,N_27911);
nor U28417 (N_28417,N_27684,N_27998);
or U28418 (N_28418,N_27977,N_27636);
or U28419 (N_28419,N_28083,N_27955);
or U28420 (N_28420,N_27702,N_28048);
xor U28421 (N_28421,N_27830,N_28094);
and U28422 (N_28422,N_28011,N_27849);
nand U28423 (N_28423,N_27710,N_27902);
xnor U28424 (N_28424,N_27791,N_27677);
or U28425 (N_28425,N_28176,N_27649);
or U28426 (N_28426,N_28001,N_28132);
nand U28427 (N_28427,N_27739,N_27766);
and U28428 (N_28428,N_28034,N_27922);
nand U28429 (N_28429,N_27862,N_27890);
xnor U28430 (N_28430,N_27872,N_27610);
nor U28431 (N_28431,N_27888,N_28039);
and U28432 (N_28432,N_28026,N_27600);
xor U28433 (N_28433,N_27675,N_27609);
xnor U28434 (N_28434,N_27884,N_28038);
nor U28435 (N_28435,N_27731,N_27944);
nand U28436 (N_28436,N_27847,N_27954);
or U28437 (N_28437,N_27742,N_27938);
or U28438 (N_28438,N_28195,N_27949);
xnor U28439 (N_28439,N_28185,N_27641);
xor U28440 (N_28440,N_28131,N_27831);
nor U28441 (N_28441,N_27724,N_28181);
nor U28442 (N_28442,N_28045,N_27947);
or U28443 (N_28443,N_27887,N_27820);
and U28444 (N_28444,N_28119,N_27871);
nor U28445 (N_28445,N_27714,N_27672);
xnor U28446 (N_28446,N_28197,N_27627);
and U28447 (N_28447,N_27637,N_27653);
nor U28448 (N_28448,N_27782,N_27940);
and U28449 (N_28449,N_28160,N_27687);
nand U28450 (N_28450,N_28170,N_27930);
or U28451 (N_28451,N_27858,N_28019);
and U28452 (N_28452,N_28178,N_27920);
nand U28453 (N_28453,N_28106,N_27816);
and U28454 (N_28454,N_27915,N_27632);
or U28455 (N_28455,N_27657,N_28110);
and U28456 (N_28456,N_28068,N_27964);
nand U28457 (N_28457,N_27953,N_27927);
or U28458 (N_28458,N_27880,N_27613);
and U28459 (N_28459,N_27711,N_27660);
xnor U28460 (N_28460,N_27728,N_28056);
nor U28461 (N_28461,N_27843,N_28135);
nand U28462 (N_28462,N_27603,N_28184);
nor U28463 (N_28463,N_27721,N_27850);
nor U28464 (N_28464,N_28078,N_27611);
nor U28465 (N_28465,N_27992,N_28049);
or U28466 (N_28466,N_27948,N_27756);
nand U28467 (N_28467,N_27787,N_27621);
nor U28468 (N_28468,N_27987,N_27932);
nand U28469 (N_28469,N_27864,N_28017);
or U28470 (N_28470,N_27983,N_27825);
and U28471 (N_28471,N_28145,N_27638);
nor U28472 (N_28472,N_28107,N_28172);
and U28473 (N_28473,N_27859,N_28147);
nor U28474 (N_28474,N_27893,N_27868);
and U28475 (N_28475,N_27716,N_27671);
and U28476 (N_28476,N_27891,N_27984);
and U28477 (N_28477,N_27952,N_27892);
or U28478 (N_28478,N_27950,N_28142);
and U28479 (N_28479,N_27988,N_28081);
nor U28480 (N_28480,N_27918,N_28188);
nand U28481 (N_28481,N_27818,N_28111);
xnor U28482 (N_28482,N_28032,N_27691);
nand U28483 (N_28483,N_27866,N_27625);
nand U28484 (N_28484,N_27832,N_28071);
or U28485 (N_28485,N_27823,N_28164);
and U28486 (N_28486,N_28158,N_27768);
xnor U28487 (N_28487,N_27622,N_27699);
xnor U28488 (N_28488,N_27670,N_27923);
and U28489 (N_28489,N_27771,N_27941);
xor U28490 (N_28490,N_28091,N_27833);
nand U28491 (N_28491,N_28109,N_27751);
nor U28492 (N_28492,N_27752,N_27919);
or U28493 (N_28493,N_27612,N_27946);
xor U28494 (N_28494,N_28154,N_27969);
or U28495 (N_28495,N_27928,N_27680);
and U28496 (N_28496,N_27798,N_27844);
nor U28497 (N_28497,N_27937,N_27873);
and U28498 (N_28498,N_28005,N_28095);
xnor U28499 (N_28499,N_27828,N_28022);
nor U28500 (N_28500,N_27821,N_28087);
and U28501 (N_28501,N_27824,N_28048);
xnor U28502 (N_28502,N_28065,N_27718);
and U28503 (N_28503,N_27853,N_27643);
and U28504 (N_28504,N_28027,N_28177);
or U28505 (N_28505,N_28041,N_28185);
and U28506 (N_28506,N_27908,N_27624);
and U28507 (N_28507,N_27693,N_27738);
and U28508 (N_28508,N_27765,N_28185);
xnor U28509 (N_28509,N_28170,N_27851);
nor U28510 (N_28510,N_27675,N_27610);
or U28511 (N_28511,N_27788,N_27632);
or U28512 (N_28512,N_27924,N_28141);
and U28513 (N_28513,N_27624,N_27600);
and U28514 (N_28514,N_27831,N_27986);
nor U28515 (N_28515,N_27689,N_27889);
or U28516 (N_28516,N_28129,N_28186);
nand U28517 (N_28517,N_27611,N_28167);
or U28518 (N_28518,N_28130,N_28084);
or U28519 (N_28519,N_27979,N_28046);
or U28520 (N_28520,N_28114,N_28027);
xnor U28521 (N_28521,N_27693,N_28078);
or U28522 (N_28522,N_27979,N_27798);
nor U28523 (N_28523,N_27812,N_27771);
nor U28524 (N_28524,N_28008,N_28003);
or U28525 (N_28525,N_27618,N_27814);
nor U28526 (N_28526,N_27849,N_27635);
nand U28527 (N_28527,N_27774,N_27659);
and U28528 (N_28528,N_27692,N_27879);
and U28529 (N_28529,N_27755,N_27678);
nor U28530 (N_28530,N_27632,N_28107);
or U28531 (N_28531,N_28103,N_27914);
and U28532 (N_28532,N_28157,N_27635);
xnor U28533 (N_28533,N_28088,N_28019);
or U28534 (N_28534,N_27704,N_27827);
nor U28535 (N_28535,N_27641,N_27820);
xnor U28536 (N_28536,N_27907,N_28097);
or U28537 (N_28537,N_28052,N_27668);
xor U28538 (N_28538,N_27682,N_27931);
xor U28539 (N_28539,N_27794,N_27861);
or U28540 (N_28540,N_27865,N_27859);
nand U28541 (N_28541,N_28139,N_27887);
nand U28542 (N_28542,N_27726,N_28134);
xor U28543 (N_28543,N_27806,N_27810);
or U28544 (N_28544,N_27653,N_27968);
xnor U28545 (N_28545,N_28089,N_28133);
and U28546 (N_28546,N_27762,N_27970);
nand U28547 (N_28547,N_27605,N_28154);
nand U28548 (N_28548,N_28076,N_27644);
xnor U28549 (N_28549,N_28161,N_27722);
and U28550 (N_28550,N_28078,N_27977);
nand U28551 (N_28551,N_27765,N_27996);
nor U28552 (N_28552,N_27633,N_28018);
or U28553 (N_28553,N_27737,N_27726);
nor U28554 (N_28554,N_27850,N_27635);
and U28555 (N_28555,N_28032,N_27774);
and U28556 (N_28556,N_27633,N_28080);
or U28557 (N_28557,N_28065,N_27994);
nand U28558 (N_28558,N_27886,N_28029);
nand U28559 (N_28559,N_27949,N_28110);
or U28560 (N_28560,N_28068,N_27730);
nor U28561 (N_28561,N_28182,N_27732);
and U28562 (N_28562,N_27947,N_27613);
or U28563 (N_28563,N_27948,N_27625);
nand U28564 (N_28564,N_27702,N_27609);
or U28565 (N_28565,N_28008,N_28160);
nand U28566 (N_28566,N_27955,N_28047);
xnor U28567 (N_28567,N_27619,N_28033);
and U28568 (N_28568,N_27979,N_27963);
and U28569 (N_28569,N_28049,N_27619);
and U28570 (N_28570,N_28074,N_27613);
nor U28571 (N_28571,N_27704,N_27602);
or U28572 (N_28572,N_27842,N_28055);
nand U28573 (N_28573,N_27943,N_27649);
xnor U28574 (N_28574,N_27615,N_27983);
nand U28575 (N_28575,N_28046,N_27816);
nor U28576 (N_28576,N_28168,N_28080);
and U28577 (N_28577,N_28111,N_27623);
xnor U28578 (N_28578,N_27752,N_27830);
nor U28579 (N_28579,N_28019,N_27706);
or U28580 (N_28580,N_27781,N_27735);
xnor U28581 (N_28581,N_28055,N_27948);
nor U28582 (N_28582,N_27730,N_27825);
or U28583 (N_28583,N_27778,N_27720);
xor U28584 (N_28584,N_27622,N_27930);
and U28585 (N_28585,N_27902,N_27609);
xnor U28586 (N_28586,N_27698,N_28171);
nor U28587 (N_28587,N_27819,N_27638);
or U28588 (N_28588,N_27708,N_27799);
nor U28589 (N_28589,N_27843,N_27704);
nor U28590 (N_28590,N_27700,N_27913);
and U28591 (N_28591,N_27824,N_27887);
or U28592 (N_28592,N_27959,N_28038);
nor U28593 (N_28593,N_27823,N_27944);
nor U28594 (N_28594,N_28168,N_27703);
or U28595 (N_28595,N_27889,N_27873);
or U28596 (N_28596,N_27619,N_27688);
or U28597 (N_28597,N_27732,N_27782);
and U28598 (N_28598,N_27731,N_28188);
xnor U28599 (N_28599,N_28102,N_27960);
or U28600 (N_28600,N_27922,N_27616);
nor U28601 (N_28601,N_27868,N_27600);
xor U28602 (N_28602,N_27747,N_27988);
and U28603 (N_28603,N_27620,N_27958);
or U28604 (N_28604,N_27954,N_27717);
xnor U28605 (N_28605,N_27937,N_27666);
nor U28606 (N_28606,N_27948,N_28007);
xnor U28607 (N_28607,N_27816,N_27764);
nor U28608 (N_28608,N_28075,N_27822);
or U28609 (N_28609,N_27985,N_27839);
xor U28610 (N_28610,N_28058,N_28008);
or U28611 (N_28611,N_27755,N_28188);
nor U28612 (N_28612,N_28139,N_27708);
xor U28613 (N_28613,N_28181,N_27807);
nor U28614 (N_28614,N_27902,N_28041);
or U28615 (N_28615,N_27876,N_27827);
or U28616 (N_28616,N_27745,N_27600);
nor U28617 (N_28617,N_28118,N_27655);
and U28618 (N_28618,N_27783,N_27654);
nand U28619 (N_28619,N_28142,N_27657);
nand U28620 (N_28620,N_27715,N_28077);
nand U28621 (N_28621,N_28083,N_27687);
or U28622 (N_28622,N_27850,N_28166);
or U28623 (N_28623,N_28189,N_28066);
nand U28624 (N_28624,N_28161,N_27646);
and U28625 (N_28625,N_27993,N_27893);
or U28626 (N_28626,N_27655,N_28022);
nor U28627 (N_28627,N_27902,N_27656);
and U28628 (N_28628,N_28014,N_27905);
xor U28629 (N_28629,N_27803,N_27839);
nand U28630 (N_28630,N_27618,N_28145);
or U28631 (N_28631,N_27622,N_28072);
and U28632 (N_28632,N_27933,N_28191);
and U28633 (N_28633,N_27934,N_28024);
xor U28634 (N_28634,N_27631,N_27986);
xnor U28635 (N_28635,N_28074,N_27673);
and U28636 (N_28636,N_27670,N_28067);
and U28637 (N_28637,N_27938,N_27674);
xnor U28638 (N_28638,N_27890,N_28153);
nand U28639 (N_28639,N_28169,N_27826);
nand U28640 (N_28640,N_27620,N_27986);
nor U28641 (N_28641,N_27965,N_27924);
or U28642 (N_28642,N_28167,N_28162);
xnor U28643 (N_28643,N_28199,N_27849);
nand U28644 (N_28644,N_27612,N_27642);
xor U28645 (N_28645,N_27867,N_27926);
or U28646 (N_28646,N_28130,N_27875);
xnor U28647 (N_28647,N_28165,N_27871);
nor U28648 (N_28648,N_28011,N_27982);
nor U28649 (N_28649,N_27924,N_27950);
or U28650 (N_28650,N_27604,N_27802);
nand U28651 (N_28651,N_27633,N_28164);
xnor U28652 (N_28652,N_28054,N_27784);
nor U28653 (N_28653,N_27897,N_27730);
nor U28654 (N_28654,N_28017,N_27603);
or U28655 (N_28655,N_27696,N_27689);
and U28656 (N_28656,N_27958,N_27971);
and U28657 (N_28657,N_28134,N_28079);
or U28658 (N_28658,N_27890,N_27915);
and U28659 (N_28659,N_27685,N_27865);
or U28660 (N_28660,N_27819,N_27632);
and U28661 (N_28661,N_27646,N_27694);
nand U28662 (N_28662,N_28129,N_28056);
nor U28663 (N_28663,N_27949,N_28141);
nor U28664 (N_28664,N_28143,N_27896);
and U28665 (N_28665,N_28047,N_28098);
xor U28666 (N_28666,N_28075,N_27932);
nand U28667 (N_28667,N_28043,N_28115);
or U28668 (N_28668,N_28049,N_28011);
xor U28669 (N_28669,N_28099,N_27896);
or U28670 (N_28670,N_27982,N_27781);
or U28671 (N_28671,N_27830,N_27918);
nand U28672 (N_28672,N_28170,N_27955);
or U28673 (N_28673,N_27914,N_27749);
nand U28674 (N_28674,N_27616,N_28151);
or U28675 (N_28675,N_27978,N_27985);
xor U28676 (N_28676,N_28106,N_27875);
and U28677 (N_28677,N_28156,N_27858);
and U28678 (N_28678,N_28197,N_27678);
and U28679 (N_28679,N_27859,N_27844);
and U28680 (N_28680,N_27837,N_27728);
nor U28681 (N_28681,N_27787,N_28177);
or U28682 (N_28682,N_28142,N_28108);
nor U28683 (N_28683,N_28103,N_28113);
nand U28684 (N_28684,N_27670,N_27906);
and U28685 (N_28685,N_27865,N_27839);
xor U28686 (N_28686,N_28164,N_27676);
and U28687 (N_28687,N_28198,N_28006);
xnor U28688 (N_28688,N_28073,N_27634);
nand U28689 (N_28689,N_28060,N_27968);
nand U28690 (N_28690,N_28014,N_27779);
nor U28691 (N_28691,N_27899,N_27867);
or U28692 (N_28692,N_27919,N_28185);
and U28693 (N_28693,N_28181,N_27769);
xor U28694 (N_28694,N_27703,N_28107);
nor U28695 (N_28695,N_27807,N_27912);
nor U28696 (N_28696,N_28090,N_27622);
nand U28697 (N_28697,N_28179,N_27867);
or U28698 (N_28698,N_27744,N_28034);
or U28699 (N_28699,N_27892,N_28181);
or U28700 (N_28700,N_28131,N_27686);
or U28701 (N_28701,N_28119,N_27938);
nor U28702 (N_28702,N_27743,N_27992);
and U28703 (N_28703,N_27862,N_27765);
xnor U28704 (N_28704,N_27797,N_27846);
nor U28705 (N_28705,N_27613,N_28162);
nand U28706 (N_28706,N_27903,N_27797);
nor U28707 (N_28707,N_28150,N_28012);
nand U28708 (N_28708,N_28174,N_27801);
and U28709 (N_28709,N_27805,N_27663);
and U28710 (N_28710,N_27783,N_28019);
xor U28711 (N_28711,N_27899,N_27848);
and U28712 (N_28712,N_28139,N_27606);
xor U28713 (N_28713,N_27964,N_27680);
xnor U28714 (N_28714,N_27991,N_27786);
nor U28715 (N_28715,N_27860,N_27847);
and U28716 (N_28716,N_27628,N_27902);
and U28717 (N_28717,N_27983,N_28070);
and U28718 (N_28718,N_27856,N_28039);
or U28719 (N_28719,N_28151,N_27603);
nor U28720 (N_28720,N_27739,N_27699);
or U28721 (N_28721,N_28098,N_27849);
nor U28722 (N_28722,N_27648,N_28165);
nor U28723 (N_28723,N_28057,N_27997);
nor U28724 (N_28724,N_27764,N_27908);
nand U28725 (N_28725,N_27747,N_27966);
and U28726 (N_28726,N_28059,N_27658);
and U28727 (N_28727,N_28157,N_27813);
nor U28728 (N_28728,N_28102,N_28058);
or U28729 (N_28729,N_27933,N_28067);
and U28730 (N_28730,N_27684,N_27689);
or U28731 (N_28731,N_27859,N_27661);
xnor U28732 (N_28732,N_27776,N_27819);
nand U28733 (N_28733,N_27838,N_28039);
or U28734 (N_28734,N_27885,N_28141);
nand U28735 (N_28735,N_27760,N_27845);
and U28736 (N_28736,N_27877,N_27745);
nand U28737 (N_28737,N_27820,N_27711);
or U28738 (N_28738,N_27700,N_27743);
xor U28739 (N_28739,N_27999,N_27963);
and U28740 (N_28740,N_28069,N_27706);
and U28741 (N_28741,N_27693,N_27976);
xor U28742 (N_28742,N_28139,N_28181);
nand U28743 (N_28743,N_27692,N_28176);
nor U28744 (N_28744,N_27819,N_27707);
or U28745 (N_28745,N_27768,N_27988);
or U28746 (N_28746,N_27664,N_27982);
and U28747 (N_28747,N_27932,N_27674);
nand U28748 (N_28748,N_27648,N_27723);
and U28749 (N_28749,N_28146,N_27977);
xnor U28750 (N_28750,N_27733,N_28161);
nand U28751 (N_28751,N_27971,N_27905);
or U28752 (N_28752,N_27945,N_27775);
xnor U28753 (N_28753,N_28056,N_27611);
and U28754 (N_28754,N_28121,N_27999);
nand U28755 (N_28755,N_27899,N_27873);
nand U28756 (N_28756,N_27751,N_27602);
nand U28757 (N_28757,N_27615,N_27833);
nand U28758 (N_28758,N_28051,N_28096);
xor U28759 (N_28759,N_27902,N_28102);
nand U28760 (N_28760,N_28162,N_27891);
nand U28761 (N_28761,N_27983,N_27680);
nand U28762 (N_28762,N_27668,N_28189);
xnor U28763 (N_28763,N_28174,N_27962);
or U28764 (N_28764,N_28134,N_27975);
nor U28765 (N_28765,N_28082,N_27695);
xor U28766 (N_28766,N_27807,N_28121);
or U28767 (N_28767,N_27623,N_28176);
and U28768 (N_28768,N_27957,N_27948);
xnor U28769 (N_28769,N_27925,N_27960);
or U28770 (N_28770,N_27618,N_28094);
or U28771 (N_28771,N_27850,N_28170);
xnor U28772 (N_28772,N_27863,N_27905);
nor U28773 (N_28773,N_28095,N_27688);
and U28774 (N_28774,N_28138,N_27872);
and U28775 (N_28775,N_27788,N_28168);
or U28776 (N_28776,N_27659,N_27992);
nand U28777 (N_28777,N_28172,N_28177);
xnor U28778 (N_28778,N_27742,N_27889);
and U28779 (N_28779,N_27785,N_27946);
or U28780 (N_28780,N_28114,N_28044);
nand U28781 (N_28781,N_27678,N_28176);
nand U28782 (N_28782,N_27940,N_27911);
or U28783 (N_28783,N_28139,N_27777);
nand U28784 (N_28784,N_27931,N_27876);
nand U28785 (N_28785,N_27997,N_28163);
nor U28786 (N_28786,N_27891,N_28037);
and U28787 (N_28787,N_28115,N_28092);
xor U28788 (N_28788,N_27849,N_28067);
xor U28789 (N_28789,N_27858,N_27608);
xor U28790 (N_28790,N_28017,N_27719);
nor U28791 (N_28791,N_28023,N_27671);
and U28792 (N_28792,N_27750,N_28079);
or U28793 (N_28793,N_27886,N_27866);
nand U28794 (N_28794,N_27910,N_27788);
xor U28795 (N_28795,N_27960,N_27980);
and U28796 (N_28796,N_27811,N_27984);
nand U28797 (N_28797,N_27708,N_28089);
nand U28798 (N_28798,N_28034,N_27656);
nand U28799 (N_28799,N_27881,N_27834);
and U28800 (N_28800,N_28248,N_28218);
xor U28801 (N_28801,N_28700,N_28259);
nand U28802 (N_28802,N_28616,N_28471);
nor U28803 (N_28803,N_28544,N_28463);
and U28804 (N_28804,N_28222,N_28518);
nor U28805 (N_28805,N_28573,N_28457);
nor U28806 (N_28806,N_28357,N_28365);
and U28807 (N_28807,N_28462,N_28226);
or U28808 (N_28808,N_28456,N_28385);
or U28809 (N_28809,N_28234,N_28630);
xor U28810 (N_28810,N_28346,N_28246);
xor U28811 (N_28811,N_28697,N_28516);
nor U28812 (N_28812,N_28481,N_28470);
xnor U28813 (N_28813,N_28599,N_28354);
and U28814 (N_28814,N_28423,N_28653);
or U28815 (N_28815,N_28435,N_28276);
nor U28816 (N_28816,N_28403,N_28310);
and U28817 (N_28817,N_28535,N_28672);
nand U28818 (N_28818,N_28315,N_28676);
or U28819 (N_28819,N_28364,N_28461);
and U28820 (N_28820,N_28796,N_28320);
or U28821 (N_28821,N_28640,N_28603);
xor U28822 (N_28822,N_28378,N_28638);
and U28823 (N_28823,N_28433,N_28398);
and U28824 (N_28824,N_28719,N_28636);
and U28825 (N_28825,N_28339,N_28219);
nor U28826 (N_28826,N_28379,N_28537);
nand U28827 (N_28827,N_28655,N_28479);
nand U28828 (N_28828,N_28529,N_28656);
nand U28829 (N_28829,N_28352,N_28689);
or U28830 (N_28830,N_28284,N_28313);
and U28831 (N_28831,N_28411,N_28649);
or U28832 (N_28832,N_28717,N_28414);
nand U28833 (N_28833,N_28244,N_28415);
nand U28834 (N_28834,N_28644,N_28776);
and U28835 (N_28835,N_28793,N_28685);
or U28836 (N_28836,N_28232,N_28449);
xor U28837 (N_28837,N_28279,N_28269);
nand U28838 (N_28838,N_28560,N_28637);
nand U28839 (N_28839,N_28517,N_28278);
or U28840 (N_28840,N_28239,N_28798);
nand U28841 (N_28841,N_28646,N_28382);
nor U28842 (N_28842,N_28417,N_28487);
and U28843 (N_28843,N_28266,N_28448);
or U28844 (N_28844,N_28250,N_28628);
or U28845 (N_28845,N_28416,N_28549);
and U28846 (N_28846,N_28752,N_28621);
or U28847 (N_28847,N_28595,N_28677);
xor U28848 (N_28848,N_28579,N_28767);
nor U28849 (N_28849,N_28572,N_28442);
nor U28850 (N_28850,N_28237,N_28756);
or U28851 (N_28851,N_28615,N_28682);
or U28852 (N_28852,N_28273,N_28507);
nand U28853 (N_28853,N_28316,N_28439);
nand U28854 (N_28854,N_28701,N_28418);
xor U28855 (N_28855,N_28642,N_28657);
and U28856 (N_28856,N_28243,N_28691);
or U28857 (N_28857,N_28305,N_28376);
nor U28858 (N_28858,N_28247,N_28394);
nor U28859 (N_28859,N_28726,N_28265);
and U28860 (N_28860,N_28440,N_28718);
nand U28861 (N_28861,N_28614,N_28322);
and U28862 (N_28862,N_28527,N_28478);
or U28863 (N_28863,N_28738,N_28468);
or U28864 (N_28864,N_28585,N_28289);
nand U28865 (N_28865,N_28400,N_28610);
and U28866 (N_28866,N_28778,N_28304);
and U28867 (N_28867,N_28201,N_28623);
nand U28868 (N_28868,N_28356,N_28667);
nor U28869 (N_28869,N_28256,N_28594);
and U28870 (N_28870,N_28762,N_28748);
nor U28871 (N_28871,N_28741,N_28484);
xnor U28872 (N_28872,N_28542,N_28450);
nor U28873 (N_28873,N_28396,N_28625);
or U28874 (N_28874,N_28541,N_28522);
and U28875 (N_28875,N_28482,N_28713);
and U28876 (N_28876,N_28794,N_28770);
xnor U28877 (N_28877,N_28506,N_28591);
xor U28878 (N_28878,N_28298,N_28792);
xnor U28879 (N_28879,N_28598,N_28335);
nand U28880 (N_28880,N_28508,N_28592);
nand U28881 (N_28881,N_28200,N_28733);
or U28882 (N_28882,N_28659,N_28410);
nor U28883 (N_28883,N_28675,N_28486);
xnor U28884 (N_28884,N_28582,N_28721);
xnor U28885 (N_28885,N_28391,N_28458);
nand U28886 (N_28886,N_28539,N_28510);
nand U28887 (N_28887,N_28281,N_28765);
and U28888 (N_28888,N_28779,N_28781);
or U28889 (N_28889,N_28453,N_28784);
nand U28890 (N_28890,N_28734,N_28666);
nand U28891 (N_28891,N_28375,N_28326);
xor U28892 (N_28892,N_28493,N_28472);
xnor U28893 (N_28893,N_28584,N_28251);
xnor U28894 (N_28894,N_28673,N_28498);
or U28895 (N_28895,N_28570,N_28490);
nor U28896 (N_28896,N_28325,N_28344);
xor U28897 (N_28897,N_28631,N_28447);
or U28898 (N_28898,N_28710,N_28728);
or U28899 (N_28899,N_28695,N_28446);
and U28900 (N_28900,N_28746,N_28562);
nand U28901 (N_28901,N_28236,N_28451);
or U28902 (N_28902,N_28327,N_28212);
xnor U28903 (N_28903,N_28293,N_28301);
xor U28904 (N_28904,N_28687,N_28291);
nand U28905 (N_28905,N_28773,N_28750);
nand U28906 (N_28906,N_28477,N_28368);
and U28907 (N_28907,N_28359,N_28377);
xor U28908 (N_28908,N_28207,N_28314);
nand U28909 (N_28909,N_28208,N_28264);
nor U28910 (N_28910,N_28520,N_28564);
and U28911 (N_28911,N_28330,N_28569);
xnor U28912 (N_28912,N_28438,N_28413);
and U28913 (N_28913,N_28611,N_28465);
nor U28914 (N_28914,N_28645,N_28679);
xnor U28915 (N_28915,N_28495,N_28589);
nor U28916 (N_28916,N_28663,N_28312);
xor U28917 (N_28917,N_28559,N_28566);
nand U28918 (N_28918,N_28369,N_28443);
xnor U28919 (N_28919,N_28780,N_28683);
nand U28920 (N_28920,N_28308,N_28355);
nor U28921 (N_28921,N_28534,N_28612);
nand U28922 (N_28922,N_28704,N_28720);
xor U28923 (N_28923,N_28444,N_28543);
nand U28924 (N_28924,N_28419,N_28736);
and U28925 (N_28925,N_28488,N_28651);
nand U28926 (N_28926,N_28300,N_28380);
and U28927 (N_28927,N_28350,N_28709);
nor U28928 (N_28928,N_28661,N_28262);
and U28929 (N_28929,N_28753,N_28577);
and U28930 (N_28930,N_28593,N_28228);
and U28931 (N_28931,N_28530,N_28771);
nand U28932 (N_28932,N_28452,N_28641);
or U28933 (N_28933,N_28213,N_28277);
nand U28934 (N_28934,N_28786,N_28216);
and U28935 (N_28935,N_28430,N_28287);
nand U28936 (N_28936,N_28203,N_28370);
and U28937 (N_28937,N_28760,N_28501);
or U28938 (N_28938,N_28583,N_28204);
or U28939 (N_28939,N_28619,N_28723);
nor U28940 (N_28940,N_28608,N_28575);
nor U28941 (N_28941,N_28241,N_28514);
nand U28942 (N_28942,N_28703,N_28654);
nand U28943 (N_28943,N_28388,N_28509);
xnor U28944 (N_28944,N_28217,N_28282);
xor U28945 (N_28945,N_28735,N_28263);
and U28946 (N_28946,N_28513,N_28684);
nor U28947 (N_28947,N_28749,N_28702);
nand U28948 (N_28948,N_28521,N_28397);
nand U28949 (N_28949,N_28650,N_28597);
xnor U28950 (N_28950,N_28620,N_28693);
and U28951 (N_28951,N_28245,N_28604);
xor U28952 (N_28952,N_28681,N_28280);
and U28953 (N_28953,N_28406,N_28485);
xor U28954 (N_28954,N_28764,N_28393);
or U28955 (N_28955,N_28224,N_28260);
and U28956 (N_28956,N_28674,N_28774);
xnor U28957 (N_28957,N_28600,N_28613);
and U28958 (N_28958,N_28240,N_28363);
nand U28959 (N_28959,N_28574,N_28639);
nand U28960 (N_28960,N_28412,N_28275);
nand U28961 (N_28961,N_28540,N_28292);
or U28962 (N_28962,N_28739,N_28769);
and U28963 (N_28963,N_28747,N_28554);
nor U28964 (N_28964,N_28556,N_28341);
xnor U28965 (N_28965,N_28467,N_28775);
or U28966 (N_28966,N_28751,N_28519);
or U28967 (N_28967,N_28669,N_28587);
and U28968 (N_28968,N_28688,N_28311);
nor U28969 (N_28969,N_28629,N_28571);
xnor U28970 (N_28970,N_28712,N_28288);
or U28971 (N_28971,N_28231,N_28635);
nor U28972 (N_28972,N_28420,N_28602);
nor U28973 (N_28973,N_28626,N_28249);
nor U28974 (N_28974,N_28445,N_28757);
and U28975 (N_28975,N_28353,N_28694);
nand U28976 (N_28976,N_28550,N_28286);
and U28977 (N_28977,N_28758,N_28772);
nor U28978 (N_28978,N_28297,N_28730);
nor U28979 (N_28979,N_28727,N_28362);
and U28980 (N_28980,N_28267,N_28551);
nor U28981 (N_28981,N_28425,N_28404);
nor U28982 (N_28982,N_28253,N_28221);
nor U28983 (N_28983,N_28586,N_28696);
and U28984 (N_28984,N_28624,N_28399);
or U28985 (N_28985,N_28743,N_28555);
nand U28986 (N_28986,N_28329,N_28690);
or U28987 (N_28987,N_28557,N_28206);
xnor U28988 (N_28988,N_28783,N_28483);
and U28989 (N_28989,N_28324,N_28337);
or U28990 (N_28990,N_28523,N_28607);
xor U28991 (N_28991,N_28214,N_28464);
nor U28992 (N_28992,N_28223,N_28525);
and U28993 (N_28993,N_28791,N_28496);
nand U28994 (N_28994,N_28536,N_28790);
or U28995 (N_28995,N_28489,N_28383);
and U28996 (N_28996,N_28401,N_28515);
or U28997 (N_28997,N_28548,N_28622);
nor U28998 (N_28998,N_28617,N_28428);
nor U28999 (N_28999,N_28524,N_28671);
and U29000 (N_29000,N_28565,N_28306);
nand U29001 (N_29001,N_28272,N_28205);
or U29002 (N_29002,N_28561,N_28553);
or U29003 (N_29003,N_28295,N_28227);
nor U29004 (N_29004,N_28552,N_28680);
nor U29005 (N_29005,N_28705,N_28698);
or U29006 (N_29006,N_28349,N_28634);
xnor U29007 (N_29007,N_28707,N_28299);
and U29008 (N_29008,N_28437,N_28643);
and U29009 (N_29009,N_28563,N_28390);
and U29010 (N_29010,N_28725,N_28469);
and U29011 (N_29011,N_28497,N_28254);
nor U29012 (N_29012,N_28699,N_28788);
and U29013 (N_29013,N_28601,N_28371);
and U29014 (N_29014,N_28426,N_28670);
nand U29015 (N_29015,N_28480,N_28476);
nand U29016 (N_29016,N_28242,N_28233);
xor U29017 (N_29017,N_28652,N_28658);
nand U29018 (N_29018,N_28381,N_28332);
or U29019 (N_29019,N_28545,N_28348);
and U29020 (N_29020,N_28318,N_28309);
nand U29021 (N_29021,N_28590,N_28473);
nand U29022 (N_29022,N_28504,N_28323);
or U29023 (N_29023,N_28334,N_28294);
and U29024 (N_29024,N_28303,N_28210);
nand U29025 (N_29025,N_28512,N_28302);
xnor U29026 (N_29026,N_28460,N_28567);
xor U29027 (N_29027,N_28366,N_28538);
nand U29028 (N_29028,N_28714,N_28787);
xor U29029 (N_29029,N_28405,N_28706);
nor U29030 (N_29030,N_28209,N_28492);
nand U29031 (N_29031,N_28494,N_28715);
and U29032 (N_29032,N_28374,N_28795);
nor U29033 (N_29033,N_28409,N_28268);
nor U29034 (N_29034,N_28660,N_28424);
nor U29035 (N_29035,N_28716,N_28402);
and U29036 (N_29036,N_28441,N_28474);
or U29037 (N_29037,N_28692,N_28580);
nand U29038 (N_29038,N_28768,N_28220);
or U29039 (N_29039,N_28358,N_28336);
or U29040 (N_29040,N_28503,N_28296);
nor U29041 (N_29041,N_28576,N_28459);
and U29042 (N_29042,N_28202,N_28340);
xor U29043 (N_29043,N_28526,N_28648);
and U29044 (N_29044,N_28475,N_28215);
and U29045 (N_29045,N_28799,N_28547);
xnor U29046 (N_29046,N_28686,N_28427);
nand U29047 (N_29047,N_28317,N_28389);
nand U29048 (N_29048,N_28434,N_28533);
nand U29049 (N_29049,N_28499,N_28285);
nand U29050 (N_29050,N_28627,N_28407);
and U29051 (N_29051,N_28283,N_28745);
and U29052 (N_29052,N_28664,N_28491);
or U29053 (N_29053,N_28436,N_28347);
or U29054 (N_29054,N_28605,N_28319);
nand U29055 (N_29055,N_28722,N_28731);
nor U29056 (N_29056,N_28274,N_28258);
nand U29057 (N_29057,N_28454,N_28588);
xor U29058 (N_29058,N_28421,N_28392);
or U29059 (N_29059,N_28455,N_28647);
nand U29060 (N_29060,N_28331,N_28606);
xor U29061 (N_29061,N_28343,N_28367);
nor U29062 (N_29062,N_28797,N_28581);
nor U29063 (N_29063,N_28785,N_28395);
or U29064 (N_29064,N_28257,N_28729);
and U29065 (N_29065,N_28351,N_28338);
nor U29066 (N_29066,N_28384,N_28737);
or U29067 (N_29067,N_28238,N_28678);
and U29068 (N_29068,N_28408,N_28500);
xor U29069 (N_29069,N_28225,N_28789);
nor U29070 (N_29070,N_28307,N_28235);
nand U29071 (N_29071,N_28252,N_28744);
nor U29072 (N_29072,N_28290,N_28270);
xnor U29073 (N_29073,N_28766,N_28665);
xnor U29074 (N_29074,N_28777,N_28568);
xor U29075 (N_29075,N_28466,N_28361);
or U29076 (N_29076,N_28229,N_28230);
nand U29077 (N_29077,N_28321,N_28782);
nand U29078 (N_29078,N_28546,N_28373);
nand U29079 (N_29079,N_28271,N_28431);
and U29080 (N_29080,N_28261,N_28432);
and U29081 (N_29081,N_28558,N_28711);
nand U29082 (N_29082,N_28761,N_28724);
nor U29083 (N_29083,N_28531,N_28342);
nand U29084 (N_29084,N_28511,N_28360);
xor U29085 (N_29085,N_28532,N_28372);
nor U29086 (N_29086,N_28609,N_28732);
nand U29087 (N_29087,N_28755,N_28578);
xor U29088 (N_29088,N_28740,N_28632);
or U29089 (N_29089,N_28668,N_28759);
or U29090 (N_29090,N_28333,N_28596);
nand U29091 (N_29091,N_28633,N_28505);
xnor U29092 (N_29092,N_28708,N_28422);
xor U29093 (N_29093,N_28754,N_28386);
xnor U29094 (N_29094,N_28528,N_28429);
nand U29095 (N_29095,N_28618,N_28255);
nor U29096 (N_29096,N_28763,N_28742);
and U29097 (N_29097,N_28387,N_28345);
xnor U29098 (N_29098,N_28211,N_28662);
nor U29099 (N_29099,N_28502,N_28328);
nor U29100 (N_29100,N_28268,N_28615);
and U29101 (N_29101,N_28596,N_28726);
nor U29102 (N_29102,N_28259,N_28227);
and U29103 (N_29103,N_28580,N_28670);
nor U29104 (N_29104,N_28678,N_28221);
nand U29105 (N_29105,N_28640,N_28271);
and U29106 (N_29106,N_28721,N_28779);
xor U29107 (N_29107,N_28475,N_28216);
nand U29108 (N_29108,N_28711,N_28435);
and U29109 (N_29109,N_28386,N_28439);
nand U29110 (N_29110,N_28557,N_28292);
nand U29111 (N_29111,N_28568,N_28483);
and U29112 (N_29112,N_28379,N_28247);
nand U29113 (N_29113,N_28249,N_28276);
nor U29114 (N_29114,N_28436,N_28319);
xor U29115 (N_29115,N_28214,N_28756);
nor U29116 (N_29116,N_28246,N_28558);
xnor U29117 (N_29117,N_28418,N_28523);
and U29118 (N_29118,N_28626,N_28603);
and U29119 (N_29119,N_28578,N_28314);
and U29120 (N_29120,N_28225,N_28211);
xnor U29121 (N_29121,N_28573,N_28756);
or U29122 (N_29122,N_28609,N_28527);
xnor U29123 (N_29123,N_28650,N_28706);
xnor U29124 (N_29124,N_28470,N_28701);
nand U29125 (N_29125,N_28484,N_28637);
xnor U29126 (N_29126,N_28696,N_28305);
xor U29127 (N_29127,N_28363,N_28241);
nor U29128 (N_29128,N_28408,N_28598);
or U29129 (N_29129,N_28390,N_28519);
or U29130 (N_29130,N_28219,N_28796);
nand U29131 (N_29131,N_28686,N_28517);
nor U29132 (N_29132,N_28300,N_28389);
xor U29133 (N_29133,N_28617,N_28229);
nor U29134 (N_29134,N_28714,N_28607);
or U29135 (N_29135,N_28603,N_28435);
nor U29136 (N_29136,N_28494,N_28565);
nand U29137 (N_29137,N_28717,N_28483);
or U29138 (N_29138,N_28517,N_28604);
and U29139 (N_29139,N_28625,N_28311);
and U29140 (N_29140,N_28743,N_28247);
or U29141 (N_29141,N_28697,N_28373);
or U29142 (N_29142,N_28420,N_28571);
nand U29143 (N_29143,N_28259,N_28360);
nand U29144 (N_29144,N_28204,N_28330);
or U29145 (N_29145,N_28612,N_28337);
or U29146 (N_29146,N_28638,N_28553);
xnor U29147 (N_29147,N_28525,N_28683);
xnor U29148 (N_29148,N_28492,N_28691);
xor U29149 (N_29149,N_28253,N_28299);
nand U29150 (N_29150,N_28504,N_28269);
nand U29151 (N_29151,N_28543,N_28713);
or U29152 (N_29152,N_28554,N_28274);
nand U29153 (N_29153,N_28746,N_28661);
or U29154 (N_29154,N_28349,N_28571);
nand U29155 (N_29155,N_28206,N_28440);
nand U29156 (N_29156,N_28434,N_28275);
and U29157 (N_29157,N_28670,N_28288);
nand U29158 (N_29158,N_28627,N_28462);
nor U29159 (N_29159,N_28576,N_28416);
nand U29160 (N_29160,N_28522,N_28215);
nor U29161 (N_29161,N_28693,N_28436);
and U29162 (N_29162,N_28480,N_28464);
xnor U29163 (N_29163,N_28787,N_28779);
nand U29164 (N_29164,N_28277,N_28792);
and U29165 (N_29165,N_28445,N_28475);
nand U29166 (N_29166,N_28451,N_28400);
and U29167 (N_29167,N_28575,N_28410);
or U29168 (N_29168,N_28355,N_28353);
nor U29169 (N_29169,N_28376,N_28356);
or U29170 (N_29170,N_28486,N_28364);
nand U29171 (N_29171,N_28585,N_28707);
nand U29172 (N_29172,N_28221,N_28390);
xor U29173 (N_29173,N_28686,N_28229);
or U29174 (N_29174,N_28648,N_28222);
nand U29175 (N_29175,N_28201,N_28359);
xor U29176 (N_29176,N_28336,N_28330);
nand U29177 (N_29177,N_28778,N_28583);
nand U29178 (N_29178,N_28771,N_28684);
xnor U29179 (N_29179,N_28566,N_28273);
xnor U29180 (N_29180,N_28270,N_28253);
or U29181 (N_29181,N_28568,N_28369);
and U29182 (N_29182,N_28205,N_28519);
nand U29183 (N_29183,N_28592,N_28363);
nand U29184 (N_29184,N_28745,N_28227);
or U29185 (N_29185,N_28796,N_28730);
nand U29186 (N_29186,N_28658,N_28428);
nand U29187 (N_29187,N_28390,N_28341);
nand U29188 (N_29188,N_28477,N_28656);
or U29189 (N_29189,N_28752,N_28662);
and U29190 (N_29190,N_28248,N_28300);
xnor U29191 (N_29191,N_28471,N_28457);
or U29192 (N_29192,N_28682,N_28316);
nand U29193 (N_29193,N_28283,N_28576);
nor U29194 (N_29194,N_28584,N_28256);
nand U29195 (N_29195,N_28577,N_28630);
or U29196 (N_29196,N_28709,N_28342);
or U29197 (N_29197,N_28768,N_28481);
and U29198 (N_29198,N_28336,N_28590);
xnor U29199 (N_29199,N_28313,N_28265);
nor U29200 (N_29200,N_28694,N_28468);
or U29201 (N_29201,N_28738,N_28799);
or U29202 (N_29202,N_28705,N_28241);
or U29203 (N_29203,N_28468,N_28556);
nand U29204 (N_29204,N_28575,N_28484);
xnor U29205 (N_29205,N_28567,N_28269);
xnor U29206 (N_29206,N_28458,N_28598);
nor U29207 (N_29207,N_28620,N_28622);
and U29208 (N_29208,N_28310,N_28424);
and U29209 (N_29209,N_28550,N_28391);
and U29210 (N_29210,N_28750,N_28253);
nor U29211 (N_29211,N_28787,N_28342);
or U29212 (N_29212,N_28203,N_28218);
and U29213 (N_29213,N_28776,N_28539);
xnor U29214 (N_29214,N_28413,N_28381);
nand U29215 (N_29215,N_28236,N_28361);
or U29216 (N_29216,N_28348,N_28423);
and U29217 (N_29217,N_28498,N_28403);
and U29218 (N_29218,N_28381,N_28628);
xor U29219 (N_29219,N_28667,N_28694);
and U29220 (N_29220,N_28520,N_28536);
xor U29221 (N_29221,N_28348,N_28265);
and U29222 (N_29222,N_28794,N_28623);
xor U29223 (N_29223,N_28460,N_28403);
nor U29224 (N_29224,N_28256,N_28553);
and U29225 (N_29225,N_28591,N_28789);
xnor U29226 (N_29226,N_28534,N_28475);
xnor U29227 (N_29227,N_28690,N_28363);
and U29228 (N_29228,N_28476,N_28429);
and U29229 (N_29229,N_28443,N_28250);
and U29230 (N_29230,N_28534,N_28213);
or U29231 (N_29231,N_28377,N_28764);
and U29232 (N_29232,N_28689,N_28264);
and U29233 (N_29233,N_28660,N_28591);
or U29234 (N_29234,N_28722,N_28692);
nor U29235 (N_29235,N_28686,N_28238);
nor U29236 (N_29236,N_28713,N_28269);
and U29237 (N_29237,N_28411,N_28767);
nor U29238 (N_29238,N_28200,N_28755);
nor U29239 (N_29239,N_28792,N_28761);
xnor U29240 (N_29240,N_28377,N_28423);
nor U29241 (N_29241,N_28315,N_28641);
and U29242 (N_29242,N_28648,N_28540);
xor U29243 (N_29243,N_28534,N_28640);
nand U29244 (N_29244,N_28703,N_28765);
nor U29245 (N_29245,N_28218,N_28401);
nor U29246 (N_29246,N_28782,N_28617);
nand U29247 (N_29247,N_28385,N_28715);
xnor U29248 (N_29248,N_28517,N_28414);
nand U29249 (N_29249,N_28646,N_28207);
nand U29250 (N_29250,N_28718,N_28790);
xnor U29251 (N_29251,N_28409,N_28399);
or U29252 (N_29252,N_28624,N_28687);
and U29253 (N_29253,N_28400,N_28233);
and U29254 (N_29254,N_28389,N_28794);
or U29255 (N_29255,N_28574,N_28521);
xnor U29256 (N_29256,N_28259,N_28235);
nand U29257 (N_29257,N_28550,N_28707);
xnor U29258 (N_29258,N_28717,N_28793);
nor U29259 (N_29259,N_28778,N_28681);
nor U29260 (N_29260,N_28664,N_28628);
and U29261 (N_29261,N_28633,N_28663);
xor U29262 (N_29262,N_28551,N_28700);
and U29263 (N_29263,N_28419,N_28524);
and U29264 (N_29264,N_28459,N_28254);
nor U29265 (N_29265,N_28351,N_28645);
nand U29266 (N_29266,N_28555,N_28376);
or U29267 (N_29267,N_28235,N_28686);
xnor U29268 (N_29268,N_28294,N_28471);
nor U29269 (N_29269,N_28650,N_28327);
xor U29270 (N_29270,N_28265,N_28398);
nor U29271 (N_29271,N_28798,N_28366);
and U29272 (N_29272,N_28433,N_28534);
and U29273 (N_29273,N_28687,N_28596);
nand U29274 (N_29274,N_28631,N_28674);
or U29275 (N_29275,N_28415,N_28436);
xor U29276 (N_29276,N_28760,N_28704);
xnor U29277 (N_29277,N_28394,N_28747);
xor U29278 (N_29278,N_28792,N_28422);
or U29279 (N_29279,N_28530,N_28339);
or U29280 (N_29280,N_28545,N_28470);
and U29281 (N_29281,N_28482,N_28205);
and U29282 (N_29282,N_28292,N_28718);
nand U29283 (N_29283,N_28214,N_28290);
and U29284 (N_29284,N_28370,N_28460);
nand U29285 (N_29285,N_28217,N_28391);
nand U29286 (N_29286,N_28264,N_28532);
or U29287 (N_29287,N_28337,N_28439);
xnor U29288 (N_29288,N_28646,N_28202);
and U29289 (N_29289,N_28400,N_28659);
and U29290 (N_29290,N_28556,N_28541);
and U29291 (N_29291,N_28235,N_28608);
nand U29292 (N_29292,N_28790,N_28496);
nor U29293 (N_29293,N_28532,N_28714);
nand U29294 (N_29294,N_28487,N_28443);
nand U29295 (N_29295,N_28760,N_28691);
and U29296 (N_29296,N_28509,N_28524);
nand U29297 (N_29297,N_28324,N_28604);
or U29298 (N_29298,N_28783,N_28633);
or U29299 (N_29299,N_28503,N_28300);
or U29300 (N_29300,N_28765,N_28715);
xor U29301 (N_29301,N_28494,N_28457);
or U29302 (N_29302,N_28326,N_28335);
nand U29303 (N_29303,N_28351,N_28553);
nand U29304 (N_29304,N_28464,N_28732);
and U29305 (N_29305,N_28742,N_28708);
xor U29306 (N_29306,N_28463,N_28610);
xnor U29307 (N_29307,N_28478,N_28306);
nand U29308 (N_29308,N_28708,N_28596);
nand U29309 (N_29309,N_28392,N_28358);
xor U29310 (N_29310,N_28286,N_28622);
xor U29311 (N_29311,N_28444,N_28437);
or U29312 (N_29312,N_28436,N_28763);
or U29313 (N_29313,N_28398,N_28683);
xnor U29314 (N_29314,N_28652,N_28436);
nor U29315 (N_29315,N_28508,N_28511);
or U29316 (N_29316,N_28265,N_28268);
and U29317 (N_29317,N_28655,N_28315);
or U29318 (N_29318,N_28627,N_28441);
nor U29319 (N_29319,N_28207,N_28525);
or U29320 (N_29320,N_28629,N_28542);
nor U29321 (N_29321,N_28776,N_28502);
or U29322 (N_29322,N_28354,N_28783);
and U29323 (N_29323,N_28448,N_28473);
or U29324 (N_29324,N_28728,N_28228);
or U29325 (N_29325,N_28455,N_28279);
nor U29326 (N_29326,N_28351,N_28262);
xnor U29327 (N_29327,N_28673,N_28200);
xor U29328 (N_29328,N_28222,N_28512);
and U29329 (N_29329,N_28770,N_28469);
xnor U29330 (N_29330,N_28290,N_28210);
and U29331 (N_29331,N_28712,N_28574);
nand U29332 (N_29332,N_28479,N_28410);
nand U29333 (N_29333,N_28291,N_28667);
xor U29334 (N_29334,N_28700,N_28742);
nand U29335 (N_29335,N_28778,N_28781);
nand U29336 (N_29336,N_28549,N_28391);
and U29337 (N_29337,N_28225,N_28726);
nand U29338 (N_29338,N_28333,N_28580);
nor U29339 (N_29339,N_28718,N_28702);
and U29340 (N_29340,N_28345,N_28551);
nor U29341 (N_29341,N_28544,N_28356);
or U29342 (N_29342,N_28240,N_28764);
and U29343 (N_29343,N_28564,N_28357);
nand U29344 (N_29344,N_28713,N_28667);
and U29345 (N_29345,N_28592,N_28693);
nor U29346 (N_29346,N_28229,N_28610);
and U29347 (N_29347,N_28360,N_28581);
and U29348 (N_29348,N_28479,N_28477);
xnor U29349 (N_29349,N_28367,N_28570);
xnor U29350 (N_29350,N_28761,N_28604);
and U29351 (N_29351,N_28558,N_28202);
nand U29352 (N_29352,N_28336,N_28770);
nor U29353 (N_29353,N_28537,N_28682);
or U29354 (N_29354,N_28796,N_28490);
xor U29355 (N_29355,N_28463,N_28264);
and U29356 (N_29356,N_28306,N_28207);
xor U29357 (N_29357,N_28283,N_28629);
xnor U29358 (N_29358,N_28634,N_28475);
xor U29359 (N_29359,N_28702,N_28365);
nor U29360 (N_29360,N_28749,N_28306);
xnor U29361 (N_29361,N_28366,N_28584);
or U29362 (N_29362,N_28448,N_28641);
xor U29363 (N_29363,N_28225,N_28560);
and U29364 (N_29364,N_28587,N_28354);
nand U29365 (N_29365,N_28540,N_28785);
nor U29366 (N_29366,N_28571,N_28683);
and U29367 (N_29367,N_28708,N_28711);
xnor U29368 (N_29368,N_28757,N_28357);
or U29369 (N_29369,N_28400,N_28739);
nand U29370 (N_29370,N_28290,N_28220);
or U29371 (N_29371,N_28587,N_28715);
or U29372 (N_29372,N_28656,N_28243);
and U29373 (N_29373,N_28658,N_28276);
nor U29374 (N_29374,N_28596,N_28791);
nand U29375 (N_29375,N_28476,N_28313);
nor U29376 (N_29376,N_28483,N_28795);
nand U29377 (N_29377,N_28510,N_28361);
nand U29378 (N_29378,N_28695,N_28457);
nand U29379 (N_29379,N_28208,N_28673);
and U29380 (N_29380,N_28464,N_28451);
xor U29381 (N_29381,N_28302,N_28401);
and U29382 (N_29382,N_28520,N_28665);
xnor U29383 (N_29383,N_28647,N_28303);
or U29384 (N_29384,N_28642,N_28508);
xor U29385 (N_29385,N_28393,N_28367);
nor U29386 (N_29386,N_28263,N_28553);
or U29387 (N_29387,N_28272,N_28284);
xnor U29388 (N_29388,N_28564,N_28779);
or U29389 (N_29389,N_28381,N_28715);
and U29390 (N_29390,N_28295,N_28483);
and U29391 (N_29391,N_28639,N_28769);
and U29392 (N_29392,N_28667,N_28669);
and U29393 (N_29393,N_28485,N_28386);
or U29394 (N_29394,N_28701,N_28420);
or U29395 (N_29395,N_28329,N_28581);
nand U29396 (N_29396,N_28308,N_28613);
nor U29397 (N_29397,N_28623,N_28542);
xnor U29398 (N_29398,N_28337,N_28248);
nand U29399 (N_29399,N_28411,N_28264);
xor U29400 (N_29400,N_28939,N_29167);
xor U29401 (N_29401,N_29259,N_28822);
xor U29402 (N_29402,N_29123,N_28920);
and U29403 (N_29403,N_29367,N_28942);
and U29404 (N_29404,N_29197,N_29256);
nor U29405 (N_29405,N_28834,N_28820);
nor U29406 (N_29406,N_29299,N_29345);
xor U29407 (N_29407,N_29108,N_29059);
xnor U29408 (N_29408,N_29229,N_29304);
nand U29409 (N_29409,N_29322,N_29252);
and U29410 (N_29410,N_29276,N_28861);
or U29411 (N_29411,N_29190,N_29036);
nor U29412 (N_29412,N_29370,N_29395);
and U29413 (N_29413,N_29151,N_29332);
nor U29414 (N_29414,N_29101,N_29194);
xor U29415 (N_29415,N_29185,N_29318);
nand U29416 (N_29416,N_28848,N_29231);
nor U29417 (N_29417,N_29355,N_28971);
and U29418 (N_29418,N_28851,N_28804);
xor U29419 (N_29419,N_29088,N_29087);
nand U29420 (N_29420,N_29300,N_29090);
xnor U29421 (N_29421,N_29104,N_29075);
nand U29422 (N_29422,N_29132,N_29309);
nand U29423 (N_29423,N_29381,N_29230);
xnor U29424 (N_29424,N_29055,N_29327);
nand U29425 (N_29425,N_28972,N_29391);
or U29426 (N_29426,N_29379,N_28899);
nor U29427 (N_29427,N_29052,N_29011);
nor U29428 (N_29428,N_29107,N_28801);
nor U29429 (N_29429,N_29016,N_29095);
nand U29430 (N_29430,N_28874,N_29277);
and U29431 (N_29431,N_29296,N_28973);
and U29432 (N_29432,N_28880,N_29002);
or U29433 (N_29433,N_29266,N_29024);
and U29434 (N_29434,N_29254,N_29189);
nand U29435 (N_29435,N_28862,N_29173);
nand U29436 (N_29436,N_28875,N_28907);
nor U29437 (N_29437,N_29073,N_28877);
nand U29438 (N_29438,N_29004,N_28807);
or U29439 (N_29439,N_29098,N_29232);
or U29440 (N_29440,N_29265,N_29093);
or U29441 (N_29441,N_29294,N_28800);
or U29442 (N_29442,N_29210,N_29312);
or U29443 (N_29443,N_28889,N_29193);
or U29444 (N_29444,N_29184,N_29074);
nor U29445 (N_29445,N_29111,N_28922);
nor U29446 (N_29446,N_28918,N_28826);
nor U29447 (N_29447,N_29091,N_29100);
or U29448 (N_29448,N_28846,N_29273);
xor U29449 (N_29449,N_29140,N_29233);
nor U29450 (N_29450,N_28982,N_29067);
xnor U29451 (N_29451,N_29038,N_28878);
xor U29452 (N_29452,N_29122,N_28959);
xor U29453 (N_29453,N_29317,N_29349);
xor U29454 (N_29454,N_29076,N_28945);
nor U29455 (N_29455,N_29035,N_28984);
nor U29456 (N_29456,N_28803,N_29031);
or U29457 (N_29457,N_29378,N_29034);
xnor U29458 (N_29458,N_28926,N_29061);
or U29459 (N_29459,N_28936,N_29281);
nor U29460 (N_29460,N_28870,N_29113);
nor U29461 (N_29461,N_29267,N_29386);
nor U29462 (N_29462,N_29143,N_29160);
nand U29463 (N_29463,N_29385,N_29212);
nor U29464 (N_29464,N_29297,N_29183);
xor U29465 (N_29465,N_29343,N_29081);
or U29466 (N_29466,N_28823,N_28838);
xnor U29467 (N_29467,N_29394,N_29175);
and U29468 (N_29468,N_29338,N_29019);
or U29469 (N_29469,N_29239,N_29295);
nor U29470 (N_29470,N_28911,N_28900);
or U29471 (N_29471,N_29136,N_28888);
or U29472 (N_29472,N_29307,N_28915);
xnor U29473 (N_29473,N_28842,N_29336);
nand U29474 (N_29474,N_28953,N_29030);
nand U29475 (N_29475,N_29375,N_28975);
nand U29476 (N_29476,N_29272,N_29365);
nand U29477 (N_29477,N_28833,N_29162);
xnor U29478 (N_29478,N_28927,N_29223);
xnor U29479 (N_29479,N_29077,N_29191);
or U29480 (N_29480,N_29166,N_28892);
or U29481 (N_29481,N_28808,N_29207);
xor U29482 (N_29482,N_29199,N_29138);
nor U29483 (N_29483,N_29202,N_29020);
xor U29484 (N_29484,N_29005,N_29240);
nor U29485 (N_29485,N_28904,N_28994);
or U29486 (N_29486,N_28992,N_29171);
xnor U29487 (N_29487,N_28817,N_29124);
and U29488 (N_29488,N_29316,N_28917);
nand U29489 (N_29489,N_28980,N_28856);
xnor U29490 (N_29490,N_29397,N_29187);
nand U29491 (N_29491,N_28997,N_29085);
xnor U29492 (N_29492,N_29246,N_28932);
or U29493 (N_29493,N_29337,N_29146);
or U29494 (N_29494,N_28865,N_29017);
nor U29495 (N_29495,N_29369,N_29131);
nand U29496 (N_29496,N_29119,N_28990);
and U29497 (N_29497,N_29039,N_29248);
nand U29498 (N_29498,N_29050,N_28983);
nor U29499 (N_29499,N_28881,N_29118);
nand U29500 (N_29500,N_29195,N_28930);
or U29501 (N_29501,N_28879,N_29208);
and U29502 (N_29502,N_29065,N_29235);
and U29503 (N_29503,N_28989,N_28876);
or U29504 (N_29504,N_29319,N_28902);
and U29505 (N_29505,N_29353,N_28863);
nand U29506 (N_29506,N_29177,N_29216);
xnor U29507 (N_29507,N_29063,N_29137);
or U29508 (N_29508,N_29043,N_29116);
nor U29509 (N_29509,N_29026,N_28893);
or U29510 (N_29510,N_29109,N_28919);
nor U29511 (N_29511,N_28859,N_28993);
nand U29512 (N_29512,N_29243,N_28956);
or U29513 (N_29513,N_29310,N_29094);
nor U29514 (N_29514,N_29306,N_29023);
nand U29515 (N_29515,N_29292,N_29013);
and U29516 (N_29516,N_29279,N_29263);
nor U29517 (N_29517,N_29176,N_28961);
xor U29518 (N_29518,N_29082,N_29214);
nor U29519 (N_29519,N_29372,N_28843);
or U29520 (N_29520,N_28949,N_28837);
nand U29521 (N_29521,N_29139,N_29335);
nand U29522 (N_29522,N_29188,N_28991);
nor U29523 (N_29523,N_28966,N_29376);
and U29524 (N_29524,N_29012,N_29298);
nand U29525 (N_29525,N_28947,N_28946);
nand U29526 (N_29526,N_28940,N_28825);
or U29527 (N_29527,N_29051,N_29147);
xnor U29528 (N_29528,N_28909,N_29334);
and U29529 (N_29529,N_29333,N_28802);
nor U29530 (N_29530,N_29287,N_29383);
nand U29531 (N_29531,N_29360,N_29289);
nand U29532 (N_29532,N_29253,N_29286);
xor U29533 (N_29533,N_29371,N_29150);
nor U29534 (N_29534,N_29398,N_29225);
xnor U29535 (N_29535,N_29127,N_29149);
and U29536 (N_29536,N_29128,N_29204);
nor U29537 (N_29537,N_29224,N_28996);
and U29538 (N_29538,N_29201,N_29222);
and U29539 (N_29539,N_28806,N_29028);
and U29540 (N_29540,N_29045,N_28908);
and U29541 (N_29541,N_29303,N_29096);
nand U29542 (N_29542,N_28913,N_28855);
and U29543 (N_29543,N_29018,N_29250);
nor U29544 (N_29544,N_28955,N_28835);
nand U29545 (N_29545,N_29341,N_29182);
or U29546 (N_29546,N_29351,N_29340);
xnor U29547 (N_29547,N_29134,N_29361);
or U29548 (N_29548,N_28854,N_29206);
xnor U29549 (N_29549,N_29155,N_29288);
xor U29550 (N_29550,N_29158,N_29325);
nor U29551 (N_29551,N_29393,N_28829);
nor U29552 (N_29552,N_28978,N_28821);
nand U29553 (N_29553,N_29196,N_28934);
or U29554 (N_29554,N_29268,N_29047);
nand U29555 (N_29555,N_28832,N_28839);
and U29556 (N_29556,N_29092,N_28867);
or U29557 (N_29557,N_28809,N_29342);
or U29558 (N_29558,N_29368,N_28810);
and U29559 (N_29559,N_29220,N_29339);
xnor U29560 (N_29560,N_29257,N_28948);
or U29561 (N_29561,N_28965,N_29198);
and U29562 (N_29562,N_29211,N_29159);
xnor U29563 (N_29563,N_28905,N_29290);
nand U29564 (N_29564,N_28831,N_28818);
or U29565 (N_29565,N_29181,N_28916);
nand U29566 (N_29566,N_29130,N_29001);
nand U29567 (N_29567,N_29121,N_29086);
nand U29568 (N_29568,N_29323,N_29058);
nor U29569 (N_29569,N_29291,N_29025);
nand U29570 (N_29570,N_29314,N_29106);
or U29571 (N_29571,N_29040,N_28824);
or U29572 (N_29572,N_29064,N_29010);
nand U29573 (N_29573,N_28828,N_28985);
xnor U29574 (N_29574,N_29237,N_29331);
or U29575 (N_29575,N_28858,N_29179);
and U29576 (N_29576,N_29129,N_29359);
nor U29577 (N_29577,N_29114,N_29046);
nand U29578 (N_29578,N_28977,N_28897);
xnor U29579 (N_29579,N_29105,N_29329);
nor U29580 (N_29580,N_28873,N_29219);
and U29581 (N_29581,N_29044,N_29380);
xor U29582 (N_29582,N_29056,N_29346);
or U29583 (N_29583,N_28883,N_28937);
and U29584 (N_29584,N_29358,N_28885);
xnor U29585 (N_29585,N_29015,N_29145);
or U29586 (N_29586,N_28849,N_29362);
nand U29587 (N_29587,N_29203,N_29363);
xnor U29588 (N_29588,N_28944,N_28995);
nor U29589 (N_29589,N_29384,N_29007);
xnor U29590 (N_29590,N_28819,N_28964);
nand U29591 (N_29591,N_28884,N_28957);
nor U29592 (N_29592,N_29320,N_29260);
or U29593 (N_29593,N_29169,N_29069);
or U29594 (N_29594,N_28901,N_28841);
and U29595 (N_29595,N_28871,N_28812);
or U29596 (N_29596,N_28868,N_29174);
xor U29597 (N_29597,N_29245,N_28906);
xor U29598 (N_29598,N_28886,N_29373);
nand U29599 (N_29599,N_29102,N_29255);
and U29600 (N_29600,N_28952,N_28894);
nor U29601 (N_29601,N_29126,N_29178);
and U29602 (N_29602,N_29099,N_29070);
or U29603 (N_29603,N_29270,N_29302);
or U29604 (N_29604,N_29305,N_29165);
nand U29605 (N_29605,N_29399,N_29278);
and U29606 (N_29606,N_28853,N_29048);
nor U29607 (N_29607,N_29228,N_28872);
nor U29608 (N_29608,N_29141,N_29097);
or U29609 (N_29609,N_29008,N_29170);
nand U29610 (N_29610,N_28912,N_29071);
or U29611 (N_29611,N_29156,N_28925);
nor U29612 (N_29612,N_29258,N_29226);
nor U29613 (N_29613,N_29022,N_28988);
or U29614 (N_29614,N_28914,N_29262);
xnor U29615 (N_29615,N_28951,N_29049);
nor U29616 (N_29616,N_29120,N_28998);
xnor U29617 (N_29617,N_29072,N_29227);
and U29618 (N_29618,N_29313,N_29213);
or U29619 (N_29619,N_28827,N_29221);
nor U29620 (N_29620,N_29168,N_28847);
xor U29621 (N_29621,N_29144,N_28895);
or U29622 (N_29622,N_29110,N_29249);
and U29623 (N_29623,N_29396,N_29078);
nand U29624 (N_29624,N_29054,N_29021);
xnor U29625 (N_29625,N_29215,N_29186);
or U29626 (N_29626,N_28814,N_29135);
or U29627 (N_29627,N_28967,N_28981);
xor U29628 (N_29628,N_29163,N_28864);
nor U29629 (N_29629,N_28931,N_29366);
nand U29630 (N_29630,N_29374,N_29103);
xnor U29631 (N_29631,N_28923,N_29244);
or U29632 (N_29632,N_28921,N_28840);
nand U29633 (N_29633,N_29347,N_29387);
xnor U29634 (N_29634,N_29027,N_29115);
nand U29635 (N_29635,N_29079,N_29172);
or U29636 (N_29636,N_29157,N_29321);
and U29637 (N_29637,N_29283,N_28950);
xnor U29638 (N_29638,N_29209,N_28830);
or U29639 (N_29639,N_29032,N_29354);
xnor U29640 (N_29640,N_29200,N_29238);
xor U29641 (N_29641,N_29269,N_29348);
nand U29642 (N_29642,N_29164,N_28898);
and U29643 (N_29643,N_29392,N_28836);
nor U29644 (N_29644,N_29242,N_29041);
or U29645 (N_29645,N_29261,N_29154);
or U29646 (N_29646,N_29352,N_28968);
or U29647 (N_29647,N_28805,N_29000);
xnor U29648 (N_29648,N_29112,N_29389);
xnor U29649 (N_29649,N_29326,N_29390);
xor U29650 (N_29650,N_29060,N_29350);
or U29651 (N_29651,N_28903,N_29029);
nand U29652 (N_29652,N_28844,N_29042);
nand U29653 (N_29653,N_28815,N_28813);
xnor U29654 (N_29654,N_29125,N_29311);
xnor U29655 (N_29655,N_28935,N_28954);
xor U29656 (N_29656,N_29014,N_28943);
xnor U29657 (N_29657,N_28987,N_29037);
nor U29658 (N_29658,N_28860,N_29344);
xnor U29659 (N_29659,N_29148,N_28941);
nand U29660 (N_29660,N_29271,N_29057);
or U29661 (N_29661,N_29282,N_29161);
nor U29662 (N_29662,N_28974,N_28969);
or U29663 (N_29663,N_29284,N_29003);
nor U29664 (N_29664,N_29084,N_28928);
nor U29665 (N_29665,N_29275,N_29089);
nor U29666 (N_29666,N_29009,N_28933);
nor U29667 (N_29667,N_29308,N_28938);
and U29668 (N_29668,N_29251,N_29080);
or U29669 (N_29669,N_29315,N_29364);
nand U29670 (N_29670,N_29377,N_28962);
or U29671 (N_29671,N_28999,N_29264);
nand U29672 (N_29672,N_28960,N_29324);
nand U29673 (N_29673,N_29330,N_29217);
nand U29674 (N_29674,N_29247,N_29293);
xor U29675 (N_29675,N_29285,N_28882);
xor U29676 (N_29676,N_29066,N_29068);
nor U29677 (N_29677,N_29142,N_29234);
xnor U29678 (N_29678,N_28891,N_28979);
and U29679 (N_29679,N_28857,N_28850);
xor U29680 (N_29680,N_29180,N_29205);
or U29681 (N_29681,N_28970,N_29152);
or U29682 (N_29682,N_29280,N_28890);
or U29683 (N_29683,N_28866,N_29328);
or U29684 (N_29684,N_28986,N_29192);
or U29685 (N_29685,N_29033,N_28852);
xor U29686 (N_29686,N_28869,N_29357);
xnor U29687 (N_29687,N_28816,N_29301);
and U29688 (N_29688,N_28811,N_29153);
nor U29689 (N_29689,N_28896,N_29006);
nand U29690 (N_29690,N_28976,N_29356);
or U29691 (N_29691,N_29241,N_29274);
nor U29692 (N_29692,N_28963,N_29083);
and U29693 (N_29693,N_28958,N_29062);
or U29694 (N_29694,N_28910,N_29117);
nand U29695 (N_29695,N_28887,N_28924);
xor U29696 (N_29696,N_28929,N_29236);
xor U29697 (N_29697,N_29133,N_29053);
and U29698 (N_29698,N_29218,N_29382);
nor U29699 (N_29699,N_29388,N_28845);
and U29700 (N_29700,N_29373,N_29337);
and U29701 (N_29701,N_29007,N_28803);
xnor U29702 (N_29702,N_29237,N_28893);
or U29703 (N_29703,N_29077,N_29360);
nand U29704 (N_29704,N_29156,N_29197);
nor U29705 (N_29705,N_29301,N_29049);
xor U29706 (N_29706,N_29242,N_29097);
or U29707 (N_29707,N_28982,N_29133);
nand U29708 (N_29708,N_28853,N_28899);
nor U29709 (N_29709,N_29018,N_29150);
and U29710 (N_29710,N_29326,N_29264);
nand U29711 (N_29711,N_29032,N_29049);
nand U29712 (N_29712,N_28816,N_28837);
or U29713 (N_29713,N_29019,N_29347);
nor U29714 (N_29714,N_28821,N_29102);
nand U29715 (N_29715,N_29086,N_29292);
nor U29716 (N_29716,N_29092,N_28839);
nand U29717 (N_29717,N_29086,N_28986);
or U29718 (N_29718,N_28834,N_28852);
or U29719 (N_29719,N_29263,N_29068);
or U29720 (N_29720,N_29186,N_29169);
xnor U29721 (N_29721,N_28950,N_29290);
nor U29722 (N_29722,N_29198,N_28860);
and U29723 (N_29723,N_28929,N_29116);
nand U29724 (N_29724,N_29272,N_29063);
and U29725 (N_29725,N_29080,N_28960);
nor U29726 (N_29726,N_28939,N_29362);
xor U29727 (N_29727,N_29075,N_28890);
nor U29728 (N_29728,N_29294,N_29187);
or U29729 (N_29729,N_29165,N_29381);
nand U29730 (N_29730,N_28981,N_28859);
and U29731 (N_29731,N_29002,N_29275);
or U29732 (N_29732,N_28977,N_28959);
nor U29733 (N_29733,N_29117,N_28855);
or U29734 (N_29734,N_28817,N_29397);
xnor U29735 (N_29735,N_29319,N_29213);
nor U29736 (N_29736,N_29231,N_29196);
nor U29737 (N_29737,N_29066,N_28830);
xnor U29738 (N_29738,N_29354,N_29364);
nand U29739 (N_29739,N_28962,N_29390);
nand U29740 (N_29740,N_28863,N_29129);
nor U29741 (N_29741,N_28959,N_29364);
xnor U29742 (N_29742,N_28921,N_29064);
nor U29743 (N_29743,N_29049,N_29002);
nor U29744 (N_29744,N_29110,N_29130);
nor U29745 (N_29745,N_29161,N_28928);
nand U29746 (N_29746,N_28892,N_29220);
nor U29747 (N_29747,N_29139,N_29083);
or U29748 (N_29748,N_29068,N_29286);
xnor U29749 (N_29749,N_29391,N_28901);
xnor U29750 (N_29750,N_28864,N_29376);
nand U29751 (N_29751,N_28968,N_29335);
nand U29752 (N_29752,N_29263,N_29381);
or U29753 (N_29753,N_28838,N_29283);
and U29754 (N_29754,N_28895,N_28845);
xor U29755 (N_29755,N_29132,N_29205);
or U29756 (N_29756,N_28924,N_29045);
or U29757 (N_29757,N_29322,N_29056);
xnor U29758 (N_29758,N_28811,N_29181);
xor U29759 (N_29759,N_29359,N_29041);
nand U29760 (N_29760,N_29236,N_29266);
or U29761 (N_29761,N_28862,N_29034);
xor U29762 (N_29762,N_28907,N_28834);
nand U29763 (N_29763,N_29363,N_28994);
or U29764 (N_29764,N_29190,N_29079);
xnor U29765 (N_29765,N_29236,N_28999);
xor U29766 (N_29766,N_29054,N_28915);
xnor U29767 (N_29767,N_28924,N_29182);
or U29768 (N_29768,N_29184,N_29339);
or U29769 (N_29769,N_29399,N_29149);
and U29770 (N_29770,N_29142,N_28997);
xnor U29771 (N_29771,N_28940,N_28855);
or U29772 (N_29772,N_28992,N_29095);
nor U29773 (N_29773,N_28813,N_29025);
and U29774 (N_29774,N_28865,N_29234);
nor U29775 (N_29775,N_29159,N_28927);
and U29776 (N_29776,N_29162,N_29120);
and U29777 (N_29777,N_29337,N_29190);
nand U29778 (N_29778,N_29030,N_29364);
xnor U29779 (N_29779,N_29366,N_28937);
or U29780 (N_29780,N_29134,N_29038);
xnor U29781 (N_29781,N_28913,N_28808);
or U29782 (N_29782,N_29153,N_29116);
nand U29783 (N_29783,N_29174,N_28861);
nand U29784 (N_29784,N_28913,N_29147);
nor U29785 (N_29785,N_29377,N_29335);
nor U29786 (N_29786,N_28928,N_28982);
xnor U29787 (N_29787,N_28802,N_29203);
xnor U29788 (N_29788,N_29092,N_28808);
nand U29789 (N_29789,N_28927,N_29212);
xnor U29790 (N_29790,N_28953,N_29047);
xor U29791 (N_29791,N_29323,N_29212);
or U29792 (N_29792,N_28906,N_29303);
and U29793 (N_29793,N_28949,N_28962);
or U29794 (N_29794,N_28843,N_28884);
xor U29795 (N_29795,N_29078,N_29220);
xor U29796 (N_29796,N_29064,N_28989);
nand U29797 (N_29797,N_29390,N_28820);
nor U29798 (N_29798,N_29236,N_29186);
xor U29799 (N_29799,N_29316,N_28892);
xor U29800 (N_29800,N_29093,N_29360);
xor U29801 (N_29801,N_29251,N_28888);
nor U29802 (N_29802,N_29362,N_28908);
or U29803 (N_29803,N_28833,N_29249);
or U29804 (N_29804,N_28863,N_28804);
nand U29805 (N_29805,N_29262,N_29307);
nor U29806 (N_29806,N_28904,N_29067);
and U29807 (N_29807,N_29145,N_28932);
and U29808 (N_29808,N_28839,N_29069);
and U29809 (N_29809,N_28803,N_29356);
nor U29810 (N_29810,N_28967,N_29389);
nand U29811 (N_29811,N_29082,N_29072);
or U29812 (N_29812,N_28996,N_28944);
or U29813 (N_29813,N_29234,N_28873);
or U29814 (N_29814,N_29285,N_29358);
or U29815 (N_29815,N_28916,N_29387);
nor U29816 (N_29816,N_29062,N_29110);
nor U29817 (N_29817,N_29312,N_28941);
and U29818 (N_29818,N_29107,N_29190);
and U29819 (N_29819,N_28824,N_28804);
xnor U29820 (N_29820,N_28835,N_29357);
or U29821 (N_29821,N_29069,N_29238);
and U29822 (N_29822,N_28950,N_29117);
nor U29823 (N_29823,N_29107,N_28999);
nand U29824 (N_29824,N_29024,N_29107);
and U29825 (N_29825,N_29294,N_29295);
xnor U29826 (N_29826,N_29247,N_29020);
nor U29827 (N_29827,N_28836,N_29376);
xor U29828 (N_29828,N_28959,N_29059);
xnor U29829 (N_29829,N_28808,N_29048);
nor U29830 (N_29830,N_28847,N_29379);
nand U29831 (N_29831,N_29309,N_28842);
nand U29832 (N_29832,N_29187,N_29125);
nor U29833 (N_29833,N_29337,N_29109);
nor U29834 (N_29834,N_29162,N_29032);
nor U29835 (N_29835,N_29375,N_28809);
or U29836 (N_29836,N_29316,N_28982);
nand U29837 (N_29837,N_28918,N_28802);
nor U29838 (N_29838,N_29265,N_28848);
nand U29839 (N_29839,N_29385,N_28883);
xnor U29840 (N_29840,N_29133,N_29156);
xor U29841 (N_29841,N_28915,N_28939);
nor U29842 (N_29842,N_29279,N_29270);
and U29843 (N_29843,N_29311,N_29392);
nor U29844 (N_29844,N_29061,N_29396);
or U29845 (N_29845,N_29353,N_29082);
nor U29846 (N_29846,N_28821,N_29188);
and U29847 (N_29847,N_28943,N_29056);
nor U29848 (N_29848,N_29080,N_29032);
and U29849 (N_29849,N_29255,N_29115);
xor U29850 (N_29850,N_29038,N_29298);
nor U29851 (N_29851,N_29113,N_28890);
and U29852 (N_29852,N_28942,N_29062);
xnor U29853 (N_29853,N_29064,N_28868);
nor U29854 (N_29854,N_29326,N_28884);
nor U29855 (N_29855,N_28958,N_29023);
or U29856 (N_29856,N_28820,N_29100);
or U29857 (N_29857,N_29127,N_29035);
xnor U29858 (N_29858,N_29100,N_29278);
and U29859 (N_29859,N_28904,N_29084);
nor U29860 (N_29860,N_28886,N_28873);
or U29861 (N_29861,N_29348,N_28919);
or U29862 (N_29862,N_28913,N_28846);
nor U29863 (N_29863,N_29201,N_29355);
nor U29864 (N_29864,N_29210,N_29103);
xnor U29865 (N_29865,N_29000,N_29122);
nor U29866 (N_29866,N_28858,N_29348);
nand U29867 (N_29867,N_29196,N_29291);
and U29868 (N_29868,N_28999,N_28911);
or U29869 (N_29869,N_29134,N_29181);
xor U29870 (N_29870,N_29299,N_29300);
or U29871 (N_29871,N_29287,N_29224);
xor U29872 (N_29872,N_28828,N_29224);
or U29873 (N_29873,N_28897,N_29074);
and U29874 (N_29874,N_29010,N_29309);
nand U29875 (N_29875,N_28920,N_29248);
or U29876 (N_29876,N_29367,N_29365);
nor U29877 (N_29877,N_29338,N_28889);
nand U29878 (N_29878,N_29216,N_29043);
or U29879 (N_29879,N_29086,N_29264);
or U29880 (N_29880,N_29048,N_29167);
nand U29881 (N_29881,N_28968,N_29202);
and U29882 (N_29882,N_29046,N_29006);
or U29883 (N_29883,N_28947,N_28852);
and U29884 (N_29884,N_29310,N_28878);
or U29885 (N_29885,N_29153,N_29393);
nand U29886 (N_29886,N_29059,N_28898);
nand U29887 (N_29887,N_29271,N_29326);
nor U29888 (N_29888,N_29068,N_29308);
nand U29889 (N_29889,N_29120,N_29230);
xor U29890 (N_29890,N_29355,N_29270);
xor U29891 (N_29891,N_29385,N_28805);
and U29892 (N_29892,N_28942,N_29187);
xnor U29893 (N_29893,N_28928,N_29125);
or U29894 (N_29894,N_28966,N_28816);
nor U29895 (N_29895,N_28995,N_29050);
nor U29896 (N_29896,N_29162,N_28898);
nand U29897 (N_29897,N_29256,N_28959);
xnor U29898 (N_29898,N_29124,N_29178);
nor U29899 (N_29899,N_29371,N_28866);
or U29900 (N_29900,N_29052,N_28992);
xor U29901 (N_29901,N_29207,N_28892);
nand U29902 (N_29902,N_29140,N_29037);
nand U29903 (N_29903,N_29174,N_29263);
nand U29904 (N_29904,N_28992,N_28880);
or U29905 (N_29905,N_29265,N_29170);
nor U29906 (N_29906,N_28833,N_29015);
and U29907 (N_29907,N_28927,N_28812);
and U29908 (N_29908,N_29332,N_29132);
nand U29909 (N_29909,N_29171,N_29083);
and U29910 (N_29910,N_29130,N_29371);
or U29911 (N_29911,N_29250,N_28890);
xor U29912 (N_29912,N_28976,N_29114);
nor U29913 (N_29913,N_29092,N_29200);
nor U29914 (N_29914,N_28945,N_29042);
nor U29915 (N_29915,N_28916,N_28838);
nand U29916 (N_29916,N_29373,N_29267);
and U29917 (N_29917,N_29038,N_29002);
xor U29918 (N_29918,N_28986,N_29289);
nand U29919 (N_29919,N_29160,N_29077);
nor U29920 (N_29920,N_28912,N_28892);
and U29921 (N_29921,N_28951,N_29022);
or U29922 (N_29922,N_29136,N_28812);
and U29923 (N_29923,N_29198,N_29263);
xor U29924 (N_29924,N_29061,N_29290);
xnor U29925 (N_29925,N_28966,N_28912);
or U29926 (N_29926,N_29095,N_28867);
nor U29927 (N_29927,N_29286,N_29078);
or U29928 (N_29928,N_29393,N_29129);
xor U29929 (N_29929,N_28978,N_29275);
nand U29930 (N_29930,N_29289,N_29219);
nand U29931 (N_29931,N_29279,N_29347);
xnor U29932 (N_29932,N_29232,N_29317);
or U29933 (N_29933,N_28986,N_29395);
nand U29934 (N_29934,N_29120,N_29004);
nor U29935 (N_29935,N_29323,N_28911);
nor U29936 (N_29936,N_29025,N_28958);
nand U29937 (N_29937,N_28939,N_29175);
or U29938 (N_29938,N_28839,N_29313);
nand U29939 (N_29939,N_29162,N_29303);
or U29940 (N_29940,N_29073,N_28917);
and U29941 (N_29941,N_28900,N_28987);
nand U29942 (N_29942,N_29307,N_28922);
or U29943 (N_29943,N_28937,N_28815);
or U29944 (N_29944,N_29133,N_29319);
and U29945 (N_29945,N_28960,N_29204);
nand U29946 (N_29946,N_28969,N_29029);
or U29947 (N_29947,N_29324,N_28949);
nor U29948 (N_29948,N_29048,N_28972);
xnor U29949 (N_29949,N_28936,N_28802);
nand U29950 (N_29950,N_28828,N_28997);
or U29951 (N_29951,N_29248,N_29227);
nor U29952 (N_29952,N_29051,N_29235);
xnor U29953 (N_29953,N_28976,N_28935);
nand U29954 (N_29954,N_28852,N_29066);
nor U29955 (N_29955,N_28943,N_29233);
or U29956 (N_29956,N_28904,N_29340);
or U29957 (N_29957,N_29355,N_29017);
or U29958 (N_29958,N_29185,N_29383);
and U29959 (N_29959,N_28804,N_28867);
nor U29960 (N_29960,N_28852,N_29144);
nor U29961 (N_29961,N_29333,N_29239);
nand U29962 (N_29962,N_28850,N_29249);
xor U29963 (N_29963,N_29171,N_29152);
nor U29964 (N_29964,N_29067,N_28925);
nor U29965 (N_29965,N_28972,N_29287);
nand U29966 (N_29966,N_28892,N_29110);
or U29967 (N_29967,N_29307,N_29018);
nor U29968 (N_29968,N_29230,N_28944);
nor U29969 (N_29969,N_29190,N_28948);
nand U29970 (N_29970,N_29264,N_29280);
nand U29971 (N_29971,N_28941,N_28962);
xnor U29972 (N_29972,N_28897,N_28910);
xnor U29973 (N_29973,N_29040,N_29094);
nand U29974 (N_29974,N_29044,N_28918);
nor U29975 (N_29975,N_28862,N_28920);
and U29976 (N_29976,N_29393,N_29381);
and U29977 (N_29977,N_28944,N_29203);
and U29978 (N_29978,N_29340,N_28808);
nand U29979 (N_29979,N_28842,N_29332);
xnor U29980 (N_29980,N_29119,N_29101);
nand U29981 (N_29981,N_28838,N_29141);
or U29982 (N_29982,N_28963,N_29375);
nand U29983 (N_29983,N_28967,N_29153);
nor U29984 (N_29984,N_29326,N_29348);
xnor U29985 (N_29985,N_29108,N_29186);
nand U29986 (N_29986,N_29334,N_29020);
and U29987 (N_29987,N_28984,N_29342);
or U29988 (N_29988,N_28841,N_29351);
nand U29989 (N_29989,N_28853,N_29039);
and U29990 (N_29990,N_29087,N_29206);
or U29991 (N_29991,N_29114,N_29234);
nand U29992 (N_29992,N_29332,N_29212);
xor U29993 (N_29993,N_29319,N_29029);
xor U29994 (N_29994,N_29320,N_29362);
and U29995 (N_29995,N_28856,N_29249);
nand U29996 (N_29996,N_29331,N_29226);
and U29997 (N_29997,N_28934,N_28808);
and U29998 (N_29998,N_28859,N_29152);
nand U29999 (N_29999,N_29376,N_29083);
or UO_0 (O_0,N_29958,N_29490);
nand UO_1 (O_1,N_29623,N_29946);
or UO_2 (O_2,N_29472,N_29901);
nor UO_3 (O_3,N_29847,N_29488);
nor UO_4 (O_4,N_29471,N_29984);
xor UO_5 (O_5,N_29758,N_29821);
nand UO_6 (O_6,N_29628,N_29625);
or UO_7 (O_7,N_29678,N_29646);
nor UO_8 (O_8,N_29943,N_29727);
nor UO_9 (O_9,N_29790,N_29426);
and UO_10 (O_10,N_29427,N_29450);
or UO_11 (O_11,N_29576,N_29467);
and UO_12 (O_12,N_29504,N_29796);
nand UO_13 (O_13,N_29859,N_29831);
or UO_14 (O_14,N_29483,N_29671);
or UO_15 (O_15,N_29825,N_29752);
nor UO_16 (O_16,N_29714,N_29698);
nand UO_17 (O_17,N_29619,N_29844);
and UO_18 (O_18,N_29889,N_29761);
nor UO_19 (O_19,N_29502,N_29663);
and UO_20 (O_20,N_29439,N_29429);
or UO_21 (O_21,N_29972,N_29498);
xnor UO_22 (O_22,N_29939,N_29590);
nand UO_23 (O_23,N_29506,N_29963);
and UO_24 (O_24,N_29622,N_29533);
xor UO_25 (O_25,N_29729,N_29688);
and UO_26 (O_26,N_29775,N_29608);
nor UO_27 (O_27,N_29469,N_29417);
nand UO_28 (O_28,N_29929,N_29945);
nand UO_29 (O_29,N_29851,N_29914);
nand UO_30 (O_30,N_29485,N_29896);
xnor UO_31 (O_31,N_29604,N_29507);
or UO_32 (O_32,N_29433,N_29876);
and UO_33 (O_33,N_29853,N_29409);
and UO_34 (O_34,N_29791,N_29589);
and UO_35 (O_35,N_29640,N_29411);
and UO_36 (O_36,N_29509,N_29815);
nand UO_37 (O_37,N_29525,N_29437);
nor UO_38 (O_38,N_29406,N_29596);
or UO_39 (O_39,N_29459,N_29559);
nand UO_40 (O_40,N_29672,N_29536);
nor UO_41 (O_41,N_29846,N_29560);
xnor UO_42 (O_42,N_29400,N_29677);
xor UO_43 (O_43,N_29618,N_29805);
nand UO_44 (O_44,N_29695,N_29738);
nand UO_45 (O_45,N_29807,N_29880);
nor UO_46 (O_46,N_29781,N_29595);
nand UO_47 (O_47,N_29440,N_29991);
nor UO_48 (O_48,N_29569,N_29523);
xor UO_49 (O_49,N_29919,N_29690);
nor UO_50 (O_50,N_29572,N_29473);
nand UO_51 (O_51,N_29541,N_29574);
nand UO_52 (O_52,N_29718,N_29863);
xor UO_53 (O_53,N_29710,N_29636);
nor UO_54 (O_54,N_29545,N_29952);
or UO_55 (O_55,N_29705,N_29477);
nand UO_56 (O_56,N_29865,N_29835);
xor UO_57 (O_57,N_29850,N_29647);
nor UO_58 (O_58,N_29616,N_29500);
xor UO_59 (O_59,N_29910,N_29558);
and UO_60 (O_60,N_29403,N_29424);
nand UO_61 (O_61,N_29848,N_29818);
and UO_62 (O_62,N_29667,N_29823);
nand UO_63 (O_63,N_29555,N_29948);
or UO_64 (O_64,N_29787,N_29598);
nor UO_65 (O_65,N_29410,N_29974);
nand UO_66 (O_66,N_29931,N_29904);
and UO_67 (O_67,N_29754,N_29734);
and UO_68 (O_68,N_29928,N_29923);
nor UO_69 (O_69,N_29529,N_29903);
xnor UO_70 (O_70,N_29909,N_29587);
and UO_71 (O_71,N_29438,N_29662);
nand UO_72 (O_72,N_29926,N_29675);
nor UO_73 (O_73,N_29693,N_29493);
nor UO_74 (O_74,N_29836,N_29534);
or UO_75 (O_75,N_29922,N_29891);
xnor UO_76 (O_76,N_29425,N_29918);
xor UO_77 (O_77,N_29711,N_29402);
xor UO_78 (O_78,N_29512,N_29819);
xor UO_79 (O_79,N_29547,N_29911);
nor UO_80 (O_80,N_29606,N_29822);
nand UO_81 (O_81,N_29994,N_29656);
or UO_82 (O_82,N_29852,N_29981);
or UO_83 (O_83,N_29947,N_29924);
xnor UO_84 (O_84,N_29601,N_29940);
or UO_85 (O_85,N_29542,N_29820);
xor UO_86 (O_86,N_29716,N_29615);
or UO_87 (O_87,N_29782,N_29873);
and UO_88 (O_88,N_29921,N_29415);
nor UO_89 (O_89,N_29780,N_29768);
nand UO_90 (O_90,N_29935,N_29933);
and UO_91 (O_91,N_29436,N_29767);
xor UO_92 (O_92,N_29737,N_29510);
and UO_93 (O_93,N_29453,N_29670);
xnor UO_94 (O_94,N_29461,N_29961);
nand UO_95 (O_95,N_29686,N_29992);
and UO_96 (O_96,N_29451,N_29573);
nor UO_97 (O_97,N_29407,N_29661);
or UO_98 (O_98,N_29624,N_29505);
or UO_99 (O_99,N_29762,N_29474);
or UO_100 (O_100,N_29913,N_29816);
or UO_101 (O_101,N_29567,N_29480);
and UO_102 (O_102,N_29912,N_29503);
nand UO_103 (O_103,N_29418,N_29811);
and UO_104 (O_104,N_29476,N_29953);
xor UO_105 (O_105,N_29941,N_29980);
nand UO_106 (O_106,N_29641,N_29588);
or UO_107 (O_107,N_29867,N_29742);
xnor UO_108 (O_108,N_29976,N_29849);
nor UO_109 (O_109,N_29659,N_29932);
and UO_110 (O_110,N_29594,N_29468);
and UO_111 (O_111,N_29783,N_29518);
nand UO_112 (O_112,N_29916,N_29637);
nor UO_113 (O_113,N_29568,N_29521);
or UO_114 (O_114,N_29703,N_29513);
xor UO_115 (O_115,N_29784,N_29522);
xnor UO_116 (O_116,N_29905,N_29757);
xnor UO_117 (O_117,N_29704,N_29538);
nand UO_118 (O_118,N_29777,N_29475);
xor UO_119 (O_119,N_29826,N_29664);
or UO_120 (O_120,N_29920,N_29829);
and UO_121 (O_121,N_29855,N_29549);
xnor UO_122 (O_122,N_29645,N_29535);
and UO_123 (O_123,N_29810,N_29803);
nor UO_124 (O_124,N_29491,N_29895);
or UO_125 (O_125,N_29756,N_29466);
nor UO_126 (O_126,N_29561,N_29650);
and UO_127 (O_127,N_29967,N_29813);
nor UO_128 (O_128,N_29499,N_29550);
nand UO_129 (O_129,N_29746,N_29795);
nand UO_130 (O_130,N_29950,N_29445);
nor UO_131 (O_131,N_29422,N_29730);
or UO_132 (O_132,N_29676,N_29987);
or UO_133 (O_133,N_29764,N_29685);
and UO_134 (O_134,N_29915,N_29539);
and UO_135 (O_135,N_29553,N_29401);
nor UO_136 (O_136,N_29717,N_29888);
xor UO_137 (O_137,N_29842,N_29448);
nand UO_138 (O_138,N_29484,N_29900);
and UO_139 (O_139,N_29626,N_29857);
nand UO_140 (O_140,N_29890,N_29883);
or UO_141 (O_141,N_29733,N_29592);
nand UO_142 (O_142,N_29827,N_29460);
nor UO_143 (O_143,N_29556,N_29897);
xor UO_144 (O_144,N_29457,N_29800);
nand UO_145 (O_145,N_29627,N_29740);
and UO_146 (O_146,N_29769,N_29612);
or UO_147 (O_147,N_29744,N_29997);
xor UO_148 (O_148,N_29828,N_29726);
xor UO_149 (O_149,N_29583,N_29494);
nor UO_150 (O_150,N_29806,N_29731);
nand UO_151 (O_151,N_29610,N_29772);
and UO_152 (O_152,N_29899,N_29870);
nor UO_153 (O_153,N_29497,N_29902);
nand UO_154 (O_154,N_29998,N_29893);
nor UO_155 (O_155,N_29487,N_29691);
nor UO_156 (O_156,N_29833,N_29966);
xor UO_157 (O_157,N_29660,N_29809);
or UO_158 (O_158,N_29814,N_29470);
nand UO_159 (O_159,N_29942,N_29706);
nor UO_160 (O_160,N_29657,N_29778);
and UO_161 (O_161,N_29620,N_29860);
nor UO_162 (O_162,N_29715,N_29580);
and UO_163 (O_163,N_29571,N_29644);
and UO_164 (O_164,N_29884,N_29428);
and UO_165 (O_165,N_29789,N_29968);
and UO_166 (O_166,N_29786,N_29412);
xor UO_167 (O_167,N_29898,N_29674);
nor UO_168 (O_168,N_29621,N_29540);
and UO_169 (O_169,N_29957,N_29985);
or UO_170 (O_170,N_29944,N_29562);
or UO_171 (O_171,N_29511,N_29954);
nor UO_172 (O_172,N_29455,N_29712);
nand UO_173 (O_173,N_29748,N_29579);
and UO_174 (O_174,N_29404,N_29515);
xor UO_175 (O_175,N_29593,N_29838);
and UO_176 (O_176,N_29463,N_29456);
or UO_177 (O_177,N_29501,N_29747);
and UO_178 (O_178,N_29959,N_29633);
or UO_179 (O_179,N_29602,N_29689);
nand UO_180 (O_180,N_29435,N_29543);
and UO_181 (O_181,N_29441,N_29804);
nor UO_182 (O_182,N_29832,N_29669);
xnor UO_183 (O_183,N_29753,N_29544);
nand UO_184 (O_184,N_29874,N_29745);
xnor UO_185 (O_185,N_29817,N_29514);
and UO_186 (O_186,N_29696,N_29699);
or UO_187 (O_187,N_29938,N_29983);
nand UO_188 (O_188,N_29708,N_29955);
nor UO_189 (O_189,N_29443,N_29681);
and UO_190 (O_190,N_29887,N_29585);
xor UO_191 (O_191,N_29546,N_29578);
xnor UO_192 (O_192,N_29839,N_29599);
nand UO_193 (O_193,N_29799,N_29908);
or UO_194 (O_194,N_29530,N_29630);
nand UO_195 (O_195,N_29871,N_29692);
nor UO_196 (O_196,N_29845,N_29707);
or UO_197 (O_197,N_29993,N_29978);
nor UO_198 (O_198,N_29629,N_29728);
nand UO_199 (O_199,N_29824,N_29917);
and UO_200 (O_200,N_29990,N_29527);
and UO_201 (O_201,N_29834,N_29591);
xor UO_202 (O_202,N_29563,N_29416);
xnor UO_203 (O_203,N_29631,N_29970);
nor UO_204 (O_204,N_29749,N_29886);
and UO_205 (O_205,N_29632,N_29841);
nor UO_206 (O_206,N_29962,N_29794);
nor UO_207 (O_207,N_29864,N_29482);
nor UO_208 (O_208,N_29875,N_29581);
nor UO_209 (O_209,N_29779,N_29802);
and UO_210 (O_210,N_29486,N_29830);
or UO_211 (O_211,N_29434,N_29638);
or UO_212 (O_212,N_29964,N_29793);
nand UO_213 (O_213,N_29774,N_29597);
and UO_214 (O_214,N_29892,N_29723);
or UO_215 (O_215,N_29881,N_29432);
nand UO_216 (O_216,N_29458,N_29537);
or UO_217 (O_217,N_29449,N_29766);
nand UO_218 (O_218,N_29413,N_29776);
nand UO_219 (O_219,N_29526,N_29687);
nand UO_220 (O_220,N_29584,N_29995);
nor UO_221 (O_221,N_29520,N_29700);
and UO_222 (O_222,N_29603,N_29858);
nand UO_223 (O_223,N_29684,N_29808);
or UO_224 (O_224,N_29570,N_29770);
xnor UO_225 (O_225,N_29524,N_29577);
nor UO_226 (O_226,N_29763,N_29532);
nand UO_227 (O_227,N_29605,N_29907);
and UO_228 (O_228,N_29788,N_29879);
and UO_229 (O_229,N_29798,N_29652);
nand UO_230 (O_230,N_29643,N_29447);
nand UO_231 (O_231,N_29421,N_29736);
and UO_232 (O_232,N_29702,N_29801);
nor UO_233 (O_233,N_29843,N_29517);
nor UO_234 (O_234,N_29725,N_29408);
and UO_235 (O_235,N_29936,N_29713);
or UO_236 (O_236,N_29885,N_29613);
or UO_237 (O_237,N_29495,N_29882);
and UO_238 (O_238,N_29750,N_29701);
and UO_239 (O_239,N_29668,N_29999);
or UO_240 (O_240,N_29655,N_29464);
and UO_241 (O_241,N_29557,N_29697);
nor UO_242 (O_242,N_29519,N_29755);
and UO_243 (O_243,N_29617,N_29759);
xnor UO_244 (O_244,N_29531,N_29986);
xor UO_245 (O_245,N_29446,N_29639);
nor UO_246 (O_246,N_29683,N_29722);
and UO_247 (O_247,N_29444,N_29977);
nand UO_248 (O_248,N_29420,N_29960);
or UO_249 (O_249,N_29837,N_29930);
nor UO_250 (O_250,N_29565,N_29956);
nor UO_251 (O_251,N_29430,N_29431);
nor UO_252 (O_252,N_29869,N_29721);
and UO_253 (O_253,N_29666,N_29996);
nand UO_254 (O_254,N_29894,N_29925);
xor UO_255 (O_255,N_29982,N_29548);
and UO_256 (O_256,N_29949,N_29680);
nor UO_257 (O_257,N_29682,N_29653);
and UO_258 (O_258,N_29508,N_29840);
nor UO_259 (O_259,N_29566,N_29479);
and UO_260 (O_260,N_29492,N_29600);
and UO_261 (O_261,N_29634,N_29872);
xnor UO_262 (O_262,N_29861,N_29452);
or UO_263 (O_263,N_29934,N_29489);
or UO_264 (O_264,N_29654,N_29658);
or UO_265 (O_265,N_29649,N_29732);
or UO_266 (O_266,N_29679,N_29454);
nor UO_267 (O_267,N_29862,N_29773);
nand UO_268 (O_268,N_29969,N_29554);
xor UO_269 (O_269,N_29694,N_29609);
nor UO_270 (O_270,N_29854,N_29989);
nor UO_271 (O_271,N_29648,N_29720);
nand UO_272 (O_272,N_29709,N_29719);
xor UO_273 (O_273,N_29866,N_29975);
and UO_274 (O_274,N_29812,N_29792);
xor UO_275 (O_275,N_29760,N_29868);
nor UO_276 (O_276,N_29582,N_29614);
xnor UO_277 (O_277,N_29478,N_29551);
nor UO_278 (O_278,N_29965,N_29724);
nor UO_279 (O_279,N_29575,N_29673);
xnor UO_280 (O_280,N_29951,N_29765);
nand UO_281 (O_281,N_29979,N_29419);
nor UO_282 (O_282,N_29405,N_29785);
or UO_283 (O_283,N_29552,N_29797);
and UO_284 (O_284,N_29743,N_29516);
nand UO_285 (O_285,N_29735,N_29906);
and UO_286 (O_286,N_29496,N_29635);
and UO_287 (O_287,N_29739,N_29937);
nand UO_288 (O_288,N_29481,N_29771);
and UO_289 (O_289,N_29651,N_29973);
nor UO_290 (O_290,N_29586,N_29462);
and UO_291 (O_291,N_29607,N_29878);
or UO_292 (O_292,N_29741,N_29465);
xnor UO_293 (O_293,N_29423,N_29988);
and UO_294 (O_294,N_29665,N_29927);
or UO_295 (O_295,N_29564,N_29442);
nor UO_296 (O_296,N_29528,N_29856);
nor UO_297 (O_297,N_29971,N_29642);
xor UO_298 (O_298,N_29611,N_29751);
xor UO_299 (O_299,N_29414,N_29877);
nor UO_300 (O_300,N_29514,N_29687);
and UO_301 (O_301,N_29712,N_29517);
and UO_302 (O_302,N_29908,N_29689);
xor UO_303 (O_303,N_29484,N_29759);
nor UO_304 (O_304,N_29836,N_29462);
and UO_305 (O_305,N_29984,N_29867);
and UO_306 (O_306,N_29662,N_29767);
or UO_307 (O_307,N_29678,N_29711);
nor UO_308 (O_308,N_29708,N_29822);
nand UO_309 (O_309,N_29839,N_29779);
xor UO_310 (O_310,N_29889,N_29592);
and UO_311 (O_311,N_29883,N_29743);
nand UO_312 (O_312,N_29630,N_29875);
nor UO_313 (O_313,N_29703,N_29697);
nand UO_314 (O_314,N_29563,N_29662);
and UO_315 (O_315,N_29473,N_29487);
or UO_316 (O_316,N_29524,N_29663);
nor UO_317 (O_317,N_29591,N_29813);
xnor UO_318 (O_318,N_29601,N_29595);
nor UO_319 (O_319,N_29991,N_29955);
xor UO_320 (O_320,N_29713,N_29702);
xnor UO_321 (O_321,N_29631,N_29434);
or UO_322 (O_322,N_29865,N_29740);
xor UO_323 (O_323,N_29550,N_29945);
nor UO_324 (O_324,N_29484,N_29575);
or UO_325 (O_325,N_29841,N_29655);
nand UO_326 (O_326,N_29973,N_29610);
nor UO_327 (O_327,N_29794,N_29486);
and UO_328 (O_328,N_29402,N_29430);
and UO_329 (O_329,N_29519,N_29809);
nor UO_330 (O_330,N_29528,N_29543);
nand UO_331 (O_331,N_29818,N_29493);
nor UO_332 (O_332,N_29538,N_29403);
and UO_333 (O_333,N_29876,N_29447);
nor UO_334 (O_334,N_29683,N_29950);
and UO_335 (O_335,N_29975,N_29729);
nand UO_336 (O_336,N_29497,N_29555);
or UO_337 (O_337,N_29556,N_29820);
or UO_338 (O_338,N_29943,N_29926);
nor UO_339 (O_339,N_29470,N_29403);
nand UO_340 (O_340,N_29656,N_29538);
nor UO_341 (O_341,N_29798,N_29861);
nor UO_342 (O_342,N_29848,N_29684);
and UO_343 (O_343,N_29861,N_29920);
nor UO_344 (O_344,N_29506,N_29689);
or UO_345 (O_345,N_29541,N_29806);
xor UO_346 (O_346,N_29418,N_29450);
and UO_347 (O_347,N_29574,N_29996);
nand UO_348 (O_348,N_29895,N_29896);
nor UO_349 (O_349,N_29477,N_29722);
xnor UO_350 (O_350,N_29678,N_29466);
nor UO_351 (O_351,N_29731,N_29594);
nand UO_352 (O_352,N_29538,N_29683);
or UO_353 (O_353,N_29973,N_29613);
nand UO_354 (O_354,N_29433,N_29935);
nor UO_355 (O_355,N_29446,N_29427);
nor UO_356 (O_356,N_29924,N_29623);
or UO_357 (O_357,N_29674,N_29402);
nor UO_358 (O_358,N_29856,N_29971);
xor UO_359 (O_359,N_29754,N_29652);
nor UO_360 (O_360,N_29534,N_29847);
xnor UO_361 (O_361,N_29869,N_29900);
and UO_362 (O_362,N_29894,N_29652);
nand UO_363 (O_363,N_29561,N_29677);
nand UO_364 (O_364,N_29769,N_29743);
and UO_365 (O_365,N_29453,N_29992);
nand UO_366 (O_366,N_29885,N_29494);
or UO_367 (O_367,N_29513,N_29521);
xnor UO_368 (O_368,N_29412,N_29860);
and UO_369 (O_369,N_29970,N_29778);
and UO_370 (O_370,N_29835,N_29724);
and UO_371 (O_371,N_29471,N_29856);
nor UO_372 (O_372,N_29858,N_29465);
or UO_373 (O_373,N_29869,N_29833);
xnor UO_374 (O_374,N_29484,N_29630);
nand UO_375 (O_375,N_29713,N_29590);
nor UO_376 (O_376,N_29909,N_29493);
xnor UO_377 (O_377,N_29991,N_29722);
and UO_378 (O_378,N_29713,N_29779);
and UO_379 (O_379,N_29691,N_29842);
xnor UO_380 (O_380,N_29600,N_29852);
and UO_381 (O_381,N_29734,N_29450);
nor UO_382 (O_382,N_29675,N_29972);
nand UO_383 (O_383,N_29462,N_29651);
or UO_384 (O_384,N_29651,N_29768);
nor UO_385 (O_385,N_29574,N_29817);
nor UO_386 (O_386,N_29523,N_29793);
nor UO_387 (O_387,N_29578,N_29953);
and UO_388 (O_388,N_29530,N_29779);
nor UO_389 (O_389,N_29516,N_29889);
nor UO_390 (O_390,N_29794,N_29496);
nand UO_391 (O_391,N_29849,N_29758);
nand UO_392 (O_392,N_29967,N_29935);
or UO_393 (O_393,N_29489,N_29884);
xnor UO_394 (O_394,N_29638,N_29658);
or UO_395 (O_395,N_29772,N_29621);
and UO_396 (O_396,N_29931,N_29935);
nand UO_397 (O_397,N_29773,N_29499);
xor UO_398 (O_398,N_29569,N_29969);
nand UO_399 (O_399,N_29500,N_29605);
nor UO_400 (O_400,N_29617,N_29897);
nand UO_401 (O_401,N_29594,N_29733);
or UO_402 (O_402,N_29400,N_29482);
nand UO_403 (O_403,N_29680,N_29770);
nor UO_404 (O_404,N_29742,N_29767);
and UO_405 (O_405,N_29793,N_29503);
nand UO_406 (O_406,N_29934,N_29476);
xnor UO_407 (O_407,N_29829,N_29728);
xor UO_408 (O_408,N_29631,N_29643);
xnor UO_409 (O_409,N_29591,N_29792);
or UO_410 (O_410,N_29986,N_29844);
and UO_411 (O_411,N_29782,N_29408);
nand UO_412 (O_412,N_29518,N_29889);
or UO_413 (O_413,N_29911,N_29805);
and UO_414 (O_414,N_29943,N_29854);
or UO_415 (O_415,N_29477,N_29803);
nand UO_416 (O_416,N_29760,N_29507);
nor UO_417 (O_417,N_29730,N_29971);
nand UO_418 (O_418,N_29785,N_29808);
nand UO_419 (O_419,N_29862,N_29752);
and UO_420 (O_420,N_29898,N_29734);
nor UO_421 (O_421,N_29435,N_29600);
and UO_422 (O_422,N_29999,N_29421);
nand UO_423 (O_423,N_29802,N_29566);
xor UO_424 (O_424,N_29446,N_29839);
or UO_425 (O_425,N_29748,N_29536);
nand UO_426 (O_426,N_29709,N_29772);
xor UO_427 (O_427,N_29733,N_29893);
or UO_428 (O_428,N_29443,N_29724);
and UO_429 (O_429,N_29998,N_29835);
nand UO_430 (O_430,N_29896,N_29831);
or UO_431 (O_431,N_29534,N_29835);
xnor UO_432 (O_432,N_29502,N_29788);
xnor UO_433 (O_433,N_29619,N_29635);
nor UO_434 (O_434,N_29874,N_29707);
or UO_435 (O_435,N_29876,N_29859);
or UO_436 (O_436,N_29890,N_29775);
xnor UO_437 (O_437,N_29565,N_29530);
nor UO_438 (O_438,N_29845,N_29644);
and UO_439 (O_439,N_29913,N_29488);
and UO_440 (O_440,N_29622,N_29892);
nor UO_441 (O_441,N_29809,N_29700);
xnor UO_442 (O_442,N_29706,N_29810);
and UO_443 (O_443,N_29447,N_29880);
and UO_444 (O_444,N_29823,N_29514);
nand UO_445 (O_445,N_29620,N_29883);
nor UO_446 (O_446,N_29678,N_29800);
nor UO_447 (O_447,N_29665,N_29411);
nand UO_448 (O_448,N_29468,N_29680);
nand UO_449 (O_449,N_29616,N_29972);
and UO_450 (O_450,N_29436,N_29525);
or UO_451 (O_451,N_29639,N_29664);
nor UO_452 (O_452,N_29681,N_29986);
xor UO_453 (O_453,N_29465,N_29582);
or UO_454 (O_454,N_29599,N_29464);
or UO_455 (O_455,N_29862,N_29539);
nand UO_456 (O_456,N_29892,N_29636);
nand UO_457 (O_457,N_29960,N_29730);
xnor UO_458 (O_458,N_29845,N_29688);
nor UO_459 (O_459,N_29804,N_29634);
and UO_460 (O_460,N_29684,N_29687);
or UO_461 (O_461,N_29863,N_29623);
and UO_462 (O_462,N_29439,N_29984);
xor UO_463 (O_463,N_29704,N_29656);
and UO_464 (O_464,N_29896,N_29845);
nor UO_465 (O_465,N_29950,N_29750);
and UO_466 (O_466,N_29714,N_29806);
nor UO_467 (O_467,N_29413,N_29755);
or UO_468 (O_468,N_29787,N_29607);
and UO_469 (O_469,N_29513,N_29510);
nor UO_470 (O_470,N_29618,N_29581);
or UO_471 (O_471,N_29827,N_29996);
xor UO_472 (O_472,N_29700,N_29451);
xnor UO_473 (O_473,N_29597,N_29571);
nor UO_474 (O_474,N_29978,N_29531);
or UO_475 (O_475,N_29893,N_29517);
nand UO_476 (O_476,N_29654,N_29434);
and UO_477 (O_477,N_29681,N_29729);
nor UO_478 (O_478,N_29566,N_29966);
nand UO_479 (O_479,N_29628,N_29626);
xor UO_480 (O_480,N_29974,N_29960);
xnor UO_481 (O_481,N_29827,N_29633);
nand UO_482 (O_482,N_29743,N_29990);
nand UO_483 (O_483,N_29621,N_29925);
xnor UO_484 (O_484,N_29433,N_29405);
nand UO_485 (O_485,N_29504,N_29986);
nor UO_486 (O_486,N_29997,N_29554);
nand UO_487 (O_487,N_29471,N_29864);
nand UO_488 (O_488,N_29465,N_29978);
nor UO_489 (O_489,N_29418,N_29810);
xnor UO_490 (O_490,N_29471,N_29427);
xnor UO_491 (O_491,N_29791,N_29980);
or UO_492 (O_492,N_29605,N_29963);
nand UO_493 (O_493,N_29929,N_29819);
nand UO_494 (O_494,N_29630,N_29478);
nor UO_495 (O_495,N_29791,N_29839);
or UO_496 (O_496,N_29918,N_29563);
nand UO_497 (O_497,N_29589,N_29527);
and UO_498 (O_498,N_29503,N_29473);
and UO_499 (O_499,N_29513,N_29595);
xor UO_500 (O_500,N_29995,N_29672);
and UO_501 (O_501,N_29732,N_29921);
nand UO_502 (O_502,N_29435,N_29855);
nor UO_503 (O_503,N_29941,N_29605);
nand UO_504 (O_504,N_29577,N_29909);
and UO_505 (O_505,N_29683,N_29859);
nand UO_506 (O_506,N_29511,N_29454);
nor UO_507 (O_507,N_29877,N_29971);
or UO_508 (O_508,N_29616,N_29628);
nand UO_509 (O_509,N_29779,N_29623);
nor UO_510 (O_510,N_29735,N_29637);
nor UO_511 (O_511,N_29999,N_29602);
xnor UO_512 (O_512,N_29493,N_29862);
nor UO_513 (O_513,N_29419,N_29566);
xor UO_514 (O_514,N_29584,N_29807);
nor UO_515 (O_515,N_29876,N_29689);
xnor UO_516 (O_516,N_29980,N_29400);
nor UO_517 (O_517,N_29964,N_29817);
xor UO_518 (O_518,N_29758,N_29464);
and UO_519 (O_519,N_29731,N_29852);
or UO_520 (O_520,N_29663,N_29612);
xor UO_521 (O_521,N_29447,N_29660);
or UO_522 (O_522,N_29464,N_29830);
xor UO_523 (O_523,N_29657,N_29429);
and UO_524 (O_524,N_29456,N_29765);
and UO_525 (O_525,N_29756,N_29508);
or UO_526 (O_526,N_29402,N_29565);
nand UO_527 (O_527,N_29529,N_29581);
nor UO_528 (O_528,N_29403,N_29845);
nand UO_529 (O_529,N_29458,N_29436);
and UO_530 (O_530,N_29839,N_29943);
and UO_531 (O_531,N_29702,N_29999);
or UO_532 (O_532,N_29547,N_29868);
or UO_533 (O_533,N_29678,N_29653);
or UO_534 (O_534,N_29488,N_29418);
nand UO_535 (O_535,N_29782,N_29991);
nand UO_536 (O_536,N_29761,N_29893);
and UO_537 (O_537,N_29789,N_29901);
and UO_538 (O_538,N_29684,N_29980);
xor UO_539 (O_539,N_29863,N_29692);
and UO_540 (O_540,N_29993,N_29647);
xnor UO_541 (O_541,N_29998,N_29786);
nor UO_542 (O_542,N_29821,N_29754);
xor UO_543 (O_543,N_29683,N_29962);
nand UO_544 (O_544,N_29842,N_29552);
xor UO_545 (O_545,N_29590,N_29715);
or UO_546 (O_546,N_29611,N_29438);
and UO_547 (O_547,N_29530,N_29963);
xor UO_548 (O_548,N_29713,N_29780);
nand UO_549 (O_549,N_29711,N_29889);
or UO_550 (O_550,N_29928,N_29620);
or UO_551 (O_551,N_29876,N_29507);
and UO_552 (O_552,N_29908,N_29510);
or UO_553 (O_553,N_29604,N_29769);
nor UO_554 (O_554,N_29569,N_29421);
and UO_555 (O_555,N_29596,N_29461);
xnor UO_556 (O_556,N_29468,N_29874);
or UO_557 (O_557,N_29900,N_29598);
xnor UO_558 (O_558,N_29784,N_29664);
and UO_559 (O_559,N_29584,N_29717);
nand UO_560 (O_560,N_29641,N_29906);
or UO_561 (O_561,N_29777,N_29785);
and UO_562 (O_562,N_29523,N_29588);
or UO_563 (O_563,N_29505,N_29871);
nor UO_564 (O_564,N_29748,N_29484);
or UO_565 (O_565,N_29550,N_29828);
nand UO_566 (O_566,N_29437,N_29554);
nand UO_567 (O_567,N_29797,N_29964);
nand UO_568 (O_568,N_29756,N_29467);
xor UO_569 (O_569,N_29879,N_29826);
nand UO_570 (O_570,N_29847,N_29427);
and UO_571 (O_571,N_29607,N_29868);
nand UO_572 (O_572,N_29674,N_29401);
nand UO_573 (O_573,N_29578,N_29533);
xor UO_574 (O_574,N_29615,N_29840);
xnor UO_575 (O_575,N_29503,N_29933);
nand UO_576 (O_576,N_29887,N_29966);
nor UO_577 (O_577,N_29921,N_29468);
or UO_578 (O_578,N_29908,N_29582);
xor UO_579 (O_579,N_29741,N_29457);
nor UO_580 (O_580,N_29428,N_29773);
nor UO_581 (O_581,N_29950,N_29967);
or UO_582 (O_582,N_29945,N_29749);
nand UO_583 (O_583,N_29705,N_29602);
nor UO_584 (O_584,N_29645,N_29572);
nand UO_585 (O_585,N_29604,N_29749);
or UO_586 (O_586,N_29489,N_29923);
or UO_587 (O_587,N_29717,N_29681);
xnor UO_588 (O_588,N_29782,N_29783);
and UO_589 (O_589,N_29490,N_29625);
nor UO_590 (O_590,N_29627,N_29828);
nor UO_591 (O_591,N_29634,N_29632);
or UO_592 (O_592,N_29492,N_29760);
xor UO_593 (O_593,N_29806,N_29688);
nand UO_594 (O_594,N_29901,N_29651);
and UO_595 (O_595,N_29953,N_29497);
nor UO_596 (O_596,N_29652,N_29732);
nand UO_597 (O_597,N_29626,N_29519);
xnor UO_598 (O_598,N_29923,N_29426);
and UO_599 (O_599,N_29842,N_29529);
and UO_600 (O_600,N_29841,N_29847);
and UO_601 (O_601,N_29657,N_29821);
or UO_602 (O_602,N_29524,N_29534);
or UO_603 (O_603,N_29673,N_29859);
or UO_604 (O_604,N_29824,N_29914);
xor UO_605 (O_605,N_29458,N_29631);
or UO_606 (O_606,N_29943,N_29799);
nor UO_607 (O_607,N_29743,N_29826);
xnor UO_608 (O_608,N_29886,N_29960);
or UO_609 (O_609,N_29434,N_29458);
nand UO_610 (O_610,N_29707,N_29609);
or UO_611 (O_611,N_29429,N_29421);
nand UO_612 (O_612,N_29987,N_29734);
and UO_613 (O_613,N_29643,N_29660);
xnor UO_614 (O_614,N_29899,N_29965);
nand UO_615 (O_615,N_29967,N_29560);
nand UO_616 (O_616,N_29521,N_29971);
or UO_617 (O_617,N_29404,N_29685);
nand UO_618 (O_618,N_29691,N_29575);
and UO_619 (O_619,N_29531,N_29669);
and UO_620 (O_620,N_29756,N_29986);
nor UO_621 (O_621,N_29629,N_29783);
xnor UO_622 (O_622,N_29719,N_29538);
or UO_623 (O_623,N_29930,N_29596);
xor UO_624 (O_624,N_29631,N_29692);
or UO_625 (O_625,N_29735,N_29494);
or UO_626 (O_626,N_29431,N_29808);
and UO_627 (O_627,N_29531,N_29479);
xor UO_628 (O_628,N_29588,N_29736);
xnor UO_629 (O_629,N_29620,N_29442);
or UO_630 (O_630,N_29907,N_29720);
and UO_631 (O_631,N_29643,N_29831);
or UO_632 (O_632,N_29772,N_29648);
and UO_633 (O_633,N_29641,N_29423);
and UO_634 (O_634,N_29415,N_29593);
nor UO_635 (O_635,N_29856,N_29723);
xor UO_636 (O_636,N_29855,N_29583);
or UO_637 (O_637,N_29678,N_29427);
nor UO_638 (O_638,N_29485,N_29465);
or UO_639 (O_639,N_29401,N_29637);
xor UO_640 (O_640,N_29637,N_29715);
or UO_641 (O_641,N_29656,N_29690);
xnor UO_642 (O_642,N_29587,N_29741);
and UO_643 (O_643,N_29775,N_29568);
xor UO_644 (O_644,N_29643,N_29477);
nor UO_645 (O_645,N_29668,N_29923);
nor UO_646 (O_646,N_29651,N_29816);
or UO_647 (O_647,N_29400,N_29846);
and UO_648 (O_648,N_29536,N_29477);
xnor UO_649 (O_649,N_29456,N_29871);
nor UO_650 (O_650,N_29769,N_29779);
xor UO_651 (O_651,N_29476,N_29987);
or UO_652 (O_652,N_29841,N_29548);
or UO_653 (O_653,N_29435,N_29954);
xor UO_654 (O_654,N_29849,N_29423);
or UO_655 (O_655,N_29944,N_29500);
nor UO_656 (O_656,N_29885,N_29918);
nand UO_657 (O_657,N_29809,N_29742);
nand UO_658 (O_658,N_29546,N_29860);
nor UO_659 (O_659,N_29525,N_29890);
nor UO_660 (O_660,N_29946,N_29768);
and UO_661 (O_661,N_29985,N_29415);
or UO_662 (O_662,N_29708,N_29939);
and UO_663 (O_663,N_29535,N_29547);
nand UO_664 (O_664,N_29657,N_29972);
nor UO_665 (O_665,N_29479,N_29930);
and UO_666 (O_666,N_29458,N_29912);
nand UO_667 (O_667,N_29754,N_29870);
and UO_668 (O_668,N_29854,N_29860);
nor UO_669 (O_669,N_29501,N_29615);
nand UO_670 (O_670,N_29735,N_29497);
nand UO_671 (O_671,N_29881,N_29658);
nand UO_672 (O_672,N_29798,N_29422);
or UO_673 (O_673,N_29644,N_29704);
xnor UO_674 (O_674,N_29434,N_29498);
nand UO_675 (O_675,N_29695,N_29847);
xor UO_676 (O_676,N_29877,N_29890);
nor UO_677 (O_677,N_29836,N_29746);
nand UO_678 (O_678,N_29831,N_29746);
nand UO_679 (O_679,N_29550,N_29870);
nand UO_680 (O_680,N_29952,N_29799);
nand UO_681 (O_681,N_29446,N_29674);
nor UO_682 (O_682,N_29879,N_29931);
xor UO_683 (O_683,N_29774,N_29770);
and UO_684 (O_684,N_29726,N_29697);
nand UO_685 (O_685,N_29522,N_29819);
and UO_686 (O_686,N_29767,N_29677);
nor UO_687 (O_687,N_29465,N_29468);
nand UO_688 (O_688,N_29429,N_29800);
and UO_689 (O_689,N_29528,N_29928);
nor UO_690 (O_690,N_29740,N_29903);
nor UO_691 (O_691,N_29489,N_29905);
or UO_692 (O_692,N_29416,N_29790);
or UO_693 (O_693,N_29454,N_29435);
nand UO_694 (O_694,N_29905,N_29415);
or UO_695 (O_695,N_29658,N_29582);
or UO_696 (O_696,N_29942,N_29841);
nand UO_697 (O_697,N_29821,N_29457);
nand UO_698 (O_698,N_29609,N_29585);
nor UO_699 (O_699,N_29726,N_29549);
and UO_700 (O_700,N_29773,N_29516);
and UO_701 (O_701,N_29808,N_29519);
nand UO_702 (O_702,N_29476,N_29741);
or UO_703 (O_703,N_29666,N_29465);
and UO_704 (O_704,N_29785,N_29730);
or UO_705 (O_705,N_29977,N_29490);
nand UO_706 (O_706,N_29574,N_29664);
nor UO_707 (O_707,N_29940,N_29490);
nand UO_708 (O_708,N_29872,N_29892);
or UO_709 (O_709,N_29740,N_29655);
nand UO_710 (O_710,N_29747,N_29500);
nor UO_711 (O_711,N_29930,N_29809);
nand UO_712 (O_712,N_29796,N_29477);
or UO_713 (O_713,N_29752,N_29596);
nand UO_714 (O_714,N_29670,N_29559);
xnor UO_715 (O_715,N_29602,N_29561);
xnor UO_716 (O_716,N_29422,N_29486);
or UO_717 (O_717,N_29465,N_29973);
xor UO_718 (O_718,N_29427,N_29906);
nand UO_719 (O_719,N_29612,N_29723);
nand UO_720 (O_720,N_29829,N_29944);
xnor UO_721 (O_721,N_29879,N_29591);
or UO_722 (O_722,N_29894,N_29656);
xnor UO_723 (O_723,N_29510,N_29925);
and UO_724 (O_724,N_29422,N_29801);
or UO_725 (O_725,N_29771,N_29723);
nand UO_726 (O_726,N_29742,N_29735);
nor UO_727 (O_727,N_29937,N_29752);
nor UO_728 (O_728,N_29626,N_29592);
xor UO_729 (O_729,N_29591,N_29730);
nor UO_730 (O_730,N_29405,N_29522);
nand UO_731 (O_731,N_29799,N_29467);
and UO_732 (O_732,N_29949,N_29643);
xnor UO_733 (O_733,N_29675,N_29934);
nor UO_734 (O_734,N_29775,N_29548);
or UO_735 (O_735,N_29909,N_29597);
nor UO_736 (O_736,N_29835,N_29642);
nand UO_737 (O_737,N_29627,N_29560);
nand UO_738 (O_738,N_29849,N_29938);
xnor UO_739 (O_739,N_29805,N_29871);
nand UO_740 (O_740,N_29733,N_29702);
nand UO_741 (O_741,N_29561,N_29604);
nand UO_742 (O_742,N_29870,N_29435);
xnor UO_743 (O_743,N_29425,N_29959);
nor UO_744 (O_744,N_29428,N_29402);
nor UO_745 (O_745,N_29896,N_29627);
nor UO_746 (O_746,N_29739,N_29548);
nand UO_747 (O_747,N_29886,N_29764);
nand UO_748 (O_748,N_29999,N_29699);
xor UO_749 (O_749,N_29701,N_29623);
nor UO_750 (O_750,N_29496,N_29459);
xor UO_751 (O_751,N_29517,N_29996);
nor UO_752 (O_752,N_29906,N_29896);
nand UO_753 (O_753,N_29529,N_29997);
and UO_754 (O_754,N_29820,N_29811);
and UO_755 (O_755,N_29884,N_29850);
nand UO_756 (O_756,N_29717,N_29444);
and UO_757 (O_757,N_29462,N_29403);
or UO_758 (O_758,N_29623,N_29411);
and UO_759 (O_759,N_29439,N_29951);
nor UO_760 (O_760,N_29619,N_29924);
nor UO_761 (O_761,N_29757,N_29804);
and UO_762 (O_762,N_29489,N_29532);
nor UO_763 (O_763,N_29882,N_29430);
nor UO_764 (O_764,N_29605,N_29530);
nor UO_765 (O_765,N_29778,N_29850);
or UO_766 (O_766,N_29495,N_29736);
nor UO_767 (O_767,N_29992,N_29662);
and UO_768 (O_768,N_29652,N_29762);
or UO_769 (O_769,N_29744,N_29629);
nor UO_770 (O_770,N_29905,N_29985);
and UO_771 (O_771,N_29762,N_29679);
nand UO_772 (O_772,N_29586,N_29830);
nand UO_773 (O_773,N_29872,N_29968);
xnor UO_774 (O_774,N_29979,N_29832);
nor UO_775 (O_775,N_29779,N_29605);
and UO_776 (O_776,N_29425,N_29465);
or UO_777 (O_777,N_29477,N_29864);
nor UO_778 (O_778,N_29735,N_29787);
xor UO_779 (O_779,N_29647,N_29483);
or UO_780 (O_780,N_29933,N_29755);
nor UO_781 (O_781,N_29774,N_29612);
and UO_782 (O_782,N_29738,N_29734);
or UO_783 (O_783,N_29800,N_29478);
or UO_784 (O_784,N_29633,N_29473);
nor UO_785 (O_785,N_29745,N_29717);
or UO_786 (O_786,N_29802,N_29481);
nand UO_787 (O_787,N_29906,N_29431);
nor UO_788 (O_788,N_29780,N_29767);
nand UO_789 (O_789,N_29820,N_29969);
xnor UO_790 (O_790,N_29555,N_29506);
xnor UO_791 (O_791,N_29541,N_29741);
nand UO_792 (O_792,N_29848,N_29643);
xnor UO_793 (O_793,N_29627,N_29423);
xor UO_794 (O_794,N_29663,N_29983);
and UO_795 (O_795,N_29659,N_29825);
and UO_796 (O_796,N_29418,N_29520);
and UO_797 (O_797,N_29530,N_29606);
nand UO_798 (O_798,N_29784,N_29465);
xnor UO_799 (O_799,N_29718,N_29990);
nand UO_800 (O_800,N_29402,N_29788);
nor UO_801 (O_801,N_29999,N_29796);
nand UO_802 (O_802,N_29676,N_29560);
or UO_803 (O_803,N_29867,N_29627);
nand UO_804 (O_804,N_29772,N_29923);
nand UO_805 (O_805,N_29624,N_29990);
nor UO_806 (O_806,N_29703,N_29633);
nand UO_807 (O_807,N_29802,N_29529);
and UO_808 (O_808,N_29542,N_29637);
xor UO_809 (O_809,N_29925,N_29440);
nor UO_810 (O_810,N_29815,N_29752);
xnor UO_811 (O_811,N_29515,N_29423);
nand UO_812 (O_812,N_29504,N_29916);
xor UO_813 (O_813,N_29468,N_29847);
xnor UO_814 (O_814,N_29914,N_29915);
and UO_815 (O_815,N_29501,N_29731);
xnor UO_816 (O_816,N_29919,N_29426);
nand UO_817 (O_817,N_29799,N_29887);
and UO_818 (O_818,N_29688,N_29978);
xnor UO_819 (O_819,N_29525,N_29840);
nor UO_820 (O_820,N_29596,N_29917);
nand UO_821 (O_821,N_29612,N_29857);
nor UO_822 (O_822,N_29560,N_29927);
and UO_823 (O_823,N_29437,N_29442);
nor UO_824 (O_824,N_29695,N_29408);
or UO_825 (O_825,N_29938,N_29783);
nor UO_826 (O_826,N_29631,N_29469);
and UO_827 (O_827,N_29437,N_29879);
or UO_828 (O_828,N_29781,N_29617);
and UO_829 (O_829,N_29814,N_29713);
nor UO_830 (O_830,N_29477,N_29403);
xnor UO_831 (O_831,N_29958,N_29649);
xnor UO_832 (O_832,N_29651,N_29585);
xnor UO_833 (O_833,N_29610,N_29676);
nand UO_834 (O_834,N_29420,N_29431);
or UO_835 (O_835,N_29522,N_29480);
nor UO_836 (O_836,N_29837,N_29917);
nand UO_837 (O_837,N_29651,N_29539);
and UO_838 (O_838,N_29864,N_29484);
or UO_839 (O_839,N_29806,N_29657);
or UO_840 (O_840,N_29659,N_29422);
and UO_841 (O_841,N_29778,N_29457);
or UO_842 (O_842,N_29856,N_29973);
nor UO_843 (O_843,N_29829,N_29939);
xor UO_844 (O_844,N_29680,N_29924);
nor UO_845 (O_845,N_29800,N_29413);
and UO_846 (O_846,N_29655,N_29476);
and UO_847 (O_847,N_29711,N_29549);
and UO_848 (O_848,N_29602,N_29620);
nand UO_849 (O_849,N_29705,N_29817);
xor UO_850 (O_850,N_29782,N_29976);
nand UO_851 (O_851,N_29451,N_29472);
nand UO_852 (O_852,N_29438,N_29772);
nand UO_853 (O_853,N_29624,N_29464);
xor UO_854 (O_854,N_29648,N_29668);
xnor UO_855 (O_855,N_29668,N_29781);
nand UO_856 (O_856,N_29926,N_29716);
nor UO_857 (O_857,N_29758,N_29711);
nor UO_858 (O_858,N_29702,N_29707);
or UO_859 (O_859,N_29757,N_29752);
xor UO_860 (O_860,N_29797,N_29425);
and UO_861 (O_861,N_29425,N_29931);
and UO_862 (O_862,N_29686,N_29468);
nand UO_863 (O_863,N_29762,N_29572);
and UO_864 (O_864,N_29798,N_29863);
or UO_865 (O_865,N_29471,N_29972);
or UO_866 (O_866,N_29517,N_29958);
and UO_867 (O_867,N_29508,N_29456);
xor UO_868 (O_868,N_29974,N_29878);
nand UO_869 (O_869,N_29816,N_29971);
nor UO_870 (O_870,N_29989,N_29741);
or UO_871 (O_871,N_29469,N_29618);
xor UO_872 (O_872,N_29860,N_29419);
nand UO_873 (O_873,N_29635,N_29582);
xor UO_874 (O_874,N_29881,N_29759);
or UO_875 (O_875,N_29849,N_29745);
xnor UO_876 (O_876,N_29790,N_29636);
or UO_877 (O_877,N_29502,N_29467);
nand UO_878 (O_878,N_29971,N_29735);
or UO_879 (O_879,N_29737,N_29511);
nand UO_880 (O_880,N_29605,N_29812);
nor UO_881 (O_881,N_29542,N_29826);
nand UO_882 (O_882,N_29528,N_29466);
or UO_883 (O_883,N_29706,N_29555);
and UO_884 (O_884,N_29576,N_29503);
nor UO_885 (O_885,N_29749,N_29401);
xor UO_886 (O_886,N_29820,N_29500);
nand UO_887 (O_887,N_29912,N_29828);
and UO_888 (O_888,N_29528,N_29653);
xor UO_889 (O_889,N_29755,N_29862);
nand UO_890 (O_890,N_29752,N_29883);
or UO_891 (O_891,N_29678,N_29700);
or UO_892 (O_892,N_29491,N_29780);
and UO_893 (O_893,N_29796,N_29659);
nand UO_894 (O_894,N_29746,N_29939);
and UO_895 (O_895,N_29901,N_29661);
nor UO_896 (O_896,N_29806,N_29984);
and UO_897 (O_897,N_29844,N_29407);
xor UO_898 (O_898,N_29546,N_29854);
nand UO_899 (O_899,N_29411,N_29491);
nor UO_900 (O_900,N_29794,N_29418);
and UO_901 (O_901,N_29635,N_29474);
nor UO_902 (O_902,N_29607,N_29465);
xor UO_903 (O_903,N_29639,N_29912);
xor UO_904 (O_904,N_29653,N_29667);
nand UO_905 (O_905,N_29777,N_29722);
or UO_906 (O_906,N_29902,N_29724);
or UO_907 (O_907,N_29514,N_29767);
nor UO_908 (O_908,N_29994,N_29472);
nand UO_909 (O_909,N_29645,N_29716);
nor UO_910 (O_910,N_29419,N_29913);
nand UO_911 (O_911,N_29709,N_29926);
and UO_912 (O_912,N_29754,N_29542);
xor UO_913 (O_913,N_29441,N_29861);
xor UO_914 (O_914,N_29856,N_29526);
xnor UO_915 (O_915,N_29432,N_29951);
nand UO_916 (O_916,N_29868,N_29588);
and UO_917 (O_917,N_29757,N_29984);
and UO_918 (O_918,N_29900,N_29496);
and UO_919 (O_919,N_29943,N_29796);
xnor UO_920 (O_920,N_29649,N_29954);
xnor UO_921 (O_921,N_29720,N_29858);
xnor UO_922 (O_922,N_29456,N_29672);
xor UO_923 (O_923,N_29808,N_29633);
and UO_924 (O_924,N_29838,N_29423);
or UO_925 (O_925,N_29839,N_29715);
nand UO_926 (O_926,N_29818,N_29830);
and UO_927 (O_927,N_29493,N_29922);
nor UO_928 (O_928,N_29408,N_29955);
nor UO_929 (O_929,N_29686,N_29590);
and UO_930 (O_930,N_29740,N_29415);
and UO_931 (O_931,N_29492,N_29628);
xor UO_932 (O_932,N_29413,N_29645);
nand UO_933 (O_933,N_29801,N_29760);
or UO_934 (O_934,N_29444,N_29447);
xnor UO_935 (O_935,N_29945,N_29817);
and UO_936 (O_936,N_29816,N_29627);
or UO_937 (O_937,N_29859,N_29559);
and UO_938 (O_938,N_29766,N_29819);
nand UO_939 (O_939,N_29499,N_29544);
xor UO_940 (O_940,N_29842,N_29650);
or UO_941 (O_941,N_29704,N_29766);
nor UO_942 (O_942,N_29608,N_29773);
nand UO_943 (O_943,N_29638,N_29655);
nand UO_944 (O_944,N_29577,N_29451);
nor UO_945 (O_945,N_29900,N_29712);
or UO_946 (O_946,N_29718,N_29801);
and UO_947 (O_947,N_29652,N_29769);
or UO_948 (O_948,N_29671,N_29447);
and UO_949 (O_949,N_29879,N_29822);
xor UO_950 (O_950,N_29481,N_29593);
and UO_951 (O_951,N_29520,N_29734);
xnor UO_952 (O_952,N_29550,N_29696);
and UO_953 (O_953,N_29938,N_29667);
nor UO_954 (O_954,N_29828,N_29596);
and UO_955 (O_955,N_29587,N_29602);
or UO_956 (O_956,N_29913,N_29641);
nand UO_957 (O_957,N_29805,N_29668);
nand UO_958 (O_958,N_29617,N_29554);
or UO_959 (O_959,N_29642,N_29768);
xor UO_960 (O_960,N_29575,N_29569);
and UO_961 (O_961,N_29871,N_29521);
xor UO_962 (O_962,N_29530,N_29783);
or UO_963 (O_963,N_29835,N_29554);
or UO_964 (O_964,N_29572,N_29537);
xnor UO_965 (O_965,N_29734,N_29969);
or UO_966 (O_966,N_29578,N_29419);
xor UO_967 (O_967,N_29578,N_29932);
xnor UO_968 (O_968,N_29964,N_29745);
xnor UO_969 (O_969,N_29490,N_29950);
nand UO_970 (O_970,N_29839,N_29738);
and UO_971 (O_971,N_29550,N_29519);
and UO_972 (O_972,N_29882,N_29785);
or UO_973 (O_973,N_29627,N_29599);
xnor UO_974 (O_974,N_29517,N_29498);
nor UO_975 (O_975,N_29788,N_29696);
nand UO_976 (O_976,N_29465,N_29686);
nand UO_977 (O_977,N_29648,N_29449);
nand UO_978 (O_978,N_29895,N_29739);
and UO_979 (O_979,N_29968,N_29769);
or UO_980 (O_980,N_29957,N_29611);
and UO_981 (O_981,N_29825,N_29459);
nand UO_982 (O_982,N_29534,N_29606);
nand UO_983 (O_983,N_29566,N_29801);
and UO_984 (O_984,N_29783,N_29983);
or UO_985 (O_985,N_29886,N_29859);
nand UO_986 (O_986,N_29487,N_29938);
or UO_987 (O_987,N_29999,N_29993);
xnor UO_988 (O_988,N_29458,N_29451);
nand UO_989 (O_989,N_29537,N_29532);
nand UO_990 (O_990,N_29601,N_29597);
nand UO_991 (O_991,N_29954,N_29840);
xnor UO_992 (O_992,N_29407,N_29927);
or UO_993 (O_993,N_29979,N_29777);
and UO_994 (O_994,N_29535,N_29758);
and UO_995 (O_995,N_29744,N_29811);
xor UO_996 (O_996,N_29518,N_29485);
nand UO_997 (O_997,N_29410,N_29734);
or UO_998 (O_998,N_29633,N_29439);
and UO_999 (O_999,N_29707,N_29941);
nand UO_1000 (O_1000,N_29760,N_29741);
xor UO_1001 (O_1001,N_29516,N_29627);
nand UO_1002 (O_1002,N_29639,N_29802);
xor UO_1003 (O_1003,N_29478,N_29405);
nor UO_1004 (O_1004,N_29837,N_29613);
xor UO_1005 (O_1005,N_29846,N_29798);
xor UO_1006 (O_1006,N_29952,N_29618);
nand UO_1007 (O_1007,N_29685,N_29585);
nor UO_1008 (O_1008,N_29407,N_29931);
and UO_1009 (O_1009,N_29408,N_29563);
xor UO_1010 (O_1010,N_29555,N_29730);
nor UO_1011 (O_1011,N_29565,N_29663);
nand UO_1012 (O_1012,N_29699,N_29790);
or UO_1013 (O_1013,N_29871,N_29895);
and UO_1014 (O_1014,N_29806,N_29963);
or UO_1015 (O_1015,N_29993,N_29909);
nand UO_1016 (O_1016,N_29704,N_29968);
nor UO_1017 (O_1017,N_29994,N_29974);
xnor UO_1018 (O_1018,N_29462,N_29833);
and UO_1019 (O_1019,N_29979,N_29439);
and UO_1020 (O_1020,N_29752,N_29429);
nand UO_1021 (O_1021,N_29441,N_29685);
nor UO_1022 (O_1022,N_29501,N_29868);
nor UO_1023 (O_1023,N_29777,N_29787);
and UO_1024 (O_1024,N_29730,N_29517);
xnor UO_1025 (O_1025,N_29776,N_29779);
nor UO_1026 (O_1026,N_29835,N_29759);
xnor UO_1027 (O_1027,N_29924,N_29963);
nand UO_1028 (O_1028,N_29544,N_29925);
nand UO_1029 (O_1029,N_29801,N_29896);
or UO_1030 (O_1030,N_29676,N_29623);
or UO_1031 (O_1031,N_29874,N_29783);
or UO_1032 (O_1032,N_29979,N_29942);
and UO_1033 (O_1033,N_29943,N_29784);
nor UO_1034 (O_1034,N_29463,N_29816);
xnor UO_1035 (O_1035,N_29408,N_29795);
xor UO_1036 (O_1036,N_29537,N_29879);
xor UO_1037 (O_1037,N_29962,N_29848);
and UO_1038 (O_1038,N_29485,N_29579);
xnor UO_1039 (O_1039,N_29885,N_29961);
nand UO_1040 (O_1040,N_29900,N_29695);
or UO_1041 (O_1041,N_29988,N_29753);
or UO_1042 (O_1042,N_29747,N_29514);
nor UO_1043 (O_1043,N_29576,N_29818);
nor UO_1044 (O_1044,N_29426,N_29639);
or UO_1045 (O_1045,N_29401,N_29722);
nor UO_1046 (O_1046,N_29452,N_29664);
or UO_1047 (O_1047,N_29445,N_29905);
or UO_1048 (O_1048,N_29876,N_29998);
xor UO_1049 (O_1049,N_29529,N_29701);
xor UO_1050 (O_1050,N_29547,N_29610);
and UO_1051 (O_1051,N_29821,N_29686);
xnor UO_1052 (O_1052,N_29858,N_29592);
nand UO_1053 (O_1053,N_29534,N_29839);
and UO_1054 (O_1054,N_29902,N_29665);
nor UO_1055 (O_1055,N_29766,N_29560);
nand UO_1056 (O_1056,N_29451,N_29881);
nor UO_1057 (O_1057,N_29406,N_29866);
and UO_1058 (O_1058,N_29556,N_29838);
or UO_1059 (O_1059,N_29437,N_29815);
nor UO_1060 (O_1060,N_29887,N_29804);
and UO_1061 (O_1061,N_29936,N_29756);
nand UO_1062 (O_1062,N_29427,N_29429);
or UO_1063 (O_1063,N_29828,N_29409);
or UO_1064 (O_1064,N_29854,N_29893);
or UO_1065 (O_1065,N_29839,N_29554);
xor UO_1066 (O_1066,N_29800,N_29805);
or UO_1067 (O_1067,N_29922,N_29467);
and UO_1068 (O_1068,N_29636,N_29414);
nand UO_1069 (O_1069,N_29822,N_29531);
nand UO_1070 (O_1070,N_29660,N_29555);
xor UO_1071 (O_1071,N_29755,N_29658);
nand UO_1072 (O_1072,N_29451,N_29805);
or UO_1073 (O_1073,N_29558,N_29759);
or UO_1074 (O_1074,N_29453,N_29489);
nor UO_1075 (O_1075,N_29895,N_29621);
and UO_1076 (O_1076,N_29932,N_29555);
and UO_1077 (O_1077,N_29560,N_29732);
xnor UO_1078 (O_1078,N_29872,N_29833);
xor UO_1079 (O_1079,N_29806,N_29732);
nor UO_1080 (O_1080,N_29790,N_29573);
xor UO_1081 (O_1081,N_29440,N_29428);
or UO_1082 (O_1082,N_29539,N_29859);
xnor UO_1083 (O_1083,N_29731,N_29789);
xor UO_1084 (O_1084,N_29596,N_29657);
nor UO_1085 (O_1085,N_29797,N_29712);
xnor UO_1086 (O_1086,N_29906,N_29985);
nor UO_1087 (O_1087,N_29898,N_29807);
and UO_1088 (O_1088,N_29978,N_29860);
nand UO_1089 (O_1089,N_29759,N_29905);
nor UO_1090 (O_1090,N_29947,N_29487);
or UO_1091 (O_1091,N_29401,N_29635);
xnor UO_1092 (O_1092,N_29502,N_29839);
xor UO_1093 (O_1093,N_29632,N_29635);
xor UO_1094 (O_1094,N_29610,N_29867);
xor UO_1095 (O_1095,N_29552,N_29670);
nand UO_1096 (O_1096,N_29747,N_29946);
nand UO_1097 (O_1097,N_29878,N_29425);
xor UO_1098 (O_1098,N_29884,N_29597);
nand UO_1099 (O_1099,N_29610,N_29546);
nand UO_1100 (O_1100,N_29524,N_29746);
nor UO_1101 (O_1101,N_29633,N_29460);
or UO_1102 (O_1102,N_29627,N_29773);
nand UO_1103 (O_1103,N_29542,N_29438);
and UO_1104 (O_1104,N_29848,N_29437);
or UO_1105 (O_1105,N_29909,N_29769);
and UO_1106 (O_1106,N_29852,N_29683);
and UO_1107 (O_1107,N_29530,N_29860);
nand UO_1108 (O_1108,N_29600,N_29489);
and UO_1109 (O_1109,N_29822,N_29787);
or UO_1110 (O_1110,N_29857,N_29836);
and UO_1111 (O_1111,N_29921,N_29682);
nand UO_1112 (O_1112,N_29912,N_29973);
or UO_1113 (O_1113,N_29940,N_29635);
or UO_1114 (O_1114,N_29665,N_29432);
nor UO_1115 (O_1115,N_29715,N_29678);
xor UO_1116 (O_1116,N_29654,N_29414);
nand UO_1117 (O_1117,N_29989,N_29950);
nand UO_1118 (O_1118,N_29850,N_29845);
nand UO_1119 (O_1119,N_29908,N_29710);
nand UO_1120 (O_1120,N_29450,N_29660);
nand UO_1121 (O_1121,N_29954,N_29799);
xor UO_1122 (O_1122,N_29903,N_29771);
and UO_1123 (O_1123,N_29604,N_29856);
or UO_1124 (O_1124,N_29908,N_29887);
or UO_1125 (O_1125,N_29843,N_29579);
nor UO_1126 (O_1126,N_29644,N_29469);
nand UO_1127 (O_1127,N_29463,N_29895);
and UO_1128 (O_1128,N_29526,N_29963);
nor UO_1129 (O_1129,N_29629,N_29419);
nor UO_1130 (O_1130,N_29652,N_29924);
nor UO_1131 (O_1131,N_29940,N_29889);
and UO_1132 (O_1132,N_29904,N_29874);
nand UO_1133 (O_1133,N_29926,N_29537);
nand UO_1134 (O_1134,N_29610,N_29822);
xnor UO_1135 (O_1135,N_29917,N_29481);
or UO_1136 (O_1136,N_29873,N_29475);
xor UO_1137 (O_1137,N_29846,N_29565);
or UO_1138 (O_1138,N_29864,N_29854);
nor UO_1139 (O_1139,N_29487,N_29920);
or UO_1140 (O_1140,N_29592,N_29488);
nand UO_1141 (O_1141,N_29730,N_29554);
or UO_1142 (O_1142,N_29955,N_29791);
xnor UO_1143 (O_1143,N_29437,N_29917);
or UO_1144 (O_1144,N_29528,N_29607);
or UO_1145 (O_1145,N_29608,N_29482);
and UO_1146 (O_1146,N_29909,N_29924);
nand UO_1147 (O_1147,N_29785,N_29585);
nand UO_1148 (O_1148,N_29460,N_29779);
nand UO_1149 (O_1149,N_29444,N_29655);
or UO_1150 (O_1150,N_29784,N_29529);
or UO_1151 (O_1151,N_29980,N_29475);
and UO_1152 (O_1152,N_29930,N_29554);
and UO_1153 (O_1153,N_29793,N_29480);
or UO_1154 (O_1154,N_29905,N_29514);
nand UO_1155 (O_1155,N_29755,N_29540);
xor UO_1156 (O_1156,N_29420,N_29463);
nand UO_1157 (O_1157,N_29734,N_29506);
nand UO_1158 (O_1158,N_29953,N_29745);
nor UO_1159 (O_1159,N_29453,N_29838);
nor UO_1160 (O_1160,N_29491,N_29683);
or UO_1161 (O_1161,N_29970,N_29993);
and UO_1162 (O_1162,N_29451,N_29654);
or UO_1163 (O_1163,N_29452,N_29531);
nor UO_1164 (O_1164,N_29649,N_29434);
and UO_1165 (O_1165,N_29575,N_29579);
or UO_1166 (O_1166,N_29716,N_29483);
and UO_1167 (O_1167,N_29458,N_29645);
nand UO_1168 (O_1168,N_29595,N_29775);
and UO_1169 (O_1169,N_29814,N_29953);
nor UO_1170 (O_1170,N_29530,N_29928);
or UO_1171 (O_1171,N_29892,N_29567);
nand UO_1172 (O_1172,N_29979,N_29786);
nand UO_1173 (O_1173,N_29859,N_29700);
nand UO_1174 (O_1174,N_29704,N_29585);
nor UO_1175 (O_1175,N_29403,N_29844);
and UO_1176 (O_1176,N_29788,N_29487);
nand UO_1177 (O_1177,N_29537,N_29453);
nor UO_1178 (O_1178,N_29810,N_29685);
xor UO_1179 (O_1179,N_29898,N_29746);
nand UO_1180 (O_1180,N_29406,N_29815);
or UO_1181 (O_1181,N_29664,N_29595);
nand UO_1182 (O_1182,N_29500,N_29568);
nor UO_1183 (O_1183,N_29467,N_29804);
nand UO_1184 (O_1184,N_29494,N_29617);
nor UO_1185 (O_1185,N_29633,N_29875);
nor UO_1186 (O_1186,N_29880,N_29728);
xnor UO_1187 (O_1187,N_29986,N_29783);
nor UO_1188 (O_1188,N_29582,N_29500);
nor UO_1189 (O_1189,N_29950,N_29892);
nand UO_1190 (O_1190,N_29559,N_29811);
xnor UO_1191 (O_1191,N_29678,N_29563);
and UO_1192 (O_1192,N_29864,N_29832);
nor UO_1193 (O_1193,N_29582,N_29581);
xnor UO_1194 (O_1194,N_29725,N_29410);
nor UO_1195 (O_1195,N_29469,N_29985);
xor UO_1196 (O_1196,N_29496,N_29551);
nor UO_1197 (O_1197,N_29966,N_29854);
or UO_1198 (O_1198,N_29649,N_29722);
or UO_1199 (O_1199,N_29999,N_29556);
nor UO_1200 (O_1200,N_29842,N_29629);
or UO_1201 (O_1201,N_29599,N_29403);
and UO_1202 (O_1202,N_29847,N_29979);
and UO_1203 (O_1203,N_29683,N_29682);
nor UO_1204 (O_1204,N_29743,N_29898);
xnor UO_1205 (O_1205,N_29537,N_29505);
xor UO_1206 (O_1206,N_29625,N_29618);
or UO_1207 (O_1207,N_29981,N_29995);
or UO_1208 (O_1208,N_29900,N_29459);
or UO_1209 (O_1209,N_29631,N_29756);
nand UO_1210 (O_1210,N_29831,N_29908);
xor UO_1211 (O_1211,N_29680,N_29467);
or UO_1212 (O_1212,N_29939,N_29578);
or UO_1213 (O_1213,N_29931,N_29964);
xor UO_1214 (O_1214,N_29782,N_29894);
nand UO_1215 (O_1215,N_29783,N_29640);
xor UO_1216 (O_1216,N_29683,N_29893);
and UO_1217 (O_1217,N_29514,N_29915);
nand UO_1218 (O_1218,N_29577,N_29613);
nand UO_1219 (O_1219,N_29721,N_29438);
nand UO_1220 (O_1220,N_29885,N_29982);
nor UO_1221 (O_1221,N_29531,N_29734);
nor UO_1222 (O_1222,N_29811,N_29779);
or UO_1223 (O_1223,N_29791,N_29435);
xor UO_1224 (O_1224,N_29579,N_29528);
and UO_1225 (O_1225,N_29761,N_29951);
nand UO_1226 (O_1226,N_29873,N_29596);
and UO_1227 (O_1227,N_29757,N_29720);
and UO_1228 (O_1228,N_29584,N_29486);
or UO_1229 (O_1229,N_29937,N_29655);
nor UO_1230 (O_1230,N_29993,N_29689);
and UO_1231 (O_1231,N_29955,N_29531);
nand UO_1232 (O_1232,N_29565,N_29681);
xnor UO_1233 (O_1233,N_29804,N_29652);
or UO_1234 (O_1234,N_29418,N_29915);
nand UO_1235 (O_1235,N_29789,N_29747);
nor UO_1236 (O_1236,N_29599,N_29785);
nor UO_1237 (O_1237,N_29704,N_29601);
xor UO_1238 (O_1238,N_29666,N_29758);
xnor UO_1239 (O_1239,N_29969,N_29931);
and UO_1240 (O_1240,N_29811,N_29455);
xor UO_1241 (O_1241,N_29683,N_29501);
nor UO_1242 (O_1242,N_29884,N_29433);
and UO_1243 (O_1243,N_29537,N_29618);
nor UO_1244 (O_1244,N_29899,N_29557);
nand UO_1245 (O_1245,N_29546,N_29607);
xnor UO_1246 (O_1246,N_29962,N_29526);
xnor UO_1247 (O_1247,N_29778,N_29591);
and UO_1248 (O_1248,N_29796,N_29628);
xor UO_1249 (O_1249,N_29838,N_29885);
or UO_1250 (O_1250,N_29983,N_29906);
nor UO_1251 (O_1251,N_29499,N_29743);
and UO_1252 (O_1252,N_29986,N_29880);
nand UO_1253 (O_1253,N_29873,N_29513);
xor UO_1254 (O_1254,N_29867,N_29580);
xnor UO_1255 (O_1255,N_29814,N_29945);
xor UO_1256 (O_1256,N_29674,N_29444);
nor UO_1257 (O_1257,N_29694,N_29898);
or UO_1258 (O_1258,N_29823,N_29739);
and UO_1259 (O_1259,N_29709,N_29903);
nor UO_1260 (O_1260,N_29459,N_29886);
or UO_1261 (O_1261,N_29516,N_29679);
xnor UO_1262 (O_1262,N_29510,N_29711);
or UO_1263 (O_1263,N_29488,N_29533);
and UO_1264 (O_1264,N_29880,N_29844);
and UO_1265 (O_1265,N_29932,N_29879);
xnor UO_1266 (O_1266,N_29781,N_29478);
nor UO_1267 (O_1267,N_29938,N_29655);
nand UO_1268 (O_1268,N_29679,N_29546);
xor UO_1269 (O_1269,N_29705,N_29708);
or UO_1270 (O_1270,N_29606,N_29699);
and UO_1271 (O_1271,N_29458,N_29779);
xnor UO_1272 (O_1272,N_29877,N_29616);
xnor UO_1273 (O_1273,N_29462,N_29990);
nor UO_1274 (O_1274,N_29833,N_29929);
or UO_1275 (O_1275,N_29874,N_29717);
and UO_1276 (O_1276,N_29490,N_29972);
nor UO_1277 (O_1277,N_29684,N_29490);
and UO_1278 (O_1278,N_29877,N_29808);
nor UO_1279 (O_1279,N_29709,N_29563);
nand UO_1280 (O_1280,N_29771,N_29764);
nand UO_1281 (O_1281,N_29866,N_29937);
nor UO_1282 (O_1282,N_29436,N_29966);
and UO_1283 (O_1283,N_29685,N_29969);
nand UO_1284 (O_1284,N_29711,N_29859);
nor UO_1285 (O_1285,N_29655,N_29489);
xnor UO_1286 (O_1286,N_29459,N_29442);
and UO_1287 (O_1287,N_29927,N_29992);
nand UO_1288 (O_1288,N_29612,N_29501);
or UO_1289 (O_1289,N_29485,N_29589);
or UO_1290 (O_1290,N_29800,N_29443);
or UO_1291 (O_1291,N_29449,N_29945);
nand UO_1292 (O_1292,N_29436,N_29415);
nand UO_1293 (O_1293,N_29965,N_29777);
or UO_1294 (O_1294,N_29584,N_29747);
nand UO_1295 (O_1295,N_29525,N_29748);
xor UO_1296 (O_1296,N_29601,N_29471);
nand UO_1297 (O_1297,N_29763,N_29719);
nand UO_1298 (O_1298,N_29497,N_29969);
or UO_1299 (O_1299,N_29584,N_29890);
and UO_1300 (O_1300,N_29654,N_29963);
or UO_1301 (O_1301,N_29456,N_29482);
nor UO_1302 (O_1302,N_29839,N_29854);
nor UO_1303 (O_1303,N_29411,N_29692);
nor UO_1304 (O_1304,N_29627,N_29403);
nand UO_1305 (O_1305,N_29975,N_29848);
or UO_1306 (O_1306,N_29563,N_29528);
or UO_1307 (O_1307,N_29768,N_29942);
or UO_1308 (O_1308,N_29677,N_29665);
or UO_1309 (O_1309,N_29727,N_29659);
xnor UO_1310 (O_1310,N_29424,N_29831);
xnor UO_1311 (O_1311,N_29592,N_29477);
and UO_1312 (O_1312,N_29405,N_29812);
nor UO_1313 (O_1313,N_29474,N_29767);
nor UO_1314 (O_1314,N_29994,N_29881);
or UO_1315 (O_1315,N_29902,N_29746);
nand UO_1316 (O_1316,N_29690,N_29932);
or UO_1317 (O_1317,N_29808,N_29793);
or UO_1318 (O_1318,N_29475,N_29806);
nor UO_1319 (O_1319,N_29478,N_29413);
and UO_1320 (O_1320,N_29427,N_29417);
and UO_1321 (O_1321,N_29732,N_29900);
or UO_1322 (O_1322,N_29760,N_29403);
nand UO_1323 (O_1323,N_29701,N_29675);
and UO_1324 (O_1324,N_29772,N_29691);
and UO_1325 (O_1325,N_29732,N_29690);
and UO_1326 (O_1326,N_29545,N_29758);
xor UO_1327 (O_1327,N_29661,N_29653);
and UO_1328 (O_1328,N_29814,N_29928);
nor UO_1329 (O_1329,N_29589,N_29883);
nand UO_1330 (O_1330,N_29791,N_29463);
nand UO_1331 (O_1331,N_29754,N_29568);
nand UO_1332 (O_1332,N_29702,N_29556);
or UO_1333 (O_1333,N_29945,N_29876);
nor UO_1334 (O_1334,N_29661,N_29716);
nand UO_1335 (O_1335,N_29757,N_29528);
nor UO_1336 (O_1336,N_29888,N_29801);
and UO_1337 (O_1337,N_29765,N_29618);
nand UO_1338 (O_1338,N_29816,N_29694);
or UO_1339 (O_1339,N_29715,N_29651);
or UO_1340 (O_1340,N_29700,N_29865);
or UO_1341 (O_1341,N_29494,N_29737);
nor UO_1342 (O_1342,N_29722,N_29482);
xnor UO_1343 (O_1343,N_29491,N_29456);
xnor UO_1344 (O_1344,N_29880,N_29969);
and UO_1345 (O_1345,N_29796,N_29717);
nor UO_1346 (O_1346,N_29600,N_29620);
nand UO_1347 (O_1347,N_29932,N_29989);
and UO_1348 (O_1348,N_29655,N_29663);
nand UO_1349 (O_1349,N_29427,N_29878);
nand UO_1350 (O_1350,N_29521,N_29472);
or UO_1351 (O_1351,N_29902,N_29913);
nand UO_1352 (O_1352,N_29467,N_29937);
xnor UO_1353 (O_1353,N_29645,N_29795);
nand UO_1354 (O_1354,N_29666,N_29489);
and UO_1355 (O_1355,N_29594,N_29701);
xor UO_1356 (O_1356,N_29720,N_29461);
nor UO_1357 (O_1357,N_29603,N_29518);
xnor UO_1358 (O_1358,N_29563,N_29587);
nand UO_1359 (O_1359,N_29418,N_29951);
xor UO_1360 (O_1360,N_29520,N_29961);
nand UO_1361 (O_1361,N_29845,N_29653);
xnor UO_1362 (O_1362,N_29968,N_29712);
and UO_1363 (O_1363,N_29718,N_29968);
nor UO_1364 (O_1364,N_29590,N_29629);
xor UO_1365 (O_1365,N_29612,N_29510);
xor UO_1366 (O_1366,N_29856,N_29997);
nand UO_1367 (O_1367,N_29947,N_29471);
and UO_1368 (O_1368,N_29987,N_29955);
xor UO_1369 (O_1369,N_29484,N_29589);
nor UO_1370 (O_1370,N_29515,N_29729);
nor UO_1371 (O_1371,N_29901,N_29992);
and UO_1372 (O_1372,N_29495,N_29510);
and UO_1373 (O_1373,N_29857,N_29789);
nand UO_1374 (O_1374,N_29856,N_29669);
and UO_1375 (O_1375,N_29709,N_29889);
and UO_1376 (O_1376,N_29896,N_29433);
nand UO_1377 (O_1377,N_29812,N_29683);
and UO_1378 (O_1378,N_29603,N_29404);
xor UO_1379 (O_1379,N_29817,N_29654);
nor UO_1380 (O_1380,N_29542,N_29965);
nor UO_1381 (O_1381,N_29888,N_29940);
and UO_1382 (O_1382,N_29644,N_29523);
nor UO_1383 (O_1383,N_29458,N_29530);
xnor UO_1384 (O_1384,N_29909,N_29505);
nor UO_1385 (O_1385,N_29781,N_29870);
nand UO_1386 (O_1386,N_29566,N_29505);
nand UO_1387 (O_1387,N_29458,N_29938);
and UO_1388 (O_1388,N_29401,N_29702);
nor UO_1389 (O_1389,N_29614,N_29927);
or UO_1390 (O_1390,N_29935,N_29659);
nor UO_1391 (O_1391,N_29943,N_29429);
nand UO_1392 (O_1392,N_29947,N_29831);
nor UO_1393 (O_1393,N_29418,N_29600);
or UO_1394 (O_1394,N_29892,N_29992);
or UO_1395 (O_1395,N_29992,N_29822);
nand UO_1396 (O_1396,N_29446,N_29505);
and UO_1397 (O_1397,N_29645,N_29474);
or UO_1398 (O_1398,N_29825,N_29433);
nand UO_1399 (O_1399,N_29497,N_29412);
nand UO_1400 (O_1400,N_29675,N_29454);
nor UO_1401 (O_1401,N_29554,N_29537);
xnor UO_1402 (O_1402,N_29958,N_29675);
nor UO_1403 (O_1403,N_29687,N_29780);
and UO_1404 (O_1404,N_29605,N_29926);
xnor UO_1405 (O_1405,N_29676,N_29506);
and UO_1406 (O_1406,N_29415,N_29490);
and UO_1407 (O_1407,N_29451,N_29526);
nand UO_1408 (O_1408,N_29611,N_29448);
nor UO_1409 (O_1409,N_29787,N_29400);
xor UO_1410 (O_1410,N_29969,N_29938);
xor UO_1411 (O_1411,N_29669,N_29778);
xnor UO_1412 (O_1412,N_29955,N_29892);
xor UO_1413 (O_1413,N_29557,N_29414);
and UO_1414 (O_1414,N_29533,N_29520);
nand UO_1415 (O_1415,N_29688,N_29565);
or UO_1416 (O_1416,N_29702,N_29568);
nor UO_1417 (O_1417,N_29635,N_29687);
xnor UO_1418 (O_1418,N_29807,N_29447);
and UO_1419 (O_1419,N_29862,N_29711);
or UO_1420 (O_1420,N_29780,N_29407);
or UO_1421 (O_1421,N_29904,N_29934);
nand UO_1422 (O_1422,N_29784,N_29928);
xor UO_1423 (O_1423,N_29582,N_29812);
nor UO_1424 (O_1424,N_29539,N_29784);
nand UO_1425 (O_1425,N_29566,N_29535);
and UO_1426 (O_1426,N_29559,N_29944);
nand UO_1427 (O_1427,N_29913,N_29640);
xnor UO_1428 (O_1428,N_29638,N_29939);
or UO_1429 (O_1429,N_29766,N_29624);
and UO_1430 (O_1430,N_29784,N_29892);
nand UO_1431 (O_1431,N_29908,N_29524);
xnor UO_1432 (O_1432,N_29528,N_29668);
nor UO_1433 (O_1433,N_29456,N_29667);
and UO_1434 (O_1434,N_29916,N_29541);
xor UO_1435 (O_1435,N_29562,N_29873);
nand UO_1436 (O_1436,N_29899,N_29814);
xor UO_1437 (O_1437,N_29656,N_29516);
nor UO_1438 (O_1438,N_29694,N_29819);
nand UO_1439 (O_1439,N_29570,N_29705);
nand UO_1440 (O_1440,N_29787,N_29980);
or UO_1441 (O_1441,N_29481,N_29652);
nand UO_1442 (O_1442,N_29531,N_29873);
nor UO_1443 (O_1443,N_29997,N_29427);
nor UO_1444 (O_1444,N_29480,N_29727);
nand UO_1445 (O_1445,N_29491,N_29777);
nand UO_1446 (O_1446,N_29758,N_29985);
nor UO_1447 (O_1447,N_29595,N_29515);
and UO_1448 (O_1448,N_29881,N_29581);
or UO_1449 (O_1449,N_29528,N_29755);
nand UO_1450 (O_1450,N_29777,N_29790);
nand UO_1451 (O_1451,N_29836,N_29796);
nand UO_1452 (O_1452,N_29975,N_29597);
nor UO_1453 (O_1453,N_29612,N_29963);
nand UO_1454 (O_1454,N_29965,N_29530);
and UO_1455 (O_1455,N_29787,N_29805);
or UO_1456 (O_1456,N_29847,N_29476);
and UO_1457 (O_1457,N_29755,N_29534);
nor UO_1458 (O_1458,N_29636,N_29807);
nand UO_1459 (O_1459,N_29490,N_29982);
or UO_1460 (O_1460,N_29920,N_29676);
or UO_1461 (O_1461,N_29412,N_29991);
nand UO_1462 (O_1462,N_29884,N_29532);
and UO_1463 (O_1463,N_29852,N_29467);
xor UO_1464 (O_1464,N_29812,N_29530);
nand UO_1465 (O_1465,N_29567,N_29641);
or UO_1466 (O_1466,N_29595,N_29514);
xor UO_1467 (O_1467,N_29661,N_29476);
and UO_1468 (O_1468,N_29934,N_29628);
and UO_1469 (O_1469,N_29864,N_29995);
nor UO_1470 (O_1470,N_29790,N_29835);
and UO_1471 (O_1471,N_29552,N_29404);
or UO_1472 (O_1472,N_29453,N_29944);
nand UO_1473 (O_1473,N_29590,N_29470);
nor UO_1474 (O_1474,N_29796,N_29557);
nor UO_1475 (O_1475,N_29463,N_29861);
nand UO_1476 (O_1476,N_29473,N_29615);
nand UO_1477 (O_1477,N_29505,N_29435);
or UO_1478 (O_1478,N_29424,N_29875);
or UO_1479 (O_1479,N_29761,N_29687);
nand UO_1480 (O_1480,N_29980,N_29680);
nor UO_1481 (O_1481,N_29957,N_29531);
nand UO_1482 (O_1482,N_29626,N_29894);
nand UO_1483 (O_1483,N_29905,N_29813);
and UO_1484 (O_1484,N_29564,N_29483);
nor UO_1485 (O_1485,N_29888,N_29506);
nand UO_1486 (O_1486,N_29945,N_29810);
and UO_1487 (O_1487,N_29645,N_29638);
and UO_1488 (O_1488,N_29872,N_29432);
and UO_1489 (O_1489,N_29752,N_29854);
and UO_1490 (O_1490,N_29970,N_29910);
nor UO_1491 (O_1491,N_29490,N_29823);
xnor UO_1492 (O_1492,N_29891,N_29787);
nand UO_1493 (O_1493,N_29807,N_29690);
and UO_1494 (O_1494,N_29658,N_29962);
nor UO_1495 (O_1495,N_29779,N_29969);
nand UO_1496 (O_1496,N_29735,N_29566);
and UO_1497 (O_1497,N_29863,N_29948);
and UO_1498 (O_1498,N_29786,N_29595);
and UO_1499 (O_1499,N_29892,N_29428);
nand UO_1500 (O_1500,N_29715,N_29438);
nor UO_1501 (O_1501,N_29910,N_29737);
xor UO_1502 (O_1502,N_29917,N_29708);
nand UO_1503 (O_1503,N_29647,N_29598);
and UO_1504 (O_1504,N_29708,N_29547);
nand UO_1505 (O_1505,N_29777,N_29976);
nand UO_1506 (O_1506,N_29484,N_29812);
xor UO_1507 (O_1507,N_29481,N_29682);
nand UO_1508 (O_1508,N_29636,N_29681);
or UO_1509 (O_1509,N_29454,N_29715);
and UO_1510 (O_1510,N_29669,N_29792);
nor UO_1511 (O_1511,N_29621,N_29554);
and UO_1512 (O_1512,N_29468,N_29432);
and UO_1513 (O_1513,N_29619,N_29495);
and UO_1514 (O_1514,N_29979,N_29940);
nand UO_1515 (O_1515,N_29805,N_29955);
and UO_1516 (O_1516,N_29574,N_29715);
nand UO_1517 (O_1517,N_29821,N_29888);
nand UO_1518 (O_1518,N_29447,N_29638);
xor UO_1519 (O_1519,N_29904,N_29632);
or UO_1520 (O_1520,N_29799,N_29769);
and UO_1521 (O_1521,N_29519,N_29662);
or UO_1522 (O_1522,N_29456,N_29459);
or UO_1523 (O_1523,N_29914,N_29923);
or UO_1524 (O_1524,N_29652,N_29653);
or UO_1525 (O_1525,N_29966,N_29613);
or UO_1526 (O_1526,N_29691,N_29615);
or UO_1527 (O_1527,N_29979,N_29611);
xor UO_1528 (O_1528,N_29438,N_29552);
xor UO_1529 (O_1529,N_29692,N_29964);
nand UO_1530 (O_1530,N_29648,N_29539);
and UO_1531 (O_1531,N_29753,N_29971);
and UO_1532 (O_1532,N_29821,N_29607);
or UO_1533 (O_1533,N_29673,N_29784);
xnor UO_1534 (O_1534,N_29747,N_29859);
or UO_1535 (O_1535,N_29737,N_29781);
or UO_1536 (O_1536,N_29904,N_29464);
and UO_1537 (O_1537,N_29891,N_29536);
and UO_1538 (O_1538,N_29615,N_29601);
and UO_1539 (O_1539,N_29980,N_29711);
or UO_1540 (O_1540,N_29558,N_29672);
nor UO_1541 (O_1541,N_29890,N_29757);
nand UO_1542 (O_1542,N_29676,N_29717);
xnor UO_1543 (O_1543,N_29546,N_29545);
nand UO_1544 (O_1544,N_29587,N_29843);
xor UO_1545 (O_1545,N_29877,N_29956);
and UO_1546 (O_1546,N_29960,N_29930);
nor UO_1547 (O_1547,N_29685,N_29565);
nor UO_1548 (O_1548,N_29412,N_29526);
nand UO_1549 (O_1549,N_29717,N_29979);
nand UO_1550 (O_1550,N_29971,N_29949);
and UO_1551 (O_1551,N_29780,N_29490);
nor UO_1552 (O_1552,N_29649,N_29897);
or UO_1553 (O_1553,N_29523,N_29572);
nor UO_1554 (O_1554,N_29644,N_29617);
nor UO_1555 (O_1555,N_29870,N_29772);
and UO_1556 (O_1556,N_29690,N_29521);
xnor UO_1557 (O_1557,N_29967,N_29410);
nand UO_1558 (O_1558,N_29566,N_29821);
xor UO_1559 (O_1559,N_29664,N_29735);
and UO_1560 (O_1560,N_29886,N_29767);
or UO_1561 (O_1561,N_29963,N_29814);
nor UO_1562 (O_1562,N_29554,N_29419);
nor UO_1563 (O_1563,N_29988,N_29750);
xor UO_1564 (O_1564,N_29579,N_29465);
nand UO_1565 (O_1565,N_29796,N_29815);
or UO_1566 (O_1566,N_29925,N_29503);
nor UO_1567 (O_1567,N_29464,N_29420);
and UO_1568 (O_1568,N_29877,N_29730);
and UO_1569 (O_1569,N_29712,N_29724);
and UO_1570 (O_1570,N_29445,N_29535);
xor UO_1571 (O_1571,N_29453,N_29824);
or UO_1572 (O_1572,N_29960,N_29764);
nor UO_1573 (O_1573,N_29836,N_29551);
or UO_1574 (O_1574,N_29688,N_29435);
xnor UO_1575 (O_1575,N_29404,N_29558);
xor UO_1576 (O_1576,N_29480,N_29583);
or UO_1577 (O_1577,N_29873,N_29563);
or UO_1578 (O_1578,N_29899,N_29980);
xor UO_1579 (O_1579,N_29510,N_29815);
or UO_1580 (O_1580,N_29863,N_29762);
nand UO_1581 (O_1581,N_29443,N_29524);
nor UO_1582 (O_1582,N_29534,N_29983);
nand UO_1583 (O_1583,N_29506,N_29484);
and UO_1584 (O_1584,N_29443,N_29649);
nand UO_1585 (O_1585,N_29681,N_29439);
xnor UO_1586 (O_1586,N_29557,N_29873);
xnor UO_1587 (O_1587,N_29735,N_29881);
nor UO_1588 (O_1588,N_29722,N_29622);
nand UO_1589 (O_1589,N_29628,N_29743);
or UO_1590 (O_1590,N_29869,N_29606);
xor UO_1591 (O_1591,N_29855,N_29640);
nand UO_1592 (O_1592,N_29825,N_29822);
or UO_1593 (O_1593,N_29952,N_29635);
nor UO_1594 (O_1594,N_29646,N_29893);
or UO_1595 (O_1595,N_29444,N_29688);
or UO_1596 (O_1596,N_29983,N_29728);
and UO_1597 (O_1597,N_29563,N_29816);
and UO_1598 (O_1598,N_29582,N_29678);
xor UO_1599 (O_1599,N_29763,N_29618);
nand UO_1600 (O_1600,N_29738,N_29584);
or UO_1601 (O_1601,N_29603,N_29859);
xnor UO_1602 (O_1602,N_29459,N_29693);
xor UO_1603 (O_1603,N_29999,N_29708);
or UO_1604 (O_1604,N_29705,N_29714);
and UO_1605 (O_1605,N_29671,N_29692);
nand UO_1606 (O_1606,N_29651,N_29559);
nand UO_1607 (O_1607,N_29819,N_29792);
xor UO_1608 (O_1608,N_29964,N_29684);
or UO_1609 (O_1609,N_29462,N_29708);
nand UO_1610 (O_1610,N_29677,N_29457);
nor UO_1611 (O_1611,N_29421,N_29518);
nand UO_1612 (O_1612,N_29948,N_29925);
xnor UO_1613 (O_1613,N_29913,N_29915);
or UO_1614 (O_1614,N_29741,N_29798);
nand UO_1615 (O_1615,N_29544,N_29767);
and UO_1616 (O_1616,N_29672,N_29767);
nand UO_1617 (O_1617,N_29483,N_29614);
or UO_1618 (O_1618,N_29436,N_29826);
and UO_1619 (O_1619,N_29590,N_29661);
and UO_1620 (O_1620,N_29956,N_29555);
nor UO_1621 (O_1621,N_29837,N_29905);
xnor UO_1622 (O_1622,N_29983,N_29750);
nand UO_1623 (O_1623,N_29691,N_29849);
and UO_1624 (O_1624,N_29602,N_29733);
or UO_1625 (O_1625,N_29449,N_29760);
and UO_1626 (O_1626,N_29978,N_29698);
xnor UO_1627 (O_1627,N_29847,N_29598);
nor UO_1628 (O_1628,N_29766,N_29489);
nor UO_1629 (O_1629,N_29788,N_29462);
and UO_1630 (O_1630,N_29562,N_29844);
and UO_1631 (O_1631,N_29731,N_29513);
nand UO_1632 (O_1632,N_29402,N_29545);
nand UO_1633 (O_1633,N_29671,N_29470);
nand UO_1634 (O_1634,N_29416,N_29721);
xnor UO_1635 (O_1635,N_29998,N_29817);
or UO_1636 (O_1636,N_29648,N_29913);
and UO_1637 (O_1637,N_29793,N_29589);
nor UO_1638 (O_1638,N_29613,N_29741);
nand UO_1639 (O_1639,N_29932,N_29854);
and UO_1640 (O_1640,N_29554,N_29483);
and UO_1641 (O_1641,N_29820,N_29836);
nor UO_1642 (O_1642,N_29647,N_29958);
and UO_1643 (O_1643,N_29719,N_29998);
and UO_1644 (O_1644,N_29727,N_29655);
xnor UO_1645 (O_1645,N_29485,N_29645);
xnor UO_1646 (O_1646,N_29728,N_29864);
xnor UO_1647 (O_1647,N_29667,N_29926);
or UO_1648 (O_1648,N_29534,N_29526);
nand UO_1649 (O_1649,N_29639,N_29644);
or UO_1650 (O_1650,N_29487,N_29630);
or UO_1651 (O_1651,N_29929,N_29886);
or UO_1652 (O_1652,N_29810,N_29656);
nor UO_1653 (O_1653,N_29978,N_29498);
nand UO_1654 (O_1654,N_29920,N_29662);
nand UO_1655 (O_1655,N_29681,N_29982);
nor UO_1656 (O_1656,N_29976,N_29481);
and UO_1657 (O_1657,N_29846,N_29764);
xnor UO_1658 (O_1658,N_29896,N_29922);
nor UO_1659 (O_1659,N_29657,N_29527);
xor UO_1660 (O_1660,N_29678,N_29451);
xnor UO_1661 (O_1661,N_29889,N_29577);
or UO_1662 (O_1662,N_29406,N_29735);
nand UO_1663 (O_1663,N_29611,N_29407);
nand UO_1664 (O_1664,N_29867,N_29758);
or UO_1665 (O_1665,N_29939,N_29691);
nor UO_1666 (O_1666,N_29628,N_29495);
nand UO_1667 (O_1667,N_29749,N_29630);
and UO_1668 (O_1668,N_29853,N_29513);
nand UO_1669 (O_1669,N_29420,N_29827);
nand UO_1670 (O_1670,N_29815,N_29897);
nor UO_1671 (O_1671,N_29630,N_29605);
xnor UO_1672 (O_1672,N_29896,N_29613);
and UO_1673 (O_1673,N_29567,N_29566);
and UO_1674 (O_1674,N_29580,N_29649);
nor UO_1675 (O_1675,N_29472,N_29571);
or UO_1676 (O_1676,N_29765,N_29739);
xnor UO_1677 (O_1677,N_29703,N_29890);
and UO_1678 (O_1678,N_29413,N_29664);
nor UO_1679 (O_1679,N_29921,N_29471);
nand UO_1680 (O_1680,N_29515,N_29873);
xnor UO_1681 (O_1681,N_29793,N_29892);
and UO_1682 (O_1682,N_29674,N_29931);
xnor UO_1683 (O_1683,N_29575,N_29967);
and UO_1684 (O_1684,N_29498,N_29469);
or UO_1685 (O_1685,N_29982,N_29559);
or UO_1686 (O_1686,N_29460,N_29900);
xor UO_1687 (O_1687,N_29955,N_29840);
or UO_1688 (O_1688,N_29715,N_29800);
nor UO_1689 (O_1689,N_29782,N_29969);
nor UO_1690 (O_1690,N_29914,N_29438);
nor UO_1691 (O_1691,N_29809,N_29685);
or UO_1692 (O_1692,N_29743,N_29865);
nand UO_1693 (O_1693,N_29410,N_29769);
and UO_1694 (O_1694,N_29930,N_29802);
nor UO_1695 (O_1695,N_29761,N_29965);
nor UO_1696 (O_1696,N_29844,N_29752);
nand UO_1697 (O_1697,N_29940,N_29428);
nor UO_1698 (O_1698,N_29452,N_29430);
xor UO_1699 (O_1699,N_29697,N_29813);
nor UO_1700 (O_1700,N_29883,N_29882);
nor UO_1701 (O_1701,N_29406,N_29774);
xnor UO_1702 (O_1702,N_29597,N_29668);
or UO_1703 (O_1703,N_29714,N_29757);
xnor UO_1704 (O_1704,N_29511,N_29599);
xor UO_1705 (O_1705,N_29917,N_29841);
or UO_1706 (O_1706,N_29417,N_29765);
or UO_1707 (O_1707,N_29870,N_29850);
nor UO_1708 (O_1708,N_29442,N_29861);
xnor UO_1709 (O_1709,N_29843,N_29607);
xnor UO_1710 (O_1710,N_29431,N_29841);
nor UO_1711 (O_1711,N_29626,N_29680);
nor UO_1712 (O_1712,N_29637,N_29402);
nand UO_1713 (O_1713,N_29634,N_29897);
nor UO_1714 (O_1714,N_29600,N_29981);
and UO_1715 (O_1715,N_29473,N_29746);
xnor UO_1716 (O_1716,N_29993,N_29838);
or UO_1717 (O_1717,N_29701,N_29553);
or UO_1718 (O_1718,N_29615,N_29692);
and UO_1719 (O_1719,N_29668,N_29624);
and UO_1720 (O_1720,N_29886,N_29563);
nand UO_1721 (O_1721,N_29596,N_29928);
nand UO_1722 (O_1722,N_29819,N_29705);
and UO_1723 (O_1723,N_29961,N_29892);
nor UO_1724 (O_1724,N_29837,N_29914);
nand UO_1725 (O_1725,N_29693,N_29831);
xnor UO_1726 (O_1726,N_29703,N_29494);
nand UO_1727 (O_1727,N_29719,N_29549);
or UO_1728 (O_1728,N_29687,N_29480);
xor UO_1729 (O_1729,N_29459,N_29595);
nand UO_1730 (O_1730,N_29579,N_29463);
nor UO_1731 (O_1731,N_29795,N_29736);
xnor UO_1732 (O_1732,N_29844,N_29855);
nand UO_1733 (O_1733,N_29642,N_29933);
nor UO_1734 (O_1734,N_29510,N_29992);
or UO_1735 (O_1735,N_29938,N_29790);
nand UO_1736 (O_1736,N_29404,N_29443);
and UO_1737 (O_1737,N_29803,N_29985);
nor UO_1738 (O_1738,N_29482,N_29801);
xnor UO_1739 (O_1739,N_29652,N_29922);
nand UO_1740 (O_1740,N_29557,N_29955);
and UO_1741 (O_1741,N_29418,N_29976);
nand UO_1742 (O_1742,N_29406,N_29767);
nor UO_1743 (O_1743,N_29969,N_29525);
nor UO_1744 (O_1744,N_29573,N_29851);
nand UO_1745 (O_1745,N_29958,N_29665);
nor UO_1746 (O_1746,N_29792,N_29836);
xnor UO_1747 (O_1747,N_29527,N_29678);
and UO_1748 (O_1748,N_29818,N_29733);
and UO_1749 (O_1749,N_29406,N_29770);
and UO_1750 (O_1750,N_29658,N_29801);
nand UO_1751 (O_1751,N_29962,N_29835);
nand UO_1752 (O_1752,N_29873,N_29929);
nand UO_1753 (O_1753,N_29682,N_29688);
or UO_1754 (O_1754,N_29479,N_29658);
nand UO_1755 (O_1755,N_29406,N_29915);
and UO_1756 (O_1756,N_29676,N_29970);
xnor UO_1757 (O_1757,N_29739,N_29958);
or UO_1758 (O_1758,N_29687,N_29845);
nand UO_1759 (O_1759,N_29435,N_29694);
and UO_1760 (O_1760,N_29519,N_29453);
xnor UO_1761 (O_1761,N_29686,N_29647);
or UO_1762 (O_1762,N_29470,N_29976);
nor UO_1763 (O_1763,N_29456,N_29722);
nor UO_1764 (O_1764,N_29547,N_29451);
nand UO_1765 (O_1765,N_29820,N_29457);
xor UO_1766 (O_1766,N_29453,N_29586);
and UO_1767 (O_1767,N_29788,N_29860);
or UO_1768 (O_1768,N_29667,N_29424);
and UO_1769 (O_1769,N_29952,N_29440);
nor UO_1770 (O_1770,N_29760,N_29616);
xor UO_1771 (O_1771,N_29712,N_29659);
nand UO_1772 (O_1772,N_29715,N_29928);
xnor UO_1773 (O_1773,N_29657,N_29663);
or UO_1774 (O_1774,N_29856,N_29586);
nor UO_1775 (O_1775,N_29700,N_29672);
nand UO_1776 (O_1776,N_29922,N_29781);
nand UO_1777 (O_1777,N_29867,N_29502);
nand UO_1778 (O_1778,N_29859,N_29898);
or UO_1779 (O_1779,N_29750,N_29593);
nor UO_1780 (O_1780,N_29641,N_29573);
and UO_1781 (O_1781,N_29798,N_29976);
xnor UO_1782 (O_1782,N_29880,N_29582);
nand UO_1783 (O_1783,N_29566,N_29413);
nor UO_1784 (O_1784,N_29503,N_29608);
or UO_1785 (O_1785,N_29844,N_29737);
xor UO_1786 (O_1786,N_29558,N_29764);
nor UO_1787 (O_1787,N_29587,N_29471);
nor UO_1788 (O_1788,N_29616,N_29403);
xor UO_1789 (O_1789,N_29471,N_29766);
or UO_1790 (O_1790,N_29466,N_29403);
nand UO_1791 (O_1791,N_29843,N_29701);
nor UO_1792 (O_1792,N_29419,N_29796);
xor UO_1793 (O_1793,N_29993,N_29418);
and UO_1794 (O_1794,N_29582,N_29779);
and UO_1795 (O_1795,N_29718,N_29508);
nand UO_1796 (O_1796,N_29606,N_29977);
xnor UO_1797 (O_1797,N_29928,N_29400);
nor UO_1798 (O_1798,N_29860,N_29770);
xor UO_1799 (O_1799,N_29797,N_29564);
nand UO_1800 (O_1800,N_29643,N_29725);
nand UO_1801 (O_1801,N_29641,N_29799);
or UO_1802 (O_1802,N_29446,N_29556);
nand UO_1803 (O_1803,N_29535,N_29792);
and UO_1804 (O_1804,N_29485,N_29534);
nor UO_1805 (O_1805,N_29435,N_29685);
nor UO_1806 (O_1806,N_29649,N_29560);
or UO_1807 (O_1807,N_29467,N_29904);
nand UO_1808 (O_1808,N_29542,N_29498);
xnor UO_1809 (O_1809,N_29855,N_29894);
nand UO_1810 (O_1810,N_29826,N_29797);
nand UO_1811 (O_1811,N_29541,N_29430);
nor UO_1812 (O_1812,N_29511,N_29429);
nor UO_1813 (O_1813,N_29585,N_29683);
or UO_1814 (O_1814,N_29935,N_29861);
nor UO_1815 (O_1815,N_29465,N_29667);
nand UO_1816 (O_1816,N_29853,N_29419);
nor UO_1817 (O_1817,N_29779,N_29888);
xnor UO_1818 (O_1818,N_29716,N_29810);
or UO_1819 (O_1819,N_29498,N_29696);
xnor UO_1820 (O_1820,N_29440,N_29777);
or UO_1821 (O_1821,N_29599,N_29953);
nor UO_1822 (O_1822,N_29570,N_29444);
nand UO_1823 (O_1823,N_29612,N_29680);
xnor UO_1824 (O_1824,N_29681,N_29828);
nor UO_1825 (O_1825,N_29459,N_29562);
nand UO_1826 (O_1826,N_29880,N_29771);
nand UO_1827 (O_1827,N_29775,N_29902);
nor UO_1828 (O_1828,N_29866,N_29915);
xnor UO_1829 (O_1829,N_29491,N_29712);
nand UO_1830 (O_1830,N_29528,N_29443);
nor UO_1831 (O_1831,N_29600,N_29942);
nor UO_1832 (O_1832,N_29851,N_29918);
and UO_1833 (O_1833,N_29971,N_29650);
and UO_1834 (O_1834,N_29523,N_29954);
or UO_1835 (O_1835,N_29766,N_29815);
xnor UO_1836 (O_1836,N_29718,N_29495);
nor UO_1837 (O_1837,N_29633,N_29426);
or UO_1838 (O_1838,N_29436,N_29935);
and UO_1839 (O_1839,N_29564,N_29994);
or UO_1840 (O_1840,N_29699,N_29933);
nand UO_1841 (O_1841,N_29652,N_29494);
nand UO_1842 (O_1842,N_29708,N_29762);
xor UO_1843 (O_1843,N_29922,N_29423);
nand UO_1844 (O_1844,N_29652,N_29998);
xnor UO_1845 (O_1845,N_29783,N_29794);
nor UO_1846 (O_1846,N_29450,N_29677);
or UO_1847 (O_1847,N_29679,N_29907);
and UO_1848 (O_1848,N_29936,N_29588);
or UO_1849 (O_1849,N_29493,N_29689);
and UO_1850 (O_1850,N_29878,N_29962);
nor UO_1851 (O_1851,N_29663,N_29453);
xnor UO_1852 (O_1852,N_29767,N_29769);
or UO_1853 (O_1853,N_29483,N_29992);
xnor UO_1854 (O_1854,N_29657,N_29564);
nand UO_1855 (O_1855,N_29586,N_29906);
or UO_1856 (O_1856,N_29813,N_29736);
and UO_1857 (O_1857,N_29872,N_29624);
and UO_1858 (O_1858,N_29942,N_29826);
and UO_1859 (O_1859,N_29418,N_29856);
nor UO_1860 (O_1860,N_29476,N_29566);
xnor UO_1861 (O_1861,N_29632,N_29616);
nor UO_1862 (O_1862,N_29728,N_29409);
nand UO_1863 (O_1863,N_29895,N_29982);
nor UO_1864 (O_1864,N_29624,N_29780);
nor UO_1865 (O_1865,N_29961,N_29863);
nor UO_1866 (O_1866,N_29680,N_29862);
nand UO_1867 (O_1867,N_29760,N_29965);
nor UO_1868 (O_1868,N_29730,N_29618);
xor UO_1869 (O_1869,N_29615,N_29745);
or UO_1870 (O_1870,N_29492,N_29885);
or UO_1871 (O_1871,N_29835,N_29832);
nor UO_1872 (O_1872,N_29976,N_29971);
or UO_1873 (O_1873,N_29527,N_29711);
or UO_1874 (O_1874,N_29568,N_29646);
nand UO_1875 (O_1875,N_29709,N_29832);
xor UO_1876 (O_1876,N_29771,N_29975);
or UO_1877 (O_1877,N_29763,N_29747);
nor UO_1878 (O_1878,N_29409,N_29463);
or UO_1879 (O_1879,N_29959,N_29435);
or UO_1880 (O_1880,N_29898,N_29673);
and UO_1881 (O_1881,N_29472,N_29794);
xor UO_1882 (O_1882,N_29850,N_29748);
nand UO_1883 (O_1883,N_29955,N_29540);
or UO_1884 (O_1884,N_29746,N_29552);
nor UO_1885 (O_1885,N_29613,N_29908);
nand UO_1886 (O_1886,N_29872,N_29454);
or UO_1887 (O_1887,N_29616,N_29965);
xnor UO_1888 (O_1888,N_29567,N_29745);
nor UO_1889 (O_1889,N_29714,N_29905);
xnor UO_1890 (O_1890,N_29403,N_29674);
nand UO_1891 (O_1891,N_29466,N_29575);
or UO_1892 (O_1892,N_29957,N_29775);
nor UO_1893 (O_1893,N_29816,N_29487);
and UO_1894 (O_1894,N_29407,N_29759);
nor UO_1895 (O_1895,N_29535,N_29963);
or UO_1896 (O_1896,N_29484,N_29822);
nor UO_1897 (O_1897,N_29496,N_29447);
nand UO_1898 (O_1898,N_29806,N_29995);
nor UO_1899 (O_1899,N_29550,N_29919);
nor UO_1900 (O_1900,N_29655,N_29730);
and UO_1901 (O_1901,N_29572,N_29891);
xor UO_1902 (O_1902,N_29726,N_29930);
nand UO_1903 (O_1903,N_29955,N_29566);
or UO_1904 (O_1904,N_29406,N_29525);
nor UO_1905 (O_1905,N_29563,N_29501);
nor UO_1906 (O_1906,N_29901,N_29712);
nand UO_1907 (O_1907,N_29971,N_29616);
nand UO_1908 (O_1908,N_29694,N_29650);
and UO_1909 (O_1909,N_29672,N_29716);
xor UO_1910 (O_1910,N_29672,N_29497);
nand UO_1911 (O_1911,N_29679,N_29603);
nand UO_1912 (O_1912,N_29994,N_29595);
xor UO_1913 (O_1913,N_29525,N_29705);
or UO_1914 (O_1914,N_29401,N_29817);
xnor UO_1915 (O_1915,N_29574,N_29446);
nor UO_1916 (O_1916,N_29645,N_29753);
xnor UO_1917 (O_1917,N_29543,N_29856);
or UO_1918 (O_1918,N_29417,N_29643);
nand UO_1919 (O_1919,N_29579,N_29742);
nand UO_1920 (O_1920,N_29869,N_29695);
nor UO_1921 (O_1921,N_29590,N_29584);
nor UO_1922 (O_1922,N_29918,N_29590);
or UO_1923 (O_1923,N_29415,N_29518);
nor UO_1924 (O_1924,N_29947,N_29782);
xor UO_1925 (O_1925,N_29588,N_29791);
and UO_1926 (O_1926,N_29972,N_29961);
nand UO_1927 (O_1927,N_29470,N_29704);
nand UO_1928 (O_1928,N_29933,N_29950);
nor UO_1929 (O_1929,N_29437,N_29883);
xor UO_1930 (O_1930,N_29552,N_29918);
nand UO_1931 (O_1931,N_29931,N_29996);
xnor UO_1932 (O_1932,N_29935,N_29900);
nor UO_1933 (O_1933,N_29739,N_29461);
and UO_1934 (O_1934,N_29450,N_29937);
xnor UO_1935 (O_1935,N_29881,N_29874);
xor UO_1936 (O_1936,N_29600,N_29582);
nor UO_1937 (O_1937,N_29828,N_29797);
nand UO_1938 (O_1938,N_29536,N_29488);
and UO_1939 (O_1939,N_29987,N_29719);
nand UO_1940 (O_1940,N_29434,N_29924);
xnor UO_1941 (O_1941,N_29737,N_29738);
nand UO_1942 (O_1942,N_29619,N_29598);
and UO_1943 (O_1943,N_29511,N_29534);
xnor UO_1944 (O_1944,N_29775,N_29469);
xor UO_1945 (O_1945,N_29711,N_29727);
nand UO_1946 (O_1946,N_29885,N_29759);
nor UO_1947 (O_1947,N_29925,N_29851);
nand UO_1948 (O_1948,N_29871,N_29657);
nand UO_1949 (O_1949,N_29684,N_29825);
and UO_1950 (O_1950,N_29729,N_29648);
or UO_1951 (O_1951,N_29441,N_29566);
nand UO_1952 (O_1952,N_29601,N_29789);
and UO_1953 (O_1953,N_29687,N_29857);
xor UO_1954 (O_1954,N_29911,N_29762);
nor UO_1955 (O_1955,N_29443,N_29522);
or UO_1956 (O_1956,N_29639,N_29577);
nor UO_1957 (O_1957,N_29999,N_29840);
nor UO_1958 (O_1958,N_29804,N_29558);
or UO_1959 (O_1959,N_29723,N_29593);
or UO_1960 (O_1960,N_29568,N_29768);
or UO_1961 (O_1961,N_29994,N_29592);
nand UO_1962 (O_1962,N_29697,N_29448);
and UO_1963 (O_1963,N_29922,N_29576);
xnor UO_1964 (O_1964,N_29852,N_29838);
and UO_1965 (O_1965,N_29511,N_29559);
xnor UO_1966 (O_1966,N_29529,N_29713);
nand UO_1967 (O_1967,N_29762,N_29602);
xnor UO_1968 (O_1968,N_29916,N_29449);
and UO_1969 (O_1969,N_29670,N_29779);
or UO_1970 (O_1970,N_29528,N_29829);
and UO_1971 (O_1971,N_29787,N_29477);
and UO_1972 (O_1972,N_29622,N_29924);
nor UO_1973 (O_1973,N_29793,N_29741);
and UO_1974 (O_1974,N_29932,N_29607);
xor UO_1975 (O_1975,N_29493,N_29633);
and UO_1976 (O_1976,N_29447,N_29466);
nand UO_1977 (O_1977,N_29763,N_29950);
nor UO_1978 (O_1978,N_29538,N_29522);
xor UO_1979 (O_1979,N_29929,N_29529);
xnor UO_1980 (O_1980,N_29830,N_29434);
nand UO_1981 (O_1981,N_29632,N_29400);
and UO_1982 (O_1982,N_29528,N_29418);
and UO_1983 (O_1983,N_29522,N_29509);
or UO_1984 (O_1984,N_29817,N_29900);
nand UO_1985 (O_1985,N_29830,N_29713);
and UO_1986 (O_1986,N_29811,N_29454);
and UO_1987 (O_1987,N_29857,N_29678);
or UO_1988 (O_1988,N_29566,N_29680);
nor UO_1989 (O_1989,N_29902,N_29580);
or UO_1990 (O_1990,N_29705,N_29523);
and UO_1991 (O_1991,N_29471,N_29418);
nor UO_1992 (O_1992,N_29732,N_29699);
and UO_1993 (O_1993,N_29431,N_29501);
nand UO_1994 (O_1994,N_29562,N_29489);
xor UO_1995 (O_1995,N_29744,N_29661);
nand UO_1996 (O_1996,N_29822,N_29713);
and UO_1997 (O_1997,N_29510,N_29851);
xor UO_1998 (O_1998,N_29605,N_29711);
or UO_1999 (O_1999,N_29792,N_29527);
xnor UO_2000 (O_2000,N_29417,N_29851);
nor UO_2001 (O_2001,N_29936,N_29753);
and UO_2002 (O_2002,N_29938,N_29438);
nor UO_2003 (O_2003,N_29680,N_29569);
xor UO_2004 (O_2004,N_29485,N_29966);
xor UO_2005 (O_2005,N_29624,N_29989);
nor UO_2006 (O_2006,N_29741,N_29585);
xnor UO_2007 (O_2007,N_29628,N_29438);
or UO_2008 (O_2008,N_29895,N_29516);
xor UO_2009 (O_2009,N_29423,N_29894);
or UO_2010 (O_2010,N_29767,N_29883);
and UO_2011 (O_2011,N_29837,N_29414);
nor UO_2012 (O_2012,N_29857,N_29611);
and UO_2013 (O_2013,N_29619,N_29477);
and UO_2014 (O_2014,N_29509,N_29855);
nand UO_2015 (O_2015,N_29641,N_29924);
xor UO_2016 (O_2016,N_29409,N_29540);
nor UO_2017 (O_2017,N_29905,N_29708);
or UO_2018 (O_2018,N_29665,N_29517);
or UO_2019 (O_2019,N_29891,N_29810);
or UO_2020 (O_2020,N_29545,N_29426);
xor UO_2021 (O_2021,N_29609,N_29751);
or UO_2022 (O_2022,N_29432,N_29874);
nor UO_2023 (O_2023,N_29729,N_29963);
nand UO_2024 (O_2024,N_29554,N_29520);
nand UO_2025 (O_2025,N_29651,N_29536);
or UO_2026 (O_2026,N_29736,N_29898);
or UO_2027 (O_2027,N_29504,N_29510);
nand UO_2028 (O_2028,N_29513,N_29988);
nor UO_2029 (O_2029,N_29932,N_29562);
nand UO_2030 (O_2030,N_29994,N_29800);
nor UO_2031 (O_2031,N_29813,N_29400);
xnor UO_2032 (O_2032,N_29724,N_29960);
and UO_2033 (O_2033,N_29894,N_29616);
nand UO_2034 (O_2034,N_29548,N_29927);
and UO_2035 (O_2035,N_29621,N_29986);
and UO_2036 (O_2036,N_29473,N_29895);
nor UO_2037 (O_2037,N_29725,N_29401);
nor UO_2038 (O_2038,N_29491,N_29509);
xor UO_2039 (O_2039,N_29882,N_29723);
xnor UO_2040 (O_2040,N_29663,N_29675);
and UO_2041 (O_2041,N_29676,N_29729);
xor UO_2042 (O_2042,N_29684,N_29771);
nor UO_2043 (O_2043,N_29480,N_29656);
xor UO_2044 (O_2044,N_29622,N_29841);
and UO_2045 (O_2045,N_29804,N_29885);
nor UO_2046 (O_2046,N_29583,N_29816);
nor UO_2047 (O_2047,N_29988,N_29817);
xor UO_2048 (O_2048,N_29605,N_29819);
and UO_2049 (O_2049,N_29954,N_29882);
nand UO_2050 (O_2050,N_29414,N_29881);
and UO_2051 (O_2051,N_29898,N_29971);
nor UO_2052 (O_2052,N_29744,N_29747);
nor UO_2053 (O_2053,N_29766,N_29962);
nor UO_2054 (O_2054,N_29734,N_29990);
nand UO_2055 (O_2055,N_29483,N_29980);
xor UO_2056 (O_2056,N_29645,N_29792);
xnor UO_2057 (O_2057,N_29765,N_29646);
nand UO_2058 (O_2058,N_29469,N_29722);
xnor UO_2059 (O_2059,N_29945,N_29737);
nor UO_2060 (O_2060,N_29618,N_29573);
nor UO_2061 (O_2061,N_29939,N_29832);
nand UO_2062 (O_2062,N_29768,N_29470);
and UO_2063 (O_2063,N_29730,N_29667);
nor UO_2064 (O_2064,N_29947,N_29675);
nand UO_2065 (O_2065,N_29842,N_29441);
nand UO_2066 (O_2066,N_29761,N_29833);
nor UO_2067 (O_2067,N_29504,N_29463);
nand UO_2068 (O_2068,N_29410,N_29742);
and UO_2069 (O_2069,N_29786,N_29545);
xor UO_2070 (O_2070,N_29977,N_29699);
and UO_2071 (O_2071,N_29918,N_29801);
and UO_2072 (O_2072,N_29972,N_29480);
xor UO_2073 (O_2073,N_29990,N_29861);
and UO_2074 (O_2074,N_29538,N_29619);
nor UO_2075 (O_2075,N_29892,N_29452);
xor UO_2076 (O_2076,N_29605,N_29808);
nor UO_2077 (O_2077,N_29701,N_29901);
or UO_2078 (O_2078,N_29852,N_29526);
or UO_2079 (O_2079,N_29506,N_29442);
nand UO_2080 (O_2080,N_29714,N_29566);
nor UO_2081 (O_2081,N_29524,N_29901);
nand UO_2082 (O_2082,N_29568,N_29709);
nor UO_2083 (O_2083,N_29802,N_29858);
nor UO_2084 (O_2084,N_29818,N_29755);
xor UO_2085 (O_2085,N_29631,N_29619);
and UO_2086 (O_2086,N_29806,N_29608);
nor UO_2087 (O_2087,N_29881,N_29439);
xor UO_2088 (O_2088,N_29627,N_29630);
xor UO_2089 (O_2089,N_29884,N_29845);
xor UO_2090 (O_2090,N_29991,N_29875);
xnor UO_2091 (O_2091,N_29543,N_29820);
nand UO_2092 (O_2092,N_29992,N_29916);
xor UO_2093 (O_2093,N_29517,N_29642);
or UO_2094 (O_2094,N_29714,N_29465);
nor UO_2095 (O_2095,N_29448,N_29445);
or UO_2096 (O_2096,N_29729,N_29822);
xnor UO_2097 (O_2097,N_29771,N_29981);
or UO_2098 (O_2098,N_29651,N_29441);
xor UO_2099 (O_2099,N_29937,N_29885);
nand UO_2100 (O_2100,N_29922,N_29732);
and UO_2101 (O_2101,N_29595,N_29981);
or UO_2102 (O_2102,N_29986,N_29794);
xnor UO_2103 (O_2103,N_29848,N_29881);
or UO_2104 (O_2104,N_29865,N_29737);
xor UO_2105 (O_2105,N_29673,N_29848);
nor UO_2106 (O_2106,N_29899,N_29437);
and UO_2107 (O_2107,N_29876,N_29532);
nor UO_2108 (O_2108,N_29919,N_29583);
nand UO_2109 (O_2109,N_29472,N_29990);
or UO_2110 (O_2110,N_29904,N_29936);
xnor UO_2111 (O_2111,N_29876,N_29678);
or UO_2112 (O_2112,N_29720,N_29597);
and UO_2113 (O_2113,N_29607,N_29707);
nor UO_2114 (O_2114,N_29474,N_29836);
or UO_2115 (O_2115,N_29998,N_29534);
and UO_2116 (O_2116,N_29458,N_29650);
and UO_2117 (O_2117,N_29465,N_29504);
nor UO_2118 (O_2118,N_29814,N_29495);
xnor UO_2119 (O_2119,N_29810,N_29581);
or UO_2120 (O_2120,N_29779,N_29971);
xnor UO_2121 (O_2121,N_29764,N_29786);
and UO_2122 (O_2122,N_29613,N_29821);
nand UO_2123 (O_2123,N_29883,N_29534);
xor UO_2124 (O_2124,N_29887,N_29535);
or UO_2125 (O_2125,N_29503,N_29451);
xor UO_2126 (O_2126,N_29761,N_29961);
xor UO_2127 (O_2127,N_29631,N_29539);
nor UO_2128 (O_2128,N_29515,N_29878);
and UO_2129 (O_2129,N_29548,N_29933);
and UO_2130 (O_2130,N_29593,N_29994);
or UO_2131 (O_2131,N_29448,N_29571);
xnor UO_2132 (O_2132,N_29599,N_29609);
and UO_2133 (O_2133,N_29496,N_29400);
and UO_2134 (O_2134,N_29880,N_29427);
or UO_2135 (O_2135,N_29955,N_29520);
and UO_2136 (O_2136,N_29856,N_29754);
or UO_2137 (O_2137,N_29981,N_29870);
nor UO_2138 (O_2138,N_29528,N_29628);
nor UO_2139 (O_2139,N_29547,N_29980);
xor UO_2140 (O_2140,N_29685,N_29416);
nor UO_2141 (O_2141,N_29494,N_29406);
and UO_2142 (O_2142,N_29734,N_29429);
and UO_2143 (O_2143,N_29447,N_29684);
and UO_2144 (O_2144,N_29599,N_29455);
nor UO_2145 (O_2145,N_29875,N_29429);
and UO_2146 (O_2146,N_29619,N_29835);
xor UO_2147 (O_2147,N_29563,N_29806);
nand UO_2148 (O_2148,N_29829,N_29466);
nor UO_2149 (O_2149,N_29857,N_29832);
and UO_2150 (O_2150,N_29872,N_29875);
xnor UO_2151 (O_2151,N_29776,N_29634);
or UO_2152 (O_2152,N_29841,N_29971);
and UO_2153 (O_2153,N_29722,N_29854);
xor UO_2154 (O_2154,N_29681,N_29531);
nor UO_2155 (O_2155,N_29946,N_29716);
nand UO_2156 (O_2156,N_29832,N_29682);
nor UO_2157 (O_2157,N_29985,N_29521);
xor UO_2158 (O_2158,N_29581,N_29977);
and UO_2159 (O_2159,N_29413,N_29467);
nor UO_2160 (O_2160,N_29839,N_29463);
nand UO_2161 (O_2161,N_29428,N_29924);
nor UO_2162 (O_2162,N_29845,N_29704);
xor UO_2163 (O_2163,N_29998,N_29586);
and UO_2164 (O_2164,N_29957,N_29948);
nand UO_2165 (O_2165,N_29801,N_29945);
xor UO_2166 (O_2166,N_29904,N_29886);
nor UO_2167 (O_2167,N_29886,N_29863);
and UO_2168 (O_2168,N_29949,N_29931);
and UO_2169 (O_2169,N_29460,N_29513);
nor UO_2170 (O_2170,N_29711,N_29500);
and UO_2171 (O_2171,N_29977,N_29897);
nand UO_2172 (O_2172,N_29754,N_29589);
nor UO_2173 (O_2173,N_29662,N_29907);
xor UO_2174 (O_2174,N_29521,N_29582);
xor UO_2175 (O_2175,N_29716,N_29605);
nand UO_2176 (O_2176,N_29971,N_29908);
nor UO_2177 (O_2177,N_29988,N_29667);
nand UO_2178 (O_2178,N_29783,N_29715);
xnor UO_2179 (O_2179,N_29714,N_29521);
nor UO_2180 (O_2180,N_29478,N_29946);
xnor UO_2181 (O_2181,N_29942,N_29846);
nand UO_2182 (O_2182,N_29752,N_29704);
xor UO_2183 (O_2183,N_29953,N_29585);
or UO_2184 (O_2184,N_29956,N_29509);
and UO_2185 (O_2185,N_29502,N_29594);
nand UO_2186 (O_2186,N_29840,N_29820);
or UO_2187 (O_2187,N_29518,N_29597);
nor UO_2188 (O_2188,N_29597,N_29442);
xor UO_2189 (O_2189,N_29838,N_29817);
xor UO_2190 (O_2190,N_29474,N_29615);
nand UO_2191 (O_2191,N_29461,N_29866);
and UO_2192 (O_2192,N_29733,N_29981);
xor UO_2193 (O_2193,N_29935,N_29701);
nand UO_2194 (O_2194,N_29404,N_29693);
or UO_2195 (O_2195,N_29867,N_29700);
nor UO_2196 (O_2196,N_29560,N_29435);
nor UO_2197 (O_2197,N_29677,N_29915);
xor UO_2198 (O_2198,N_29542,N_29930);
or UO_2199 (O_2199,N_29968,N_29661);
nand UO_2200 (O_2200,N_29727,N_29475);
xor UO_2201 (O_2201,N_29966,N_29768);
nand UO_2202 (O_2202,N_29609,N_29542);
xor UO_2203 (O_2203,N_29786,N_29962);
xnor UO_2204 (O_2204,N_29474,N_29914);
or UO_2205 (O_2205,N_29577,N_29456);
xnor UO_2206 (O_2206,N_29798,N_29558);
nor UO_2207 (O_2207,N_29516,N_29581);
nor UO_2208 (O_2208,N_29533,N_29846);
nor UO_2209 (O_2209,N_29711,N_29484);
or UO_2210 (O_2210,N_29442,N_29878);
nand UO_2211 (O_2211,N_29876,N_29960);
xor UO_2212 (O_2212,N_29607,N_29532);
and UO_2213 (O_2213,N_29706,N_29972);
nand UO_2214 (O_2214,N_29574,N_29726);
or UO_2215 (O_2215,N_29844,N_29807);
and UO_2216 (O_2216,N_29805,N_29602);
and UO_2217 (O_2217,N_29960,N_29638);
and UO_2218 (O_2218,N_29611,N_29883);
nor UO_2219 (O_2219,N_29864,N_29802);
xor UO_2220 (O_2220,N_29421,N_29687);
xnor UO_2221 (O_2221,N_29433,N_29408);
nand UO_2222 (O_2222,N_29727,N_29950);
and UO_2223 (O_2223,N_29911,N_29550);
xor UO_2224 (O_2224,N_29914,N_29549);
xnor UO_2225 (O_2225,N_29819,N_29511);
or UO_2226 (O_2226,N_29812,N_29791);
nor UO_2227 (O_2227,N_29522,N_29427);
nor UO_2228 (O_2228,N_29991,N_29633);
xor UO_2229 (O_2229,N_29470,N_29734);
and UO_2230 (O_2230,N_29458,N_29465);
xnor UO_2231 (O_2231,N_29829,N_29729);
nor UO_2232 (O_2232,N_29617,N_29608);
nor UO_2233 (O_2233,N_29709,N_29560);
nand UO_2234 (O_2234,N_29861,N_29586);
nand UO_2235 (O_2235,N_29707,N_29943);
and UO_2236 (O_2236,N_29603,N_29593);
xnor UO_2237 (O_2237,N_29778,N_29582);
and UO_2238 (O_2238,N_29407,N_29781);
nand UO_2239 (O_2239,N_29420,N_29752);
nand UO_2240 (O_2240,N_29672,N_29593);
xor UO_2241 (O_2241,N_29632,N_29972);
nand UO_2242 (O_2242,N_29690,N_29794);
xor UO_2243 (O_2243,N_29776,N_29451);
nand UO_2244 (O_2244,N_29681,N_29454);
or UO_2245 (O_2245,N_29851,N_29569);
xnor UO_2246 (O_2246,N_29879,N_29782);
nand UO_2247 (O_2247,N_29637,N_29994);
or UO_2248 (O_2248,N_29741,N_29554);
xor UO_2249 (O_2249,N_29460,N_29911);
nor UO_2250 (O_2250,N_29678,N_29407);
and UO_2251 (O_2251,N_29929,N_29461);
xnor UO_2252 (O_2252,N_29797,N_29409);
or UO_2253 (O_2253,N_29957,N_29903);
and UO_2254 (O_2254,N_29792,N_29770);
and UO_2255 (O_2255,N_29525,N_29929);
xor UO_2256 (O_2256,N_29619,N_29857);
nor UO_2257 (O_2257,N_29447,N_29589);
and UO_2258 (O_2258,N_29511,N_29487);
nand UO_2259 (O_2259,N_29635,N_29468);
nor UO_2260 (O_2260,N_29425,N_29743);
nor UO_2261 (O_2261,N_29407,N_29461);
or UO_2262 (O_2262,N_29751,N_29938);
nand UO_2263 (O_2263,N_29709,N_29669);
xor UO_2264 (O_2264,N_29500,N_29961);
nor UO_2265 (O_2265,N_29960,N_29481);
or UO_2266 (O_2266,N_29945,N_29474);
and UO_2267 (O_2267,N_29829,N_29849);
xor UO_2268 (O_2268,N_29463,N_29996);
nand UO_2269 (O_2269,N_29894,N_29583);
nor UO_2270 (O_2270,N_29610,N_29497);
nor UO_2271 (O_2271,N_29613,N_29673);
nand UO_2272 (O_2272,N_29437,N_29938);
nand UO_2273 (O_2273,N_29720,N_29501);
nor UO_2274 (O_2274,N_29618,N_29931);
nor UO_2275 (O_2275,N_29861,N_29639);
nand UO_2276 (O_2276,N_29628,N_29705);
nand UO_2277 (O_2277,N_29839,N_29690);
nor UO_2278 (O_2278,N_29782,N_29795);
nand UO_2279 (O_2279,N_29943,N_29437);
and UO_2280 (O_2280,N_29689,N_29725);
nor UO_2281 (O_2281,N_29875,N_29541);
and UO_2282 (O_2282,N_29933,N_29421);
or UO_2283 (O_2283,N_29780,N_29422);
nor UO_2284 (O_2284,N_29855,N_29795);
or UO_2285 (O_2285,N_29504,N_29989);
or UO_2286 (O_2286,N_29873,N_29619);
xor UO_2287 (O_2287,N_29677,N_29529);
nand UO_2288 (O_2288,N_29846,N_29492);
nand UO_2289 (O_2289,N_29764,N_29464);
or UO_2290 (O_2290,N_29871,N_29630);
and UO_2291 (O_2291,N_29781,N_29623);
nor UO_2292 (O_2292,N_29667,N_29421);
xnor UO_2293 (O_2293,N_29846,N_29574);
xnor UO_2294 (O_2294,N_29638,N_29485);
nor UO_2295 (O_2295,N_29711,N_29825);
or UO_2296 (O_2296,N_29487,N_29439);
nor UO_2297 (O_2297,N_29678,N_29741);
and UO_2298 (O_2298,N_29792,N_29844);
and UO_2299 (O_2299,N_29795,N_29577);
nand UO_2300 (O_2300,N_29707,N_29767);
or UO_2301 (O_2301,N_29655,N_29680);
nor UO_2302 (O_2302,N_29897,N_29891);
xnor UO_2303 (O_2303,N_29939,N_29597);
nand UO_2304 (O_2304,N_29482,N_29672);
or UO_2305 (O_2305,N_29653,N_29860);
xnor UO_2306 (O_2306,N_29708,N_29595);
nor UO_2307 (O_2307,N_29952,N_29472);
nand UO_2308 (O_2308,N_29543,N_29561);
nor UO_2309 (O_2309,N_29585,N_29737);
nand UO_2310 (O_2310,N_29643,N_29559);
nor UO_2311 (O_2311,N_29755,N_29465);
nand UO_2312 (O_2312,N_29532,N_29449);
or UO_2313 (O_2313,N_29403,N_29597);
and UO_2314 (O_2314,N_29482,N_29530);
or UO_2315 (O_2315,N_29510,N_29814);
nor UO_2316 (O_2316,N_29486,N_29416);
or UO_2317 (O_2317,N_29963,N_29756);
nor UO_2318 (O_2318,N_29994,N_29832);
nand UO_2319 (O_2319,N_29999,N_29454);
nor UO_2320 (O_2320,N_29957,N_29852);
nor UO_2321 (O_2321,N_29655,N_29717);
nor UO_2322 (O_2322,N_29849,N_29800);
and UO_2323 (O_2323,N_29479,N_29841);
xor UO_2324 (O_2324,N_29541,N_29557);
or UO_2325 (O_2325,N_29707,N_29736);
nor UO_2326 (O_2326,N_29874,N_29947);
or UO_2327 (O_2327,N_29427,N_29950);
nand UO_2328 (O_2328,N_29996,N_29722);
nor UO_2329 (O_2329,N_29966,N_29489);
or UO_2330 (O_2330,N_29941,N_29711);
and UO_2331 (O_2331,N_29974,N_29520);
and UO_2332 (O_2332,N_29750,N_29614);
nand UO_2333 (O_2333,N_29498,N_29442);
and UO_2334 (O_2334,N_29720,N_29600);
and UO_2335 (O_2335,N_29796,N_29804);
xor UO_2336 (O_2336,N_29900,N_29518);
nor UO_2337 (O_2337,N_29586,N_29657);
and UO_2338 (O_2338,N_29995,N_29911);
and UO_2339 (O_2339,N_29880,N_29495);
and UO_2340 (O_2340,N_29835,N_29882);
or UO_2341 (O_2341,N_29749,N_29568);
and UO_2342 (O_2342,N_29965,N_29801);
and UO_2343 (O_2343,N_29982,N_29958);
xor UO_2344 (O_2344,N_29478,N_29598);
xor UO_2345 (O_2345,N_29663,N_29914);
or UO_2346 (O_2346,N_29507,N_29557);
xor UO_2347 (O_2347,N_29594,N_29826);
or UO_2348 (O_2348,N_29473,N_29997);
and UO_2349 (O_2349,N_29429,N_29946);
nor UO_2350 (O_2350,N_29907,N_29655);
and UO_2351 (O_2351,N_29479,N_29578);
and UO_2352 (O_2352,N_29882,N_29708);
or UO_2353 (O_2353,N_29711,N_29861);
and UO_2354 (O_2354,N_29823,N_29558);
xor UO_2355 (O_2355,N_29655,N_29637);
xnor UO_2356 (O_2356,N_29992,N_29779);
and UO_2357 (O_2357,N_29468,N_29602);
nand UO_2358 (O_2358,N_29812,N_29947);
nor UO_2359 (O_2359,N_29651,N_29799);
nand UO_2360 (O_2360,N_29664,N_29427);
nor UO_2361 (O_2361,N_29557,N_29648);
nand UO_2362 (O_2362,N_29545,N_29632);
nor UO_2363 (O_2363,N_29823,N_29772);
or UO_2364 (O_2364,N_29854,N_29526);
nand UO_2365 (O_2365,N_29981,N_29607);
nand UO_2366 (O_2366,N_29924,N_29545);
or UO_2367 (O_2367,N_29623,N_29838);
and UO_2368 (O_2368,N_29746,N_29529);
or UO_2369 (O_2369,N_29983,N_29446);
nor UO_2370 (O_2370,N_29455,N_29913);
xnor UO_2371 (O_2371,N_29996,N_29672);
nand UO_2372 (O_2372,N_29819,N_29513);
nand UO_2373 (O_2373,N_29965,N_29815);
nand UO_2374 (O_2374,N_29481,N_29561);
nand UO_2375 (O_2375,N_29772,N_29705);
and UO_2376 (O_2376,N_29588,N_29528);
nor UO_2377 (O_2377,N_29979,N_29791);
nor UO_2378 (O_2378,N_29597,N_29686);
and UO_2379 (O_2379,N_29751,N_29437);
and UO_2380 (O_2380,N_29956,N_29975);
nand UO_2381 (O_2381,N_29489,N_29788);
xnor UO_2382 (O_2382,N_29888,N_29847);
nand UO_2383 (O_2383,N_29719,N_29954);
nand UO_2384 (O_2384,N_29950,N_29769);
nor UO_2385 (O_2385,N_29561,N_29875);
nor UO_2386 (O_2386,N_29867,N_29596);
or UO_2387 (O_2387,N_29725,N_29895);
nor UO_2388 (O_2388,N_29843,N_29944);
xor UO_2389 (O_2389,N_29852,N_29565);
nor UO_2390 (O_2390,N_29916,N_29532);
or UO_2391 (O_2391,N_29701,N_29642);
and UO_2392 (O_2392,N_29473,N_29725);
xor UO_2393 (O_2393,N_29405,N_29604);
nand UO_2394 (O_2394,N_29726,N_29556);
and UO_2395 (O_2395,N_29817,N_29753);
nand UO_2396 (O_2396,N_29544,N_29867);
nor UO_2397 (O_2397,N_29667,N_29613);
xor UO_2398 (O_2398,N_29679,N_29784);
nand UO_2399 (O_2399,N_29947,N_29999);
and UO_2400 (O_2400,N_29835,N_29641);
or UO_2401 (O_2401,N_29686,N_29584);
nand UO_2402 (O_2402,N_29601,N_29469);
or UO_2403 (O_2403,N_29538,N_29921);
nand UO_2404 (O_2404,N_29947,N_29862);
nand UO_2405 (O_2405,N_29785,N_29799);
and UO_2406 (O_2406,N_29413,N_29439);
and UO_2407 (O_2407,N_29577,N_29581);
or UO_2408 (O_2408,N_29453,N_29636);
or UO_2409 (O_2409,N_29485,N_29944);
nand UO_2410 (O_2410,N_29865,N_29811);
nor UO_2411 (O_2411,N_29914,N_29898);
and UO_2412 (O_2412,N_29904,N_29733);
or UO_2413 (O_2413,N_29812,N_29681);
and UO_2414 (O_2414,N_29898,N_29516);
xnor UO_2415 (O_2415,N_29417,N_29844);
or UO_2416 (O_2416,N_29845,N_29945);
or UO_2417 (O_2417,N_29532,N_29503);
and UO_2418 (O_2418,N_29790,N_29934);
nor UO_2419 (O_2419,N_29511,N_29793);
nor UO_2420 (O_2420,N_29861,N_29624);
xnor UO_2421 (O_2421,N_29501,N_29702);
and UO_2422 (O_2422,N_29951,N_29918);
nor UO_2423 (O_2423,N_29943,N_29472);
or UO_2424 (O_2424,N_29896,N_29589);
nand UO_2425 (O_2425,N_29782,N_29822);
xnor UO_2426 (O_2426,N_29751,N_29711);
and UO_2427 (O_2427,N_29762,N_29979);
and UO_2428 (O_2428,N_29656,N_29995);
nand UO_2429 (O_2429,N_29621,N_29449);
and UO_2430 (O_2430,N_29976,N_29455);
nand UO_2431 (O_2431,N_29663,N_29571);
nor UO_2432 (O_2432,N_29442,N_29883);
nor UO_2433 (O_2433,N_29405,N_29455);
nor UO_2434 (O_2434,N_29631,N_29975);
nand UO_2435 (O_2435,N_29924,N_29872);
or UO_2436 (O_2436,N_29604,N_29645);
or UO_2437 (O_2437,N_29926,N_29698);
and UO_2438 (O_2438,N_29698,N_29708);
and UO_2439 (O_2439,N_29929,N_29577);
nor UO_2440 (O_2440,N_29931,N_29540);
or UO_2441 (O_2441,N_29669,N_29911);
nor UO_2442 (O_2442,N_29462,N_29996);
xor UO_2443 (O_2443,N_29563,N_29534);
nor UO_2444 (O_2444,N_29981,N_29562);
or UO_2445 (O_2445,N_29501,N_29416);
nand UO_2446 (O_2446,N_29688,N_29403);
nand UO_2447 (O_2447,N_29937,N_29511);
nor UO_2448 (O_2448,N_29641,N_29581);
xor UO_2449 (O_2449,N_29423,N_29526);
nand UO_2450 (O_2450,N_29648,N_29414);
xnor UO_2451 (O_2451,N_29838,N_29823);
and UO_2452 (O_2452,N_29534,N_29743);
and UO_2453 (O_2453,N_29734,N_29872);
or UO_2454 (O_2454,N_29431,N_29810);
nor UO_2455 (O_2455,N_29540,N_29662);
or UO_2456 (O_2456,N_29737,N_29747);
and UO_2457 (O_2457,N_29605,N_29608);
nor UO_2458 (O_2458,N_29850,N_29802);
or UO_2459 (O_2459,N_29762,N_29569);
or UO_2460 (O_2460,N_29443,N_29775);
nand UO_2461 (O_2461,N_29655,N_29520);
nor UO_2462 (O_2462,N_29976,N_29902);
xor UO_2463 (O_2463,N_29763,N_29952);
nor UO_2464 (O_2464,N_29749,N_29595);
nand UO_2465 (O_2465,N_29534,N_29539);
and UO_2466 (O_2466,N_29420,N_29851);
and UO_2467 (O_2467,N_29520,N_29885);
nand UO_2468 (O_2468,N_29919,N_29975);
nor UO_2469 (O_2469,N_29660,N_29723);
and UO_2470 (O_2470,N_29838,N_29428);
or UO_2471 (O_2471,N_29436,N_29496);
or UO_2472 (O_2472,N_29743,N_29489);
xnor UO_2473 (O_2473,N_29557,N_29532);
nor UO_2474 (O_2474,N_29831,N_29449);
nand UO_2475 (O_2475,N_29423,N_29668);
xnor UO_2476 (O_2476,N_29983,N_29626);
nand UO_2477 (O_2477,N_29579,N_29586);
and UO_2478 (O_2478,N_29542,N_29751);
and UO_2479 (O_2479,N_29472,N_29658);
xnor UO_2480 (O_2480,N_29595,N_29722);
or UO_2481 (O_2481,N_29806,N_29641);
xnor UO_2482 (O_2482,N_29771,N_29927);
and UO_2483 (O_2483,N_29865,N_29471);
nand UO_2484 (O_2484,N_29944,N_29888);
or UO_2485 (O_2485,N_29648,N_29880);
and UO_2486 (O_2486,N_29803,N_29739);
or UO_2487 (O_2487,N_29681,N_29517);
nor UO_2488 (O_2488,N_29740,N_29537);
or UO_2489 (O_2489,N_29605,N_29975);
xor UO_2490 (O_2490,N_29755,N_29994);
nor UO_2491 (O_2491,N_29780,N_29833);
xor UO_2492 (O_2492,N_29635,N_29508);
nand UO_2493 (O_2493,N_29970,N_29786);
and UO_2494 (O_2494,N_29585,N_29499);
nand UO_2495 (O_2495,N_29908,N_29803);
and UO_2496 (O_2496,N_29756,N_29856);
xor UO_2497 (O_2497,N_29855,N_29888);
nand UO_2498 (O_2498,N_29705,N_29910);
xnor UO_2499 (O_2499,N_29983,N_29876);
or UO_2500 (O_2500,N_29536,N_29811);
or UO_2501 (O_2501,N_29730,N_29549);
or UO_2502 (O_2502,N_29489,N_29851);
and UO_2503 (O_2503,N_29431,N_29418);
nor UO_2504 (O_2504,N_29668,N_29580);
or UO_2505 (O_2505,N_29506,N_29798);
nor UO_2506 (O_2506,N_29619,N_29745);
and UO_2507 (O_2507,N_29670,N_29426);
or UO_2508 (O_2508,N_29926,N_29522);
nor UO_2509 (O_2509,N_29739,N_29651);
nor UO_2510 (O_2510,N_29561,N_29605);
nor UO_2511 (O_2511,N_29561,N_29925);
or UO_2512 (O_2512,N_29551,N_29675);
nand UO_2513 (O_2513,N_29844,N_29664);
xor UO_2514 (O_2514,N_29608,N_29648);
nand UO_2515 (O_2515,N_29565,N_29634);
or UO_2516 (O_2516,N_29952,N_29485);
nor UO_2517 (O_2517,N_29579,N_29810);
and UO_2518 (O_2518,N_29572,N_29467);
nand UO_2519 (O_2519,N_29460,N_29926);
nand UO_2520 (O_2520,N_29836,N_29421);
nor UO_2521 (O_2521,N_29780,N_29639);
nand UO_2522 (O_2522,N_29600,N_29692);
nor UO_2523 (O_2523,N_29820,N_29786);
nor UO_2524 (O_2524,N_29425,N_29421);
and UO_2525 (O_2525,N_29582,N_29739);
xor UO_2526 (O_2526,N_29795,N_29804);
xnor UO_2527 (O_2527,N_29772,N_29795);
xnor UO_2528 (O_2528,N_29907,N_29790);
nand UO_2529 (O_2529,N_29922,N_29968);
nor UO_2530 (O_2530,N_29933,N_29838);
nor UO_2531 (O_2531,N_29910,N_29845);
nand UO_2532 (O_2532,N_29971,N_29684);
and UO_2533 (O_2533,N_29426,N_29597);
xor UO_2534 (O_2534,N_29869,N_29679);
nand UO_2535 (O_2535,N_29657,N_29830);
or UO_2536 (O_2536,N_29830,N_29403);
nand UO_2537 (O_2537,N_29423,N_29807);
and UO_2538 (O_2538,N_29996,N_29719);
xnor UO_2539 (O_2539,N_29517,N_29613);
xnor UO_2540 (O_2540,N_29621,N_29845);
nand UO_2541 (O_2541,N_29843,N_29976);
nor UO_2542 (O_2542,N_29513,N_29599);
nand UO_2543 (O_2543,N_29612,N_29495);
nand UO_2544 (O_2544,N_29682,N_29441);
and UO_2545 (O_2545,N_29841,N_29682);
nor UO_2546 (O_2546,N_29637,N_29927);
or UO_2547 (O_2547,N_29963,N_29866);
and UO_2548 (O_2548,N_29852,N_29806);
nor UO_2549 (O_2549,N_29836,N_29485);
nand UO_2550 (O_2550,N_29923,N_29869);
and UO_2551 (O_2551,N_29715,N_29797);
or UO_2552 (O_2552,N_29516,N_29687);
nor UO_2553 (O_2553,N_29625,N_29922);
xor UO_2554 (O_2554,N_29627,N_29722);
xnor UO_2555 (O_2555,N_29684,N_29661);
nor UO_2556 (O_2556,N_29882,N_29646);
or UO_2557 (O_2557,N_29404,N_29582);
and UO_2558 (O_2558,N_29766,N_29945);
nor UO_2559 (O_2559,N_29825,N_29483);
xor UO_2560 (O_2560,N_29737,N_29513);
xnor UO_2561 (O_2561,N_29928,N_29465);
xor UO_2562 (O_2562,N_29830,N_29455);
xnor UO_2563 (O_2563,N_29673,N_29678);
nor UO_2564 (O_2564,N_29660,N_29595);
or UO_2565 (O_2565,N_29813,N_29931);
or UO_2566 (O_2566,N_29870,N_29576);
xnor UO_2567 (O_2567,N_29615,N_29668);
and UO_2568 (O_2568,N_29542,N_29727);
nor UO_2569 (O_2569,N_29445,N_29544);
nor UO_2570 (O_2570,N_29891,N_29448);
xnor UO_2571 (O_2571,N_29954,N_29887);
nand UO_2572 (O_2572,N_29738,N_29804);
and UO_2573 (O_2573,N_29618,N_29532);
nor UO_2574 (O_2574,N_29705,N_29752);
nor UO_2575 (O_2575,N_29782,N_29810);
nand UO_2576 (O_2576,N_29945,N_29590);
nand UO_2577 (O_2577,N_29721,N_29420);
and UO_2578 (O_2578,N_29668,N_29690);
or UO_2579 (O_2579,N_29446,N_29665);
nor UO_2580 (O_2580,N_29761,N_29978);
or UO_2581 (O_2581,N_29903,N_29501);
or UO_2582 (O_2582,N_29431,N_29899);
xnor UO_2583 (O_2583,N_29419,N_29870);
or UO_2584 (O_2584,N_29918,N_29534);
and UO_2585 (O_2585,N_29439,N_29482);
or UO_2586 (O_2586,N_29793,N_29838);
nor UO_2587 (O_2587,N_29793,N_29901);
xor UO_2588 (O_2588,N_29698,N_29950);
nand UO_2589 (O_2589,N_29979,N_29753);
or UO_2590 (O_2590,N_29419,N_29995);
or UO_2591 (O_2591,N_29931,N_29998);
nand UO_2592 (O_2592,N_29765,N_29560);
nand UO_2593 (O_2593,N_29668,N_29407);
xnor UO_2594 (O_2594,N_29977,N_29859);
xnor UO_2595 (O_2595,N_29723,N_29990);
xor UO_2596 (O_2596,N_29529,N_29494);
nand UO_2597 (O_2597,N_29749,N_29743);
nand UO_2598 (O_2598,N_29806,N_29935);
and UO_2599 (O_2599,N_29959,N_29830);
nand UO_2600 (O_2600,N_29606,N_29928);
nand UO_2601 (O_2601,N_29568,N_29920);
and UO_2602 (O_2602,N_29574,N_29645);
and UO_2603 (O_2603,N_29735,N_29568);
or UO_2604 (O_2604,N_29556,N_29564);
and UO_2605 (O_2605,N_29833,N_29465);
or UO_2606 (O_2606,N_29890,N_29471);
nor UO_2607 (O_2607,N_29481,N_29511);
and UO_2608 (O_2608,N_29470,N_29428);
or UO_2609 (O_2609,N_29527,N_29902);
or UO_2610 (O_2610,N_29851,N_29461);
nor UO_2611 (O_2611,N_29912,N_29765);
and UO_2612 (O_2612,N_29755,N_29460);
or UO_2613 (O_2613,N_29472,N_29568);
nor UO_2614 (O_2614,N_29457,N_29649);
or UO_2615 (O_2615,N_29411,N_29790);
or UO_2616 (O_2616,N_29635,N_29661);
nand UO_2617 (O_2617,N_29622,N_29420);
nand UO_2618 (O_2618,N_29620,N_29419);
and UO_2619 (O_2619,N_29449,N_29829);
or UO_2620 (O_2620,N_29754,N_29613);
nand UO_2621 (O_2621,N_29458,N_29459);
or UO_2622 (O_2622,N_29917,N_29879);
and UO_2623 (O_2623,N_29924,N_29882);
xnor UO_2624 (O_2624,N_29528,N_29724);
or UO_2625 (O_2625,N_29782,N_29687);
nand UO_2626 (O_2626,N_29757,N_29648);
nor UO_2627 (O_2627,N_29512,N_29435);
and UO_2628 (O_2628,N_29704,N_29701);
nor UO_2629 (O_2629,N_29638,N_29867);
and UO_2630 (O_2630,N_29910,N_29767);
xor UO_2631 (O_2631,N_29515,N_29473);
or UO_2632 (O_2632,N_29480,N_29834);
or UO_2633 (O_2633,N_29468,N_29882);
xor UO_2634 (O_2634,N_29632,N_29842);
or UO_2635 (O_2635,N_29517,N_29798);
xor UO_2636 (O_2636,N_29824,N_29991);
xor UO_2637 (O_2637,N_29964,N_29764);
or UO_2638 (O_2638,N_29492,N_29704);
or UO_2639 (O_2639,N_29802,N_29859);
and UO_2640 (O_2640,N_29778,N_29769);
and UO_2641 (O_2641,N_29712,N_29679);
nor UO_2642 (O_2642,N_29567,N_29853);
and UO_2643 (O_2643,N_29738,N_29972);
and UO_2644 (O_2644,N_29603,N_29831);
and UO_2645 (O_2645,N_29576,N_29541);
nand UO_2646 (O_2646,N_29937,N_29793);
nand UO_2647 (O_2647,N_29750,N_29981);
nand UO_2648 (O_2648,N_29531,N_29893);
and UO_2649 (O_2649,N_29598,N_29732);
nand UO_2650 (O_2650,N_29597,N_29947);
or UO_2651 (O_2651,N_29593,N_29512);
xnor UO_2652 (O_2652,N_29751,N_29495);
or UO_2653 (O_2653,N_29905,N_29885);
or UO_2654 (O_2654,N_29426,N_29441);
or UO_2655 (O_2655,N_29869,N_29436);
nor UO_2656 (O_2656,N_29720,N_29788);
nand UO_2657 (O_2657,N_29725,N_29882);
xnor UO_2658 (O_2658,N_29588,N_29729);
or UO_2659 (O_2659,N_29534,N_29550);
xor UO_2660 (O_2660,N_29832,N_29840);
or UO_2661 (O_2661,N_29531,N_29430);
nor UO_2662 (O_2662,N_29758,N_29423);
and UO_2663 (O_2663,N_29587,N_29719);
nand UO_2664 (O_2664,N_29854,N_29646);
nand UO_2665 (O_2665,N_29427,N_29930);
nor UO_2666 (O_2666,N_29890,N_29671);
xnor UO_2667 (O_2667,N_29701,N_29903);
nor UO_2668 (O_2668,N_29593,N_29934);
nor UO_2669 (O_2669,N_29425,N_29790);
nor UO_2670 (O_2670,N_29682,N_29987);
xnor UO_2671 (O_2671,N_29660,N_29954);
or UO_2672 (O_2672,N_29792,N_29687);
or UO_2673 (O_2673,N_29621,N_29853);
nand UO_2674 (O_2674,N_29729,N_29923);
and UO_2675 (O_2675,N_29406,N_29577);
and UO_2676 (O_2676,N_29418,N_29772);
nor UO_2677 (O_2677,N_29863,N_29981);
and UO_2678 (O_2678,N_29583,N_29848);
nand UO_2679 (O_2679,N_29642,N_29481);
and UO_2680 (O_2680,N_29819,N_29688);
or UO_2681 (O_2681,N_29440,N_29530);
and UO_2682 (O_2682,N_29438,N_29875);
nand UO_2683 (O_2683,N_29762,N_29827);
nand UO_2684 (O_2684,N_29831,N_29516);
nor UO_2685 (O_2685,N_29859,N_29431);
nor UO_2686 (O_2686,N_29743,N_29683);
nor UO_2687 (O_2687,N_29546,N_29714);
and UO_2688 (O_2688,N_29859,N_29543);
nor UO_2689 (O_2689,N_29883,N_29423);
or UO_2690 (O_2690,N_29443,N_29783);
or UO_2691 (O_2691,N_29817,N_29869);
xnor UO_2692 (O_2692,N_29426,N_29882);
or UO_2693 (O_2693,N_29421,N_29725);
nor UO_2694 (O_2694,N_29643,N_29748);
and UO_2695 (O_2695,N_29792,N_29439);
nand UO_2696 (O_2696,N_29572,N_29550);
and UO_2697 (O_2697,N_29601,N_29933);
and UO_2698 (O_2698,N_29892,N_29905);
xor UO_2699 (O_2699,N_29626,N_29547);
xor UO_2700 (O_2700,N_29685,N_29846);
nor UO_2701 (O_2701,N_29545,N_29880);
and UO_2702 (O_2702,N_29447,N_29658);
or UO_2703 (O_2703,N_29870,N_29917);
or UO_2704 (O_2704,N_29659,N_29420);
nor UO_2705 (O_2705,N_29544,N_29839);
and UO_2706 (O_2706,N_29503,N_29712);
nand UO_2707 (O_2707,N_29593,N_29699);
and UO_2708 (O_2708,N_29855,N_29582);
nor UO_2709 (O_2709,N_29483,N_29524);
nand UO_2710 (O_2710,N_29929,N_29801);
and UO_2711 (O_2711,N_29436,N_29954);
nand UO_2712 (O_2712,N_29468,N_29984);
and UO_2713 (O_2713,N_29839,N_29978);
xnor UO_2714 (O_2714,N_29550,N_29834);
nor UO_2715 (O_2715,N_29829,N_29517);
nor UO_2716 (O_2716,N_29798,N_29766);
xor UO_2717 (O_2717,N_29924,N_29977);
or UO_2718 (O_2718,N_29493,N_29458);
xor UO_2719 (O_2719,N_29917,N_29719);
and UO_2720 (O_2720,N_29604,N_29617);
nor UO_2721 (O_2721,N_29833,N_29694);
xor UO_2722 (O_2722,N_29790,N_29605);
and UO_2723 (O_2723,N_29755,N_29829);
or UO_2724 (O_2724,N_29825,N_29533);
xnor UO_2725 (O_2725,N_29556,N_29787);
and UO_2726 (O_2726,N_29861,N_29484);
nand UO_2727 (O_2727,N_29539,N_29486);
and UO_2728 (O_2728,N_29645,N_29684);
nand UO_2729 (O_2729,N_29427,N_29792);
xor UO_2730 (O_2730,N_29428,N_29729);
nand UO_2731 (O_2731,N_29607,N_29412);
xor UO_2732 (O_2732,N_29976,N_29974);
nor UO_2733 (O_2733,N_29839,N_29720);
xnor UO_2734 (O_2734,N_29706,N_29860);
nand UO_2735 (O_2735,N_29791,N_29892);
nor UO_2736 (O_2736,N_29724,N_29682);
nand UO_2737 (O_2737,N_29741,N_29589);
and UO_2738 (O_2738,N_29967,N_29864);
nor UO_2739 (O_2739,N_29986,N_29694);
or UO_2740 (O_2740,N_29504,N_29646);
and UO_2741 (O_2741,N_29464,N_29691);
xor UO_2742 (O_2742,N_29793,N_29651);
and UO_2743 (O_2743,N_29459,N_29413);
nor UO_2744 (O_2744,N_29726,N_29620);
xor UO_2745 (O_2745,N_29890,N_29413);
nand UO_2746 (O_2746,N_29922,N_29527);
and UO_2747 (O_2747,N_29844,N_29943);
or UO_2748 (O_2748,N_29650,N_29448);
xnor UO_2749 (O_2749,N_29875,N_29618);
or UO_2750 (O_2750,N_29850,N_29970);
or UO_2751 (O_2751,N_29959,N_29951);
nand UO_2752 (O_2752,N_29894,N_29876);
and UO_2753 (O_2753,N_29674,N_29992);
or UO_2754 (O_2754,N_29732,N_29899);
nor UO_2755 (O_2755,N_29601,N_29509);
nor UO_2756 (O_2756,N_29685,N_29903);
xor UO_2757 (O_2757,N_29836,N_29995);
nor UO_2758 (O_2758,N_29982,N_29488);
or UO_2759 (O_2759,N_29989,N_29506);
nand UO_2760 (O_2760,N_29732,N_29600);
or UO_2761 (O_2761,N_29467,N_29503);
nor UO_2762 (O_2762,N_29462,N_29561);
and UO_2763 (O_2763,N_29938,N_29651);
and UO_2764 (O_2764,N_29453,N_29913);
nand UO_2765 (O_2765,N_29652,N_29440);
nand UO_2766 (O_2766,N_29757,N_29693);
or UO_2767 (O_2767,N_29787,N_29895);
or UO_2768 (O_2768,N_29523,N_29852);
and UO_2769 (O_2769,N_29431,N_29990);
nand UO_2770 (O_2770,N_29666,N_29435);
xor UO_2771 (O_2771,N_29750,N_29557);
nor UO_2772 (O_2772,N_29672,N_29852);
and UO_2773 (O_2773,N_29609,N_29922);
nor UO_2774 (O_2774,N_29487,N_29720);
xor UO_2775 (O_2775,N_29461,N_29573);
or UO_2776 (O_2776,N_29442,N_29519);
nand UO_2777 (O_2777,N_29504,N_29477);
xor UO_2778 (O_2778,N_29984,N_29803);
and UO_2779 (O_2779,N_29889,N_29767);
nand UO_2780 (O_2780,N_29724,N_29537);
xnor UO_2781 (O_2781,N_29863,N_29609);
nor UO_2782 (O_2782,N_29875,N_29742);
or UO_2783 (O_2783,N_29626,N_29786);
xor UO_2784 (O_2784,N_29664,N_29785);
xor UO_2785 (O_2785,N_29878,N_29557);
nand UO_2786 (O_2786,N_29473,N_29926);
xnor UO_2787 (O_2787,N_29732,N_29913);
xor UO_2788 (O_2788,N_29663,N_29648);
xnor UO_2789 (O_2789,N_29802,N_29951);
nor UO_2790 (O_2790,N_29690,N_29903);
nor UO_2791 (O_2791,N_29792,N_29412);
xor UO_2792 (O_2792,N_29736,N_29701);
nand UO_2793 (O_2793,N_29699,N_29972);
or UO_2794 (O_2794,N_29572,N_29500);
and UO_2795 (O_2795,N_29462,N_29581);
nand UO_2796 (O_2796,N_29781,N_29715);
nor UO_2797 (O_2797,N_29857,N_29898);
xor UO_2798 (O_2798,N_29505,N_29961);
nor UO_2799 (O_2799,N_29567,N_29934);
or UO_2800 (O_2800,N_29983,N_29947);
nand UO_2801 (O_2801,N_29936,N_29869);
nand UO_2802 (O_2802,N_29504,N_29542);
and UO_2803 (O_2803,N_29971,N_29967);
or UO_2804 (O_2804,N_29726,N_29866);
nor UO_2805 (O_2805,N_29841,N_29545);
nand UO_2806 (O_2806,N_29483,N_29702);
nand UO_2807 (O_2807,N_29897,N_29585);
or UO_2808 (O_2808,N_29672,N_29414);
and UO_2809 (O_2809,N_29767,N_29447);
nand UO_2810 (O_2810,N_29786,N_29950);
or UO_2811 (O_2811,N_29836,N_29414);
nand UO_2812 (O_2812,N_29962,N_29556);
nor UO_2813 (O_2813,N_29559,N_29409);
nand UO_2814 (O_2814,N_29978,N_29748);
nor UO_2815 (O_2815,N_29440,N_29961);
nand UO_2816 (O_2816,N_29728,N_29906);
nor UO_2817 (O_2817,N_29999,N_29920);
and UO_2818 (O_2818,N_29737,N_29923);
xor UO_2819 (O_2819,N_29966,N_29838);
or UO_2820 (O_2820,N_29526,N_29406);
nor UO_2821 (O_2821,N_29682,N_29472);
or UO_2822 (O_2822,N_29667,N_29866);
nor UO_2823 (O_2823,N_29456,N_29738);
nand UO_2824 (O_2824,N_29790,N_29918);
or UO_2825 (O_2825,N_29839,N_29817);
or UO_2826 (O_2826,N_29816,N_29575);
nand UO_2827 (O_2827,N_29849,N_29793);
xnor UO_2828 (O_2828,N_29665,N_29832);
and UO_2829 (O_2829,N_29921,N_29847);
xnor UO_2830 (O_2830,N_29522,N_29711);
nand UO_2831 (O_2831,N_29811,N_29999);
and UO_2832 (O_2832,N_29925,N_29609);
or UO_2833 (O_2833,N_29832,N_29946);
xor UO_2834 (O_2834,N_29694,N_29977);
and UO_2835 (O_2835,N_29720,N_29558);
xor UO_2836 (O_2836,N_29907,N_29846);
nor UO_2837 (O_2837,N_29754,N_29563);
or UO_2838 (O_2838,N_29940,N_29619);
and UO_2839 (O_2839,N_29646,N_29908);
nor UO_2840 (O_2840,N_29850,N_29687);
or UO_2841 (O_2841,N_29707,N_29741);
and UO_2842 (O_2842,N_29965,N_29751);
nand UO_2843 (O_2843,N_29504,N_29503);
xor UO_2844 (O_2844,N_29462,N_29720);
or UO_2845 (O_2845,N_29982,N_29461);
or UO_2846 (O_2846,N_29799,N_29822);
and UO_2847 (O_2847,N_29553,N_29729);
or UO_2848 (O_2848,N_29986,N_29923);
nand UO_2849 (O_2849,N_29485,N_29491);
nand UO_2850 (O_2850,N_29459,N_29809);
nand UO_2851 (O_2851,N_29468,N_29837);
nor UO_2852 (O_2852,N_29921,N_29855);
nand UO_2853 (O_2853,N_29428,N_29767);
xor UO_2854 (O_2854,N_29418,N_29844);
or UO_2855 (O_2855,N_29405,N_29653);
or UO_2856 (O_2856,N_29560,N_29961);
or UO_2857 (O_2857,N_29784,N_29741);
or UO_2858 (O_2858,N_29930,N_29859);
or UO_2859 (O_2859,N_29516,N_29651);
or UO_2860 (O_2860,N_29569,N_29831);
and UO_2861 (O_2861,N_29925,N_29626);
nand UO_2862 (O_2862,N_29677,N_29688);
nand UO_2863 (O_2863,N_29770,N_29611);
nor UO_2864 (O_2864,N_29826,N_29507);
or UO_2865 (O_2865,N_29680,N_29981);
nand UO_2866 (O_2866,N_29964,N_29999);
nand UO_2867 (O_2867,N_29534,N_29842);
and UO_2868 (O_2868,N_29826,N_29730);
xnor UO_2869 (O_2869,N_29854,N_29894);
nor UO_2870 (O_2870,N_29646,N_29724);
and UO_2871 (O_2871,N_29986,N_29989);
and UO_2872 (O_2872,N_29991,N_29609);
xor UO_2873 (O_2873,N_29485,N_29775);
xnor UO_2874 (O_2874,N_29797,N_29602);
and UO_2875 (O_2875,N_29901,N_29813);
nor UO_2876 (O_2876,N_29566,N_29575);
or UO_2877 (O_2877,N_29808,N_29792);
xor UO_2878 (O_2878,N_29840,N_29870);
nand UO_2879 (O_2879,N_29452,N_29887);
or UO_2880 (O_2880,N_29718,N_29480);
nand UO_2881 (O_2881,N_29882,N_29898);
and UO_2882 (O_2882,N_29928,N_29437);
or UO_2883 (O_2883,N_29588,N_29955);
nand UO_2884 (O_2884,N_29544,N_29743);
xor UO_2885 (O_2885,N_29757,N_29658);
nor UO_2886 (O_2886,N_29691,N_29604);
or UO_2887 (O_2887,N_29763,N_29934);
or UO_2888 (O_2888,N_29638,N_29806);
xnor UO_2889 (O_2889,N_29747,N_29749);
xnor UO_2890 (O_2890,N_29771,N_29407);
or UO_2891 (O_2891,N_29455,N_29662);
nand UO_2892 (O_2892,N_29801,N_29457);
xor UO_2893 (O_2893,N_29791,N_29777);
xnor UO_2894 (O_2894,N_29991,N_29642);
nor UO_2895 (O_2895,N_29607,N_29963);
and UO_2896 (O_2896,N_29770,N_29676);
xnor UO_2897 (O_2897,N_29755,N_29541);
nor UO_2898 (O_2898,N_29919,N_29941);
and UO_2899 (O_2899,N_29736,N_29453);
or UO_2900 (O_2900,N_29759,N_29966);
or UO_2901 (O_2901,N_29923,N_29856);
xor UO_2902 (O_2902,N_29500,N_29529);
and UO_2903 (O_2903,N_29659,N_29914);
and UO_2904 (O_2904,N_29538,N_29846);
xnor UO_2905 (O_2905,N_29537,N_29928);
or UO_2906 (O_2906,N_29411,N_29901);
and UO_2907 (O_2907,N_29804,N_29719);
nor UO_2908 (O_2908,N_29595,N_29475);
and UO_2909 (O_2909,N_29868,N_29785);
xor UO_2910 (O_2910,N_29455,N_29636);
xnor UO_2911 (O_2911,N_29729,N_29848);
and UO_2912 (O_2912,N_29911,N_29410);
or UO_2913 (O_2913,N_29489,N_29756);
and UO_2914 (O_2914,N_29999,N_29492);
nor UO_2915 (O_2915,N_29407,N_29536);
or UO_2916 (O_2916,N_29546,N_29652);
nand UO_2917 (O_2917,N_29606,N_29870);
and UO_2918 (O_2918,N_29824,N_29835);
or UO_2919 (O_2919,N_29504,N_29540);
or UO_2920 (O_2920,N_29503,N_29859);
nand UO_2921 (O_2921,N_29923,N_29977);
or UO_2922 (O_2922,N_29905,N_29608);
or UO_2923 (O_2923,N_29501,N_29636);
or UO_2924 (O_2924,N_29450,N_29668);
and UO_2925 (O_2925,N_29999,N_29525);
or UO_2926 (O_2926,N_29667,N_29760);
and UO_2927 (O_2927,N_29977,N_29478);
or UO_2928 (O_2928,N_29665,N_29848);
xnor UO_2929 (O_2929,N_29955,N_29495);
nor UO_2930 (O_2930,N_29625,N_29621);
xor UO_2931 (O_2931,N_29663,N_29948);
nand UO_2932 (O_2932,N_29733,N_29492);
xnor UO_2933 (O_2933,N_29553,N_29963);
or UO_2934 (O_2934,N_29620,N_29528);
nand UO_2935 (O_2935,N_29945,N_29904);
xnor UO_2936 (O_2936,N_29889,N_29704);
and UO_2937 (O_2937,N_29493,N_29695);
xor UO_2938 (O_2938,N_29421,N_29853);
nand UO_2939 (O_2939,N_29579,N_29536);
nand UO_2940 (O_2940,N_29440,N_29702);
or UO_2941 (O_2941,N_29846,N_29537);
xor UO_2942 (O_2942,N_29574,N_29441);
nor UO_2943 (O_2943,N_29470,N_29543);
nor UO_2944 (O_2944,N_29951,N_29565);
nor UO_2945 (O_2945,N_29679,N_29801);
xnor UO_2946 (O_2946,N_29538,N_29643);
nand UO_2947 (O_2947,N_29486,N_29453);
and UO_2948 (O_2948,N_29472,N_29669);
xnor UO_2949 (O_2949,N_29917,N_29628);
or UO_2950 (O_2950,N_29684,N_29882);
nand UO_2951 (O_2951,N_29434,N_29864);
nor UO_2952 (O_2952,N_29754,N_29678);
and UO_2953 (O_2953,N_29436,N_29920);
or UO_2954 (O_2954,N_29849,N_29655);
nand UO_2955 (O_2955,N_29607,N_29605);
nor UO_2956 (O_2956,N_29404,N_29821);
xor UO_2957 (O_2957,N_29980,N_29743);
nand UO_2958 (O_2958,N_29536,N_29487);
and UO_2959 (O_2959,N_29968,N_29535);
or UO_2960 (O_2960,N_29937,N_29582);
nand UO_2961 (O_2961,N_29927,N_29553);
or UO_2962 (O_2962,N_29832,N_29451);
nor UO_2963 (O_2963,N_29825,N_29984);
xor UO_2964 (O_2964,N_29846,N_29747);
and UO_2965 (O_2965,N_29703,N_29618);
nor UO_2966 (O_2966,N_29503,N_29903);
xor UO_2967 (O_2967,N_29451,N_29692);
and UO_2968 (O_2968,N_29999,N_29876);
and UO_2969 (O_2969,N_29756,N_29640);
or UO_2970 (O_2970,N_29906,N_29663);
and UO_2971 (O_2971,N_29409,N_29423);
nor UO_2972 (O_2972,N_29471,N_29835);
xor UO_2973 (O_2973,N_29462,N_29950);
xor UO_2974 (O_2974,N_29976,N_29425);
xnor UO_2975 (O_2975,N_29465,N_29944);
or UO_2976 (O_2976,N_29784,N_29560);
nor UO_2977 (O_2977,N_29957,N_29443);
or UO_2978 (O_2978,N_29443,N_29888);
xnor UO_2979 (O_2979,N_29739,N_29992);
xor UO_2980 (O_2980,N_29422,N_29914);
xor UO_2981 (O_2981,N_29872,N_29733);
xnor UO_2982 (O_2982,N_29576,N_29783);
and UO_2983 (O_2983,N_29742,N_29559);
nand UO_2984 (O_2984,N_29941,N_29819);
nand UO_2985 (O_2985,N_29618,N_29412);
and UO_2986 (O_2986,N_29969,N_29698);
nand UO_2987 (O_2987,N_29636,N_29555);
or UO_2988 (O_2988,N_29659,N_29901);
or UO_2989 (O_2989,N_29473,N_29917);
xnor UO_2990 (O_2990,N_29756,N_29859);
or UO_2991 (O_2991,N_29437,N_29870);
or UO_2992 (O_2992,N_29506,N_29544);
or UO_2993 (O_2993,N_29658,N_29495);
xor UO_2994 (O_2994,N_29713,N_29613);
and UO_2995 (O_2995,N_29937,N_29714);
and UO_2996 (O_2996,N_29829,N_29606);
xnor UO_2997 (O_2997,N_29632,N_29413);
xor UO_2998 (O_2998,N_29435,N_29547);
nor UO_2999 (O_2999,N_29929,N_29549);
nor UO_3000 (O_3000,N_29577,N_29560);
xnor UO_3001 (O_3001,N_29870,N_29653);
nand UO_3002 (O_3002,N_29461,N_29746);
and UO_3003 (O_3003,N_29721,N_29584);
nand UO_3004 (O_3004,N_29413,N_29422);
xnor UO_3005 (O_3005,N_29559,N_29618);
or UO_3006 (O_3006,N_29442,N_29480);
xor UO_3007 (O_3007,N_29500,N_29617);
or UO_3008 (O_3008,N_29710,N_29490);
nand UO_3009 (O_3009,N_29840,N_29472);
nor UO_3010 (O_3010,N_29887,N_29700);
and UO_3011 (O_3011,N_29907,N_29665);
xnor UO_3012 (O_3012,N_29518,N_29549);
or UO_3013 (O_3013,N_29891,N_29903);
nor UO_3014 (O_3014,N_29764,N_29632);
or UO_3015 (O_3015,N_29703,N_29838);
or UO_3016 (O_3016,N_29706,N_29804);
or UO_3017 (O_3017,N_29987,N_29730);
and UO_3018 (O_3018,N_29956,N_29625);
xnor UO_3019 (O_3019,N_29772,N_29787);
xnor UO_3020 (O_3020,N_29799,N_29481);
xor UO_3021 (O_3021,N_29741,N_29787);
nor UO_3022 (O_3022,N_29627,N_29800);
and UO_3023 (O_3023,N_29877,N_29481);
and UO_3024 (O_3024,N_29553,N_29614);
nand UO_3025 (O_3025,N_29812,N_29837);
nand UO_3026 (O_3026,N_29897,N_29485);
nor UO_3027 (O_3027,N_29659,N_29730);
nand UO_3028 (O_3028,N_29677,N_29492);
nand UO_3029 (O_3029,N_29789,N_29579);
nand UO_3030 (O_3030,N_29897,N_29416);
or UO_3031 (O_3031,N_29743,N_29565);
nor UO_3032 (O_3032,N_29747,N_29725);
nand UO_3033 (O_3033,N_29766,N_29495);
xor UO_3034 (O_3034,N_29906,N_29504);
nand UO_3035 (O_3035,N_29472,N_29797);
nor UO_3036 (O_3036,N_29987,N_29742);
xnor UO_3037 (O_3037,N_29548,N_29536);
xnor UO_3038 (O_3038,N_29759,N_29591);
nor UO_3039 (O_3039,N_29585,N_29559);
or UO_3040 (O_3040,N_29886,N_29439);
or UO_3041 (O_3041,N_29883,N_29915);
nor UO_3042 (O_3042,N_29522,N_29603);
nor UO_3043 (O_3043,N_29739,N_29805);
and UO_3044 (O_3044,N_29772,N_29897);
or UO_3045 (O_3045,N_29916,N_29404);
nor UO_3046 (O_3046,N_29608,N_29737);
xor UO_3047 (O_3047,N_29956,N_29900);
nor UO_3048 (O_3048,N_29999,N_29888);
or UO_3049 (O_3049,N_29711,N_29912);
or UO_3050 (O_3050,N_29762,N_29612);
nand UO_3051 (O_3051,N_29475,N_29560);
or UO_3052 (O_3052,N_29934,N_29806);
or UO_3053 (O_3053,N_29703,N_29609);
nor UO_3054 (O_3054,N_29627,N_29542);
nor UO_3055 (O_3055,N_29470,N_29532);
and UO_3056 (O_3056,N_29692,N_29577);
and UO_3057 (O_3057,N_29791,N_29998);
xnor UO_3058 (O_3058,N_29492,N_29468);
nor UO_3059 (O_3059,N_29663,N_29587);
xnor UO_3060 (O_3060,N_29598,N_29689);
and UO_3061 (O_3061,N_29709,N_29762);
or UO_3062 (O_3062,N_29866,N_29582);
and UO_3063 (O_3063,N_29633,N_29442);
nor UO_3064 (O_3064,N_29498,N_29580);
or UO_3065 (O_3065,N_29608,N_29951);
nor UO_3066 (O_3066,N_29869,N_29441);
nand UO_3067 (O_3067,N_29838,N_29414);
nand UO_3068 (O_3068,N_29942,N_29531);
and UO_3069 (O_3069,N_29840,N_29591);
and UO_3070 (O_3070,N_29761,N_29996);
or UO_3071 (O_3071,N_29552,N_29810);
xor UO_3072 (O_3072,N_29854,N_29947);
nand UO_3073 (O_3073,N_29881,N_29614);
and UO_3074 (O_3074,N_29523,N_29738);
nand UO_3075 (O_3075,N_29719,N_29541);
nor UO_3076 (O_3076,N_29626,N_29469);
nand UO_3077 (O_3077,N_29539,N_29971);
xnor UO_3078 (O_3078,N_29449,N_29653);
xnor UO_3079 (O_3079,N_29566,N_29746);
xnor UO_3080 (O_3080,N_29686,N_29908);
and UO_3081 (O_3081,N_29483,N_29631);
or UO_3082 (O_3082,N_29963,N_29455);
or UO_3083 (O_3083,N_29918,N_29466);
or UO_3084 (O_3084,N_29753,N_29940);
or UO_3085 (O_3085,N_29835,N_29814);
nand UO_3086 (O_3086,N_29856,N_29936);
xnor UO_3087 (O_3087,N_29769,N_29878);
nor UO_3088 (O_3088,N_29749,N_29976);
nor UO_3089 (O_3089,N_29618,N_29475);
and UO_3090 (O_3090,N_29537,N_29952);
xnor UO_3091 (O_3091,N_29929,N_29476);
nor UO_3092 (O_3092,N_29822,N_29727);
nor UO_3093 (O_3093,N_29591,N_29499);
nor UO_3094 (O_3094,N_29430,N_29865);
or UO_3095 (O_3095,N_29422,N_29713);
or UO_3096 (O_3096,N_29595,N_29567);
nand UO_3097 (O_3097,N_29581,N_29923);
and UO_3098 (O_3098,N_29448,N_29540);
nand UO_3099 (O_3099,N_29901,N_29424);
and UO_3100 (O_3100,N_29459,N_29951);
or UO_3101 (O_3101,N_29539,N_29535);
and UO_3102 (O_3102,N_29646,N_29887);
nand UO_3103 (O_3103,N_29867,N_29510);
nand UO_3104 (O_3104,N_29555,N_29463);
or UO_3105 (O_3105,N_29436,N_29544);
nand UO_3106 (O_3106,N_29997,N_29735);
nor UO_3107 (O_3107,N_29465,N_29828);
nor UO_3108 (O_3108,N_29516,N_29744);
nand UO_3109 (O_3109,N_29669,N_29849);
xor UO_3110 (O_3110,N_29684,N_29642);
nand UO_3111 (O_3111,N_29568,N_29639);
or UO_3112 (O_3112,N_29717,N_29855);
nor UO_3113 (O_3113,N_29896,N_29942);
nand UO_3114 (O_3114,N_29589,N_29415);
and UO_3115 (O_3115,N_29681,N_29954);
nor UO_3116 (O_3116,N_29526,N_29979);
and UO_3117 (O_3117,N_29564,N_29534);
or UO_3118 (O_3118,N_29569,N_29910);
nor UO_3119 (O_3119,N_29747,N_29706);
xor UO_3120 (O_3120,N_29941,N_29440);
nor UO_3121 (O_3121,N_29587,N_29475);
and UO_3122 (O_3122,N_29524,N_29590);
xnor UO_3123 (O_3123,N_29836,N_29646);
xor UO_3124 (O_3124,N_29725,N_29963);
and UO_3125 (O_3125,N_29609,N_29725);
nor UO_3126 (O_3126,N_29884,N_29496);
nor UO_3127 (O_3127,N_29709,N_29910);
and UO_3128 (O_3128,N_29686,N_29834);
nor UO_3129 (O_3129,N_29598,N_29690);
xor UO_3130 (O_3130,N_29760,N_29911);
and UO_3131 (O_3131,N_29794,N_29871);
or UO_3132 (O_3132,N_29729,N_29538);
and UO_3133 (O_3133,N_29736,N_29820);
xor UO_3134 (O_3134,N_29855,N_29519);
and UO_3135 (O_3135,N_29477,N_29814);
xnor UO_3136 (O_3136,N_29609,N_29486);
and UO_3137 (O_3137,N_29970,N_29797);
nor UO_3138 (O_3138,N_29758,N_29403);
or UO_3139 (O_3139,N_29648,N_29882);
nand UO_3140 (O_3140,N_29726,N_29501);
nand UO_3141 (O_3141,N_29804,N_29582);
or UO_3142 (O_3142,N_29656,N_29685);
xor UO_3143 (O_3143,N_29648,N_29922);
xnor UO_3144 (O_3144,N_29489,N_29641);
nor UO_3145 (O_3145,N_29932,N_29469);
or UO_3146 (O_3146,N_29693,N_29932);
nor UO_3147 (O_3147,N_29491,N_29973);
nand UO_3148 (O_3148,N_29600,N_29429);
xor UO_3149 (O_3149,N_29969,N_29519);
and UO_3150 (O_3150,N_29446,N_29576);
and UO_3151 (O_3151,N_29808,N_29765);
xnor UO_3152 (O_3152,N_29758,N_29900);
nor UO_3153 (O_3153,N_29660,N_29862);
xor UO_3154 (O_3154,N_29907,N_29432);
and UO_3155 (O_3155,N_29968,N_29427);
xnor UO_3156 (O_3156,N_29409,N_29969);
or UO_3157 (O_3157,N_29448,N_29670);
xnor UO_3158 (O_3158,N_29739,N_29712);
nor UO_3159 (O_3159,N_29869,N_29772);
xor UO_3160 (O_3160,N_29569,N_29538);
or UO_3161 (O_3161,N_29769,N_29435);
nor UO_3162 (O_3162,N_29709,N_29670);
or UO_3163 (O_3163,N_29842,N_29766);
nand UO_3164 (O_3164,N_29994,N_29590);
xor UO_3165 (O_3165,N_29794,N_29536);
xor UO_3166 (O_3166,N_29467,N_29560);
nand UO_3167 (O_3167,N_29745,N_29778);
nand UO_3168 (O_3168,N_29725,N_29726);
or UO_3169 (O_3169,N_29695,N_29792);
xnor UO_3170 (O_3170,N_29946,N_29836);
xnor UO_3171 (O_3171,N_29860,N_29486);
or UO_3172 (O_3172,N_29569,N_29875);
xnor UO_3173 (O_3173,N_29465,N_29893);
nand UO_3174 (O_3174,N_29762,N_29953);
and UO_3175 (O_3175,N_29715,N_29997);
xor UO_3176 (O_3176,N_29785,N_29971);
or UO_3177 (O_3177,N_29524,N_29836);
xor UO_3178 (O_3178,N_29563,N_29669);
xnor UO_3179 (O_3179,N_29588,N_29903);
nor UO_3180 (O_3180,N_29660,N_29578);
nor UO_3181 (O_3181,N_29844,N_29459);
or UO_3182 (O_3182,N_29733,N_29674);
nor UO_3183 (O_3183,N_29709,N_29472);
or UO_3184 (O_3184,N_29506,N_29977);
and UO_3185 (O_3185,N_29747,N_29667);
nor UO_3186 (O_3186,N_29966,N_29762);
nor UO_3187 (O_3187,N_29696,N_29616);
xor UO_3188 (O_3188,N_29556,N_29538);
xor UO_3189 (O_3189,N_29516,N_29969);
xor UO_3190 (O_3190,N_29470,N_29812);
nand UO_3191 (O_3191,N_29866,N_29545);
nor UO_3192 (O_3192,N_29682,N_29433);
and UO_3193 (O_3193,N_29670,N_29444);
nor UO_3194 (O_3194,N_29462,N_29538);
nand UO_3195 (O_3195,N_29897,N_29574);
nand UO_3196 (O_3196,N_29685,N_29457);
or UO_3197 (O_3197,N_29794,N_29807);
and UO_3198 (O_3198,N_29603,N_29855);
nand UO_3199 (O_3199,N_29939,N_29703);
nor UO_3200 (O_3200,N_29934,N_29528);
nor UO_3201 (O_3201,N_29529,N_29994);
or UO_3202 (O_3202,N_29965,N_29448);
or UO_3203 (O_3203,N_29740,N_29561);
nor UO_3204 (O_3204,N_29868,N_29748);
xnor UO_3205 (O_3205,N_29733,N_29846);
nand UO_3206 (O_3206,N_29843,N_29644);
nand UO_3207 (O_3207,N_29768,N_29705);
nor UO_3208 (O_3208,N_29423,N_29577);
xnor UO_3209 (O_3209,N_29848,N_29439);
xnor UO_3210 (O_3210,N_29433,N_29834);
nor UO_3211 (O_3211,N_29406,N_29754);
nor UO_3212 (O_3212,N_29638,N_29741);
nand UO_3213 (O_3213,N_29476,N_29678);
xor UO_3214 (O_3214,N_29944,N_29900);
nor UO_3215 (O_3215,N_29748,N_29769);
nor UO_3216 (O_3216,N_29983,N_29412);
nand UO_3217 (O_3217,N_29858,N_29855);
nand UO_3218 (O_3218,N_29887,N_29984);
nor UO_3219 (O_3219,N_29729,N_29616);
or UO_3220 (O_3220,N_29916,N_29726);
or UO_3221 (O_3221,N_29677,N_29653);
nand UO_3222 (O_3222,N_29550,N_29559);
and UO_3223 (O_3223,N_29853,N_29936);
xnor UO_3224 (O_3224,N_29850,N_29554);
and UO_3225 (O_3225,N_29830,N_29758);
xor UO_3226 (O_3226,N_29959,N_29406);
or UO_3227 (O_3227,N_29694,N_29597);
or UO_3228 (O_3228,N_29470,N_29946);
nand UO_3229 (O_3229,N_29949,N_29599);
and UO_3230 (O_3230,N_29832,N_29995);
nand UO_3231 (O_3231,N_29422,N_29406);
and UO_3232 (O_3232,N_29544,N_29653);
xnor UO_3233 (O_3233,N_29642,N_29614);
and UO_3234 (O_3234,N_29953,N_29607);
or UO_3235 (O_3235,N_29531,N_29922);
and UO_3236 (O_3236,N_29452,N_29501);
xnor UO_3237 (O_3237,N_29898,N_29532);
xor UO_3238 (O_3238,N_29543,N_29803);
or UO_3239 (O_3239,N_29665,N_29754);
nor UO_3240 (O_3240,N_29636,N_29488);
or UO_3241 (O_3241,N_29837,N_29911);
nor UO_3242 (O_3242,N_29955,N_29672);
and UO_3243 (O_3243,N_29594,N_29930);
or UO_3244 (O_3244,N_29700,N_29685);
and UO_3245 (O_3245,N_29448,N_29913);
xor UO_3246 (O_3246,N_29801,N_29724);
xnor UO_3247 (O_3247,N_29829,N_29866);
or UO_3248 (O_3248,N_29444,N_29528);
or UO_3249 (O_3249,N_29793,N_29966);
nor UO_3250 (O_3250,N_29666,N_29660);
nand UO_3251 (O_3251,N_29910,N_29790);
or UO_3252 (O_3252,N_29542,N_29671);
or UO_3253 (O_3253,N_29710,N_29956);
nor UO_3254 (O_3254,N_29879,N_29451);
xor UO_3255 (O_3255,N_29460,N_29992);
nor UO_3256 (O_3256,N_29695,N_29683);
and UO_3257 (O_3257,N_29542,N_29652);
nand UO_3258 (O_3258,N_29865,N_29500);
nor UO_3259 (O_3259,N_29631,N_29438);
xnor UO_3260 (O_3260,N_29863,N_29817);
nor UO_3261 (O_3261,N_29844,N_29479);
xor UO_3262 (O_3262,N_29676,N_29885);
xnor UO_3263 (O_3263,N_29538,N_29949);
nand UO_3264 (O_3264,N_29820,N_29621);
xor UO_3265 (O_3265,N_29999,N_29470);
and UO_3266 (O_3266,N_29866,N_29619);
nand UO_3267 (O_3267,N_29538,N_29810);
nand UO_3268 (O_3268,N_29935,N_29794);
xnor UO_3269 (O_3269,N_29446,N_29657);
and UO_3270 (O_3270,N_29651,N_29928);
xor UO_3271 (O_3271,N_29404,N_29533);
or UO_3272 (O_3272,N_29632,N_29636);
or UO_3273 (O_3273,N_29509,N_29454);
xor UO_3274 (O_3274,N_29697,N_29817);
or UO_3275 (O_3275,N_29530,N_29535);
nor UO_3276 (O_3276,N_29923,N_29809);
nand UO_3277 (O_3277,N_29850,N_29447);
xnor UO_3278 (O_3278,N_29436,N_29647);
or UO_3279 (O_3279,N_29708,N_29664);
xnor UO_3280 (O_3280,N_29710,N_29728);
xor UO_3281 (O_3281,N_29757,N_29578);
nand UO_3282 (O_3282,N_29619,N_29984);
nand UO_3283 (O_3283,N_29690,N_29846);
and UO_3284 (O_3284,N_29780,N_29998);
and UO_3285 (O_3285,N_29794,N_29680);
and UO_3286 (O_3286,N_29507,N_29779);
nor UO_3287 (O_3287,N_29618,N_29925);
nand UO_3288 (O_3288,N_29845,N_29685);
xor UO_3289 (O_3289,N_29488,N_29439);
nand UO_3290 (O_3290,N_29735,N_29538);
or UO_3291 (O_3291,N_29749,N_29524);
nand UO_3292 (O_3292,N_29567,N_29944);
or UO_3293 (O_3293,N_29704,N_29805);
and UO_3294 (O_3294,N_29432,N_29830);
xor UO_3295 (O_3295,N_29608,N_29581);
nand UO_3296 (O_3296,N_29749,N_29628);
xnor UO_3297 (O_3297,N_29715,N_29854);
or UO_3298 (O_3298,N_29448,N_29816);
nand UO_3299 (O_3299,N_29786,N_29619);
xor UO_3300 (O_3300,N_29967,N_29500);
xor UO_3301 (O_3301,N_29500,N_29585);
nor UO_3302 (O_3302,N_29566,N_29616);
nand UO_3303 (O_3303,N_29536,N_29675);
or UO_3304 (O_3304,N_29687,N_29712);
and UO_3305 (O_3305,N_29427,N_29756);
nand UO_3306 (O_3306,N_29705,N_29861);
and UO_3307 (O_3307,N_29404,N_29656);
xor UO_3308 (O_3308,N_29421,N_29642);
nand UO_3309 (O_3309,N_29707,N_29629);
nand UO_3310 (O_3310,N_29868,N_29691);
nor UO_3311 (O_3311,N_29611,N_29426);
and UO_3312 (O_3312,N_29925,N_29468);
and UO_3313 (O_3313,N_29560,N_29406);
or UO_3314 (O_3314,N_29891,N_29930);
xor UO_3315 (O_3315,N_29587,N_29588);
or UO_3316 (O_3316,N_29545,N_29773);
or UO_3317 (O_3317,N_29618,N_29605);
and UO_3318 (O_3318,N_29905,N_29702);
xor UO_3319 (O_3319,N_29750,N_29711);
nand UO_3320 (O_3320,N_29843,N_29600);
xor UO_3321 (O_3321,N_29484,N_29849);
and UO_3322 (O_3322,N_29508,N_29549);
nand UO_3323 (O_3323,N_29483,N_29956);
nand UO_3324 (O_3324,N_29656,N_29629);
xor UO_3325 (O_3325,N_29798,N_29463);
or UO_3326 (O_3326,N_29461,N_29506);
and UO_3327 (O_3327,N_29889,N_29941);
and UO_3328 (O_3328,N_29506,N_29856);
nor UO_3329 (O_3329,N_29521,N_29420);
and UO_3330 (O_3330,N_29849,N_29825);
or UO_3331 (O_3331,N_29682,N_29739);
nor UO_3332 (O_3332,N_29916,N_29427);
and UO_3333 (O_3333,N_29484,N_29860);
xor UO_3334 (O_3334,N_29594,N_29861);
or UO_3335 (O_3335,N_29750,N_29767);
and UO_3336 (O_3336,N_29460,N_29830);
and UO_3337 (O_3337,N_29844,N_29448);
or UO_3338 (O_3338,N_29818,N_29873);
nor UO_3339 (O_3339,N_29738,N_29967);
and UO_3340 (O_3340,N_29881,N_29455);
xor UO_3341 (O_3341,N_29539,N_29633);
and UO_3342 (O_3342,N_29804,N_29453);
and UO_3343 (O_3343,N_29828,N_29993);
or UO_3344 (O_3344,N_29974,N_29665);
nor UO_3345 (O_3345,N_29746,N_29873);
nand UO_3346 (O_3346,N_29681,N_29773);
nand UO_3347 (O_3347,N_29462,N_29835);
or UO_3348 (O_3348,N_29895,N_29974);
or UO_3349 (O_3349,N_29743,N_29729);
and UO_3350 (O_3350,N_29572,N_29883);
xor UO_3351 (O_3351,N_29535,N_29665);
nor UO_3352 (O_3352,N_29545,N_29490);
xor UO_3353 (O_3353,N_29448,N_29958);
or UO_3354 (O_3354,N_29934,N_29715);
or UO_3355 (O_3355,N_29500,N_29492);
and UO_3356 (O_3356,N_29649,N_29514);
nand UO_3357 (O_3357,N_29401,N_29713);
xnor UO_3358 (O_3358,N_29590,N_29834);
and UO_3359 (O_3359,N_29411,N_29581);
nand UO_3360 (O_3360,N_29825,N_29745);
xnor UO_3361 (O_3361,N_29888,N_29726);
or UO_3362 (O_3362,N_29426,N_29472);
nor UO_3363 (O_3363,N_29933,N_29684);
or UO_3364 (O_3364,N_29886,N_29858);
or UO_3365 (O_3365,N_29658,N_29736);
or UO_3366 (O_3366,N_29701,N_29418);
nor UO_3367 (O_3367,N_29484,N_29644);
nor UO_3368 (O_3368,N_29903,N_29775);
or UO_3369 (O_3369,N_29409,N_29530);
nor UO_3370 (O_3370,N_29540,N_29800);
or UO_3371 (O_3371,N_29812,N_29562);
or UO_3372 (O_3372,N_29858,N_29889);
and UO_3373 (O_3373,N_29935,N_29693);
xor UO_3374 (O_3374,N_29840,N_29641);
nand UO_3375 (O_3375,N_29925,N_29858);
nor UO_3376 (O_3376,N_29464,N_29635);
nor UO_3377 (O_3377,N_29952,N_29529);
and UO_3378 (O_3378,N_29988,N_29883);
nor UO_3379 (O_3379,N_29626,N_29920);
nand UO_3380 (O_3380,N_29419,N_29889);
nand UO_3381 (O_3381,N_29704,N_29431);
nor UO_3382 (O_3382,N_29722,N_29940);
nor UO_3383 (O_3383,N_29586,N_29957);
nor UO_3384 (O_3384,N_29973,N_29918);
and UO_3385 (O_3385,N_29851,N_29602);
nand UO_3386 (O_3386,N_29709,N_29610);
nand UO_3387 (O_3387,N_29678,N_29848);
xnor UO_3388 (O_3388,N_29825,N_29772);
and UO_3389 (O_3389,N_29763,N_29654);
nand UO_3390 (O_3390,N_29459,N_29636);
nor UO_3391 (O_3391,N_29944,N_29503);
nand UO_3392 (O_3392,N_29573,N_29858);
nor UO_3393 (O_3393,N_29873,N_29543);
nand UO_3394 (O_3394,N_29777,N_29953);
nor UO_3395 (O_3395,N_29916,N_29969);
xnor UO_3396 (O_3396,N_29921,N_29909);
and UO_3397 (O_3397,N_29661,N_29770);
nand UO_3398 (O_3398,N_29404,N_29702);
xnor UO_3399 (O_3399,N_29687,N_29702);
and UO_3400 (O_3400,N_29468,N_29463);
nand UO_3401 (O_3401,N_29562,N_29754);
or UO_3402 (O_3402,N_29624,N_29625);
and UO_3403 (O_3403,N_29690,N_29573);
xnor UO_3404 (O_3404,N_29479,N_29643);
nand UO_3405 (O_3405,N_29966,N_29810);
nand UO_3406 (O_3406,N_29792,N_29618);
or UO_3407 (O_3407,N_29999,N_29625);
nand UO_3408 (O_3408,N_29984,N_29976);
xor UO_3409 (O_3409,N_29734,N_29705);
or UO_3410 (O_3410,N_29698,N_29768);
nor UO_3411 (O_3411,N_29563,N_29919);
or UO_3412 (O_3412,N_29434,N_29931);
xnor UO_3413 (O_3413,N_29613,N_29605);
xor UO_3414 (O_3414,N_29410,N_29583);
or UO_3415 (O_3415,N_29642,N_29502);
nand UO_3416 (O_3416,N_29543,N_29556);
and UO_3417 (O_3417,N_29858,N_29893);
and UO_3418 (O_3418,N_29688,N_29407);
xor UO_3419 (O_3419,N_29934,N_29623);
and UO_3420 (O_3420,N_29407,N_29804);
xor UO_3421 (O_3421,N_29900,N_29542);
nor UO_3422 (O_3422,N_29954,N_29585);
nor UO_3423 (O_3423,N_29645,N_29878);
or UO_3424 (O_3424,N_29517,N_29773);
and UO_3425 (O_3425,N_29750,N_29564);
xor UO_3426 (O_3426,N_29768,N_29931);
xor UO_3427 (O_3427,N_29542,N_29670);
nor UO_3428 (O_3428,N_29759,N_29661);
nand UO_3429 (O_3429,N_29520,N_29653);
nor UO_3430 (O_3430,N_29709,N_29497);
nor UO_3431 (O_3431,N_29743,N_29482);
and UO_3432 (O_3432,N_29631,N_29730);
and UO_3433 (O_3433,N_29748,N_29976);
and UO_3434 (O_3434,N_29795,N_29465);
nand UO_3435 (O_3435,N_29824,N_29967);
and UO_3436 (O_3436,N_29878,N_29481);
and UO_3437 (O_3437,N_29807,N_29684);
and UO_3438 (O_3438,N_29723,N_29605);
nand UO_3439 (O_3439,N_29783,N_29953);
nand UO_3440 (O_3440,N_29917,N_29829);
or UO_3441 (O_3441,N_29766,N_29993);
nand UO_3442 (O_3442,N_29627,N_29556);
nand UO_3443 (O_3443,N_29698,N_29840);
xor UO_3444 (O_3444,N_29563,N_29532);
or UO_3445 (O_3445,N_29455,N_29957);
and UO_3446 (O_3446,N_29952,N_29527);
and UO_3447 (O_3447,N_29624,N_29858);
nand UO_3448 (O_3448,N_29651,N_29403);
and UO_3449 (O_3449,N_29502,N_29538);
and UO_3450 (O_3450,N_29712,N_29816);
nand UO_3451 (O_3451,N_29717,N_29617);
nor UO_3452 (O_3452,N_29588,N_29884);
nor UO_3453 (O_3453,N_29675,N_29870);
and UO_3454 (O_3454,N_29470,N_29711);
nor UO_3455 (O_3455,N_29562,N_29793);
nor UO_3456 (O_3456,N_29800,N_29714);
nand UO_3457 (O_3457,N_29516,N_29818);
nor UO_3458 (O_3458,N_29806,N_29492);
nand UO_3459 (O_3459,N_29743,N_29929);
xnor UO_3460 (O_3460,N_29404,N_29880);
or UO_3461 (O_3461,N_29917,N_29443);
nor UO_3462 (O_3462,N_29662,N_29706);
nor UO_3463 (O_3463,N_29526,N_29436);
or UO_3464 (O_3464,N_29889,N_29671);
and UO_3465 (O_3465,N_29878,N_29430);
nand UO_3466 (O_3466,N_29761,N_29523);
nor UO_3467 (O_3467,N_29573,N_29867);
and UO_3468 (O_3468,N_29706,N_29485);
nand UO_3469 (O_3469,N_29778,N_29502);
nand UO_3470 (O_3470,N_29611,N_29860);
xnor UO_3471 (O_3471,N_29971,N_29915);
and UO_3472 (O_3472,N_29410,N_29810);
nand UO_3473 (O_3473,N_29791,N_29502);
and UO_3474 (O_3474,N_29991,N_29864);
or UO_3475 (O_3475,N_29589,N_29985);
and UO_3476 (O_3476,N_29537,N_29910);
and UO_3477 (O_3477,N_29754,N_29569);
nand UO_3478 (O_3478,N_29668,N_29710);
nand UO_3479 (O_3479,N_29750,N_29846);
xor UO_3480 (O_3480,N_29505,N_29456);
xnor UO_3481 (O_3481,N_29920,N_29531);
nor UO_3482 (O_3482,N_29594,N_29791);
nor UO_3483 (O_3483,N_29738,N_29994);
and UO_3484 (O_3484,N_29785,N_29590);
nand UO_3485 (O_3485,N_29882,N_29916);
nor UO_3486 (O_3486,N_29656,N_29626);
or UO_3487 (O_3487,N_29770,N_29537);
or UO_3488 (O_3488,N_29988,N_29939);
nor UO_3489 (O_3489,N_29580,N_29463);
xnor UO_3490 (O_3490,N_29717,N_29826);
and UO_3491 (O_3491,N_29729,N_29801);
or UO_3492 (O_3492,N_29779,N_29407);
xnor UO_3493 (O_3493,N_29466,N_29880);
nand UO_3494 (O_3494,N_29607,N_29722);
nand UO_3495 (O_3495,N_29966,N_29637);
nand UO_3496 (O_3496,N_29716,N_29729);
nor UO_3497 (O_3497,N_29905,N_29625);
and UO_3498 (O_3498,N_29674,N_29793);
and UO_3499 (O_3499,N_29784,N_29934);
endmodule